module basic_2500_25000_3000_10_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_767,In_625);
nor U1 (N_1,In_872,In_680);
and U2 (N_2,In_180,In_27);
nand U3 (N_3,In_1840,In_2440);
nand U4 (N_4,In_2297,In_945);
nand U5 (N_5,In_2024,In_2030);
nand U6 (N_6,In_371,In_1105);
and U7 (N_7,In_2266,In_276);
or U8 (N_8,In_1759,In_1790);
or U9 (N_9,In_2122,In_666);
and U10 (N_10,In_85,In_1011);
nand U11 (N_11,In_498,In_636);
or U12 (N_12,In_1073,In_275);
nand U13 (N_13,In_1742,In_120);
or U14 (N_14,In_2354,In_1543);
and U15 (N_15,In_173,In_1128);
nand U16 (N_16,In_259,In_379);
or U17 (N_17,In_2281,In_964);
or U18 (N_18,In_1715,In_2326);
nor U19 (N_19,In_1679,In_393);
nand U20 (N_20,In_732,In_1692);
and U21 (N_21,In_1556,In_1960);
or U22 (N_22,In_1406,In_1347);
or U23 (N_23,In_1839,In_1313);
nand U24 (N_24,In_1366,In_594);
nor U25 (N_25,In_2260,In_1405);
nor U26 (N_26,In_410,In_423);
nand U27 (N_27,In_2275,In_1417);
and U28 (N_28,In_1953,In_1254);
or U29 (N_29,In_854,In_144);
or U30 (N_30,In_2080,In_1411);
nor U31 (N_31,In_1546,In_2119);
or U32 (N_32,In_165,In_207);
or U33 (N_33,In_1090,In_1232);
nor U34 (N_34,In_1442,In_1928);
nor U35 (N_35,In_1272,In_2114);
and U36 (N_36,In_2120,In_1233);
nand U37 (N_37,In_1104,In_642);
nand U38 (N_38,In_2382,In_2203);
nand U39 (N_39,In_2320,In_1358);
or U40 (N_40,In_1631,In_282);
or U41 (N_41,In_2201,In_2363);
or U42 (N_42,In_1798,In_279);
nor U43 (N_43,In_364,In_557);
nand U44 (N_44,In_2476,In_2091);
nand U45 (N_45,In_1460,In_995);
nand U46 (N_46,In_373,In_991);
and U47 (N_47,In_527,In_2288);
nor U48 (N_48,In_653,In_109);
nor U49 (N_49,In_1147,In_1842);
xor U50 (N_50,In_1564,In_1588);
nand U51 (N_51,In_89,In_792);
nand U52 (N_52,In_1414,In_2093);
or U53 (N_53,In_2362,In_2443);
nand U54 (N_54,In_1628,In_696);
and U55 (N_55,In_997,In_1419);
nand U56 (N_56,In_358,In_419);
or U57 (N_57,In_1671,In_2498);
nand U58 (N_58,In_2347,In_936);
nand U59 (N_59,In_2360,In_29);
nor U60 (N_60,In_1736,In_1365);
or U61 (N_61,In_359,In_1046);
nor U62 (N_62,In_895,In_2349);
nor U63 (N_63,In_645,In_130);
nand U64 (N_64,In_1424,In_168);
nor U65 (N_65,In_1107,In_510);
nor U66 (N_66,In_682,In_1784);
and U67 (N_67,In_707,In_2283);
and U68 (N_68,In_1506,In_2046);
nand U69 (N_69,In_1923,In_1894);
or U70 (N_70,In_1727,In_1970);
nand U71 (N_71,In_2238,In_1587);
and U72 (N_72,In_1827,In_1328);
nor U73 (N_73,In_980,In_274);
or U74 (N_74,In_2135,In_690);
or U75 (N_75,In_939,In_1093);
nor U76 (N_76,In_783,In_1271);
and U77 (N_77,In_1648,In_82);
nor U78 (N_78,In_129,In_2265);
and U79 (N_79,In_1226,In_491);
nand U80 (N_80,In_1268,In_2366);
and U81 (N_81,In_710,In_1244);
nand U82 (N_82,In_2333,In_2337);
nor U83 (N_83,In_1101,In_2167);
nor U84 (N_84,In_1067,In_1998);
nand U85 (N_85,In_1608,In_236);
nor U86 (N_86,In_2469,In_1126);
or U87 (N_87,In_2481,In_1463);
and U88 (N_88,In_1984,In_2494);
nand U89 (N_89,In_1224,In_64);
nor U90 (N_90,In_385,In_102);
or U91 (N_91,In_838,In_1377);
nor U92 (N_92,In_1934,In_238);
nand U93 (N_93,In_1799,In_2392);
or U94 (N_94,In_189,In_1973);
nor U95 (N_95,In_533,In_2218);
nand U96 (N_96,In_867,In_1797);
or U97 (N_97,In_965,In_979);
or U98 (N_98,In_2401,In_197);
and U99 (N_99,In_2132,In_567);
and U100 (N_100,In_1513,In_992);
and U101 (N_101,In_839,In_1555);
or U102 (N_102,In_1156,In_1431);
nand U103 (N_103,In_656,In_2215);
and U104 (N_104,In_1976,In_1999);
or U105 (N_105,In_996,In_1844);
and U106 (N_106,In_1082,In_2426);
nand U107 (N_107,In_813,In_1075);
and U108 (N_108,In_1275,In_2035);
nor U109 (N_109,In_2403,In_678);
or U110 (N_110,In_1372,In_1416);
nor U111 (N_111,In_249,In_1178);
nand U112 (N_112,In_2313,In_1114);
nand U113 (N_113,In_1155,In_1214);
and U114 (N_114,In_2386,In_815);
xnor U115 (N_115,In_488,In_758);
or U116 (N_116,In_472,In_2451);
nand U117 (N_117,In_906,In_864);
and U118 (N_118,In_1944,In_2131);
and U119 (N_119,In_460,In_232);
or U120 (N_120,In_225,In_622);
or U121 (N_121,In_1758,In_1367);
or U122 (N_122,In_1192,In_341);
nor U123 (N_123,In_2027,In_855);
and U124 (N_124,In_1814,In_1488);
nor U125 (N_125,In_2126,In_1451);
nand U126 (N_126,In_1712,In_1522);
nor U127 (N_127,In_2061,In_1884);
xor U128 (N_128,In_51,In_1455);
or U129 (N_129,In_729,In_2213);
nor U130 (N_130,In_632,In_1108);
nand U131 (N_131,In_1489,In_2009);
nand U132 (N_132,In_988,In_188);
nor U133 (N_133,In_1326,In_2235);
nand U134 (N_134,In_1318,In_427);
or U135 (N_135,In_1332,In_2474);
or U136 (N_136,In_1935,In_628);
nor U137 (N_137,In_1693,In_493);
nand U138 (N_138,In_1145,In_2322);
and U139 (N_139,In_426,In_1299);
nand U140 (N_140,In_94,In_1913);
nor U141 (N_141,In_1403,In_1824);
or U142 (N_142,In_35,In_791);
nor U143 (N_143,In_1535,In_908);
and U144 (N_144,In_1660,In_564);
or U145 (N_145,In_1512,In_2277);
nor U146 (N_146,In_730,In_301);
nand U147 (N_147,In_1948,In_552);
nand U148 (N_148,In_148,In_289);
nand U149 (N_149,In_689,In_1203);
nor U150 (N_150,In_288,In_568);
or U151 (N_151,In_1070,In_1245);
xnor U152 (N_152,In_607,In_747);
or U153 (N_153,In_612,In_1330);
and U154 (N_154,In_389,In_749);
nor U155 (N_155,In_1753,In_1634);
and U156 (N_156,In_194,In_829);
and U157 (N_157,In_386,In_4);
nor U158 (N_158,In_1293,In_571);
nand U159 (N_159,In_2019,In_1949);
nand U160 (N_160,In_1127,In_1282);
nand U161 (N_161,In_1346,In_950);
or U162 (N_162,In_2318,In_1468);
or U163 (N_163,In_3,In_11);
nand U164 (N_164,In_2471,In_2129);
nand U165 (N_165,In_2000,In_2196);
nor U166 (N_166,In_1558,In_2043);
nor U167 (N_167,In_1576,In_2107);
nor U168 (N_168,In_775,In_1164);
nand U169 (N_169,In_2197,In_47);
nor U170 (N_170,In_1118,In_1172);
or U171 (N_171,In_596,In_2279);
or U172 (N_172,In_699,In_366);
nor U173 (N_173,In_1012,In_1670);
nor U174 (N_174,In_1335,In_1925);
nand U175 (N_175,In_750,In_1601);
and U176 (N_176,In_2017,In_1922);
nand U177 (N_177,In_2383,In_86);
and U178 (N_178,In_993,In_2368);
and U179 (N_179,In_1499,In_530);
or U180 (N_180,In_849,In_489);
and U181 (N_181,In_526,In_1698);
nor U182 (N_182,In_576,In_1765);
nor U183 (N_183,In_1937,In_941);
nor U184 (N_184,In_1287,In_1109);
or U185 (N_185,In_952,In_445);
or U186 (N_186,In_2087,In_181);
or U187 (N_187,In_743,In_1874);
and U188 (N_188,In_81,In_91);
or U189 (N_189,In_1135,In_528);
xnor U190 (N_190,In_1462,In_496);
and U191 (N_191,In_1408,In_442);
and U192 (N_192,In_2071,In_659);
nor U193 (N_193,In_2488,In_2435);
nor U194 (N_194,In_2141,In_1866);
and U195 (N_195,In_1062,In_212);
nand U196 (N_196,In_2356,In_1154);
nand U197 (N_197,In_1015,In_416);
and U198 (N_198,In_2078,In_208);
nor U199 (N_199,In_1452,In_1096);
xnor U200 (N_200,In_810,In_331);
and U201 (N_201,In_2136,In_322);
or U202 (N_202,In_725,In_1484);
and U203 (N_203,In_164,In_2490);
nor U204 (N_204,In_638,In_591);
or U205 (N_205,In_721,In_344);
and U206 (N_206,In_1017,In_2444);
and U207 (N_207,In_2365,In_1688);
nor U208 (N_208,In_1672,In_819);
nor U209 (N_209,In_1741,In_874);
and U210 (N_210,In_615,In_1606);
and U211 (N_211,In_1028,In_1051);
nand U212 (N_212,In_1746,In_1324);
nor U213 (N_213,In_1166,In_1722);
and U214 (N_214,In_1952,In_1032);
nand U215 (N_215,In_2355,In_2237);
and U216 (N_216,In_1965,In_2121);
nand U217 (N_217,In_1355,In_1354);
or U218 (N_218,In_1927,In_2202);
and U219 (N_219,In_1781,In_2045);
and U220 (N_220,In_869,In_1078);
nand U221 (N_221,In_948,In_1153);
or U222 (N_222,In_2467,In_1767);
or U223 (N_223,In_1151,In_337);
and U224 (N_224,In_1225,In_161);
and U225 (N_225,In_2003,In_1450);
or U226 (N_226,In_79,In_114);
nand U227 (N_227,In_1482,In_318);
and U228 (N_228,In_132,In_842);
nor U229 (N_229,In_695,In_953);
nor U230 (N_230,In_56,In_420);
and U231 (N_231,In_2343,In_676);
nand U232 (N_232,In_2060,In_408);
nor U233 (N_233,In_1505,In_283);
or U234 (N_234,In_1989,In_298);
nor U235 (N_235,In_692,In_740);
or U236 (N_236,In_1921,In_2329);
nand U237 (N_237,In_1918,In_1885);
nand U238 (N_238,In_1149,In_1880);
nor U239 (N_239,In_1071,In_1896);
nand U240 (N_240,In_326,In_1349);
and U241 (N_241,In_1407,In_1764);
and U242 (N_242,In_1751,In_314);
or U243 (N_243,In_1184,In_1750);
nand U244 (N_244,In_2190,In_1124);
or U245 (N_245,In_932,In_159);
or U246 (N_246,In_2258,In_2262);
or U247 (N_247,In_346,In_1723);
nand U248 (N_248,In_1074,In_820);
or U249 (N_249,In_2424,In_1585);
nor U250 (N_250,In_1507,In_1562);
and U251 (N_251,In_2187,In_1158);
nand U252 (N_252,In_16,In_943);
nand U253 (N_253,In_1009,In_1402);
or U254 (N_254,In_973,In_2259);
or U255 (N_255,In_316,In_1503);
and U256 (N_256,In_1357,In_1069);
or U257 (N_257,In_1130,In_2004);
nor U258 (N_258,In_2461,In_1709);
or U259 (N_259,In_800,In_1390);
or U260 (N_260,In_816,In_608);
and U261 (N_261,In_1899,In_975);
and U262 (N_262,In_2397,In_2147);
or U263 (N_263,In_0,In_1316);
nand U264 (N_264,In_403,In_2088);
xor U265 (N_265,In_994,In_1384);
nand U266 (N_266,In_2475,In_2282);
nand U267 (N_267,In_2040,In_1851);
and U268 (N_268,In_2064,In_1681);
nor U269 (N_269,In_938,In_2252);
nor U270 (N_270,In_866,In_34);
and U271 (N_271,In_265,In_580);
nand U272 (N_272,In_1199,In_1175);
or U273 (N_273,In_2072,In_2056);
nor U274 (N_274,In_978,In_1168);
nand U275 (N_275,In_1963,In_1539);
and U276 (N_276,In_1187,In_1337);
nand U277 (N_277,In_773,In_2089);
and U278 (N_278,In_2303,In_1530);
xor U279 (N_279,In_2206,In_913);
or U280 (N_280,In_417,In_2211);
nor U281 (N_281,In_387,In_762);
and U282 (N_282,In_1286,In_1196);
nand U283 (N_283,In_80,In_1491);
nand U284 (N_284,In_1834,In_2497);
nand U285 (N_285,In_59,In_837);
or U286 (N_286,In_158,In_302);
and U287 (N_287,In_2034,In_798);
nor U288 (N_288,In_1205,In_2348);
nor U289 (N_289,In_2033,In_790);
or U290 (N_290,In_1964,In_1435);
or U291 (N_291,In_2094,In_2150);
nor U292 (N_292,In_492,In_1718);
xnor U293 (N_293,In_579,In_2044);
and U294 (N_294,In_2344,In_1152);
and U295 (N_295,In_904,In_990);
and U296 (N_296,In_616,In_769);
nor U297 (N_297,In_186,In_1911);
nor U298 (N_298,In_446,In_1210);
nand U299 (N_299,In_777,In_39);
and U300 (N_300,In_443,In_2325);
nor U301 (N_301,In_354,In_903);
nor U302 (N_302,In_565,In_119);
and U303 (N_303,In_1375,In_1296);
or U304 (N_304,In_1230,In_2410);
and U305 (N_305,In_1443,In_1983);
and U306 (N_306,In_1622,In_362);
and U307 (N_307,In_1023,In_143);
nor U308 (N_308,In_1289,In_1768);
nor U309 (N_309,In_1000,In_2458);
and U310 (N_310,In_2417,In_586);
or U311 (N_311,In_629,In_698);
nor U312 (N_312,In_1242,In_2395);
nor U313 (N_313,In_428,In_940);
and U314 (N_314,In_2178,In_1720);
and U315 (N_315,In_2070,In_327);
nor U316 (N_316,In_2143,In_930);
nand U317 (N_317,In_1321,In_296);
and U318 (N_318,In_1083,In_834);
and U319 (N_319,In_1818,In_2371);
nand U320 (N_320,In_541,In_87);
nand U321 (N_321,In_2384,In_2012);
nand U322 (N_322,In_483,In_1053);
nand U323 (N_323,In_520,In_2117);
and U324 (N_324,In_424,In_1967);
or U325 (N_325,In_824,In_734);
nor U326 (N_326,In_10,In_2406);
or U327 (N_327,In_2229,In_2242);
nand U328 (N_328,In_1122,In_641);
nor U329 (N_329,In_2264,In_280);
nor U330 (N_330,In_1620,In_947);
or U331 (N_331,In_1027,In_556);
and U332 (N_332,In_270,In_2307);
and U333 (N_333,In_1030,In_1426);
nand U334 (N_334,In_1700,In_706);
or U335 (N_335,In_860,In_2057);
and U336 (N_336,In_95,In_83);
nand U337 (N_337,In_240,In_2128);
or U338 (N_338,In_1730,In_634);
or U339 (N_339,In_1778,In_1902);
and U340 (N_340,In_1255,In_2418);
or U341 (N_341,In_286,In_1529);
or U342 (N_342,In_1234,In_2407);
nand U343 (N_343,In_343,In_210);
nor U344 (N_344,In_1541,In_848);
or U345 (N_345,In_630,In_668);
or U346 (N_346,In_342,In_1301);
and U347 (N_347,In_717,In_1959);
xnor U348 (N_348,In_673,In_871);
and U349 (N_349,In_1094,In_779);
and U350 (N_350,In_720,In_1095);
nor U351 (N_351,In_2416,In_142);
and U352 (N_352,In_9,In_1803);
nor U353 (N_353,In_1991,In_2250);
nor U354 (N_354,In_703,In_1705);
nand U355 (N_355,In_1914,In_2367);
or U356 (N_356,In_141,In_48);
nand U357 (N_357,In_910,In_2387);
nand U358 (N_358,In_501,In_1534);
and U359 (N_359,In_1183,In_1055);
or U360 (N_360,In_1855,In_2209);
nor U361 (N_361,In_1815,In_1992);
nand U362 (N_362,In_218,In_170);
nor U363 (N_363,In_1605,In_1081);
or U364 (N_364,In_1072,In_1089);
or U365 (N_365,In_1604,In_2184);
nor U366 (N_366,In_479,In_2075);
nor U367 (N_367,In_701,In_922);
nor U368 (N_368,In_1662,In_759);
and U369 (N_369,In_2018,In_1769);
nand U370 (N_370,In_2021,In_2241);
nand U371 (N_371,In_1573,In_1550);
or U372 (N_372,In_1551,In_1932);
nor U373 (N_373,In_60,In_620);
xor U374 (N_374,In_1630,In_1439);
and U375 (N_375,In_1941,In_1651);
nor U376 (N_376,In_1602,In_889);
nor U377 (N_377,In_1415,In_78);
nand U378 (N_378,In_217,In_1859);
or U379 (N_379,In_1962,In_2472);
nand U380 (N_380,In_1434,In_1441);
xor U381 (N_381,In_2134,In_481);
nand U382 (N_382,In_1413,In_1777);
nand U383 (N_383,In_1058,In_1554);
nand U384 (N_384,In_900,In_2321);
nor U385 (N_385,In_2449,In_1616);
nor U386 (N_386,In_2376,In_516);
and U387 (N_387,In_915,In_1305);
nand U388 (N_388,In_2463,In_2351);
nand U389 (N_389,In_99,In_672);
and U390 (N_390,In_1352,In_2152);
and U391 (N_391,In_1956,In_2224);
and U392 (N_392,In_1676,In_951);
and U393 (N_393,In_431,In_989);
or U394 (N_394,In_55,In_1873);
nor U395 (N_395,In_2011,In_394);
nor U396 (N_396,In_2293,In_2358);
nand U397 (N_397,In_1170,In_1760);
nor U398 (N_398,In_2331,In_439);
nor U399 (N_399,In_914,In_18);
nor U400 (N_400,In_20,In_687);
nand U401 (N_401,In_738,In_755);
nor U402 (N_402,In_1930,In_2272);
nor U403 (N_403,In_1290,In_765);
or U404 (N_404,In_495,In_970);
or U405 (N_405,In_2340,In_23);
nand U406 (N_406,In_2050,In_826);
nor U407 (N_407,In_2186,In_1303);
or U408 (N_408,In_1888,In_1878);
nand U409 (N_409,In_1780,In_1821);
and U410 (N_410,In_681,In_1785);
nand U411 (N_411,In_511,In_31);
or U412 (N_412,In_2442,In_1227);
xor U413 (N_413,In_133,In_2290);
and U414 (N_414,In_1481,In_646);
nor U415 (N_415,In_2074,In_1486);
nor U416 (N_416,In_1861,In_1532);
nand U417 (N_417,In_2254,In_817);
nand U418 (N_418,In_177,In_1117);
nand U419 (N_419,In_2154,In_1915);
nand U420 (N_420,In_469,In_2300);
nand U421 (N_421,In_1137,In_1238);
nor U422 (N_422,In_558,In_1382);
or U423 (N_423,In_780,In_2062);
or U424 (N_424,In_2427,In_2137);
or U425 (N_425,In_1646,In_1438);
or U426 (N_426,In_2109,In_1707);
or U427 (N_427,In_399,In_310);
and U428 (N_428,In_976,In_1836);
and U429 (N_429,In_1643,In_320);
nor U430 (N_430,In_795,In_67);
nand U431 (N_431,In_868,In_1449);
and U432 (N_432,In_437,In_821);
nand U433 (N_433,In_355,In_253);
nor U434 (N_434,In_675,In_2248);
nor U435 (N_435,In_329,In_1910);
and U436 (N_436,In_1248,In_1278);
nor U437 (N_437,In_1779,In_1483);
nor U438 (N_438,In_1938,In_193);
and U439 (N_439,In_1013,In_2415);
nor U440 (N_440,In_1586,In_1552);
nand U441 (N_441,In_1054,In_804);
nand U442 (N_442,In_2172,In_2276);
nand U443 (N_443,In_1674,In_21);
and U444 (N_444,In_1860,In_1036);
nand U445 (N_445,In_1446,In_623);
and U446 (N_446,In_2068,In_2139);
nand U447 (N_447,In_215,In_1193);
nor U448 (N_448,In_2316,In_1867);
nand U449 (N_449,In_1615,In_1945);
or U450 (N_450,In_2470,In_1565);
nand U451 (N_451,In_1659,In_1575);
xnor U452 (N_452,In_933,In_573);
nor U453 (N_453,In_438,In_1958);
or U454 (N_454,In_156,In_1749);
nand U455 (N_455,In_2176,In_1624);
nor U456 (N_456,In_293,In_986);
nor U457 (N_457,In_771,In_1906);
nand U458 (N_458,In_1563,In_1189);
nand U459 (N_459,In_833,In_532);
or U460 (N_460,In_500,In_248);
or U461 (N_461,In_1487,In_1080);
nand U462 (N_462,In_1498,In_772);
nor U463 (N_463,In_313,In_1079);
and U464 (N_464,In_1497,In_169);
or U465 (N_465,In_1207,In_984);
nor U466 (N_466,In_2308,In_2140);
or U467 (N_467,In_474,In_106);
and U468 (N_468,In_590,In_19);
nor U469 (N_469,In_201,In_1881);
and U470 (N_470,In_665,In_312);
or U471 (N_471,In_883,In_1454);
nor U472 (N_472,In_890,In_844);
nor U473 (N_473,In_75,In_1381);
nor U474 (N_474,In_1350,In_2492);
or U475 (N_475,In_2496,In_2287);
or U476 (N_476,In_1047,In_234);
or U477 (N_477,In_2170,In_1292);
xor U478 (N_478,In_1285,In_2037);
nor U479 (N_479,In_1239,In_353);
nor U480 (N_480,In_1668,In_1120);
xnor U481 (N_481,In_432,In_348);
xor U482 (N_482,In_1900,In_263);
and U483 (N_483,In_2342,In_2023);
and U484 (N_484,In_1895,In_397);
or U485 (N_485,In_2175,In_836);
or U486 (N_486,In_2465,In_1389);
or U487 (N_487,In_2437,In_325);
nand U488 (N_488,In_1174,In_1314);
or U489 (N_489,In_1858,In_856);
or U490 (N_490,In_482,In_825);
and U491 (N_491,In_686,In_985);
nor U492 (N_492,In_37,In_614);
nor U493 (N_493,In_1592,In_2106);
or U494 (N_494,In_163,In_2200);
nor U495 (N_495,In_583,In_1857);
nand U496 (N_496,In_919,In_1360);
xnor U497 (N_497,In_1584,In_2460);
nand U498 (N_498,In_542,In_1173);
nor U499 (N_499,In_1162,In_1252);
or U500 (N_500,In_1582,In_69);
nor U501 (N_501,In_2221,In_1950);
nor U502 (N_502,In_1209,In_1086);
or U503 (N_503,In_1946,In_853);
nor U504 (N_504,In_2031,In_221);
nor U505 (N_505,In_2433,In_202);
nor U506 (N_506,In_693,In_733);
nand U507 (N_507,In_880,In_1283);
and U508 (N_508,In_661,In_1571);
nand U509 (N_509,In_1979,In_1022);
nand U510 (N_510,In_807,In_2285);
xor U511 (N_511,In_409,In_1150);
or U512 (N_512,In_1853,In_2079);
and U513 (N_513,In_476,In_2385);
nor U514 (N_514,In_2160,In_1801);
or U515 (N_515,In_2353,In_581);
nor U516 (N_516,In_388,In_832);
and U517 (N_517,In_136,In_63);
or U518 (N_518,In_213,In_2127);
or U519 (N_519,In_330,In_506);
nor U520 (N_520,In_1480,In_2189);
or U521 (N_521,In_778,In_1845);
nand U522 (N_522,In_1270,In_1100);
nor U523 (N_523,In_1087,In_806);
and U524 (N_524,In_999,In_1869);
nand U525 (N_525,In_1106,In_62);
and U526 (N_526,In_1501,In_649);
or U527 (N_527,In_519,In_2317);
and U528 (N_528,In_1206,In_300);
nand U529 (N_529,In_88,In_96);
and U530 (N_530,In_1590,In_1247);
nor U531 (N_531,In_846,In_307);
and U532 (N_532,In_726,In_1644);
or U533 (N_533,In_1835,In_852);
or U534 (N_534,In_2102,In_1929);
or U535 (N_535,In_1796,In_335);
nor U536 (N_536,In_1447,In_667);
and U537 (N_537,In_1638,In_1837);
nand U538 (N_538,In_1533,In_1972);
nand U539 (N_539,In_1008,In_1831);
or U540 (N_540,In_2292,In_17);
nor U541 (N_541,In_1437,In_2099);
nor U542 (N_542,In_237,In_1887);
nor U543 (N_543,In_2038,In_1469);
or U544 (N_544,In_2243,In_1448);
nor U545 (N_545,In_361,In_1745);
nor U546 (N_546,In_2408,In_2273);
xor U547 (N_547,In_1025,In_512);
nor U548 (N_548,In_1598,In_324);
or U549 (N_549,In_1775,In_505);
nand U550 (N_550,In_1059,In_1810);
and U551 (N_551,In_1772,In_233);
nor U552 (N_552,In_2454,In_338);
nand U553 (N_553,In_1329,In_444);
nand U554 (N_554,In_851,In_2239);
and U555 (N_555,In_105,In_2049);
and U556 (N_556,In_2378,In_1721);
nand U557 (N_557,In_73,In_150);
nand U558 (N_558,In_360,In_451);
or U559 (N_559,In_1841,In_662);
nor U560 (N_560,In_1273,In_58);
nand U561 (N_561,In_1735,In_1988);
nor U562 (N_562,In_1589,In_2);
nor U563 (N_563,In_468,In_477);
nor U564 (N_564,In_1171,In_561);
and U565 (N_565,In_2234,In_1312);
and U566 (N_566,In_1031,In_954);
or U567 (N_567,In_2446,In_1276);
or U568 (N_568,In_2151,In_1545);
or U569 (N_569,In_962,In_484);
nor U570 (N_570,In_651,In_76);
nand U571 (N_571,In_1395,In_185);
and U572 (N_572,In_1773,In_793);
and U573 (N_573,In_670,In_1811);
or U574 (N_574,In_1143,In_98);
nor U575 (N_575,In_2380,In_184);
and U576 (N_576,In_268,In_1280);
nor U577 (N_577,In_1509,In_77);
nor U578 (N_578,In_768,In_1904);
and U579 (N_579,In_1961,In_1762);
nor U580 (N_580,In_1696,In_174);
or U581 (N_581,In_308,In_2216);
or U582 (N_582,In_1739,In_2188);
and U583 (N_583,In_1065,In_6);
or U584 (N_584,In_635,In_172);
or U585 (N_585,In_1323,In_176);
xor U586 (N_586,In_1627,In_1669);
nand U587 (N_587,In_2101,In_562);
and U588 (N_588,In_1547,In_1331);
or U589 (N_589,In_1368,In_2425);
xnor U590 (N_590,In_1005,In_2332);
nor U591 (N_591,In_1655,In_1342);
nor U592 (N_592,In_402,In_2240);
nand U593 (N_593,In_1274,In_7);
nor U594 (N_594,In_2390,In_2352);
and U595 (N_595,In_38,In_539);
nand U596 (N_596,In_1430,In_2041);
nand U597 (N_597,In_1392,In_931);
and U598 (N_598,In_1099,In_1043);
nor U599 (N_599,In_1876,In_2053);
nor U600 (N_600,In_640,In_497);
nor U601 (N_601,In_1578,In_862);
and U602 (N_602,In_794,In_1726);
nand U603 (N_603,In_1477,In_894);
or U604 (N_604,In_2400,In_728);
and U605 (N_605,In_1664,In_357);
and U606 (N_606,In_2205,In_1186);
xor U607 (N_607,In_1579,In_117);
nand U608 (N_608,In_714,In_830);
and U609 (N_609,In_1146,In_550);
nor U610 (N_610,In_1237,In_1444);
and U611 (N_611,In_924,In_257);
nor U612 (N_612,In_1115,In_2309);
and U613 (N_613,In_1987,In_458);
nand U614 (N_614,In_1163,In_1816);
nand U615 (N_615,In_1212,In_452);
nor U616 (N_616,In_396,In_1516);
or U617 (N_617,In_823,In_1982);
nor U618 (N_618,In_1097,In_811);
nand U619 (N_619,In_269,In_1596);
nor U620 (N_620,In_2207,In_537);
or U621 (N_621,In_2335,In_1319);
or U622 (N_622,In_572,In_1974);
nor U623 (N_623,In_674,In_447);
and U624 (N_624,In_927,In_192);
and U625 (N_625,In_1198,In_284);
nor U626 (N_626,In_2379,In_742);
or U627 (N_627,In_885,In_1421);
xnor U628 (N_628,In_1531,In_896);
and U629 (N_629,In_1445,In_1378);
and U630 (N_630,In_1854,In_1400);
nor U631 (N_631,In_224,In_2028);
nand U632 (N_632,In_1076,In_1370);
and U633 (N_633,In_245,In_1466);
nand U634 (N_634,In_1057,In_1257);
nor U635 (N_635,In_1258,In_1436);
and U636 (N_636,In_2231,In_149);
and U637 (N_637,In_1640,In_1320);
nor U638 (N_638,In_957,In_1216);
nand U639 (N_639,In_278,In_1182);
or U640 (N_640,In_1716,In_731);
or U641 (N_641,In_367,In_1684);
or U642 (N_642,In_1068,In_239);
and U643 (N_643,In_140,In_691);
nor U644 (N_644,In_392,In_128);
nand U645 (N_645,In_1453,In_1295);
nor U646 (N_646,In_372,In_650);
or U647 (N_647,In_418,In_781);
nor U648 (N_648,In_1757,In_2346);
and U649 (N_649,In_1309,In_2092);
and U650 (N_650,In_1609,In_770);
or U651 (N_651,In_1422,In_2161);
and U652 (N_652,In_1340,In_840);
or U653 (N_653,In_1939,In_1393);
and U654 (N_654,In_2261,In_2069);
nand U655 (N_655,In_753,In_899);
nand U656 (N_656,In_599,In_1495);
or U657 (N_657,In_272,In_1577);
nor U658 (N_658,In_723,In_15);
or U659 (N_659,In_376,In_2148);
and U660 (N_660,In_1694,In_1363);
nor U661 (N_661,In_1642,In_1217);
and U662 (N_662,In_1593,In_407);
and U663 (N_663,In_2409,In_466);
or U664 (N_664,In_524,In_1731);
and U665 (N_665,In_1800,In_763);
and U666 (N_666,In_2479,In_2414);
nand U667 (N_667,In_1066,In_2473);
nand U668 (N_668,In_2270,In_22);
nand U669 (N_669,In_1474,In_574);
and U670 (N_670,In_712,In_700);
or U671 (N_671,In_1830,In_2339);
and U672 (N_672,In_103,In_1675);
nor U673 (N_673,In_1636,In_1308);
nor U674 (N_674,In_937,In_2289);
or U675 (N_675,In_2047,In_704);
or U676 (N_676,In_370,In_2156);
nand U677 (N_677,In_688,In_1903);
nand U678 (N_678,In_818,In_211);
or U679 (N_679,In_2077,In_1905);
nor U680 (N_680,In_1159,In_1056);
nor U681 (N_681,In_739,In_1912);
nor U682 (N_682,In_1298,In_2422);
or U683 (N_683,In_2284,In_1253);
nor U684 (N_684,In_1754,In_124);
and U685 (N_685,In_1410,In_1591);
nand U686 (N_686,In_406,In_708);
nand U687 (N_687,In_2245,In_290);
nand U688 (N_688,In_1353,In_1425);
nor U689 (N_689,In_974,In_2491);
nor U690 (N_690,In_2484,In_1663);
or U691 (N_691,In_2432,In_926);
and U692 (N_692,In_544,In_1889);
nor U693 (N_693,In_24,In_1542);
or U694 (N_694,In_766,In_1536);
or U695 (N_695,In_944,In_465);
nor U696 (N_696,In_1429,In_786);
nand U697 (N_697,In_1695,In_929);
or U698 (N_698,In_982,In_264);
nor U699 (N_699,In_2179,In_2373);
nand U700 (N_700,In_1061,In_2445);
nand U701 (N_701,In_514,In_697);
nand U702 (N_702,In_400,In_2008);
and U703 (N_703,In_50,In_1907);
and U704 (N_704,In_1102,In_513);
or U705 (N_705,In_205,In_1623);
xnor U706 (N_706,In_107,In_116);
nor U707 (N_707,In_1465,In_1527);
nor U708 (N_708,In_1617,In_110);
nor U709 (N_709,In_1865,In_1024);
nand U710 (N_710,In_1618,In_610);
nor U711 (N_711,In_2010,In_2486);
or U712 (N_712,In_2225,In_998);
or U713 (N_713,In_1817,In_1266);
or U714 (N_714,In_784,In_2398);
or U715 (N_715,In_1740,In_1849);
or U716 (N_716,In_1711,In_182);
nor U717 (N_717,In_1996,In_381);
and U718 (N_718,In_1269,In_633);
nand U719 (N_719,In_606,In_72);
nor U720 (N_720,In_1467,In_621);
or U721 (N_721,In_1222,In_415);
nor U722 (N_722,In_303,In_1048);
or U723 (N_723,In_2459,In_122);
or U724 (N_724,In_2301,In_1897);
nor U725 (N_725,In_1661,In_1391);
or U726 (N_726,In_2097,In_291);
nor U727 (N_727,In_1875,In_705);
and U728 (N_728,In_1561,In_504);
and U729 (N_729,In_412,In_1138);
nor U730 (N_730,In_1010,In_1901);
and U731 (N_731,In_1064,In_1687);
nor U732 (N_732,In_1806,In_1607);
and U733 (N_733,In_509,In_1194);
or U734 (N_734,In_345,In_1204);
or U735 (N_735,In_2098,In_1518);
nor U736 (N_736,In_1829,In_2464);
nor U737 (N_737,In_137,In_1181);
nor U738 (N_738,In_2162,In_2381);
or U739 (N_739,In_737,In_1014);
and U740 (N_740,In_946,In_761);
or U741 (N_741,In_2267,In_595);
nand U742 (N_742,In_736,In_2468);
nand U743 (N_743,In_1045,In_2456);
and U744 (N_744,In_480,In_2311);
nor U745 (N_745,In_1141,In_1215);
and U746 (N_746,In_1748,In_455);
nor U747 (N_747,In_230,In_1362);
and U748 (N_748,In_1743,In_2306);
xnor U749 (N_749,In_131,In_1995);
xnor U750 (N_750,In_175,In_981);
or U751 (N_751,In_1197,In_2350);
and U752 (N_752,In_677,In_2480);
and U753 (N_753,In_457,In_578);
xor U754 (N_754,In_639,In_135);
xnor U755 (N_755,In_754,In_917);
nor U756 (N_756,In_71,In_1334);
xnor U757 (N_757,In_350,In_1185);
or U758 (N_758,In_1523,In_1626);
nor U759 (N_759,In_1847,In_1110);
nor U760 (N_760,In_2298,In_2104);
nor U761 (N_761,In_2374,In_14);
nor U762 (N_762,In_1202,In_375);
and U763 (N_763,In_760,In_1398);
nor U764 (N_764,In_1990,In_1478);
or U765 (N_765,In_1597,In_1470);
and U766 (N_766,In_1883,In_535);
nand U767 (N_767,In_555,In_2214);
or U768 (N_768,In_2022,In_1020);
or U769 (N_769,In_1256,In_305);
or U770 (N_770,In_1044,In_1891);
xnor U771 (N_771,In_187,In_1490);
nand U772 (N_772,In_847,In_475);
nand U773 (N_773,In_190,In_1882);
xor U774 (N_774,In_746,In_1240);
or U775 (N_775,In_809,In_802);
nand U776 (N_776,In_285,In_2084);
and U777 (N_777,In_33,In_1954);
and U778 (N_778,In_1734,In_540);
or U779 (N_779,In_1993,In_1947);
nand U780 (N_780,In_1580,In_1228);
nor U781 (N_781,In_1610,In_1632);
and U782 (N_782,In_2169,In_2327);
and U783 (N_783,In_1981,In_624);
nor U784 (N_784,In_473,In_1500);
and U785 (N_785,In_2001,In_664);
nand U786 (N_786,In_2164,In_2402);
and U787 (N_787,In_152,In_413);
nor U788 (N_788,In_422,In_2236);
nor U789 (N_789,In_587,In_1333);
or U790 (N_790,In_1786,In_2466);
nor U791 (N_791,In_861,In_2103);
and U792 (N_792,In_1619,In_1699);
nand U793 (N_793,In_968,In_2294);
and U794 (N_794,In_2182,In_1085);
or U795 (N_795,In_921,In_909);
or U796 (N_796,In_198,In_1502);
or U797 (N_797,In_709,In_1807);
and U798 (N_798,In_1063,In_2493);
nand U799 (N_799,In_797,In_955);
nor U800 (N_800,In_235,In_845);
and U801 (N_801,In_2113,In_191);
nor U802 (N_802,In_2142,In_1264);
nor U803 (N_803,In_1737,In_138);
nor U804 (N_804,In_1160,In_1211);
nand U805 (N_805,In_1476,In_1761);
and U806 (N_806,In_891,In_2251);
nor U807 (N_807,In_799,In_1600);
nor U808 (N_808,In_2462,In_1689);
or U809 (N_809,In_2364,In_1139);
nand U810 (N_810,In_1683,In_507);
nand U811 (N_811,In_395,In_554);
or U812 (N_812,In_757,In_2429);
or U813 (N_813,In_125,In_1394);
nor U814 (N_814,In_1710,In_2222);
nand U815 (N_815,In_1037,In_1994);
and U816 (N_816,In_1300,In_1213);
or U817 (N_817,In_776,In_332);
nand U818 (N_818,In_46,In_336);
xor U819 (N_819,In_227,In_2073);
and U820 (N_820,In_969,In_787);
and U821 (N_821,In_2489,In_1376);
or U822 (N_822,In_1783,In_1440);
nor U823 (N_823,In_884,In_2420);
nor U824 (N_824,In_1650,In_905);
xor U825 (N_825,In_2163,In_1339);
nor U826 (N_826,In_2391,In_1569);
or U827 (N_827,In_1348,In_684);
nand U828 (N_828,In_44,In_774);
nor U829 (N_829,In_2312,In_1310);
or U830 (N_830,In_470,In_471);
nand U831 (N_831,In_1485,In_2124);
nor U832 (N_832,In_534,In_963);
nand U833 (N_833,In_231,In_1304);
and U834 (N_834,In_1971,In_2052);
nand U835 (N_835,In_461,In_967);
and U836 (N_836,In_2198,In_401);
nand U837 (N_837,In_2105,In_13);
nand U838 (N_838,In_2138,In_1524);
nand U839 (N_839,In_1459,In_745);
nand U840 (N_840,In_1871,In_1594);
nor U841 (N_841,In_956,In_881);
nor U842 (N_842,In_2413,In_1060);
and U843 (N_843,In_1732,In_1635);
and U844 (N_844,In_2054,In_334);
and U845 (N_845,In_1241,In_517);
or U846 (N_846,In_2372,In_1886);
nand U847 (N_847,In_878,In_1926);
and U848 (N_848,In_602,In_1788);
nor U849 (N_849,In_2125,In_2083);
or U850 (N_850,In_1042,In_2423);
or U851 (N_851,In_2020,In_1464);
and U852 (N_852,In_2195,In_1121);
nor U853 (N_853,In_256,In_456);
or U854 (N_854,In_1892,In_1396);
nor U855 (N_855,In_887,In_1980);
or U856 (N_856,In_657,In_2111);
or U857 (N_857,In_822,In_2112);
and U858 (N_858,In_1195,In_801);
and U859 (N_859,In_1261,In_250);
nor U860 (N_860,In_2310,In_679);
or U861 (N_861,In_592,In_1177);
or U862 (N_862,In_2191,In_2388);
or U863 (N_863,In_1528,In_115);
nor U864 (N_864,In_1251,In_2302);
nand U865 (N_865,In_2171,In_1933);
nor U866 (N_866,In_2452,In_1714);
or U867 (N_867,In_384,In_1098);
nor U868 (N_868,In_508,In_570);
nand U869 (N_869,In_898,In_1595);
and U870 (N_870,In_26,In_317);
and U871 (N_871,In_589,In_1572);
nand U872 (N_872,In_751,In_2286);
nand U873 (N_873,In_1220,In_2278);
nor U874 (N_874,In_183,In_112);
and U875 (N_875,In_1461,In_702);
nor U876 (N_876,In_1771,In_228);
and U877 (N_877,In_1678,In_1514);
nor U878 (N_878,In_1752,In_785);
and U879 (N_879,In_340,In_1029);
nor U880 (N_880,In_1908,In_907);
nor U881 (N_881,In_1200,In_1599);
or U882 (N_882,In_972,In_1581);
or U883 (N_883,In_206,In_1658);
or U884 (N_884,In_1129,In_888);
and U885 (N_885,In_430,In_315);
or U886 (N_886,In_1864,In_2412);
nand U887 (N_887,In_1361,In_1026);
nor U888 (N_888,In_2450,In_2180);
and U889 (N_889,In_1621,In_719);
and U890 (N_890,In_1420,In_2330);
or U891 (N_891,In_545,In_803);
and U892 (N_892,In_902,In_252);
or U893 (N_893,In_1511,In_494);
nand U894 (N_894,In_347,In_873);
nor U895 (N_895,In_1336,In_1427);
nor U896 (N_896,In_1639,In_328);
nor U897 (N_897,In_1148,In_549);
nand U898 (N_898,In_577,In_1549);
or U899 (N_899,In_1359,In_1776);
or U900 (N_900,In_127,In_1924);
nand U901 (N_901,In_2419,In_942);
and U902 (N_902,In_5,In_2082);
or U903 (N_903,In_216,In_859);
nand U904 (N_904,In_2244,In_831);
nor U905 (N_905,In_865,In_582);
nand U906 (N_906,In_1936,In_2081);
nand U907 (N_907,In_2421,In_1281);
nand U908 (N_908,In_1260,In_1052);
or U909 (N_909,In_1515,In_490);
or U910 (N_910,In_195,In_875);
and U911 (N_911,In_2166,In_2048);
nor U912 (N_912,In_1633,In_1221);
xor U913 (N_913,In_569,In_1327);
nor U914 (N_914,In_1428,In_2223);
or U915 (N_915,In_49,In_1113);
or U916 (N_916,In_671,In_655);
or U917 (N_917,In_1344,In_365);
nand U918 (N_918,In_1373,In_1540);
nand U919 (N_919,In_601,In_1942);
nand U920 (N_920,In_1691,In_101);
nand U921 (N_921,In_2193,In_2228);
or U922 (N_922,In_258,In_1049);
or U923 (N_923,In_2173,In_722);
xnor U924 (N_924,In_960,In_2396);
nor U925 (N_925,In_2226,In_247);
or U926 (N_926,In_146,In_525);
and U927 (N_927,In_1898,In_547);
and U928 (N_928,In_157,In_893);
nor U929 (N_929,In_521,In_2208);
or U930 (N_930,In_613,In_1084);
and U931 (N_931,In_2146,In_2324);
nor U932 (N_932,In_2448,In_2029);
nor U933 (N_933,In_958,In_1766);
nor U934 (N_934,In_8,In_2487);
nor U935 (N_935,In_1103,In_718);
nor U936 (N_936,In_1433,In_1704);
nor U937 (N_937,In_1125,In_74);
nand U938 (N_938,In_1846,In_66);
and U939 (N_939,In_857,In_2067);
nand U940 (N_940,In_1890,In_1144);
and U941 (N_941,In_126,In_449);
xnor U942 (N_942,In_436,In_459);
or U943 (N_943,In_619,In_934);
nor U944 (N_944,In_219,In_789);
nand U945 (N_945,In_2455,In_2483);
nor U946 (N_946,In_1302,In_1508);
and U947 (N_947,In_1525,In_566);
or U948 (N_948,In_45,In_84);
nand U949 (N_949,In_1116,In_2280);
nor U950 (N_950,In_553,In_1645);
xnor U951 (N_951,In_421,In_1223);
and U952 (N_952,In_2269,In_54);
nor U953 (N_953,In_1038,In_1978);
nor U954 (N_954,In_153,In_2212);
nand U955 (N_955,In_1003,In_1157);
or U956 (N_956,In_1169,In_1231);
or U957 (N_957,In_1496,In_43);
nor U958 (N_958,In_782,In_654);
nand U959 (N_959,In_1649,In_162);
or U960 (N_960,In_2100,In_1560);
nor U961 (N_961,In_1,In_2085);
and U962 (N_962,In_2336,In_57);
nand U963 (N_963,In_752,In_1548);
nand U964 (N_964,In_1504,In_2177);
nor U965 (N_965,In_1088,In_923);
xnor U966 (N_966,In_450,In_139);
xnor U967 (N_967,In_2377,In_1782);
nand U968 (N_968,In_1041,In_2118);
nand U969 (N_969,In_1161,In_886);
and U970 (N_970,In_515,In_53);
nand U971 (N_971,In_1744,In_1322);
nand U972 (N_972,In_2192,In_2123);
nand U973 (N_973,In_1706,In_1828);
nor U974 (N_974,In_40,In_2014);
nor U975 (N_975,In_1006,In_935);
xor U976 (N_976,In_1656,In_598);
nand U977 (N_977,In_1473,In_1092);
and U978 (N_978,In_2210,In_916);
and U979 (N_979,In_2305,In_487);
nand U980 (N_980,In_229,In_1423);
or U981 (N_981,In_2263,In_28);
and U982 (N_982,In_1190,In_151);
and U983 (N_983,In_1603,In_1409);
or U984 (N_984,In_251,In_1729);
and U985 (N_985,In_1909,In_648);
and U986 (N_986,In_1040,In_644);
nor U987 (N_987,In_405,In_1510);
and U988 (N_988,In_2247,In_2485);
and U989 (N_989,In_2149,In_1018);
and U990 (N_990,In_563,In_2334);
and U991 (N_991,In_178,In_1492);
nand U992 (N_992,In_1033,In_892);
nand U993 (N_993,In_877,In_1016);
nor U994 (N_994,In_2253,In_304);
or U995 (N_995,In_241,In_2059);
and U996 (N_996,In_1201,In_2436);
nor U997 (N_997,In_2315,In_2323);
nand U998 (N_998,In_584,In_1931);
nand U999 (N_999,In_543,In_1188);
nor U1000 (N_1000,In_382,In_1077);
and U1001 (N_1001,In_627,In_2328);
or U1002 (N_1002,In_1418,In_1386);
and U1003 (N_1003,In_2338,In_2295);
nand U1004 (N_1004,In_1613,In_1637);
nor U1005 (N_1005,In_1975,In_204);
xor U1006 (N_1006,In_1702,In_1625);
and U1007 (N_1007,In_850,In_65);
and U1008 (N_1008,In_2375,In_716);
nor U1009 (N_1009,In_724,In_1838);
nor U1010 (N_1010,In_2255,In_1397);
nor U1011 (N_1011,In_2168,In_1119);
and U1012 (N_1012,In_1236,In_222);
or U1013 (N_1013,In_814,In_2181);
nand U1014 (N_1014,In_200,In_1826);
or U1015 (N_1015,In_1612,In_277);
xnor U1016 (N_1016,In_1191,In_748);
and U1017 (N_1017,In_1341,In_2055);
nor U1018 (N_1018,In_1793,In_1034);
or U1019 (N_1019,In_548,In_2499);
nand U1020 (N_1020,In_604,In_756);
nor U1021 (N_1021,In_380,In_1677);
nor U1022 (N_1022,In_2411,In_97);
and U1023 (N_1023,In_306,In_179);
and U1024 (N_1024,In_1035,In_260);
nor U1025 (N_1025,In_987,In_1665);
nor U1026 (N_1026,In_2183,In_1325);
nor U1027 (N_1027,In_1856,In_1458);
and U1028 (N_1028,In_2478,In_1136);
and U1029 (N_1029,In_2065,In_1985);
or U1030 (N_1030,In_559,In_966);
nor U1031 (N_1031,In_2025,In_42);
or U1032 (N_1032,In_658,In_1356);
and U1033 (N_1033,In_1812,In_1315);
or U1034 (N_1034,In_1218,In_1297);
nand U1035 (N_1035,In_155,In_2096);
or U1036 (N_1036,In_486,In_2007);
and U1037 (N_1037,In_1690,In_1553);
nand U1038 (N_1038,In_1568,In_1872);
nor U1039 (N_1039,In_1176,In_1385);
xnor U1040 (N_1040,In_1802,In_267);
nor U1041 (N_1041,In_2256,In_1795);
nor U1042 (N_1042,In_1208,In_1957);
nand U1043 (N_1043,In_374,In_715);
nand U1044 (N_1044,In_2026,In_1557);
nand U1045 (N_1045,In_209,In_1870);
or U1046 (N_1046,In_1879,In_2090);
and U1047 (N_1047,In_2439,In_1747);
xor U1048 (N_1048,In_2249,In_2145);
or U1049 (N_1049,In_2304,In_145);
or U1050 (N_1050,In_398,In_262);
and U1051 (N_1051,In_2005,In_841);
nor U1052 (N_1052,In_1789,In_828);
and U1053 (N_1053,In_2194,In_104);
nand U1054 (N_1054,In_1311,In_575);
and U1055 (N_1055,In_882,In_1916);
or U1056 (N_1056,In_977,In_266);
nand U1057 (N_1057,In_485,In_203);
and U1058 (N_1058,In_2039,In_2155);
or U1059 (N_1059,In_1673,In_1364);
nand U1060 (N_1060,In_1813,In_2036);
and U1061 (N_1061,In_1713,In_531);
or U1062 (N_1062,In_160,In_1808);
and U1063 (N_1063,In_1493,In_1920);
nor U1064 (N_1064,In_863,In_2361);
or U1065 (N_1065,In_1133,In_522);
xor U1066 (N_1066,In_1848,In_669);
and U1067 (N_1067,In_1246,In_808);
or U1068 (N_1068,In_2217,In_600);
and U1069 (N_1069,In_949,In_2116);
and U1070 (N_1070,In_1235,In_1629);
and U1071 (N_1071,In_378,In_2066);
nor U1072 (N_1072,In_1641,In_2482);
and U1073 (N_1073,In_2144,In_523);
or U1074 (N_1074,In_2006,In_1685);
and U1075 (N_1075,In_897,In_287);
and U1076 (N_1076,In_2257,In_1850);
nor U1077 (N_1077,In_529,In_1968);
nand U1078 (N_1078,In_2438,In_1345);
and U1079 (N_1079,In_1142,In_1940);
and U1080 (N_1080,In_429,In_2227);
and U1081 (N_1081,In_2219,In_928);
and U1082 (N_1082,In_441,In_1520);
and U1083 (N_1083,In_1019,In_1371);
and U1084 (N_1084,In_1794,In_1653);
and U1085 (N_1085,In_32,In_2369);
and U1086 (N_1086,In_2133,In_1804);
nand U1087 (N_1087,In_167,In_1697);
nor U1088 (N_1088,In_925,In_1111);
or U1089 (N_1089,In_2447,In_1756);
or U1090 (N_1090,In_1719,In_271);
or U1091 (N_1091,In_2341,In_68);
and U1092 (N_1092,In_1369,In_2232);
or U1093 (N_1093,In_478,In_660);
nor U1094 (N_1094,In_835,In_220);
nand U1095 (N_1095,In_261,In_377);
nand U1096 (N_1096,In_2357,In_796);
nand U1097 (N_1097,In_685,In_2157);
nand U1098 (N_1098,In_1654,In_242);
nand U1099 (N_1099,In_1997,In_983);
and U1100 (N_1100,In_2032,In_435);
nand U1101 (N_1101,In_1521,In_647);
and U1102 (N_1102,In_1412,In_603);
or U1103 (N_1103,In_1001,In_1471);
nand U1104 (N_1104,In_2158,In_1180);
or U1105 (N_1105,In_448,In_618);
xor U1106 (N_1106,In_255,In_1284);
nor U1107 (N_1107,In_1007,In_404);
or U1108 (N_1108,In_1791,In_52);
nand U1109 (N_1109,In_339,In_1432);
nor U1110 (N_1110,In_2115,In_2428);
nor U1111 (N_1111,In_1267,In_1574);
nor U1112 (N_1112,In_1456,In_1570);
nand U1113 (N_1113,In_694,In_1401);
or U1114 (N_1114,In_1050,In_311);
nor U1115 (N_1115,In_1021,In_2389);
and U1116 (N_1116,In_788,In_383);
nor U1117 (N_1117,In_2204,In_1833);
and U1118 (N_1118,In_1526,In_1134);
xor U1119 (N_1119,In_713,In_2013);
nand U1120 (N_1120,In_920,In_1123);
nor U1121 (N_1121,In_113,In_1399);
and U1122 (N_1122,In_918,In_368);
nand U1123 (N_1123,In_462,In_1986);
or U1124 (N_1124,In_1249,In_912);
nor U1125 (N_1125,In_2015,In_118);
nor U1126 (N_1126,In_626,In_605);
nand U1127 (N_1127,In_764,In_1703);
or U1128 (N_1128,In_2063,In_551);
and U1129 (N_1129,In_352,In_1728);
nand U1130 (N_1130,In_2199,In_92);
or U1131 (N_1131,In_333,In_735);
and U1132 (N_1132,In_1250,In_1919);
or U1133 (N_1133,In_2399,In_2405);
xor U1134 (N_1134,In_1165,In_805);
or U1135 (N_1135,In_2086,In_243);
or U1136 (N_1136,In_454,In_100);
nor U1137 (N_1137,In_1132,In_2271);
and U1138 (N_1138,In_1583,In_1701);
or U1139 (N_1139,In_1265,In_1140);
or U1140 (N_1140,In_585,In_411);
nand U1141 (N_1141,In_36,In_1519);
or U1142 (N_1142,In_2274,In_166);
and U1143 (N_1143,In_1877,In_1288);
and U1144 (N_1144,In_309,In_1666);
nand U1145 (N_1145,In_1380,In_2441);
and U1146 (N_1146,In_1823,In_440);
and U1147 (N_1147,In_214,In_2319);
nand U1148 (N_1148,In_727,In_744);
and U1149 (N_1149,In_2220,In_121);
nor U1150 (N_1150,In_518,In_876);
nor U1151 (N_1151,In_2291,In_2110);
nor U1152 (N_1152,In_588,In_244);
nand U1153 (N_1153,In_292,In_2174);
and U1154 (N_1154,In_1279,In_1724);
nand U1155 (N_1155,In_827,In_1567);
nor U1156 (N_1156,In_1374,In_1647);
nor U1157 (N_1157,In_226,In_351);
and U1158 (N_1158,In_711,In_631);
nand U1159 (N_1159,In_1680,In_41);
nor U1160 (N_1160,In_1755,In_25);
nor U1161 (N_1161,In_959,In_499);
nand U1162 (N_1162,In_652,In_323);
nor U1163 (N_1163,In_1843,In_295);
nor U1164 (N_1164,In_1472,In_901);
nor U1165 (N_1165,In_123,In_502);
or U1166 (N_1166,In_961,In_349);
nor U1167 (N_1167,In_199,In_643);
nor U1168 (N_1168,In_2130,In_2393);
nor U1169 (N_1169,In_2431,In_93);
and U1170 (N_1170,In_911,In_2095);
and U1171 (N_1171,In_1317,In_299);
nor U1172 (N_1172,In_663,In_1862);
nand U1173 (N_1173,In_434,In_1951);
nand U1174 (N_1174,In_70,In_1733);
xnor U1175 (N_1175,In_1277,In_1822);
or U1176 (N_1176,In_1294,In_1229);
and U1177 (N_1177,In_321,In_1343);
nor U1178 (N_1178,In_147,In_536);
or U1179 (N_1179,In_154,In_12);
and U1180 (N_1180,In_2058,In_90);
xor U1181 (N_1181,In_2404,In_281);
and U1182 (N_1182,In_108,In_1863);
nand U1183 (N_1183,In_2185,In_1167);
and U1184 (N_1184,In_2477,In_1338);
or U1185 (N_1185,In_1943,In_246);
and U1186 (N_1186,In_2153,In_1686);
and U1187 (N_1187,In_1657,In_1538);
nor U1188 (N_1188,In_1112,In_1262);
or U1189 (N_1189,In_1667,In_2495);
and U1190 (N_1190,In_2457,In_463);
or U1191 (N_1191,In_1263,In_538);
or U1192 (N_1192,In_1792,In_61);
and U1193 (N_1193,In_30,In_363);
or U1194 (N_1194,In_1537,In_2314);
or U1195 (N_1195,In_319,In_414);
nor U1196 (N_1196,In_858,In_1819);
or U1197 (N_1197,In_1774,In_1917);
nand U1198 (N_1198,In_2233,In_467);
nor U1199 (N_1199,In_1259,In_2165);
nand U1200 (N_1200,In_1475,In_637);
or U1201 (N_1201,In_1770,In_879);
nor U1202 (N_1202,In_2296,In_1966);
nand U1203 (N_1203,In_1955,In_2370);
or U1204 (N_1204,In_1852,In_390);
and U1205 (N_1205,In_2394,In_2246);
and U1206 (N_1206,In_1388,In_196);
nor U1207 (N_1207,In_1243,In_1517);
nor U1208 (N_1208,In_1179,In_294);
and U1209 (N_1209,In_611,In_2230);
or U1210 (N_1210,In_1825,In_2268);
and U1211 (N_1211,In_111,In_1977);
nand U1212 (N_1212,In_2434,In_134);
nand U1213 (N_1213,In_546,In_297);
nand U1214 (N_1214,In_1219,In_971);
nand U1215 (N_1215,In_609,In_1404);
xnor U1216 (N_1216,In_1725,In_1611);
nor U1217 (N_1217,In_1893,In_1832);
and U1218 (N_1218,In_593,In_741);
nand U1219 (N_1219,In_2076,In_1614);
or U1220 (N_1220,In_870,In_1383);
nor U1221 (N_1221,In_1291,In_2453);
nor U1222 (N_1222,In_1738,In_843);
nand U1223 (N_1223,In_2345,In_1002);
nor U1224 (N_1224,In_2108,In_560);
or U1225 (N_1225,In_433,In_597);
nor U1226 (N_1226,In_1387,In_1039);
nor U1227 (N_1227,In_503,In_683);
and U1228 (N_1228,In_1969,In_1787);
xor U1229 (N_1229,In_1566,In_1457);
nand U1230 (N_1230,In_1131,In_1479);
or U1231 (N_1231,In_1805,In_369);
or U1232 (N_1232,In_2359,In_617);
nand U1233 (N_1233,In_391,In_812);
nor U1234 (N_1234,In_1307,In_1494);
or U1235 (N_1235,In_1868,In_171);
and U1236 (N_1236,In_1708,In_254);
or U1237 (N_1237,In_1820,In_1763);
nor U1238 (N_1238,In_2159,In_273);
or U1239 (N_1239,In_1004,In_1717);
nor U1240 (N_1240,In_1379,In_453);
or U1241 (N_1241,In_2016,In_2042);
or U1242 (N_1242,In_1351,In_1091);
and U1243 (N_1243,In_425,In_464);
nand U1244 (N_1244,In_1809,In_1544);
nor U1245 (N_1245,In_2430,In_356);
or U1246 (N_1246,In_1682,In_1306);
nor U1247 (N_1247,In_1559,In_2002);
or U1248 (N_1248,In_2299,In_223);
or U1249 (N_1249,In_2051,In_1652);
and U1250 (N_1250,In_190,In_320);
nor U1251 (N_1251,In_2399,In_1861);
nand U1252 (N_1252,In_659,In_2437);
nor U1253 (N_1253,In_1462,In_1131);
nand U1254 (N_1254,In_35,In_1645);
and U1255 (N_1255,In_604,In_1804);
and U1256 (N_1256,In_1967,In_1679);
nor U1257 (N_1257,In_1404,In_2051);
and U1258 (N_1258,In_2170,In_2141);
nand U1259 (N_1259,In_1343,In_73);
nand U1260 (N_1260,In_2454,In_864);
or U1261 (N_1261,In_722,In_1375);
or U1262 (N_1262,In_572,In_1363);
nand U1263 (N_1263,In_1464,In_2156);
nor U1264 (N_1264,In_2157,In_527);
and U1265 (N_1265,In_2334,In_887);
or U1266 (N_1266,In_1435,In_343);
and U1267 (N_1267,In_2016,In_2247);
and U1268 (N_1268,In_1691,In_549);
nand U1269 (N_1269,In_2422,In_1092);
nand U1270 (N_1270,In_1048,In_1190);
nand U1271 (N_1271,In_651,In_2348);
nand U1272 (N_1272,In_545,In_1687);
nand U1273 (N_1273,In_1288,In_1817);
nor U1274 (N_1274,In_76,In_1016);
or U1275 (N_1275,In_483,In_427);
nor U1276 (N_1276,In_1576,In_241);
or U1277 (N_1277,In_1631,In_142);
nand U1278 (N_1278,In_136,In_1156);
nor U1279 (N_1279,In_2331,In_165);
nor U1280 (N_1280,In_2306,In_2130);
or U1281 (N_1281,In_549,In_627);
nand U1282 (N_1282,In_342,In_2401);
and U1283 (N_1283,In_1040,In_645);
and U1284 (N_1284,In_1695,In_1929);
and U1285 (N_1285,In_1059,In_2135);
or U1286 (N_1286,In_2036,In_1539);
nand U1287 (N_1287,In_721,In_1611);
xnor U1288 (N_1288,In_1372,In_1811);
nor U1289 (N_1289,In_829,In_1365);
nor U1290 (N_1290,In_2441,In_2014);
nand U1291 (N_1291,In_390,In_1470);
and U1292 (N_1292,In_781,In_2418);
nor U1293 (N_1293,In_2302,In_945);
nor U1294 (N_1294,In_1387,In_1862);
nand U1295 (N_1295,In_955,In_784);
xnor U1296 (N_1296,In_602,In_731);
nand U1297 (N_1297,In_1828,In_1890);
or U1298 (N_1298,In_969,In_836);
nor U1299 (N_1299,In_1153,In_554);
or U1300 (N_1300,In_985,In_1988);
nor U1301 (N_1301,In_262,In_1154);
and U1302 (N_1302,In_670,In_901);
nor U1303 (N_1303,In_93,In_1043);
nand U1304 (N_1304,In_547,In_308);
or U1305 (N_1305,In_435,In_579);
nand U1306 (N_1306,In_91,In_1991);
nor U1307 (N_1307,In_109,In_2485);
nor U1308 (N_1308,In_2166,In_347);
or U1309 (N_1309,In_2488,In_31);
or U1310 (N_1310,In_1302,In_2461);
or U1311 (N_1311,In_1881,In_1070);
nand U1312 (N_1312,In_813,In_2080);
or U1313 (N_1313,In_801,In_529);
or U1314 (N_1314,In_2275,In_1284);
nor U1315 (N_1315,In_699,In_2405);
or U1316 (N_1316,In_440,In_1763);
nor U1317 (N_1317,In_2420,In_3);
or U1318 (N_1318,In_983,In_585);
nor U1319 (N_1319,In_1862,In_1537);
and U1320 (N_1320,In_784,In_1589);
nand U1321 (N_1321,In_17,In_1778);
or U1322 (N_1322,In_1571,In_1840);
nor U1323 (N_1323,In_2240,In_1998);
nor U1324 (N_1324,In_1648,In_553);
nor U1325 (N_1325,In_2361,In_971);
nand U1326 (N_1326,In_538,In_370);
and U1327 (N_1327,In_1852,In_604);
and U1328 (N_1328,In_1056,In_869);
nand U1329 (N_1329,In_1537,In_2348);
nor U1330 (N_1330,In_2273,In_2219);
nand U1331 (N_1331,In_1855,In_1846);
xnor U1332 (N_1332,In_1996,In_253);
or U1333 (N_1333,In_2472,In_2477);
or U1334 (N_1334,In_1519,In_2440);
nand U1335 (N_1335,In_989,In_54);
nand U1336 (N_1336,In_2300,In_62);
and U1337 (N_1337,In_313,In_159);
nand U1338 (N_1338,In_636,In_2146);
and U1339 (N_1339,In_190,In_1878);
or U1340 (N_1340,In_2436,In_933);
or U1341 (N_1341,In_1481,In_2080);
nand U1342 (N_1342,In_2416,In_473);
or U1343 (N_1343,In_2204,In_209);
or U1344 (N_1344,In_2106,In_271);
nand U1345 (N_1345,In_185,In_1861);
or U1346 (N_1346,In_2263,In_1542);
nor U1347 (N_1347,In_404,In_700);
and U1348 (N_1348,In_860,In_2069);
and U1349 (N_1349,In_40,In_879);
nand U1350 (N_1350,In_1866,In_155);
nand U1351 (N_1351,In_199,In_1314);
nand U1352 (N_1352,In_505,In_20);
nand U1353 (N_1353,In_13,In_371);
nor U1354 (N_1354,In_1661,In_1313);
or U1355 (N_1355,In_1644,In_406);
or U1356 (N_1356,In_589,In_1996);
or U1357 (N_1357,In_2266,In_61);
nand U1358 (N_1358,In_1342,In_287);
or U1359 (N_1359,In_2419,In_2210);
and U1360 (N_1360,In_846,In_2370);
and U1361 (N_1361,In_53,In_1008);
nand U1362 (N_1362,In_769,In_208);
or U1363 (N_1363,In_860,In_57);
xor U1364 (N_1364,In_2366,In_1560);
nor U1365 (N_1365,In_1967,In_489);
and U1366 (N_1366,In_768,In_1316);
nor U1367 (N_1367,In_2058,In_2223);
and U1368 (N_1368,In_1230,In_180);
nor U1369 (N_1369,In_1860,In_2352);
or U1370 (N_1370,In_1747,In_1379);
or U1371 (N_1371,In_1358,In_885);
xor U1372 (N_1372,In_2328,In_1135);
nand U1373 (N_1373,In_1842,In_1526);
nand U1374 (N_1374,In_613,In_881);
xnor U1375 (N_1375,In_1344,In_77);
nand U1376 (N_1376,In_532,In_2040);
or U1377 (N_1377,In_1677,In_1211);
nor U1378 (N_1378,In_1810,In_1104);
or U1379 (N_1379,In_178,In_1696);
xnor U1380 (N_1380,In_75,In_582);
or U1381 (N_1381,In_1665,In_1811);
and U1382 (N_1382,In_2485,In_14);
and U1383 (N_1383,In_698,In_2132);
and U1384 (N_1384,In_1761,In_1568);
nor U1385 (N_1385,In_1111,In_1287);
or U1386 (N_1386,In_1036,In_1945);
or U1387 (N_1387,In_27,In_1713);
or U1388 (N_1388,In_2001,In_911);
and U1389 (N_1389,In_391,In_330);
xor U1390 (N_1390,In_758,In_73);
and U1391 (N_1391,In_713,In_728);
xnor U1392 (N_1392,In_2099,In_972);
nand U1393 (N_1393,In_2373,In_616);
nor U1394 (N_1394,In_1552,In_586);
nor U1395 (N_1395,In_460,In_1664);
nand U1396 (N_1396,In_2254,In_1741);
nor U1397 (N_1397,In_2346,In_1907);
and U1398 (N_1398,In_2205,In_55);
nand U1399 (N_1399,In_743,In_1224);
and U1400 (N_1400,In_2204,In_707);
nor U1401 (N_1401,In_1547,In_741);
nor U1402 (N_1402,In_934,In_1939);
nor U1403 (N_1403,In_496,In_454);
or U1404 (N_1404,In_1438,In_920);
nand U1405 (N_1405,In_1614,In_6);
and U1406 (N_1406,In_2137,In_332);
and U1407 (N_1407,In_1911,In_2413);
and U1408 (N_1408,In_1362,In_843);
nand U1409 (N_1409,In_362,In_2283);
nand U1410 (N_1410,In_419,In_58);
nor U1411 (N_1411,In_135,In_2283);
nor U1412 (N_1412,In_962,In_1308);
nor U1413 (N_1413,In_610,In_935);
xor U1414 (N_1414,In_1295,In_1010);
or U1415 (N_1415,In_2457,In_326);
and U1416 (N_1416,In_157,In_1262);
and U1417 (N_1417,In_1103,In_593);
or U1418 (N_1418,In_783,In_1448);
and U1419 (N_1419,In_2224,In_1591);
xnor U1420 (N_1420,In_334,In_2087);
nor U1421 (N_1421,In_1378,In_126);
nor U1422 (N_1422,In_1681,In_532);
nor U1423 (N_1423,In_34,In_1397);
xnor U1424 (N_1424,In_83,In_991);
nand U1425 (N_1425,In_1245,In_384);
and U1426 (N_1426,In_1194,In_1203);
nor U1427 (N_1427,In_1479,In_1849);
nor U1428 (N_1428,In_1977,In_1013);
nor U1429 (N_1429,In_764,In_924);
nor U1430 (N_1430,In_355,In_528);
and U1431 (N_1431,In_2129,In_915);
or U1432 (N_1432,In_1628,In_85);
nand U1433 (N_1433,In_1202,In_1489);
nor U1434 (N_1434,In_1869,In_971);
and U1435 (N_1435,In_1114,In_2130);
and U1436 (N_1436,In_817,In_1685);
nor U1437 (N_1437,In_1069,In_2165);
and U1438 (N_1438,In_973,In_2204);
and U1439 (N_1439,In_313,In_1889);
and U1440 (N_1440,In_1363,In_1318);
nand U1441 (N_1441,In_1704,In_2307);
nand U1442 (N_1442,In_613,In_543);
and U1443 (N_1443,In_858,In_2126);
or U1444 (N_1444,In_48,In_1110);
nand U1445 (N_1445,In_1174,In_2364);
nor U1446 (N_1446,In_648,In_1566);
and U1447 (N_1447,In_1947,In_1003);
or U1448 (N_1448,In_1707,In_1295);
or U1449 (N_1449,In_789,In_1037);
and U1450 (N_1450,In_2138,In_283);
and U1451 (N_1451,In_656,In_727);
or U1452 (N_1452,In_485,In_625);
nand U1453 (N_1453,In_1686,In_2227);
nand U1454 (N_1454,In_55,In_68);
nor U1455 (N_1455,In_1020,In_2185);
or U1456 (N_1456,In_2340,In_2233);
or U1457 (N_1457,In_1957,In_1657);
and U1458 (N_1458,In_1909,In_560);
and U1459 (N_1459,In_573,In_819);
and U1460 (N_1460,In_1770,In_1521);
or U1461 (N_1461,In_2183,In_252);
nand U1462 (N_1462,In_1395,In_311);
nor U1463 (N_1463,In_1686,In_1348);
or U1464 (N_1464,In_1551,In_653);
and U1465 (N_1465,In_1715,In_175);
and U1466 (N_1466,In_743,In_1997);
and U1467 (N_1467,In_746,In_639);
and U1468 (N_1468,In_375,In_1748);
nand U1469 (N_1469,In_180,In_654);
or U1470 (N_1470,In_2207,In_1896);
nand U1471 (N_1471,In_764,In_2103);
nor U1472 (N_1472,In_1529,In_1707);
and U1473 (N_1473,In_150,In_1622);
nand U1474 (N_1474,In_1265,In_972);
or U1475 (N_1475,In_951,In_493);
nand U1476 (N_1476,In_1086,In_2116);
nand U1477 (N_1477,In_1448,In_522);
nand U1478 (N_1478,In_2204,In_358);
or U1479 (N_1479,In_2441,In_2335);
and U1480 (N_1480,In_584,In_339);
nor U1481 (N_1481,In_1227,In_2037);
nand U1482 (N_1482,In_1142,In_946);
nand U1483 (N_1483,In_1567,In_2211);
nor U1484 (N_1484,In_104,In_1482);
and U1485 (N_1485,In_1775,In_291);
and U1486 (N_1486,In_775,In_284);
nor U1487 (N_1487,In_2174,In_729);
nor U1488 (N_1488,In_196,In_1581);
nor U1489 (N_1489,In_930,In_2489);
nor U1490 (N_1490,In_2196,In_2350);
nand U1491 (N_1491,In_2102,In_1334);
and U1492 (N_1492,In_273,In_852);
nor U1493 (N_1493,In_313,In_2488);
nor U1494 (N_1494,In_808,In_2170);
nand U1495 (N_1495,In_926,In_1830);
and U1496 (N_1496,In_1335,In_671);
and U1497 (N_1497,In_1506,In_1752);
nand U1498 (N_1498,In_1614,In_1176);
nand U1499 (N_1499,In_1689,In_1452);
nand U1500 (N_1500,In_826,In_775);
and U1501 (N_1501,In_2120,In_337);
or U1502 (N_1502,In_1414,In_1471);
and U1503 (N_1503,In_1985,In_556);
nor U1504 (N_1504,In_318,In_681);
and U1505 (N_1505,In_95,In_59);
nand U1506 (N_1506,In_334,In_1180);
nor U1507 (N_1507,In_1184,In_95);
and U1508 (N_1508,In_157,In_1350);
and U1509 (N_1509,In_1962,In_1378);
nand U1510 (N_1510,In_1474,In_709);
or U1511 (N_1511,In_783,In_84);
or U1512 (N_1512,In_102,In_555);
and U1513 (N_1513,In_2010,In_2257);
nor U1514 (N_1514,In_1719,In_1522);
and U1515 (N_1515,In_2135,In_500);
or U1516 (N_1516,In_931,In_486);
nor U1517 (N_1517,In_1690,In_103);
xnor U1518 (N_1518,In_474,In_56);
nor U1519 (N_1519,In_473,In_562);
nand U1520 (N_1520,In_412,In_935);
or U1521 (N_1521,In_1288,In_1675);
nor U1522 (N_1522,In_2266,In_1673);
nand U1523 (N_1523,In_1647,In_1775);
nor U1524 (N_1524,In_770,In_185);
nand U1525 (N_1525,In_1655,In_1755);
or U1526 (N_1526,In_1284,In_1414);
nand U1527 (N_1527,In_1915,In_1945);
nor U1528 (N_1528,In_1220,In_1148);
or U1529 (N_1529,In_2239,In_1184);
or U1530 (N_1530,In_1799,In_1091);
nand U1531 (N_1531,In_2431,In_2144);
and U1532 (N_1532,In_1366,In_1623);
nor U1533 (N_1533,In_1394,In_1472);
and U1534 (N_1534,In_1951,In_2481);
nor U1535 (N_1535,In_2248,In_1064);
nor U1536 (N_1536,In_461,In_2054);
and U1537 (N_1537,In_101,In_985);
and U1538 (N_1538,In_1271,In_771);
or U1539 (N_1539,In_2241,In_1395);
nand U1540 (N_1540,In_2295,In_855);
nor U1541 (N_1541,In_2210,In_1810);
and U1542 (N_1542,In_937,In_1293);
or U1543 (N_1543,In_1643,In_1761);
and U1544 (N_1544,In_382,In_2336);
nor U1545 (N_1545,In_2012,In_1668);
nand U1546 (N_1546,In_801,In_858);
nor U1547 (N_1547,In_1359,In_900);
nand U1548 (N_1548,In_1660,In_790);
nand U1549 (N_1549,In_2013,In_1465);
and U1550 (N_1550,In_1301,In_317);
and U1551 (N_1551,In_1499,In_545);
and U1552 (N_1552,In_1394,In_52);
or U1553 (N_1553,In_1955,In_1091);
nor U1554 (N_1554,In_610,In_1889);
xnor U1555 (N_1555,In_1101,In_298);
or U1556 (N_1556,In_2022,In_143);
nand U1557 (N_1557,In_31,In_1123);
nor U1558 (N_1558,In_631,In_546);
and U1559 (N_1559,In_2482,In_696);
or U1560 (N_1560,In_1976,In_1158);
or U1561 (N_1561,In_1311,In_1537);
nand U1562 (N_1562,In_2381,In_2261);
xnor U1563 (N_1563,In_2004,In_1798);
and U1564 (N_1564,In_922,In_809);
or U1565 (N_1565,In_1434,In_148);
xnor U1566 (N_1566,In_3,In_1528);
nor U1567 (N_1567,In_66,In_1128);
and U1568 (N_1568,In_1710,In_1075);
and U1569 (N_1569,In_390,In_744);
nand U1570 (N_1570,In_2441,In_2333);
or U1571 (N_1571,In_1363,In_977);
or U1572 (N_1572,In_848,In_799);
or U1573 (N_1573,In_1447,In_1410);
nor U1574 (N_1574,In_1328,In_316);
or U1575 (N_1575,In_1519,In_631);
nor U1576 (N_1576,In_612,In_2097);
or U1577 (N_1577,In_1544,In_383);
and U1578 (N_1578,In_1550,In_1467);
and U1579 (N_1579,In_1500,In_386);
nor U1580 (N_1580,In_937,In_161);
nor U1581 (N_1581,In_1011,In_1796);
and U1582 (N_1582,In_2385,In_497);
and U1583 (N_1583,In_325,In_1087);
nor U1584 (N_1584,In_718,In_109);
nand U1585 (N_1585,In_1898,In_687);
nand U1586 (N_1586,In_386,In_1605);
nand U1587 (N_1587,In_186,In_1162);
and U1588 (N_1588,In_516,In_1555);
nand U1589 (N_1589,In_1067,In_1203);
nor U1590 (N_1590,In_485,In_1258);
and U1591 (N_1591,In_1475,In_1038);
xor U1592 (N_1592,In_2427,In_1900);
nand U1593 (N_1593,In_822,In_174);
nand U1594 (N_1594,In_1488,In_1002);
xor U1595 (N_1595,In_210,In_866);
nand U1596 (N_1596,In_448,In_1553);
nor U1597 (N_1597,In_1430,In_895);
nor U1598 (N_1598,In_671,In_1115);
nand U1599 (N_1599,In_50,In_2404);
or U1600 (N_1600,In_1081,In_58);
nand U1601 (N_1601,In_1400,In_2410);
or U1602 (N_1602,In_1703,In_660);
nor U1603 (N_1603,In_454,In_1083);
nor U1604 (N_1604,In_805,In_676);
nor U1605 (N_1605,In_105,In_855);
nor U1606 (N_1606,In_1420,In_1148);
and U1607 (N_1607,In_2285,In_67);
and U1608 (N_1608,In_827,In_1799);
or U1609 (N_1609,In_2327,In_2103);
or U1610 (N_1610,In_1814,In_1767);
nor U1611 (N_1611,In_1286,In_1683);
and U1612 (N_1612,In_2378,In_2181);
and U1613 (N_1613,In_1436,In_2050);
and U1614 (N_1614,In_335,In_21);
nor U1615 (N_1615,In_515,In_160);
and U1616 (N_1616,In_2451,In_1695);
nor U1617 (N_1617,In_1356,In_2495);
xor U1618 (N_1618,In_1164,In_804);
nor U1619 (N_1619,In_1286,In_466);
nand U1620 (N_1620,In_537,In_1220);
or U1621 (N_1621,In_2193,In_867);
nor U1622 (N_1622,In_1330,In_1177);
nand U1623 (N_1623,In_1810,In_908);
and U1624 (N_1624,In_263,In_765);
nor U1625 (N_1625,In_128,In_755);
or U1626 (N_1626,In_1101,In_2131);
nand U1627 (N_1627,In_1475,In_1981);
or U1628 (N_1628,In_2345,In_1352);
nor U1629 (N_1629,In_116,In_1236);
and U1630 (N_1630,In_1709,In_1815);
and U1631 (N_1631,In_2065,In_1468);
xnor U1632 (N_1632,In_480,In_1075);
nor U1633 (N_1633,In_215,In_702);
nand U1634 (N_1634,In_2178,In_828);
or U1635 (N_1635,In_954,In_1818);
and U1636 (N_1636,In_1337,In_2155);
xnor U1637 (N_1637,In_751,In_512);
and U1638 (N_1638,In_770,In_194);
xor U1639 (N_1639,In_277,In_71);
or U1640 (N_1640,In_692,In_68);
nor U1641 (N_1641,In_757,In_2040);
or U1642 (N_1642,In_1154,In_1647);
nor U1643 (N_1643,In_2206,In_882);
and U1644 (N_1644,In_618,In_1650);
nand U1645 (N_1645,In_2155,In_1916);
nand U1646 (N_1646,In_2022,In_2436);
nor U1647 (N_1647,In_1808,In_684);
and U1648 (N_1648,In_137,In_839);
nand U1649 (N_1649,In_2430,In_398);
and U1650 (N_1650,In_1747,In_1242);
and U1651 (N_1651,In_1953,In_292);
and U1652 (N_1652,In_837,In_1881);
nor U1653 (N_1653,In_705,In_241);
and U1654 (N_1654,In_368,In_153);
and U1655 (N_1655,In_632,In_658);
and U1656 (N_1656,In_1210,In_426);
or U1657 (N_1657,In_1714,In_968);
or U1658 (N_1658,In_1535,In_1611);
and U1659 (N_1659,In_1865,In_2144);
nand U1660 (N_1660,In_174,In_577);
nor U1661 (N_1661,In_2263,In_1360);
nor U1662 (N_1662,In_1670,In_2149);
nand U1663 (N_1663,In_1811,In_1925);
nor U1664 (N_1664,In_778,In_1375);
nand U1665 (N_1665,In_1551,In_1209);
and U1666 (N_1666,In_2104,In_2286);
and U1667 (N_1667,In_848,In_1548);
nand U1668 (N_1668,In_377,In_798);
nand U1669 (N_1669,In_2128,In_252);
nand U1670 (N_1670,In_872,In_2215);
nand U1671 (N_1671,In_1364,In_2347);
nor U1672 (N_1672,In_2059,In_604);
and U1673 (N_1673,In_2059,In_524);
and U1674 (N_1674,In_2347,In_675);
or U1675 (N_1675,In_481,In_496);
nor U1676 (N_1676,In_483,In_1393);
and U1677 (N_1677,In_261,In_1084);
and U1678 (N_1678,In_309,In_629);
or U1679 (N_1679,In_1166,In_455);
nor U1680 (N_1680,In_1572,In_2250);
or U1681 (N_1681,In_206,In_1512);
and U1682 (N_1682,In_1808,In_1088);
nor U1683 (N_1683,In_1104,In_1068);
and U1684 (N_1684,In_1056,In_1597);
or U1685 (N_1685,In_259,In_139);
and U1686 (N_1686,In_766,In_357);
nor U1687 (N_1687,In_730,In_1056);
and U1688 (N_1688,In_1329,In_1481);
xor U1689 (N_1689,In_2144,In_1425);
nor U1690 (N_1690,In_1976,In_2250);
nor U1691 (N_1691,In_591,In_2029);
nor U1692 (N_1692,In_2108,In_2450);
nor U1693 (N_1693,In_1295,In_1082);
and U1694 (N_1694,In_1002,In_1452);
or U1695 (N_1695,In_1739,In_1915);
and U1696 (N_1696,In_2069,In_1460);
nand U1697 (N_1697,In_1453,In_2168);
and U1698 (N_1698,In_4,In_2335);
or U1699 (N_1699,In_1060,In_2139);
nand U1700 (N_1700,In_2315,In_491);
or U1701 (N_1701,In_2283,In_2374);
nor U1702 (N_1702,In_640,In_1276);
and U1703 (N_1703,In_1108,In_2411);
and U1704 (N_1704,In_1666,In_1106);
or U1705 (N_1705,In_1534,In_2327);
nand U1706 (N_1706,In_518,In_667);
nand U1707 (N_1707,In_828,In_929);
and U1708 (N_1708,In_1168,In_501);
or U1709 (N_1709,In_191,In_100);
or U1710 (N_1710,In_1532,In_827);
or U1711 (N_1711,In_14,In_1336);
nand U1712 (N_1712,In_2420,In_283);
and U1713 (N_1713,In_1634,In_1015);
and U1714 (N_1714,In_1093,In_554);
or U1715 (N_1715,In_1703,In_456);
nor U1716 (N_1716,In_2089,In_1234);
nor U1717 (N_1717,In_2164,In_51);
and U1718 (N_1718,In_1908,In_805);
nand U1719 (N_1719,In_1558,In_902);
or U1720 (N_1720,In_1467,In_1966);
nor U1721 (N_1721,In_349,In_1039);
nor U1722 (N_1722,In_1660,In_340);
nand U1723 (N_1723,In_415,In_327);
and U1724 (N_1724,In_1466,In_1739);
or U1725 (N_1725,In_2054,In_2089);
nor U1726 (N_1726,In_540,In_1039);
nand U1727 (N_1727,In_2385,In_1956);
and U1728 (N_1728,In_375,In_2479);
nor U1729 (N_1729,In_525,In_1657);
or U1730 (N_1730,In_2172,In_1488);
and U1731 (N_1731,In_567,In_2299);
and U1732 (N_1732,In_2068,In_1340);
or U1733 (N_1733,In_2101,In_814);
nor U1734 (N_1734,In_429,In_1536);
nor U1735 (N_1735,In_2109,In_843);
and U1736 (N_1736,In_718,In_1566);
nor U1737 (N_1737,In_439,In_1409);
nand U1738 (N_1738,In_219,In_2181);
nand U1739 (N_1739,In_482,In_1413);
or U1740 (N_1740,In_686,In_1145);
nand U1741 (N_1741,In_867,In_1892);
nor U1742 (N_1742,In_1259,In_1099);
nor U1743 (N_1743,In_1052,In_2247);
nor U1744 (N_1744,In_1890,In_239);
and U1745 (N_1745,In_812,In_143);
nor U1746 (N_1746,In_1431,In_1104);
and U1747 (N_1747,In_1386,In_903);
nor U1748 (N_1748,In_626,In_837);
and U1749 (N_1749,In_1241,In_233);
nor U1750 (N_1750,In_883,In_1775);
or U1751 (N_1751,In_1608,In_1075);
nand U1752 (N_1752,In_2135,In_355);
and U1753 (N_1753,In_710,In_1036);
and U1754 (N_1754,In_1060,In_760);
nand U1755 (N_1755,In_218,In_1406);
and U1756 (N_1756,In_1268,In_1106);
or U1757 (N_1757,In_1099,In_2401);
or U1758 (N_1758,In_42,In_1060);
nand U1759 (N_1759,In_2231,In_818);
nor U1760 (N_1760,In_1762,In_1984);
nand U1761 (N_1761,In_76,In_1165);
and U1762 (N_1762,In_1143,In_1330);
or U1763 (N_1763,In_1119,In_621);
and U1764 (N_1764,In_1939,In_697);
and U1765 (N_1765,In_1642,In_1940);
and U1766 (N_1766,In_1496,In_204);
nand U1767 (N_1767,In_1979,In_908);
and U1768 (N_1768,In_2058,In_239);
or U1769 (N_1769,In_1787,In_249);
nand U1770 (N_1770,In_1028,In_115);
or U1771 (N_1771,In_482,In_1572);
and U1772 (N_1772,In_21,In_784);
or U1773 (N_1773,In_2271,In_2258);
nand U1774 (N_1774,In_1532,In_546);
nand U1775 (N_1775,In_2273,In_82);
or U1776 (N_1776,In_2392,In_1497);
and U1777 (N_1777,In_169,In_2150);
xnor U1778 (N_1778,In_1270,In_1444);
nor U1779 (N_1779,In_1484,In_1057);
nor U1780 (N_1780,In_12,In_330);
and U1781 (N_1781,In_652,In_1505);
or U1782 (N_1782,In_1037,In_1556);
or U1783 (N_1783,In_2252,In_836);
and U1784 (N_1784,In_2104,In_506);
nand U1785 (N_1785,In_1520,In_2095);
or U1786 (N_1786,In_2134,In_596);
and U1787 (N_1787,In_268,In_858);
or U1788 (N_1788,In_2251,In_1385);
or U1789 (N_1789,In_264,In_1359);
nand U1790 (N_1790,In_1462,In_1897);
nand U1791 (N_1791,In_1365,In_1791);
or U1792 (N_1792,In_2425,In_2111);
or U1793 (N_1793,In_1446,In_1057);
or U1794 (N_1794,In_374,In_1388);
nand U1795 (N_1795,In_2142,In_1241);
nor U1796 (N_1796,In_855,In_1268);
nand U1797 (N_1797,In_1634,In_851);
nor U1798 (N_1798,In_1055,In_1671);
nand U1799 (N_1799,In_495,In_227);
nor U1800 (N_1800,In_435,In_1659);
or U1801 (N_1801,In_1142,In_860);
or U1802 (N_1802,In_450,In_2173);
or U1803 (N_1803,In_1058,In_168);
and U1804 (N_1804,In_735,In_2208);
or U1805 (N_1805,In_2429,In_243);
xor U1806 (N_1806,In_2013,In_1357);
nand U1807 (N_1807,In_1031,In_2051);
nand U1808 (N_1808,In_650,In_802);
and U1809 (N_1809,In_1867,In_2474);
or U1810 (N_1810,In_1250,In_1808);
nand U1811 (N_1811,In_294,In_345);
and U1812 (N_1812,In_2300,In_1832);
nor U1813 (N_1813,In_1749,In_382);
or U1814 (N_1814,In_459,In_795);
or U1815 (N_1815,In_859,In_980);
or U1816 (N_1816,In_1021,In_574);
or U1817 (N_1817,In_2110,In_1626);
nor U1818 (N_1818,In_2208,In_2112);
and U1819 (N_1819,In_2221,In_1520);
xor U1820 (N_1820,In_2264,In_2396);
or U1821 (N_1821,In_1072,In_1369);
or U1822 (N_1822,In_1480,In_279);
nor U1823 (N_1823,In_2053,In_301);
nand U1824 (N_1824,In_1725,In_1588);
xor U1825 (N_1825,In_1113,In_972);
and U1826 (N_1826,In_2442,In_956);
nor U1827 (N_1827,In_752,In_1156);
nand U1828 (N_1828,In_2249,In_1276);
nand U1829 (N_1829,In_1219,In_156);
nand U1830 (N_1830,In_816,In_247);
nor U1831 (N_1831,In_553,In_1892);
or U1832 (N_1832,In_1449,In_457);
xor U1833 (N_1833,In_2238,In_984);
nand U1834 (N_1834,In_1743,In_417);
or U1835 (N_1835,In_1264,In_1613);
and U1836 (N_1836,In_2148,In_348);
and U1837 (N_1837,In_2437,In_1347);
and U1838 (N_1838,In_1990,In_1887);
nor U1839 (N_1839,In_1075,In_2040);
nand U1840 (N_1840,In_654,In_83);
and U1841 (N_1841,In_1465,In_685);
nand U1842 (N_1842,In_116,In_1848);
nor U1843 (N_1843,In_341,In_134);
and U1844 (N_1844,In_196,In_2082);
and U1845 (N_1845,In_323,In_2418);
nor U1846 (N_1846,In_771,In_313);
and U1847 (N_1847,In_253,In_1310);
and U1848 (N_1848,In_1832,In_1226);
and U1849 (N_1849,In_638,In_1841);
or U1850 (N_1850,In_1903,In_1535);
or U1851 (N_1851,In_2322,In_1329);
nor U1852 (N_1852,In_2399,In_2051);
and U1853 (N_1853,In_1154,In_254);
or U1854 (N_1854,In_43,In_2107);
nor U1855 (N_1855,In_1320,In_2396);
and U1856 (N_1856,In_639,In_179);
nand U1857 (N_1857,In_2431,In_2218);
and U1858 (N_1858,In_530,In_1687);
nand U1859 (N_1859,In_1246,In_1827);
nor U1860 (N_1860,In_2135,In_1050);
nor U1861 (N_1861,In_2450,In_1966);
nand U1862 (N_1862,In_2359,In_494);
or U1863 (N_1863,In_2229,In_1617);
and U1864 (N_1864,In_149,In_1947);
nor U1865 (N_1865,In_1134,In_919);
nor U1866 (N_1866,In_426,In_1758);
xor U1867 (N_1867,In_2272,In_1710);
nand U1868 (N_1868,In_926,In_2337);
nor U1869 (N_1869,In_81,In_145);
and U1870 (N_1870,In_692,In_2478);
or U1871 (N_1871,In_498,In_1841);
or U1872 (N_1872,In_890,In_168);
nor U1873 (N_1873,In_1834,In_471);
and U1874 (N_1874,In_2377,In_977);
xnor U1875 (N_1875,In_117,In_477);
xor U1876 (N_1876,In_810,In_898);
nand U1877 (N_1877,In_293,In_707);
nor U1878 (N_1878,In_1397,In_1885);
nand U1879 (N_1879,In_728,In_161);
nand U1880 (N_1880,In_1313,In_1522);
nor U1881 (N_1881,In_1999,In_341);
or U1882 (N_1882,In_1387,In_435);
nand U1883 (N_1883,In_2288,In_1173);
nor U1884 (N_1884,In_2279,In_2464);
or U1885 (N_1885,In_1167,In_1266);
nor U1886 (N_1886,In_1140,In_1077);
and U1887 (N_1887,In_1272,In_2228);
nor U1888 (N_1888,In_2350,In_1162);
nor U1889 (N_1889,In_584,In_1831);
or U1890 (N_1890,In_1743,In_847);
or U1891 (N_1891,In_1782,In_131);
nand U1892 (N_1892,In_456,In_1010);
nor U1893 (N_1893,In_1083,In_921);
xor U1894 (N_1894,In_1628,In_2100);
and U1895 (N_1895,In_1118,In_1474);
or U1896 (N_1896,In_1013,In_2048);
nor U1897 (N_1897,In_1262,In_2031);
and U1898 (N_1898,In_2408,In_170);
and U1899 (N_1899,In_86,In_874);
or U1900 (N_1900,In_2137,In_227);
or U1901 (N_1901,In_58,In_1937);
nand U1902 (N_1902,In_732,In_1576);
nand U1903 (N_1903,In_1967,In_165);
or U1904 (N_1904,In_2417,In_1804);
nand U1905 (N_1905,In_505,In_2203);
nand U1906 (N_1906,In_1262,In_688);
nand U1907 (N_1907,In_2005,In_1789);
or U1908 (N_1908,In_2174,In_818);
nor U1909 (N_1909,In_1620,In_1957);
nor U1910 (N_1910,In_1835,In_728);
nand U1911 (N_1911,In_1755,In_65);
nand U1912 (N_1912,In_1491,In_1267);
nor U1913 (N_1913,In_663,In_885);
nor U1914 (N_1914,In_1252,In_1067);
nor U1915 (N_1915,In_339,In_106);
nor U1916 (N_1916,In_48,In_2333);
nand U1917 (N_1917,In_1160,In_350);
and U1918 (N_1918,In_584,In_827);
and U1919 (N_1919,In_1299,In_706);
nand U1920 (N_1920,In_1434,In_1682);
and U1921 (N_1921,In_992,In_557);
and U1922 (N_1922,In_1986,In_758);
or U1923 (N_1923,In_548,In_1630);
and U1924 (N_1924,In_734,In_649);
or U1925 (N_1925,In_23,In_375);
nand U1926 (N_1926,In_254,In_1122);
and U1927 (N_1927,In_1751,In_292);
nor U1928 (N_1928,In_2253,In_73);
or U1929 (N_1929,In_641,In_135);
nand U1930 (N_1930,In_256,In_370);
nor U1931 (N_1931,In_1265,In_591);
nand U1932 (N_1932,In_485,In_989);
nand U1933 (N_1933,In_289,In_1332);
nor U1934 (N_1934,In_1200,In_316);
nor U1935 (N_1935,In_2492,In_2117);
and U1936 (N_1936,In_1201,In_381);
nor U1937 (N_1937,In_246,In_2151);
and U1938 (N_1938,In_2366,In_1483);
nor U1939 (N_1939,In_869,In_1798);
or U1940 (N_1940,In_863,In_1130);
and U1941 (N_1941,In_667,In_1960);
nor U1942 (N_1942,In_2342,In_2234);
nand U1943 (N_1943,In_1794,In_221);
and U1944 (N_1944,In_1789,In_2227);
and U1945 (N_1945,In_2155,In_1693);
nand U1946 (N_1946,In_873,In_1180);
nand U1947 (N_1947,In_2435,In_1992);
or U1948 (N_1948,In_1071,In_474);
and U1949 (N_1949,In_166,In_1439);
nand U1950 (N_1950,In_983,In_2280);
nor U1951 (N_1951,In_1922,In_2251);
and U1952 (N_1952,In_953,In_1882);
or U1953 (N_1953,In_1294,In_709);
xnor U1954 (N_1954,In_14,In_1128);
nand U1955 (N_1955,In_2337,In_106);
nor U1956 (N_1956,In_1112,In_8);
and U1957 (N_1957,In_2218,In_555);
and U1958 (N_1958,In_1916,In_2370);
and U1959 (N_1959,In_2261,In_861);
nand U1960 (N_1960,In_2316,In_2399);
nor U1961 (N_1961,In_1691,In_1226);
and U1962 (N_1962,In_467,In_799);
nand U1963 (N_1963,In_1103,In_664);
and U1964 (N_1964,In_1424,In_265);
nand U1965 (N_1965,In_1463,In_569);
nand U1966 (N_1966,In_1323,In_1495);
nand U1967 (N_1967,In_2399,In_1404);
nor U1968 (N_1968,In_267,In_1415);
and U1969 (N_1969,In_1209,In_2430);
or U1970 (N_1970,In_746,In_514);
and U1971 (N_1971,In_1334,In_1988);
or U1972 (N_1972,In_981,In_1131);
nand U1973 (N_1973,In_1658,In_263);
nor U1974 (N_1974,In_1715,In_888);
and U1975 (N_1975,In_2029,In_1802);
nand U1976 (N_1976,In_375,In_1952);
xnor U1977 (N_1977,In_144,In_536);
nand U1978 (N_1978,In_618,In_2291);
nor U1979 (N_1979,In_1041,In_343);
nor U1980 (N_1980,In_1011,In_1130);
and U1981 (N_1981,In_1891,In_1965);
nor U1982 (N_1982,In_1223,In_920);
nor U1983 (N_1983,In_1499,In_846);
or U1984 (N_1984,In_1896,In_586);
nor U1985 (N_1985,In_1810,In_420);
nor U1986 (N_1986,In_2434,In_1234);
or U1987 (N_1987,In_1654,In_2094);
and U1988 (N_1988,In_2332,In_2440);
nand U1989 (N_1989,In_2131,In_1095);
nand U1990 (N_1990,In_1378,In_1759);
or U1991 (N_1991,In_1299,In_931);
nand U1992 (N_1992,In_728,In_2220);
nand U1993 (N_1993,In_1672,In_1004);
and U1994 (N_1994,In_2103,In_1744);
and U1995 (N_1995,In_94,In_2086);
and U1996 (N_1996,In_596,In_900);
nor U1997 (N_1997,In_1306,In_1884);
nand U1998 (N_1998,In_1016,In_615);
or U1999 (N_1999,In_395,In_1265);
nor U2000 (N_2000,In_2428,In_1204);
nor U2001 (N_2001,In_562,In_1562);
nor U2002 (N_2002,In_1599,In_1950);
or U2003 (N_2003,In_834,In_1876);
and U2004 (N_2004,In_1988,In_2349);
nand U2005 (N_2005,In_128,In_152);
or U2006 (N_2006,In_141,In_1457);
nand U2007 (N_2007,In_303,In_460);
and U2008 (N_2008,In_1344,In_587);
nor U2009 (N_2009,In_961,In_1768);
or U2010 (N_2010,In_64,In_98);
and U2011 (N_2011,In_849,In_2282);
and U2012 (N_2012,In_457,In_1896);
nor U2013 (N_2013,In_306,In_731);
and U2014 (N_2014,In_1597,In_1836);
and U2015 (N_2015,In_784,In_2233);
nor U2016 (N_2016,In_1591,In_1720);
nor U2017 (N_2017,In_952,In_47);
xnor U2018 (N_2018,In_1296,In_351);
and U2019 (N_2019,In_2431,In_1854);
and U2020 (N_2020,In_2361,In_1662);
and U2021 (N_2021,In_188,In_1371);
or U2022 (N_2022,In_1626,In_962);
nor U2023 (N_2023,In_1584,In_2187);
and U2024 (N_2024,In_1814,In_1522);
nand U2025 (N_2025,In_610,In_711);
and U2026 (N_2026,In_713,In_1176);
nand U2027 (N_2027,In_2125,In_1744);
and U2028 (N_2028,In_2004,In_1290);
nor U2029 (N_2029,In_2124,In_1975);
or U2030 (N_2030,In_1138,In_839);
or U2031 (N_2031,In_1610,In_152);
nand U2032 (N_2032,In_179,In_636);
nand U2033 (N_2033,In_1280,In_437);
nand U2034 (N_2034,In_2372,In_381);
and U2035 (N_2035,In_279,In_939);
and U2036 (N_2036,In_1364,In_1304);
and U2037 (N_2037,In_1499,In_705);
nor U2038 (N_2038,In_1206,In_1575);
nand U2039 (N_2039,In_715,In_506);
or U2040 (N_2040,In_1345,In_1424);
or U2041 (N_2041,In_220,In_1364);
or U2042 (N_2042,In_1264,In_1603);
and U2043 (N_2043,In_1874,In_862);
or U2044 (N_2044,In_2301,In_1475);
or U2045 (N_2045,In_431,In_843);
nor U2046 (N_2046,In_545,In_1466);
nor U2047 (N_2047,In_1851,In_508);
and U2048 (N_2048,In_2159,In_1193);
nand U2049 (N_2049,In_1500,In_899);
nor U2050 (N_2050,In_935,In_607);
and U2051 (N_2051,In_1919,In_1544);
or U2052 (N_2052,In_206,In_226);
and U2053 (N_2053,In_1527,In_2483);
nor U2054 (N_2054,In_889,In_1932);
nor U2055 (N_2055,In_1744,In_2315);
nand U2056 (N_2056,In_1060,In_2309);
and U2057 (N_2057,In_1390,In_2381);
nor U2058 (N_2058,In_1922,In_2286);
nor U2059 (N_2059,In_2485,In_2113);
nor U2060 (N_2060,In_2025,In_1566);
nor U2061 (N_2061,In_344,In_688);
or U2062 (N_2062,In_2379,In_1923);
nor U2063 (N_2063,In_913,In_2075);
nand U2064 (N_2064,In_2354,In_2147);
or U2065 (N_2065,In_2280,In_746);
and U2066 (N_2066,In_1837,In_973);
or U2067 (N_2067,In_1306,In_1400);
or U2068 (N_2068,In_218,In_1350);
xor U2069 (N_2069,In_409,In_935);
and U2070 (N_2070,In_1697,In_1964);
nor U2071 (N_2071,In_1283,In_1850);
nand U2072 (N_2072,In_1877,In_375);
and U2073 (N_2073,In_2274,In_290);
or U2074 (N_2074,In_486,In_560);
or U2075 (N_2075,In_2111,In_2008);
or U2076 (N_2076,In_1678,In_625);
or U2077 (N_2077,In_800,In_1334);
nor U2078 (N_2078,In_2186,In_349);
and U2079 (N_2079,In_1135,In_498);
or U2080 (N_2080,In_655,In_648);
nor U2081 (N_2081,In_104,In_1566);
or U2082 (N_2082,In_301,In_1319);
or U2083 (N_2083,In_2257,In_1197);
or U2084 (N_2084,In_1169,In_25);
or U2085 (N_2085,In_2095,In_2078);
and U2086 (N_2086,In_2399,In_1100);
nor U2087 (N_2087,In_2375,In_2279);
and U2088 (N_2088,In_59,In_1985);
or U2089 (N_2089,In_525,In_415);
nor U2090 (N_2090,In_184,In_3);
nor U2091 (N_2091,In_175,In_2387);
nor U2092 (N_2092,In_1430,In_355);
and U2093 (N_2093,In_2112,In_2155);
nand U2094 (N_2094,In_2256,In_927);
nor U2095 (N_2095,In_407,In_504);
and U2096 (N_2096,In_227,In_147);
or U2097 (N_2097,In_1374,In_1460);
or U2098 (N_2098,In_1424,In_1668);
and U2099 (N_2099,In_453,In_883);
nor U2100 (N_2100,In_2086,In_1959);
nor U2101 (N_2101,In_259,In_1019);
and U2102 (N_2102,In_1368,In_733);
or U2103 (N_2103,In_2394,In_711);
xor U2104 (N_2104,In_1269,In_563);
nor U2105 (N_2105,In_958,In_686);
or U2106 (N_2106,In_1544,In_2196);
nand U2107 (N_2107,In_2126,In_1777);
or U2108 (N_2108,In_1006,In_1140);
or U2109 (N_2109,In_41,In_1363);
nand U2110 (N_2110,In_2484,In_764);
and U2111 (N_2111,In_901,In_2143);
or U2112 (N_2112,In_1924,In_795);
and U2113 (N_2113,In_12,In_1449);
nand U2114 (N_2114,In_1695,In_2082);
and U2115 (N_2115,In_1184,In_1858);
or U2116 (N_2116,In_559,In_1162);
and U2117 (N_2117,In_1642,In_1116);
nand U2118 (N_2118,In_1202,In_1453);
nor U2119 (N_2119,In_2004,In_2230);
nand U2120 (N_2120,In_1210,In_1660);
and U2121 (N_2121,In_1890,In_1793);
nand U2122 (N_2122,In_496,In_2130);
nand U2123 (N_2123,In_1266,In_1832);
nand U2124 (N_2124,In_288,In_1079);
or U2125 (N_2125,In_715,In_2269);
and U2126 (N_2126,In_1990,In_1135);
nor U2127 (N_2127,In_604,In_383);
or U2128 (N_2128,In_1869,In_864);
nor U2129 (N_2129,In_2061,In_1998);
nand U2130 (N_2130,In_1276,In_905);
and U2131 (N_2131,In_1352,In_1681);
or U2132 (N_2132,In_1763,In_1125);
nand U2133 (N_2133,In_2227,In_2367);
and U2134 (N_2134,In_1436,In_2005);
or U2135 (N_2135,In_898,In_53);
nor U2136 (N_2136,In_1183,In_673);
nor U2137 (N_2137,In_1178,In_745);
and U2138 (N_2138,In_2052,In_978);
nor U2139 (N_2139,In_62,In_733);
or U2140 (N_2140,In_728,In_111);
nor U2141 (N_2141,In_525,In_1274);
nand U2142 (N_2142,In_1690,In_883);
or U2143 (N_2143,In_170,In_1734);
and U2144 (N_2144,In_1614,In_1833);
or U2145 (N_2145,In_439,In_328);
and U2146 (N_2146,In_1593,In_621);
nor U2147 (N_2147,In_631,In_90);
and U2148 (N_2148,In_1019,In_1214);
xor U2149 (N_2149,In_1006,In_1363);
nor U2150 (N_2150,In_2308,In_460);
nand U2151 (N_2151,In_2269,In_1444);
and U2152 (N_2152,In_998,In_263);
nand U2153 (N_2153,In_352,In_1858);
or U2154 (N_2154,In_1706,In_1315);
nand U2155 (N_2155,In_1788,In_2004);
nand U2156 (N_2156,In_682,In_770);
or U2157 (N_2157,In_1927,In_381);
or U2158 (N_2158,In_183,In_1470);
and U2159 (N_2159,In_535,In_461);
and U2160 (N_2160,In_2144,In_2180);
or U2161 (N_2161,In_1472,In_355);
or U2162 (N_2162,In_1746,In_2414);
nand U2163 (N_2163,In_1001,In_2013);
and U2164 (N_2164,In_2285,In_2089);
and U2165 (N_2165,In_1554,In_1152);
nand U2166 (N_2166,In_1914,In_734);
or U2167 (N_2167,In_382,In_222);
and U2168 (N_2168,In_2077,In_1933);
or U2169 (N_2169,In_2308,In_1130);
xnor U2170 (N_2170,In_2007,In_1872);
and U2171 (N_2171,In_610,In_1848);
nand U2172 (N_2172,In_1507,In_645);
or U2173 (N_2173,In_219,In_254);
nor U2174 (N_2174,In_1892,In_1905);
nor U2175 (N_2175,In_1056,In_762);
nor U2176 (N_2176,In_2379,In_477);
nor U2177 (N_2177,In_178,In_315);
and U2178 (N_2178,In_547,In_2151);
nor U2179 (N_2179,In_914,In_237);
or U2180 (N_2180,In_1415,In_761);
and U2181 (N_2181,In_54,In_1108);
nand U2182 (N_2182,In_2288,In_1436);
nand U2183 (N_2183,In_1007,In_2303);
nand U2184 (N_2184,In_1933,In_2379);
nor U2185 (N_2185,In_901,In_1734);
or U2186 (N_2186,In_1066,In_1826);
or U2187 (N_2187,In_513,In_1478);
and U2188 (N_2188,In_1605,In_2281);
nand U2189 (N_2189,In_220,In_1313);
or U2190 (N_2190,In_1170,In_701);
nand U2191 (N_2191,In_1491,In_1439);
or U2192 (N_2192,In_2257,In_2240);
or U2193 (N_2193,In_90,In_532);
nor U2194 (N_2194,In_1166,In_1982);
nor U2195 (N_2195,In_1695,In_2207);
nor U2196 (N_2196,In_438,In_2194);
and U2197 (N_2197,In_1589,In_1024);
and U2198 (N_2198,In_1467,In_780);
nor U2199 (N_2199,In_1291,In_743);
nand U2200 (N_2200,In_799,In_1137);
and U2201 (N_2201,In_1843,In_824);
and U2202 (N_2202,In_2263,In_2276);
and U2203 (N_2203,In_1068,In_1288);
or U2204 (N_2204,In_550,In_301);
nor U2205 (N_2205,In_930,In_2219);
nand U2206 (N_2206,In_78,In_1745);
and U2207 (N_2207,In_2114,In_1617);
nor U2208 (N_2208,In_2418,In_654);
nand U2209 (N_2209,In_2212,In_2026);
and U2210 (N_2210,In_862,In_516);
or U2211 (N_2211,In_407,In_1280);
or U2212 (N_2212,In_90,In_1816);
nor U2213 (N_2213,In_1020,In_1665);
or U2214 (N_2214,In_2324,In_1569);
nand U2215 (N_2215,In_286,In_2403);
or U2216 (N_2216,In_2460,In_240);
and U2217 (N_2217,In_1897,In_317);
and U2218 (N_2218,In_939,In_1682);
nand U2219 (N_2219,In_304,In_1063);
or U2220 (N_2220,In_838,In_204);
xnor U2221 (N_2221,In_302,In_1351);
or U2222 (N_2222,In_2322,In_827);
nor U2223 (N_2223,In_2397,In_2353);
or U2224 (N_2224,In_2251,In_1205);
nor U2225 (N_2225,In_1729,In_1581);
nor U2226 (N_2226,In_173,In_784);
nand U2227 (N_2227,In_917,In_1572);
nor U2228 (N_2228,In_1251,In_2311);
nor U2229 (N_2229,In_774,In_931);
or U2230 (N_2230,In_980,In_2238);
or U2231 (N_2231,In_25,In_1180);
and U2232 (N_2232,In_2225,In_2111);
or U2233 (N_2233,In_38,In_275);
or U2234 (N_2234,In_2003,In_1001);
nor U2235 (N_2235,In_2090,In_269);
or U2236 (N_2236,In_2164,In_2128);
nand U2237 (N_2237,In_1681,In_1123);
and U2238 (N_2238,In_2201,In_140);
nor U2239 (N_2239,In_2388,In_1368);
nor U2240 (N_2240,In_1902,In_1873);
xnor U2241 (N_2241,In_1117,In_1823);
nand U2242 (N_2242,In_2181,In_1620);
nand U2243 (N_2243,In_895,In_1519);
nor U2244 (N_2244,In_1789,In_2182);
and U2245 (N_2245,In_73,In_2194);
nand U2246 (N_2246,In_782,In_7);
nand U2247 (N_2247,In_364,In_828);
nand U2248 (N_2248,In_696,In_539);
or U2249 (N_2249,In_1040,In_2119);
nand U2250 (N_2250,In_22,In_862);
or U2251 (N_2251,In_2443,In_489);
or U2252 (N_2252,In_14,In_2352);
or U2253 (N_2253,In_1102,In_141);
and U2254 (N_2254,In_525,In_1627);
nor U2255 (N_2255,In_1960,In_328);
nand U2256 (N_2256,In_2439,In_2058);
nand U2257 (N_2257,In_952,In_546);
nand U2258 (N_2258,In_1271,In_31);
or U2259 (N_2259,In_424,In_2357);
nand U2260 (N_2260,In_1743,In_644);
or U2261 (N_2261,In_301,In_1244);
nor U2262 (N_2262,In_1854,In_2283);
or U2263 (N_2263,In_2488,In_929);
nor U2264 (N_2264,In_317,In_1129);
nor U2265 (N_2265,In_764,In_86);
and U2266 (N_2266,In_1911,In_519);
nor U2267 (N_2267,In_2246,In_1161);
or U2268 (N_2268,In_2090,In_1891);
nand U2269 (N_2269,In_2441,In_2196);
nand U2270 (N_2270,In_2394,In_523);
nor U2271 (N_2271,In_2435,In_1767);
and U2272 (N_2272,In_1528,In_1393);
nand U2273 (N_2273,In_96,In_1595);
and U2274 (N_2274,In_2048,In_889);
nor U2275 (N_2275,In_1405,In_134);
nor U2276 (N_2276,In_34,In_351);
nand U2277 (N_2277,In_249,In_2130);
xnor U2278 (N_2278,In_1844,In_156);
xor U2279 (N_2279,In_2490,In_1632);
nand U2280 (N_2280,In_1432,In_1446);
nand U2281 (N_2281,In_1045,In_143);
or U2282 (N_2282,In_1647,In_1146);
and U2283 (N_2283,In_195,In_2299);
or U2284 (N_2284,In_1102,In_2123);
and U2285 (N_2285,In_2333,In_594);
nor U2286 (N_2286,In_911,In_499);
nor U2287 (N_2287,In_904,In_1140);
or U2288 (N_2288,In_567,In_2117);
nor U2289 (N_2289,In_591,In_2426);
nand U2290 (N_2290,In_345,In_2139);
or U2291 (N_2291,In_995,In_1298);
nor U2292 (N_2292,In_1855,In_1178);
nor U2293 (N_2293,In_1009,In_2236);
nand U2294 (N_2294,In_1724,In_1061);
nor U2295 (N_2295,In_556,In_1534);
and U2296 (N_2296,In_1647,In_571);
and U2297 (N_2297,In_2229,In_306);
nand U2298 (N_2298,In_918,In_1834);
nand U2299 (N_2299,In_785,In_835);
and U2300 (N_2300,In_1007,In_1016);
and U2301 (N_2301,In_315,In_1795);
and U2302 (N_2302,In_2157,In_821);
or U2303 (N_2303,In_1573,In_1404);
nor U2304 (N_2304,In_1721,In_746);
and U2305 (N_2305,In_1429,In_2063);
xnor U2306 (N_2306,In_931,In_221);
or U2307 (N_2307,In_164,In_1547);
nand U2308 (N_2308,In_2402,In_1846);
or U2309 (N_2309,In_1802,In_1758);
and U2310 (N_2310,In_1802,In_1578);
nor U2311 (N_2311,In_1297,In_2479);
nor U2312 (N_2312,In_1049,In_313);
or U2313 (N_2313,In_482,In_538);
and U2314 (N_2314,In_125,In_1931);
or U2315 (N_2315,In_841,In_112);
or U2316 (N_2316,In_2069,In_762);
or U2317 (N_2317,In_2406,In_2441);
xor U2318 (N_2318,In_2243,In_683);
nand U2319 (N_2319,In_1518,In_1058);
nor U2320 (N_2320,In_2275,In_1433);
nor U2321 (N_2321,In_1060,In_1603);
nand U2322 (N_2322,In_215,In_1649);
nand U2323 (N_2323,In_378,In_1762);
and U2324 (N_2324,In_97,In_1323);
nand U2325 (N_2325,In_933,In_1101);
and U2326 (N_2326,In_1825,In_2089);
or U2327 (N_2327,In_917,In_426);
nor U2328 (N_2328,In_1010,In_2486);
nor U2329 (N_2329,In_709,In_2201);
or U2330 (N_2330,In_1745,In_2171);
or U2331 (N_2331,In_1112,In_1330);
nor U2332 (N_2332,In_1769,In_846);
nand U2333 (N_2333,In_210,In_2132);
nand U2334 (N_2334,In_710,In_958);
nor U2335 (N_2335,In_893,In_284);
nor U2336 (N_2336,In_1958,In_579);
and U2337 (N_2337,In_341,In_1049);
nor U2338 (N_2338,In_1521,In_235);
and U2339 (N_2339,In_94,In_974);
nor U2340 (N_2340,In_2057,In_2186);
nand U2341 (N_2341,In_116,In_2300);
nand U2342 (N_2342,In_340,In_2015);
and U2343 (N_2343,In_570,In_590);
or U2344 (N_2344,In_9,In_1887);
nand U2345 (N_2345,In_1836,In_9);
nand U2346 (N_2346,In_990,In_2403);
nor U2347 (N_2347,In_678,In_474);
or U2348 (N_2348,In_141,In_155);
nor U2349 (N_2349,In_994,In_651);
xor U2350 (N_2350,In_2228,In_670);
nand U2351 (N_2351,In_1705,In_22);
nand U2352 (N_2352,In_1034,In_97);
or U2353 (N_2353,In_389,In_688);
and U2354 (N_2354,In_1647,In_1580);
xnor U2355 (N_2355,In_1711,In_2298);
nand U2356 (N_2356,In_2262,In_526);
xor U2357 (N_2357,In_1597,In_2449);
and U2358 (N_2358,In_514,In_1396);
and U2359 (N_2359,In_1898,In_1351);
or U2360 (N_2360,In_1051,In_1340);
nand U2361 (N_2361,In_951,In_664);
nand U2362 (N_2362,In_27,In_1632);
xor U2363 (N_2363,In_1528,In_365);
or U2364 (N_2364,In_237,In_1521);
or U2365 (N_2365,In_602,In_2198);
nor U2366 (N_2366,In_1567,In_2495);
or U2367 (N_2367,In_644,In_2287);
or U2368 (N_2368,In_1366,In_80);
nand U2369 (N_2369,In_305,In_671);
and U2370 (N_2370,In_1267,In_2229);
or U2371 (N_2371,In_706,In_127);
or U2372 (N_2372,In_612,In_817);
and U2373 (N_2373,In_405,In_1865);
or U2374 (N_2374,In_1003,In_2378);
or U2375 (N_2375,In_951,In_1950);
or U2376 (N_2376,In_2399,In_10);
or U2377 (N_2377,In_58,In_1643);
or U2378 (N_2378,In_1559,In_604);
nor U2379 (N_2379,In_1067,In_903);
nor U2380 (N_2380,In_1876,In_603);
nand U2381 (N_2381,In_801,In_1059);
or U2382 (N_2382,In_869,In_805);
nand U2383 (N_2383,In_628,In_2171);
nor U2384 (N_2384,In_1956,In_2163);
and U2385 (N_2385,In_2474,In_1099);
nor U2386 (N_2386,In_2460,In_869);
xor U2387 (N_2387,In_1806,In_88);
and U2388 (N_2388,In_231,In_1221);
xnor U2389 (N_2389,In_2219,In_411);
nor U2390 (N_2390,In_1316,In_1674);
nand U2391 (N_2391,In_613,In_1198);
or U2392 (N_2392,In_530,In_475);
nor U2393 (N_2393,In_2023,In_1939);
and U2394 (N_2394,In_98,In_104);
nand U2395 (N_2395,In_2205,In_897);
nand U2396 (N_2396,In_1488,In_530);
nor U2397 (N_2397,In_1680,In_872);
and U2398 (N_2398,In_174,In_667);
or U2399 (N_2399,In_846,In_2284);
nand U2400 (N_2400,In_933,In_1264);
or U2401 (N_2401,In_835,In_2393);
and U2402 (N_2402,In_352,In_1014);
nor U2403 (N_2403,In_338,In_1346);
and U2404 (N_2404,In_1864,In_1756);
or U2405 (N_2405,In_1451,In_2155);
nor U2406 (N_2406,In_1308,In_797);
and U2407 (N_2407,In_1546,In_765);
or U2408 (N_2408,In_2173,In_1192);
or U2409 (N_2409,In_1215,In_2461);
or U2410 (N_2410,In_1339,In_81);
nand U2411 (N_2411,In_427,In_1208);
nor U2412 (N_2412,In_1918,In_76);
nand U2413 (N_2413,In_2006,In_816);
and U2414 (N_2414,In_1420,In_1223);
or U2415 (N_2415,In_2234,In_2110);
xnor U2416 (N_2416,In_108,In_358);
nand U2417 (N_2417,In_1353,In_227);
xnor U2418 (N_2418,In_1176,In_2190);
nor U2419 (N_2419,In_2088,In_1446);
nand U2420 (N_2420,In_1080,In_2043);
and U2421 (N_2421,In_1402,In_1675);
and U2422 (N_2422,In_286,In_842);
or U2423 (N_2423,In_1597,In_1066);
nor U2424 (N_2424,In_157,In_364);
nand U2425 (N_2425,In_609,In_249);
or U2426 (N_2426,In_1548,In_103);
and U2427 (N_2427,In_138,In_1530);
nand U2428 (N_2428,In_967,In_590);
nand U2429 (N_2429,In_1111,In_324);
xnor U2430 (N_2430,In_2446,In_237);
nor U2431 (N_2431,In_2221,In_1976);
nor U2432 (N_2432,In_1901,In_915);
nor U2433 (N_2433,In_1557,In_2459);
and U2434 (N_2434,In_732,In_809);
nand U2435 (N_2435,In_324,In_1250);
nor U2436 (N_2436,In_185,In_432);
or U2437 (N_2437,In_261,In_2132);
or U2438 (N_2438,In_412,In_1237);
nor U2439 (N_2439,In_684,In_1822);
or U2440 (N_2440,In_1809,In_1218);
and U2441 (N_2441,In_1600,In_1456);
nand U2442 (N_2442,In_1065,In_1870);
nand U2443 (N_2443,In_2395,In_802);
nand U2444 (N_2444,In_78,In_1809);
or U2445 (N_2445,In_1470,In_1266);
and U2446 (N_2446,In_974,In_576);
nor U2447 (N_2447,In_1254,In_703);
and U2448 (N_2448,In_1095,In_129);
nand U2449 (N_2449,In_757,In_1543);
and U2450 (N_2450,In_805,In_1225);
nor U2451 (N_2451,In_1124,In_1886);
and U2452 (N_2452,In_980,In_1287);
xor U2453 (N_2453,In_1544,In_2224);
nand U2454 (N_2454,In_2335,In_161);
or U2455 (N_2455,In_1288,In_1626);
nor U2456 (N_2456,In_1374,In_1299);
or U2457 (N_2457,In_1479,In_688);
or U2458 (N_2458,In_2192,In_1393);
nor U2459 (N_2459,In_1040,In_1493);
and U2460 (N_2460,In_225,In_1437);
or U2461 (N_2461,In_341,In_1323);
or U2462 (N_2462,In_2299,In_1249);
or U2463 (N_2463,In_1067,In_1278);
or U2464 (N_2464,In_2067,In_2312);
nand U2465 (N_2465,In_2203,In_2340);
nor U2466 (N_2466,In_1947,In_2060);
nand U2467 (N_2467,In_1837,In_291);
and U2468 (N_2468,In_1793,In_1817);
and U2469 (N_2469,In_1590,In_1689);
and U2470 (N_2470,In_715,In_254);
xnor U2471 (N_2471,In_1864,In_836);
and U2472 (N_2472,In_1514,In_424);
nand U2473 (N_2473,In_1512,In_1436);
nand U2474 (N_2474,In_919,In_1922);
and U2475 (N_2475,In_2421,In_879);
xnor U2476 (N_2476,In_554,In_1484);
or U2477 (N_2477,In_1662,In_739);
nand U2478 (N_2478,In_2062,In_228);
or U2479 (N_2479,In_1841,In_1831);
nor U2480 (N_2480,In_2028,In_573);
and U2481 (N_2481,In_2405,In_2190);
xnor U2482 (N_2482,In_31,In_643);
nor U2483 (N_2483,In_2399,In_646);
nand U2484 (N_2484,In_1609,In_1457);
nand U2485 (N_2485,In_971,In_220);
and U2486 (N_2486,In_1986,In_1724);
nor U2487 (N_2487,In_223,In_1209);
or U2488 (N_2488,In_954,In_1672);
or U2489 (N_2489,In_1658,In_2370);
nor U2490 (N_2490,In_2489,In_1959);
nor U2491 (N_2491,In_856,In_1700);
xnor U2492 (N_2492,In_1965,In_1932);
and U2493 (N_2493,In_607,In_1965);
and U2494 (N_2494,In_1035,In_1589);
or U2495 (N_2495,In_1461,In_2312);
and U2496 (N_2496,In_1029,In_1126);
nand U2497 (N_2497,In_748,In_396);
nor U2498 (N_2498,In_1922,In_627);
nand U2499 (N_2499,In_2463,In_407);
nand U2500 (N_2500,N_1283,N_104);
or U2501 (N_2501,N_521,N_1452);
and U2502 (N_2502,N_1091,N_1641);
xnor U2503 (N_2503,N_1726,N_998);
or U2504 (N_2504,N_2067,N_2143);
and U2505 (N_2505,N_60,N_2017);
and U2506 (N_2506,N_1660,N_1623);
nand U2507 (N_2507,N_562,N_1097);
nor U2508 (N_2508,N_2379,N_668);
or U2509 (N_2509,N_428,N_1948);
nand U2510 (N_2510,N_1177,N_1650);
nor U2511 (N_2511,N_673,N_1043);
nor U2512 (N_2512,N_1227,N_2223);
xnor U2513 (N_2513,N_553,N_651);
and U2514 (N_2514,N_1932,N_1632);
nor U2515 (N_2515,N_638,N_692);
nand U2516 (N_2516,N_603,N_1147);
nand U2517 (N_2517,N_1699,N_2176);
nand U2518 (N_2518,N_1139,N_504);
and U2519 (N_2519,N_2162,N_1661);
nand U2520 (N_2520,N_2027,N_2006);
nand U2521 (N_2521,N_759,N_279);
nor U2522 (N_2522,N_415,N_1507);
and U2523 (N_2523,N_302,N_169);
or U2524 (N_2524,N_1930,N_462);
and U2525 (N_2525,N_377,N_1820);
or U2526 (N_2526,N_807,N_1517);
nor U2527 (N_2527,N_1908,N_1395);
or U2528 (N_2528,N_316,N_2383);
nor U2529 (N_2529,N_1612,N_1727);
or U2530 (N_2530,N_2330,N_137);
xnor U2531 (N_2531,N_448,N_1947);
and U2532 (N_2532,N_992,N_724);
or U2533 (N_2533,N_1827,N_982);
nand U2534 (N_2534,N_480,N_980);
nand U2535 (N_2535,N_1459,N_669);
or U2536 (N_2536,N_1071,N_2008);
and U2537 (N_2537,N_2018,N_787);
and U2538 (N_2538,N_825,N_1214);
or U2539 (N_2539,N_2249,N_2);
nand U2540 (N_2540,N_901,N_2253);
or U2541 (N_2541,N_664,N_2174);
nor U2542 (N_2542,N_867,N_1281);
nand U2543 (N_2543,N_2054,N_1552);
and U2544 (N_2544,N_461,N_177);
nor U2545 (N_2545,N_1870,N_1659);
or U2546 (N_2546,N_1473,N_1925);
and U2547 (N_2547,N_290,N_347);
xnor U2548 (N_2548,N_1157,N_1083);
and U2549 (N_2549,N_1423,N_146);
and U2550 (N_2550,N_1942,N_2228);
and U2551 (N_2551,N_1633,N_2127);
and U2552 (N_2552,N_626,N_554);
or U2553 (N_2553,N_326,N_2108);
or U2554 (N_2554,N_624,N_1330);
and U2555 (N_2555,N_178,N_612);
nand U2556 (N_2556,N_1701,N_129);
nor U2557 (N_2557,N_1263,N_1831);
and U2558 (N_2558,N_667,N_878);
or U2559 (N_2559,N_1983,N_161);
or U2560 (N_2560,N_372,N_911);
and U2561 (N_2561,N_21,N_2132);
xor U2562 (N_2562,N_1367,N_1357);
and U2563 (N_2563,N_792,N_1738);
xor U2564 (N_2564,N_1314,N_307);
nand U2565 (N_2565,N_418,N_446);
or U2566 (N_2566,N_2191,N_709);
nor U2567 (N_2567,N_454,N_1736);
and U2568 (N_2568,N_56,N_1915);
xor U2569 (N_2569,N_2110,N_1411);
and U2570 (N_2570,N_955,N_305);
nor U2571 (N_2571,N_2063,N_1079);
or U2572 (N_2572,N_2263,N_165);
nand U2573 (N_2573,N_103,N_2112);
nor U2574 (N_2574,N_747,N_1592);
and U2575 (N_2575,N_2277,N_826);
nand U2576 (N_2576,N_1107,N_1654);
and U2577 (N_2577,N_239,N_2157);
or U2578 (N_2578,N_989,N_2393);
or U2579 (N_2579,N_2084,N_647);
and U2580 (N_2580,N_493,N_1628);
nor U2581 (N_2581,N_1687,N_170);
or U2582 (N_2582,N_384,N_64);
or U2583 (N_2583,N_730,N_318);
and U2584 (N_2584,N_1640,N_1418);
nor U2585 (N_2585,N_35,N_863);
or U2586 (N_2586,N_606,N_1880);
and U2587 (N_2587,N_1321,N_996);
nand U2588 (N_2588,N_1643,N_1457);
or U2589 (N_2589,N_2152,N_2270);
or U2590 (N_2590,N_4,N_923);
nand U2591 (N_2591,N_868,N_1233);
nor U2592 (N_2592,N_1444,N_650);
xnor U2593 (N_2593,N_840,N_1519);
xnor U2594 (N_2594,N_597,N_2012);
nor U2595 (N_2595,N_1994,N_2248);
nand U2596 (N_2596,N_2107,N_78);
or U2597 (N_2597,N_885,N_544);
or U2598 (N_2598,N_2398,N_166);
nand U2599 (N_2599,N_958,N_528);
nor U2600 (N_2600,N_1226,N_1340);
xor U2601 (N_2601,N_1860,N_1469);
xor U2602 (N_2602,N_1719,N_1535);
nand U2603 (N_2603,N_2432,N_1521);
and U2604 (N_2604,N_1311,N_164);
nor U2605 (N_2605,N_1338,N_2011);
nand U2606 (N_2606,N_6,N_1167);
or U2607 (N_2607,N_978,N_550);
xnor U2608 (N_2608,N_2233,N_257);
nor U2609 (N_2609,N_808,N_156);
nand U2610 (N_2610,N_128,N_2453);
or U2611 (N_2611,N_585,N_780);
and U2612 (N_2612,N_700,N_436);
nand U2613 (N_2613,N_79,N_2070);
nor U2614 (N_2614,N_1431,N_2172);
or U2615 (N_2615,N_1998,N_338);
and U2616 (N_2616,N_817,N_2311);
nand U2617 (N_2617,N_1721,N_2224);
nor U2618 (N_2618,N_80,N_2032);
nor U2619 (N_2619,N_1876,N_385);
nor U2620 (N_2620,N_140,N_2103);
or U2621 (N_2621,N_1448,N_1974);
nand U2622 (N_2622,N_230,N_2036);
or U2623 (N_2623,N_1501,N_27);
nand U2624 (N_2624,N_145,N_1931);
or U2625 (N_2625,N_2299,N_713);
nor U2626 (N_2626,N_1645,N_502);
nand U2627 (N_2627,N_367,N_1387);
nand U2628 (N_2628,N_2349,N_424);
nor U2629 (N_2629,N_1581,N_1818);
nor U2630 (N_2630,N_860,N_698);
and U2631 (N_2631,N_779,N_1292);
nand U2632 (N_2632,N_2150,N_365);
xor U2633 (N_2633,N_52,N_360);
nor U2634 (N_2634,N_2167,N_96);
and U2635 (N_2635,N_162,N_2258);
and U2636 (N_2636,N_558,N_2305);
and U2637 (N_2637,N_2354,N_527);
nand U2638 (N_2638,N_2433,N_632);
and U2639 (N_2639,N_1746,N_1379);
or U2640 (N_2640,N_2335,N_444);
nand U2641 (N_2641,N_2345,N_382);
or U2642 (N_2642,N_74,N_2049);
and U2643 (N_2643,N_1176,N_2227);
and U2644 (N_2644,N_468,N_2370);
nor U2645 (N_2645,N_1953,N_2475);
nand U2646 (N_2646,N_1905,N_1759);
nor U2647 (N_2647,N_846,N_2251);
and U2648 (N_2648,N_1788,N_293);
nand U2649 (N_2649,N_2386,N_1248);
or U2650 (N_2650,N_1713,N_703);
nand U2651 (N_2651,N_34,N_539);
or U2652 (N_2652,N_2064,N_495);
and U2653 (N_2653,N_2368,N_2028);
or U2654 (N_2654,N_816,N_2374);
or U2655 (N_2655,N_1583,N_551);
or U2656 (N_2656,N_701,N_2343);
nor U2657 (N_2657,N_1234,N_820);
nand U2658 (N_2658,N_2175,N_1258);
and U2659 (N_2659,N_2088,N_524);
or U2660 (N_2660,N_598,N_2105);
nor U2661 (N_2661,N_1450,N_1825);
xor U2662 (N_2662,N_987,N_84);
or U2663 (N_2663,N_1490,N_2231);
and U2664 (N_2664,N_706,N_805);
and U2665 (N_2665,N_715,N_16);
or U2666 (N_2666,N_2169,N_1951);
nand U2667 (N_2667,N_1879,N_218);
and U2668 (N_2668,N_1426,N_1815);
nand U2669 (N_2669,N_1035,N_247);
or U2670 (N_2670,N_1391,N_339);
and U2671 (N_2671,N_1346,N_1481);
nand U2672 (N_2672,N_1203,N_1074);
or U2673 (N_2673,N_2493,N_39);
or U2674 (N_2674,N_297,N_1580);
nor U2675 (N_2675,N_1279,N_2187);
nor U2676 (N_2676,N_2003,N_195);
nor U2677 (N_2677,N_934,N_2361);
nand U2678 (N_2678,N_1752,N_657);
and U2679 (N_2679,N_2392,N_1364);
nand U2680 (N_2680,N_232,N_2288);
and U2681 (N_2681,N_2436,N_561);
nor U2682 (N_2682,N_2164,N_639);
and U2683 (N_2683,N_1978,N_1047);
nand U2684 (N_2684,N_320,N_2295);
and U2685 (N_2685,N_686,N_1454);
and U2686 (N_2686,N_1337,N_378);
nor U2687 (N_2687,N_834,N_731);
and U2688 (N_2688,N_742,N_941);
and U2689 (N_2689,N_1048,N_1239);
nand U2690 (N_2690,N_1836,N_1038);
and U2691 (N_2691,N_2483,N_1491);
nand U2692 (N_2692,N_1209,N_1003);
nor U2693 (N_2693,N_2306,N_175);
nor U2694 (N_2694,N_716,N_100);
nor U2695 (N_2695,N_1184,N_2087);
nor U2696 (N_2696,N_2225,N_1272);
nor U2697 (N_2697,N_499,N_1156);
nand U2698 (N_2698,N_1064,N_306);
and U2699 (N_2699,N_2146,N_2417);
nor U2700 (N_2700,N_2252,N_938);
nor U2701 (N_2701,N_1101,N_1121);
and U2702 (N_2702,N_51,N_1275);
nand U2703 (N_2703,N_192,N_1779);
or U2704 (N_2704,N_2029,N_1414);
nor U2705 (N_2705,N_1262,N_1875);
nor U2706 (N_2706,N_1786,N_1253);
or U2707 (N_2707,N_602,N_2055);
nand U2708 (N_2708,N_803,N_1862);
and U2709 (N_2709,N_2309,N_1560);
nand U2710 (N_2710,N_1839,N_2426);
and U2711 (N_2711,N_42,N_1251);
or U2712 (N_2712,N_1682,N_1028);
nor U2713 (N_2713,N_61,N_2066);
and U2714 (N_2714,N_2069,N_2056);
and U2715 (N_2715,N_2043,N_1175);
nor U2716 (N_2716,N_1559,N_903);
and U2717 (N_2717,N_395,N_1822);
or U2718 (N_2718,N_2238,N_2294);
nor U2719 (N_2719,N_2016,N_2131);
nand U2720 (N_2720,N_2470,N_908);
or U2721 (N_2721,N_1575,N_1445);
nand U2722 (N_2722,N_355,N_298);
nor U2723 (N_2723,N_1955,N_2437);
or U2724 (N_2724,N_1053,N_1658);
nor U2725 (N_2725,N_235,N_1664);
nand U2726 (N_2726,N_2239,N_2271);
nand U2727 (N_2727,N_2114,N_2302);
and U2728 (N_2728,N_97,N_1724);
nand U2729 (N_2729,N_463,N_909);
nand U2730 (N_2730,N_1689,N_1608);
xor U2731 (N_2731,N_2355,N_2473);
or U2732 (N_2732,N_2010,N_1551);
and U2733 (N_2733,N_1816,N_1402);
nand U2734 (N_2734,N_679,N_29);
nand U2735 (N_2735,N_1540,N_1052);
nor U2736 (N_2736,N_1888,N_973);
and U2737 (N_2737,N_1183,N_2362);
and U2738 (N_2738,N_1196,N_1604);
nand U2739 (N_2739,N_836,N_2357);
or U2740 (N_2740,N_2356,N_774);
nand U2741 (N_2741,N_1812,N_112);
nand U2742 (N_2742,N_691,N_895);
nor U2743 (N_2743,N_1057,N_2117);
nand U2744 (N_2744,N_1773,N_464);
nand U2745 (N_2745,N_848,N_183);
xor U2746 (N_2746,N_1056,N_1518);
nor U2747 (N_2747,N_2323,N_1784);
or U2748 (N_2748,N_1909,N_2428);
and U2749 (N_2749,N_41,N_2073);
or U2750 (N_2750,N_621,N_295);
nor U2751 (N_2751,N_1200,N_2081);
nand U2752 (N_2752,N_2100,N_1168);
nor U2753 (N_2753,N_500,N_1396);
nor U2754 (N_2754,N_1415,N_340);
nor U2755 (N_2755,N_1902,N_2274);
nor U2756 (N_2756,N_2179,N_352);
or U2757 (N_2757,N_501,N_361);
and U2758 (N_2758,N_40,N_2047);
nor U2759 (N_2759,N_2111,N_92);
nor U2760 (N_2760,N_2236,N_1138);
and U2761 (N_2761,N_1462,N_1565);
and U2762 (N_2762,N_1131,N_2441);
or U2763 (N_2763,N_1790,N_1158);
nor U2764 (N_2764,N_1971,N_1322);
nor U2765 (N_2765,N_99,N_1528);
nor U2766 (N_2766,N_718,N_1458);
and U2767 (N_2767,N_1170,N_656);
nor U2768 (N_2768,N_1690,N_234);
nand U2769 (N_2769,N_124,N_1576);
or U2770 (N_2770,N_1144,N_102);
and U2771 (N_2771,N_1384,N_605);
or U2772 (N_2772,N_1720,N_2468);
and U2773 (N_2773,N_750,N_2421);
and U2774 (N_2774,N_2405,N_1989);
nand U2775 (N_2775,N_689,N_1707);
nor U2776 (N_2776,N_2463,N_1004);
nor U2777 (N_2777,N_1480,N_1162);
nand U2778 (N_2778,N_745,N_32);
nand U2779 (N_2779,N_1392,N_1068);
nand U2780 (N_2780,N_2412,N_2275);
nor U2781 (N_2781,N_2109,N_1085);
or U2782 (N_2782,N_1073,N_1914);
or U2783 (N_2783,N_1141,N_2209);
nor U2784 (N_2784,N_738,N_1212);
nand U2785 (N_2785,N_1696,N_753);
nor U2786 (N_2786,N_966,N_59);
and U2787 (N_2787,N_2030,N_333);
nand U2788 (N_2788,N_144,N_2206);
nor U2789 (N_2789,N_304,N_1694);
nand U2790 (N_2790,N_619,N_2021);
nor U2791 (N_2791,N_969,N_1897);
nor U2792 (N_2792,N_1336,N_1446);
xor U2793 (N_2793,N_1103,N_683);
nand U2794 (N_2794,N_2353,N_1465);
nor U2795 (N_2795,N_1344,N_213);
and U2796 (N_2796,N_1276,N_2397);
and U2797 (N_2797,N_2234,N_55);
nand U2798 (N_2798,N_1164,N_1742);
nor U2799 (N_2799,N_2020,N_2431);
nor U2800 (N_2800,N_1342,N_1553);
or U2801 (N_2801,N_1350,N_1090);
and U2802 (N_2802,N_1671,N_2267);
and U2803 (N_2803,N_1115,N_572);
nor U2804 (N_2804,N_560,N_810);
or U2805 (N_2805,N_2488,N_366);
xor U2806 (N_2806,N_712,N_1265);
nor U2807 (N_2807,N_1401,N_1656);
nand U2808 (N_2808,N_1408,N_1325);
nand U2809 (N_2809,N_777,N_1901);
or U2810 (N_2810,N_2486,N_2075);
xnor U2811 (N_2811,N_1882,N_150);
xnor U2812 (N_2812,N_2147,N_680);
nand U2813 (N_2813,N_1892,N_961);
and U2814 (N_2814,N_1536,N_1929);
and U2815 (N_2815,N_1478,N_1832);
nand U2816 (N_2816,N_628,N_949);
or U2817 (N_2817,N_114,N_1728);
nor U2818 (N_2818,N_1009,N_1749);
nor U2819 (N_2819,N_48,N_121);
or U2820 (N_2820,N_335,N_336);
nand U2821 (N_2821,N_798,N_1590);
nor U2822 (N_2822,N_1296,N_2245);
or U2823 (N_2823,N_2264,N_858);
xor U2824 (N_2824,N_2050,N_1717);
and U2825 (N_2825,N_390,N_350);
nor U2826 (N_2826,N_1748,N_1061);
nor U2827 (N_2827,N_1735,N_1268);
or U2828 (N_2828,N_2422,N_1451);
or U2829 (N_2829,N_497,N_1700);
and U2830 (N_2830,N_2447,N_1143);
or U2831 (N_2831,N_2448,N_1018);
nand U2832 (N_2832,N_243,N_1142);
and U2833 (N_2833,N_1310,N_159);
nand U2834 (N_2834,N_107,N_696);
nor U2835 (N_2835,N_1443,N_199);
nor U2836 (N_2836,N_400,N_1877);
nand U2837 (N_2837,N_173,N_1406);
nand U2838 (N_2838,N_228,N_1800);
nor U2839 (N_2839,N_287,N_1821);
and U2840 (N_2840,N_1471,N_1783);
nand U2841 (N_2841,N_132,N_2487);
nand U2842 (N_2842,N_1383,N_453);
nor U2843 (N_2843,N_2165,N_1838);
nor U2844 (N_2844,N_904,N_705);
nand U2845 (N_2845,N_474,N_1343);
and U2846 (N_2846,N_138,N_725);
or U2847 (N_2847,N_1685,N_890);
nor U2848 (N_2848,N_2196,N_1084);
nor U2849 (N_2849,N_1125,N_1460);
and U2850 (N_2850,N_615,N_2315);
nand U2851 (N_2851,N_2138,N_1544);
nor U2852 (N_2852,N_1377,N_1649);
nor U2853 (N_2853,N_756,N_1274);
nor U2854 (N_2854,N_1747,N_1309);
and U2855 (N_2855,N_2325,N_2401);
or U2856 (N_2856,N_842,N_1150);
and U2857 (N_2857,N_2472,N_2192);
and U2858 (N_2858,N_930,N_313);
and U2859 (N_2859,N_945,N_1351);
nand U2860 (N_2860,N_1070,N_1136);
nand U2861 (N_2861,N_555,N_1938);
and U2862 (N_2862,N_1864,N_2254);
nand U2863 (N_2863,N_1264,N_1494);
nand U2864 (N_2864,N_511,N_2272);
nor U2865 (N_2865,N_1197,N_1045);
or U2866 (N_2866,N_2439,N_2474);
and U2867 (N_2867,N_872,N_1674);
and U2868 (N_2868,N_1966,N_2045);
or U2869 (N_2869,N_1792,N_1390);
xor U2870 (N_2870,N_126,N_19);
nor U2871 (N_2871,N_1944,N_63);
nand U2872 (N_2872,N_1113,N_1532);
or U2873 (N_2873,N_1372,N_1596);
nor U2874 (N_2874,N_763,N_2237);
nor U2875 (N_2875,N_1844,N_2443);
nand U2876 (N_2876,N_265,N_1841);
nand U2877 (N_2877,N_376,N_1005);
or U2878 (N_2878,N_654,N_2170);
and U2879 (N_2879,N_284,N_1291);
nand U2880 (N_2880,N_548,N_2166);
or U2881 (N_2881,N_449,N_1472);
and U2882 (N_2882,N_75,N_1767);
nand U2883 (N_2883,N_1716,N_586);
nor U2884 (N_2884,N_1352,N_1564);
nor U2885 (N_2885,N_36,N_12);
nor U2886 (N_2886,N_2026,N_1970);
nor U2887 (N_2887,N_2051,N_1960);
nand U2888 (N_2888,N_726,N_1934);
or U2889 (N_2889,N_929,N_2390);
nor U2890 (N_2890,N_425,N_1271);
nor U2891 (N_2891,N_2160,N_2438);
or U2892 (N_2892,N_1075,N_321);
nor U2893 (N_2893,N_273,N_452);
xor U2894 (N_2894,N_2136,N_1119);
nor U2895 (N_2895,N_465,N_205);
nand U2896 (N_2896,N_1542,N_1328);
nand U2897 (N_2897,N_503,N_1250);
nand U2898 (N_2898,N_1127,N_1851);
or U2899 (N_2899,N_1729,N_1202);
xnor U2900 (N_2900,N_2492,N_570);
nor U2901 (N_2901,N_1111,N_1059);
or U2902 (N_2902,N_197,N_1795);
nor U2903 (N_2903,N_1964,N_676);
nand U2904 (N_2904,N_154,N_821);
nor U2905 (N_2905,N_421,N_1793);
nor U2906 (N_2906,N_957,N_1801);
nand U2907 (N_2907,N_1243,N_364);
and U2908 (N_2908,N_439,N_1631);
and U2909 (N_2909,N_1405,N_2292);
nor U2910 (N_2910,N_2221,N_1733);
nor U2911 (N_2911,N_221,N_466);
nor U2912 (N_2912,N_1850,N_1904);
nor U2913 (N_2913,N_671,N_323);
or U2914 (N_2914,N_933,N_702);
and U2915 (N_2915,N_947,N_1872);
nor U2916 (N_2916,N_1163,N_1739);
nand U2917 (N_2917,N_920,N_1305);
xor U2918 (N_2918,N_1422,N_1506);
nand U2919 (N_2919,N_974,N_1573);
or U2920 (N_2920,N_1684,N_959);
nor U2921 (N_2921,N_1269,N_1598);
nand U2922 (N_2922,N_475,N_1116);
and U2923 (N_2923,N_1096,N_1019);
nand U2924 (N_2924,N_1549,N_2415);
and U2925 (N_2925,N_1438,N_2246);
or U2926 (N_2926,N_962,N_658);
or U2927 (N_2927,N_1927,N_1207);
and U2928 (N_2928,N_1348,N_2489);
or U2929 (N_2929,N_196,N_2380);
or U2930 (N_2930,N_1315,N_964);
and U2931 (N_2931,N_580,N_592);
and U2932 (N_2932,N_1657,N_1524);
or U2933 (N_2933,N_417,N_2340);
and U2934 (N_2934,N_785,N_1543);
and U2935 (N_2935,N_1201,N_547);
nand U2936 (N_2936,N_892,N_440);
and U2937 (N_2937,N_1678,N_388);
nand U2938 (N_2938,N_1956,N_1607);
or U2939 (N_2939,N_1531,N_1722);
or U2940 (N_2940,N_1776,N_1312);
nand U2941 (N_2941,N_179,N_2048);
and U2942 (N_2942,N_1781,N_515);
and U2943 (N_2943,N_369,N_1928);
nor U2944 (N_2944,N_311,N_708);
or U2945 (N_2945,N_2203,N_1630);
and U2946 (N_2946,N_850,N_1199);
nand U2947 (N_2947,N_2389,N_2243);
and U2948 (N_2948,N_300,N_1488);
and U2949 (N_2949,N_1854,N_1898);
nand U2950 (N_2950,N_94,N_1353);
and U2951 (N_2951,N_263,N_83);
and U2952 (N_2952,N_1007,N_1867);
and U2953 (N_2953,N_976,N_2313);
nor U2954 (N_2954,N_2304,N_1359);
nor U2955 (N_2955,N_1318,N_1208);
nand U2956 (N_2956,N_697,N_2148);
and U2957 (N_2957,N_1282,N_211);
nor U2958 (N_2958,N_936,N_732);
and U2959 (N_2959,N_1099,N_2185);
or U2960 (N_2960,N_1740,N_1252);
and U2961 (N_2961,N_1605,N_13);
and U2962 (N_2962,N_2076,N_608);
nor U2963 (N_2963,N_2019,N_481);
or U2964 (N_2964,N_447,N_677);
or U2965 (N_2965,N_182,N_105);
or U2966 (N_2966,N_1026,N_1358);
nor U2967 (N_2967,N_670,N_1789);
nand U2968 (N_2968,N_1132,N_2052);
nand U2969 (N_2969,N_152,N_143);
and U2970 (N_2970,N_912,N_1062);
and U2971 (N_2971,N_1436,N_902);
or U2972 (N_2972,N_2015,N_546);
nand U2973 (N_2973,N_1609,N_661);
or U2974 (N_2974,N_1417,N_1525);
nand U2975 (N_2975,N_2467,N_2014);
and U2976 (N_2976,N_1618,N_1824);
nor U2977 (N_2977,N_2096,N_2151);
nor U2978 (N_2978,N_498,N_133);
and U2979 (N_2979,N_2024,N_1219);
nor U2980 (N_2980,N_717,N_2074);
nor U2981 (N_2981,N_797,N_244);
and U2982 (N_2982,N_507,N_2477);
and U2983 (N_2983,N_1180,N_879);
or U2984 (N_2984,N_310,N_1247);
nor U2985 (N_2985,N_2285,N_1509);
or U2986 (N_2986,N_319,N_1151);
nor U2987 (N_2987,N_433,N_242);
or U2988 (N_2988,N_204,N_1246);
or U2989 (N_2989,N_1171,N_286);
or U2990 (N_2990,N_1081,N_393);
nor U2991 (N_2991,N_236,N_2359);
and U2992 (N_2992,N_250,N_261);
xor U2993 (N_2993,N_2255,N_299);
and U2994 (N_2994,N_1610,N_1847);
nor U2995 (N_2995,N_2348,N_1320);
or U2996 (N_2996,N_2139,N_2161);
and U2997 (N_2997,N_180,N_1484);
or U2998 (N_2998,N_1259,N_308);
and U2999 (N_2999,N_531,N_1750);
nor U3000 (N_3000,N_505,N_1129);
xnor U3001 (N_3001,N_217,N_1435);
nand U3002 (N_3002,N_862,N_1677);
or U3003 (N_3003,N_472,N_829);
nor U3004 (N_3004,N_1261,N_1906);
nand U3005 (N_3005,N_1903,N_398);
nand U3006 (N_3006,N_516,N_1412);
nand U3007 (N_3007,N_88,N_1122);
nand U3008 (N_3008,N_1987,N_2068);
nor U3009 (N_3009,N_662,N_216);
nand U3010 (N_3010,N_411,N_760);
nor U3011 (N_3011,N_1770,N_2301);
nand U3012 (N_3012,N_54,N_981);
or U3013 (N_3013,N_2465,N_1668);
and U3014 (N_3014,N_1334,N_735);
nor U3015 (N_3015,N_1811,N_1893);
xnor U3016 (N_3016,N_1845,N_435);
and U3017 (N_3017,N_1146,N_995);
and U3018 (N_3018,N_1493,N_1049);
nor U3019 (N_3019,N_754,N_1257);
nor U3020 (N_3020,N_109,N_2387);
nor U3021 (N_3021,N_788,N_430);
or U3022 (N_3022,N_1731,N_510);
nand U3023 (N_3023,N_1333,N_1709);
nand U3024 (N_3024,N_1194,N_1);
and U3025 (N_3025,N_1124,N_2002);
nand U3026 (N_3026,N_1662,N_875);
xnor U3027 (N_3027,N_490,N_5);
or U3028 (N_3028,N_983,N_2446);
nand U3029 (N_3029,N_1218,N_2180);
or U3030 (N_3030,N_869,N_210);
or U3031 (N_3031,N_1629,N_2418);
and U3032 (N_3032,N_2391,N_2135);
nor U3033 (N_3033,N_741,N_838);
xnor U3034 (N_3034,N_694,N_1008);
nand U3035 (N_3035,N_1295,N_806);
or U3036 (N_3036,N_46,N_2218);
xnor U3037 (N_3037,N_1385,N_1266);
and U3038 (N_3038,N_186,N_871);
nor U3039 (N_3039,N_729,N_583);
xor U3040 (N_3040,N_1743,N_1307);
nor U3041 (N_3041,N_2211,N_2186);
nand U3042 (N_3042,N_220,N_1582);
xor U3043 (N_3043,N_1873,N_2189);
nand U3044 (N_3044,N_2041,N_2424);
and U3045 (N_3045,N_591,N_833);
and U3046 (N_3046,N_2079,N_2038);
or U3047 (N_3047,N_1919,N_520);
nand U3048 (N_3048,N_926,N_758);
nor U3049 (N_3049,N_1686,N_482);
nand U3050 (N_3050,N_1849,N_1229);
and U3051 (N_3051,N_1267,N_1922);
and U3052 (N_3052,N_419,N_1277);
nor U3053 (N_3053,N_722,N_1945);
or U3054 (N_3054,N_168,N_1585);
nand U3055 (N_3055,N_282,N_2430);
nor U3056 (N_3056,N_134,N_1810);
nor U3057 (N_3057,N_1884,N_832);
xor U3058 (N_3058,N_545,N_704);
and U3059 (N_3059,N_95,N_2130);
or U3060 (N_3060,N_1673,N_1033);
and U3061 (N_3061,N_1058,N_970);
nor U3062 (N_3062,N_723,N_2482);
nor U3063 (N_3063,N_1255,N_781);
and U3064 (N_3064,N_744,N_2229);
or U3065 (N_3065,N_2022,N_49);
nor U3066 (N_3066,N_1014,N_270);
or U3067 (N_3067,N_1533,N_2204);
nor U3068 (N_3068,N_477,N_392);
and U3069 (N_3069,N_1149,N_1496);
and U3070 (N_3070,N_1619,N_460);
nand U3071 (N_3071,N_645,N_348);
and U3072 (N_3072,N_1428,N_1399);
nand U3073 (N_3073,N_190,N_420);
and U3074 (N_3074,N_2235,N_1853);
and U3075 (N_3075,N_574,N_719);
and U3076 (N_3076,N_1695,N_828);
nor U3077 (N_3077,N_208,N_886);
and U3078 (N_3078,N_2326,N_1077);
or U3079 (N_3079,N_2065,N_1361);
and U3080 (N_3080,N_1326,N_209);
nand U3081 (N_3081,N_770,N_841);
and U3082 (N_3082,N_1977,N_148);
nand U3083 (N_3083,N_975,N_2440);
or U3084 (N_3084,N_1530,N_1920);
or U3085 (N_3085,N_1464,N_1297);
and U3086 (N_3086,N_1615,N_260);
nand U3087 (N_3087,N_1787,N_494);
or U3088 (N_3088,N_1804,N_2458);
or U3089 (N_3089,N_1468,N_1123);
nand U3090 (N_3090,N_1991,N_93);
nor U3091 (N_3091,N_1702,N_1732);
and U3092 (N_3092,N_120,N_928);
xor U3093 (N_3093,N_1982,N_487);
or U3094 (N_3094,N_1210,N_720);
nor U3095 (N_3095,N_262,N_1486);
nand U3096 (N_3096,N_404,N_324);
or U3097 (N_3097,N_887,N_101);
xnor U3098 (N_3098,N_2344,N_2078);
and U3099 (N_3099,N_2257,N_1807);
and U3100 (N_3100,N_2371,N_1368);
nor U3101 (N_3101,N_831,N_918);
and U3102 (N_3102,N_768,N_2282);
or U3103 (N_3103,N_2399,N_1456);
or U3104 (N_3104,N_1244,N_775);
nand U3105 (N_3105,N_2296,N_2230);
nand U3106 (N_3106,N_1497,N_2300);
or U3107 (N_3107,N_913,N_1188);
and U3108 (N_3108,N_85,N_403);
and U3109 (N_3109,N_1675,N_2316);
or U3110 (N_3110,N_1441,N_529);
and U3111 (N_3111,N_824,N_916);
nor U3112 (N_3112,N_1301,N_2145);
nor U3113 (N_3113,N_682,N_241);
and U3114 (N_3114,N_2149,N_391);
and U3115 (N_3115,N_1316,N_2101);
and U3116 (N_3116,N_1958,N_1260);
nand U3117 (N_3117,N_1237,N_188);
xor U3118 (N_3118,N_1588,N_535);
nand U3119 (N_3119,N_1676,N_993);
nor U3120 (N_3120,N_1635,N_2452);
and U3121 (N_3121,N_325,N_2342);
nand U3122 (N_3122,N_946,N_772);
nor U3123 (N_3123,N_1923,N_231);
nand U3124 (N_3124,N_66,N_1245);
and U3125 (N_3125,N_1324,N_484);
or U3126 (N_3126,N_1562,N_1570);
nor U3127 (N_3127,N_240,N_1148);
or U3128 (N_3128,N_1794,N_1600);
nor U3129 (N_3129,N_386,N_1771);
or U3130 (N_3130,N_275,N_789);
nand U3131 (N_3131,N_1894,N_2382);
nor U3132 (N_3132,N_843,N_2459);
and U3133 (N_3133,N_512,N_765);
nor U3134 (N_3134,N_2480,N_1140);
nand U3135 (N_3135,N_556,N_2128);
nor U3136 (N_3136,N_2193,N_2321);
xor U3137 (N_3137,N_567,N_1775);
nand U3138 (N_3138,N_1545,N_776);
or U3139 (N_3139,N_1036,N_329);
nor U3140 (N_3140,N_1510,N_149);
nand U3141 (N_3141,N_371,N_1397);
and U3142 (N_3142,N_312,N_751);
nor U3143 (N_3143,N_429,N_223);
and U3144 (N_3144,N_2144,N_442);
nand U3145 (N_3145,N_1890,N_237);
and U3146 (N_3146,N_136,N_637);
or U3147 (N_3147,N_1537,N_489);
and U3148 (N_3148,N_1681,N_852);
xor U3149 (N_3149,N_2214,N_986);
or U3150 (N_3150,N_1782,N_1409);
and U3151 (N_3151,N_584,N_925);
nor U3152 (N_3152,N_1041,N_881);
and U3153 (N_3153,N_1249,N_940);
nor U3154 (N_3154,N_893,N_1959);
and U3155 (N_3155,N_563,N_1155);
and U3156 (N_3156,N_1624,N_518);
and U3157 (N_3157,N_2481,N_2046);
nand U3158 (N_3158,N_660,N_264);
and U3159 (N_3159,N_89,N_2314);
or U3160 (N_3160,N_845,N_883);
nor U3161 (N_3161,N_2407,N_283);
and U3162 (N_3162,N_1883,N_1204);
nor U3163 (N_3163,N_341,N_2097);
and U3164 (N_3164,N_1511,N_1968);
nand U3165 (N_3165,N_2256,N_2435);
and U3166 (N_3166,N_1670,N_1482);
nand U3167 (N_3167,N_1843,N_422);
or U3168 (N_3168,N_301,N_519);
and U3169 (N_3169,N_2266,N_1737);
or U3170 (N_3170,N_389,N_1706);
nand U3171 (N_3171,N_73,N_849);
or U3172 (N_3172,N_1606,N_2007);
nand U3173 (N_3173,N_752,N_1190);
nand U3174 (N_3174,N_76,N_1529);
nand U3175 (N_3175,N_1466,N_2455);
and U3176 (N_3176,N_630,N_414);
and U3177 (N_3177,N_1766,N_578);
or U3178 (N_3178,N_1160,N_117);
nor U3179 (N_3179,N_2142,N_907);
and U3180 (N_3180,N_399,N_1221);
nor U3181 (N_3181,N_1055,N_2190);
nor U3182 (N_3182,N_269,N_1425);
or U3183 (N_3183,N_2090,N_58);
nor U3184 (N_3184,N_1652,N_2334);
nor U3185 (N_3185,N_1487,N_288);
or U3186 (N_3186,N_317,N_127);
or U3187 (N_3187,N_358,N_1601);
nand U3188 (N_3188,N_1360,N_693);
or U3189 (N_3189,N_130,N_1345);
nor U3190 (N_3190,N_791,N_457);
or U3191 (N_3191,N_2378,N_1895);
or U3192 (N_3192,N_2322,N_1015);
nand U3193 (N_3193,N_1120,N_71);
nor U3194 (N_3194,N_649,N_513);
nand U3195 (N_3195,N_1718,N_1741);
nand U3196 (N_3196,N_1105,N_33);
or U3197 (N_3197,N_1889,N_801);
nand U3198 (N_3198,N_952,N_1976);
or U3199 (N_3199,N_748,N_1546);
nand U3200 (N_3200,N_1913,N_618);
and U3201 (N_3201,N_246,N_2464);
and U3202 (N_3202,N_1917,N_2416);
nor U3203 (N_3203,N_292,N_2469);
and U3204 (N_3204,N_1040,N_1830);
and U3205 (N_3205,N_1622,N_526);
or U3206 (N_3206,N_172,N_455);
or U3207 (N_3207,N_1764,N_1758);
nor U3208 (N_3208,N_616,N_576);
nand U3209 (N_3209,N_967,N_2198);
nor U3210 (N_3210,N_837,N_839);
nand U3211 (N_3211,N_160,N_1768);
nand U3212 (N_3212,N_2278,N_564);
or U3213 (N_3213,N_207,N_342);
nand U3214 (N_3214,N_1933,N_1023);
nor U3215 (N_3215,N_796,N_11);
nor U3216 (N_3216,N_950,N_1683);
nand U3217 (N_3217,N_1637,N_1054);
xor U3218 (N_3218,N_53,N_1969);
or U3219 (N_3219,N_1037,N_2173);
xnor U3220 (N_3220,N_935,N_857);
nor U3221 (N_3221,N_1017,N_363);
and U3222 (N_3222,N_2479,N_2291);
and U3223 (N_3223,N_252,N_1745);
nand U3224 (N_3224,N_736,N_607);
nor U3225 (N_3225,N_1753,N_919);
and U3226 (N_3226,N_108,N_674);
nand U3227 (N_3227,N_2195,N_1187);
or U3228 (N_3228,N_665,N_2384);
or U3229 (N_3229,N_1181,N_1523);
and U3230 (N_3230,N_458,N_965);
and U3231 (N_3231,N_1106,N_1440);
nor U3232 (N_3232,N_1679,N_1937);
nor U3233 (N_3233,N_644,N_536);
nand U3234 (N_3234,N_1287,N_125);
or U3235 (N_3235,N_884,N_517);
nor U3236 (N_3236,N_2140,N_2269);
nand U3237 (N_3237,N_767,N_82);
and U3238 (N_3238,N_1626,N_2336);
nand U3239 (N_3239,N_1335,N_802);
nor U3240 (N_3240,N_994,N_1613);
nand U3241 (N_3241,N_2268,N_2338);
nand U3242 (N_3242,N_113,N_1985);
nor U3243 (N_3243,N_2158,N_2121);
and U3244 (N_3244,N_739,N_206);
and U3245 (N_3245,N_68,N_1066);
nand U3246 (N_3246,N_7,N_1433);
nor U3247 (N_3247,N_1461,N_2013);
or U3248 (N_3248,N_119,N_542);
nand U3249 (N_3249,N_2327,N_98);
or U3250 (N_3250,N_1193,N_1648);
nor U3251 (N_3251,N_1711,N_827);
or U3252 (N_3252,N_1093,N_1306);
or U3253 (N_3253,N_678,N_122);
and U3254 (N_3254,N_1474,N_337);
nor U3255 (N_3255,N_2373,N_2290);
nand U3256 (N_3256,N_189,N_1802);
or U3257 (N_3257,N_1388,N_1323);
xor U3258 (N_3258,N_1134,N_2126);
or U3259 (N_3259,N_280,N_1503);
and U3260 (N_3260,N_2466,N_1572);
and U3261 (N_3261,N_1861,N_1950);
or U3262 (N_3262,N_648,N_2406);
and U3263 (N_3263,N_1561,N_1828);
nand U3264 (N_3264,N_1407,N_2337);
nor U3265 (N_3265,N_2163,N_894);
nand U3266 (N_3266,N_1972,N_1254);
nand U3267 (N_3267,N_1620,N_2210);
or U3268 (N_3268,N_10,N_1512);
nor U3269 (N_3269,N_1118,N_1072);
and U3270 (N_3270,N_1192,N_577);
nand U3271 (N_3271,N_2071,N_587);
or U3272 (N_3272,N_2040,N_814);
nor U3273 (N_3273,N_2347,N_971);
nor U3274 (N_3274,N_1642,N_1602);
nand U3275 (N_3275,N_2402,N_1479);
or U3276 (N_3276,N_90,N_118);
nor U3277 (N_3277,N_2034,N_642);
nand U3278 (N_3278,N_727,N_1453);
or U3279 (N_3279,N_506,N_1042);
nand U3280 (N_3280,N_1534,N_1869);
and U3281 (N_3281,N_2120,N_408);
nor U3282 (N_3282,N_412,N_1102);
or U3283 (N_3283,N_984,N_1761);
or U3284 (N_3284,N_888,N_2425);
nor U3285 (N_3285,N_1666,N_1527);
nand U3286 (N_3286,N_695,N_226);
and U3287 (N_3287,N_1538,N_1161);
and U3288 (N_3288,N_866,N_2461);
nand U3289 (N_3289,N_1878,N_819);
nand U3290 (N_3290,N_2023,N_1981);
or U3291 (N_3291,N_2450,N_2217);
or U3292 (N_3292,N_1191,N_1852);
nor U3293 (N_3293,N_1999,N_549);
or U3294 (N_3294,N_456,N_141);
nor U3295 (N_3295,N_1725,N_508);
nand U3296 (N_3296,N_1698,N_1386);
or U3297 (N_3297,N_1371,N_2080);
nand U3298 (N_3298,N_2286,N_2320);
and U3299 (N_3299,N_956,N_625);
nand U3300 (N_3300,N_1489,N_728);
nand U3301 (N_3301,N_559,N_18);
and U3302 (N_3302,N_309,N_999);
xnor U3303 (N_3303,N_910,N_2042);
nand U3304 (N_3304,N_1848,N_861);
nand U3305 (N_3305,N_1755,N_1376);
and U3306 (N_3306,N_2454,N_2159);
and U3307 (N_3307,N_91,N_1439);
nor U3308 (N_3308,N_1463,N_147);
nand U3309 (N_3309,N_343,N_537);
nand U3310 (N_3310,N_1691,N_2381);
and U3311 (N_3311,N_931,N_663);
and U3312 (N_3312,N_1710,N_1104);
and U3313 (N_3313,N_2033,N_1963);
nor U3314 (N_3314,N_924,N_1508);
and U3315 (N_3315,N_2122,N_1051);
nand U3316 (N_3316,N_1421,N_328);
and U3317 (N_3317,N_1012,N_1178);
nand U3318 (N_3318,N_368,N_1137);
or U3319 (N_3319,N_557,N_977);
nor U3320 (N_3320,N_1434,N_353);
and U3321 (N_3321,N_1327,N_1757);
or U3322 (N_3322,N_479,N_1505);
and U3323 (N_3323,N_2062,N_8);
nand U3324 (N_3324,N_932,N_870);
and U3325 (N_3325,N_86,N_357);
and U3326 (N_3326,N_1996,N_1366);
and U3327 (N_3327,N_2181,N_248);
and U3328 (N_3328,N_1427,N_1921);
and U3329 (N_3329,N_1858,N_1857);
nand U3330 (N_3330,N_1294,N_2442);
and U3331 (N_3331,N_921,N_1001);
or U3332 (N_3332,N_1437,N_854);
nand U3333 (N_3333,N_1300,N_1152);
and U3334 (N_3334,N_2404,N_291);
or U3335 (N_3335,N_1751,N_800);
or U3336 (N_3336,N_2215,N_1065);
and U3337 (N_3337,N_1704,N_891);
nand U3338 (N_3338,N_1080,N_2365);
nand U3339 (N_3339,N_634,N_2244);
and U3340 (N_3340,N_200,N_569);
nand U3341 (N_3341,N_491,N_2449);
or U3342 (N_3342,N_1621,N_2184);
or U3343 (N_3343,N_2154,N_2411);
or U3344 (N_3344,N_985,N_57);
or U3345 (N_3345,N_1855,N_2053);
nand U3346 (N_3346,N_258,N_2118);
or U3347 (N_3347,N_523,N_1403);
nor U3348 (N_3348,N_1347,N_566);
nand U3349 (N_3349,N_331,N_2129);
nor U3350 (N_3350,N_1571,N_2093);
nand U3351 (N_3351,N_2491,N_1492);
nor U3352 (N_3352,N_2329,N_1502);
nand U3353 (N_3353,N_533,N_2276);
and U3354 (N_3354,N_2499,N_922);
nand U3355 (N_3355,N_2241,N_1088);
or U3356 (N_3356,N_1597,N_1769);
nor U3357 (N_3357,N_997,N_2072);
and U3358 (N_3358,N_1513,N_1574);
and U3359 (N_3359,N_1016,N_356);
nor U3360 (N_3360,N_1173,N_135);
or U3361 (N_3361,N_951,N_737);
nor U3362 (N_3362,N_1498,N_1774);
nand U3363 (N_3363,N_1242,N_795);
nor U3364 (N_3364,N_766,N_2057);
nor U3365 (N_3365,N_185,N_2498);
nand U3366 (N_3366,N_1220,N_1416);
nand U3367 (N_3367,N_2318,N_699);
nand U3368 (N_3368,N_2279,N_2297);
or U3369 (N_3369,N_743,N_1910);
nor U3370 (N_3370,N_794,N_2035);
nand U3371 (N_3371,N_157,N_1429);
and U3372 (N_3372,N_25,N_238);
and U3373 (N_3373,N_2141,N_2460);
and U3374 (N_3374,N_972,N_1082);
or U3375 (N_3375,N_413,N_707);
or U3376 (N_3376,N_1557,N_1413);
nor U3377 (N_3377,N_2375,N_1646);
or U3378 (N_3378,N_1109,N_581);
or U3379 (N_3379,N_1639,N_646);
nand U3380 (N_3380,N_1547,N_470);
and U3381 (N_3381,N_346,N_1515);
or U3382 (N_3382,N_2310,N_1092);
nand U3383 (N_3383,N_1589,N_1697);
or U3384 (N_3384,N_757,N_473);
and U3385 (N_3385,N_1419,N_1834);
nor U3386 (N_3386,N_2201,N_1031);
and U3387 (N_3387,N_1217,N_1232);
nor U3388 (N_3388,N_1859,N_681);
xor U3389 (N_3389,N_2485,N_534);
nor U3390 (N_3390,N_2094,N_2124);
nand U3391 (N_3391,N_407,N_2134);
nor U3392 (N_3392,N_1339,N_2328);
and U3393 (N_3393,N_375,N_70);
and U3394 (N_3394,N_23,N_2490);
or U3395 (N_3395,N_2363,N_396);
xor U3396 (N_3396,N_873,N_1962);
or U3397 (N_3397,N_2242,N_1625);
nand U3398 (N_3398,N_2457,N_530);
and U3399 (N_3399,N_1911,N_1224);
or U3400 (N_3400,N_734,N_2312);
nor U3401 (N_3401,N_214,N_1997);
nor U3402 (N_3402,N_2085,N_509);
and U3403 (N_3403,N_330,N_514);
nand U3404 (N_3404,N_1647,N_406);
nor U3405 (N_3405,N_437,N_374);
nor U3406 (N_3406,N_2319,N_1034);
nor U3407 (N_3407,N_589,N_110);
xnor U3408 (N_3408,N_714,N_459);
nor U3409 (N_3409,N_1655,N_2484);
nor U3410 (N_3410,N_1723,N_2385);
nor U3411 (N_3411,N_483,N_1837);
or U3412 (N_3412,N_2494,N_864);
and U3413 (N_3413,N_1813,N_2434);
nor U3414 (N_3414,N_1587,N_1370);
nand U3415 (N_3415,N_1189,N_1653);
nand U3416 (N_3416,N_1814,N_2396);
nor U3417 (N_3417,N_1550,N_245);
and U3418 (N_3418,N_2423,N_749);
nand U3419 (N_3419,N_818,N_1304);
nor U3420 (N_3420,N_1734,N_1331);
nor U3421 (N_3421,N_155,N_540);
nand U3422 (N_3422,N_960,N_2031);
and U3423 (N_3423,N_2058,N_582);
or U3424 (N_3424,N_2200,N_31);
nand U3425 (N_3425,N_1159,N_212);
nand U3426 (N_3426,N_1988,N_2082);
and U3427 (N_3427,N_2213,N_2178);
nand U3428 (N_3428,N_1135,N_565);
nand U3429 (N_3429,N_2194,N_2332);
or U3430 (N_3430,N_631,N_2414);
or U3431 (N_3431,N_281,N_1500);
and U3432 (N_3432,N_1290,N_783);
nor U3433 (N_3433,N_809,N_588);
and U3434 (N_3434,N_2095,N_67);
nor U3435 (N_3435,N_823,N_1128);
nor U3436 (N_3436,N_874,N_1868);
nor U3437 (N_3437,N_485,N_1298);
nor U3438 (N_3438,N_1593,N_87);
nor U3439 (N_3439,N_379,N_1943);
and U3440 (N_3440,N_1899,N_72);
nor U3441 (N_3441,N_1288,N_383);
nor U3442 (N_3442,N_1025,N_2216);
and U3443 (N_3443,N_271,N_111);
nor U3444 (N_3444,N_2259,N_1599);
and U3445 (N_3445,N_471,N_1114);
or U3446 (N_3446,N_123,N_1069);
nand U3447 (N_3447,N_769,N_784);
and U3448 (N_3448,N_254,N_450);
or U3449 (N_3449,N_2408,N_1907);
nor U3450 (N_3450,N_2039,N_1577);
and U3451 (N_3451,N_2360,N_1293);
and U3452 (N_3452,N_1455,N_847);
and U3453 (N_3453,N_968,N_1754);
and U3454 (N_3454,N_443,N_397);
and U3455 (N_3455,N_1541,N_2183);
nand U3456 (N_3456,N_2283,N_799);
or U3457 (N_3457,N_2462,N_1949);
and U3458 (N_3458,N_1313,N_1627);
and U3459 (N_3459,N_1400,N_1712);
or U3460 (N_3460,N_77,N_201);
and U3461 (N_3461,N_1030,N_28);
and U3462 (N_3462,N_786,N_1846);
nor U3463 (N_3463,N_9,N_1760);
and U3464 (N_3464,N_2317,N_1863);
nand U3465 (N_3465,N_1317,N_1094);
and U3466 (N_3466,N_2331,N_1356);
or U3467 (N_3467,N_401,N_2451);
nor U3468 (N_3468,N_1389,N_1108);
nor U3469 (N_3469,N_2265,N_943);
nand U3470 (N_3470,N_1778,N_1578);
or U3471 (N_3471,N_2496,N_2471);
or U3472 (N_3472,N_1667,N_1228);
and U3473 (N_3473,N_2001,N_1165);
and U3474 (N_3474,N_778,N_1499);
and U3475 (N_3475,N_1100,N_2220);
xor U3476 (N_3476,N_274,N_253);
or U3477 (N_3477,N_370,N_1285);
or U3478 (N_3478,N_1797,N_1993);
nand U3479 (N_3479,N_2222,N_1616);
or U3480 (N_3480,N_1896,N_2086);
and U3481 (N_3481,N_2366,N_1881);
or U3482 (N_3482,N_1011,N_153);
nor U3483 (N_3483,N_2284,N_1174);
and U3484 (N_3484,N_1935,N_944);
nand U3485 (N_3485,N_991,N_1780);
or U3486 (N_3486,N_1182,N_793);
nor U3487 (N_3487,N_2025,N_1520);
nor U3488 (N_3488,N_1584,N_2367);
nand U3489 (N_3489,N_362,N_617);
nor U3490 (N_3490,N_595,N_139);
nand U3491 (N_3491,N_666,N_2171);
nand U3492 (N_3492,N_2429,N_2089);
or U3493 (N_3493,N_203,N_2273);
nand U3494 (N_3494,N_445,N_773);
and U3495 (N_3495,N_771,N_1803);
xor U3496 (N_3496,N_552,N_1117);
and U3497 (N_3497,N_1223,N_47);
and U3498 (N_3498,N_1130,N_568);
nor U3499 (N_3499,N_2497,N_194);
and U3500 (N_3500,N_2188,N_2298);
nand U3501 (N_3501,N_296,N_2376);
nor U3502 (N_3502,N_1024,N_815);
nand U3503 (N_3503,N_1010,N_1195);
xnor U3504 (N_3504,N_905,N_1856);
nor U3505 (N_3505,N_2351,N_2293);
and U3506 (N_3506,N_1169,N_2308);
nor U3507 (N_3507,N_623,N_1586);
and U3508 (N_3508,N_855,N_1078);
nor U3509 (N_3509,N_1235,N_277);
nor U3510 (N_3510,N_2199,N_740);
nor U3511 (N_3511,N_476,N_2240);
or U3512 (N_3512,N_1591,N_1225);
nand U3513 (N_3513,N_601,N_1808);
and U3514 (N_3514,N_2333,N_1526);
nand U3515 (N_3515,N_215,N_1730);
nand U3516 (N_3516,N_2205,N_1172);
and U3517 (N_3517,N_543,N_979);
or U3518 (N_3518,N_373,N_2394);
nor U3519 (N_3519,N_469,N_990);
and U3520 (N_3520,N_1885,N_1809);
and U3521 (N_3521,N_1286,N_2495);
and U3522 (N_3522,N_684,N_1617);
nand U3523 (N_3523,N_2061,N_710);
nor U3524 (N_3524,N_1179,N_2289);
nor U3525 (N_3525,N_255,N_2413);
nor U3526 (N_3526,N_1032,N_1046);
or U3527 (N_3527,N_2092,N_614);
and U3528 (N_3528,N_1975,N_620);
or U3529 (N_3529,N_2476,N_1021);
nand U3530 (N_3530,N_2262,N_2358);
and U3531 (N_3531,N_1603,N_2119);
or U3532 (N_3532,N_1961,N_633);
and U3533 (N_3533,N_2009,N_927);
or U3534 (N_3534,N_915,N_2091);
nor U3535 (N_3535,N_191,N_1222);
or U3536 (N_3536,N_822,N_1185);
nor U3537 (N_3537,N_416,N_627);
nor U3538 (N_3538,N_896,N_1772);
or U3539 (N_3539,N_1984,N_1539);
nand U3540 (N_3540,N_268,N_579);
nand U3541 (N_3541,N_954,N_2324);
or U3542 (N_3542,N_690,N_423);
or U3543 (N_3543,N_441,N_1865);
nand U3544 (N_3544,N_2125,N_1638);
and U3545 (N_3545,N_2202,N_596);
nor U3546 (N_3546,N_1424,N_2123);
nand U3547 (N_3547,N_69,N_193);
and U3548 (N_3548,N_303,N_2156);
and U3549 (N_3549,N_1374,N_1833);
nand U3550 (N_3550,N_44,N_1240);
nor U3551 (N_3551,N_1420,N_1886);
or U3552 (N_3552,N_2364,N_853);
or U3553 (N_3553,N_426,N_2410);
or U3554 (N_3554,N_1823,N_2350);
or U3555 (N_3555,N_687,N_880);
nand U3556 (N_3556,N_1205,N_1133);
or U3557 (N_3557,N_1714,N_1302);
nor U3558 (N_3558,N_590,N_2247);
nand U3559 (N_3559,N_643,N_259);
nor U3560 (N_3560,N_2099,N_1089);
and U3561 (N_3561,N_1992,N_359);
nor U3562 (N_3562,N_635,N_1842);
nand U3563 (N_3563,N_942,N_1153);
nor U3564 (N_3564,N_1086,N_294);
or U3565 (N_3565,N_1299,N_1912);
nand U3566 (N_3566,N_1556,N_2115);
nand U3567 (N_3567,N_865,N_764);
nand U3568 (N_3568,N_640,N_1215);
nand U3569 (N_3569,N_1611,N_115);
and U3570 (N_3570,N_1050,N_1382);
nand U3571 (N_3571,N_1284,N_45);
or U3572 (N_3572,N_1819,N_1483);
or U3573 (N_3573,N_835,N_427);
or U3574 (N_3574,N_1319,N_1946);
and U3575 (N_3575,N_1198,N_1941);
or U3576 (N_3576,N_575,N_142);
or U3577 (N_3577,N_2400,N_2044);
nor U3578 (N_3578,N_525,N_844);
nand U3579 (N_3579,N_1394,N_224);
or U3580 (N_3580,N_1567,N_1470);
nand U3581 (N_3581,N_532,N_1569);
or U3582 (N_3582,N_1112,N_1432);
and U3583 (N_3583,N_3,N_1430);
nor U3584 (N_3584,N_15,N_1614);
nand U3585 (N_3585,N_176,N_1280);
nand U3586 (N_3586,N_711,N_1663);
or U3587 (N_3587,N_2250,N_813);
or U3588 (N_3588,N_1634,N_1447);
or U3589 (N_3589,N_1680,N_622);
nand U3590 (N_3590,N_1236,N_882);
nor U3591 (N_3591,N_1688,N_1965);
or U3592 (N_3592,N_655,N_2104);
nor U3593 (N_3593,N_761,N_1477);
or U3594 (N_3594,N_600,N_2004);
xnor U3595 (N_3595,N_1449,N_174);
nor U3596 (N_3596,N_2339,N_1256);
nor U3597 (N_3597,N_1744,N_2352);
or U3598 (N_3598,N_1829,N_782);
or U3599 (N_3599,N_611,N_538);
nand U3600 (N_3600,N_1349,N_2106);
nand U3601 (N_3601,N_906,N_1308);
or U3602 (N_3602,N_790,N_30);
nor U3603 (N_3603,N_953,N_314);
and U3604 (N_3604,N_184,N_1918);
nor U3605 (N_3605,N_897,N_721);
nand U3606 (N_3606,N_387,N_1241);
nand U3607 (N_3607,N_65,N_1022);
nand U3608 (N_3608,N_1952,N_812);
nor U3609 (N_3609,N_432,N_2113);
and U3610 (N_3610,N_272,N_1940);
nand U3611 (N_3611,N_1467,N_1278);
and U3612 (N_3612,N_22,N_571);
nor U3613 (N_3613,N_1476,N_2153);
and U3614 (N_3614,N_1835,N_2137);
and U3615 (N_3615,N_354,N_492);
and U3616 (N_3616,N_1516,N_1672);
and U3617 (N_3617,N_1514,N_2182);
and U3618 (N_3618,N_1887,N_2177);
nor U3619 (N_3619,N_1442,N_1926);
or U3620 (N_3620,N_229,N_2037);
nand U3621 (N_3621,N_2395,N_2102);
and U3622 (N_3622,N_613,N_917);
nor U3623 (N_3623,N_1504,N_2307);
nand U3624 (N_3624,N_478,N_2280);
nand U3625 (N_3625,N_1095,N_202);
and U3626 (N_3626,N_1329,N_106);
nand U3627 (N_3627,N_2226,N_1303);
nor U3628 (N_3628,N_2409,N_1900);
nor U3629 (N_3629,N_158,N_1029);
nor U3630 (N_3630,N_1186,N_2208);
or U3631 (N_3631,N_266,N_1039);
and U3632 (N_3632,N_1145,N_1777);
or U3633 (N_3633,N_856,N_278);
and U3634 (N_3634,N_1213,N_1967);
nand U3635 (N_3635,N_1380,N_187);
nand U3636 (N_3636,N_1669,N_26);
or U3637 (N_3637,N_2260,N_1939);
or U3638 (N_3638,N_1866,N_2060);
and U3639 (N_3639,N_830,N_1798);
and U3640 (N_3640,N_762,N_876);
nor U3641 (N_3641,N_1087,N_62);
nor U3642 (N_3642,N_486,N_431);
nand U3643 (N_3643,N_1354,N_1595);
nand U3644 (N_3644,N_438,N_496);
or U3645 (N_3645,N_1826,N_1230);
xor U3646 (N_3646,N_2287,N_609);
or U3647 (N_3647,N_222,N_1579);
and U3648 (N_3648,N_227,N_163);
nor U3649 (N_3649,N_1044,N_541);
nand U3650 (N_3650,N_1063,N_899);
or U3651 (N_3651,N_636,N_289);
nand U3652 (N_3652,N_2456,N_1891);
nor U3653 (N_3653,N_1791,N_2098);
and U3654 (N_3654,N_1651,N_593);
and U3655 (N_3655,N_1369,N_2420);
nor U3656 (N_3656,N_1805,N_1126);
nor U3657 (N_3657,N_2403,N_1060);
nand U3658 (N_3658,N_1211,N_889);
and U3659 (N_3659,N_1076,N_1475);
and U3660 (N_3660,N_1363,N_688);
nand U3661 (N_3661,N_1238,N_2155);
nand U3662 (N_3662,N_20,N_1273);
nor U3663 (N_3663,N_629,N_17);
and U3664 (N_3664,N_24,N_225);
and U3665 (N_3665,N_0,N_653);
and U3666 (N_3666,N_402,N_451);
or U3667 (N_3667,N_2232,N_249);
nand U3668 (N_3668,N_1393,N_2427);
or U3669 (N_3669,N_2419,N_1362);
nand U3670 (N_3670,N_488,N_345);
nand U3671 (N_3671,N_1289,N_2377);
and U3672 (N_3672,N_1936,N_1206);
and U3673 (N_3673,N_1763,N_1027);
or U3674 (N_3674,N_1756,N_1558);
xor U3675 (N_3675,N_939,N_198);
nand U3676 (N_3676,N_2388,N_1973);
nor U3677 (N_3677,N_900,N_131);
nand U3678 (N_3678,N_948,N_2207);
or U3679 (N_3679,N_594,N_1566);
or U3680 (N_3680,N_2197,N_1693);
or U3681 (N_3681,N_2346,N_1002);
or U3682 (N_3682,N_1270,N_276);
and U3683 (N_3683,N_1708,N_1166);
and U3684 (N_3684,N_937,N_1636);
and U3685 (N_3685,N_349,N_604);
and U3686 (N_3686,N_1013,N_332);
or U3687 (N_3687,N_43,N_1995);
nor U3688 (N_3688,N_672,N_1692);
or U3689 (N_3689,N_1703,N_1410);
and U3690 (N_3690,N_1765,N_1924);
and U3691 (N_3691,N_380,N_14);
or U3692 (N_3692,N_641,N_2478);
or U3693 (N_3693,N_1665,N_1762);
nor U3694 (N_3694,N_811,N_37);
nor U3695 (N_3695,N_1522,N_233);
nand U3696 (N_3696,N_167,N_1806);
nand U3697 (N_3697,N_859,N_1216);
nand U3698 (N_3698,N_1715,N_351);
nand U3699 (N_3699,N_116,N_409);
nor U3700 (N_3700,N_1817,N_522);
or U3701 (N_3701,N_1871,N_733);
or U3702 (N_3702,N_1355,N_1378);
and U3703 (N_3703,N_1785,N_1957);
nor U3704 (N_3704,N_1563,N_1020);
nand U3705 (N_3705,N_2083,N_2303);
nor U3706 (N_3706,N_1341,N_410);
and U3707 (N_3707,N_1404,N_2212);
nand U3708 (N_3708,N_1398,N_1568);
xnor U3709 (N_3709,N_171,N_2444);
or U3710 (N_3710,N_2000,N_1840);
nor U3711 (N_3711,N_1006,N_1874);
nor U3712 (N_3712,N_1373,N_2116);
nor U3713 (N_3713,N_1799,N_1154);
nand U3714 (N_3714,N_1485,N_2445);
or U3715 (N_3715,N_610,N_1980);
or U3716 (N_3716,N_2005,N_1916);
nor U3717 (N_3717,N_81,N_898);
nor U3718 (N_3718,N_914,N_251);
nor U3719 (N_3719,N_2059,N_652);
nor U3720 (N_3720,N_434,N_2168);
nand U3721 (N_3721,N_2341,N_1954);
and U3722 (N_3722,N_1495,N_322);
nor U3723 (N_3723,N_1332,N_659);
and U3724 (N_3724,N_1554,N_2369);
nand U3725 (N_3725,N_1705,N_1796);
or U3726 (N_3726,N_381,N_1555);
nand U3727 (N_3727,N_405,N_2281);
nor U3728 (N_3728,N_256,N_1098);
nand U3729 (N_3729,N_344,N_1231);
nor U3730 (N_3730,N_877,N_2261);
nor U3731 (N_3731,N_804,N_1000);
or U3732 (N_3732,N_334,N_755);
or U3733 (N_3733,N_2372,N_1594);
nor U3734 (N_3734,N_219,N_1644);
nor U3735 (N_3735,N_1381,N_2077);
nor U3736 (N_3736,N_2133,N_151);
and U3737 (N_3737,N_1365,N_1067);
nand U3738 (N_3738,N_851,N_746);
nand U3739 (N_3739,N_327,N_2219);
nand U3740 (N_3740,N_1986,N_315);
nand U3741 (N_3741,N_50,N_267);
nand U3742 (N_3742,N_181,N_285);
and U3743 (N_3743,N_573,N_963);
nor U3744 (N_3744,N_1110,N_467);
and U3745 (N_3745,N_1990,N_1979);
nand U3746 (N_3746,N_1548,N_394);
nand U3747 (N_3747,N_1375,N_685);
nand U3748 (N_3748,N_599,N_675);
nor U3749 (N_3749,N_38,N_988);
nor U3750 (N_3750,N_1238,N_487);
nor U3751 (N_3751,N_71,N_946);
nor U3752 (N_3752,N_94,N_1610);
or U3753 (N_3753,N_2206,N_585);
nor U3754 (N_3754,N_791,N_2044);
nor U3755 (N_3755,N_1037,N_259);
nand U3756 (N_3756,N_421,N_2496);
nand U3757 (N_3757,N_2090,N_1040);
nor U3758 (N_3758,N_1501,N_65);
nand U3759 (N_3759,N_1320,N_136);
or U3760 (N_3760,N_2007,N_12);
nand U3761 (N_3761,N_242,N_1276);
or U3762 (N_3762,N_1880,N_845);
or U3763 (N_3763,N_1583,N_697);
or U3764 (N_3764,N_889,N_1428);
nand U3765 (N_3765,N_1698,N_1054);
and U3766 (N_3766,N_436,N_1846);
nand U3767 (N_3767,N_2205,N_2018);
nand U3768 (N_3768,N_1965,N_1244);
nor U3769 (N_3769,N_1343,N_1764);
or U3770 (N_3770,N_628,N_700);
or U3771 (N_3771,N_691,N_1630);
or U3772 (N_3772,N_124,N_404);
nor U3773 (N_3773,N_1683,N_1012);
or U3774 (N_3774,N_354,N_731);
or U3775 (N_3775,N_673,N_1636);
nor U3776 (N_3776,N_246,N_2214);
nand U3777 (N_3777,N_1411,N_1973);
and U3778 (N_3778,N_1385,N_320);
nand U3779 (N_3779,N_247,N_143);
or U3780 (N_3780,N_404,N_1483);
and U3781 (N_3781,N_1155,N_786);
nand U3782 (N_3782,N_583,N_2299);
or U3783 (N_3783,N_1718,N_565);
and U3784 (N_3784,N_1252,N_27);
nand U3785 (N_3785,N_2406,N_338);
or U3786 (N_3786,N_767,N_208);
and U3787 (N_3787,N_1222,N_1016);
nand U3788 (N_3788,N_2129,N_1896);
or U3789 (N_3789,N_487,N_1871);
nand U3790 (N_3790,N_1499,N_1650);
or U3791 (N_3791,N_336,N_324);
nand U3792 (N_3792,N_901,N_1738);
nand U3793 (N_3793,N_1211,N_563);
and U3794 (N_3794,N_95,N_2376);
or U3795 (N_3795,N_2123,N_1149);
and U3796 (N_3796,N_1466,N_1698);
nand U3797 (N_3797,N_2136,N_1158);
nor U3798 (N_3798,N_19,N_2337);
nor U3799 (N_3799,N_1880,N_1164);
nor U3800 (N_3800,N_2203,N_1664);
nand U3801 (N_3801,N_1004,N_1152);
and U3802 (N_3802,N_1544,N_2278);
nand U3803 (N_3803,N_932,N_1008);
nor U3804 (N_3804,N_1359,N_2333);
nor U3805 (N_3805,N_1039,N_2107);
nand U3806 (N_3806,N_1046,N_1742);
nand U3807 (N_3807,N_1811,N_2305);
nor U3808 (N_3808,N_1478,N_895);
nand U3809 (N_3809,N_1263,N_215);
nand U3810 (N_3810,N_1491,N_205);
or U3811 (N_3811,N_1117,N_710);
nor U3812 (N_3812,N_2329,N_2231);
or U3813 (N_3813,N_1682,N_1309);
nand U3814 (N_3814,N_2290,N_2143);
and U3815 (N_3815,N_1071,N_143);
nand U3816 (N_3816,N_1015,N_1033);
or U3817 (N_3817,N_849,N_2227);
or U3818 (N_3818,N_2467,N_974);
nand U3819 (N_3819,N_1386,N_301);
nand U3820 (N_3820,N_612,N_13);
or U3821 (N_3821,N_1974,N_1877);
and U3822 (N_3822,N_108,N_1167);
nand U3823 (N_3823,N_1735,N_2482);
and U3824 (N_3824,N_1992,N_2131);
nand U3825 (N_3825,N_1940,N_820);
nand U3826 (N_3826,N_222,N_1183);
nand U3827 (N_3827,N_2016,N_2318);
and U3828 (N_3828,N_9,N_161);
nand U3829 (N_3829,N_2151,N_174);
and U3830 (N_3830,N_2003,N_1914);
nor U3831 (N_3831,N_482,N_1618);
or U3832 (N_3832,N_2447,N_712);
nand U3833 (N_3833,N_1092,N_669);
nand U3834 (N_3834,N_1176,N_1764);
or U3835 (N_3835,N_485,N_96);
nor U3836 (N_3836,N_551,N_1261);
nor U3837 (N_3837,N_664,N_2479);
and U3838 (N_3838,N_333,N_2193);
nor U3839 (N_3839,N_2054,N_1480);
and U3840 (N_3840,N_1418,N_578);
and U3841 (N_3841,N_1642,N_159);
nor U3842 (N_3842,N_2140,N_1969);
nand U3843 (N_3843,N_2321,N_1174);
and U3844 (N_3844,N_2152,N_2032);
and U3845 (N_3845,N_927,N_898);
and U3846 (N_3846,N_864,N_1407);
or U3847 (N_3847,N_2202,N_1117);
nor U3848 (N_3848,N_2292,N_1216);
and U3849 (N_3849,N_826,N_806);
nor U3850 (N_3850,N_168,N_813);
and U3851 (N_3851,N_1788,N_580);
nor U3852 (N_3852,N_962,N_90);
and U3853 (N_3853,N_876,N_1496);
or U3854 (N_3854,N_533,N_1180);
and U3855 (N_3855,N_784,N_629);
or U3856 (N_3856,N_2332,N_1476);
and U3857 (N_3857,N_1133,N_576);
nand U3858 (N_3858,N_507,N_829);
or U3859 (N_3859,N_345,N_113);
nor U3860 (N_3860,N_1539,N_192);
nand U3861 (N_3861,N_1143,N_2474);
nor U3862 (N_3862,N_533,N_689);
and U3863 (N_3863,N_98,N_2218);
and U3864 (N_3864,N_2469,N_1319);
or U3865 (N_3865,N_60,N_1816);
or U3866 (N_3866,N_975,N_323);
nand U3867 (N_3867,N_1899,N_1498);
nor U3868 (N_3868,N_1134,N_1461);
or U3869 (N_3869,N_1373,N_825);
or U3870 (N_3870,N_2040,N_946);
or U3871 (N_3871,N_1739,N_334);
nor U3872 (N_3872,N_302,N_466);
nand U3873 (N_3873,N_2498,N_2279);
or U3874 (N_3874,N_831,N_1385);
nand U3875 (N_3875,N_199,N_2196);
or U3876 (N_3876,N_148,N_130);
or U3877 (N_3877,N_179,N_2198);
nand U3878 (N_3878,N_166,N_946);
and U3879 (N_3879,N_1376,N_1484);
and U3880 (N_3880,N_793,N_355);
or U3881 (N_3881,N_2498,N_693);
or U3882 (N_3882,N_286,N_2016);
or U3883 (N_3883,N_1838,N_1557);
nor U3884 (N_3884,N_1974,N_1761);
nand U3885 (N_3885,N_9,N_2167);
nand U3886 (N_3886,N_1844,N_1240);
or U3887 (N_3887,N_1724,N_440);
xor U3888 (N_3888,N_1265,N_1097);
nand U3889 (N_3889,N_815,N_1975);
nand U3890 (N_3890,N_1260,N_1484);
or U3891 (N_3891,N_2123,N_110);
nor U3892 (N_3892,N_1507,N_1658);
and U3893 (N_3893,N_1461,N_1634);
or U3894 (N_3894,N_2436,N_1811);
nand U3895 (N_3895,N_1014,N_243);
or U3896 (N_3896,N_1043,N_2240);
or U3897 (N_3897,N_2401,N_1683);
nor U3898 (N_3898,N_816,N_1069);
or U3899 (N_3899,N_1378,N_1661);
and U3900 (N_3900,N_704,N_56);
xnor U3901 (N_3901,N_2080,N_2394);
and U3902 (N_3902,N_1835,N_1070);
nor U3903 (N_3903,N_1670,N_1889);
and U3904 (N_3904,N_1014,N_968);
nor U3905 (N_3905,N_1767,N_1276);
or U3906 (N_3906,N_1347,N_444);
nand U3907 (N_3907,N_1068,N_924);
nor U3908 (N_3908,N_2387,N_193);
and U3909 (N_3909,N_1625,N_195);
nand U3910 (N_3910,N_805,N_214);
nor U3911 (N_3911,N_1561,N_1591);
nand U3912 (N_3912,N_1929,N_1348);
nand U3913 (N_3913,N_1780,N_929);
nand U3914 (N_3914,N_1742,N_197);
or U3915 (N_3915,N_1012,N_1105);
or U3916 (N_3916,N_92,N_2170);
nand U3917 (N_3917,N_2327,N_761);
nand U3918 (N_3918,N_1561,N_1656);
or U3919 (N_3919,N_1313,N_1501);
or U3920 (N_3920,N_443,N_2040);
and U3921 (N_3921,N_188,N_579);
and U3922 (N_3922,N_639,N_68);
nand U3923 (N_3923,N_873,N_2245);
nor U3924 (N_3924,N_739,N_1083);
and U3925 (N_3925,N_1432,N_2344);
nor U3926 (N_3926,N_811,N_1524);
nor U3927 (N_3927,N_268,N_815);
or U3928 (N_3928,N_1452,N_1036);
and U3929 (N_3929,N_2123,N_1181);
and U3930 (N_3930,N_1605,N_200);
nor U3931 (N_3931,N_1715,N_1779);
and U3932 (N_3932,N_2001,N_2065);
nor U3933 (N_3933,N_693,N_119);
and U3934 (N_3934,N_1349,N_1970);
or U3935 (N_3935,N_1070,N_502);
and U3936 (N_3936,N_1501,N_195);
nand U3937 (N_3937,N_1802,N_572);
and U3938 (N_3938,N_1589,N_1663);
nand U3939 (N_3939,N_1693,N_1712);
nand U3940 (N_3940,N_678,N_606);
or U3941 (N_3941,N_2309,N_1245);
nand U3942 (N_3942,N_679,N_286);
and U3943 (N_3943,N_1761,N_813);
and U3944 (N_3944,N_973,N_1417);
nor U3945 (N_3945,N_1892,N_370);
nand U3946 (N_3946,N_2234,N_1652);
and U3947 (N_3947,N_859,N_168);
and U3948 (N_3948,N_648,N_175);
nand U3949 (N_3949,N_2368,N_1412);
nor U3950 (N_3950,N_301,N_1874);
or U3951 (N_3951,N_2119,N_2190);
nor U3952 (N_3952,N_724,N_520);
xnor U3953 (N_3953,N_2296,N_927);
and U3954 (N_3954,N_1706,N_1760);
nor U3955 (N_3955,N_809,N_187);
nand U3956 (N_3956,N_1131,N_1541);
nor U3957 (N_3957,N_1444,N_2354);
or U3958 (N_3958,N_602,N_525);
xor U3959 (N_3959,N_100,N_508);
nor U3960 (N_3960,N_1809,N_2418);
nor U3961 (N_3961,N_1354,N_1960);
or U3962 (N_3962,N_1143,N_2479);
nand U3963 (N_3963,N_906,N_2218);
and U3964 (N_3964,N_1483,N_869);
nand U3965 (N_3965,N_2158,N_1512);
nand U3966 (N_3966,N_1158,N_1829);
and U3967 (N_3967,N_596,N_888);
and U3968 (N_3968,N_791,N_2201);
nand U3969 (N_3969,N_274,N_1486);
nand U3970 (N_3970,N_50,N_814);
and U3971 (N_3971,N_123,N_1200);
and U3972 (N_3972,N_1835,N_731);
and U3973 (N_3973,N_2357,N_911);
nor U3974 (N_3974,N_178,N_634);
and U3975 (N_3975,N_273,N_2404);
nand U3976 (N_3976,N_1791,N_1129);
and U3977 (N_3977,N_2479,N_1865);
nor U3978 (N_3978,N_1697,N_261);
and U3979 (N_3979,N_640,N_853);
and U3980 (N_3980,N_1811,N_2311);
xnor U3981 (N_3981,N_1638,N_1525);
nand U3982 (N_3982,N_2141,N_281);
or U3983 (N_3983,N_1651,N_2145);
and U3984 (N_3984,N_522,N_972);
or U3985 (N_3985,N_364,N_1980);
or U3986 (N_3986,N_900,N_1242);
nor U3987 (N_3987,N_1668,N_1639);
and U3988 (N_3988,N_2186,N_1397);
nor U3989 (N_3989,N_1835,N_1855);
nand U3990 (N_3990,N_1868,N_1919);
and U3991 (N_3991,N_348,N_934);
nor U3992 (N_3992,N_1770,N_1923);
or U3993 (N_3993,N_1550,N_2004);
nor U3994 (N_3994,N_390,N_1032);
nand U3995 (N_3995,N_320,N_1991);
nand U3996 (N_3996,N_2301,N_1944);
nand U3997 (N_3997,N_2197,N_475);
nor U3998 (N_3998,N_756,N_1923);
nor U3999 (N_3999,N_1209,N_268);
or U4000 (N_4000,N_2450,N_969);
and U4001 (N_4001,N_840,N_1784);
nand U4002 (N_4002,N_478,N_2349);
nor U4003 (N_4003,N_2053,N_80);
and U4004 (N_4004,N_2095,N_1161);
xor U4005 (N_4005,N_204,N_523);
nor U4006 (N_4006,N_152,N_2155);
nor U4007 (N_4007,N_1254,N_755);
or U4008 (N_4008,N_1191,N_899);
and U4009 (N_4009,N_618,N_724);
and U4010 (N_4010,N_1277,N_1329);
nor U4011 (N_4011,N_1303,N_1351);
xnor U4012 (N_4012,N_2300,N_2177);
and U4013 (N_4013,N_2269,N_75);
nand U4014 (N_4014,N_1221,N_111);
and U4015 (N_4015,N_1457,N_2110);
nor U4016 (N_4016,N_439,N_512);
xnor U4017 (N_4017,N_1205,N_542);
nand U4018 (N_4018,N_685,N_476);
and U4019 (N_4019,N_22,N_1144);
or U4020 (N_4020,N_940,N_1876);
and U4021 (N_4021,N_822,N_1331);
nor U4022 (N_4022,N_2212,N_462);
or U4023 (N_4023,N_1252,N_686);
nand U4024 (N_4024,N_2488,N_1404);
and U4025 (N_4025,N_273,N_2014);
nor U4026 (N_4026,N_1962,N_1530);
nor U4027 (N_4027,N_2076,N_2214);
nor U4028 (N_4028,N_1887,N_1040);
nand U4029 (N_4029,N_1462,N_17);
or U4030 (N_4030,N_1933,N_1430);
or U4031 (N_4031,N_1066,N_1709);
and U4032 (N_4032,N_1490,N_2361);
and U4033 (N_4033,N_1185,N_858);
or U4034 (N_4034,N_2278,N_979);
or U4035 (N_4035,N_2091,N_645);
nor U4036 (N_4036,N_1049,N_407);
nand U4037 (N_4037,N_762,N_1016);
nor U4038 (N_4038,N_1624,N_1616);
and U4039 (N_4039,N_1,N_1878);
nand U4040 (N_4040,N_1183,N_1640);
nand U4041 (N_4041,N_681,N_2253);
or U4042 (N_4042,N_1406,N_862);
or U4043 (N_4043,N_1795,N_2284);
and U4044 (N_4044,N_1324,N_2042);
and U4045 (N_4045,N_1268,N_1445);
nand U4046 (N_4046,N_1556,N_1157);
and U4047 (N_4047,N_1471,N_2164);
nand U4048 (N_4048,N_1125,N_2437);
and U4049 (N_4049,N_1527,N_2203);
nor U4050 (N_4050,N_2221,N_2476);
nand U4051 (N_4051,N_89,N_2429);
and U4052 (N_4052,N_1950,N_2369);
and U4053 (N_4053,N_1104,N_1508);
or U4054 (N_4054,N_812,N_943);
and U4055 (N_4055,N_1042,N_421);
and U4056 (N_4056,N_713,N_1030);
and U4057 (N_4057,N_1539,N_1320);
nor U4058 (N_4058,N_2336,N_170);
nand U4059 (N_4059,N_2064,N_780);
or U4060 (N_4060,N_764,N_1228);
nand U4061 (N_4061,N_1585,N_1583);
or U4062 (N_4062,N_804,N_60);
nand U4063 (N_4063,N_1114,N_1716);
nor U4064 (N_4064,N_1899,N_1835);
or U4065 (N_4065,N_1232,N_288);
nand U4066 (N_4066,N_1267,N_1845);
or U4067 (N_4067,N_1440,N_637);
or U4068 (N_4068,N_1061,N_1588);
and U4069 (N_4069,N_2454,N_1229);
or U4070 (N_4070,N_1041,N_1798);
and U4071 (N_4071,N_45,N_2243);
nor U4072 (N_4072,N_1438,N_337);
nand U4073 (N_4073,N_1459,N_1249);
nor U4074 (N_4074,N_1879,N_2498);
and U4075 (N_4075,N_1944,N_1572);
nand U4076 (N_4076,N_1222,N_900);
and U4077 (N_4077,N_965,N_1441);
and U4078 (N_4078,N_1376,N_547);
or U4079 (N_4079,N_1788,N_2498);
or U4080 (N_4080,N_2254,N_1741);
nand U4081 (N_4081,N_2310,N_1819);
nor U4082 (N_4082,N_793,N_139);
nand U4083 (N_4083,N_1415,N_378);
and U4084 (N_4084,N_2,N_1211);
or U4085 (N_4085,N_1712,N_2230);
or U4086 (N_4086,N_1402,N_1373);
and U4087 (N_4087,N_1945,N_1768);
or U4088 (N_4088,N_1453,N_1668);
or U4089 (N_4089,N_906,N_396);
or U4090 (N_4090,N_515,N_126);
nor U4091 (N_4091,N_2218,N_558);
and U4092 (N_4092,N_1706,N_2083);
nor U4093 (N_4093,N_130,N_2260);
nor U4094 (N_4094,N_817,N_99);
or U4095 (N_4095,N_805,N_1363);
and U4096 (N_4096,N_1601,N_84);
or U4097 (N_4097,N_1467,N_1640);
and U4098 (N_4098,N_1896,N_1545);
nand U4099 (N_4099,N_2147,N_547);
nor U4100 (N_4100,N_1592,N_2334);
nand U4101 (N_4101,N_503,N_1329);
nor U4102 (N_4102,N_1839,N_1963);
and U4103 (N_4103,N_2204,N_161);
nor U4104 (N_4104,N_680,N_2320);
and U4105 (N_4105,N_496,N_253);
nor U4106 (N_4106,N_1097,N_2048);
and U4107 (N_4107,N_1747,N_1146);
nand U4108 (N_4108,N_1258,N_1035);
or U4109 (N_4109,N_1687,N_220);
nand U4110 (N_4110,N_1844,N_1925);
nand U4111 (N_4111,N_1497,N_439);
and U4112 (N_4112,N_1702,N_1412);
nand U4113 (N_4113,N_2062,N_922);
nor U4114 (N_4114,N_924,N_1985);
nand U4115 (N_4115,N_1172,N_461);
and U4116 (N_4116,N_71,N_1520);
or U4117 (N_4117,N_674,N_1506);
nor U4118 (N_4118,N_880,N_1557);
nor U4119 (N_4119,N_1454,N_2202);
nand U4120 (N_4120,N_2475,N_1672);
nor U4121 (N_4121,N_8,N_2387);
nor U4122 (N_4122,N_1797,N_601);
and U4123 (N_4123,N_2281,N_1538);
and U4124 (N_4124,N_1122,N_1120);
and U4125 (N_4125,N_1859,N_753);
and U4126 (N_4126,N_1354,N_308);
nand U4127 (N_4127,N_132,N_776);
nor U4128 (N_4128,N_402,N_2283);
or U4129 (N_4129,N_2078,N_18);
or U4130 (N_4130,N_1265,N_1034);
nand U4131 (N_4131,N_810,N_867);
and U4132 (N_4132,N_2207,N_1843);
or U4133 (N_4133,N_667,N_1754);
or U4134 (N_4134,N_718,N_524);
nand U4135 (N_4135,N_919,N_859);
nor U4136 (N_4136,N_2213,N_2283);
nor U4137 (N_4137,N_1152,N_2385);
nand U4138 (N_4138,N_2023,N_1528);
nor U4139 (N_4139,N_623,N_2049);
and U4140 (N_4140,N_1110,N_2489);
or U4141 (N_4141,N_2213,N_781);
or U4142 (N_4142,N_1229,N_1628);
nand U4143 (N_4143,N_1657,N_1913);
nor U4144 (N_4144,N_591,N_473);
nand U4145 (N_4145,N_2048,N_378);
nor U4146 (N_4146,N_495,N_602);
and U4147 (N_4147,N_759,N_2295);
and U4148 (N_4148,N_1022,N_461);
nand U4149 (N_4149,N_297,N_1538);
nor U4150 (N_4150,N_1687,N_1859);
or U4151 (N_4151,N_994,N_634);
and U4152 (N_4152,N_1709,N_1967);
nand U4153 (N_4153,N_2331,N_1566);
nand U4154 (N_4154,N_1276,N_1657);
and U4155 (N_4155,N_207,N_285);
nand U4156 (N_4156,N_794,N_1927);
or U4157 (N_4157,N_1471,N_2069);
nor U4158 (N_4158,N_362,N_2142);
nor U4159 (N_4159,N_440,N_1814);
and U4160 (N_4160,N_958,N_1150);
and U4161 (N_4161,N_1666,N_1690);
nand U4162 (N_4162,N_424,N_1459);
and U4163 (N_4163,N_1128,N_1328);
and U4164 (N_4164,N_698,N_973);
nor U4165 (N_4165,N_1790,N_1640);
nand U4166 (N_4166,N_259,N_2397);
and U4167 (N_4167,N_330,N_1276);
nor U4168 (N_4168,N_399,N_234);
or U4169 (N_4169,N_2099,N_1706);
nor U4170 (N_4170,N_2009,N_2058);
nand U4171 (N_4171,N_1861,N_582);
nand U4172 (N_4172,N_1591,N_1831);
nand U4173 (N_4173,N_933,N_1469);
or U4174 (N_4174,N_2121,N_88);
xnor U4175 (N_4175,N_2221,N_551);
nor U4176 (N_4176,N_731,N_322);
nor U4177 (N_4177,N_1839,N_393);
nor U4178 (N_4178,N_112,N_1112);
nand U4179 (N_4179,N_2395,N_1609);
nand U4180 (N_4180,N_1663,N_518);
nand U4181 (N_4181,N_616,N_190);
nor U4182 (N_4182,N_1327,N_2340);
and U4183 (N_4183,N_955,N_104);
or U4184 (N_4184,N_2110,N_13);
and U4185 (N_4185,N_1287,N_2006);
or U4186 (N_4186,N_2005,N_1039);
or U4187 (N_4187,N_2296,N_88);
and U4188 (N_4188,N_596,N_1839);
or U4189 (N_4189,N_1703,N_1801);
or U4190 (N_4190,N_820,N_2333);
nand U4191 (N_4191,N_2123,N_543);
and U4192 (N_4192,N_23,N_503);
nor U4193 (N_4193,N_544,N_1752);
nand U4194 (N_4194,N_2050,N_649);
or U4195 (N_4195,N_950,N_1929);
xor U4196 (N_4196,N_2013,N_1496);
and U4197 (N_4197,N_794,N_900);
nand U4198 (N_4198,N_1489,N_494);
and U4199 (N_4199,N_2216,N_1446);
or U4200 (N_4200,N_410,N_741);
nor U4201 (N_4201,N_462,N_412);
nand U4202 (N_4202,N_1075,N_900);
nand U4203 (N_4203,N_125,N_2139);
nand U4204 (N_4204,N_1666,N_864);
or U4205 (N_4205,N_421,N_655);
nand U4206 (N_4206,N_958,N_648);
and U4207 (N_4207,N_1861,N_42);
xnor U4208 (N_4208,N_123,N_1848);
and U4209 (N_4209,N_681,N_682);
or U4210 (N_4210,N_10,N_1744);
nand U4211 (N_4211,N_2274,N_48);
nor U4212 (N_4212,N_812,N_1804);
nand U4213 (N_4213,N_496,N_1203);
or U4214 (N_4214,N_266,N_1242);
nand U4215 (N_4215,N_873,N_482);
and U4216 (N_4216,N_2491,N_1670);
nand U4217 (N_4217,N_1732,N_1536);
and U4218 (N_4218,N_1934,N_1884);
nand U4219 (N_4219,N_2263,N_431);
nand U4220 (N_4220,N_1340,N_1113);
nor U4221 (N_4221,N_545,N_1327);
nor U4222 (N_4222,N_2072,N_2236);
and U4223 (N_4223,N_1001,N_296);
nand U4224 (N_4224,N_1918,N_1676);
or U4225 (N_4225,N_69,N_1962);
nor U4226 (N_4226,N_161,N_755);
nor U4227 (N_4227,N_1051,N_736);
nand U4228 (N_4228,N_1654,N_2300);
nand U4229 (N_4229,N_1048,N_1356);
and U4230 (N_4230,N_345,N_285);
nand U4231 (N_4231,N_536,N_453);
or U4232 (N_4232,N_1051,N_404);
nor U4233 (N_4233,N_618,N_1561);
and U4234 (N_4234,N_2278,N_1720);
or U4235 (N_4235,N_2228,N_611);
or U4236 (N_4236,N_528,N_1778);
or U4237 (N_4237,N_635,N_782);
nor U4238 (N_4238,N_2370,N_1193);
nor U4239 (N_4239,N_2261,N_1378);
or U4240 (N_4240,N_607,N_2360);
nand U4241 (N_4241,N_2018,N_1901);
nand U4242 (N_4242,N_1805,N_200);
or U4243 (N_4243,N_1004,N_726);
or U4244 (N_4244,N_1239,N_1702);
or U4245 (N_4245,N_1314,N_1478);
nor U4246 (N_4246,N_2333,N_2286);
nand U4247 (N_4247,N_1579,N_1150);
or U4248 (N_4248,N_888,N_496);
nor U4249 (N_4249,N_836,N_2334);
nor U4250 (N_4250,N_1417,N_566);
or U4251 (N_4251,N_1809,N_1615);
nor U4252 (N_4252,N_1753,N_720);
and U4253 (N_4253,N_2366,N_1371);
and U4254 (N_4254,N_491,N_876);
nand U4255 (N_4255,N_735,N_631);
nand U4256 (N_4256,N_783,N_980);
nor U4257 (N_4257,N_1882,N_1050);
nand U4258 (N_4258,N_1480,N_993);
nor U4259 (N_4259,N_886,N_620);
nand U4260 (N_4260,N_151,N_2064);
and U4261 (N_4261,N_1928,N_1299);
or U4262 (N_4262,N_1966,N_2112);
nand U4263 (N_4263,N_2225,N_1797);
nor U4264 (N_4264,N_1753,N_387);
nor U4265 (N_4265,N_1577,N_377);
or U4266 (N_4266,N_48,N_2353);
or U4267 (N_4267,N_882,N_700);
or U4268 (N_4268,N_496,N_2421);
nand U4269 (N_4269,N_2073,N_1201);
nor U4270 (N_4270,N_1847,N_2397);
nor U4271 (N_4271,N_547,N_1126);
nand U4272 (N_4272,N_1497,N_2260);
xor U4273 (N_4273,N_1956,N_1856);
or U4274 (N_4274,N_385,N_1073);
nor U4275 (N_4275,N_1532,N_2137);
nand U4276 (N_4276,N_1814,N_661);
and U4277 (N_4277,N_1763,N_209);
xor U4278 (N_4278,N_1829,N_1868);
or U4279 (N_4279,N_852,N_1527);
nor U4280 (N_4280,N_1355,N_450);
and U4281 (N_4281,N_937,N_843);
nand U4282 (N_4282,N_255,N_2246);
and U4283 (N_4283,N_435,N_1645);
or U4284 (N_4284,N_1682,N_1399);
or U4285 (N_4285,N_704,N_458);
nand U4286 (N_4286,N_42,N_543);
nand U4287 (N_4287,N_999,N_2118);
nor U4288 (N_4288,N_108,N_1044);
nor U4289 (N_4289,N_649,N_2277);
nor U4290 (N_4290,N_1420,N_2419);
or U4291 (N_4291,N_159,N_177);
or U4292 (N_4292,N_2006,N_1821);
nand U4293 (N_4293,N_2452,N_2154);
nand U4294 (N_4294,N_1830,N_2339);
or U4295 (N_4295,N_2050,N_643);
or U4296 (N_4296,N_2381,N_2316);
nor U4297 (N_4297,N_2151,N_1252);
nor U4298 (N_4298,N_187,N_2274);
nor U4299 (N_4299,N_1643,N_1711);
xnor U4300 (N_4300,N_995,N_594);
nor U4301 (N_4301,N_707,N_1110);
nand U4302 (N_4302,N_1305,N_1635);
or U4303 (N_4303,N_1516,N_1621);
or U4304 (N_4304,N_1213,N_1160);
or U4305 (N_4305,N_1182,N_1749);
nor U4306 (N_4306,N_16,N_2256);
nand U4307 (N_4307,N_1174,N_1051);
nand U4308 (N_4308,N_1327,N_1113);
nor U4309 (N_4309,N_884,N_242);
nand U4310 (N_4310,N_1185,N_745);
nand U4311 (N_4311,N_42,N_2461);
and U4312 (N_4312,N_1199,N_342);
nor U4313 (N_4313,N_1798,N_1539);
nand U4314 (N_4314,N_715,N_979);
or U4315 (N_4315,N_314,N_348);
and U4316 (N_4316,N_1950,N_753);
nor U4317 (N_4317,N_1645,N_249);
and U4318 (N_4318,N_2455,N_1748);
nor U4319 (N_4319,N_2267,N_593);
nor U4320 (N_4320,N_1556,N_878);
nor U4321 (N_4321,N_643,N_2175);
and U4322 (N_4322,N_205,N_1747);
nor U4323 (N_4323,N_1910,N_835);
and U4324 (N_4324,N_1578,N_288);
or U4325 (N_4325,N_618,N_1346);
nor U4326 (N_4326,N_1400,N_130);
nand U4327 (N_4327,N_307,N_639);
or U4328 (N_4328,N_370,N_1789);
or U4329 (N_4329,N_20,N_803);
and U4330 (N_4330,N_1671,N_818);
nand U4331 (N_4331,N_1988,N_1576);
and U4332 (N_4332,N_403,N_722);
nor U4333 (N_4333,N_2193,N_2184);
nand U4334 (N_4334,N_2,N_1155);
nand U4335 (N_4335,N_266,N_634);
nor U4336 (N_4336,N_706,N_811);
nand U4337 (N_4337,N_536,N_2047);
or U4338 (N_4338,N_1871,N_671);
or U4339 (N_4339,N_1507,N_432);
nand U4340 (N_4340,N_928,N_389);
nand U4341 (N_4341,N_1174,N_578);
nand U4342 (N_4342,N_1303,N_1370);
nor U4343 (N_4343,N_2232,N_1433);
nor U4344 (N_4344,N_1240,N_931);
xor U4345 (N_4345,N_251,N_1479);
and U4346 (N_4346,N_2308,N_633);
or U4347 (N_4347,N_2423,N_2080);
or U4348 (N_4348,N_1998,N_1186);
and U4349 (N_4349,N_2145,N_536);
and U4350 (N_4350,N_692,N_1811);
nor U4351 (N_4351,N_1419,N_2202);
nor U4352 (N_4352,N_425,N_1188);
or U4353 (N_4353,N_2351,N_2321);
or U4354 (N_4354,N_2081,N_828);
or U4355 (N_4355,N_1535,N_1449);
nor U4356 (N_4356,N_223,N_2097);
or U4357 (N_4357,N_106,N_2145);
nor U4358 (N_4358,N_472,N_2275);
nand U4359 (N_4359,N_81,N_1422);
or U4360 (N_4360,N_110,N_995);
and U4361 (N_4361,N_2440,N_1329);
nor U4362 (N_4362,N_342,N_2189);
or U4363 (N_4363,N_1656,N_586);
nand U4364 (N_4364,N_1233,N_1951);
or U4365 (N_4365,N_241,N_1093);
nand U4366 (N_4366,N_1588,N_1331);
or U4367 (N_4367,N_1551,N_2446);
and U4368 (N_4368,N_2045,N_50);
nor U4369 (N_4369,N_807,N_2239);
nand U4370 (N_4370,N_1762,N_361);
nor U4371 (N_4371,N_776,N_2185);
and U4372 (N_4372,N_1796,N_1458);
or U4373 (N_4373,N_1369,N_157);
xnor U4374 (N_4374,N_2443,N_1902);
xor U4375 (N_4375,N_48,N_1528);
nor U4376 (N_4376,N_1867,N_2321);
nand U4377 (N_4377,N_445,N_2357);
nand U4378 (N_4378,N_1424,N_2435);
or U4379 (N_4379,N_685,N_1445);
and U4380 (N_4380,N_2113,N_1793);
nor U4381 (N_4381,N_1511,N_1092);
nor U4382 (N_4382,N_1767,N_1733);
or U4383 (N_4383,N_2439,N_481);
nor U4384 (N_4384,N_434,N_1124);
or U4385 (N_4385,N_1926,N_94);
nand U4386 (N_4386,N_1167,N_110);
and U4387 (N_4387,N_1421,N_1052);
and U4388 (N_4388,N_467,N_1724);
nand U4389 (N_4389,N_2491,N_991);
and U4390 (N_4390,N_1897,N_526);
nand U4391 (N_4391,N_1414,N_1960);
nand U4392 (N_4392,N_366,N_93);
and U4393 (N_4393,N_1027,N_617);
and U4394 (N_4394,N_1085,N_201);
or U4395 (N_4395,N_1912,N_802);
nor U4396 (N_4396,N_131,N_814);
and U4397 (N_4397,N_2314,N_1661);
or U4398 (N_4398,N_2457,N_823);
or U4399 (N_4399,N_387,N_1051);
xnor U4400 (N_4400,N_1888,N_1934);
and U4401 (N_4401,N_567,N_684);
nor U4402 (N_4402,N_1261,N_2169);
nor U4403 (N_4403,N_337,N_257);
xnor U4404 (N_4404,N_1919,N_379);
nand U4405 (N_4405,N_449,N_1719);
or U4406 (N_4406,N_1187,N_201);
nand U4407 (N_4407,N_786,N_611);
xnor U4408 (N_4408,N_1586,N_1938);
or U4409 (N_4409,N_429,N_1132);
and U4410 (N_4410,N_2304,N_1773);
and U4411 (N_4411,N_1888,N_763);
or U4412 (N_4412,N_2424,N_1747);
nor U4413 (N_4413,N_1903,N_1513);
nand U4414 (N_4414,N_417,N_1252);
and U4415 (N_4415,N_1471,N_824);
nand U4416 (N_4416,N_279,N_1224);
nor U4417 (N_4417,N_709,N_213);
nand U4418 (N_4418,N_2021,N_2103);
xor U4419 (N_4419,N_384,N_1171);
and U4420 (N_4420,N_1587,N_532);
and U4421 (N_4421,N_1108,N_126);
nor U4422 (N_4422,N_2326,N_1327);
or U4423 (N_4423,N_834,N_2180);
or U4424 (N_4424,N_1954,N_1007);
or U4425 (N_4425,N_2251,N_1246);
nand U4426 (N_4426,N_2030,N_2337);
nand U4427 (N_4427,N_826,N_1239);
nand U4428 (N_4428,N_1716,N_2281);
nand U4429 (N_4429,N_688,N_1977);
nor U4430 (N_4430,N_1177,N_1538);
nand U4431 (N_4431,N_2425,N_101);
and U4432 (N_4432,N_1131,N_156);
or U4433 (N_4433,N_873,N_1210);
nand U4434 (N_4434,N_1698,N_952);
nand U4435 (N_4435,N_1056,N_422);
nand U4436 (N_4436,N_1065,N_1428);
nand U4437 (N_4437,N_1577,N_2405);
nand U4438 (N_4438,N_972,N_1787);
nand U4439 (N_4439,N_1102,N_857);
nand U4440 (N_4440,N_1819,N_1294);
nand U4441 (N_4441,N_2036,N_464);
and U4442 (N_4442,N_1009,N_1720);
or U4443 (N_4443,N_110,N_1482);
and U4444 (N_4444,N_1277,N_810);
nor U4445 (N_4445,N_1962,N_879);
and U4446 (N_4446,N_647,N_677);
nor U4447 (N_4447,N_2016,N_1978);
or U4448 (N_4448,N_262,N_2049);
nor U4449 (N_4449,N_2283,N_391);
nor U4450 (N_4450,N_539,N_526);
or U4451 (N_4451,N_373,N_2069);
nand U4452 (N_4452,N_2359,N_571);
and U4453 (N_4453,N_2478,N_534);
and U4454 (N_4454,N_2074,N_58);
or U4455 (N_4455,N_409,N_1870);
nor U4456 (N_4456,N_2146,N_2450);
or U4457 (N_4457,N_1956,N_1118);
or U4458 (N_4458,N_868,N_42);
nor U4459 (N_4459,N_320,N_613);
or U4460 (N_4460,N_716,N_1889);
or U4461 (N_4461,N_1791,N_693);
xor U4462 (N_4462,N_2300,N_761);
nor U4463 (N_4463,N_837,N_409);
nor U4464 (N_4464,N_632,N_751);
and U4465 (N_4465,N_477,N_372);
nor U4466 (N_4466,N_1279,N_2377);
or U4467 (N_4467,N_489,N_340);
nor U4468 (N_4468,N_874,N_1411);
nor U4469 (N_4469,N_865,N_2408);
nand U4470 (N_4470,N_1209,N_1768);
nor U4471 (N_4471,N_2448,N_1712);
nand U4472 (N_4472,N_138,N_543);
or U4473 (N_4473,N_658,N_393);
or U4474 (N_4474,N_105,N_1253);
and U4475 (N_4475,N_2032,N_2145);
nand U4476 (N_4476,N_2444,N_690);
nand U4477 (N_4477,N_2387,N_2237);
or U4478 (N_4478,N_1249,N_1445);
or U4479 (N_4479,N_221,N_2302);
nor U4480 (N_4480,N_1762,N_2099);
or U4481 (N_4481,N_6,N_1434);
or U4482 (N_4482,N_1547,N_1774);
nand U4483 (N_4483,N_2206,N_2046);
and U4484 (N_4484,N_1216,N_1703);
or U4485 (N_4485,N_2091,N_2013);
and U4486 (N_4486,N_1202,N_2197);
nor U4487 (N_4487,N_1495,N_1416);
nor U4488 (N_4488,N_1607,N_2449);
and U4489 (N_4489,N_1993,N_58);
or U4490 (N_4490,N_2432,N_1351);
and U4491 (N_4491,N_198,N_138);
nor U4492 (N_4492,N_874,N_2204);
nor U4493 (N_4493,N_1322,N_1952);
nor U4494 (N_4494,N_409,N_476);
and U4495 (N_4495,N_849,N_2300);
or U4496 (N_4496,N_1308,N_1231);
or U4497 (N_4497,N_309,N_352);
and U4498 (N_4498,N_574,N_228);
xor U4499 (N_4499,N_1937,N_1874);
nor U4500 (N_4500,N_1832,N_1732);
and U4501 (N_4501,N_1026,N_78);
or U4502 (N_4502,N_896,N_1832);
nor U4503 (N_4503,N_1015,N_1031);
and U4504 (N_4504,N_2389,N_1741);
and U4505 (N_4505,N_353,N_2208);
and U4506 (N_4506,N_247,N_1004);
or U4507 (N_4507,N_74,N_1118);
nand U4508 (N_4508,N_1934,N_1834);
nor U4509 (N_4509,N_1333,N_744);
or U4510 (N_4510,N_1012,N_2112);
nor U4511 (N_4511,N_1456,N_874);
and U4512 (N_4512,N_36,N_2485);
nand U4513 (N_4513,N_1441,N_176);
nor U4514 (N_4514,N_2386,N_50);
or U4515 (N_4515,N_963,N_2178);
nand U4516 (N_4516,N_1975,N_654);
xnor U4517 (N_4517,N_45,N_520);
or U4518 (N_4518,N_2136,N_1487);
and U4519 (N_4519,N_1000,N_1143);
xnor U4520 (N_4520,N_365,N_1808);
and U4521 (N_4521,N_771,N_2167);
nand U4522 (N_4522,N_1609,N_1983);
nand U4523 (N_4523,N_1715,N_436);
nand U4524 (N_4524,N_1976,N_1678);
or U4525 (N_4525,N_2352,N_93);
nand U4526 (N_4526,N_562,N_1319);
nand U4527 (N_4527,N_397,N_954);
or U4528 (N_4528,N_1444,N_326);
or U4529 (N_4529,N_957,N_2033);
nand U4530 (N_4530,N_831,N_555);
nand U4531 (N_4531,N_665,N_793);
or U4532 (N_4532,N_1410,N_3);
nor U4533 (N_4533,N_1297,N_62);
nor U4534 (N_4534,N_1350,N_1397);
and U4535 (N_4535,N_767,N_576);
or U4536 (N_4536,N_248,N_1694);
nor U4537 (N_4537,N_1559,N_1755);
or U4538 (N_4538,N_685,N_824);
and U4539 (N_4539,N_1394,N_2352);
and U4540 (N_4540,N_2480,N_1014);
nor U4541 (N_4541,N_740,N_1913);
nor U4542 (N_4542,N_202,N_2460);
or U4543 (N_4543,N_471,N_1394);
or U4544 (N_4544,N_2111,N_1669);
nand U4545 (N_4545,N_310,N_919);
or U4546 (N_4546,N_1405,N_983);
or U4547 (N_4547,N_2269,N_525);
and U4548 (N_4548,N_312,N_1844);
nor U4549 (N_4549,N_2122,N_1182);
or U4550 (N_4550,N_364,N_2427);
nand U4551 (N_4551,N_2149,N_1049);
and U4552 (N_4552,N_2446,N_131);
nand U4553 (N_4553,N_473,N_1049);
nand U4554 (N_4554,N_2222,N_2247);
and U4555 (N_4555,N_144,N_2364);
nand U4556 (N_4556,N_1434,N_1237);
or U4557 (N_4557,N_1989,N_1254);
nand U4558 (N_4558,N_139,N_32);
nand U4559 (N_4559,N_1044,N_804);
or U4560 (N_4560,N_1461,N_1089);
and U4561 (N_4561,N_1520,N_73);
and U4562 (N_4562,N_568,N_750);
and U4563 (N_4563,N_266,N_713);
nand U4564 (N_4564,N_1083,N_373);
nor U4565 (N_4565,N_2195,N_1685);
nor U4566 (N_4566,N_313,N_2478);
nor U4567 (N_4567,N_1791,N_1087);
and U4568 (N_4568,N_2308,N_1660);
nor U4569 (N_4569,N_2390,N_1924);
nor U4570 (N_4570,N_1061,N_99);
or U4571 (N_4571,N_1495,N_326);
and U4572 (N_4572,N_993,N_2213);
and U4573 (N_4573,N_1820,N_210);
or U4574 (N_4574,N_1452,N_2273);
nand U4575 (N_4575,N_1454,N_729);
nor U4576 (N_4576,N_1801,N_1205);
nor U4577 (N_4577,N_917,N_478);
nand U4578 (N_4578,N_64,N_178);
nor U4579 (N_4579,N_1221,N_2278);
xor U4580 (N_4580,N_1206,N_1765);
nand U4581 (N_4581,N_2359,N_114);
and U4582 (N_4582,N_483,N_978);
nor U4583 (N_4583,N_27,N_2199);
and U4584 (N_4584,N_2379,N_334);
nor U4585 (N_4585,N_96,N_409);
or U4586 (N_4586,N_1318,N_230);
or U4587 (N_4587,N_1741,N_947);
nand U4588 (N_4588,N_2178,N_1508);
nand U4589 (N_4589,N_1941,N_211);
or U4590 (N_4590,N_115,N_1356);
nand U4591 (N_4591,N_518,N_1753);
nand U4592 (N_4592,N_212,N_1554);
nor U4593 (N_4593,N_570,N_1273);
or U4594 (N_4594,N_1171,N_1568);
and U4595 (N_4595,N_220,N_504);
or U4596 (N_4596,N_1803,N_632);
or U4597 (N_4597,N_741,N_307);
nand U4598 (N_4598,N_857,N_1881);
or U4599 (N_4599,N_974,N_1399);
and U4600 (N_4600,N_730,N_200);
nor U4601 (N_4601,N_464,N_778);
nor U4602 (N_4602,N_2134,N_1757);
and U4603 (N_4603,N_641,N_1039);
nor U4604 (N_4604,N_1290,N_1328);
nor U4605 (N_4605,N_2480,N_342);
nand U4606 (N_4606,N_877,N_2311);
or U4607 (N_4607,N_1448,N_535);
nand U4608 (N_4608,N_330,N_1697);
nand U4609 (N_4609,N_550,N_2463);
nor U4610 (N_4610,N_752,N_352);
or U4611 (N_4611,N_804,N_1385);
nand U4612 (N_4612,N_1243,N_1596);
nor U4613 (N_4613,N_2043,N_192);
nor U4614 (N_4614,N_1036,N_731);
nand U4615 (N_4615,N_1641,N_1765);
and U4616 (N_4616,N_1975,N_206);
xor U4617 (N_4617,N_1153,N_1938);
nor U4618 (N_4618,N_2242,N_2333);
and U4619 (N_4619,N_1402,N_287);
nand U4620 (N_4620,N_1718,N_410);
or U4621 (N_4621,N_1981,N_710);
nor U4622 (N_4622,N_2463,N_1916);
and U4623 (N_4623,N_1660,N_1444);
and U4624 (N_4624,N_818,N_1209);
nor U4625 (N_4625,N_1831,N_12);
nor U4626 (N_4626,N_586,N_1419);
or U4627 (N_4627,N_902,N_264);
nor U4628 (N_4628,N_1025,N_837);
nor U4629 (N_4629,N_760,N_2005);
or U4630 (N_4630,N_481,N_983);
and U4631 (N_4631,N_53,N_689);
nor U4632 (N_4632,N_2464,N_1341);
nor U4633 (N_4633,N_2463,N_1063);
nand U4634 (N_4634,N_2304,N_1341);
and U4635 (N_4635,N_664,N_2169);
or U4636 (N_4636,N_1081,N_1830);
nand U4637 (N_4637,N_1620,N_1299);
and U4638 (N_4638,N_2285,N_2485);
or U4639 (N_4639,N_1903,N_1272);
or U4640 (N_4640,N_897,N_1341);
nor U4641 (N_4641,N_2496,N_643);
nor U4642 (N_4642,N_705,N_2206);
nor U4643 (N_4643,N_311,N_1532);
nor U4644 (N_4644,N_499,N_1633);
nand U4645 (N_4645,N_1288,N_1465);
nor U4646 (N_4646,N_372,N_2105);
nand U4647 (N_4647,N_1436,N_1506);
or U4648 (N_4648,N_1596,N_2434);
nand U4649 (N_4649,N_191,N_539);
and U4650 (N_4650,N_1931,N_1653);
nand U4651 (N_4651,N_317,N_1858);
nor U4652 (N_4652,N_503,N_734);
nor U4653 (N_4653,N_1362,N_770);
nor U4654 (N_4654,N_931,N_750);
or U4655 (N_4655,N_1053,N_1706);
and U4656 (N_4656,N_200,N_507);
and U4657 (N_4657,N_2089,N_1004);
nand U4658 (N_4658,N_1807,N_2151);
and U4659 (N_4659,N_144,N_1794);
or U4660 (N_4660,N_2366,N_1139);
nor U4661 (N_4661,N_1204,N_1525);
nand U4662 (N_4662,N_1996,N_309);
nor U4663 (N_4663,N_2197,N_426);
nor U4664 (N_4664,N_1812,N_1085);
or U4665 (N_4665,N_1929,N_1753);
and U4666 (N_4666,N_1046,N_1694);
or U4667 (N_4667,N_1719,N_397);
nor U4668 (N_4668,N_1181,N_1488);
nor U4669 (N_4669,N_2277,N_206);
nand U4670 (N_4670,N_2354,N_507);
and U4671 (N_4671,N_301,N_1699);
or U4672 (N_4672,N_1115,N_1509);
or U4673 (N_4673,N_1947,N_705);
nor U4674 (N_4674,N_1907,N_2114);
nor U4675 (N_4675,N_552,N_1126);
nor U4676 (N_4676,N_2368,N_978);
nand U4677 (N_4677,N_1257,N_2218);
and U4678 (N_4678,N_1953,N_2075);
and U4679 (N_4679,N_1687,N_1169);
nand U4680 (N_4680,N_1324,N_684);
nand U4681 (N_4681,N_705,N_1478);
nand U4682 (N_4682,N_748,N_1990);
and U4683 (N_4683,N_752,N_421);
or U4684 (N_4684,N_1288,N_1036);
and U4685 (N_4685,N_867,N_180);
or U4686 (N_4686,N_175,N_228);
or U4687 (N_4687,N_996,N_427);
nand U4688 (N_4688,N_565,N_1366);
nor U4689 (N_4689,N_1310,N_2433);
or U4690 (N_4690,N_1036,N_814);
and U4691 (N_4691,N_2184,N_2030);
or U4692 (N_4692,N_831,N_1658);
or U4693 (N_4693,N_1216,N_2397);
nand U4694 (N_4694,N_530,N_2260);
nand U4695 (N_4695,N_1711,N_630);
or U4696 (N_4696,N_513,N_1633);
nor U4697 (N_4697,N_428,N_202);
xor U4698 (N_4698,N_150,N_1369);
nand U4699 (N_4699,N_2003,N_2026);
or U4700 (N_4700,N_1405,N_1295);
nor U4701 (N_4701,N_707,N_656);
or U4702 (N_4702,N_2107,N_956);
and U4703 (N_4703,N_1727,N_1561);
nand U4704 (N_4704,N_612,N_703);
nand U4705 (N_4705,N_1947,N_150);
and U4706 (N_4706,N_1722,N_1182);
and U4707 (N_4707,N_273,N_2281);
or U4708 (N_4708,N_603,N_1576);
nand U4709 (N_4709,N_1194,N_1090);
nand U4710 (N_4710,N_694,N_1769);
or U4711 (N_4711,N_1039,N_1738);
or U4712 (N_4712,N_1203,N_1510);
nand U4713 (N_4713,N_325,N_522);
and U4714 (N_4714,N_1020,N_2228);
nand U4715 (N_4715,N_1928,N_2076);
or U4716 (N_4716,N_1926,N_2289);
and U4717 (N_4717,N_1415,N_8);
or U4718 (N_4718,N_1391,N_1191);
nand U4719 (N_4719,N_2355,N_1239);
nand U4720 (N_4720,N_2460,N_2026);
or U4721 (N_4721,N_2144,N_2074);
and U4722 (N_4722,N_1401,N_232);
nor U4723 (N_4723,N_123,N_864);
or U4724 (N_4724,N_960,N_161);
and U4725 (N_4725,N_2163,N_1629);
nor U4726 (N_4726,N_64,N_877);
or U4727 (N_4727,N_2130,N_2003);
or U4728 (N_4728,N_592,N_540);
nor U4729 (N_4729,N_2309,N_2412);
nand U4730 (N_4730,N_2185,N_716);
and U4731 (N_4731,N_541,N_1944);
and U4732 (N_4732,N_449,N_878);
and U4733 (N_4733,N_1770,N_1204);
nor U4734 (N_4734,N_681,N_1434);
nand U4735 (N_4735,N_1531,N_729);
and U4736 (N_4736,N_900,N_517);
or U4737 (N_4737,N_2199,N_696);
nor U4738 (N_4738,N_1121,N_1219);
nand U4739 (N_4739,N_225,N_529);
nor U4740 (N_4740,N_1455,N_1876);
nand U4741 (N_4741,N_1493,N_1441);
nand U4742 (N_4742,N_617,N_536);
nand U4743 (N_4743,N_1364,N_1211);
or U4744 (N_4744,N_2290,N_83);
or U4745 (N_4745,N_1565,N_1706);
or U4746 (N_4746,N_659,N_1348);
nor U4747 (N_4747,N_1521,N_2081);
nor U4748 (N_4748,N_944,N_1739);
or U4749 (N_4749,N_1327,N_660);
nor U4750 (N_4750,N_802,N_628);
and U4751 (N_4751,N_1795,N_568);
or U4752 (N_4752,N_2405,N_1477);
and U4753 (N_4753,N_1921,N_785);
nor U4754 (N_4754,N_1429,N_506);
or U4755 (N_4755,N_339,N_687);
or U4756 (N_4756,N_1433,N_1386);
and U4757 (N_4757,N_369,N_93);
and U4758 (N_4758,N_1517,N_1308);
and U4759 (N_4759,N_586,N_2372);
nand U4760 (N_4760,N_1395,N_1548);
or U4761 (N_4761,N_137,N_2197);
or U4762 (N_4762,N_835,N_1036);
or U4763 (N_4763,N_1207,N_1187);
or U4764 (N_4764,N_1795,N_331);
nor U4765 (N_4765,N_53,N_2294);
and U4766 (N_4766,N_1420,N_2102);
nor U4767 (N_4767,N_713,N_2211);
or U4768 (N_4768,N_156,N_1243);
and U4769 (N_4769,N_715,N_2171);
and U4770 (N_4770,N_797,N_617);
or U4771 (N_4771,N_571,N_809);
nor U4772 (N_4772,N_2435,N_10);
or U4773 (N_4773,N_237,N_800);
nand U4774 (N_4774,N_415,N_2405);
nand U4775 (N_4775,N_15,N_1274);
or U4776 (N_4776,N_1332,N_1799);
or U4777 (N_4777,N_263,N_1198);
and U4778 (N_4778,N_2338,N_1617);
nor U4779 (N_4779,N_990,N_1572);
nor U4780 (N_4780,N_1218,N_1117);
nor U4781 (N_4781,N_1287,N_1955);
and U4782 (N_4782,N_2246,N_1219);
xnor U4783 (N_4783,N_1592,N_786);
or U4784 (N_4784,N_553,N_996);
and U4785 (N_4785,N_606,N_2388);
nand U4786 (N_4786,N_186,N_1438);
nand U4787 (N_4787,N_725,N_574);
nand U4788 (N_4788,N_826,N_948);
nor U4789 (N_4789,N_756,N_1285);
or U4790 (N_4790,N_1841,N_1681);
and U4791 (N_4791,N_330,N_1076);
or U4792 (N_4792,N_364,N_1376);
and U4793 (N_4793,N_1640,N_504);
nor U4794 (N_4794,N_798,N_741);
nor U4795 (N_4795,N_561,N_671);
and U4796 (N_4796,N_1476,N_659);
nand U4797 (N_4797,N_1303,N_2364);
and U4798 (N_4798,N_525,N_1223);
nand U4799 (N_4799,N_1932,N_1326);
nor U4800 (N_4800,N_422,N_102);
nor U4801 (N_4801,N_1062,N_2022);
or U4802 (N_4802,N_1698,N_1583);
and U4803 (N_4803,N_2428,N_2245);
nor U4804 (N_4804,N_2199,N_137);
nor U4805 (N_4805,N_678,N_1007);
and U4806 (N_4806,N_2361,N_586);
nor U4807 (N_4807,N_660,N_483);
nand U4808 (N_4808,N_1466,N_507);
nand U4809 (N_4809,N_2382,N_907);
nand U4810 (N_4810,N_1373,N_861);
and U4811 (N_4811,N_1101,N_2002);
nand U4812 (N_4812,N_1829,N_818);
and U4813 (N_4813,N_2215,N_516);
and U4814 (N_4814,N_1208,N_1756);
nor U4815 (N_4815,N_1602,N_465);
or U4816 (N_4816,N_659,N_1378);
xnor U4817 (N_4817,N_2013,N_1907);
nand U4818 (N_4818,N_1283,N_218);
xor U4819 (N_4819,N_1306,N_1708);
nor U4820 (N_4820,N_1686,N_2476);
nor U4821 (N_4821,N_1866,N_1084);
nor U4822 (N_4822,N_836,N_309);
and U4823 (N_4823,N_1170,N_1806);
or U4824 (N_4824,N_598,N_853);
and U4825 (N_4825,N_600,N_1998);
or U4826 (N_4826,N_2451,N_160);
or U4827 (N_4827,N_484,N_1665);
nor U4828 (N_4828,N_2170,N_2372);
or U4829 (N_4829,N_814,N_2137);
or U4830 (N_4830,N_760,N_1365);
and U4831 (N_4831,N_42,N_539);
and U4832 (N_4832,N_1996,N_2139);
or U4833 (N_4833,N_14,N_1517);
nor U4834 (N_4834,N_92,N_2287);
xor U4835 (N_4835,N_1687,N_1332);
nand U4836 (N_4836,N_1826,N_429);
and U4837 (N_4837,N_53,N_2100);
or U4838 (N_4838,N_2368,N_1103);
or U4839 (N_4839,N_1019,N_585);
nor U4840 (N_4840,N_1505,N_1578);
nand U4841 (N_4841,N_1174,N_1359);
and U4842 (N_4842,N_985,N_2084);
nor U4843 (N_4843,N_231,N_418);
and U4844 (N_4844,N_343,N_1328);
and U4845 (N_4845,N_597,N_2245);
nand U4846 (N_4846,N_670,N_2068);
nor U4847 (N_4847,N_939,N_618);
nor U4848 (N_4848,N_1800,N_1323);
and U4849 (N_4849,N_947,N_2215);
xor U4850 (N_4850,N_1048,N_190);
xor U4851 (N_4851,N_178,N_987);
or U4852 (N_4852,N_2381,N_1103);
and U4853 (N_4853,N_9,N_2004);
or U4854 (N_4854,N_1872,N_620);
nor U4855 (N_4855,N_1473,N_1045);
and U4856 (N_4856,N_516,N_1641);
and U4857 (N_4857,N_2411,N_926);
nand U4858 (N_4858,N_866,N_1250);
and U4859 (N_4859,N_1404,N_192);
nor U4860 (N_4860,N_1484,N_1916);
or U4861 (N_4861,N_1443,N_1773);
nor U4862 (N_4862,N_492,N_2321);
nor U4863 (N_4863,N_1770,N_1439);
nand U4864 (N_4864,N_509,N_1792);
or U4865 (N_4865,N_1635,N_1282);
and U4866 (N_4866,N_1496,N_262);
nor U4867 (N_4867,N_1162,N_1351);
nand U4868 (N_4868,N_1390,N_2014);
nand U4869 (N_4869,N_797,N_1704);
nand U4870 (N_4870,N_2001,N_1489);
nand U4871 (N_4871,N_666,N_1342);
nand U4872 (N_4872,N_1748,N_746);
nor U4873 (N_4873,N_320,N_2152);
and U4874 (N_4874,N_1767,N_1788);
and U4875 (N_4875,N_1855,N_1314);
and U4876 (N_4876,N_1385,N_453);
or U4877 (N_4877,N_342,N_2428);
xnor U4878 (N_4878,N_2042,N_1024);
and U4879 (N_4879,N_258,N_0);
and U4880 (N_4880,N_42,N_1266);
and U4881 (N_4881,N_1892,N_2263);
or U4882 (N_4882,N_867,N_154);
and U4883 (N_4883,N_1370,N_2258);
and U4884 (N_4884,N_1541,N_1179);
and U4885 (N_4885,N_1276,N_886);
and U4886 (N_4886,N_867,N_1758);
and U4887 (N_4887,N_2149,N_1932);
nand U4888 (N_4888,N_194,N_2272);
nor U4889 (N_4889,N_1047,N_1314);
and U4890 (N_4890,N_781,N_809);
xor U4891 (N_4891,N_552,N_29);
or U4892 (N_4892,N_1539,N_1202);
or U4893 (N_4893,N_883,N_350);
and U4894 (N_4894,N_1541,N_816);
nor U4895 (N_4895,N_1618,N_947);
or U4896 (N_4896,N_2214,N_963);
and U4897 (N_4897,N_442,N_1228);
nand U4898 (N_4898,N_2251,N_775);
nor U4899 (N_4899,N_1337,N_705);
or U4900 (N_4900,N_810,N_1048);
xnor U4901 (N_4901,N_2129,N_1982);
and U4902 (N_4902,N_1838,N_1987);
nor U4903 (N_4903,N_462,N_908);
xor U4904 (N_4904,N_439,N_1402);
or U4905 (N_4905,N_340,N_1587);
nor U4906 (N_4906,N_1089,N_182);
and U4907 (N_4907,N_1239,N_1009);
nor U4908 (N_4908,N_130,N_1424);
and U4909 (N_4909,N_2304,N_2287);
nor U4910 (N_4910,N_2149,N_782);
nor U4911 (N_4911,N_1538,N_123);
and U4912 (N_4912,N_964,N_2289);
nor U4913 (N_4913,N_502,N_1218);
and U4914 (N_4914,N_28,N_2269);
nand U4915 (N_4915,N_942,N_2006);
nand U4916 (N_4916,N_1669,N_2210);
and U4917 (N_4917,N_2074,N_1905);
nand U4918 (N_4918,N_943,N_1025);
nand U4919 (N_4919,N_1126,N_2020);
nand U4920 (N_4920,N_2038,N_1810);
nor U4921 (N_4921,N_2000,N_408);
and U4922 (N_4922,N_1896,N_277);
nor U4923 (N_4923,N_1771,N_845);
and U4924 (N_4924,N_2398,N_2365);
or U4925 (N_4925,N_1334,N_915);
nor U4926 (N_4926,N_811,N_25);
and U4927 (N_4927,N_1573,N_2306);
nand U4928 (N_4928,N_1594,N_1437);
nand U4929 (N_4929,N_2010,N_1068);
or U4930 (N_4930,N_416,N_464);
nor U4931 (N_4931,N_2001,N_985);
nand U4932 (N_4932,N_2481,N_846);
and U4933 (N_4933,N_295,N_1273);
nor U4934 (N_4934,N_1962,N_181);
nand U4935 (N_4935,N_1349,N_338);
or U4936 (N_4936,N_178,N_584);
and U4937 (N_4937,N_1974,N_1207);
or U4938 (N_4938,N_1004,N_64);
nand U4939 (N_4939,N_350,N_1400);
nand U4940 (N_4940,N_969,N_2314);
nor U4941 (N_4941,N_642,N_191);
nor U4942 (N_4942,N_2276,N_146);
nor U4943 (N_4943,N_359,N_345);
nand U4944 (N_4944,N_642,N_2225);
nand U4945 (N_4945,N_1991,N_229);
and U4946 (N_4946,N_1282,N_2127);
or U4947 (N_4947,N_1425,N_1572);
or U4948 (N_4948,N_1685,N_807);
and U4949 (N_4949,N_2009,N_413);
nor U4950 (N_4950,N_1342,N_399);
or U4951 (N_4951,N_2189,N_419);
and U4952 (N_4952,N_1520,N_905);
or U4953 (N_4953,N_20,N_2164);
nor U4954 (N_4954,N_2264,N_420);
or U4955 (N_4955,N_2376,N_750);
nor U4956 (N_4956,N_920,N_1006);
or U4957 (N_4957,N_222,N_1427);
and U4958 (N_4958,N_156,N_940);
and U4959 (N_4959,N_232,N_675);
or U4960 (N_4960,N_2176,N_550);
or U4961 (N_4961,N_923,N_1372);
nor U4962 (N_4962,N_907,N_1776);
and U4963 (N_4963,N_1870,N_760);
and U4964 (N_4964,N_1939,N_1604);
and U4965 (N_4965,N_2113,N_1457);
and U4966 (N_4966,N_654,N_1243);
nand U4967 (N_4967,N_920,N_1382);
and U4968 (N_4968,N_2182,N_2177);
nor U4969 (N_4969,N_1216,N_1864);
xnor U4970 (N_4970,N_252,N_2232);
or U4971 (N_4971,N_2387,N_325);
xnor U4972 (N_4972,N_2278,N_2120);
or U4973 (N_4973,N_118,N_405);
or U4974 (N_4974,N_791,N_1181);
or U4975 (N_4975,N_1009,N_2347);
nand U4976 (N_4976,N_1419,N_2471);
nor U4977 (N_4977,N_1914,N_940);
nor U4978 (N_4978,N_2139,N_1064);
or U4979 (N_4979,N_1551,N_1980);
nor U4980 (N_4980,N_848,N_1128);
and U4981 (N_4981,N_1914,N_2169);
or U4982 (N_4982,N_2451,N_2062);
xor U4983 (N_4983,N_2255,N_1991);
or U4984 (N_4984,N_4,N_1434);
or U4985 (N_4985,N_1301,N_37);
and U4986 (N_4986,N_798,N_1067);
nor U4987 (N_4987,N_1943,N_1162);
nor U4988 (N_4988,N_1162,N_164);
xor U4989 (N_4989,N_64,N_1698);
or U4990 (N_4990,N_2012,N_1947);
nor U4991 (N_4991,N_1347,N_2462);
xor U4992 (N_4992,N_1882,N_704);
nand U4993 (N_4993,N_2220,N_1475);
and U4994 (N_4994,N_827,N_1100);
nand U4995 (N_4995,N_2218,N_1058);
nor U4996 (N_4996,N_760,N_1896);
nor U4997 (N_4997,N_472,N_2461);
nor U4998 (N_4998,N_1210,N_2057);
nand U4999 (N_4999,N_529,N_1960);
or U5000 (N_5000,N_3385,N_3606);
nand U5001 (N_5001,N_3642,N_4214);
or U5002 (N_5002,N_3375,N_2926);
or U5003 (N_5003,N_3810,N_2549);
nor U5004 (N_5004,N_3872,N_2629);
nand U5005 (N_5005,N_3163,N_3292);
or U5006 (N_5006,N_4216,N_2608);
or U5007 (N_5007,N_4783,N_3782);
nor U5008 (N_5008,N_3035,N_4217);
nor U5009 (N_5009,N_2686,N_4606);
and U5010 (N_5010,N_4863,N_3156);
or U5011 (N_5011,N_3837,N_4736);
or U5012 (N_5012,N_2957,N_3641);
nor U5013 (N_5013,N_3229,N_4945);
nand U5014 (N_5014,N_2746,N_2538);
and U5015 (N_5015,N_3317,N_3135);
nor U5016 (N_5016,N_4170,N_4349);
and U5017 (N_5017,N_4177,N_2670);
xor U5018 (N_5018,N_3728,N_3057);
nand U5019 (N_5019,N_3732,N_3380);
and U5020 (N_5020,N_4907,N_3090);
nand U5021 (N_5021,N_4448,N_3526);
and U5022 (N_5022,N_3643,N_3315);
nor U5023 (N_5023,N_4062,N_4430);
nand U5024 (N_5024,N_4145,N_4888);
nand U5025 (N_5025,N_3879,N_3992);
nand U5026 (N_5026,N_4687,N_3011);
nor U5027 (N_5027,N_4047,N_3362);
and U5028 (N_5028,N_3816,N_4238);
and U5029 (N_5029,N_3536,N_3186);
or U5030 (N_5030,N_4360,N_3275);
nand U5031 (N_5031,N_3657,N_4971);
nor U5032 (N_5032,N_3333,N_2831);
nor U5033 (N_5033,N_4308,N_4837);
and U5034 (N_5034,N_4056,N_4543);
or U5035 (N_5035,N_2758,N_4610);
nand U5036 (N_5036,N_3040,N_3861);
and U5037 (N_5037,N_2572,N_2666);
or U5038 (N_5038,N_2952,N_4143);
and U5039 (N_5039,N_2569,N_2505);
or U5040 (N_5040,N_4402,N_3258);
and U5041 (N_5041,N_3755,N_4532);
and U5042 (N_5042,N_2515,N_3123);
or U5043 (N_5043,N_3870,N_4635);
nand U5044 (N_5044,N_3891,N_4223);
or U5045 (N_5045,N_4972,N_3271);
nor U5046 (N_5046,N_2921,N_4642);
or U5047 (N_5047,N_4188,N_3354);
and U5048 (N_5048,N_4439,N_3935);
or U5049 (N_5049,N_3668,N_4626);
nand U5050 (N_5050,N_3136,N_3149);
and U5051 (N_5051,N_4748,N_3559);
and U5052 (N_5052,N_3045,N_4459);
nor U5053 (N_5053,N_4637,N_3640);
or U5054 (N_5054,N_2547,N_4664);
xor U5055 (N_5055,N_3570,N_2790);
nor U5056 (N_5056,N_4706,N_2979);
nand U5057 (N_5057,N_3002,N_4695);
nor U5058 (N_5058,N_4284,N_3304);
xnor U5059 (N_5059,N_3554,N_3975);
xnor U5060 (N_5060,N_3478,N_2688);
nand U5061 (N_5061,N_4785,N_4374);
xnor U5062 (N_5062,N_4844,N_4862);
or U5063 (N_5063,N_4488,N_2615);
nand U5064 (N_5064,N_4113,N_4613);
or U5065 (N_5065,N_3051,N_4717);
and U5066 (N_5066,N_3639,N_3082);
and U5067 (N_5067,N_4507,N_2668);
nand U5068 (N_5068,N_4832,N_3028);
and U5069 (N_5069,N_3916,N_2700);
nor U5070 (N_5070,N_2847,N_3137);
and U5071 (N_5071,N_4629,N_4497);
and U5072 (N_5072,N_2747,N_3415);
or U5073 (N_5073,N_4319,N_4701);
nand U5074 (N_5074,N_3153,N_4782);
or U5075 (N_5075,N_4949,N_3340);
or U5076 (N_5076,N_4006,N_3994);
or U5077 (N_5077,N_3813,N_2981);
or U5078 (N_5078,N_4141,N_3144);
or U5079 (N_5079,N_4833,N_4994);
or U5080 (N_5080,N_4363,N_4568);
nand U5081 (N_5081,N_4347,N_3902);
and U5082 (N_5082,N_2685,N_4152);
and U5083 (N_5083,N_4154,N_4764);
nor U5084 (N_5084,N_3052,N_4481);
or U5085 (N_5085,N_2945,N_3998);
nor U5086 (N_5086,N_4373,N_3131);
nor U5087 (N_5087,N_3704,N_4108);
and U5088 (N_5088,N_4622,N_3190);
or U5089 (N_5089,N_2646,N_2743);
nor U5090 (N_5090,N_3330,N_3392);
nor U5091 (N_5091,N_2617,N_4632);
nor U5092 (N_5092,N_3750,N_4253);
nor U5093 (N_5093,N_4416,N_3503);
nand U5094 (N_5094,N_3681,N_3308);
and U5095 (N_5095,N_2680,N_2794);
or U5096 (N_5096,N_3164,N_2533);
nor U5097 (N_5097,N_4352,N_2837);
nor U5098 (N_5098,N_4132,N_3637);
or U5099 (N_5099,N_4825,N_2920);
and U5100 (N_5100,N_4100,N_4151);
and U5101 (N_5101,N_3949,N_3276);
nor U5102 (N_5102,N_4175,N_3847);
and U5103 (N_5103,N_2932,N_4137);
nand U5104 (N_5104,N_4322,N_3351);
or U5105 (N_5105,N_3405,N_4546);
and U5106 (N_5106,N_3029,N_4400);
nor U5107 (N_5107,N_4130,N_2958);
or U5108 (N_5108,N_3513,N_3714);
nor U5109 (N_5109,N_3421,N_3845);
nor U5110 (N_5110,N_3284,N_2712);
nor U5111 (N_5111,N_4963,N_3169);
nor U5112 (N_5112,N_4368,N_3587);
and U5113 (N_5113,N_3698,N_4544);
and U5114 (N_5114,N_3202,N_3635);
nand U5115 (N_5115,N_3147,N_4298);
or U5116 (N_5116,N_4902,N_2554);
nand U5117 (N_5117,N_3341,N_2673);
nor U5118 (N_5118,N_4735,N_4570);
nand U5119 (N_5119,N_3107,N_4127);
or U5120 (N_5120,N_4234,N_4650);
xnor U5121 (N_5121,N_2718,N_3316);
nor U5122 (N_5122,N_4958,N_4725);
or U5123 (N_5123,N_2883,N_3841);
and U5124 (N_5124,N_2571,N_2527);
nand U5125 (N_5125,N_2600,N_3099);
and U5126 (N_5126,N_2587,N_4818);
or U5127 (N_5127,N_3967,N_4112);
nand U5128 (N_5128,N_4796,N_3623);
or U5129 (N_5129,N_2756,N_2730);
or U5130 (N_5130,N_4116,N_4657);
xnor U5131 (N_5131,N_3571,N_3314);
nor U5132 (N_5132,N_3900,N_3962);
and U5133 (N_5133,N_4817,N_4104);
nor U5134 (N_5134,N_3464,N_3961);
and U5135 (N_5135,N_4337,N_4277);
nand U5136 (N_5136,N_4072,N_4729);
nand U5137 (N_5137,N_4265,N_3644);
nor U5138 (N_5138,N_3208,N_2777);
or U5139 (N_5139,N_4752,N_4128);
nand U5140 (N_5140,N_3287,N_4342);
nor U5141 (N_5141,N_4569,N_4315);
nor U5142 (N_5142,N_4290,N_4683);
and U5143 (N_5143,N_3226,N_4566);
or U5144 (N_5144,N_3826,N_4375);
or U5145 (N_5145,N_4335,N_4280);
nor U5146 (N_5146,N_3209,N_4351);
or U5147 (N_5147,N_3656,N_3022);
nor U5148 (N_5148,N_2787,N_3778);
and U5149 (N_5149,N_2930,N_3007);
and U5150 (N_5150,N_4479,N_4634);
nand U5151 (N_5151,N_4719,N_3966);
or U5152 (N_5152,N_3734,N_4680);
nand U5153 (N_5153,N_3302,N_2934);
nor U5154 (N_5154,N_3990,N_4032);
and U5155 (N_5155,N_4089,N_2725);
nor U5156 (N_5156,N_3146,N_4530);
nor U5157 (N_5157,N_3827,N_3427);
or U5158 (N_5158,N_4625,N_3924);
nand U5159 (N_5159,N_2509,N_3168);
nand U5160 (N_5160,N_4466,N_3461);
nand U5161 (N_5161,N_3636,N_4462);
and U5162 (N_5162,N_3471,N_3013);
nand U5163 (N_5163,N_2836,N_2536);
or U5164 (N_5164,N_2601,N_4394);
nand U5165 (N_5165,N_2633,N_4336);
or U5166 (N_5166,N_3372,N_4604);
nand U5167 (N_5167,N_4079,N_4565);
and U5168 (N_5168,N_3970,N_4774);
and U5169 (N_5169,N_4326,N_3983);
and U5170 (N_5170,N_3999,N_3551);
nor U5171 (N_5171,N_4082,N_4457);
or U5172 (N_5172,N_3412,N_3181);
nor U5173 (N_5173,N_3555,N_2563);
nand U5174 (N_5174,N_3905,N_4976);
and U5175 (N_5175,N_4547,N_4918);
and U5176 (N_5176,N_2899,N_4854);
nor U5177 (N_5177,N_2690,N_2654);
or U5178 (N_5178,N_2842,N_2828);
and U5179 (N_5179,N_2558,N_2908);
nand U5180 (N_5180,N_4283,N_4895);
nor U5181 (N_5181,N_3723,N_3538);
nand U5182 (N_5182,N_2868,N_3758);
and U5183 (N_5183,N_3746,N_2887);
nor U5184 (N_5184,N_3824,N_4251);
or U5185 (N_5185,N_3987,N_4898);
nor U5186 (N_5186,N_4829,N_4811);
nand U5187 (N_5187,N_2895,N_2839);
nand U5188 (N_5188,N_2624,N_4867);
or U5189 (N_5189,N_3094,N_4668);
or U5190 (N_5190,N_4919,N_3669);
nand U5191 (N_5191,N_3675,N_3420);
and U5192 (N_5192,N_4377,N_3516);
nor U5193 (N_5193,N_3222,N_3610);
and U5194 (N_5194,N_4126,N_3880);
nand U5195 (N_5195,N_2812,N_3865);
nor U5196 (N_5196,N_3436,N_4185);
and U5197 (N_5197,N_3194,N_3466);
and U5198 (N_5198,N_3871,N_3006);
and U5199 (N_5199,N_2915,N_4696);
nor U5200 (N_5200,N_3005,N_4069);
or U5201 (N_5201,N_2693,N_4519);
nor U5202 (N_5202,N_4172,N_3470);
nand U5203 (N_5203,N_3066,N_3134);
xnor U5204 (N_5204,N_3701,N_3577);
nand U5205 (N_5205,N_3139,N_4969);
and U5206 (N_5206,N_4327,N_3702);
nor U5207 (N_5207,N_3976,N_2635);
nand U5208 (N_5208,N_3449,N_4313);
nand U5209 (N_5209,N_3991,N_2692);
and U5210 (N_5210,N_3798,N_3350);
or U5211 (N_5211,N_2864,N_3625);
nand U5212 (N_5212,N_2622,N_3337);
nor U5213 (N_5213,N_4615,N_4376);
and U5214 (N_5214,N_2590,N_3580);
nor U5215 (N_5215,N_4076,N_4094);
and U5216 (N_5216,N_3697,N_2826);
or U5217 (N_5217,N_3207,N_4876);
nor U5218 (N_5218,N_2516,N_4926);
nand U5219 (N_5219,N_2927,N_3482);
and U5220 (N_5220,N_4449,N_4429);
and U5221 (N_5221,N_4762,N_4150);
nor U5222 (N_5222,N_3024,N_3326);
nand U5223 (N_5223,N_3390,N_3525);
nand U5224 (N_5224,N_2785,N_3901);
or U5225 (N_5225,N_4574,N_2924);
nor U5226 (N_5226,N_2944,N_4821);
and U5227 (N_5227,N_4011,N_2805);
nand U5228 (N_5228,N_3632,N_3799);
nor U5229 (N_5229,N_3522,N_4297);
nor U5230 (N_5230,N_4523,N_2827);
nor U5231 (N_5231,N_2851,N_4779);
nand U5232 (N_5232,N_2704,N_4886);
and U5233 (N_5233,N_3821,N_4043);
nand U5234 (N_5234,N_2922,N_3026);
nand U5235 (N_5235,N_4968,N_3150);
and U5236 (N_5236,N_4845,N_3398);
and U5237 (N_5237,N_2745,N_3012);
nand U5238 (N_5238,N_2644,N_4630);
nand U5239 (N_5239,N_3709,N_4339);
and U5240 (N_5240,N_4765,N_3058);
and U5241 (N_5241,N_4077,N_2998);
nor U5242 (N_5242,N_2925,N_4598);
or U5243 (N_5243,N_4178,N_2573);
nand U5244 (N_5244,N_3004,N_3454);
nand U5245 (N_5245,N_4745,N_3437);
nand U5246 (N_5246,N_2948,N_4667);
nor U5247 (N_5247,N_3106,N_3439);
and U5248 (N_5248,N_3882,N_4215);
nor U5249 (N_5249,N_4623,N_4751);
and U5250 (N_5250,N_3739,N_4401);
and U5251 (N_5251,N_4105,N_3878);
or U5252 (N_5252,N_4200,N_3592);
nor U5253 (N_5253,N_4866,N_2714);
nor U5254 (N_5254,N_3620,N_3576);
nand U5255 (N_5255,N_3059,N_2970);
or U5256 (N_5256,N_4279,N_3568);
nand U5257 (N_5257,N_3433,N_2872);
or U5258 (N_5258,N_3469,N_4219);
and U5259 (N_5259,N_3025,N_3187);
nand U5260 (N_5260,N_4161,N_3815);
nand U5261 (N_5261,N_3027,N_4766);
nand U5262 (N_5262,N_4987,N_2506);
nand U5263 (N_5263,N_2556,N_3786);
or U5264 (N_5264,N_3130,N_4658);
nand U5265 (N_5265,N_3129,N_4900);
nand U5266 (N_5266,N_3797,N_3745);
or U5267 (N_5267,N_2893,N_4853);
and U5268 (N_5268,N_3868,N_3018);
nand U5269 (N_5269,N_3829,N_2859);
and U5270 (N_5270,N_2542,N_2738);
and U5271 (N_5271,N_3173,N_4605);
nor U5272 (N_5272,N_4474,N_3706);
and U5273 (N_5273,N_2882,N_3230);
nand U5274 (N_5274,N_3291,N_2795);
and U5275 (N_5275,N_3023,N_3850);
nor U5276 (N_5276,N_2963,N_4808);
nor U5277 (N_5277,N_3196,N_2551);
or U5278 (N_5278,N_4482,N_4260);
nor U5279 (N_5279,N_4620,N_2763);
or U5280 (N_5280,N_2656,N_4757);
and U5281 (N_5281,N_4292,N_4688);
nand U5282 (N_5282,N_4916,N_4274);
nor U5283 (N_5283,N_2512,N_3176);
nand U5284 (N_5284,N_4978,N_4885);
nand U5285 (N_5285,N_3856,N_3456);
and U5286 (N_5286,N_2698,N_4831);
and U5287 (N_5287,N_2820,N_4645);
or U5288 (N_5288,N_3553,N_3157);
or U5289 (N_5289,N_4189,N_3825);
or U5290 (N_5290,N_2645,N_3959);
nor U5291 (N_5291,N_4858,N_4982);
or U5292 (N_5292,N_3740,N_2679);
or U5293 (N_5293,N_4588,N_3852);
nand U5294 (N_5294,N_4852,N_2636);
or U5295 (N_5295,N_3583,N_4381);
and U5296 (N_5296,N_2620,N_3397);
nand U5297 (N_5297,N_4691,N_3273);
and U5298 (N_5298,N_4048,N_4996);
and U5299 (N_5299,N_4017,N_3960);
nand U5300 (N_5300,N_3529,N_2562);
nor U5301 (N_5301,N_3549,N_3319);
and U5302 (N_5302,N_3851,N_3406);
nand U5303 (N_5303,N_4961,N_3184);
and U5304 (N_5304,N_2736,N_3659);
or U5305 (N_5305,N_3424,N_2584);
nand U5306 (N_5306,N_4358,N_4052);
or U5307 (N_5307,N_4515,N_2732);
and U5308 (N_5308,N_4021,N_3805);
xor U5309 (N_5309,N_4295,N_3492);
and U5310 (N_5310,N_3743,N_4797);
xor U5311 (N_5311,N_2655,N_3682);
and U5312 (N_5312,N_4596,N_4518);
or U5313 (N_5313,N_4301,N_3175);
and U5314 (N_5314,N_2540,N_4597);
and U5315 (N_5315,N_3696,N_2613);
nand U5316 (N_5316,N_3790,N_4504);
nor U5317 (N_5317,N_3459,N_3820);
nand U5318 (N_5318,N_4934,N_3050);
or U5319 (N_5319,N_3996,N_3507);
or U5320 (N_5320,N_4289,N_4097);
and U5321 (N_5321,N_2570,N_2876);
nor U5322 (N_5322,N_4018,N_2996);
nand U5323 (N_5323,N_3977,N_3263);
and U5324 (N_5324,N_3925,N_3543);
or U5325 (N_5325,N_3744,N_3044);
and U5326 (N_5326,N_4164,N_4550);
and U5327 (N_5327,N_3360,N_3498);
nand U5328 (N_5328,N_4204,N_3217);
or U5329 (N_5329,N_4266,N_2508);
nand U5330 (N_5330,N_3270,N_3691);
or U5331 (N_5331,N_3748,N_4428);
nor U5332 (N_5332,N_3122,N_3769);
and U5333 (N_5333,N_4511,N_2610);
or U5334 (N_5334,N_2776,N_4795);
nand U5335 (N_5335,N_2760,N_4192);
or U5336 (N_5336,N_3085,N_4503);
or U5337 (N_5337,N_2535,N_3590);
and U5338 (N_5338,N_4988,N_4372);
or U5339 (N_5339,N_4035,N_4698);
or U5340 (N_5340,N_3835,N_3000);
and U5341 (N_5341,N_3947,N_2696);
nor U5342 (N_5342,N_4311,N_4830);
nand U5343 (N_5343,N_3678,N_2802);
nor U5344 (N_5344,N_3355,N_3067);
and U5345 (N_5345,N_4475,N_4201);
and U5346 (N_5346,N_4387,N_3544);
or U5347 (N_5347,N_3465,N_3930);
nor U5348 (N_5348,N_3227,N_4676);
or U5349 (N_5349,N_3649,N_3567);
nand U5350 (N_5350,N_2875,N_3191);
nand U5351 (N_5351,N_3545,N_4710);
and U5352 (N_5352,N_2817,N_3602);
or U5353 (N_5353,N_4659,N_4564);
nand U5354 (N_5354,N_3228,N_3694);
nor U5355 (N_5355,N_2733,N_4526);
and U5356 (N_5356,N_4396,N_2650);
or U5357 (N_5357,N_2742,N_2751);
nand U5358 (N_5358,N_2721,N_3411);
nor U5359 (N_5359,N_3854,N_3952);
nand U5360 (N_5360,N_2514,N_3448);
and U5361 (N_5361,N_4158,N_3695);
or U5362 (N_5362,N_4554,N_3773);
nand U5363 (N_5363,N_4524,N_4771);
nand U5364 (N_5364,N_3760,N_2757);
nand U5365 (N_5365,N_4212,N_4925);
or U5366 (N_5366,N_4222,N_4302);
nor U5367 (N_5367,N_3328,N_4397);
or U5368 (N_5368,N_2834,N_4573);
and U5369 (N_5369,N_3908,N_3352);
or U5370 (N_5370,N_4784,N_4002);
nor U5371 (N_5371,N_2560,N_2748);
nor U5372 (N_5372,N_3838,N_4619);
nor U5373 (N_5373,N_3289,N_4914);
nor U5374 (N_5374,N_3846,N_2701);
or U5375 (N_5375,N_4495,N_4560);
nand U5376 (N_5376,N_3972,N_2781);
or U5377 (N_5377,N_3599,N_4258);
and U5378 (N_5378,N_3113,N_4835);
nor U5379 (N_5379,N_3237,N_3515);
or U5380 (N_5380,N_4226,N_3906);
or U5381 (N_5381,N_3020,N_4577);
and U5382 (N_5382,N_2792,N_3586);
or U5383 (N_5383,N_2699,N_4276);
nand U5384 (N_5384,N_2967,N_4191);
or U5385 (N_5385,N_2797,N_4741);
and U5386 (N_5386,N_4707,N_3096);
nor U5387 (N_5387,N_4148,N_3738);
nand U5388 (N_5388,N_3251,N_4425);
or U5389 (N_5389,N_4468,N_4979);
nor U5390 (N_5390,N_3761,N_3788);
or U5391 (N_5391,N_3775,N_4897);
nor U5392 (N_5392,N_4559,N_2914);
nand U5393 (N_5393,N_2898,N_4792);
nand U5394 (N_5394,N_4587,N_3776);
or U5395 (N_5395,N_4552,N_4271);
or U5396 (N_5396,N_4672,N_2607);
or U5397 (N_5397,N_4165,N_4927);
nand U5398 (N_5398,N_3777,N_4010);
nand U5399 (N_5399,N_3384,N_3517);
or U5400 (N_5400,N_2648,N_4241);
and U5401 (N_5401,N_2521,N_4293);
or U5402 (N_5402,N_4548,N_2722);
nor U5403 (N_5403,N_3303,N_4663);
and U5404 (N_5404,N_4412,N_3578);
nand U5405 (N_5405,N_3034,N_3512);
and U5406 (N_5406,N_2943,N_4628);
nand U5407 (N_5407,N_4029,N_3312);
nor U5408 (N_5408,N_3105,N_3366);
nand U5409 (N_5409,N_4964,N_4730);
and U5410 (N_5410,N_4436,N_4404);
or U5411 (N_5411,N_2773,N_2999);
xor U5412 (N_5412,N_4465,N_4044);
or U5413 (N_5413,N_3626,N_2539);
or U5414 (N_5414,N_3888,N_4937);
or U5415 (N_5415,N_3876,N_4364);
and U5416 (N_5416,N_4936,N_2510);
and U5417 (N_5417,N_2994,N_3299);
nand U5418 (N_5418,N_4344,N_4159);
or U5419 (N_5419,N_3386,N_3347);
or U5420 (N_5420,N_2578,N_4405);
nand U5421 (N_5421,N_2923,N_3918);
nor U5422 (N_5422,N_4814,N_2591);
nor U5423 (N_5423,N_4003,N_2749);
nand U5424 (N_5424,N_3814,N_3460);
nor U5425 (N_5425,N_4064,N_2741);
nor U5426 (N_5426,N_3313,N_3864);
nand U5427 (N_5427,N_4367,N_2965);
xor U5428 (N_5428,N_4753,N_3754);
nand U5429 (N_5429,N_3087,N_3542);
or U5430 (N_5430,N_3402,N_4001);
or U5431 (N_5431,N_2709,N_3686);
nor U5432 (N_5432,N_4561,N_2818);
and U5433 (N_5433,N_3383,N_3489);
nor U5434 (N_5434,N_4884,N_2577);
and U5435 (N_5435,N_3032,N_4860);
xor U5436 (N_5436,N_2564,N_3982);
and U5437 (N_5437,N_4286,N_2596);
nor U5438 (N_5438,N_3774,N_4539);
and U5439 (N_5439,N_3611,N_4102);
and U5440 (N_5440,N_3371,N_4330);
nand U5441 (N_5441,N_2843,N_2774);
or U5442 (N_5442,N_3408,N_4306);
and U5443 (N_5443,N_2676,N_2857);
and U5444 (N_5444,N_4486,N_2772);
nor U5445 (N_5445,N_3496,N_4157);
nor U5446 (N_5446,N_4173,N_4180);
nand U5447 (N_5447,N_4910,N_3546);
and U5448 (N_5448,N_3409,N_4960);
nor U5449 (N_5449,N_2822,N_2545);
nor U5450 (N_5450,N_4060,N_3484);
nor U5451 (N_5451,N_3565,N_3633);
and U5452 (N_5452,N_4849,N_3839);
nor U5453 (N_5453,N_3016,N_2737);
nand U5454 (N_5454,N_2936,N_4174);
or U5455 (N_5455,N_3365,N_4567);
nand U5456 (N_5456,N_3800,N_3345);
or U5457 (N_5457,N_3737,N_4492);
nand U5458 (N_5458,N_4231,N_4601);
and U5459 (N_5459,N_3429,N_2766);
or U5460 (N_5460,N_3892,N_3662);
and U5461 (N_5461,N_3680,N_4847);
or U5462 (N_5462,N_3631,N_3223);
nand U5463 (N_5463,N_4822,N_4438);
or U5464 (N_5464,N_3894,N_3225);
or U5465 (N_5465,N_3417,N_2580);
nor U5466 (N_5466,N_4183,N_2678);
and U5467 (N_5467,N_2630,N_4882);
nand U5468 (N_5468,N_2659,N_4304);
and U5469 (N_5469,N_2912,N_3540);
and U5470 (N_5470,N_2603,N_3765);
and U5471 (N_5471,N_2838,N_3628);
nand U5472 (N_5472,N_4197,N_4815);
and U5473 (N_5473,N_2684,N_3717);
nand U5474 (N_5474,N_3121,N_3250);
and U5475 (N_5475,N_4230,N_4646);
or U5476 (N_5476,N_3564,N_3652);
and U5477 (N_5477,N_4700,N_3497);
nand U5478 (N_5478,N_3843,N_2529);
nor U5479 (N_5479,N_2582,N_2829);
nand U5480 (N_5480,N_3603,N_2705);
nor U5481 (N_5481,N_3591,N_3807);
nor U5482 (N_5482,N_4681,N_3205);
or U5483 (N_5483,N_3376,N_4660);
or U5484 (N_5484,N_3183,N_4464);
xor U5485 (N_5485,N_4262,N_3811);
nand U5486 (N_5486,N_3699,N_3110);
and U5487 (N_5487,N_4022,N_2768);
and U5488 (N_5488,N_4321,N_4013);
and U5489 (N_5489,N_3098,N_4407);
nor U5490 (N_5490,N_4242,N_3895);
nor U5491 (N_5491,N_3883,N_4312);
nand U5492 (N_5492,N_2885,N_4708);
nor U5493 (N_5493,N_3294,N_2977);
nor U5494 (N_5494,N_4555,N_2697);
xor U5495 (N_5495,N_4788,N_4506);
or U5496 (N_5496,N_4618,N_4585);
and U5497 (N_5497,N_3689,N_3957);
xor U5498 (N_5498,N_3311,N_2968);
and U5499 (N_5499,N_3306,N_3056);
or U5500 (N_5500,N_2900,N_2810);
nand U5501 (N_5501,N_3458,N_4140);
nand U5502 (N_5502,N_4210,N_3574);
or U5503 (N_5503,N_4602,N_3092);
nand U5504 (N_5504,N_3180,N_3071);
and U5505 (N_5505,N_4122,N_4278);
and U5506 (N_5506,N_2513,N_4036);
nand U5507 (N_5507,N_3419,N_4582);
nor U5508 (N_5508,N_2652,N_4747);
and U5509 (N_5509,N_3446,N_3898);
and U5510 (N_5510,N_4168,N_4758);
or U5511 (N_5511,N_3653,N_2980);
nor U5512 (N_5512,N_4865,N_4611);
nand U5513 (N_5513,N_4702,N_3242);
or U5514 (N_5514,N_2976,N_3581);
nand U5515 (N_5515,N_3008,N_4699);
nand U5516 (N_5516,N_4643,N_3995);
and U5517 (N_5517,N_3595,N_3951);
nor U5518 (N_5518,N_2755,N_2565);
nand U5519 (N_5519,N_4133,N_3182);
and U5520 (N_5520,N_3455,N_2647);
nand U5521 (N_5521,N_4943,N_3053);
or U5522 (N_5522,N_3500,N_3479);
or U5523 (N_5523,N_2771,N_4955);
and U5524 (N_5524,N_4440,N_4494);
nor U5525 (N_5525,N_3929,N_3387);
or U5526 (N_5526,N_3795,N_3725);
and U5527 (N_5527,N_3037,N_3081);
nor U5528 (N_5528,N_3014,N_2989);
or U5529 (N_5529,N_3486,N_4786);
nand U5530 (N_5530,N_3001,N_3869);
or U5531 (N_5531,N_4087,N_3462);
and U5532 (N_5532,N_4254,N_3844);
xor U5533 (N_5533,N_4692,N_3757);
xor U5534 (N_5534,N_4843,N_4983);
or U5535 (N_5535,N_4644,N_4000);
nand U5536 (N_5536,N_3527,N_3309);
nand U5537 (N_5537,N_4746,N_4944);
or U5538 (N_5538,N_2585,N_3033);
or U5539 (N_5539,N_3965,N_4513);
and U5540 (N_5540,N_4435,N_3942);
nand U5541 (N_5541,N_2561,N_3812);
or U5542 (N_5542,N_3166,N_2939);
and U5543 (N_5543,N_3323,N_4186);
nor U5544 (N_5544,N_3600,N_4073);
or U5545 (N_5545,N_3700,N_3480);
or U5546 (N_5546,N_4163,N_3508);
nand U5547 (N_5547,N_4731,N_4928);
and U5548 (N_5548,N_3069,N_4913);
nand U5549 (N_5549,N_4827,N_4422);
nor U5550 (N_5550,N_2660,N_2519);
nand U5551 (N_5551,N_4096,N_3256);
and U5552 (N_5552,N_3391,N_4763);
nor U5553 (N_5553,N_3444,N_4962);
and U5554 (N_5554,N_4307,N_3434);
and U5555 (N_5555,N_3676,N_2507);
nor U5556 (N_5556,N_3719,N_2502);
nor U5557 (N_5557,N_3189,N_3556);
nor U5558 (N_5558,N_4129,N_2595);
and U5559 (N_5559,N_4328,N_3934);
nand U5560 (N_5560,N_3809,N_3818);
or U5561 (N_5561,N_3487,N_3715);
and U5562 (N_5562,N_4156,N_3231);
nand U5563 (N_5563,N_3793,N_4107);
xor U5564 (N_5564,N_4353,N_4472);
nor U5565 (N_5565,N_2675,N_4004);
or U5566 (N_5566,N_4841,N_3684);
nand U5567 (N_5567,N_4477,N_2956);
or U5568 (N_5568,N_3651,N_4023);
nand U5569 (N_5569,N_4420,N_3440);
and U5570 (N_5570,N_3585,N_3441);
nor U5571 (N_5571,N_3198,N_3519);
or U5572 (N_5572,N_3054,N_3243);
or U5573 (N_5573,N_2778,N_3070);
nor U5574 (N_5574,N_3938,N_4727);
or U5575 (N_5575,N_4235,N_2931);
and U5576 (N_5576,N_4749,N_4614);
or U5577 (N_5577,N_2767,N_2671);
nor U5578 (N_5578,N_4389,N_3922);
or U5579 (N_5579,N_2504,N_4732);
nand U5580 (N_5580,N_3203,N_3569);
xor U5581 (N_5581,N_3979,N_3502);
and U5582 (N_5582,N_2664,N_3296);
nand U5583 (N_5583,N_4496,N_4742);
nand U5584 (N_5584,N_3241,N_3060);
nor U5585 (N_5585,N_3624,N_3566);
or U5586 (N_5586,N_3727,N_4441);
nand U5587 (N_5587,N_3617,N_3781);
nor U5588 (N_5588,N_3216,N_4446);
nand U5589 (N_5589,N_4090,N_4921);
and U5590 (N_5590,N_4379,N_3572);
and U5591 (N_5591,N_3363,N_3667);
nor U5592 (N_5592,N_3802,N_4693);
nor U5593 (N_5593,N_4923,N_4538);
nand U5594 (N_5594,N_2602,N_3831);
or U5595 (N_5595,N_3505,N_3331);
nand U5596 (N_5596,N_4591,N_3335);
nand U5597 (N_5597,N_4607,N_4093);
and U5598 (N_5598,N_3562,N_3445);
xnor U5599 (N_5599,N_4670,N_3065);
or U5600 (N_5600,N_4531,N_2770);
nor U5601 (N_5601,N_4046,N_3148);
and U5602 (N_5602,N_4810,N_4716);
and U5603 (N_5603,N_4576,N_4859);
nor U5604 (N_5604,N_4008,N_3654);
nand U5605 (N_5605,N_3622,N_3932);
nand U5606 (N_5606,N_3240,N_3716);
nand U5607 (N_5607,N_3161,N_3224);
and U5608 (N_5608,N_3254,N_3504);
nor U5609 (N_5609,N_4252,N_4679);
and U5610 (N_5610,N_3579,N_2942);
or U5611 (N_5611,N_2726,N_2858);
or U5612 (N_5612,N_2752,N_4967);
nor U5613 (N_5613,N_3467,N_3560);
or U5614 (N_5614,N_2870,N_3055);
nor U5615 (N_5615,N_3213,N_2744);
nand U5616 (N_5616,N_4331,N_4873);
nand U5617 (N_5617,N_3946,N_3749);
nor U5618 (N_5618,N_3931,N_4684);
nand U5619 (N_5619,N_3655,N_3944);
or U5620 (N_5620,N_3860,N_4640);
and U5621 (N_5621,N_4456,N_3233);
nand U5622 (N_5622,N_2850,N_4805);
and U5623 (N_5623,N_4155,N_4065);
nor U5624 (N_5624,N_4267,N_3188);
and U5625 (N_5625,N_4469,N_4755);
and U5626 (N_5626,N_4303,N_2727);
nor U5627 (N_5627,N_4124,N_4789);
or U5628 (N_5628,N_3679,N_3780);
nand U5629 (N_5629,N_3819,N_4869);
nor U5630 (N_5630,N_2574,N_3115);
and U5631 (N_5631,N_2806,N_3613);
nor U5632 (N_5632,N_3890,N_3178);
and U5633 (N_5633,N_2543,N_3660);
and U5634 (N_5634,N_3393,N_4600);
xnor U5635 (N_5635,N_3248,N_2871);
nand U5636 (N_5636,N_4998,N_4224);
nor U5637 (N_5637,N_4648,N_4080);
or U5638 (N_5638,N_2691,N_4268);
nand U5639 (N_5639,N_3605,N_3152);
and U5640 (N_5640,N_4119,N_4933);
nor U5641 (N_5641,N_4638,N_2500);
nand U5642 (N_5642,N_3558,N_3266);
nor U5643 (N_5643,N_4190,N_4842);
or U5644 (N_5644,N_4391,N_2935);
nand U5645 (N_5645,N_3041,N_3561);
nor U5646 (N_5646,N_3255,N_4509);
nand U5647 (N_5647,N_4992,N_2642);
and U5648 (N_5648,N_3803,N_3080);
nor U5649 (N_5649,N_2824,N_3359);
or U5650 (N_5650,N_4361,N_4616);
nand U5651 (N_5651,N_3768,N_2555);
or U5652 (N_5652,N_2604,N_3741);
and U5653 (N_5653,N_2788,N_3320);
or U5654 (N_5654,N_4399,N_3245);
nor U5655 (N_5655,N_4540,N_3074);
or U5656 (N_5656,N_2626,N_2974);
or U5657 (N_5657,N_2634,N_4609);
nor U5658 (N_5658,N_3974,N_4879);
nor U5659 (N_5659,N_3801,N_4502);
and U5660 (N_5660,N_3141,N_4535);
and U5661 (N_5661,N_4649,N_4750);
nand U5662 (N_5662,N_3109,N_3683);
nand U5663 (N_5663,N_4366,N_3855);
and U5664 (N_5664,N_2581,N_3435);
and U5665 (N_5665,N_3563,N_4593);
or U5666 (N_5666,N_2910,N_3638);
and U5667 (N_5667,N_3510,N_3936);
or U5668 (N_5668,N_3783,N_2983);
or U5669 (N_5669,N_4179,N_3661);
nor U5670 (N_5670,N_4718,N_4499);
or U5671 (N_5671,N_3817,N_4990);
nor U5672 (N_5672,N_4453,N_2579);
nor U5673 (N_5673,N_3221,N_4426);
nand U5674 (N_5674,N_2984,N_4227);
nand U5675 (N_5675,N_3290,N_3370);
nand U5676 (N_5676,N_3630,N_3666);
nand U5677 (N_5677,N_4229,N_3971);
and U5678 (N_5678,N_3984,N_3418);
nor U5679 (N_5679,N_4024,N_4300);
nor U5680 (N_5680,N_3866,N_3729);
nand U5681 (N_5681,N_4054,N_3753);
nand U5682 (N_5682,N_4948,N_3926);
nand U5683 (N_5683,N_3937,N_4458);
and U5684 (N_5684,N_3432,N_2643);
and U5685 (N_5685,N_3172,N_3808);
or U5686 (N_5686,N_2884,N_4309);
nand U5687 (N_5687,N_3073,N_4678);
and U5688 (N_5688,N_4516,N_4355);
nand U5689 (N_5689,N_2694,N_3463);
and U5690 (N_5690,N_3127,N_3557);
nor U5691 (N_5691,N_4893,N_3249);
and U5692 (N_5692,N_4917,N_4798);
or U5693 (N_5693,N_4655,N_4121);
or U5694 (N_5694,N_4166,N_4483);
and U5695 (N_5695,N_2933,N_4848);
nor U5696 (N_5696,N_3038,N_2661);
nor U5697 (N_5697,N_2511,N_4633);
and U5698 (N_5698,N_4202,N_2779);
nand U5699 (N_5699,N_4434,N_2557);
or U5700 (N_5700,N_2841,N_2867);
or U5701 (N_5701,N_2960,N_2576);
nand U5702 (N_5702,N_3764,N_4739);
nor U5703 (N_5703,N_3722,N_2821);
and U5704 (N_5704,N_2729,N_4999);
or U5705 (N_5705,N_3511,N_2750);
nor U5706 (N_5706,N_4142,N_4802);
or U5707 (N_5707,N_3283,N_2892);
nand U5708 (N_5708,N_2840,N_3101);
nor U5709 (N_5709,N_4819,N_3945);
nand U5710 (N_5710,N_4878,N_2552);
or U5711 (N_5711,N_3167,N_4380);
nand U5712 (N_5712,N_3766,N_4641);
and U5713 (N_5713,N_2854,N_2716);
nand U5714 (N_5714,N_3903,N_3112);
and U5715 (N_5715,N_4333,N_4639);
nor U5716 (N_5716,N_4666,N_4533);
and U5717 (N_5717,N_2961,N_4704);
nor U5718 (N_5718,N_2677,N_3428);
or U5719 (N_5719,N_4196,N_2663);
nand U5720 (N_5720,N_3343,N_3236);
nand U5721 (N_5721,N_3621,N_4790);
and U5722 (N_5722,N_2780,N_3368);
xor U5723 (N_5723,N_4595,N_3200);
nor U5724 (N_5724,N_4444,N_3031);
and U5725 (N_5725,N_4395,N_4673);
nor U5726 (N_5726,N_2845,N_4030);
nand U5727 (N_5727,N_2501,N_4371);
nand U5728 (N_5728,N_3881,N_3215);
and U5729 (N_5729,N_4887,N_2860);
and U5730 (N_5730,N_2717,N_2583);
and U5731 (N_5731,N_3321,N_3452);
and U5732 (N_5732,N_3956,N_2753);
and U5733 (N_5733,N_4500,N_3003);
nor U5734 (N_5734,N_2969,N_2973);
nor U5735 (N_5735,N_3747,N_3634);
or U5736 (N_5736,N_3842,N_3307);
nand U5737 (N_5737,N_4807,N_3353);
nand U5738 (N_5738,N_3039,N_3278);
nor U5739 (N_5739,N_4287,N_4162);
or U5740 (N_5740,N_2651,N_3400);
nand U5741 (N_5741,N_4915,N_2653);
nand U5742 (N_5742,N_2711,N_3804);
or U5743 (N_5743,N_4206,N_3832);
or U5744 (N_5744,N_2940,N_3477);
nand U5745 (N_5745,N_2526,N_3874);
nor U5746 (N_5746,N_4904,N_2833);
and U5747 (N_5747,N_3162,N_2995);
nor U5748 (N_5748,N_3378,N_4721);
nor U5749 (N_5749,N_3756,N_4450);
nand U5750 (N_5750,N_3095,N_3524);
and U5751 (N_5751,N_2575,N_4099);
nand U5752 (N_5752,N_3886,N_4343);
or U5753 (N_5753,N_3410,N_4443);
or U5754 (N_5754,N_2775,N_3751);
or U5755 (N_5755,N_4669,N_4872);
or U5756 (N_5756,N_4111,N_3015);
nand U5757 (N_5757,N_4671,N_4317);
nand U5758 (N_5758,N_3614,N_3896);
nor U5759 (N_5759,N_3648,N_4775);
and U5760 (N_5760,N_2594,N_4726);
nand U5761 (N_5761,N_4318,N_4016);
nand U5762 (N_5762,N_4256,N_4557);
xnor U5763 (N_5763,N_3382,N_3533);
and U5764 (N_5764,N_4370,N_3796);
nand U5765 (N_5765,N_3859,N_2901);
or U5766 (N_5766,N_4282,N_3849);
or U5767 (N_5767,N_4045,N_3887);
xnor U5768 (N_5768,N_3091,N_2951);
or U5769 (N_5769,N_2782,N_4864);
nor U5770 (N_5770,N_4038,N_3049);
and U5771 (N_5771,N_4993,N_3920);
or U5772 (N_5772,N_3142,N_4768);
nor U5773 (N_5773,N_3784,N_4690);
or U5774 (N_5774,N_4661,N_4039);
nand U5775 (N_5775,N_4259,N_4744);
nor U5776 (N_5776,N_2906,N_4432);
nand U5777 (N_5777,N_4037,N_2681);
nor U5778 (N_5778,N_4244,N_2846);
nor U5779 (N_5779,N_4930,N_3584);
nand U5780 (N_5780,N_3019,N_4883);
or U5781 (N_5781,N_4946,N_2865);
and U5782 (N_5782,N_2523,N_3265);
nand U5783 (N_5783,N_3076,N_2605);
or U5784 (N_5784,N_4711,N_3963);
and U5785 (N_5785,N_3730,N_2762);
and U5786 (N_5786,N_3118,N_3195);
nor U5787 (N_5787,N_3939,N_3483);
and U5788 (N_5788,N_2953,N_4118);
nor U5789 (N_5789,N_4627,N_2713);
nand U5790 (N_5790,N_3438,N_4553);
or U5791 (N_5791,N_4437,N_4409);
and U5792 (N_5792,N_4207,N_2658);
or U5793 (N_5793,N_3604,N_4652);
or U5794 (N_5794,N_4269,N_4147);
or U5795 (N_5795,N_3928,N_3179);
nor U5796 (N_5796,N_2702,N_3550);
and U5797 (N_5797,N_4586,N_3528);
and U5798 (N_5798,N_3119,N_2723);
nand U5799 (N_5799,N_4737,N_4951);
or U5800 (N_5800,N_3252,N_4106);
xnor U5801 (N_5801,N_4176,N_4071);
and U5802 (N_5802,N_4985,N_3670);
or U5803 (N_5803,N_2611,N_4041);
and U5804 (N_5804,N_4050,N_3547);
or U5805 (N_5805,N_3833,N_4986);
nand U5806 (N_5806,N_3862,N_2966);
nor U5807 (N_5807,N_3955,N_3618);
nand U5808 (N_5808,N_4491,N_4724);
nor U5809 (N_5809,N_3541,N_4485);
and U5810 (N_5810,N_2784,N_2532);
or U5811 (N_5811,N_3357,N_2878);
and U5812 (N_5812,N_4575,N_4583);
and U5813 (N_5813,N_2835,N_3358);
nor U5814 (N_5814,N_4261,N_4187);
nor U5815 (N_5815,N_4305,N_4417);
or U5816 (N_5816,N_4193,N_3128);
and U5817 (N_5817,N_4498,N_4793);
or U5818 (N_5818,N_4647,N_4599);
or U5819 (N_5819,N_4362,N_4086);
and U5820 (N_5820,N_3720,N_2568);
and U5821 (N_5821,N_4460,N_3759);
nand U5822 (N_5822,N_3204,N_4320);
nand U5823 (N_5823,N_2609,N_2559);
nor U5824 (N_5824,N_4257,N_4490);
or U5825 (N_5825,N_4542,N_4922);
nor U5826 (N_5826,N_3672,N_3506);
or U5827 (N_5827,N_4406,N_3885);
nor U5828 (N_5828,N_3272,N_4419);
or U5829 (N_5829,N_4249,N_4480);
nor U5830 (N_5830,N_3084,N_2890);
and U5831 (N_5831,N_3373,N_3009);
nor U5832 (N_5832,N_4068,N_2990);
nand U5833 (N_5833,N_2550,N_2525);
and U5834 (N_5834,N_3475,N_3980);
nand U5835 (N_5835,N_3485,N_4115);
nand U5836 (N_5836,N_4232,N_2528);
nor U5837 (N_5837,N_4199,N_2641);
nand U5838 (N_5838,N_3601,N_3451);
nand U5839 (N_5839,N_4467,N_2544);
nor U5840 (N_5840,N_3509,N_4421);
nand U5841 (N_5841,N_4579,N_4901);
nor U5842 (N_5842,N_3160,N_3899);
and U5843 (N_5843,N_4813,N_4194);
and U5844 (N_5844,N_3915,N_4463);
nor U5845 (N_5845,N_3532,N_2852);
and U5846 (N_5846,N_2855,N_3369);
or U5847 (N_5847,N_2631,N_3736);
or U5848 (N_5848,N_3165,N_3779);
nand U5849 (N_5849,N_4912,N_3615);
nor U5850 (N_5850,N_2789,N_4941);
nand U5851 (N_5851,N_4388,N_3117);
and U5852 (N_5852,N_3154,N_3379);
and U5853 (N_5853,N_2597,N_4034);
and U5854 (N_5854,N_3629,N_4451);
and U5855 (N_5855,N_4015,N_3132);
or U5856 (N_5856,N_3713,N_3884);
nor U5857 (N_5857,N_2861,N_3261);
nand U5858 (N_5858,N_3262,N_4773);
or U5859 (N_5859,N_3552,N_4057);
nor U5860 (N_5860,N_4255,N_4505);
and U5861 (N_5861,N_4682,N_4685);
or U5862 (N_5862,N_3907,N_2988);
nand U5863 (N_5863,N_4911,N_4135);
nor U5864 (N_5864,N_3170,N_4493);
nor U5865 (N_5865,N_2804,N_4952);
and U5866 (N_5866,N_2674,N_2759);
and U5867 (N_5867,N_3921,N_2830);
or U5868 (N_5868,N_4521,N_3244);
or U5869 (N_5869,N_4131,N_4074);
and U5870 (N_5870,N_3277,N_3711);
nand U5871 (N_5871,N_4019,N_4957);
nand U5872 (N_5872,N_3822,N_4489);
or U5873 (N_5873,N_2886,N_2589);
or U5874 (N_5874,N_3548,N_3985);
and U5875 (N_5875,N_3234,N_3318);
nand U5876 (N_5876,N_3177,N_3158);
and U5877 (N_5877,N_4675,N_2913);
and U5878 (N_5878,N_4812,N_3494);
or U5879 (N_5879,N_4720,N_2992);
nand U5880 (N_5880,N_4563,N_2807);
or U5881 (N_5881,N_3520,N_3210);
nand U5882 (N_5882,N_4723,N_3414);
and U5883 (N_5883,N_3377,N_4760);
or U5884 (N_5884,N_2672,N_3401);
and U5885 (N_5885,N_4846,N_4942);
nor U5886 (N_5886,N_4534,N_3036);
and U5887 (N_5887,N_4769,N_4929);
and U5888 (N_5888,N_4572,N_3269);
nand U5889 (N_5889,N_3958,N_2720);
nand U5890 (N_5890,N_3645,N_3997);
nor U5891 (N_5891,N_4947,N_4350);
nor U5892 (N_5892,N_4804,N_2928);
nor U5893 (N_5893,N_4078,N_3274);
and U5894 (N_5894,N_3218,N_4677);
or U5895 (N_5895,N_4954,N_2710);
nand U5896 (N_5896,N_4213,N_3889);
and U5897 (N_5897,N_2687,N_3650);
xnor U5898 (N_5898,N_3338,N_3863);
and U5899 (N_5899,N_4908,N_3647);
and U5900 (N_5900,N_4386,N_3214);
or U5901 (N_5901,N_4323,N_3597);
nand U5902 (N_5902,N_3940,N_3493);
and U5903 (N_5903,N_4525,N_3612);
or U5904 (N_5904,N_4508,N_4794);
or U5905 (N_5905,N_2849,N_3282);
nand U5906 (N_5906,N_3677,N_3442);
nand U5907 (N_5907,N_4665,N_3361);
or U5908 (N_5908,N_4031,N_3285);
nor U5909 (N_5909,N_2588,N_3246);
nor U5910 (N_5910,N_2503,N_2881);
or U5911 (N_5911,N_4608,N_4991);
nor U5912 (N_5912,N_3616,N_4780);
or U5913 (N_5913,N_3791,N_3501);
nor U5914 (N_5914,N_4995,N_4651);
nor U5915 (N_5915,N_3344,N_3422);
or U5916 (N_5916,N_2546,N_3785);
nand U5917 (N_5917,N_4236,N_3708);
and U5918 (N_5918,N_3364,N_4903);
or U5919 (N_5919,N_4316,N_4636);
nor U5920 (N_5920,N_2955,N_3324);
nor U5921 (N_5921,N_2632,N_3718);
or U5922 (N_5922,N_3171,N_4110);
and U5923 (N_5923,N_3912,N_4899);
nor U5924 (N_5924,N_3619,N_3910);
xnor U5925 (N_5925,N_4061,N_2592);
nand U5926 (N_5926,N_4722,N_4123);
and U5927 (N_5927,N_2662,N_3575);
nor U5928 (N_5928,N_3447,N_3943);
nand U5929 (N_5929,N_3431,N_4767);
or U5930 (N_5930,N_3986,N_3381);
nand U5931 (N_5931,N_4875,N_3426);
nor U5932 (N_5932,N_3295,N_3665);
nand U5933 (N_5933,N_3257,N_4025);
nor U5934 (N_5934,N_3933,N_4334);
or U5935 (N_5935,N_2903,N_2880);
nor U5936 (N_5936,N_4346,N_4528);
and U5937 (N_5937,N_2905,N_4756);
nand U5938 (N_5938,N_3787,N_3140);
and U5939 (N_5939,N_3927,N_2902);
nand U5940 (N_5940,N_3443,N_4058);
nand U5941 (N_5941,N_3794,N_3735);
or U5942 (N_5942,N_3367,N_4411);
nand U5943 (N_5943,N_3627,N_4776);
nor U5944 (N_5944,N_4447,N_2618);
or U5945 (N_5945,N_4855,N_3473);
nor U5946 (N_5946,N_2593,N_4012);
xnor U5947 (N_5947,N_3293,N_2832);
and U5948 (N_5948,N_4932,N_2619);
and U5949 (N_5949,N_3062,N_4703);
nand U5950 (N_5950,N_3989,N_4085);
and U5951 (N_5951,N_3093,N_3151);
and U5952 (N_5952,N_4026,N_4423);
or U5953 (N_5953,N_4454,N_4512);
or U5954 (N_5954,N_2649,N_2918);
or U5955 (N_5955,N_4338,N_3457);
nor U5956 (N_5956,N_3267,N_4171);
nand U5957 (N_5957,N_4167,N_2897);
and U5958 (N_5958,N_3968,N_3403);
nand U5959 (N_5959,N_3663,N_4989);
or U5960 (N_5960,N_4868,N_3911);
nand U5961 (N_5961,N_3124,N_3671);
nand U5962 (N_5962,N_2894,N_3836);
nand U5963 (N_5963,N_3192,N_3138);
or U5964 (N_5964,N_2975,N_4806);
nand U5965 (N_5965,N_3712,N_3332);
or U5966 (N_5966,N_2606,N_4770);
and U5967 (N_5967,N_4091,N_3232);
nor U5968 (N_5968,N_4712,N_4938);
or U5969 (N_5969,N_4759,N_4027);
or U5970 (N_5970,N_3125,N_3102);
nor U5971 (N_5971,N_4624,N_3286);
and U5972 (N_5972,N_4529,N_4415);
nor U5973 (N_5973,N_3043,N_3301);
or U5974 (N_5974,N_2530,N_3063);
nand U5975 (N_5975,N_3253,N_4551);
and U5976 (N_5976,N_2761,N_3079);
and U5977 (N_5977,N_2524,N_3268);
and U5978 (N_5978,N_4040,N_4896);
or U5979 (N_5979,N_3685,N_3212);
xor U5980 (N_5980,N_4674,N_4631);
nor U5981 (N_5981,N_4966,N_4270);
nand U5982 (N_5982,N_3394,N_4007);
and U5983 (N_5983,N_3919,N_4836);
and U5984 (N_5984,N_3111,N_3521);
or U5985 (N_5985,N_4617,N_4083);
nand U5986 (N_5986,N_3077,N_4578);
nand U5987 (N_5987,N_3078,N_2724);
or U5988 (N_5988,N_4880,N_2791);
or U5989 (N_5989,N_4340,N_4839);
and U5990 (N_5990,N_4612,N_2879);
nand U5991 (N_5991,N_3103,N_4520);
xor U5992 (N_5992,N_3909,N_4861);
nand U5993 (N_5993,N_4556,N_4117);
nand U5994 (N_5994,N_3133,N_2754);
nand U5995 (N_5995,N_3211,N_4874);
and U5996 (N_5996,N_4953,N_3305);
and U5997 (N_5997,N_4211,N_3220);
nor U5998 (N_5998,N_4354,N_4777);
nor U5999 (N_5999,N_4470,N_2949);
xnor U6000 (N_6000,N_4838,N_4359);
nand U6001 (N_6001,N_4487,N_2823);
nand U6002 (N_6002,N_4101,N_3707);
and U6003 (N_6003,N_4431,N_4296);
and U6004 (N_6004,N_4146,N_4042);
nor U6005 (N_6005,N_4081,N_3742);
nand U6006 (N_6006,N_2640,N_2916);
and U6007 (N_6007,N_4590,N_4894);
nor U6008 (N_6008,N_3126,N_4689);
or U6009 (N_6009,N_2938,N_3848);
nor U6010 (N_6010,N_4134,N_2682);
and U6011 (N_6011,N_2809,N_4820);
or U6012 (N_6012,N_2548,N_2614);
and U6013 (N_6013,N_3830,N_4028);
or U6014 (N_6014,N_3064,N_3097);
nand U6015 (N_6015,N_3523,N_4738);
and U6016 (N_6016,N_4891,N_4545);
nor U6017 (N_6017,N_3867,N_4823);
nand U6018 (N_6018,N_4471,N_4418);
nand U6019 (N_6019,N_2917,N_2874);
nand U6020 (N_6020,N_3495,N_3724);
nand U6021 (N_6021,N_3954,N_3792);
and U6022 (N_6022,N_3193,N_4761);
or U6023 (N_6023,N_3374,N_2707);
nand U6024 (N_6024,N_3913,N_3046);
and U6025 (N_6025,N_2866,N_4088);
and U6026 (N_6026,N_3771,N_2639);
and U6027 (N_6027,N_3017,N_3030);
nor U6028 (N_6028,N_4965,N_4809);
nor U6029 (N_6029,N_3857,N_3806);
and U6030 (N_6030,N_2627,N_4005);
and U6031 (N_6031,N_3423,N_4997);
xor U6032 (N_6032,N_2734,N_4589);
and U6033 (N_6033,N_3534,N_2667);
nor U6034 (N_6034,N_2719,N_4114);
nor U6035 (N_6035,N_4120,N_3853);
or U6036 (N_6036,N_4294,N_4959);
xnor U6037 (N_6037,N_3710,N_4169);
nand U6038 (N_6038,N_4935,N_2911);
nand U6039 (N_6039,N_2783,N_4754);
nand U6040 (N_6040,N_2844,N_3476);
nand U6041 (N_6041,N_4383,N_4398);
nand U6042 (N_6042,N_2814,N_3772);
or U6043 (N_6043,N_3413,N_2993);
nand U6044 (N_6044,N_3300,N_4221);
nand U6045 (N_6045,N_4059,N_3430);
and U6046 (N_6046,N_4153,N_4584);
and U6047 (N_6047,N_4324,N_4109);
nor U6048 (N_6048,N_4275,N_4452);
or U6049 (N_6049,N_3339,N_2971);
nor U6050 (N_6050,N_2904,N_2941);
nand U6051 (N_6051,N_4709,N_2919);
nand U6052 (N_6052,N_2715,N_3877);
nor U6053 (N_6053,N_4205,N_2695);
nand U6054 (N_6054,N_4603,N_4049);
nand U6055 (N_6055,N_2946,N_2997);
nand U6056 (N_6056,N_4410,N_2638);
and U6057 (N_6057,N_2862,N_3114);
nand U6058 (N_6058,N_4403,N_4931);
and U6059 (N_6059,N_4973,N_3348);
or U6060 (N_6060,N_3472,N_4714);
nand U6061 (N_6061,N_3823,N_3721);
nor U6062 (N_6062,N_4713,N_4098);
and U6063 (N_6063,N_4501,N_3239);
nand U6064 (N_6064,N_4571,N_4218);
or U6065 (N_6065,N_2869,N_2907);
nand U6066 (N_6066,N_3329,N_4478);
nand U6067 (N_6067,N_4517,N_3664);
or U6068 (N_6068,N_3589,N_3336);
or U6069 (N_6069,N_4250,N_2534);
and U6070 (N_6070,N_4033,N_4920);
nand U6071 (N_6071,N_3969,N_3687);
or U6072 (N_6072,N_2964,N_4558);
nor U6073 (N_6073,N_4909,N_3416);
nor U6074 (N_6074,N_3310,N_2972);
or U6075 (N_6075,N_3917,N_2657);
xnor U6076 (N_6076,N_3705,N_4272);
nor U6077 (N_6077,N_4778,N_4382);
and U6078 (N_6078,N_4136,N_2819);
nand U6079 (N_6079,N_3155,N_4414);
and U6080 (N_6080,N_4144,N_2520);
nand U6081 (N_6081,N_3488,N_4273);
nand U6082 (N_6082,N_3828,N_3281);
and U6083 (N_6083,N_4981,N_2793);
or U6084 (N_6084,N_4139,N_2873);
nand U6085 (N_6085,N_2628,N_3490);
nand U6086 (N_6086,N_4549,N_4247);
and U6087 (N_6087,N_4182,N_4803);
and U6088 (N_6088,N_3450,N_3048);
nand U6089 (N_6089,N_4233,N_4580);
or U6090 (N_6090,N_4455,N_4392);
nor U6091 (N_6091,N_4541,N_3763);
nand U6092 (N_6092,N_4905,N_2517);
nor U6093 (N_6093,N_3349,N_4621);
or U6094 (N_6094,N_4393,N_2987);
or U6095 (N_6095,N_2541,N_2803);
and U6096 (N_6096,N_4053,N_3950);
or U6097 (N_6097,N_3072,N_4522);
or U6098 (N_6098,N_2950,N_2739);
or U6099 (N_6099,N_4066,N_3596);
and U6100 (N_6100,N_3174,N_4203);
and U6101 (N_6101,N_4281,N_2801);
nand U6102 (N_6102,N_3199,N_4288);
nor U6103 (N_6103,N_3116,N_4009);
nor U6104 (N_6104,N_4184,N_2813);
or U6105 (N_6105,N_3399,N_3973);
xor U6106 (N_6106,N_4856,N_4581);
nor U6107 (N_6107,N_3674,N_4733);
nor U6108 (N_6108,N_2798,N_4728);
nand U6109 (N_6109,N_4209,N_3873);
or U6110 (N_6110,N_2764,N_3356);
and U6111 (N_6111,N_3247,N_2877);
nor U6112 (N_6112,N_4662,N_3083);
nand U6113 (N_6113,N_2786,N_4977);
nand U6114 (N_6114,N_4892,N_3264);
nand U6115 (N_6115,N_2796,N_4975);
and U6116 (N_6116,N_2637,N_4799);
and U6117 (N_6117,N_4592,N_2888);
and U6118 (N_6118,N_4906,N_4332);
nor U6119 (N_6119,N_4345,N_4537);
or U6120 (N_6120,N_4653,N_3260);
nand U6121 (N_6121,N_2731,N_4881);
nand U6122 (N_6122,N_4246,N_3840);
nor U6123 (N_6123,N_3327,N_3100);
nor U6124 (N_6124,N_4715,N_2708);
and U6125 (N_6125,N_3075,N_3298);
nor U6126 (N_6126,N_3981,N_2518);
and U6127 (N_6127,N_2985,N_4594);
or U6128 (N_6128,N_3235,N_4851);
nand U6129 (N_6129,N_3941,N_4974);
nor U6130 (N_6130,N_4299,N_2853);
nor U6131 (N_6131,N_4442,N_4149);
and U6132 (N_6132,N_4051,N_2947);
or U6133 (N_6133,N_3608,N_4871);
nor U6134 (N_6134,N_3042,N_3104);
nor U6135 (N_6135,N_4889,N_3407);
or U6136 (N_6136,N_3731,N_3068);
and U6137 (N_6137,N_3086,N_4801);
nand U6138 (N_6138,N_3537,N_4427);
nor U6139 (N_6139,N_4980,N_3573);
nand U6140 (N_6140,N_4285,N_3770);
nor U6141 (N_6141,N_4325,N_3259);
and U6142 (N_6142,N_4433,N_2929);
and U6143 (N_6143,N_4743,N_4950);
and U6144 (N_6144,N_2991,N_2891);
nor U6145 (N_6145,N_3673,N_4181);
and U6146 (N_6146,N_4138,N_4562);
nor U6147 (N_6147,N_2825,N_4656);
and U6148 (N_6148,N_2735,N_4527);
nor U6149 (N_6149,N_4476,N_4939);
nor U6150 (N_6150,N_3752,N_3593);
and U6151 (N_6151,N_2537,N_4413);
or U6152 (N_6152,N_3404,N_2815);
or U6153 (N_6153,N_4075,N_4826);
nand U6154 (N_6154,N_4870,N_4800);
xnor U6155 (N_6155,N_3061,N_3396);
or U6156 (N_6156,N_2800,N_4160);
or U6157 (N_6157,N_4473,N_2706);
xor U6158 (N_6158,N_3875,N_3322);
nor U6159 (N_6159,N_2616,N_3530);
and U6160 (N_6160,N_3288,N_4378);
nor U6161 (N_6161,N_3609,N_3021);
and U6162 (N_6162,N_2598,N_3988);
nand U6163 (N_6163,N_3474,N_4055);
or U6164 (N_6164,N_2856,N_3726);
or U6165 (N_6165,N_3607,N_2665);
and U6166 (N_6166,N_4694,N_4536);
or U6167 (N_6167,N_2848,N_4824);
or U6168 (N_6168,N_3143,N_3297);
nand U6169 (N_6169,N_3201,N_2669);
nand U6170 (N_6170,N_4014,N_4239);
or U6171 (N_6171,N_2986,N_4125);
nor U6172 (N_6172,N_4291,N_4195);
nor U6173 (N_6173,N_4384,N_4828);
or U6174 (N_6174,N_3948,N_4816);
or U6175 (N_6175,N_3993,N_4424);
nand U6176 (N_6176,N_4686,N_4220);
nand U6177 (N_6177,N_2889,N_3491);
nand U6178 (N_6178,N_4240,N_3120);
nor U6179 (N_6179,N_3767,N_3481);
nand U6180 (N_6180,N_4787,N_2612);
nor U6181 (N_6181,N_2808,N_4956);
nor U6182 (N_6182,N_4510,N_4940);
and U6183 (N_6183,N_2740,N_4314);
nor U6184 (N_6184,N_3279,N_4850);
nand U6185 (N_6185,N_4084,N_3159);
nand U6186 (N_6186,N_4484,N_3703);
xor U6187 (N_6187,N_2553,N_2703);
nor U6188 (N_6188,N_4070,N_2811);
nand U6189 (N_6189,N_3789,N_3145);
nor U6190 (N_6190,N_4095,N_2623);
nand U6191 (N_6191,N_4356,N_3468);
and U6192 (N_6192,N_2566,N_4924);
or U6193 (N_6193,N_3693,N_4840);
nand U6194 (N_6194,N_3964,N_4772);
and U6195 (N_6195,N_2621,N_4357);
and U6196 (N_6196,N_4877,N_4245);
nor U6197 (N_6197,N_3688,N_2765);
and U6198 (N_6198,N_3334,N_2567);
nor U6199 (N_6199,N_2863,N_4020);
and U6200 (N_6200,N_4740,N_3539);
or U6201 (N_6201,N_4198,N_3518);
or U6202 (N_6202,N_3588,N_4734);
and U6203 (N_6203,N_4208,N_3197);
nand U6204 (N_6204,N_3219,N_3904);
and U6205 (N_6205,N_3499,N_4834);
or U6206 (N_6206,N_4514,N_3453);
and U6207 (N_6207,N_3582,N_3953);
nand U6208 (N_6208,N_3089,N_3206);
or U6209 (N_6209,N_2959,N_3108);
nor U6210 (N_6210,N_2962,N_3280);
and U6211 (N_6211,N_4237,N_4092);
nor U6212 (N_6212,N_3762,N_3389);
nand U6213 (N_6213,N_2978,N_4697);
nor U6214 (N_6214,N_4890,N_3395);
or U6215 (N_6215,N_3088,N_4243);
and U6216 (N_6216,N_3346,N_4791);
and U6217 (N_6217,N_2769,N_4461);
nand U6218 (N_6218,N_4390,N_4263);
nor U6219 (N_6219,N_4365,N_3531);
or U6220 (N_6220,N_2909,N_2982);
and U6221 (N_6221,N_4310,N_3010);
or U6222 (N_6222,N_3690,N_3425);
and U6223 (N_6223,N_3834,N_2531);
and U6224 (N_6224,N_4341,N_4408);
nor U6225 (N_6225,N_2522,N_4264);
and U6226 (N_6226,N_3978,N_2683);
or U6227 (N_6227,N_4248,N_3692);
nand U6228 (N_6228,N_2896,N_3594);
and U6229 (N_6229,N_4063,N_3646);
or U6230 (N_6230,N_2937,N_3535);
and U6231 (N_6231,N_2586,N_4970);
or U6232 (N_6232,N_4781,N_2625);
and U6233 (N_6233,N_4228,N_3185);
nor U6234 (N_6234,N_4369,N_3238);
nor U6235 (N_6235,N_3923,N_3914);
or U6236 (N_6236,N_3342,N_4067);
nand U6237 (N_6237,N_3893,N_4445);
nand U6238 (N_6238,N_4329,N_2728);
or U6239 (N_6239,N_3598,N_3514);
nor U6240 (N_6240,N_3897,N_4654);
or U6241 (N_6241,N_3733,N_4225);
nor U6242 (N_6242,N_4857,N_2689);
or U6243 (N_6243,N_4348,N_3325);
and U6244 (N_6244,N_2599,N_2816);
or U6245 (N_6245,N_4705,N_4984);
nor U6246 (N_6246,N_3858,N_3658);
and U6247 (N_6247,N_4103,N_3388);
nor U6248 (N_6248,N_2799,N_3047);
nor U6249 (N_6249,N_2954,N_4385);
and U6250 (N_6250,N_2564,N_3480);
nand U6251 (N_6251,N_4643,N_3089);
nand U6252 (N_6252,N_3105,N_3820);
nand U6253 (N_6253,N_2757,N_4969);
nand U6254 (N_6254,N_3932,N_4781);
and U6255 (N_6255,N_4152,N_4453);
nor U6256 (N_6256,N_4042,N_3630);
nor U6257 (N_6257,N_4902,N_4830);
nand U6258 (N_6258,N_4185,N_3794);
nor U6259 (N_6259,N_3903,N_4519);
nand U6260 (N_6260,N_2585,N_2554);
nand U6261 (N_6261,N_4959,N_4963);
or U6262 (N_6262,N_4448,N_3837);
or U6263 (N_6263,N_3846,N_4993);
xor U6264 (N_6264,N_4307,N_3227);
and U6265 (N_6265,N_3523,N_4875);
nor U6266 (N_6266,N_2607,N_4024);
nor U6267 (N_6267,N_4025,N_2846);
xor U6268 (N_6268,N_3087,N_4065);
nand U6269 (N_6269,N_2840,N_2529);
nand U6270 (N_6270,N_2686,N_4159);
or U6271 (N_6271,N_2695,N_2932);
xor U6272 (N_6272,N_3425,N_4222);
nor U6273 (N_6273,N_4391,N_4100);
or U6274 (N_6274,N_3226,N_3111);
nand U6275 (N_6275,N_4415,N_4236);
or U6276 (N_6276,N_2587,N_4146);
nand U6277 (N_6277,N_4870,N_4700);
nor U6278 (N_6278,N_3988,N_3233);
or U6279 (N_6279,N_3509,N_4771);
and U6280 (N_6280,N_4796,N_2581);
nand U6281 (N_6281,N_4396,N_2887);
or U6282 (N_6282,N_4062,N_3239);
and U6283 (N_6283,N_3470,N_3919);
nor U6284 (N_6284,N_4178,N_3825);
and U6285 (N_6285,N_4615,N_4484);
nand U6286 (N_6286,N_2705,N_4309);
nor U6287 (N_6287,N_2517,N_3988);
xor U6288 (N_6288,N_4415,N_4028);
nand U6289 (N_6289,N_2806,N_3976);
nand U6290 (N_6290,N_2513,N_3429);
and U6291 (N_6291,N_3307,N_4326);
nand U6292 (N_6292,N_2658,N_2836);
nand U6293 (N_6293,N_4171,N_3482);
nand U6294 (N_6294,N_3968,N_3978);
and U6295 (N_6295,N_4735,N_3343);
and U6296 (N_6296,N_2740,N_4066);
or U6297 (N_6297,N_4897,N_3111);
nand U6298 (N_6298,N_4848,N_4654);
nor U6299 (N_6299,N_4292,N_3164);
nor U6300 (N_6300,N_3197,N_3787);
nor U6301 (N_6301,N_4975,N_4331);
nand U6302 (N_6302,N_2934,N_2647);
xnor U6303 (N_6303,N_3250,N_4246);
or U6304 (N_6304,N_3915,N_3855);
nor U6305 (N_6305,N_2691,N_3209);
nor U6306 (N_6306,N_4481,N_2651);
nor U6307 (N_6307,N_3589,N_3325);
nand U6308 (N_6308,N_3872,N_2657);
or U6309 (N_6309,N_4735,N_2984);
or U6310 (N_6310,N_4736,N_4302);
nor U6311 (N_6311,N_3544,N_3063);
nor U6312 (N_6312,N_3347,N_3039);
and U6313 (N_6313,N_2838,N_4687);
and U6314 (N_6314,N_4080,N_3724);
nor U6315 (N_6315,N_4150,N_2890);
and U6316 (N_6316,N_2638,N_2591);
nor U6317 (N_6317,N_2719,N_2933);
and U6318 (N_6318,N_4636,N_3714);
or U6319 (N_6319,N_4646,N_4606);
nand U6320 (N_6320,N_3425,N_4396);
nor U6321 (N_6321,N_2697,N_4488);
nor U6322 (N_6322,N_4666,N_4701);
nor U6323 (N_6323,N_3824,N_3508);
xor U6324 (N_6324,N_3669,N_3402);
and U6325 (N_6325,N_3662,N_4319);
and U6326 (N_6326,N_3061,N_3176);
nand U6327 (N_6327,N_3447,N_3961);
and U6328 (N_6328,N_3259,N_4482);
nand U6329 (N_6329,N_2760,N_3375);
nand U6330 (N_6330,N_3536,N_4571);
and U6331 (N_6331,N_4477,N_4248);
nand U6332 (N_6332,N_3159,N_3870);
nor U6333 (N_6333,N_2761,N_4376);
nor U6334 (N_6334,N_4384,N_4876);
nor U6335 (N_6335,N_3976,N_2622);
or U6336 (N_6336,N_4272,N_3003);
and U6337 (N_6337,N_4127,N_4562);
nor U6338 (N_6338,N_4456,N_3812);
or U6339 (N_6339,N_3614,N_4551);
and U6340 (N_6340,N_4339,N_4662);
xnor U6341 (N_6341,N_4444,N_2952);
and U6342 (N_6342,N_4691,N_3363);
and U6343 (N_6343,N_2749,N_3701);
nand U6344 (N_6344,N_2802,N_3134);
nand U6345 (N_6345,N_2780,N_2955);
nand U6346 (N_6346,N_2853,N_3709);
and U6347 (N_6347,N_4086,N_2805);
nor U6348 (N_6348,N_2692,N_2894);
nor U6349 (N_6349,N_3852,N_4111);
nand U6350 (N_6350,N_4850,N_3953);
nor U6351 (N_6351,N_3103,N_2990);
or U6352 (N_6352,N_2667,N_2896);
or U6353 (N_6353,N_4287,N_4524);
or U6354 (N_6354,N_2500,N_4073);
or U6355 (N_6355,N_4151,N_4540);
nor U6356 (N_6356,N_3766,N_2709);
or U6357 (N_6357,N_3198,N_4772);
and U6358 (N_6358,N_3245,N_3727);
or U6359 (N_6359,N_4869,N_4617);
nand U6360 (N_6360,N_3748,N_4051);
xor U6361 (N_6361,N_3385,N_4916);
and U6362 (N_6362,N_3451,N_3920);
nor U6363 (N_6363,N_3345,N_3177);
nor U6364 (N_6364,N_3898,N_4132);
nand U6365 (N_6365,N_3572,N_4041);
nor U6366 (N_6366,N_3638,N_4767);
nand U6367 (N_6367,N_2878,N_2777);
and U6368 (N_6368,N_3316,N_4627);
or U6369 (N_6369,N_3697,N_2869);
or U6370 (N_6370,N_3254,N_4411);
and U6371 (N_6371,N_3933,N_4055);
and U6372 (N_6372,N_3261,N_4116);
or U6373 (N_6373,N_4933,N_3622);
nand U6374 (N_6374,N_3325,N_4245);
nand U6375 (N_6375,N_4561,N_3957);
or U6376 (N_6376,N_3814,N_2609);
nand U6377 (N_6377,N_4499,N_4884);
nand U6378 (N_6378,N_4041,N_4730);
or U6379 (N_6379,N_4156,N_4290);
and U6380 (N_6380,N_4452,N_3644);
nand U6381 (N_6381,N_4063,N_2917);
nand U6382 (N_6382,N_3912,N_3215);
or U6383 (N_6383,N_3531,N_4638);
and U6384 (N_6384,N_3379,N_2557);
xnor U6385 (N_6385,N_3119,N_4947);
or U6386 (N_6386,N_3601,N_2753);
nor U6387 (N_6387,N_3747,N_3388);
or U6388 (N_6388,N_3908,N_3952);
nor U6389 (N_6389,N_4636,N_4525);
or U6390 (N_6390,N_2880,N_3172);
nand U6391 (N_6391,N_4236,N_2975);
or U6392 (N_6392,N_2557,N_3743);
or U6393 (N_6393,N_4184,N_4305);
or U6394 (N_6394,N_4302,N_3713);
or U6395 (N_6395,N_2541,N_3463);
and U6396 (N_6396,N_3550,N_3088);
or U6397 (N_6397,N_2576,N_2980);
nor U6398 (N_6398,N_3473,N_4965);
nand U6399 (N_6399,N_4481,N_4102);
and U6400 (N_6400,N_3298,N_4236);
or U6401 (N_6401,N_4965,N_4011);
or U6402 (N_6402,N_4723,N_3489);
nand U6403 (N_6403,N_4418,N_2531);
or U6404 (N_6404,N_3167,N_4755);
and U6405 (N_6405,N_4425,N_4632);
nor U6406 (N_6406,N_2825,N_3984);
and U6407 (N_6407,N_4602,N_4923);
nor U6408 (N_6408,N_4537,N_4740);
nor U6409 (N_6409,N_4441,N_3205);
nor U6410 (N_6410,N_3799,N_3237);
nor U6411 (N_6411,N_2872,N_4872);
and U6412 (N_6412,N_3603,N_3513);
nor U6413 (N_6413,N_3573,N_2634);
and U6414 (N_6414,N_4812,N_4380);
or U6415 (N_6415,N_4176,N_3506);
and U6416 (N_6416,N_3914,N_3965);
nand U6417 (N_6417,N_4307,N_3848);
or U6418 (N_6418,N_3394,N_4418);
nor U6419 (N_6419,N_2800,N_2711);
or U6420 (N_6420,N_3318,N_3036);
and U6421 (N_6421,N_4059,N_2843);
and U6422 (N_6422,N_4907,N_2542);
nor U6423 (N_6423,N_3656,N_4951);
and U6424 (N_6424,N_4892,N_3029);
and U6425 (N_6425,N_2988,N_4899);
or U6426 (N_6426,N_4032,N_4478);
nor U6427 (N_6427,N_2908,N_3661);
or U6428 (N_6428,N_3443,N_2510);
and U6429 (N_6429,N_3402,N_4626);
and U6430 (N_6430,N_3435,N_3952);
or U6431 (N_6431,N_3671,N_4227);
and U6432 (N_6432,N_4160,N_2588);
and U6433 (N_6433,N_3916,N_2707);
nor U6434 (N_6434,N_3907,N_3170);
and U6435 (N_6435,N_2777,N_3771);
nand U6436 (N_6436,N_3846,N_2675);
or U6437 (N_6437,N_4243,N_4493);
or U6438 (N_6438,N_2856,N_3014);
or U6439 (N_6439,N_3475,N_4399);
or U6440 (N_6440,N_3458,N_2733);
xor U6441 (N_6441,N_4098,N_4668);
nand U6442 (N_6442,N_3763,N_4987);
xor U6443 (N_6443,N_4859,N_3963);
or U6444 (N_6444,N_4470,N_4109);
or U6445 (N_6445,N_4710,N_3265);
or U6446 (N_6446,N_3039,N_4553);
or U6447 (N_6447,N_4226,N_3140);
and U6448 (N_6448,N_4994,N_3900);
nor U6449 (N_6449,N_3322,N_3024);
and U6450 (N_6450,N_4724,N_2861);
or U6451 (N_6451,N_3142,N_2906);
or U6452 (N_6452,N_4267,N_3057);
and U6453 (N_6453,N_4695,N_3137);
and U6454 (N_6454,N_2579,N_3228);
nor U6455 (N_6455,N_3688,N_4999);
nor U6456 (N_6456,N_3436,N_3686);
and U6457 (N_6457,N_4579,N_4363);
nor U6458 (N_6458,N_4984,N_3638);
or U6459 (N_6459,N_3523,N_4615);
xor U6460 (N_6460,N_4538,N_3038);
xnor U6461 (N_6461,N_4019,N_2699);
or U6462 (N_6462,N_2661,N_3514);
or U6463 (N_6463,N_4073,N_3650);
nor U6464 (N_6464,N_2950,N_3277);
nand U6465 (N_6465,N_3867,N_2639);
or U6466 (N_6466,N_3293,N_3916);
xnor U6467 (N_6467,N_3625,N_4706);
nor U6468 (N_6468,N_4566,N_4400);
and U6469 (N_6469,N_2776,N_3704);
nand U6470 (N_6470,N_4995,N_4334);
xor U6471 (N_6471,N_2798,N_4229);
or U6472 (N_6472,N_2760,N_4059);
or U6473 (N_6473,N_3275,N_3859);
nand U6474 (N_6474,N_3806,N_4741);
nor U6475 (N_6475,N_2689,N_3827);
and U6476 (N_6476,N_4001,N_3304);
nand U6477 (N_6477,N_2981,N_2938);
nor U6478 (N_6478,N_3883,N_2640);
and U6479 (N_6479,N_4599,N_4471);
nor U6480 (N_6480,N_3845,N_4063);
and U6481 (N_6481,N_4603,N_3855);
or U6482 (N_6482,N_4974,N_2953);
nor U6483 (N_6483,N_4874,N_3414);
or U6484 (N_6484,N_3655,N_4754);
nand U6485 (N_6485,N_2955,N_3685);
nand U6486 (N_6486,N_2731,N_3157);
nor U6487 (N_6487,N_3882,N_3051);
nor U6488 (N_6488,N_4724,N_3173);
nor U6489 (N_6489,N_4606,N_3188);
and U6490 (N_6490,N_3386,N_4250);
and U6491 (N_6491,N_4367,N_2687);
nand U6492 (N_6492,N_4452,N_4408);
and U6493 (N_6493,N_3994,N_2841);
or U6494 (N_6494,N_4096,N_3236);
nor U6495 (N_6495,N_2535,N_2628);
nor U6496 (N_6496,N_3142,N_4469);
nand U6497 (N_6497,N_3722,N_4245);
or U6498 (N_6498,N_4019,N_2702);
xor U6499 (N_6499,N_3232,N_2899);
nor U6500 (N_6500,N_3975,N_4879);
nand U6501 (N_6501,N_2631,N_2618);
and U6502 (N_6502,N_3802,N_3002);
or U6503 (N_6503,N_3780,N_2965);
nor U6504 (N_6504,N_2698,N_2559);
nor U6505 (N_6505,N_3454,N_3282);
nand U6506 (N_6506,N_4981,N_3454);
nand U6507 (N_6507,N_3706,N_3509);
and U6508 (N_6508,N_4530,N_3137);
nand U6509 (N_6509,N_3336,N_2756);
and U6510 (N_6510,N_4604,N_4994);
nor U6511 (N_6511,N_3907,N_4229);
nand U6512 (N_6512,N_4430,N_2758);
or U6513 (N_6513,N_3844,N_3358);
nor U6514 (N_6514,N_4806,N_3275);
nand U6515 (N_6515,N_3446,N_2969);
or U6516 (N_6516,N_3359,N_3826);
or U6517 (N_6517,N_4771,N_2923);
or U6518 (N_6518,N_3957,N_4749);
and U6519 (N_6519,N_4659,N_3277);
or U6520 (N_6520,N_3916,N_4149);
and U6521 (N_6521,N_3852,N_3809);
nor U6522 (N_6522,N_4040,N_3891);
nand U6523 (N_6523,N_4743,N_3516);
nor U6524 (N_6524,N_4556,N_3553);
nor U6525 (N_6525,N_4707,N_3864);
nor U6526 (N_6526,N_4309,N_4790);
nand U6527 (N_6527,N_3548,N_4442);
and U6528 (N_6528,N_4373,N_3110);
or U6529 (N_6529,N_3529,N_4170);
nand U6530 (N_6530,N_4136,N_4745);
nor U6531 (N_6531,N_2859,N_2981);
and U6532 (N_6532,N_2741,N_3218);
nor U6533 (N_6533,N_3856,N_3786);
nor U6534 (N_6534,N_3683,N_3552);
nor U6535 (N_6535,N_3061,N_3938);
or U6536 (N_6536,N_3994,N_4041);
or U6537 (N_6537,N_2971,N_4401);
or U6538 (N_6538,N_2799,N_4833);
or U6539 (N_6539,N_2890,N_4660);
nor U6540 (N_6540,N_3476,N_4028);
and U6541 (N_6541,N_4821,N_2995);
and U6542 (N_6542,N_3970,N_3225);
nor U6543 (N_6543,N_3447,N_2516);
xnor U6544 (N_6544,N_3024,N_3553);
or U6545 (N_6545,N_2790,N_2882);
nand U6546 (N_6546,N_3743,N_3859);
and U6547 (N_6547,N_4802,N_2687);
nor U6548 (N_6548,N_2662,N_4958);
and U6549 (N_6549,N_4144,N_4138);
or U6550 (N_6550,N_4741,N_4392);
nor U6551 (N_6551,N_4799,N_3825);
nor U6552 (N_6552,N_4907,N_4471);
and U6553 (N_6553,N_2937,N_4872);
or U6554 (N_6554,N_2972,N_3752);
or U6555 (N_6555,N_2832,N_4046);
or U6556 (N_6556,N_4121,N_4087);
nand U6557 (N_6557,N_2943,N_3840);
nand U6558 (N_6558,N_4940,N_3241);
and U6559 (N_6559,N_4879,N_2706);
nand U6560 (N_6560,N_3741,N_4597);
or U6561 (N_6561,N_3910,N_4643);
nand U6562 (N_6562,N_2732,N_4200);
and U6563 (N_6563,N_4980,N_4511);
or U6564 (N_6564,N_3137,N_2508);
nand U6565 (N_6565,N_3921,N_3404);
nand U6566 (N_6566,N_4139,N_4893);
and U6567 (N_6567,N_4081,N_3654);
nand U6568 (N_6568,N_4848,N_4305);
or U6569 (N_6569,N_2822,N_2595);
nor U6570 (N_6570,N_2693,N_3474);
nand U6571 (N_6571,N_4952,N_3030);
or U6572 (N_6572,N_4799,N_3741);
nand U6573 (N_6573,N_3618,N_3404);
nand U6574 (N_6574,N_3384,N_3297);
nor U6575 (N_6575,N_3066,N_4845);
nand U6576 (N_6576,N_2642,N_4618);
and U6577 (N_6577,N_3115,N_3247);
and U6578 (N_6578,N_4367,N_4560);
and U6579 (N_6579,N_3590,N_3064);
and U6580 (N_6580,N_4807,N_3694);
nor U6581 (N_6581,N_3806,N_4570);
and U6582 (N_6582,N_3170,N_4824);
nor U6583 (N_6583,N_4894,N_4749);
or U6584 (N_6584,N_3982,N_3736);
nor U6585 (N_6585,N_3551,N_4410);
nor U6586 (N_6586,N_3196,N_2601);
or U6587 (N_6587,N_3730,N_3313);
nand U6588 (N_6588,N_4038,N_4450);
nor U6589 (N_6589,N_4651,N_2971);
or U6590 (N_6590,N_4897,N_2544);
nor U6591 (N_6591,N_4510,N_4639);
nor U6592 (N_6592,N_3314,N_4897);
nor U6593 (N_6593,N_3292,N_3387);
nor U6594 (N_6594,N_3073,N_3916);
nand U6595 (N_6595,N_2925,N_4814);
or U6596 (N_6596,N_4876,N_4141);
and U6597 (N_6597,N_4550,N_2571);
nor U6598 (N_6598,N_2666,N_2926);
or U6599 (N_6599,N_4676,N_4458);
nand U6600 (N_6600,N_4630,N_4537);
nor U6601 (N_6601,N_3634,N_4961);
or U6602 (N_6602,N_4215,N_4170);
and U6603 (N_6603,N_3756,N_3142);
or U6604 (N_6604,N_4782,N_4549);
nor U6605 (N_6605,N_3220,N_3344);
or U6606 (N_6606,N_3010,N_4716);
nand U6607 (N_6607,N_2959,N_3877);
or U6608 (N_6608,N_3631,N_4326);
or U6609 (N_6609,N_3738,N_4159);
or U6610 (N_6610,N_3581,N_4920);
nor U6611 (N_6611,N_3057,N_3828);
nand U6612 (N_6612,N_4723,N_3754);
or U6613 (N_6613,N_4848,N_2747);
nand U6614 (N_6614,N_4199,N_3096);
nand U6615 (N_6615,N_4025,N_3003);
nor U6616 (N_6616,N_3166,N_3773);
and U6617 (N_6617,N_3067,N_3101);
and U6618 (N_6618,N_2849,N_2660);
or U6619 (N_6619,N_4655,N_3295);
or U6620 (N_6620,N_4304,N_3074);
xor U6621 (N_6621,N_3766,N_3806);
or U6622 (N_6622,N_4153,N_2680);
nor U6623 (N_6623,N_4621,N_4758);
nand U6624 (N_6624,N_4042,N_2875);
and U6625 (N_6625,N_3233,N_4171);
nor U6626 (N_6626,N_3750,N_3182);
nor U6627 (N_6627,N_4320,N_2762);
and U6628 (N_6628,N_4830,N_4510);
or U6629 (N_6629,N_4634,N_4256);
nand U6630 (N_6630,N_4115,N_4334);
or U6631 (N_6631,N_3536,N_2736);
or U6632 (N_6632,N_2676,N_4470);
nand U6633 (N_6633,N_4346,N_3635);
and U6634 (N_6634,N_4042,N_4607);
xor U6635 (N_6635,N_4184,N_4443);
and U6636 (N_6636,N_2524,N_3562);
and U6637 (N_6637,N_3973,N_2629);
or U6638 (N_6638,N_3423,N_2992);
or U6639 (N_6639,N_4997,N_3219);
nor U6640 (N_6640,N_3528,N_2674);
nand U6641 (N_6641,N_2983,N_4485);
or U6642 (N_6642,N_2562,N_3054);
nand U6643 (N_6643,N_4374,N_2649);
or U6644 (N_6644,N_4710,N_3440);
nor U6645 (N_6645,N_3959,N_3404);
and U6646 (N_6646,N_3263,N_3657);
nand U6647 (N_6647,N_3665,N_2700);
nor U6648 (N_6648,N_3752,N_4140);
or U6649 (N_6649,N_2687,N_2635);
nor U6650 (N_6650,N_3338,N_3279);
and U6651 (N_6651,N_3191,N_4243);
nand U6652 (N_6652,N_3479,N_4510);
and U6653 (N_6653,N_3251,N_3335);
xor U6654 (N_6654,N_4790,N_2645);
nand U6655 (N_6655,N_4134,N_2985);
nand U6656 (N_6656,N_2889,N_4492);
nor U6657 (N_6657,N_4286,N_3679);
nand U6658 (N_6658,N_3593,N_3033);
nor U6659 (N_6659,N_2955,N_2908);
and U6660 (N_6660,N_4777,N_2788);
nand U6661 (N_6661,N_2742,N_4145);
nor U6662 (N_6662,N_4861,N_2709);
and U6663 (N_6663,N_3591,N_3597);
nand U6664 (N_6664,N_4533,N_2773);
nor U6665 (N_6665,N_4093,N_3848);
and U6666 (N_6666,N_2721,N_3227);
nor U6667 (N_6667,N_4277,N_3173);
or U6668 (N_6668,N_4767,N_3558);
or U6669 (N_6669,N_2720,N_4328);
and U6670 (N_6670,N_4041,N_4322);
or U6671 (N_6671,N_4170,N_3442);
or U6672 (N_6672,N_3665,N_4452);
nor U6673 (N_6673,N_4556,N_3001);
and U6674 (N_6674,N_4560,N_3616);
and U6675 (N_6675,N_4938,N_3110);
or U6676 (N_6676,N_3430,N_2524);
and U6677 (N_6677,N_4074,N_3558);
nor U6678 (N_6678,N_4448,N_3458);
xnor U6679 (N_6679,N_4090,N_3855);
nor U6680 (N_6680,N_4667,N_3792);
and U6681 (N_6681,N_3727,N_4282);
nand U6682 (N_6682,N_4814,N_2624);
and U6683 (N_6683,N_3567,N_3915);
xnor U6684 (N_6684,N_3242,N_4185);
nand U6685 (N_6685,N_3390,N_3946);
nand U6686 (N_6686,N_4498,N_2822);
nand U6687 (N_6687,N_2513,N_4673);
nor U6688 (N_6688,N_3624,N_3641);
and U6689 (N_6689,N_3312,N_3811);
nand U6690 (N_6690,N_3326,N_2765);
nand U6691 (N_6691,N_2789,N_3686);
nand U6692 (N_6692,N_3933,N_4702);
nand U6693 (N_6693,N_3485,N_2833);
or U6694 (N_6694,N_4982,N_2526);
nand U6695 (N_6695,N_4584,N_3310);
and U6696 (N_6696,N_4941,N_3340);
nor U6697 (N_6697,N_2710,N_3428);
and U6698 (N_6698,N_2760,N_3616);
nand U6699 (N_6699,N_3099,N_2826);
and U6700 (N_6700,N_4703,N_2699);
nor U6701 (N_6701,N_3767,N_3022);
or U6702 (N_6702,N_4578,N_4221);
nor U6703 (N_6703,N_3702,N_3845);
nor U6704 (N_6704,N_4718,N_2626);
or U6705 (N_6705,N_4888,N_4993);
nor U6706 (N_6706,N_4716,N_3774);
nand U6707 (N_6707,N_3236,N_3216);
and U6708 (N_6708,N_2544,N_2854);
and U6709 (N_6709,N_3489,N_4639);
or U6710 (N_6710,N_3080,N_4633);
nand U6711 (N_6711,N_3886,N_3739);
or U6712 (N_6712,N_2840,N_2548);
or U6713 (N_6713,N_4259,N_3676);
or U6714 (N_6714,N_4259,N_3527);
and U6715 (N_6715,N_3256,N_2690);
and U6716 (N_6716,N_4141,N_2868);
or U6717 (N_6717,N_3855,N_4361);
nor U6718 (N_6718,N_4488,N_2880);
nand U6719 (N_6719,N_4461,N_4360);
or U6720 (N_6720,N_4807,N_4953);
nor U6721 (N_6721,N_4689,N_4642);
nor U6722 (N_6722,N_3753,N_3685);
or U6723 (N_6723,N_2532,N_2701);
and U6724 (N_6724,N_2945,N_4429);
nor U6725 (N_6725,N_4746,N_3622);
or U6726 (N_6726,N_3020,N_4298);
or U6727 (N_6727,N_3540,N_4458);
nand U6728 (N_6728,N_2819,N_4352);
or U6729 (N_6729,N_4204,N_4679);
and U6730 (N_6730,N_2640,N_3650);
nand U6731 (N_6731,N_3635,N_3318);
nand U6732 (N_6732,N_4844,N_4216);
or U6733 (N_6733,N_4194,N_4284);
or U6734 (N_6734,N_4250,N_3080);
nand U6735 (N_6735,N_4341,N_4618);
nor U6736 (N_6736,N_3508,N_3020);
nor U6737 (N_6737,N_3517,N_3765);
nor U6738 (N_6738,N_3434,N_3845);
nand U6739 (N_6739,N_3668,N_4566);
nand U6740 (N_6740,N_2713,N_3781);
or U6741 (N_6741,N_2773,N_3919);
nor U6742 (N_6742,N_4844,N_4287);
nand U6743 (N_6743,N_3818,N_3598);
nor U6744 (N_6744,N_4562,N_2744);
or U6745 (N_6745,N_3185,N_4022);
nor U6746 (N_6746,N_4488,N_3166);
and U6747 (N_6747,N_3963,N_4045);
and U6748 (N_6748,N_4969,N_4102);
xor U6749 (N_6749,N_3549,N_4964);
nand U6750 (N_6750,N_3135,N_3002);
nand U6751 (N_6751,N_3409,N_3257);
and U6752 (N_6752,N_4855,N_3690);
or U6753 (N_6753,N_2825,N_3336);
and U6754 (N_6754,N_3224,N_4807);
xnor U6755 (N_6755,N_3636,N_2610);
or U6756 (N_6756,N_4727,N_4000);
or U6757 (N_6757,N_3156,N_3953);
nor U6758 (N_6758,N_3431,N_2790);
or U6759 (N_6759,N_4493,N_2822);
or U6760 (N_6760,N_3593,N_2892);
xor U6761 (N_6761,N_2844,N_4130);
and U6762 (N_6762,N_4529,N_3218);
nor U6763 (N_6763,N_3204,N_3239);
and U6764 (N_6764,N_3489,N_3247);
nand U6765 (N_6765,N_3768,N_4227);
and U6766 (N_6766,N_3532,N_4601);
nand U6767 (N_6767,N_4853,N_4896);
nand U6768 (N_6768,N_3550,N_3727);
or U6769 (N_6769,N_3677,N_4425);
and U6770 (N_6770,N_3871,N_4129);
xnor U6771 (N_6771,N_4718,N_3070);
or U6772 (N_6772,N_2974,N_4524);
or U6773 (N_6773,N_3685,N_3516);
nand U6774 (N_6774,N_2500,N_3200);
nor U6775 (N_6775,N_4288,N_2946);
and U6776 (N_6776,N_3972,N_4301);
nand U6777 (N_6777,N_4710,N_3927);
nor U6778 (N_6778,N_2954,N_3365);
or U6779 (N_6779,N_4435,N_2632);
or U6780 (N_6780,N_4490,N_3636);
nand U6781 (N_6781,N_3116,N_3333);
nand U6782 (N_6782,N_3682,N_4050);
nor U6783 (N_6783,N_3178,N_4405);
nor U6784 (N_6784,N_3373,N_3545);
nand U6785 (N_6785,N_2703,N_2799);
and U6786 (N_6786,N_3645,N_4371);
nor U6787 (N_6787,N_2834,N_3241);
nor U6788 (N_6788,N_3954,N_3213);
nor U6789 (N_6789,N_4014,N_4142);
nand U6790 (N_6790,N_4917,N_4843);
or U6791 (N_6791,N_3987,N_3393);
or U6792 (N_6792,N_4580,N_3269);
xnor U6793 (N_6793,N_3023,N_4185);
nand U6794 (N_6794,N_3223,N_3462);
and U6795 (N_6795,N_3009,N_4262);
nand U6796 (N_6796,N_3720,N_3063);
and U6797 (N_6797,N_3233,N_3855);
nor U6798 (N_6798,N_2512,N_3147);
xnor U6799 (N_6799,N_3213,N_2614);
and U6800 (N_6800,N_2980,N_2720);
and U6801 (N_6801,N_4778,N_3491);
nand U6802 (N_6802,N_2924,N_2507);
or U6803 (N_6803,N_3820,N_3595);
or U6804 (N_6804,N_3888,N_2529);
nand U6805 (N_6805,N_4919,N_4461);
nor U6806 (N_6806,N_3185,N_3167);
or U6807 (N_6807,N_3370,N_2880);
nor U6808 (N_6808,N_4899,N_4924);
nand U6809 (N_6809,N_4079,N_3766);
nor U6810 (N_6810,N_3944,N_2532);
or U6811 (N_6811,N_2966,N_4058);
and U6812 (N_6812,N_3312,N_4836);
nor U6813 (N_6813,N_4397,N_2526);
or U6814 (N_6814,N_4473,N_2629);
and U6815 (N_6815,N_3373,N_4253);
and U6816 (N_6816,N_3772,N_2868);
nand U6817 (N_6817,N_2707,N_3731);
xor U6818 (N_6818,N_4879,N_3704);
or U6819 (N_6819,N_2694,N_2731);
or U6820 (N_6820,N_4025,N_3890);
and U6821 (N_6821,N_3784,N_3444);
nand U6822 (N_6822,N_3235,N_3964);
or U6823 (N_6823,N_4947,N_4836);
and U6824 (N_6824,N_3770,N_4764);
and U6825 (N_6825,N_4325,N_3009);
or U6826 (N_6826,N_4341,N_4811);
and U6827 (N_6827,N_3156,N_4983);
and U6828 (N_6828,N_2888,N_4737);
nor U6829 (N_6829,N_2658,N_2707);
nor U6830 (N_6830,N_2843,N_4848);
nand U6831 (N_6831,N_4615,N_4778);
and U6832 (N_6832,N_2521,N_4966);
and U6833 (N_6833,N_4535,N_2636);
nand U6834 (N_6834,N_3890,N_2653);
or U6835 (N_6835,N_2774,N_3071);
and U6836 (N_6836,N_2582,N_3330);
or U6837 (N_6837,N_4287,N_2541);
and U6838 (N_6838,N_2812,N_2811);
or U6839 (N_6839,N_3766,N_2896);
and U6840 (N_6840,N_4979,N_4399);
or U6841 (N_6841,N_4141,N_3026);
nand U6842 (N_6842,N_4345,N_4045);
nand U6843 (N_6843,N_3331,N_4134);
nor U6844 (N_6844,N_4312,N_3676);
and U6845 (N_6845,N_3525,N_4906);
nand U6846 (N_6846,N_4047,N_4499);
and U6847 (N_6847,N_3623,N_4118);
nand U6848 (N_6848,N_2797,N_2950);
and U6849 (N_6849,N_3939,N_3430);
nor U6850 (N_6850,N_2609,N_4957);
or U6851 (N_6851,N_4419,N_3018);
or U6852 (N_6852,N_4965,N_3695);
nand U6853 (N_6853,N_3972,N_3803);
and U6854 (N_6854,N_2542,N_2701);
nand U6855 (N_6855,N_4030,N_3316);
or U6856 (N_6856,N_3269,N_3089);
and U6857 (N_6857,N_2551,N_4840);
or U6858 (N_6858,N_2975,N_3097);
nor U6859 (N_6859,N_4835,N_3053);
nand U6860 (N_6860,N_3581,N_3482);
and U6861 (N_6861,N_2732,N_4472);
and U6862 (N_6862,N_3434,N_2770);
xnor U6863 (N_6863,N_2522,N_4117);
xnor U6864 (N_6864,N_4634,N_3517);
nand U6865 (N_6865,N_3438,N_3868);
and U6866 (N_6866,N_2602,N_3795);
and U6867 (N_6867,N_3820,N_4059);
nor U6868 (N_6868,N_4644,N_4741);
nand U6869 (N_6869,N_2644,N_3475);
nor U6870 (N_6870,N_3491,N_4970);
nor U6871 (N_6871,N_2817,N_3171);
or U6872 (N_6872,N_3901,N_2610);
nand U6873 (N_6873,N_3066,N_4783);
and U6874 (N_6874,N_4806,N_3860);
or U6875 (N_6875,N_3113,N_4194);
and U6876 (N_6876,N_4472,N_4752);
nor U6877 (N_6877,N_4954,N_4969);
nor U6878 (N_6878,N_2762,N_4359);
and U6879 (N_6879,N_4049,N_3568);
or U6880 (N_6880,N_2954,N_2915);
nor U6881 (N_6881,N_4516,N_3680);
and U6882 (N_6882,N_3665,N_3297);
nor U6883 (N_6883,N_3057,N_3839);
nor U6884 (N_6884,N_3105,N_2996);
nand U6885 (N_6885,N_4392,N_3808);
or U6886 (N_6886,N_4080,N_4371);
nand U6887 (N_6887,N_2639,N_4126);
and U6888 (N_6888,N_4611,N_3591);
and U6889 (N_6889,N_2958,N_3834);
nand U6890 (N_6890,N_4794,N_3695);
nor U6891 (N_6891,N_4142,N_4632);
nor U6892 (N_6892,N_3619,N_3090);
nor U6893 (N_6893,N_4190,N_3613);
and U6894 (N_6894,N_2949,N_4996);
nand U6895 (N_6895,N_4112,N_4653);
or U6896 (N_6896,N_3697,N_4433);
nor U6897 (N_6897,N_4327,N_4971);
and U6898 (N_6898,N_3790,N_4320);
nor U6899 (N_6899,N_3064,N_3269);
or U6900 (N_6900,N_4943,N_3325);
or U6901 (N_6901,N_4390,N_3138);
nor U6902 (N_6902,N_3699,N_4464);
nor U6903 (N_6903,N_4109,N_4585);
nor U6904 (N_6904,N_3620,N_4392);
and U6905 (N_6905,N_4905,N_3850);
nor U6906 (N_6906,N_3794,N_2906);
nor U6907 (N_6907,N_2832,N_3203);
xnor U6908 (N_6908,N_2827,N_3176);
or U6909 (N_6909,N_4333,N_4035);
or U6910 (N_6910,N_4430,N_3607);
nor U6911 (N_6911,N_4848,N_4681);
nand U6912 (N_6912,N_2786,N_4726);
nor U6913 (N_6913,N_3803,N_4942);
nand U6914 (N_6914,N_3556,N_4580);
or U6915 (N_6915,N_2935,N_4951);
nor U6916 (N_6916,N_2813,N_3025);
nand U6917 (N_6917,N_3875,N_3673);
nand U6918 (N_6918,N_3427,N_3823);
or U6919 (N_6919,N_3318,N_4834);
or U6920 (N_6920,N_4179,N_4660);
or U6921 (N_6921,N_3964,N_2607);
nor U6922 (N_6922,N_3921,N_2792);
nand U6923 (N_6923,N_3958,N_4878);
nand U6924 (N_6924,N_4782,N_3846);
or U6925 (N_6925,N_3448,N_3332);
and U6926 (N_6926,N_2541,N_3553);
nand U6927 (N_6927,N_4007,N_4232);
or U6928 (N_6928,N_2569,N_4902);
nor U6929 (N_6929,N_4484,N_2729);
or U6930 (N_6930,N_3745,N_2606);
nor U6931 (N_6931,N_4234,N_2770);
and U6932 (N_6932,N_4465,N_2852);
and U6933 (N_6933,N_2670,N_2790);
nor U6934 (N_6934,N_3313,N_3252);
nand U6935 (N_6935,N_3133,N_4323);
nand U6936 (N_6936,N_3257,N_2527);
and U6937 (N_6937,N_3145,N_2714);
nor U6938 (N_6938,N_4759,N_2646);
and U6939 (N_6939,N_2983,N_2959);
and U6940 (N_6940,N_4738,N_2924);
nor U6941 (N_6941,N_3423,N_3526);
nand U6942 (N_6942,N_3146,N_4963);
nor U6943 (N_6943,N_3072,N_2918);
nand U6944 (N_6944,N_4339,N_4816);
nand U6945 (N_6945,N_3712,N_3595);
and U6946 (N_6946,N_3318,N_2672);
and U6947 (N_6947,N_3128,N_4937);
or U6948 (N_6948,N_3649,N_3177);
or U6949 (N_6949,N_4407,N_3519);
and U6950 (N_6950,N_3987,N_4565);
nor U6951 (N_6951,N_4049,N_4493);
and U6952 (N_6952,N_2634,N_3020);
nand U6953 (N_6953,N_3540,N_3644);
nand U6954 (N_6954,N_4864,N_4293);
and U6955 (N_6955,N_2588,N_4377);
nor U6956 (N_6956,N_3388,N_3318);
nor U6957 (N_6957,N_3551,N_4798);
nor U6958 (N_6958,N_3272,N_3973);
and U6959 (N_6959,N_3040,N_3229);
and U6960 (N_6960,N_4672,N_2593);
and U6961 (N_6961,N_4911,N_3151);
nor U6962 (N_6962,N_4506,N_2868);
nor U6963 (N_6963,N_2503,N_3031);
nand U6964 (N_6964,N_3792,N_3288);
nor U6965 (N_6965,N_3465,N_2542);
and U6966 (N_6966,N_4796,N_3124);
nor U6967 (N_6967,N_3322,N_4096);
or U6968 (N_6968,N_2567,N_4996);
nor U6969 (N_6969,N_4469,N_3738);
and U6970 (N_6970,N_3642,N_3300);
and U6971 (N_6971,N_4802,N_4300);
xor U6972 (N_6972,N_3819,N_3699);
xnor U6973 (N_6973,N_2598,N_2670);
and U6974 (N_6974,N_3750,N_4567);
and U6975 (N_6975,N_3253,N_3914);
nand U6976 (N_6976,N_2503,N_2675);
or U6977 (N_6977,N_3770,N_4661);
nand U6978 (N_6978,N_4153,N_3748);
and U6979 (N_6979,N_3895,N_4175);
nand U6980 (N_6980,N_2932,N_4031);
and U6981 (N_6981,N_4723,N_2515);
nor U6982 (N_6982,N_3793,N_4346);
nand U6983 (N_6983,N_3858,N_4199);
nor U6984 (N_6984,N_2722,N_3226);
and U6985 (N_6985,N_2598,N_3841);
nand U6986 (N_6986,N_4325,N_3531);
nor U6987 (N_6987,N_4791,N_2687);
nand U6988 (N_6988,N_2777,N_3206);
nand U6989 (N_6989,N_4416,N_4626);
nand U6990 (N_6990,N_3457,N_4865);
or U6991 (N_6991,N_3915,N_2822);
nor U6992 (N_6992,N_4771,N_4547);
nor U6993 (N_6993,N_2964,N_3170);
nor U6994 (N_6994,N_3256,N_2946);
nand U6995 (N_6995,N_3710,N_3049);
nand U6996 (N_6996,N_3238,N_3798);
or U6997 (N_6997,N_4260,N_4883);
or U6998 (N_6998,N_3577,N_3906);
nand U6999 (N_6999,N_3354,N_3443);
or U7000 (N_7000,N_4487,N_2822);
nand U7001 (N_7001,N_3457,N_3514);
nand U7002 (N_7002,N_3959,N_4536);
nand U7003 (N_7003,N_4579,N_4711);
or U7004 (N_7004,N_4292,N_3399);
nor U7005 (N_7005,N_3981,N_4692);
nand U7006 (N_7006,N_4165,N_4304);
nor U7007 (N_7007,N_3536,N_2607);
xnor U7008 (N_7008,N_2533,N_4128);
nor U7009 (N_7009,N_3108,N_2581);
or U7010 (N_7010,N_3094,N_3168);
and U7011 (N_7011,N_4664,N_4157);
nand U7012 (N_7012,N_4795,N_2818);
nand U7013 (N_7013,N_3808,N_3107);
and U7014 (N_7014,N_3539,N_3487);
nand U7015 (N_7015,N_3094,N_3907);
or U7016 (N_7016,N_3626,N_4523);
or U7017 (N_7017,N_3089,N_2528);
and U7018 (N_7018,N_2804,N_3124);
xor U7019 (N_7019,N_2932,N_2883);
or U7020 (N_7020,N_4669,N_3565);
or U7021 (N_7021,N_2943,N_3566);
nand U7022 (N_7022,N_3408,N_4599);
or U7023 (N_7023,N_2913,N_3065);
nand U7024 (N_7024,N_4450,N_3664);
or U7025 (N_7025,N_2799,N_2784);
or U7026 (N_7026,N_3642,N_4995);
and U7027 (N_7027,N_4129,N_3143);
and U7028 (N_7028,N_3463,N_3892);
nor U7029 (N_7029,N_3736,N_2945);
and U7030 (N_7030,N_3582,N_4414);
and U7031 (N_7031,N_4125,N_4775);
and U7032 (N_7032,N_4884,N_4635);
nor U7033 (N_7033,N_4147,N_3205);
and U7034 (N_7034,N_4998,N_2982);
nand U7035 (N_7035,N_3405,N_2737);
and U7036 (N_7036,N_4374,N_3371);
or U7037 (N_7037,N_2901,N_2579);
and U7038 (N_7038,N_4892,N_4538);
or U7039 (N_7039,N_2918,N_3936);
and U7040 (N_7040,N_3274,N_3779);
and U7041 (N_7041,N_2847,N_3365);
nand U7042 (N_7042,N_4181,N_3832);
xor U7043 (N_7043,N_2934,N_4994);
nor U7044 (N_7044,N_3445,N_2843);
or U7045 (N_7045,N_4344,N_3676);
or U7046 (N_7046,N_4879,N_3675);
nand U7047 (N_7047,N_4671,N_4896);
and U7048 (N_7048,N_3070,N_3068);
nand U7049 (N_7049,N_3883,N_4904);
or U7050 (N_7050,N_3614,N_3650);
and U7051 (N_7051,N_2727,N_3012);
nor U7052 (N_7052,N_3593,N_3252);
nand U7053 (N_7053,N_3078,N_3480);
nand U7054 (N_7054,N_2657,N_3016);
nor U7055 (N_7055,N_4717,N_3629);
nor U7056 (N_7056,N_3543,N_3973);
and U7057 (N_7057,N_4361,N_2614);
nand U7058 (N_7058,N_4687,N_3710);
xnor U7059 (N_7059,N_2681,N_4465);
nor U7060 (N_7060,N_4479,N_3979);
nand U7061 (N_7061,N_3016,N_2796);
nor U7062 (N_7062,N_3007,N_2612);
or U7063 (N_7063,N_3143,N_3808);
or U7064 (N_7064,N_3970,N_3583);
and U7065 (N_7065,N_3606,N_3114);
and U7066 (N_7066,N_4584,N_4526);
nand U7067 (N_7067,N_3448,N_3925);
or U7068 (N_7068,N_4861,N_2916);
nand U7069 (N_7069,N_3478,N_4007);
and U7070 (N_7070,N_4777,N_3453);
nor U7071 (N_7071,N_3569,N_2679);
or U7072 (N_7072,N_4041,N_3620);
or U7073 (N_7073,N_4825,N_4329);
nand U7074 (N_7074,N_4801,N_3923);
and U7075 (N_7075,N_3274,N_4634);
or U7076 (N_7076,N_2898,N_4588);
nor U7077 (N_7077,N_4157,N_3251);
nor U7078 (N_7078,N_3680,N_2924);
nand U7079 (N_7079,N_3544,N_3447);
nand U7080 (N_7080,N_4298,N_2763);
nand U7081 (N_7081,N_3497,N_3752);
and U7082 (N_7082,N_2979,N_4176);
and U7083 (N_7083,N_4688,N_4693);
nor U7084 (N_7084,N_4640,N_4066);
nor U7085 (N_7085,N_4966,N_4482);
and U7086 (N_7086,N_3262,N_3862);
nor U7087 (N_7087,N_2816,N_4166);
nand U7088 (N_7088,N_3023,N_3291);
or U7089 (N_7089,N_3620,N_2748);
and U7090 (N_7090,N_3857,N_3559);
or U7091 (N_7091,N_4387,N_2855);
nand U7092 (N_7092,N_4802,N_4886);
and U7093 (N_7093,N_4545,N_3485);
xnor U7094 (N_7094,N_4011,N_3140);
nand U7095 (N_7095,N_4629,N_2898);
and U7096 (N_7096,N_4533,N_2547);
nor U7097 (N_7097,N_4235,N_3810);
nand U7098 (N_7098,N_4787,N_4087);
or U7099 (N_7099,N_3447,N_2831);
nand U7100 (N_7100,N_4651,N_3441);
nor U7101 (N_7101,N_4573,N_4366);
nand U7102 (N_7102,N_4377,N_4069);
nor U7103 (N_7103,N_2577,N_4508);
and U7104 (N_7104,N_4649,N_2691);
and U7105 (N_7105,N_4812,N_4084);
nand U7106 (N_7106,N_2814,N_3149);
nand U7107 (N_7107,N_3558,N_3280);
nand U7108 (N_7108,N_3713,N_3359);
xor U7109 (N_7109,N_3967,N_4583);
and U7110 (N_7110,N_2777,N_2873);
or U7111 (N_7111,N_4167,N_4917);
nor U7112 (N_7112,N_3286,N_4466);
or U7113 (N_7113,N_4857,N_4583);
nor U7114 (N_7114,N_3778,N_4548);
and U7115 (N_7115,N_3053,N_3763);
nor U7116 (N_7116,N_3655,N_3581);
nand U7117 (N_7117,N_3765,N_4252);
xor U7118 (N_7118,N_3939,N_2821);
nand U7119 (N_7119,N_2559,N_2515);
nand U7120 (N_7120,N_4154,N_3651);
nor U7121 (N_7121,N_3764,N_2789);
and U7122 (N_7122,N_4555,N_3794);
and U7123 (N_7123,N_4891,N_4929);
and U7124 (N_7124,N_2793,N_4670);
or U7125 (N_7125,N_3598,N_4942);
or U7126 (N_7126,N_3606,N_3981);
nor U7127 (N_7127,N_3765,N_4952);
nand U7128 (N_7128,N_3485,N_3738);
or U7129 (N_7129,N_4625,N_4419);
or U7130 (N_7130,N_3490,N_3793);
nand U7131 (N_7131,N_3759,N_3843);
nor U7132 (N_7132,N_3079,N_3395);
nor U7133 (N_7133,N_2720,N_2773);
xnor U7134 (N_7134,N_4672,N_4740);
or U7135 (N_7135,N_3701,N_4154);
nor U7136 (N_7136,N_2986,N_4580);
nand U7137 (N_7137,N_4401,N_4564);
nor U7138 (N_7138,N_4791,N_3226);
or U7139 (N_7139,N_4875,N_3129);
nor U7140 (N_7140,N_3925,N_3843);
nand U7141 (N_7141,N_3049,N_3556);
nand U7142 (N_7142,N_4860,N_3704);
nand U7143 (N_7143,N_3237,N_3747);
and U7144 (N_7144,N_3475,N_3420);
and U7145 (N_7145,N_4288,N_4728);
nand U7146 (N_7146,N_3795,N_3490);
nor U7147 (N_7147,N_2735,N_3550);
nand U7148 (N_7148,N_4193,N_3732);
and U7149 (N_7149,N_3294,N_3573);
or U7150 (N_7150,N_2823,N_4272);
nor U7151 (N_7151,N_3097,N_4708);
and U7152 (N_7152,N_4295,N_4199);
or U7153 (N_7153,N_3938,N_4431);
and U7154 (N_7154,N_2624,N_2742);
and U7155 (N_7155,N_3616,N_3495);
nand U7156 (N_7156,N_3726,N_3236);
or U7157 (N_7157,N_3853,N_4315);
and U7158 (N_7158,N_2867,N_3625);
nor U7159 (N_7159,N_4556,N_3715);
nand U7160 (N_7160,N_3390,N_4334);
nor U7161 (N_7161,N_3488,N_3093);
and U7162 (N_7162,N_4379,N_3523);
and U7163 (N_7163,N_3921,N_2766);
or U7164 (N_7164,N_2578,N_3529);
or U7165 (N_7165,N_3538,N_4212);
nor U7166 (N_7166,N_4358,N_3818);
and U7167 (N_7167,N_3687,N_4102);
nor U7168 (N_7168,N_3675,N_4055);
xor U7169 (N_7169,N_3247,N_3796);
or U7170 (N_7170,N_3345,N_3244);
xnor U7171 (N_7171,N_4793,N_3456);
nand U7172 (N_7172,N_4245,N_4443);
nor U7173 (N_7173,N_3526,N_3778);
and U7174 (N_7174,N_4974,N_4825);
or U7175 (N_7175,N_4339,N_4158);
xnor U7176 (N_7176,N_4784,N_3076);
and U7177 (N_7177,N_3484,N_2922);
nor U7178 (N_7178,N_4920,N_4850);
and U7179 (N_7179,N_3053,N_4952);
nand U7180 (N_7180,N_3199,N_3837);
nand U7181 (N_7181,N_2671,N_4698);
or U7182 (N_7182,N_3435,N_3731);
or U7183 (N_7183,N_4946,N_3285);
nor U7184 (N_7184,N_3702,N_3245);
and U7185 (N_7185,N_4763,N_4854);
nand U7186 (N_7186,N_3296,N_4343);
nor U7187 (N_7187,N_3204,N_4634);
or U7188 (N_7188,N_2518,N_4148);
and U7189 (N_7189,N_4904,N_4651);
or U7190 (N_7190,N_4004,N_3997);
nand U7191 (N_7191,N_3507,N_2660);
nand U7192 (N_7192,N_2898,N_3074);
and U7193 (N_7193,N_4989,N_4661);
and U7194 (N_7194,N_3667,N_4009);
and U7195 (N_7195,N_3951,N_3688);
and U7196 (N_7196,N_3970,N_4750);
nand U7197 (N_7197,N_4959,N_3069);
nand U7198 (N_7198,N_4464,N_4087);
nand U7199 (N_7199,N_2957,N_3076);
nor U7200 (N_7200,N_2517,N_4773);
and U7201 (N_7201,N_3192,N_4511);
nand U7202 (N_7202,N_3161,N_2601);
nor U7203 (N_7203,N_4394,N_3543);
nand U7204 (N_7204,N_3081,N_4651);
and U7205 (N_7205,N_3092,N_3270);
or U7206 (N_7206,N_3440,N_3586);
or U7207 (N_7207,N_3205,N_2717);
and U7208 (N_7208,N_3031,N_3563);
and U7209 (N_7209,N_4620,N_3222);
and U7210 (N_7210,N_4168,N_3543);
nand U7211 (N_7211,N_4090,N_4347);
nand U7212 (N_7212,N_4456,N_4406);
xnor U7213 (N_7213,N_3640,N_3179);
or U7214 (N_7214,N_3320,N_4621);
nor U7215 (N_7215,N_4751,N_4745);
and U7216 (N_7216,N_2686,N_4031);
nand U7217 (N_7217,N_3193,N_4082);
and U7218 (N_7218,N_3511,N_4280);
and U7219 (N_7219,N_4274,N_3218);
or U7220 (N_7220,N_4484,N_3508);
and U7221 (N_7221,N_3052,N_2898);
nor U7222 (N_7222,N_3305,N_3233);
or U7223 (N_7223,N_4397,N_3849);
nor U7224 (N_7224,N_2723,N_4837);
nand U7225 (N_7225,N_2797,N_4167);
nand U7226 (N_7226,N_4657,N_4135);
and U7227 (N_7227,N_2678,N_4161);
or U7228 (N_7228,N_3785,N_3783);
nand U7229 (N_7229,N_3255,N_3302);
or U7230 (N_7230,N_3076,N_4301);
or U7231 (N_7231,N_4330,N_3842);
or U7232 (N_7232,N_3910,N_4626);
nand U7233 (N_7233,N_3897,N_4852);
or U7234 (N_7234,N_3338,N_4934);
nor U7235 (N_7235,N_2679,N_4297);
nand U7236 (N_7236,N_3155,N_4359);
nor U7237 (N_7237,N_4259,N_3118);
nor U7238 (N_7238,N_4856,N_4147);
and U7239 (N_7239,N_4846,N_2639);
nor U7240 (N_7240,N_3337,N_3721);
or U7241 (N_7241,N_2821,N_4346);
nor U7242 (N_7242,N_2925,N_3585);
nor U7243 (N_7243,N_2552,N_4633);
nor U7244 (N_7244,N_3020,N_3625);
nand U7245 (N_7245,N_3254,N_2744);
nand U7246 (N_7246,N_2728,N_4266);
or U7247 (N_7247,N_3011,N_3165);
xor U7248 (N_7248,N_2923,N_3619);
nand U7249 (N_7249,N_3926,N_2979);
nor U7250 (N_7250,N_3627,N_2704);
and U7251 (N_7251,N_4539,N_3186);
nand U7252 (N_7252,N_4414,N_3427);
nand U7253 (N_7253,N_3957,N_4712);
nor U7254 (N_7254,N_3320,N_4588);
xnor U7255 (N_7255,N_3007,N_2749);
nor U7256 (N_7256,N_2657,N_4221);
or U7257 (N_7257,N_4923,N_2543);
xor U7258 (N_7258,N_4935,N_3820);
nor U7259 (N_7259,N_3628,N_3703);
nor U7260 (N_7260,N_3602,N_3672);
and U7261 (N_7261,N_4761,N_3425);
or U7262 (N_7262,N_3528,N_3770);
nor U7263 (N_7263,N_4047,N_4947);
nor U7264 (N_7264,N_2740,N_3323);
or U7265 (N_7265,N_2650,N_2817);
and U7266 (N_7266,N_4186,N_3601);
or U7267 (N_7267,N_3441,N_2875);
or U7268 (N_7268,N_3912,N_4974);
xor U7269 (N_7269,N_3699,N_3572);
nand U7270 (N_7270,N_3885,N_3984);
nand U7271 (N_7271,N_4112,N_2797);
or U7272 (N_7272,N_4244,N_4220);
or U7273 (N_7273,N_3790,N_2559);
or U7274 (N_7274,N_2528,N_4101);
and U7275 (N_7275,N_3554,N_4711);
and U7276 (N_7276,N_4807,N_4637);
or U7277 (N_7277,N_3800,N_3964);
nor U7278 (N_7278,N_2589,N_3457);
nand U7279 (N_7279,N_3505,N_3164);
nand U7280 (N_7280,N_3117,N_3167);
and U7281 (N_7281,N_2583,N_3034);
and U7282 (N_7282,N_3449,N_3015);
or U7283 (N_7283,N_4460,N_2539);
nand U7284 (N_7284,N_2888,N_4629);
or U7285 (N_7285,N_3442,N_4147);
and U7286 (N_7286,N_3105,N_4855);
or U7287 (N_7287,N_4204,N_3389);
xor U7288 (N_7288,N_3218,N_3002);
nand U7289 (N_7289,N_4111,N_3616);
nand U7290 (N_7290,N_4838,N_3258);
and U7291 (N_7291,N_4174,N_3984);
or U7292 (N_7292,N_3006,N_4994);
and U7293 (N_7293,N_3502,N_4879);
and U7294 (N_7294,N_2780,N_3911);
xnor U7295 (N_7295,N_4374,N_4571);
nand U7296 (N_7296,N_2994,N_3462);
nor U7297 (N_7297,N_3092,N_4372);
or U7298 (N_7298,N_2743,N_4937);
or U7299 (N_7299,N_2835,N_4106);
and U7300 (N_7300,N_2664,N_3076);
nor U7301 (N_7301,N_4531,N_3008);
or U7302 (N_7302,N_4483,N_4092);
or U7303 (N_7303,N_4850,N_4434);
nor U7304 (N_7304,N_3417,N_4211);
nor U7305 (N_7305,N_3778,N_3638);
nor U7306 (N_7306,N_3139,N_3400);
nor U7307 (N_7307,N_2775,N_4525);
and U7308 (N_7308,N_4885,N_4333);
or U7309 (N_7309,N_3163,N_2801);
nor U7310 (N_7310,N_4962,N_2946);
nor U7311 (N_7311,N_3626,N_2835);
or U7312 (N_7312,N_2700,N_3357);
nor U7313 (N_7313,N_4866,N_2917);
and U7314 (N_7314,N_4843,N_4303);
nand U7315 (N_7315,N_4306,N_2655);
nor U7316 (N_7316,N_4342,N_4512);
or U7317 (N_7317,N_2702,N_4935);
nand U7318 (N_7318,N_3599,N_4139);
nand U7319 (N_7319,N_4107,N_2957);
nand U7320 (N_7320,N_3058,N_3656);
or U7321 (N_7321,N_4442,N_4976);
or U7322 (N_7322,N_2638,N_4110);
or U7323 (N_7323,N_3790,N_4590);
xor U7324 (N_7324,N_2722,N_3852);
and U7325 (N_7325,N_4436,N_3909);
or U7326 (N_7326,N_4008,N_3812);
nor U7327 (N_7327,N_2670,N_2587);
nor U7328 (N_7328,N_3522,N_4986);
nand U7329 (N_7329,N_3972,N_4807);
nor U7330 (N_7330,N_2810,N_4869);
and U7331 (N_7331,N_3892,N_4047);
nor U7332 (N_7332,N_3768,N_4709);
or U7333 (N_7333,N_4604,N_4939);
nand U7334 (N_7334,N_4794,N_4245);
nand U7335 (N_7335,N_2862,N_2957);
xor U7336 (N_7336,N_4135,N_4570);
xor U7337 (N_7337,N_4902,N_3233);
nand U7338 (N_7338,N_3134,N_4795);
nor U7339 (N_7339,N_4192,N_2548);
and U7340 (N_7340,N_4496,N_4916);
or U7341 (N_7341,N_4228,N_4642);
nor U7342 (N_7342,N_2660,N_4061);
or U7343 (N_7343,N_4836,N_3755);
nand U7344 (N_7344,N_3428,N_4780);
and U7345 (N_7345,N_3841,N_4104);
and U7346 (N_7346,N_3614,N_2639);
nor U7347 (N_7347,N_4813,N_4416);
nor U7348 (N_7348,N_3622,N_3617);
nand U7349 (N_7349,N_4360,N_2874);
and U7350 (N_7350,N_3423,N_4024);
and U7351 (N_7351,N_2568,N_4782);
and U7352 (N_7352,N_2505,N_4547);
and U7353 (N_7353,N_3218,N_2684);
or U7354 (N_7354,N_3748,N_3450);
or U7355 (N_7355,N_3795,N_3670);
nand U7356 (N_7356,N_3371,N_2633);
or U7357 (N_7357,N_3455,N_4844);
nor U7358 (N_7358,N_3592,N_2575);
and U7359 (N_7359,N_2759,N_2857);
nand U7360 (N_7360,N_2709,N_4448);
and U7361 (N_7361,N_3841,N_3167);
and U7362 (N_7362,N_3624,N_4815);
and U7363 (N_7363,N_2968,N_3159);
or U7364 (N_7364,N_3344,N_3121);
and U7365 (N_7365,N_3364,N_3281);
and U7366 (N_7366,N_4908,N_4400);
nor U7367 (N_7367,N_4076,N_4369);
nor U7368 (N_7368,N_2737,N_2969);
or U7369 (N_7369,N_4009,N_3912);
nand U7370 (N_7370,N_3511,N_4730);
nor U7371 (N_7371,N_3698,N_4586);
nand U7372 (N_7372,N_2634,N_3983);
nand U7373 (N_7373,N_3829,N_3352);
or U7374 (N_7374,N_3650,N_4149);
nand U7375 (N_7375,N_3057,N_4935);
nor U7376 (N_7376,N_4677,N_2777);
and U7377 (N_7377,N_3360,N_4831);
nor U7378 (N_7378,N_4240,N_2903);
and U7379 (N_7379,N_4169,N_3687);
nor U7380 (N_7380,N_3178,N_3710);
nand U7381 (N_7381,N_2565,N_4728);
nand U7382 (N_7382,N_2966,N_3426);
nand U7383 (N_7383,N_4002,N_3800);
and U7384 (N_7384,N_4172,N_4340);
nor U7385 (N_7385,N_4486,N_3476);
and U7386 (N_7386,N_2692,N_4276);
or U7387 (N_7387,N_2789,N_3657);
nand U7388 (N_7388,N_4081,N_4448);
and U7389 (N_7389,N_3454,N_4657);
and U7390 (N_7390,N_3778,N_3143);
nor U7391 (N_7391,N_2763,N_3716);
nand U7392 (N_7392,N_3587,N_3655);
or U7393 (N_7393,N_4878,N_3018);
xnor U7394 (N_7394,N_4790,N_3413);
or U7395 (N_7395,N_3444,N_3810);
and U7396 (N_7396,N_3289,N_3043);
nor U7397 (N_7397,N_3959,N_2799);
or U7398 (N_7398,N_3263,N_3415);
nand U7399 (N_7399,N_2650,N_4506);
nor U7400 (N_7400,N_3986,N_2679);
nand U7401 (N_7401,N_2778,N_4177);
nand U7402 (N_7402,N_2836,N_4973);
nor U7403 (N_7403,N_4015,N_2539);
or U7404 (N_7404,N_3424,N_4368);
and U7405 (N_7405,N_4622,N_2983);
xnor U7406 (N_7406,N_4952,N_4165);
and U7407 (N_7407,N_3142,N_4128);
nor U7408 (N_7408,N_4142,N_3240);
nand U7409 (N_7409,N_4502,N_3019);
nor U7410 (N_7410,N_3615,N_3297);
and U7411 (N_7411,N_4915,N_4520);
nor U7412 (N_7412,N_2508,N_3733);
nor U7413 (N_7413,N_4843,N_2928);
nand U7414 (N_7414,N_3866,N_4976);
and U7415 (N_7415,N_4346,N_4551);
and U7416 (N_7416,N_4320,N_3580);
or U7417 (N_7417,N_4398,N_4698);
and U7418 (N_7418,N_3726,N_4707);
nand U7419 (N_7419,N_3365,N_2974);
and U7420 (N_7420,N_2768,N_2728);
or U7421 (N_7421,N_2906,N_4918);
nand U7422 (N_7422,N_2701,N_3182);
and U7423 (N_7423,N_3051,N_4787);
nor U7424 (N_7424,N_2903,N_3892);
nor U7425 (N_7425,N_3991,N_3540);
and U7426 (N_7426,N_4725,N_2890);
nand U7427 (N_7427,N_3888,N_2984);
and U7428 (N_7428,N_2704,N_3230);
or U7429 (N_7429,N_3918,N_4925);
and U7430 (N_7430,N_4275,N_3979);
nand U7431 (N_7431,N_4061,N_4387);
nand U7432 (N_7432,N_3303,N_4079);
nor U7433 (N_7433,N_3775,N_3484);
and U7434 (N_7434,N_3357,N_4130);
or U7435 (N_7435,N_2952,N_4804);
nor U7436 (N_7436,N_4459,N_4885);
or U7437 (N_7437,N_4262,N_3907);
nor U7438 (N_7438,N_3741,N_3250);
or U7439 (N_7439,N_2917,N_4603);
nand U7440 (N_7440,N_3373,N_3010);
or U7441 (N_7441,N_2741,N_4354);
nor U7442 (N_7442,N_3607,N_4315);
and U7443 (N_7443,N_2520,N_2925);
or U7444 (N_7444,N_2868,N_3329);
nor U7445 (N_7445,N_4106,N_3104);
nor U7446 (N_7446,N_4778,N_4579);
nor U7447 (N_7447,N_4495,N_4164);
and U7448 (N_7448,N_3530,N_4792);
and U7449 (N_7449,N_4462,N_3137);
or U7450 (N_7450,N_3891,N_2828);
nand U7451 (N_7451,N_4204,N_3628);
or U7452 (N_7452,N_2528,N_2814);
and U7453 (N_7453,N_2883,N_2717);
or U7454 (N_7454,N_2803,N_3704);
or U7455 (N_7455,N_4469,N_3734);
xor U7456 (N_7456,N_2804,N_4062);
and U7457 (N_7457,N_3467,N_4134);
or U7458 (N_7458,N_3369,N_4843);
nor U7459 (N_7459,N_2726,N_4785);
nor U7460 (N_7460,N_4404,N_3528);
nor U7461 (N_7461,N_2566,N_3064);
nor U7462 (N_7462,N_2927,N_4251);
and U7463 (N_7463,N_4179,N_3811);
and U7464 (N_7464,N_2927,N_4190);
or U7465 (N_7465,N_2889,N_3752);
nand U7466 (N_7466,N_3600,N_4202);
or U7467 (N_7467,N_3634,N_4934);
and U7468 (N_7468,N_4240,N_3862);
nor U7469 (N_7469,N_4201,N_2747);
and U7470 (N_7470,N_3299,N_4893);
nor U7471 (N_7471,N_2709,N_4556);
nand U7472 (N_7472,N_3514,N_4679);
or U7473 (N_7473,N_3044,N_3735);
nand U7474 (N_7474,N_3930,N_4322);
and U7475 (N_7475,N_2776,N_4934);
nand U7476 (N_7476,N_2760,N_2911);
nor U7477 (N_7477,N_3224,N_4498);
and U7478 (N_7478,N_4133,N_3422);
nor U7479 (N_7479,N_2517,N_2725);
nor U7480 (N_7480,N_3867,N_4682);
or U7481 (N_7481,N_4970,N_2703);
nor U7482 (N_7482,N_2805,N_3893);
nand U7483 (N_7483,N_2716,N_3549);
nor U7484 (N_7484,N_2682,N_4335);
nand U7485 (N_7485,N_3533,N_4077);
or U7486 (N_7486,N_2656,N_4863);
and U7487 (N_7487,N_4164,N_4190);
and U7488 (N_7488,N_3111,N_3081);
and U7489 (N_7489,N_4947,N_4841);
nand U7490 (N_7490,N_4474,N_3766);
and U7491 (N_7491,N_3931,N_2635);
and U7492 (N_7492,N_2759,N_2998);
nor U7493 (N_7493,N_2912,N_4168);
nor U7494 (N_7494,N_3571,N_4019);
nand U7495 (N_7495,N_4155,N_3651);
nand U7496 (N_7496,N_3918,N_2744);
nand U7497 (N_7497,N_3404,N_3557);
nand U7498 (N_7498,N_2946,N_4562);
or U7499 (N_7499,N_4298,N_3839);
and U7500 (N_7500,N_7262,N_6604);
or U7501 (N_7501,N_5638,N_6237);
and U7502 (N_7502,N_5240,N_5797);
xor U7503 (N_7503,N_7415,N_5479);
or U7504 (N_7504,N_6578,N_5072);
or U7505 (N_7505,N_7128,N_6505);
nand U7506 (N_7506,N_5192,N_6636);
or U7507 (N_7507,N_5695,N_6534);
nor U7508 (N_7508,N_6934,N_6542);
and U7509 (N_7509,N_7086,N_6721);
nand U7510 (N_7510,N_6343,N_6651);
nor U7511 (N_7511,N_6995,N_5074);
nand U7512 (N_7512,N_7364,N_7179);
or U7513 (N_7513,N_7202,N_7399);
nand U7514 (N_7514,N_7337,N_6277);
nand U7515 (N_7515,N_5759,N_5398);
nor U7516 (N_7516,N_6949,N_5238);
nor U7517 (N_7517,N_5308,N_5891);
or U7518 (N_7518,N_6445,N_6801);
nand U7519 (N_7519,N_7455,N_6839);
nor U7520 (N_7520,N_6361,N_6427);
nand U7521 (N_7521,N_5813,N_6381);
nand U7522 (N_7522,N_5449,N_6051);
nand U7523 (N_7523,N_6832,N_5447);
nor U7524 (N_7524,N_5288,N_7053);
and U7525 (N_7525,N_5836,N_7037);
nand U7526 (N_7526,N_6073,N_6002);
or U7527 (N_7527,N_7171,N_5597);
nor U7528 (N_7528,N_6273,N_6777);
nor U7529 (N_7529,N_6570,N_5041);
nand U7530 (N_7530,N_7453,N_7347);
and U7531 (N_7531,N_6559,N_5877);
nand U7532 (N_7532,N_5027,N_5939);
nand U7533 (N_7533,N_6853,N_7191);
or U7534 (N_7534,N_5468,N_7088);
nand U7535 (N_7535,N_5576,N_5421);
nand U7536 (N_7536,N_5665,N_7106);
or U7537 (N_7537,N_5451,N_5102);
nand U7538 (N_7538,N_5352,N_7494);
and U7539 (N_7539,N_5431,N_5679);
and U7540 (N_7540,N_6883,N_6618);
nor U7541 (N_7541,N_5965,N_5754);
or U7542 (N_7542,N_7110,N_6911);
nor U7543 (N_7543,N_6720,N_5146);
nand U7544 (N_7544,N_6018,N_6300);
nand U7545 (N_7545,N_6345,N_7094);
nand U7546 (N_7546,N_6201,N_6518);
nand U7547 (N_7547,N_6411,N_6414);
or U7548 (N_7548,N_7416,N_7411);
nand U7549 (N_7549,N_5198,N_6535);
and U7550 (N_7550,N_7165,N_7275);
or U7551 (N_7551,N_7158,N_5795);
or U7552 (N_7552,N_6962,N_6096);
or U7553 (N_7553,N_7184,N_7019);
or U7554 (N_7554,N_5129,N_7488);
and U7555 (N_7555,N_5315,N_7427);
or U7556 (N_7556,N_5881,N_6066);
nand U7557 (N_7557,N_7187,N_6887);
nor U7558 (N_7558,N_6819,N_7002);
nand U7559 (N_7559,N_6019,N_6866);
nand U7560 (N_7560,N_6267,N_7402);
nand U7561 (N_7561,N_7318,N_5310);
nor U7562 (N_7562,N_6010,N_5437);
or U7563 (N_7563,N_5219,N_5339);
and U7564 (N_7564,N_5271,N_5211);
and U7565 (N_7565,N_6617,N_7324);
nor U7566 (N_7566,N_5770,N_5247);
or U7567 (N_7567,N_6101,N_7480);
nand U7568 (N_7568,N_6791,N_5483);
nor U7569 (N_7569,N_5212,N_6841);
nor U7570 (N_7570,N_5716,N_6288);
or U7571 (N_7571,N_6067,N_5751);
nand U7572 (N_7572,N_5208,N_7109);
nand U7573 (N_7573,N_6403,N_6211);
nand U7574 (N_7574,N_5189,N_6616);
and U7575 (N_7575,N_5166,N_6865);
and U7576 (N_7576,N_5739,N_7119);
nand U7577 (N_7577,N_5486,N_5096);
or U7578 (N_7578,N_6392,N_6823);
nand U7579 (N_7579,N_7495,N_5251);
and U7580 (N_7580,N_5843,N_7290);
or U7581 (N_7581,N_5426,N_5188);
nor U7582 (N_7582,N_6289,N_5897);
nor U7583 (N_7583,N_5320,N_5345);
or U7584 (N_7584,N_7349,N_5856);
nand U7585 (N_7585,N_7295,N_5017);
or U7586 (N_7586,N_6528,N_6407);
nor U7587 (N_7587,N_6303,N_6961);
nand U7588 (N_7588,N_7172,N_5623);
nor U7589 (N_7589,N_5839,N_6881);
and U7590 (N_7590,N_5557,N_6703);
or U7591 (N_7591,N_7438,N_7242);
nand U7592 (N_7592,N_7093,N_5454);
and U7593 (N_7593,N_5349,N_5976);
nand U7594 (N_7594,N_5996,N_6146);
and U7595 (N_7595,N_5299,N_5061);
or U7596 (N_7596,N_6382,N_6847);
and U7597 (N_7597,N_6647,N_6863);
and U7598 (N_7598,N_6362,N_6608);
and U7599 (N_7599,N_6488,N_5448);
nand U7600 (N_7600,N_6151,N_6170);
and U7601 (N_7601,N_6149,N_6543);
and U7602 (N_7602,N_5190,N_6432);
or U7603 (N_7603,N_5572,N_5667);
or U7604 (N_7604,N_7247,N_7439);
or U7605 (N_7605,N_6610,N_5579);
xor U7606 (N_7606,N_5379,N_7329);
nor U7607 (N_7607,N_5408,N_6972);
nand U7608 (N_7608,N_5539,N_6276);
and U7609 (N_7609,N_5782,N_5199);
nor U7610 (N_7610,N_5956,N_7291);
nor U7611 (N_7611,N_6590,N_5776);
and U7612 (N_7612,N_5478,N_5809);
nand U7613 (N_7613,N_7099,N_5039);
nor U7614 (N_7614,N_6351,N_5159);
and U7615 (N_7615,N_6918,N_5276);
nor U7616 (N_7616,N_6661,N_5917);
nand U7617 (N_7617,N_5140,N_6491);
xnor U7618 (N_7618,N_6372,N_6127);
nor U7619 (N_7619,N_5955,N_5921);
nand U7620 (N_7620,N_6592,N_5442);
or U7621 (N_7621,N_5714,N_5158);
nand U7622 (N_7622,N_7479,N_5849);
or U7623 (N_7623,N_5831,N_5825);
nand U7624 (N_7624,N_5684,N_7205);
nor U7625 (N_7625,N_6633,N_5535);
nor U7626 (N_7626,N_5174,N_5974);
nand U7627 (N_7627,N_5960,N_7293);
nand U7628 (N_7628,N_5293,N_5472);
and U7629 (N_7629,N_7029,N_7007);
or U7630 (N_7630,N_5092,N_5270);
xor U7631 (N_7631,N_6199,N_7294);
nor U7632 (N_7632,N_6249,N_5551);
nand U7633 (N_7633,N_5812,N_6475);
nor U7634 (N_7634,N_7154,N_6397);
nor U7635 (N_7635,N_5182,N_6412);
and U7636 (N_7636,N_5936,N_6363);
or U7637 (N_7637,N_5047,N_6932);
nor U7638 (N_7638,N_6166,N_6973);
or U7639 (N_7639,N_7100,N_7199);
nor U7640 (N_7640,N_6510,N_7194);
xnor U7641 (N_7641,N_7392,N_5136);
nor U7642 (N_7642,N_5499,N_5765);
or U7643 (N_7643,N_5866,N_7430);
and U7644 (N_7644,N_7424,N_5979);
and U7645 (N_7645,N_6283,N_5169);
or U7646 (N_7646,N_6481,N_6272);
and U7647 (N_7647,N_5547,N_5727);
nand U7648 (N_7648,N_5006,N_5793);
or U7649 (N_7649,N_6649,N_6433);
and U7650 (N_7650,N_5123,N_6483);
or U7651 (N_7651,N_6890,N_7227);
nand U7652 (N_7652,N_5151,N_7079);
nand U7653 (N_7653,N_7476,N_6733);
nand U7654 (N_7654,N_6341,N_6682);
and U7655 (N_7655,N_6728,N_5111);
xnor U7656 (N_7656,N_6844,N_6696);
nor U7657 (N_7657,N_6487,N_6873);
nand U7658 (N_7658,N_7313,N_6097);
nor U7659 (N_7659,N_7000,N_5729);
or U7660 (N_7660,N_6831,N_5640);
and U7661 (N_7661,N_5053,N_5469);
or U7662 (N_7662,N_6614,N_7446);
nand U7663 (N_7663,N_5014,N_6266);
and U7664 (N_7664,N_7193,N_6077);
or U7665 (N_7665,N_7045,N_5787);
nand U7666 (N_7666,N_6336,N_5402);
nand U7667 (N_7667,N_6848,N_5330);
and U7668 (N_7668,N_6092,N_5767);
or U7669 (N_7669,N_7175,N_7139);
or U7670 (N_7670,N_5099,N_5626);
nor U7671 (N_7671,N_6321,N_5707);
and U7672 (N_7672,N_5544,N_7285);
nor U7673 (N_7673,N_5459,N_5200);
and U7674 (N_7674,N_6558,N_6955);
and U7675 (N_7675,N_7006,N_5083);
nor U7676 (N_7676,N_5513,N_6192);
or U7677 (N_7677,N_6259,N_5057);
nor U7678 (N_7678,N_7047,N_5800);
xor U7679 (N_7679,N_6260,N_6282);
xor U7680 (N_7680,N_6484,N_6223);
and U7681 (N_7681,N_7015,N_6920);
and U7682 (N_7682,N_7405,N_6595);
nand U7683 (N_7683,N_6552,N_5923);
nand U7684 (N_7684,N_6744,N_6425);
and U7685 (N_7685,N_5945,N_5060);
nor U7686 (N_7686,N_6385,N_5914);
nor U7687 (N_7687,N_5711,N_7268);
or U7688 (N_7688,N_6786,N_5217);
nor U7689 (N_7689,N_7073,N_6511);
nor U7690 (N_7690,N_5884,N_5346);
nor U7691 (N_7691,N_6401,N_6016);
nand U7692 (N_7692,N_6900,N_6624);
nor U7693 (N_7693,N_6554,N_7140);
nand U7694 (N_7694,N_7487,N_6766);
nand U7695 (N_7695,N_6723,N_6286);
or U7696 (N_7696,N_6985,N_5370);
or U7697 (N_7697,N_5062,N_6325);
and U7698 (N_7698,N_6409,N_6384);
nor U7699 (N_7699,N_5000,N_7363);
nor U7700 (N_7700,N_6956,N_6125);
nand U7701 (N_7701,N_7482,N_6557);
or U7702 (N_7702,N_6037,N_5197);
and U7703 (N_7703,N_6461,N_7148);
nand U7704 (N_7704,N_6340,N_5020);
nand U7705 (N_7705,N_6891,N_6098);
nor U7706 (N_7706,N_5734,N_6431);
and U7707 (N_7707,N_6971,N_5781);
and U7708 (N_7708,N_6364,N_6868);
or U7709 (N_7709,N_6908,N_5387);
or U7710 (N_7710,N_6959,N_7155);
or U7711 (N_7711,N_7125,N_5086);
or U7712 (N_7712,N_5703,N_7027);
or U7713 (N_7713,N_6117,N_6760);
nand U7714 (N_7714,N_7071,N_6027);
or U7715 (N_7715,N_7330,N_6026);
nor U7716 (N_7716,N_6515,N_5692);
xor U7717 (N_7717,N_5995,N_5772);
nand U7718 (N_7718,N_5927,N_7388);
and U7719 (N_7719,N_5242,N_5231);
and U7720 (N_7720,N_5930,N_6085);
nand U7721 (N_7721,N_5113,N_5878);
nor U7722 (N_7722,N_5842,N_7390);
nand U7723 (N_7723,N_7266,N_6583);
and U7724 (N_7724,N_6022,N_7008);
nor U7725 (N_7725,N_6992,N_6417);
and U7726 (N_7726,N_6568,N_5420);
or U7727 (N_7727,N_7447,N_5657);
or U7728 (N_7728,N_6834,N_6088);
nor U7729 (N_7729,N_5161,N_7210);
and U7730 (N_7730,N_6304,N_5746);
and U7731 (N_7731,N_5329,N_6928);
nand U7732 (N_7732,N_6547,N_7342);
or U7733 (N_7733,N_5433,N_6279);
and U7734 (N_7734,N_6619,N_5080);
and U7735 (N_7735,N_6912,N_5430);
or U7736 (N_7736,N_5562,N_6296);
or U7737 (N_7737,N_5491,N_6105);
and U7738 (N_7738,N_5350,N_6563);
or U7739 (N_7739,N_7168,N_5528);
nor U7740 (N_7740,N_6825,N_7201);
nand U7741 (N_7741,N_5802,N_6448);
or U7742 (N_7742,N_7458,N_6710);
nor U7743 (N_7743,N_7108,N_7124);
nor U7744 (N_7744,N_7360,N_7491);
or U7745 (N_7745,N_6792,N_5970);
and U7746 (N_7746,N_6337,N_5646);
nor U7747 (N_7747,N_6242,N_6056);
or U7748 (N_7748,N_6525,N_6013);
and U7749 (N_7749,N_6391,N_5961);
or U7750 (N_7750,N_5994,N_5128);
nor U7751 (N_7751,N_5404,N_5065);
nand U7752 (N_7752,N_5032,N_5620);
nor U7753 (N_7753,N_7009,N_7215);
or U7754 (N_7754,N_5835,N_5973);
nand U7755 (N_7755,N_7457,N_6631);
nor U7756 (N_7756,N_6545,N_5785);
nor U7757 (N_7757,N_7425,N_7223);
nand U7758 (N_7758,N_7032,N_5023);
nand U7759 (N_7759,N_6731,N_5569);
nor U7760 (N_7760,N_5394,N_7080);
nor U7761 (N_7761,N_6311,N_6986);
nand U7762 (N_7762,N_6817,N_6135);
and U7763 (N_7763,N_6870,N_7338);
or U7764 (N_7764,N_5456,N_5419);
nand U7765 (N_7765,N_6808,N_6196);
nand U7766 (N_7766,N_6875,N_6057);
nand U7767 (N_7767,N_6164,N_7429);
and U7768 (N_7768,N_5131,N_6157);
and U7769 (N_7769,N_7260,N_6441);
xor U7770 (N_7770,N_5326,N_5105);
nand U7771 (N_7771,N_5618,N_5063);
nand U7772 (N_7772,N_6291,N_5689);
nand U7773 (N_7773,N_6255,N_5514);
and U7774 (N_7774,N_6496,N_7412);
and U7775 (N_7775,N_6121,N_6726);
or U7776 (N_7776,N_5107,N_7448);
nor U7777 (N_7777,N_6204,N_6280);
nand U7778 (N_7778,N_7063,N_6679);
and U7779 (N_7779,N_5989,N_7061);
xnor U7780 (N_7780,N_6526,N_7287);
or U7781 (N_7781,N_6113,N_6235);
nor U7782 (N_7782,N_5031,N_6686);
nor U7783 (N_7783,N_6241,N_6925);
nor U7784 (N_7784,N_5152,N_7211);
or U7785 (N_7785,N_6087,N_7166);
xnor U7786 (N_7786,N_5333,N_5899);
or U7787 (N_7787,N_7343,N_7132);
and U7788 (N_7788,N_6306,N_5386);
nor U7789 (N_7789,N_5301,N_5347);
or U7790 (N_7790,N_6377,N_6724);
nor U7791 (N_7791,N_6634,N_7145);
nand U7792 (N_7792,N_5325,N_7170);
or U7793 (N_7793,N_6118,N_5500);
and U7794 (N_7794,N_6184,N_5762);
nand U7795 (N_7795,N_5580,N_6025);
nand U7796 (N_7796,N_7209,N_5069);
or U7797 (N_7797,N_6860,N_6793);
nor U7798 (N_7798,N_5221,N_7389);
nor U7799 (N_7799,N_6533,N_6987);
nor U7800 (N_7800,N_6675,N_5134);
nand U7801 (N_7801,N_5311,N_7230);
or U7802 (N_7802,N_6406,N_5611);
and U7803 (N_7803,N_6588,N_6804);
and U7804 (N_7804,N_6323,N_5266);
and U7805 (N_7805,N_7257,N_6339);
nand U7806 (N_7806,N_5991,N_5706);
nor U7807 (N_7807,N_7234,N_6938);
nor U7808 (N_7808,N_5552,N_5972);
and U7809 (N_7809,N_5207,N_5385);
or U7810 (N_7810,N_6083,N_7011);
nand U7811 (N_7811,N_5196,N_5411);
nor U7812 (N_7812,N_7180,N_7279);
nand U7813 (N_7813,N_5808,N_6852);
nand U7814 (N_7814,N_7451,N_6232);
or U7815 (N_7815,N_6247,N_5735);
nor U7816 (N_7816,N_5229,N_6115);
nand U7817 (N_7817,N_5715,N_5794);
nand U7818 (N_7818,N_6376,N_6740);
nand U7819 (N_7819,N_5122,N_5249);
nand U7820 (N_7820,N_5222,N_6958);
and U7821 (N_7821,N_5819,N_5204);
nor U7822 (N_7822,N_6327,N_6522);
or U7823 (N_7823,N_7339,N_5928);
nor U7824 (N_7824,N_5149,N_6898);
or U7825 (N_7825,N_5521,N_5837);
or U7826 (N_7826,N_6416,N_7310);
nor U7827 (N_7827,N_6606,N_5944);
nand U7828 (N_7828,N_5774,N_5892);
nand U7829 (N_7829,N_5250,N_6375);
xnor U7830 (N_7830,N_6318,N_5538);
and U7831 (N_7831,N_7307,N_7200);
or U7832 (N_7832,N_6882,N_5438);
xnor U7833 (N_7833,N_5636,N_6830);
nor U7834 (N_7834,N_5811,N_6556);
or U7835 (N_7835,N_5697,N_6916);
and U7836 (N_7836,N_5591,N_7018);
or U7837 (N_7837,N_5476,N_5348);
nand U7838 (N_7838,N_6435,N_5252);
nor U7839 (N_7839,N_5365,N_5850);
and U7840 (N_7840,N_5596,N_5088);
and U7841 (N_7841,N_7244,N_6152);
or U7842 (N_7842,N_6292,N_6773);
and U7843 (N_7843,N_6671,N_5399);
nor U7844 (N_7844,N_6126,N_6641);
or U7845 (N_7845,N_7466,N_5567);
nor U7846 (N_7846,N_5443,N_6694);
and U7847 (N_7847,N_5473,N_5648);
and U7848 (N_7848,N_5034,N_6456);
or U7849 (N_7849,N_5296,N_6090);
nand U7850 (N_7850,N_6350,N_5671);
or U7851 (N_7851,N_6569,N_6380);
nor U7852 (N_7852,N_5705,N_6331);
xor U7853 (N_7853,N_6840,N_6423);
nor U7854 (N_7854,N_7243,N_6031);
nand U7855 (N_7855,N_6978,N_6869);
or U7856 (N_7856,N_5601,N_7253);
nor U7857 (N_7857,N_7010,N_6393);
nand U7858 (N_7858,N_7024,N_7286);
nor U7859 (N_7859,N_5680,N_6996);
and U7860 (N_7860,N_7303,N_6897);
and U7861 (N_7861,N_5821,N_6131);
nand U7862 (N_7862,N_6460,N_6937);
or U7863 (N_7863,N_6443,N_7102);
and U7864 (N_7864,N_6017,N_6993);
nand U7865 (N_7865,N_7323,N_6173);
nor U7866 (N_7866,N_5823,N_7147);
and U7867 (N_7867,N_7252,N_5467);
or U7868 (N_7868,N_6532,N_5205);
nand U7869 (N_7869,N_5415,N_6449);
or U7870 (N_7870,N_7400,N_6892);
or U7871 (N_7871,N_5699,N_5678);
nand U7872 (N_7872,N_6253,N_6356);
and U7873 (N_7873,N_7115,N_7229);
nor U7874 (N_7874,N_5202,N_6234);
nand U7875 (N_7875,N_5076,N_5949);
nand U7876 (N_7876,N_6240,N_5790);
and U7877 (N_7877,N_6422,N_7426);
xor U7878 (N_7878,N_6219,N_5520);
or U7879 (N_7879,N_7492,N_5510);
nor U7880 (N_7880,N_5931,N_5418);
nand U7881 (N_7881,N_5561,N_5589);
nand U7882 (N_7882,N_5798,N_5957);
nand U7883 (N_7883,N_5924,N_6821);
xor U7884 (N_7884,N_5745,N_6188);
nor U7885 (N_7885,N_5650,N_5303);
or U7886 (N_7886,N_6948,N_7443);
or U7887 (N_7887,N_6594,N_5354);
and U7888 (N_7888,N_7049,N_5397);
or U7889 (N_7889,N_5543,N_6764);
and U7890 (N_7890,N_5488,N_7043);
and U7891 (N_7891,N_5026,N_5210);
nand U7892 (N_7892,N_6389,N_6787);
nor U7893 (N_7893,N_6815,N_7344);
and U7894 (N_7894,N_5361,N_5712);
or U7895 (N_7895,N_7112,N_7397);
nand U7896 (N_7896,N_6370,N_7192);
nand U7897 (N_7897,N_5461,N_6779);
and U7898 (N_7898,N_5982,N_6100);
or U7899 (N_7899,N_5658,N_7273);
nand U7900 (N_7900,N_5030,N_6565);
and U7901 (N_7901,N_5805,N_6153);
or U7902 (N_7902,N_6107,N_5992);
nor U7903 (N_7903,N_6444,N_5104);
nor U7904 (N_7904,N_5452,N_7233);
nand U7905 (N_7905,N_7327,N_7219);
nor U7906 (N_7906,N_6319,N_6645);
nor U7907 (N_7907,N_6975,N_5369);
nand U7908 (N_7908,N_6623,N_6603);
and U7909 (N_7909,N_6745,N_5465);
or U7910 (N_7910,N_7152,N_5933);
nor U7911 (N_7911,N_5911,N_6656);
or U7912 (N_7912,N_5554,N_5693);
and U7913 (N_7913,N_6725,N_5815);
or U7914 (N_7914,N_5389,N_6269);
or U7915 (N_7915,N_6413,N_7305);
nand U7916 (N_7916,N_5838,N_7134);
or U7917 (N_7917,N_6575,N_5133);
or U7918 (N_7918,N_5827,N_5214);
nand U7919 (N_7919,N_7246,N_6539);
and U7920 (N_7920,N_6669,N_5726);
nor U7921 (N_7921,N_5645,N_5356);
nor U7922 (N_7922,N_6564,N_5816);
and U7923 (N_7923,N_5602,N_6353);
nor U7924 (N_7924,N_7144,N_7142);
nor U7925 (N_7925,N_5463,N_7326);
nand U7926 (N_7926,N_5336,N_5292);
nor U7927 (N_7927,N_7022,N_5291);
and U7928 (N_7928,N_7241,N_5959);
or U7929 (N_7929,N_5713,N_7272);
nand U7930 (N_7930,N_5545,N_6347);
and U7931 (N_7931,N_6529,N_7410);
and U7932 (N_7932,N_6111,N_5142);
nand U7933 (N_7933,N_5236,N_5373);
and U7934 (N_7934,N_6867,N_7283);
and U7935 (N_7935,N_6906,N_6775);
and U7936 (N_7936,N_6765,N_5470);
nor U7937 (N_7937,N_5590,N_7003);
nor U7938 (N_7938,N_5144,N_5559);
xnor U7939 (N_7939,N_5977,N_5300);
nor U7940 (N_7940,N_6313,N_5593);
nand U7941 (N_7941,N_7117,N_6951);
and U7942 (N_7942,N_5542,N_5244);
nand U7943 (N_7943,N_6006,N_7316);
nand U7944 (N_7944,N_6776,N_5568);
nand U7945 (N_7945,N_6673,N_5832);
nand U7946 (N_7946,N_6719,N_6806);
nor U7947 (N_7947,N_5858,N_6506);
or U7948 (N_7948,N_5077,N_6239);
nor U7949 (N_7949,N_6683,N_6226);
nand U7950 (N_7950,N_6257,N_5852);
nor U7951 (N_7951,N_7445,N_6795);
xnor U7952 (N_7952,N_5553,N_6655);
and U7953 (N_7953,N_6216,N_5254);
nor U7954 (N_7954,N_5778,N_6687);
nor U7955 (N_7955,N_5135,N_7382);
nor U7956 (N_7956,N_7302,N_6601);
and U7957 (N_7957,N_6957,N_6179);
or U7958 (N_7958,N_6069,N_7196);
and U7959 (N_7959,N_6386,N_5390);
nand U7960 (N_7960,N_7278,N_7331);
and U7961 (N_7961,N_5287,N_6530);
or U7962 (N_7962,N_6877,N_7204);
or U7963 (N_7963,N_6212,N_6156);
nor U7964 (N_7964,N_7036,N_7042);
and U7965 (N_7965,N_5239,N_5530);
nand U7966 (N_7966,N_5127,N_6677);
nor U7967 (N_7967,N_5256,N_6607);
nor U7968 (N_7968,N_5297,N_7058);
and U7969 (N_7969,N_6952,N_5038);
and U7970 (N_7970,N_5922,N_6082);
and U7971 (N_7971,N_6663,N_6812);
nand U7972 (N_7972,N_5890,N_5672);
nand U7973 (N_7973,N_7467,N_6089);
or U7974 (N_7974,N_6368,N_5533);
nor U7975 (N_7975,N_6322,N_6560);
and U7976 (N_7976,N_5382,N_6309);
nand U7977 (N_7977,N_5051,N_5642);
and U7978 (N_7978,N_5529,N_6501);
nand U7979 (N_7979,N_7437,N_6471);
nand U7980 (N_7980,N_6454,N_6822);
or U7981 (N_7981,N_6034,N_6238);
and U7982 (N_7982,N_6243,N_6312);
or U7983 (N_7983,N_6290,N_7357);
or U7984 (N_7984,N_5833,N_6509);
or U7985 (N_7985,N_6281,N_6976);
nand U7986 (N_7986,N_5028,N_5477);
and U7987 (N_7987,N_6301,N_5749);
or U7988 (N_7988,N_5425,N_5938);
or U7989 (N_7989,N_7282,N_6208);
or U7990 (N_7990,N_6797,N_7078);
nand U7991 (N_7991,N_6921,N_7190);
or U7992 (N_7992,N_5784,N_6662);
or U7993 (N_7993,N_6480,N_5964);
nand U7994 (N_7994,N_6478,N_6537);
or U7995 (N_7995,N_5901,N_7114);
nand U7996 (N_7996,N_5600,N_6463);
and U7997 (N_7997,N_7428,N_5584);
and U7998 (N_7998,N_6181,N_5285);
nand U7999 (N_7999,N_6043,N_5147);
nand U8000 (N_8000,N_7432,N_6155);
nor U8001 (N_8001,N_6140,N_5777);
or U8002 (N_8002,N_5265,N_5342);
nor U8003 (N_8003,N_5779,N_6546);
or U8004 (N_8004,N_5082,N_7486);
or U8005 (N_8005,N_5275,N_6803);
nand U8006 (N_8006,N_6730,N_5963);
nand U8007 (N_8007,N_5864,N_6763);
nand U8008 (N_8008,N_6969,N_7376);
nand U8009 (N_8009,N_7475,N_6849);
or U8010 (N_8010,N_5810,N_5457);
and U8011 (N_8011,N_5025,N_6221);
and U8012 (N_8012,N_5048,N_5164);
nor U8013 (N_8013,N_6134,N_5040);
nor U8014 (N_8014,N_7040,N_6360);
or U8015 (N_8015,N_5625,N_5694);
nor U8016 (N_8016,N_6622,N_7055);
nand U8017 (N_8017,N_7419,N_6833);
xnor U8018 (N_8018,N_7026,N_6741);
nand U8019 (N_8019,N_5616,N_5013);
and U8020 (N_8020,N_5985,N_7409);
or U8021 (N_8021,N_7493,N_6109);
nand U8022 (N_8022,N_6383,N_7387);
nand U8023 (N_8023,N_5487,N_5704);
nor U8024 (N_8024,N_5953,N_5246);
and U8025 (N_8025,N_7336,N_5516);
nor U8026 (N_8026,N_5183,N_6613);
nand U8027 (N_8027,N_6917,N_6161);
or U8028 (N_8028,N_7375,N_6344);
or U8029 (N_8029,N_6182,N_6202);
or U8030 (N_8030,N_5983,N_5845);
nor U8031 (N_8031,N_5844,N_7136);
nor U8032 (N_8032,N_6566,N_6538);
nor U8033 (N_8033,N_5950,N_6298);
nor U8034 (N_8034,N_6145,N_6346);
or U8035 (N_8035,N_5067,N_6648);
and U8036 (N_8036,N_5518,N_7121);
and U8037 (N_8037,N_6746,N_7391);
nand U8038 (N_8038,N_6625,N_5733);
or U8039 (N_8039,N_6864,N_6408);
or U8040 (N_8040,N_6095,N_6246);
xor U8041 (N_8041,N_6732,N_6465);
xnor U8042 (N_8042,N_5056,N_5132);
xnor U8043 (N_8043,N_6215,N_6653);
or U8044 (N_8044,N_5255,N_5156);
nor U8045 (N_8045,N_6218,N_7351);
nand U8046 (N_8046,N_5830,N_5525);
nand U8047 (N_8047,N_7133,N_7352);
and U8048 (N_8048,N_5464,N_7090);
nand U8049 (N_8049,N_6584,N_7284);
nand U8050 (N_8050,N_5791,N_5295);
and U8051 (N_8051,N_5124,N_5388);
nor U8052 (N_8052,N_6142,N_6024);
nand U8053 (N_8053,N_5241,N_7356);
nor U8054 (N_8054,N_5540,N_7081);
nor U8055 (N_8055,N_6206,N_6038);
or U8056 (N_8056,N_6637,N_6665);
nand U8057 (N_8057,N_5087,N_7362);
nand U8058 (N_8058,N_5257,N_6843);
nand U8059 (N_8059,N_5458,N_5937);
or U8060 (N_8060,N_5171,N_5138);
nand U8061 (N_8061,N_6264,N_5608);
and U8062 (N_8062,N_7435,N_5359);
nand U8063 (N_8063,N_7012,N_6561);
nand U8064 (N_8064,N_5003,N_5141);
xor U8065 (N_8065,N_5619,N_5226);
and U8066 (N_8066,N_6050,N_5148);
or U8067 (N_8067,N_5380,N_5676);
or U8068 (N_8068,N_7436,N_5903);
and U8069 (N_8069,N_7288,N_6842);
nand U8070 (N_8070,N_7182,N_7245);
nand U8071 (N_8071,N_6195,N_5012);
or U8072 (N_8072,N_6667,N_5916);
nor U8073 (N_8073,N_6981,N_6122);
nand U8074 (N_8074,N_5441,N_5710);
or U8075 (N_8075,N_6357,N_7098);
or U8076 (N_8076,N_7271,N_6738);
nor U8077 (N_8077,N_5515,N_5337);
nor U8078 (N_8078,N_6452,N_5817);
nand U8079 (N_8079,N_5180,N_6778);
or U8080 (N_8080,N_6472,N_6941);
nor U8081 (N_8081,N_6854,N_7417);
nand U8082 (N_8082,N_6418,N_6580);
and U8083 (N_8083,N_5410,N_6358);
nand U8084 (N_8084,N_5796,N_6718);
and U8085 (N_8085,N_5286,N_7146);
and U8086 (N_8086,N_5075,N_6944);
nand U8087 (N_8087,N_6977,N_6837);
nand U8088 (N_8088,N_5125,N_7463);
and U8089 (N_8089,N_6338,N_5717);
or U8090 (N_8090,N_5341,N_7300);
and U8091 (N_8091,N_7251,N_6758);
or U8092 (N_8092,N_6003,N_5050);
xnor U8093 (N_8093,N_6130,N_5137);
or U8094 (N_8094,N_7385,N_6330);
or U8095 (N_8095,N_5688,N_6693);
nand U8096 (N_8096,N_6189,N_5177);
and U8097 (N_8097,N_7014,N_5243);
nand U8098 (N_8098,N_5377,N_7469);
or U8099 (N_8099,N_6964,N_7274);
or U8100 (N_8100,N_7335,N_5971);
nor U8101 (N_8101,N_5245,N_5068);
nand U8102 (N_8102,N_7276,N_6988);
or U8103 (N_8103,N_6602,N_6742);
and U8104 (N_8104,N_6587,N_7420);
and U8105 (N_8105,N_6102,N_5764);
nand U8106 (N_8106,N_7025,N_5358);
nor U8107 (N_8107,N_6536,N_5362);
and U8108 (N_8108,N_5095,N_6520);
nand U8109 (N_8109,N_6593,N_6229);
and U8110 (N_8110,N_5351,N_5259);
nor U8111 (N_8111,N_5637,N_5604);
nand U8112 (N_8112,N_5885,N_6880);
nand U8113 (N_8113,N_7373,N_6691);
nand U8114 (N_8114,N_5851,N_7236);
nor U8115 (N_8115,N_6676,N_6737);
nand U8116 (N_8116,N_6342,N_5033);
nand U8117 (N_8117,N_7384,N_5738);
nand U8118 (N_8118,N_7353,N_6227);
or U8119 (N_8119,N_5999,N_6222);
xor U8120 (N_8120,N_7280,N_5374);
nand U8121 (N_8121,N_5175,N_5423);
nor U8122 (N_8122,N_6473,N_5383);
nand U8123 (N_8123,N_6688,N_6954);
and U8124 (N_8124,N_5268,N_6945);
nand U8125 (N_8125,N_7226,N_5112);
nand U8126 (N_8126,N_6695,N_6252);
nor U8127 (N_8127,N_7046,N_6698);
nor U8128 (N_8128,N_7198,N_5854);
nand U8129 (N_8129,N_5913,N_5681);
and U8130 (N_8130,N_5422,N_6394);
xor U8131 (N_8131,N_5573,N_6681);
nor U8132 (N_8132,N_7143,N_5634);
nor U8133 (N_8133,N_6893,N_6567);
nor U8134 (N_8134,N_6931,N_5632);
or U8135 (N_8135,N_5564,N_5306);
and U8136 (N_8136,N_6838,N_7379);
nor U8137 (N_8137,N_6168,N_6103);
or U8138 (N_8138,N_6850,N_6147);
nor U8139 (N_8139,N_6194,N_6929);
nor U8140 (N_8140,N_5353,N_6500);
and U8141 (N_8141,N_7345,N_6349);
or U8142 (N_8142,N_5453,N_5070);
and U8143 (N_8143,N_6704,N_5857);
or U8144 (N_8144,N_5314,N_5355);
nand U8145 (N_8145,N_7167,N_7481);
nor U8146 (N_8146,N_6180,N_7346);
and U8147 (N_8147,N_5305,N_7095);
or U8148 (N_8148,N_7460,N_6494);
or U8149 (N_8149,N_5185,N_6049);
nor U8150 (N_8150,N_5644,N_6058);
or U8151 (N_8151,N_6129,N_7369);
or U8152 (N_8152,N_7113,N_7450);
nand U8153 (N_8153,N_6398,N_5577);
nor U8154 (N_8154,N_5085,N_5743);
nand U8155 (N_8155,N_5768,N_6664);
nor U8156 (N_8156,N_5879,N_6713);
nand U8157 (N_8157,N_7380,N_6007);
and U8158 (N_8158,N_6611,N_6150);
and U8159 (N_8159,N_7394,N_5829);
nand U8160 (N_8160,N_5228,N_5054);
or U8161 (N_8161,N_7059,N_5001);
and U8162 (N_8162,N_6924,N_5876);
nand U8163 (N_8163,N_7225,N_6599);
xor U8164 (N_8164,N_6374,N_6660);
nor U8165 (N_8165,N_5595,N_5263);
nor U8166 (N_8166,N_7076,N_6984);
nand U8167 (N_8167,N_6263,N_5687);
and U8168 (N_8168,N_5763,N_6966);
nand U8169 (N_8169,N_7401,N_5323);
nor U8170 (N_8170,N_7068,N_6666);
or U8171 (N_8171,N_5489,N_7431);
or U8172 (N_8172,N_5073,N_5381);
nand U8173 (N_8173,N_5818,N_6799);
nand U8174 (N_8174,N_5635,N_7013);
and U8175 (N_8175,N_5496,N_6084);
nand U8176 (N_8176,N_7470,N_6573);
or U8177 (N_8177,N_5670,N_6757);
and U8178 (N_8178,N_5880,N_6450);
nand U8179 (N_8179,N_5624,N_7383);
nor U8180 (N_8180,N_5090,N_7214);
and U8181 (N_8181,N_7333,N_6540);
nand U8182 (N_8182,N_6783,N_6589);
nor U8183 (N_8183,N_7281,N_6748);
nand U8184 (N_8184,N_5507,N_7372);
nand U8185 (N_8185,N_6466,N_6005);
and U8186 (N_8186,N_5371,N_6369);
nor U8187 (N_8187,N_6788,N_6274);
nand U8188 (N_8188,N_7178,N_6236);
and U8189 (N_8189,N_5728,N_7087);
or U8190 (N_8190,N_6523,N_7408);
and U8191 (N_8191,N_5109,N_5783);
and U8192 (N_8192,N_7065,N_6979);
or U8193 (N_8193,N_6571,N_6205);
nor U8194 (N_8194,N_7195,N_7296);
or U8195 (N_8195,N_6160,N_6334);
nor U8196 (N_8196,N_6680,N_6919);
nor U8197 (N_8197,N_6598,N_7407);
nand U8198 (N_8198,N_7277,N_6750);
nand U8199 (N_8199,N_5011,N_5546);
nor U8200 (N_8200,N_6256,N_7089);
nand U8201 (N_8201,N_7122,N_5427);
nand U8202 (N_8202,N_5114,N_7354);
and U8203 (N_8203,N_7398,N_7023);
or U8204 (N_8204,N_7496,N_5523);
nor U8205 (N_8205,N_6387,N_6207);
and U8206 (N_8206,N_5064,N_5641);
and U8207 (N_8207,N_6752,N_6248);
nor U8208 (N_8208,N_5460,N_6670);
nor U8209 (N_8209,N_6642,N_7485);
and U8210 (N_8210,N_5193,N_5824);
and U8211 (N_8211,N_6139,N_5775);
nand U8212 (N_8212,N_7157,N_5902);
and U8213 (N_8213,N_6354,N_7220);
or U8214 (N_8214,N_6998,N_6659);
or U8215 (N_8215,N_6714,N_6857);
or U8216 (N_8216,N_5607,N_5757);
nor U8217 (N_8217,N_5046,N_5571);
nor U8218 (N_8218,N_7378,N_5583);
or U8219 (N_8219,N_6244,N_6712);
nor U8220 (N_8220,N_5509,N_5432);
nor U8221 (N_8221,N_7164,N_5788);
nor U8222 (N_8222,N_5375,N_5725);
nor U8223 (N_8223,N_6621,N_5558);
nor U8224 (N_8224,N_7030,N_6258);
and U8225 (N_8225,N_5215,N_5984);
and U8226 (N_8226,N_6798,N_6579);
and U8227 (N_8227,N_6458,N_7096);
nand U8228 (N_8228,N_5853,N_6032);
nor U8229 (N_8229,N_7107,N_5363);
nor U8230 (N_8230,N_7054,N_6317);
nor U8231 (N_8231,N_6320,N_6447);
or U8232 (N_8232,N_5106,N_5429);
nor U8233 (N_8233,N_5392,N_6415);
nor U8234 (N_8234,N_6582,N_6497);
nor U8235 (N_8235,N_6820,N_7321);
or U8236 (N_8236,N_5406,N_5277);
nand U8237 (N_8237,N_6809,N_7461);
nor U8238 (N_8238,N_6489,N_5614);
and U8239 (N_8239,N_6175,N_6190);
and U8240 (N_8240,N_7159,N_6275);
nor U8241 (N_8241,N_6968,N_5043);
or U8242 (N_8242,N_6046,N_5378);
xor U8243 (N_8243,N_5234,N_5022);
and U8244 (N_8244,N_6172,N_7069);
or U8245 (N_8245,N_5975,N_5586);
nand U8246 (N_8246,N_5908,N_6761);
nor U8247 (N_8247,N_6933,N_7464);
or U8248 (N_8248,N_5436,N_7149);
nand U8249 (N_8249,N_5701,N_6555);
nor U8250 (N_8250,N_6326,N_6112);
nor U8251 (N_8251,N_6294,N_6462);
xnor U8252 (N_8252,N_6805,N_6652);
nor U8253 (N_8253,N_5631,N_6033);
xnor U8254 (N_8254,N_5042,N_6261);
nand U8255 (N_8255,N_7224,N_5360);
nor U8256 (N_8256,N_7355,N_5581);
xnor U8257 (N_8257,N_5615,N_5103);
and U8258 (N_8258,N_7255,N_7249);
nand U8259 (N_8259,N_6054,N_5071);
and U8260 (N_8260,N_5522,N_5588);
nand U8261 (N_8261,N_7365,N_5673);
or U8262 (N_8262,N_6446,N_6440);
nor U8263 (N_8263,N_5167,N_6824);
nand U8264 (N_8264,N_5621,N_6541);
or U8265 (N_8265,N_6562,N_5224);
nand U8266 (N_8266,N_5407,N_6378);
nor U8267 (N_8267,N_5417,N_5279);
nor U8268 (N_8268,N_7176,N_5160);
nand U8269 (N_8269,N_5321,N_6430);
and U8270 (N_8270,N_6884,N_7062);
or U8271 (N_8271,N_5894,N_5344);
and U8272 (N_8272,N_6136,N_5541);
nand U8273 (N_8273,N_5920,N_5505);
nand U8274 (N_8274,N_6591,N_6644);
and U8275 (N_8275,N_7468,N_5609);
and U8276 (N_8276,N_6041,N_6442);
or U8277 (N_8277,N_6635,N_6685);
nand U8278 (N_8278,N_7396,N_6627);
or U8279 (N_8279,N_5267,N_7297);
nor U8280 (N_8280,N_5317,N_7218);
nor U8281 (N_8281,N_5331,N_6527);
or U8282 (N_8282,N_5343,N_5907);
and U8283 (N_8283,N_6609,N_6749);
and U8284 (N_8284,N_5718,N_6295);
nor U8285 (N_8285,N_5652,N_7237);
nand U8286 (N_8286,N_5414,N_6901);
and U8287 (N_8287,N_6544,N_6071);
and U8288 (N_8288,N_6989,N_7358);
nor U8289 (N_8289,N_6650,N_5742);
or U8290 (N_8290,N_6855,N_6388);
and U8291 (N_8291,N_5574,N_6699);
nand U8292 (N_8292,N_5582,N_6549);
nand U8293 (N_8293,N_5570,N_6055);
nor U8294 (N_8294,N_6768,N_5753);
or U8295 (N_8295,N_5594,N_5036);
and U8296 (N_8296,N_6771,N_5312);
or U8297 (N_8297,N_6308,N_6245);
nor U8298 (N_8298,N_6935,N_5661);
nand U8299 (N_8299,N_6894,N_6639);
and U8300 (N_8300,N_6983,N_7074);
or U8301 (N_8301,N_7206,N_5121);
nor U8302 (N_8302,N_6193,N_5685);
or U8303 (N_8303,N_7473,N_5480);
nand U8304 (N_8304,N_5861,N_6052);
nor U8305 (N_8305,N_7440,N_6991);
nand U8306 (N_8306,N_6872,N_5780);
or U8307 (N_8307,N_5988,N_5893);
and U8308 (N_8308,N_6436,N_5435);
or U8309 (N_8309,N_7004,N_5424);
or U8310 (N_8310,N_5059,N_6517);
xor U8311 (N_8311,N_5290,N_7235);
or U8312 (N_8312,N_5501,N_7138);
and U8313 (N_8313,N_5269,N_7270);
nor U8314 (N_8314,N_6233,N_5935);
or U8315 (N_8315,N_5863,N_5340);
nand U8316 (N_8316,N_5663,N_7449);
nand U8317 (N_8317,N_5391,N_6504);
nor U8318 (N_8318,N_7038,N_6020);
nor U8319 (N_8319,N_5926,N_5094);
or U8320 (N_8320,N_5366,N_5803);
and U8321 (N_8321,N_6278,N_5822);
nand U8322 (N_8322,N_5035,N_5690);
nor U8323 (N_8323,N_6094,N_7130);
nand U8324 (N_8324,N_6285,N_7304);
nor U8325 (N_8325,N_6626,N_5942);
nor U8326 (N_8326,N_5281,N_6782);
and U8327 (N_8327,N_5428,N_7371);
nor U8328 (N_8328,N_5723,N_5186);
and U8329 (N_8329,N_6428,N_7320);
or U8330 (N_8330,N_5203,N_5237);
nand U8331 (N_8331,N_6927,N_6332);
or U8332 (N_8332,N_6047,N_6735);
nand U8333 (N_8333,N_5905,N_5934);
and U8334 (N_8334,N_5248,N_6366);
and U8335 (N_8335,N_6469,N_5534);
nor U8336 (N_8336,N_5900,N_5958);
nand U8337 (N_8337,N_5283,N_6705);
or U8338 (N_8338,N_6485,N_5912);
nor U8339 (N_8339,N_6270,N_5444);
or U8340 (N_8340,N_5962,N_7239);
or U8341 (N_8341,N_6287,N_5037);
nand U8342 (N_8342,N_6063,N_7497);
nand U8343 (N_8343,N_6503,N_6000);
nor U8344 (N_8344,N_7423,N_7232);
nand U8345 (N_8345,N_5409,N_6643);
or U8346 (N_8346,N_6514,N_6551);
nor U8347 (N_8347,N_5807,N_5302);
nor U8348 (N_8348,N_6674,N_7341);
nor U8349 (N_8349,N_6297,N_5376);
xnor U8350 (N_8350,N_5997,N_6913);
xor U8351 (N_8351,N_5179,N_7348);
and U8352 (N_8352,N_5004,N_7048);
nor U8353 (N_8353,N_6177,N_6895);
and U8354 (N_8354,N_6672,N_6507);
and U8355 (N_8355,N_6400,N_6072);
and U8356 (N_8356,N_5490,N_7315);
nand U8357 (N_8357,N_7197,N_5143);
nand U8358 (N_8358,N_7261,N_6990);
nand U8359 (N_8359,N_7309,N_5393);
nand U8360 (N_8360,N_7471,N_5462);
nand U8361 (N_8361,N_5058,N_5126);
and U8362 (N_8362,N_6060,N_6213);
nor U8363 (N_8363,N_7083,N_6846);
nor U8364 (N_8364,N_6531,N_6284);
nor U8365 (N_8365,N_5736,N_6859);
or U8366 (N_8366,N_6835,N_6225);
nor U8367 (N_8367,N_5168,N_6729);
and U8368 (N_8368,N_7050,N_6715);
nor U8369 (N_8369,N_7181,N_7311);
nand U8370 (N_8370,N_6615,N_5502);
and U8371 (N_8371,N_5954,N_5005);
or U8372 (N_8372,N_5826,N_6490);
or U8373 (N_8373,N_5550,N_5405);
nand U8374 (N_8374,N_5018,N_5846);
or U8375 (N_8375,N_5744,N_5655);
or U8376 (N_8376,N_5948,N_6254);
nor U8377 (N_8377,N_6600,N_7150);
and U8378 (N_8378,N_6596,N_5682);
nand U8379 (N_8379,N_7203,N_6638);
nand U8380 (N_8380,N_5946,N_5886);
nand U8381 (N_8381,N_7028,N_7444);
nor U8382 (N_8382,N_6014,N_6813);
nor U8383 (N_8383,N_7289,N_7489);
nor U8384 (N_8384,N_5258,N_5117);
nor U8385 (N_8385,N_6210,N_5497);
nor U8386 (N_8386,N_6879,N_5560);
or U8387 (N_8387,N_5882,N_7156);
nor U8388 (N_8388,N_5191,N_6076);
or U8389 (N_8389,N_6116,N_6023);
nand U8390 (N_8390,N_7433,N_6075);
or U8391 (N_8391,N_6011,N_6909);
nand U8392 (N_8392,N_6717,N_6200);
and U8393 (N_8393,N_5862,N_6114);
nor U8394 (N_8394,N_6743,N_6922);
or U8395 (N_8395,N_5508,N_6065);
and U8396 (N_8396,N_5605,N_6646);
or U8397 (N_8397,N_5875,N_6008);
and U8398 (N_8398,N_5235,N_6068);
nand U8399 (N_8399,N_5556,N_5367);
and U8400 (N_8400,N_6474,N_5978);
nor U8401 (N_8401,N_6781,N_6163);
and U8402 (N_8402,N_6802,N_6769);
and U8403 (N_8403,N_7070,N_5756);
or U8404 (N_8404,N_6251,N_5372);
nor U8405 (N_8405,N_6708,N_5494);
and U8406 (N_8406,N_6459,N_6576);
or U8407 (N_8407,N_5966,N_5100);
or U8408 (N_8408,N_6093,N_6889);
nand U8409 (N_8409,N_5773,N_6348);
and U8410 (N_8410,N_6926,N_5218);
xor U8411 (N_8411,N_6419,N_6477);
nand U8412 (N_8412,N_5606,N_7422);
nor U8413 (N_8413,N_5184,N_5115);
and U8414 (N_8414,N_6630,N_6640);
nand U8415 (N_8415,N_7314,N_6162);
nand U8416 (N_8416,N_5598,N_5201);
nor U8417 (N_8417,N_6876,N_6856);
or U8418 (N_8418,N_5548,N_7370);
nor U8419 (N_8419,N_5872,N_7216);
or U8420 (N_8420,N_5002,N_5799);
and U8421 (N_8421,N_5748,N_6519);
or U8422 (N_8422,N_7035,N_6755);
or U8423 (N_8423,N_5526,N_6780);
or U8424 (N_8424,N_6739,N_5338);
and U8425 (N_8425,N_5653,N_5834);
nor U8426 (N_8426,N_6183,N_5078);
or U8427 (N_8427,N_6035,N_7186);
nand U8428 (N_8428,N_7017,N_6209);
or U8429 (N_8429,N_7033,N_6851);
nand U8430 (N_8430,N_7418,N_6464);
and U8431 (N_8431,N_5686,N_5328);
or U8432 (N_8432,N_5698,N_6220);
nor U8433 (N_8433,N_7386,N_6045);
and U8434 (N_8434,N_6574,N_6404);
and U8435 (N_8435,N_6079,N_5482);
xnor U8436 (N_8436,N_6141,N_5952);
nand U8437 (N_8437,N_5130,N_7414);
or U8438 (N_8438,N_5613,N_6521);
nand U8439 (N_8439,N_6654,N_6217);
nand U8440 (N_8440,N_6762,N_6796);
or U8441 (N_8441,N_6482,N_5503);
nand U8442 (N_8442,N_6513,N_6548);
nor U8443 (N_8443,N_5563,N_5868);
nand U8444 (N_8444,N_7077,N_5980);
or U8445 (N_8445,N_5139,N_6885);
or U8446 (N_8446,N_5750,N_5627);
and U8447 (N_8447,N_5450,N_6316);
or U8448 (N_8448,N_5910,N_5549);
nand U8449 (N_8449,N_7207,N_6811);
nor U8450 (N_8450,N_7308,N_5622);
or U8451 (N_8451,N_5664,N_6753);
and U8452 (N_8452,N_5968,N_7060);
and U8453 (N_8453,N_5307,N_6128);
and U8454 (N_8454,N_6365,N_6498);
nand U8455 (N_8455,N_5493,N_6426);
and U8456 (N_8456,N_5055,N_7129);
and U8457 (N_8457,N_7127,N_6438);
or U8458 (N_8458,N_7474,N_7085);
nand U8459 (N_8459,N_5322,N_5181);
or U8460 (N_8460,N_7367,N_7021);
nor U8461 (N_8461,N_6751,N_6457);
or U8462 (N_8462,N_7263,N_5747);
or U8463 (N_8463,N_5909,N_5045);
nor U8464 (N_8464,N_7477,N_7072);
nor U8465 (N_8465,N_6963,N_5264);
nand U8466 (N_8466,N_5446,N_5730);
nor U8467 (N_8467,N_6302,N_6091);
nor U8468 (N_8468,N_5659,N_7306);
nand U8469 (N_8469,N_6994,N_5769);
or U8470 (N_8470,N_6476,N_5384);
or U8471 (N_8471,N_5220,N_6572);
xor U8472 (N_8472,N_7240,N_5702);
and U8473 (N_8473,N_6424,N_7484);
and U8474 (N_8474,N_7067,N_5691);
nor U8475 (N_8475,N_5118,N_6904);
and U8476 (N_8476,N_5101,N_7120);
nor U8477 (N_8477,N_6896,N_6553);
and U8478 (N_8478,N_6455,N_5683);
nor U8479 (N_8479,N_7248,N_6176);
nand U8480 (N_8480,N_5860,N_5566);
nor U8481 (N_8481,N_6828,N_5108);
nand U8482 (N_8482,N_5895,N_6329);
nor U8483 (N_8483,N_7301,N_7104);
nor U8484 (N_8484,N_5700,N_5519);
and U8485 (N_8485,N_6186,N_5599);
and U8486 (N_8486,N_7123,N_6790);
nor U8487 (N_8487,N_7368,N_6352);
and U8488 (N_8488,N_7465,N_6187);
nor U8489 (N_8489,N_6794,N_6692);
nor U8490 (N_8490,N_5969,N_5674);
nor U8491 (N_8491,N_5859,N_5145);
and U8492 (N_8492,N_5294,N_6437);
or U8493 (N_8493,N_5708,N_5786);
nand U8494 (N_8494,N_6800,N_6878);
nor U8495 (N_8495,N_5084,N_6434);
nand U8496 (N_8496,N_6826,N_5150);
or U8497 (N_8497,N_6104,N_7212);
nand U8498 (N_8498,N_6701,N_5639);
nand U8499 (N_8499,N_5771,N_5731);
nand U8500 (N_8500,N_6980,N_5225);
nor U8501 (N_8501,N_5696,N_6396);
nor U8502 (N_8502,N_5170,N_7267);
and U8503 (N_8503,N_6577,N_7238);
nor U8504 (N_8504,N_7322,N_5660);
or U8505 (N_8505,N_6271,N_6262);
or U8506 (N_8506,N_5455,N_6914);
and U8507 (N_8507,N_7082,N_7153);
or U8508 (N_8508,N_7403,N_6486);
or U8509 (N_8509,N_7312,N_5260);
and U8510 (N_8510,N_6405,N_7490);
nand U8511 (N_8511,N_5172,N_7174);
nor U8512 (N_8512,N_6059,N_6265);
nand U8513 (N_8513,N_7421,N_7377);
or U8514 (N_8514,N_5481,N_6706);
or U8515 (N_8515,N_6965,N_6021);
or U8516 (N_8516,N_7173,N_5485);
nor U8517 (N_8517,N_7066,N_6399);
nor U8518 (N_8518,N_5801,N_5758);
nand U8519 (N_8519,N_5888,N_6810);
nand U8520 (N_8520,N_6108,N_7177);
or U8521 (N_8521,N_7317,N_6119);
and U8522 (N_8522,N_6829,N_6324);
nand U8523 (N_8523,N_6159,N_7183);
or U8524 (N_8524,N_7041,N_5585);
and U8525 (N_8525,N_5162,N_6767);
nor U8526 (N_8526,N_7258,N_5284);
nand U8527 (N_8527,N_7413,N_6044);
xor U8528 (N_8528,N_6328,N_6144);
or U8529 (N_8529,N_7091,N_5941);
and U8530 (N_8530,N_7075,N_6512);
nand U8531 (N_8531,N_5213,N_5873);
nand U8532 (N_8532,N_6982,N_5178);
nor U8533 (N_8533,N_6862,N_5316);
or U8534 (N_8534,N_5755,N_7161);
or U8535 (N_8535,N_5029,N_7231);
or U8536 (N_8536,N_6178,N_6709);
and U8537 (N_8537,N_5932,N_6736);
nor U8538 (N_8538,N_5766,N_6947);
and U8539 (N_8539,N_5019,N_6086);
and U8540 (N_8540,N_5719,N_7366);
and U8541 (N_8541,N_5947,N_6657);
and U8542 (N_8542,N_7001,N_6231);
nor U8543 (N_8543,N_5536,N_6902);
or U8544 (N_8544,N_5049,N_6858);
nand U8545 (N_8545,N_6070,N_6581);
and U8546 (N_8546,N_5466,N_6940);
or U8547 (N_8547,N_6214,N_5021);
nand U8548 (N_8548,N_5915,N_6064);
nor U8549 (N_8549,N_7292,N_7269);
or U8550 (N_8550,N_7350,N_6910);
and U8551 (N_8551,N_6169,N_6081);
and U8552 (N_8552,N_6702,N_7221);
nand U8553 (N_8553,N_5720,N_5282);
nor U8554 (N_8554,N_7101,N_7084);
nor U8555 (N_8555,N_7328,N_5227);
nand U8556 (N_8556,N_5010,N_7034);
and U8557 (N_8557,N_5334,N_6203);
or U8558 (N_8558,N_7118,N_5806);
or U8559 (N_8559,N_7454,N_5009);
or U8560 (N_8560,N_7228,N_5760);
and U8561 (N_8561,N_6410,N_5841);
nand U8562 (N_8562,N_6930,N_5412);
or U8563 (N_8563,N_5840,N_7160);
nand U8564 (N_8564,N_5223,N_5887);
nand U8565 (N_8565,N_7298,N_6974);
nor U8566 (N_8566,N_6936,N_6550);
nand U8567 (N_8567,N_6467,N_6943);
and U8568 (N_8568,N_5052,N_6716);
nor U8569 (N_8569,N_6586,N_5814);
nand U8570 (N_8570,N_5732,N_5091);
nor U8571 (N_8571,N_6061,N_6333);
or U8572 (N_8572,N_5669,N_5531);
and U8573 (N_8573,N_5940,N_6493);
nand U8574 (N_8574,N_5668,N_5575);
nor U8575 (N_8575,N_7340,N_5110);
and U8576 (N_8576,N_6727,N_7459);
nor U8577 (N_8577,N_7456,N_6785);
nand U8578 (N_8578,N_5318,N_5603);
or U8579 (N_8579,N_5289,N_5504);
nor U8580 (N_8580,N_5537,N_6310);
and U8581 (N_8581,N_5555,N_5870);
or U8582 (N_8582,N_7299,N_7319);
or U8583 (N_8583,N_5471,N_5273);
or U8584 (N_8584,N_5324,N_6167);
nand U8585 (N_8585,N_7256,N_7039);
nor U8586 (N_8586,N_5628,N_5400);
nor U8587 (N_8587,N_5015,N_7188);
nor U8588 (N_8588,N_7442,N_7483);
nor U8589 (N_8589,N_5925,N_5262);
and U8590 (N_8590,N_5709,N_7097);
or U8591 (N_8591,N_6395,N_5883);
nand U8592 (N_8592,N_5527,N_5274);
and U8593 (N_8593,N_5610,N_5484);
nor U8594 (N_8594,N_5662,N_6678);
or U8595 (N_8595,N_5439,N_7213);
nor U8596 (N_8596,N_6029,N_7374);
nand U8597 (N_8597,N_6165,N_5677);
and U8598 (N_8598,N_6479,N_6939);
or U8599 (N_8599,N_6001,N_7056);
or U8600 (N_8600,N_6429,N_6470);
or U8601 (N_8601,N_6632,N_5578);
and U8602 (N_8602,N_5176,N_5532);
nor U8603 (N_8603,N_6028,N_6845);
and U8604 (N_8604,N_7250,N_5403);
and U8605 (N_8605,N_7325,N_5741);
nand U8606 (N_8606,N_5309,N_5592);
nor U8607 (N_8607,N_6754,N_6373);
or U8608 (N_8608,N_5724,N_5990);
nor U8609 (N_8609,N_5675,N_5740);
or U8610 (N_8610,N_6827,N_6468);
nor U8611 (N_8611,N_6305,N_5066);
and U8612 (N_8612,N_5492,N_5874);
xnor U8613 (N_8613,N_7016,N_6807);
nand U8614 (N_8614,N_6759,N_6228);
nor U8615 (N_8615,N_5233,N_6133);
nand U8616 (N_8616,N_6185,N_5792);
or U8617 (N_8617,N_6524,N_5651);
or U8618 (N_8618,N_5918,N_6106);
or U8619 (N_8619,N_5643,N_5721);
nand U8620 (N_8620,N_6314,N_5804);
or U8621 (N_8621,N_5194,N_6359);
and U8622 (N_8622,N_7264,N_6390);
and U8623 (N_8623,N_5666,N_6970);
nor U8624 (N_8624,N_5820,N_5475);
nand U8625 (N_8625,N_5511,N_5981);
nand U8626 (N_8626,N_6628,N_6495);
and U8627 (N_8627,N_6903,N_5524);
nor U8628 (N_8628,N_6138,N_7005);
and U8629 (N_8629,N_6814,N_5304);
or U8630 (N_8630,N_5517,N_6042);
and U8631 (N_8631,N_6439,N_5163);
or U8632 (N_8632,N_5319,N_6997);
nand U8633 (N_8633,N_6508,N_6658);
nor U8634 (N_8634,N_6905,N_5943);
nand U8635 (N_8635,N_6355,N_5313);
and U8636 (N_8636,N_5647,N_6707);
and U8637 (N_8637,N_5008,N_6942);
nand U8638 (N_8638,N_5630,N_7116);
and U8639 (N_8639,N_7452,N_6907);
nor U8640 (N_8640,N_6039,N_5093);
nand U8641 (N_8641,N_6198,N_7051);
and U8642 (N_8642,N_6230,N_6078);
and U8643 (N_8643,N_5335,N_6888);
nor U8644 (N_8644,N_5512,N_7208);
nand U8645 (N_8645,N_7141,N_5633);
nor U8646 (N_8646,N_5896,N_5395);
and U8647 (N_8647,N_6293,N_6148);
nand U8648 (N_8648,N_6585,N_5629);
or U8649 (N_8649,N_7361,N_6923);
and U8650 (N_8650,N_5173,N_5157);
and U8651 (N_8651,N_6137,N_5848);
nor U8652 (N_8652,N_5120,N_5871);
nor U8653 (N_8653,N_5413,N_5079);
nand U8654 (N_8654,N_5993,N_5847);
or U8655 (N_8655,N_6420,N_5498);
xnor U8656 (N_8656,N_6953,N_6451);
nor U8657 (N_8657,N_6899,N_7441);
and U8658 (N_8658,N_5044,N_5906);
nand U8659 (N_8659,N_7151,N_7472);
nor U8660 (N_8660,N_7189,N_5987);
or U8661 (N_8661,N_6960,N_6099);
and U8662 (N_8662,N_6315,N_6191);
nand U8663 (N_8663,N_7393,N_6379);
and U8664 (N_8664,N_5828,N_7498);
and U8665 (N_8665,N_7020,N_5612);
nor U8666 (N_8666,N_5368,N_6722);
nor U8667 (N_8667,N_6711,N_5154);
and U8668 (N_8668,N_7163,N_7126);
nand U8669 (N_8669,N_5904,N_6874);
or U8670 (N_8670,N_6080,N_7332);
nand U8671 (N_8671,N_7131,N_5951);
nand U8672 (N_8672,N_5416,N_6015);
or U8673 (N_8673,N_6110,N_5216);
xor U8674 (N_8674,N_7381,N_6268);
or U8675 (N_8675,N_7265,N_5617);
nor U8676 (N_8676,N_6967,N_6772);
and U8677 (N_8677,N_5272,N_5919);
and U8678 (N_8678,N_6030,N_5016);
and U8679 (N_8679,N_5898,N_5195);
or U8680 (N_8680,N_5855,N_5656);
or U8681 (N_8681,N_7137,N_5357);
nand U8682 (N_8682,N_7105,N_6053);
or U8683 (N_8683,N_6036,N_6074);
nor U8684 (N_8684,N_6048,N_6605);
nand U8685 (N_8685,N_5119,N_6453);
or U8686 (N_8686,N_7404,N_6946);
or U8687 (N_8687,N_5396,N_5867);
or U8688 (N_8688,N_6299,N_6516);
nand U8689 (N_8689,N_5209,N_6668);
nand U8690 (N_8690,N_6816,N_6062);
or U8691 (N_8691,N_6915,N_5278);
and U8692 (N_8692,N_5565,N_6999);
nor U8693 (N_8693,N_5253,N_5967);
nand U8694 (N_8694,N_5889,N_5230);
nor U8695 (N_8695,N_6307,N_6836);
and U8696 (N_8696,N_7434,N_5206);
xnor U8697 (N_8697,N_6502,N_6371);
and U8698 (N_8698,N_5869,N_5153);
or U8699 (N_8699,N_5998,N_7222);
or U8700 (N_8700,N_6629,N_5440);
or U8701 (N_8701,N_6123,N_6684);
or U8702 (N_8702,N_5401,N_6689);
nor U8703 (N_8703,N_6770,N_6124);
and U8704 (N_8704,N_5187,N_6335);
nand U8705 (N_8705,N_7259,N_6492);
nor U8706 (N_8706,N_6040,N_6158);
nand U8707 (N_8707,N_6784,N_5587);
or U8708 (N_8708,N_6250,N_6154);
and U8709 (N_8709,N_7254,N_5232);
and U8710 (N_8710,N_6620,N_7103);
or U8711 (N_8711,N_7064,N_6950);
nand U8712 (N_8712,N_6197,N_7111);
and U8713 (N_8713,N_5722,N_6499);
nand U8714 (N_8714,N_5155,N_5098);
and U8715 (N_8715,N_6171,N_7217);
nand U8716 (N_8716,N_6174,N_6224);
nand U8717 (N_8717,N_7052,N_5097);
or U8718 (N_8718,N_5737,N_7135);
nand U8719 (N_8719,N_5024,N_5007);
and U8720 (N_8720,N_5495,N_5364);
or U8721 (N_8721,N_7031,N_5654);
nor U8722 (N_8722,N_6421,N_5506);
nor U8723 (N_8723,N_5434,N_5081);
or U8724 (N_8724,N_6886,N_5929);
nor U8725 (N_8725,N_7395,N_5327);
or U8726 (N_8726,N_6597,N_6789);
and U8727 (N_8727,N_7462,N_6861);
nand U8728 (N_8728,N_6009,N_5752);
nand U8729 (N_8729,N_6612,N_7169);
or U8730 (N_8730,N_5116,N_7162);
nand U8731 (N_8731,N_6402,N_7185);
nand U8732 (N_8732,N_6818,N_5298);
and U8733 (N_8733,N_7092,N_6143);
nor U8734 (N_8734,N_6690,N_5089);
nor U8735 (N_8735,N_5261,N_6734);
and U8736 (N_8736,N_6871,N_6367);
nor U8737 (N_8737,N_6774,N_5986);
nor U8738 (N_8738,N_5761,N_7057);
nand U8739 (N_8739,N_7044,N_5332);
and U8740 (N_8740,N_5789,N_7406);
and U8741 (N_8741,N_5649,N_6747);
nor U8742 (N_8742,N_6012,N_6004);
or U8743 (N_8743,N_5165,N_5865);
and U8744 (N_8744,N_5445,N_7478);
xor U8745 (N_8745,N_7359,N_5280);
and U8746 (N_8746,N_6132,N_7499);
or U8747 (N_8747,N_6700,N_5474);
or U8748 (N_8748,N_6756,N_7334);
nor U8749 (N_8749,N_6120,N_6697);
nand U8750 (N_8750,N_5168,N_6366);
nand U8751 (N_8751,N_6025,N_6241);
or U8752 (N_8752,N_6568,N_5879);
nand U8753 (N_8753,N_5333,N_5759);
nor U8754 (N_8754,N_5619,N_5304);
or U8755 (N_8755,N_7051,N_6977);
or U8756 (N_8756,N_6508,N_5292);
or U8757 (N_8757,N_7052,N_5507);
nor U8758 (N_8758,N_6122,N_7066);
nor U8759 (N_8759,N_6593,N_7447);
or U8760 (N_8760,N_6629,N_6051);
or U8761 (N_8761,N_5075,N_5666);
nor U8762 (N_8762,N_5302,N_5484);
or U8763 (N_8763,N_7147,N_7372);
nand U8764 (N_8764,N_6510,N_5902);
nor U8765 (N_8765,N_5807,N_6240);
nor U8766 (N_8766,N_6391,N_6688);
and U8767 (N_8767,N_6115,N_7011);
nor U8768 (N_8768,N_5930,N_5066);
or U8769 (N_8769,N_5700,N_7280);
nor U8770 (N_8770,N_5600,N_7075);
or U8771 (N_8771,N_6359,N_6377);
and U8772 (N_8772,N_5617,N_7118);
nor U8773 (N_8773,N_7039,N_7483);
nand U8774 (N_8774,N_5981,N_6405);
and U8775 (N_8775,N_5963,N_5724);
nor U8776 (N_8776,N_6972,N_7105);
or U8777 (N_8777,N_5437,N_6120);
and U8778 (N_8778,N_5743,N_5511);
nand U8779 (N_8779,N_5471,N_6842);
nand U8780 (N_8780,N_5384,N_5934);
and U8781 (N_8781,N_5482,N_6643);
nor U8782 (N_8782,N_6053,N_7212);
or U8783 (N_8783,N_6111,N_7041);
xnor U8784 (N_8784,N_6623,N_6635);
and U8785 (N_8785,N_5533,N_5576);
and U8786 (N_8786,N_5542,N_6279);
nor U8787 (N_8787,N_5875,N_7277);
nor U8788 (N_8788,N_5535,N_6698);
and U8789 (N_8789,N_5403,N_5073);
nor U8790 (N_8790,N_5343,N_7369);
nand U8791 (N_8791,N_7046,N_7319);
nor U8792 (N_8792,N_5074,N_5252);
and U8793 (N_8793,N_6697,N_6872);
xor U8794 (N_8794,N_5070,N_7039);
nand U8795 (N_8795,N_6133,N_7024);
nand U8796 (N_8796,N_6292,N_5663);
or U8797 (N_8797,N_7142,N_5913);
and U8798 (N_8798,N_5863,N_5843);
and U8799 (N_8799,N_6221,N_5876);
nor U8800 (N_8800,N_7143,N_6689);
nand U8801 (N_8801,N_7392,N_7187);
nand U8802 (N_8802,N_7276,N_5911);
nand U8803 (N_8803,N_6728,N_5657);
and U8804 (N_8804,N_7162,N_5700);
or U8805 (N_8805,N_6293,N_5070);
or U8806 (N_8806,N_7012,N_5733);
nor U8807 (N_8807,N_5103,N_5800);
or U8808 (N_8808,N_5805,N_7251);
or U8809 (N_8809,N_6085,N_5622);
nor U8810 (N_8810,N_6181,N_5119);
xor U8811 (N_8811,N_5136,N_6430);
nand U8812 (N_8812,N_7270,N_6393);
and U8813 (N_8813,N_6357,N_6342);
nor U8814 (N_8814,N_7217,N_6954);
nor U8815 (N_8815,N_6269,N_6477);
nand U8816 (N_8816,N_6814,N_6864);
nand U8817 (N_8817,N_5506,N_7413);
or U8818 (N_8818,N_7076,N_6496);
or U8819 (N_8819,N_5236,N_7352);
nand U8820 (N_8820,N_5643,N_6157);
or U8821 (N_8821,N_6543,N_6259);
nand U8822 (N_8822,N_5667,N_5114);
nor U8823 (N_8823,N_5039,N_6694);
and U8824 (N_8824,N_5242,N_6313);
or U8825 (N_8825,N_6540,N_7475);
nor U8826 (N_8826,N_5054,N_6593);
and U8827 (N_8827,N_6551,N_5928);
nand U8828 (N_8828,N_6069,N_5097);
xor U8829 (N_8829,N_6786,N_6138);
nor U8830 (N_8830,N_6049,N_6423);
nor U8831 (N_8831,N_6995,N_5137);
and U8832 (N_8832,N_7115,N_5443);
nand U8833 (N_8833,N_7346,N_7260);
nand U8834 (N_8834,N_7449,N_5734);
nor U8835 (N_8835,N_6081,N_7480);
nand U8836 (N_8836,N_5079,N_5792);
and U8837 (N_8837,N_7431,N_6015);
nor U8838 (N_8838,N_6042,N_5253);
or U8839 (N_8839,N_5309,N_5974);
nand U8840 (N_8840,N_5233,N_7286);
nand U8841 (N_8841,N_6075,N_7412);
and U8842 (N_8842,N_6785,N_5506);
and U8843 (N_8843,N_6482,N_6969);
or U8844 (N_8844,N_6434,N_5053);
nor U8845 (N_8845,N_5826,N_6202);
or U8846 (N_8846,N_6022,N_6368);
nand U8847 (N_8847,N_6329,N_7197);
nand U8848 (N_8848,N_7044,N_5845);
and U8849 (N_8849,N_6636,N_5026);
nand U8850 (N_8850,N_7489,N_5909);
xnor U8851 (N_8851,N_5505,N_6318);
and U8852 (N_8852,N_6160,N_6641);
nor U8853 (N_8853,N_6901,N_7430);
nor U8854 (N_8854,N_6776,N_5348);
nand U8855 (N_8855,N_7486,N_6707);
or U8856 (N_8856,N_5367,N_5571);
nand U8857 (N_8857,N_5715,N_6623);
and U8858 (N_8858,N_6828,N_6647);
nor U8859 (N_8859,N_5317,N_6505);
or U8860 (N_8860,N_5784,N_6332);
and U8861 (N_8861,N_7249,N_6032);
and U8862 (N_8862,N_7222,N_5355);
or U8863 (N_8863,N_7042,N_5508);
nor U8864 (N_8864,N_7154,N_5463);
nor U8865 (N_8865,N_6906,N_7420);
nor U8866 (N_8866,N_6150,N_5774);
and U8867 (N_8867,N_7257,N_7184);
and U8868 (N_8868,N_5786,N_7005);
nor U8869 (N_8869,N_6015,N_5492);
nor U8870 (N_8870,N_6822,N_5067);
nor U8871 (N_8871,N_6999,N_6844);
nand U8872 (N_8872,N_5008,N_5608);
nor U8873 (N_8873,N_5902,N_7016);
nor U8874 (N_8874,N_6664,N_7150);
nor U8875 (N_8875,N_6531,N_5164);
and U8876 (N_8876,N_5308,N_5154);
nor U8877 (N_8877,N_5647,N_5056);
nor U8878 (N_8878,N_5834,N_7398);
and U8879 (N_8879,N_5218,N_6395);
nand U8880 (N_8880,N_6755,N_5969);
nand U8881 (N_8881,N_6590,N_5201);
nor U8882 (N_8882,N_6528,N_6396);
nor U8883 (N_8883,N_7061,N_5835);
and U8884 (N_8884,N_6163,N_5843);
nor U8885 (N_8885,N_5743,N_7255);
nand U8886 (N_8886,N_5871,N_7348);
nor U8887 (N_8887,N_6340,N_7418);
nand U8888 (N_8888,N_5326,N_5729);
nor U8889 (N_8889,N_7312,N_7232);
or U8890 (N_8890,N_5247,N_6207);
and U8891 (N_8891,N_7172,N_6940);
nor U8892 (N_8892,N_7391,N_7449);
nand U8893 (N_8893,N_6382,N_5177);
or U8894 (N_8894,N_5243,N_6156);
nand U8895 (N_8895,N_7054,N_7022);
nand U8896 (N_8896,N_5351,N_5938);
and U8897 (N_8897,N_5318,N_7124);
nor U8898 (N_8898,N_6318,N_7213);
and U8899 (N_8899,N_7326,N_6794);
or U8900 (N_8900,N_6019,N_7111);
or U8901 (N_8901,N_6500,N_5972);
and U8902 (N_8902,N_7393,N_6444);
or U8903 (N_8903,N_7114,N_5577);
or U8904 (N_8904,N_7224,N_7482);
nand U8905 (N_8905,N_5094,N_7037);
nand U8906 (N_8906,N_6817,N_6062);
or U8907 (N_8907,N_6677,N_5693);
and U8908 (N_8908,N_6762,N_7119);
nand U8909 (N_8909,N_5029,N_5230);
nand U8910 (N_8910,N_5724,N_7414);
xnor U8911 (N_8911,N_5830,N_5090);
nand U8912 (N_8912,N_6699,N_7205);
nand U8913 (N_8913,N_6196,N_6835);
xor U8914 (N_8914,N_6007,N_6896);
and U8915 (N_8915,N_5421,N_5251);
nand U8916 (N_8916,N_5861,N_7434);
nand U8917 (N_8917,N_5388,N_6042);
nor U8918 (N_8918,N_6543,N_6444);
nor U8919 (N_8919,N_5393,N_6926);
nand U8920 (N_8920,N_7086,N_5864);
nand U8921 (N_8921,N_6555,N_6223);
or U8922 (N_8922,N_5917,N_6084);
xor U8923 (N_8923,N_6985,N_6942);
nand U8924 (N_8924,N_5423,N_6022);
nand U8925 (N_8925,N_6086,N_7357);
nor U8926 (N_8926,N_6704,N_6049);
nand U8927 (N_8927,N_6899,N_7050);
nor U8928 (N_8928,N_7478,N_7038);
or U8929 (N_8929,N_5231,N_6281);
nand U8930 (N_8930,N_7083,N_5733);
and U8931 (N_8931,N_7454,N_5742);
nor U8932 (N_8932,N_5258,N_6580);
nand U8933 (N_8933,N_7122,N_5789);
nand U8934 (N_8934,N_6970,N_5310);
nor U8935 (N_8935,N_7094,N_6924);
or U8936 (N_8936,N_5763,N_7459);
nand U8937 (N_8937,N_5444,N_6314);
and U8938 (N_8938,N_6697,N_6827);
and U8939 (N_8939,N_6994,N_6257);
and U8940 (N_8940,N_6133,N_6350);
and U8941 (N_8941,N_7194,N_6041);
or U8942 (N_8942,N_5590,N_5042);
nor U8943 (N_8943,N_5699,N_5471);
nand U8944 (N_8944,N_6688,N_6547);
nor U8945 (N_8945,N_6313,N_6440);
nor U8946 (N_8946,N_6656,N_5563);
nor U8947 (N_8947,N_7018,N_7259);
and U8948 (N_8948,N_6285,N_6976);
nand U8949 (N_8949,N_6813,N_5434);
or U8950 (N_8950,N_6009,N_7124);
and U8951 (N_8951,N_6529,N_6628);
nand U8952 (N_8952,N_7027,N_5482);
and U8953 (N_8953,N_5181,N_6380);
and U8954 (N_8954,N_6227,N_5702);
nand U8955 (N_8955,N_7394,N_6570);
nor U8956 (N_8956,N_6410,N_7078);
and U8957 (N_8957,N_7048,N_5153);
nand U8958 (N_8958,N_7091,N_5384);
nor U8959 (N_8959,N_6454,N_7186);
or U8960 (N_8960,N_6201,N_6035);
and U8961 (N_8961,N_7329,N_5991);
nand U8962 (N_8962,N_5752,N_5187);
or U8963 (N_8963,N_7134,N_6271);
nand U8964 (N_8964,N_7232,N_6721);
nor U8965 (N_8965,N_7388,N_5804);
or U8966 (N_8966,N_5363,N_6266);
nor U8967 (N_8967,N_7493,N_5662);
nand U8968 (N_8968,N_5062,N_6613);
or U8969 (N_8969,N_6619,N_6587);
and U8970 (N_8970,N_7270,N_7126);
nand U8971 (N_8971,N_7224,N_6171);
nor U8972 (N_8972,N_5338,N_7077);
nor U8973 (N_8973,N_5500,N_6925);
and U8974 (N_8974,N_5006,N_5990);
nor U8975 (N_8975,N_6467,N_5632);
and U8976 (N_8976,N_5569,N_7298);
or U8977 (N_8977,N_5156,N_6609);
nand U8978 (N_8978,N_7297,N_6404);
and U8979 (N_8979,N_7103,N_5081);
nand U8980 (N_8980,N_6015,N_6917);
nand U8981 (N_8981,N_5529,N_5117);
or U8982 (N_8982,N_5269,N_5330);
nand U8983 (N_8983,N_6191,N_6304);
or U8984 (N_8984,N_5222,N_6048);
and U8985 (N_8985,N_7086,N_5301);
nor U8986 (N_8986,N_5184,N_6992);
nand U8987 (N_8987,N_5701,N_5973);
or U8988 (N_8988,N_5040,N_6977);
nor U8989 (N_8989,N_5824,N_6460);
nand U8990 (N_8990,N_5389,N_6968);
nand U8991 (N_8991,N_5285,N_5683);
nor U8992 (N_8992,N_6826,N_7463);
nor U8993 (N_8993,N_5031,N_6546);
or U8994 (N_8994,N_7392,N_6296);
nor U8995 (N_8995,N_6776,N_6227);
nor U8996 (N_8996,N_6292,N_7065);
or U8997 (N_8997,N_5363,N_5189);
and U8998 (N_8998,N_6996,N_5062);
or U8999 (N_8999,N_5405,N_5400);
nor U9000 (N_9000,N_6197,N_5732);
or U9001 (N_9001,N_5050,N_6387);
or U9002 (N_9002,N_6706,N_6308);
and U9003 (N_9003,N_5978,N_6640);
or U9004 (N_9004,N_5844,N_6425);
and U9005 (N_9005,N_7307,N_5450);
nand U9006 (N_9006,N_7388,N_5319);
or U9007 (N_9007,N_5971,N_6290);
and U9008 (N_9008,N_5884,N_5415);
nand U9009 (N_9009,N_5124,N_6532);
and U9010 (N_9010,N_6639,N_6570);
nor U9011 (N_9011,N_6568,N_7196);
nand U9012 (N_9012,N_7270,N_6951);
nor U9013 (N_9013,N_5696,N_7070);
and U9014 (N_9014,N_6708,N_5464);
or U9015 (N_9015,N_5845,N_7326);
nand U9016 (N_9016,N_6820,N_6007);
nor U9017 (N_9017,N_5818,N_7273);
and U9018 (N_9018,N_6834,N_7257);
or U9019 (N_9019,N_6439,N_7179);
nand U9020 (N_9020,N_6125,N_6193);
and U9021 (N_9021,N_5474,N_6621);
and U9022 (N_9022,N_5600,N_5496);
and U9023 (N_9023,N_5200,N_7136);
nor U9024 (N_9024,N_6604,N_5481);
nand U9025 (N_9025,N_6549,N_6736);
nand U9026 (N_9026,N_6758,N_5558);
nand U9027 (N_9027,N_6375,N_7230);
and U9028 (N_9028,N_6071,N_5631);
nand U9029 (N_9029,N_7235,N_5939);
xnor U9030 (N_9030,N_6538,N_7235);
or U9031 (N_9031,N_5415,N_6138);
nand U9032 (N_9032,N_5226,N_5119);
nor U9033 (N_9033,N_5639,N_5277);
nand U9034 (N_9034,N_5990,N_6142);
nor U9035 (N_9035,N_7291,N_6956);
or U9036 (N_9036,N_6138,N_6845);
nand U9037 (N_9037,N_7115,N_6586);
nand U9038 (N_9038,N_6616,N_6543);
or U9039 (N_9039,N_6970,N_6801);
and U9040 (N_9040,N_6711,N_5514);
and U9041 (N_9041,N_5564,N_6731);
nand U9042 (N_9042,N_5098,N_6099);
nor U9043 (N_9043,N_7489,N_6182);
and U9044 (N_9044,N_5243,N_7198);
or U9045 (N_9045,N_5396,N_7363);
or U9046 (N_9046,N_7031,N_7444);
and U9047 (N_9047,N_7251,N_6808);
xor U9048 (N_9048,N_6645,N_6562);
nand U9049 (N_9049,N_6315,N_5782);
nand U9050 (N_9050,N_6946,N_6220);
nand U9051 (N_9051,N_6451,N_6470);
or U9052 (N_9052,N_6883,N_5198);
nand U9053 (N_9053,N_6662,N_7191);
or U9054 (N_9054,N_7198,N_5109);
nand U9055 (N_9055,N_5547,N_7066);
or U9056 (N_9056,N_5753,N_7429);
nand U9057 (N_9057,N_5202,N_5727);
nor U9058 (N_9058,N_6160,N_5482);
or U9059 (N_9059,N_6992,N_6374);
nand U9060 (N_9060,N_5898,N_6463);
nand U9061 (N_9061,N_5644,N_5478);
nand U9062 (N_9062,N_5801,N_6217);
or U9063 (N_9063,N_7430,N_7312);
nand U9064 (N_9064,N_5925,N_6749);
and U9065 (N_9065,N_7264,N_6775);
nand U9066 (N_9066,N_6003,N_7258);
nand U9067 (N_9067,N_7136,N_5751);
or U9068 (N_9068,N_7362,N_6740);
and U9069 (N_9069,N_6831,N_5900);
nor U9070 (N_9070,N_5876,N_7459);
nor U9071 (N_9071,N_6793,N_6062);
or U9072 (N_9072,N_6315,N_5427);
or U9073 (N_9073,N_6810,N_6665);
and U9074 (N_9074,N_5653,N_6014);
nand U9075 (N_9075,N_6615,N_5615);
nor U9076 (N_9076,N_5715,N_5421);
or U9077 (N_9077,N_5412,N_5183);
or U9078 (N_9078,N_6750,N_5926);
or U9079 (N_9079,N_6060,N_7265);
nand U9080 (N_9080,N_6007,N_6890);
or U9081 (N_9081,N_6376,N_5276);
and U9082 (N_9082,N_6126,N_5009);
nand U9083 (N_9083,N_5712,N_5215);
nand U9084 (N_9084,N_6988,N_7321);
nand U9085 (N_9085,N_7218,N_7187);
or U9086 (N_9086,N_6561,N_7206);
or U9087 (N_9087,N_5141,N_5881);
and U9088 (N_9088,N_5013,N_7144);
and U9089 (N_9089,N_6723,N_5240);
nor U9090 (N_9090,N_5593,N_5883);
or U9091 (N_9091,N_6535,N_5504);
nand U9092 (N_9092,N_5684,N_6736);
and U9093 (N_9093,N_5434,N_6977);
and U9094 (N_9094,N_7168,N_5880);
nor U9095 (N_9095,N_6855,N_7221);
nor U9096 (N_9096,N_5268,N_5534);
nand U9097 (N_9097,N_6794,N_6080);
nor U9098 (N_9098,N_6582,N_7081);
nand U9099 (N_9099,N_5136,N_6557);
nand U9100 (N_9100,N_5137,N_6979);
nor U9101 (N_9101,N_5790,N_5777);
nand U9102 (N_9102,N_7135,N_7429);
nand U9103 (N_9103,N_6371,N_5587);
and U9104 (N_9104,N_6932,N_5639);
or U9105 (N_9105,N_6097,N_6868);
or U9106 (N_9106,N_6195,N_6643);
nand U9107 (N_9107,N_5789,N_5332);
and U9108 (N_9108,N_7275,N_5515);
nor U9109 (N_9109,N_6520,N_6578);
nand U9110 (N_9110,N_5233,N_5578);
nor U9111 (N_9111,N_5527,N_6103);
nand U9112 (N_9112,N_5848,N_6033);
and U9113 (N_9113,N_6395,N_6510);
or U9114 (N_9114,N_6313,N_7218);
or U9115 (N_9115,N_5888,N_6314);
or U9116 (N_9116,N_5608,N_5874);
nor U9117 (N_9117,N_6351,N_5447);
or U9118 (N_9118,N_7389,N_7267);
nor U9119 (N_9119,N_7099,N_6446);
and U9120 (N_9120,N_6224,N_6085);
and U9121 (N_9121,N_5755,N_6430);
nor U9122 (N_9122,N_6321,N_6020);
nor U9123 (N_9123,N_7400,N_6777);
nand U9124 (N_9124,N_6832,N_7494);
or U9125 (N_9125,N_5138,N_6341);
nor U9126 (N_9126,N_6537,N_6306);
nand U9127 (N_9127,N_5873,N_5461);
nor U9128 (N_9128,N_6611,N_6395);
or U9129 (N_9129,N_6256,N_5289);
nor U9130 (N_9130,N_5861,N_5761);
or U9131 (N_9131,N_6212,N_5082);
nand U9132 (N_9132,N_5472,N_7032);
nor U9133 (N_9133,N_5538,N_5663);
nor U9134 (N_9134,N_7399,N_5708);
or U9135 (N_9135,N_6132,N_5563);
and U9136 (N_9136,N_5956,N_6240);
and U9137 (N_9137,N_5439,N_7215);
or U9138 (N_9138,N_7073,N_5151);
xnor U9139 (N_9139,N_5970,N_6571);
nand U9140 (N_9140,N_5367,N_5066);
nand U9141 (N_9141,N_5959,N_6346);
nand U9142 (N_9142,N_7313,N_5966);
nor U9143 (N_9143,N_5178,N_5182);
and U9144 (N_9144,N_5118,N_6088);
nor U9145 (N_9145,N_6302,N_6144);
or U9146 (N_9146,N_5739,N_6772);
and U9147 (N_9147,N_7001,N_7057);
nor U9148 (N_9148,N_5325,N_6503);
nand U9149 (N_9149,N_6119,N_5450);
and U9150 (N_9150,N_7133,N_5986);
or U9151 (N_9151,N_5170,N_6357);
nor U9152 (N_9152,N_5028,N_5407);
or U9153 (N_9153,N_6867,N_7070);
or U9154 (N_9154,N_6833,N_7123);
and U9155 (N_9155,N_6448,N_6277);
or U9156 (N_9156,N_7292,N_5105);
xor U9157 (N_9157,N_5685,N_7192);
nor U9158 (N_9158,N_5963,N_6272);
nand U9159 (N_9159,N_6175,N_7044);
nor U9160 (N_9160,N_7133,N_5551);
and U9161 (N_9161,N_5273,N_5347);
and U9162 (N_9162,N_6000,N_5498);
nor U9163 (N_9163,N_7448,N_5280);
nor U9164 (N_9164,N_6089,N_5202);
nor U9165 (N_9165,N_7261,N_6735);
nor U9166 (N_9166,N_5134,N_6724);
nand U9167 (N_9167,N_5037,N_7488);
and U9168 (N_9168,N_6093,N_6954);
and U9169 (N_9169,N_5536,N_5370);
and U9170 (N_9170,N_6956,N_5139);
nor U9171 (N_9171,N_5761,N_5890);
and U9172 (N_9172,N_5845,N_5270);
nand U9173 (N_9173,N_5537,N_6725);
or U9174 (N_9174,N_7145,N_7460);
nand U9175 (N_9175,N_7430,N_6484);
nor U9176 (N_9176,N_5198,N_6716);
nand U9177 (N_9177,N_6894,N_5833);
nand U9178 (N_9178,N_6729,N_6683);
xor U9179 (N_9179,N_5505,N_7315);
nand U9180 (N_9180,N_6980,N_6720);
nor U9181 (N_9181,N_5828,N_5974);
nor U9182 (N_9182,N_5455,N_7285);
or U9183 (N_9183,N_6845,N_5820);
or U9184 (N_9184,N_7219,N_6950);
or U9185 (N_9185,N_6183,N_6233);
nand U9186 (N_9186,N_7439,N_7308);
nor U9187 (N_9187,N_6118,N_5864);
and U9188 (N_9188,N_7006,N_7314);
nor U9189 (N_9189,N_6357,N_5235);
xnor U9190 (N_9190,N_6773,N_7200);
and U9191 (N_9191,N_5342,N_6236);
nand U9192 (N_9192,N_7352,N_6011);
nor U9193 (N_9193,N_5996,N_6050);
nand U9194 (N_9194,N_5064,N_5446);
nor U9195 (N_9195,N_6687,N_6892);
and U9196 (N_9196,N_7081,N_6896);
nor U9197 (N_9197,N_6971,N_5150);
nor U9198 (N_9198,N_6237,N_7244);
nor U9199 (N_9199,N_7393,N_5847);
xnor U9200 (N_9200,N_5017,N_5163);
nand U9201 (N_9201,N_7015,N_5993);
nand U9202 (N_9202,N_6767,N_6207);
or U9203 (N_9203,N_5579,N_6626);
nand U9204 (N_9204,N_7160,N_5527);
nand U9205 (N_9205,N_7182,N_7379);
nand U9206 (N_9206,N_6518,N_6233);
and U9207 (N_9207,N_5786,N_5630);
nor U9208 (N_9208,N_7381,N_7273);
or U9209 (N_9209,N_7253,N_5078);
and U9210 (N_9210,N_6651,N_6346);
and U9211 (N_9211,N_5219,N_5723);
nand U9212 (N_9212,N_6329,N_7130);
nand U9213 (N_9213,N_6442,N_5073);
nor U9214 (N_9214,N_6370,N_6222);
nand U9215 (N_9215,N_5104,N_7458);
nand U9216 (N_9216,N_6436,N_6132);
and U9217 (N_9217,N_5205,N_6892);
and U9218 (N_9218,N_5602,N_5474);
nand U9219 (N_9219,N_5362,N_6348);
or U9220 (N_9220,N_6884,N_5484);
nor U9221 (N_9221,N_6012,N_6586);
or U9222 (N_9222,N_5358,N_5486);
and U9223 (N_9223,N_7224,N_7416);
nand U9224 (N_9224,N_7292,N_6055);
or U9225 (N_9225,N_6625,N_7244);
or U9226 (N_9226,N_6770,N_6942);
nand U9227 (N_9227,N_5231,N_7413);
or U9228 (N_9228,N_6647,N_6609);
and U9229 (N_9229,N_5467,N_6626);
or U9230 (N_9230,N_5165,N_5871);
or U9231 (N_9231,N_6417,N_5066);
or U9232 (N_9232,N_5416,N_5963);
and U9233 (N_9233,N_5317,N_6973);
nand U9234 (N_9234,N_6850,N_5525);
or U9235 (N_9235,N_5146,N_5562);
and U9236 (N_9236,N_5814,N_5752);
and U9237 (N_9237,N_7022,N_6950);
nand U9238 (N_9238,N_6687,N_5623);
or U9239 (N_9239,N_5497,N_5130);
and U9240 (N_9240,N_5419,N_6146);
nor U9241 (N_9241,N_5124,N_7044);
and U9242 (N_9242,N_5477,N_7390);
nor U9243 (N_9243,N_7282,N_5448);
nor U9244 (N_9244,N_6176,N_5359);
and U9245 (N_9245,N_5959,N_6945);
nand U9246 (N_9246,N_7204,N_6549);
nor U9247 (N_9247,N_5806,N_6298);
nor U9248 (N_9248,N_5205,N_5240);
and U9249 (N_9249,N_5099,N_6175);
or U9250 (N_9250,N_7262,N_6845);
or U9251 (N_9251,N_6501,N_5922);
xor U9252 (N_9252,N_6365,N_7184);
nor U9253 (N_9253,N_6469,N_6611);
and U9254 (N_9254,N_5508,N_5851);
nor U9255 (N_9255,N_6201,N_7359);
nand U9256 (N_9256,N_6586,N_5061);
nand U9257 (N_9257,N_6059,N_5341);
nor U9258 (N_9258,N_6619,N_6926);
and U9259 (N_9259,N_6750,N_5728);
nor U9260 (N_9260,N_6505,N_5528);
or U9261 (N_9261,N_7223,N_5650);
or U9262 (N_9262,N_5177,N_7182);
and U9263 (N_9263,N_6112,N_7102);
or U9264 (N_9264,N_6351,N_6273);
and U9265 (N_9265,N_6942,N_6420);
and U9266 (N_9266,N_5727,N_5686);
or U9267 (N_9267,N_5141,N_6932);
nand U9268 (N_9268,N_5881,N_7073);
nor U9269 (N_9269,N_6758,N_6164);
or U9270 (N_9270,N_6758,N_6048);
nor U9271 (N_9271,N_5907,N_5254);
and U9272 (N_9272,N_6906,N_5067);
and U9273 (N_9273,N_7101,N_6829);
or U9274 (N_9274,N_6281,N_6714);
nand U9275 (N_9275,N_5943,N_5522);
nand U9276 (N_9276,N_7171,N_6002);
nor U9277 (N_9277,N_7218,N_6341);
and U9278 (N_9278,N_5117,N_5551);
nor U9279 (N_9279,N_5412,N_6948);
or U9280 (N_9280,N_7367,N_7181);
or U9281 (N_9281,N_5742,N_6545);
nand U9282 (N_9282,N_7341,N_5020);
nand U9283 (N_9283,N_7063,N_5399);
and U9284 (N_9284,N_5214,N_5429);
and U9285 (N_9285,N_5597,N_5404);
nand U9286 (N_9286,N_5027,N_6108);
or U9287 (N_9287,N_7180,N_5532);
xor U9288 (N_9288,N_5025,N_5649);
nand U9289 (N_9289,N_7395,N_5035);
or U9290 (N_9290,N_5289,N_6360);
nor U9291 (N_9291,N_5458,N_6666);
nor U9292 (N_9292,N_5309,N_7485);
or U9293 (N_9293,N_7457,N_6034);
nand U9294 (N_9294,N_6529,N_5846);
or U9295 (N_9295,N_6231,N_7211);
nand U9296 (N_9296,N_6571,N_5077);
xor U9297 (N_9297,N_7184,N_7130);
or U9298 (N_9298,N_5403,N_6117);
and U9299 (N_9299,N_5744,N_6059);
nand U9300 (N_9300,N_7119,N_6935);
or U9301 (N_9301,N_6777,N_7027);
and U9302 (N_9302,N_5612,N_5656);
and U9303 (N_9303,N_6224,N_5445);
and U9304 (N_9304,N_5567,N_5167);
nand U9305 (N_9305,N_6132,N_5732);
and U9306 (N_9306,N_5274,N_6113);
and U9307 (N_9307,N_7191,N_6234);
nand U9308 (N_9308,N_6809,N_7346);
nor U9309 (N_9309,N_5290,N_5039);
nor U9310 (N_9310,N_7414,N_7015);
and U9311 (N_9311,N_6435,N_5406);
and U9312 (N_9312,N_5001,N_7243);
nand U9313 (N_9313,N_6989,N_6395);
nor U9314 (N_9314,N_6285,N_6631);
or U9315 (N_9315,N_6890,N_5795);
or U9316 (N_9316,N_6417,N_6105);
and U9317 (N_9317,N_6865,N_7076);
nor U9318 (N_9318,N_6387,N_6186);
nand U9319 (N_9319,N_6651,N_5754);
nor U9320 (N_9320,N_6641,N_5301);
or U9321 (N_9321,N_5288,N_5914);
and U9322 (N_9322,N_5561,N_6210);
and U9323 (N_9323,N_6256,N_6476);
or U9324 (N_9324,N_6113,N_5605);
or U9325 (N_9325,N_5852,N_6551);
nand U9326 (N_9326,N_6675,N_6949);
and U9327 (N_9327,N_7257,N_5387);
xnor U9328 (N_9328,N_6737,N_6653);
nand U9329 (N_9329,N_6843,N_5372);
and U9330 (N_9330,N_5415,N_6636);
nand U9331 (N_9331,N_5265,N_5260);
or U9332 (N_9332,N_5400,N_6409);
nor U9333 (N_9333,N_5663,N_6281);
nor U9334 (N_9334,N_7018,N_5141);
and U9335 (N_9335,N_5650,N_5029);
and U9336 (N_9336,N_6143,N_6721);
or U9337 (N_9337,N_5211,N_6412);
xnor U9338 (N_9338,N_5037,N_5910);
nand U9339 (N_9339,N_6151,N_6048);
nor U9340 (N_9340,N_7431,N_5632);
or U9341 (N_9341,N_5721,N_6051);
nor U9342 (N_9342,N_5096,N_6314);
nand U9343 (N_9343,N_6757,N_5071);
nor U9344 (N_9344,N_5275,N_6065);
nand U9345 (N_9345,N_6775,N_6102);
nor U9346 (N_9346,N_5982,N_5852);
and U9347 (N_9347,N_5993,N_6821);
or U9348 (N_9348,N_5537,N_6797);
and U9349 (N_9349,N_5724,N_5001);
and U9350 (N_9350,N_5409,N_5138);
or U9351 (N_9351,N_5513,N_5617);
and U9352 (N_9352,N_5805,N_5890);
nor U9353 (N_9353,N_5076,N_5979);
nand U9354 (N_9354,N_5134,N_5828);
and U9355 (N_9355,N_7260,N_7243);
nand U9356 (N_9356,N_5043,N_6336);
nor U9357 (N_9357,N_6743,N_5483);
nand U9358 (N_9358,N_5419,N_6050);
xor U9359 (N_9359,N_6500,N_6973);
nor U9360 (N_9360,N_7378,N_5947);
or U9361 (N_9361,N_7211,N_5792);
nor U9362 (N_9362,N_6355,N_6495);
or U9363 (N_9363,N_5927,N_6685);
nor U9364 (N_9364,N_5387,N_6866);
nor U9365 (N_9365,N_6685,N_5420);
or U9366 (N_9366,N_5193,N_6544);
xnor U9367 (N_9367,N_5229,N_5976);
or U9368 (N_9368,N_6294,N_5013);
and U9369 (N_9369,N_5184,N_5691);
nand U9370 (N_9370,N_5002,N_5842);
and U9371 (N_9371,N_5187,N_5611);
or U9372 (N_9372,N_6576,N_6489);
and U9373 (N_9373,N_6527,N_6862);
nor U9374 (N_9374,N_5303,N_6797);
and U9375 (N_9375,N_6881,N_5024);
and U9376 (N_9376,N_6201,N_7160);
xnor U9377 (N_9377,N_7354,N_6745);
nor U9378 (N_9378,N_6688,N_5442);
and U9379 (N_9379,N_5823,N_6558);
nand U9380 (N_9380,N_6457,N_6943);
or U9381 (N_9381,N_6974,N_5527);
nor U9382 (N_9382,N_6193,N_6501);
and U9383 (N_9383,N_5383,N_7247);
or U9384 (N_9384,N_6440,N_7140);
nor U9385 (N_9385,N_5755,N_7208);
and U9386 (N_9386,N_7258,N_7058);
or U9387 (N_9387,N_5176,N_5027);
or U9388 (N_9388,N_6928,N_6236);
nor U9389 (N_9389,N_5419,N_5704);
nor U9390 (N_9390,N_6319,N_5220);
and U9391 (N_9391,N_6855,N_6048);
nand U9392 (N_9392,N_5173,N_6915);
or U9393 (N_9393,N_6483,N_6957);
and U9394 (N_9394,N_6715,N_6732);
or U9395 (N_9395,N_5593,N_6583);
nand U9396 (N_9396,N_7208,N_5960);
nand U9397 (N_9397,N_7294,N_5955);
nand U9398 (N_9398,N_7394,N_5416);
nor U9399 (N_9399,N_5151,N_7049);
nand U9400 (N_9400,N_6233,N_6234);
and U9401 (N_9401,N_5709,N_5248);
nand U9402 (N_9402,N_6034,N_7042);
and U9403 (N_9403,N_5918,N_5608);
nor U9404 (N_9404,N_5113,N_6536);
and U9405 (N_9405,N_6090,N_5006);
or U9406 (N_9406,N_7057,N_6770);
and U9407 (N_9407,N_7425,N_7089);
nand U9408 (N_9408,N_6863,N_5683);
or U9409 (N_9409,N_5195,N_7422);
and U9410 (N_9410,N_5953,N_7210);
or U9411 (N_9411,N_5367,N_5837);
and U9412 (N_9412,N_5021,N_5240);
nor U9413 (N_9413,N_6524,N_6380);
nor U9414 (N_9414,N_6231,N_6601);
nor U9415 (N_9415,N_6056,N_5169);
or U9416 (N_9416,N_7211,N_7262);
nor U9417 (N_9417,N_5280,N_5252);
nand U9418 (N_9418,N_5714,N_7053);
or U9419 (N_9419,N_7194,N_5446);
and U9420 (N_9420,N_6912,N_7017);
nor U9421 (N_9421,N_5663,N_6064);
and U9422 (N_9422,N_6496,N_5325);
or U9423 (N_9423,N_5927,N_6251);
nor U9424 (N_9424,N_6679,N_5783);
nor U9425 (N_9425,N_6814,N_7249);
nor U9426 (N_9426,N_7387,N_6943);
and U9427 (N_9427,N_7308,N_5531);
nand U9428 (N_9428,N_6014,N_6522);
nand U9429 (N_9429,N_5284,N_5018);
nor U9430 (N_9430,N_5093,N_7153);
and U9431 (N_9431,N_6452,N_5094);
nor U9432 (N_9432,N_5810,N_6340);
nand U9433 (N_9433,N_7404,N_7366);
and U9434 (N_9434,N_7167,N_5114);
nor U9435 (N_9435,N_6447,N_5633);
nand U9436 (N_9436,N_5419,N_7491);
and U9437 (N_9437,N_5909,N_6161);
nor U9438 (N_9438,N_7113,N_6903);
xnor U9439 (N_9439,N_6034,N_7267);
and U9440 (N_9440,N_5942,N_5569);
and U9441 (N_9441,N_7498,N_6875);
and U9442 (N_9442,N_6363,N_6845);
or U9443 (N_9443,N_6798,N_5486);
nor U9444 (N_9444,N_5527,N_5792);
or U9445 (N_9445,N_6170,N_5239);
and U9446 (N_9446,N_5463,N_6969);
or U9447 (N_9447,N_5759,N_5271);
or U9448 (N_9448,N_6018,N_5221);
and U9449 (N_9449,N_7319,N_5712);
nand U9450 (N_9450,N_6564,N_6269);
and U9451 (N_9451,N_6329,N_6697);
or U9452 (N_9452,N_5399,N_5343);
and U9453 (N_9453,N_5185,N_5181);
or U9454 (N_9454,N_6504,N_6369);
nand U9455 (N_9455,N_5494,N_5844);
nor U9456 (N_9456,N_5395,N_5903);
or U9457 (N_9457,N_5677,N_6820);
nor U9458 (N_9458,N_5722,N_5276);
nand U9459 (N_9459,N_6164,N_6367);
nor U9460 (N_9460,N_6260,N_5022);
and U9461 (N_9461,N_6452,N_7320);
nand U9462 (N_9462,N_6461,N_5143);
nor U9463 (N_9463,N_5960,N_7158);
nand U9464 (N_9464,N_6406,N_6588);
or U9465 (N_9465,N_7129,N_7359);
or U9466 (N_9466,N_5183,N_7479);
nor U9467 (N_9467,N_5638,N_7063);
nor U9468 (N_9468,N_6436,N_6112);
nor U9469 (N_9469,N_6170,N_5515);
xnor U9470 (N_9470,N_6399,N_5650);
nand U9471 (N_9471,N_7227,N_5188);
or U9472 (N_9472,N_5860,N_7472);
nor U9473 (N_9473,N_6934,N_5725);
or U9474 (N_9474,N_7309,N_6295);
nand U9475 (N_9475,N_6552,N_6715);
nor U9476 (N_9476,N_6892,N_5194);
nand U9477 (N_9477,N_6060,N_7156);
xnor U9478 (N_9478,N_5354,N_7425);
and U9479 (N_9479,N_7441,N_7083);
nand U9480 (N_9480,N_5702,N_7137);
or U9481 (N_9481,N_6928,N_6577);
and U9482 (N_9482,N_5400,N_6191);
or U9483 (N_9483,N_5428,N_6443);
and U9484 (N_9484,N_6249,N_6016);
nor U9485 (N_9485,N_6996,N_5121);
nand U9486 (N_9486,N_5992,N_5678);
and U9487 (N_9487,N_6794,N_6824);
or U9488 (N_9488,N_7316,N_6664);
or U9489 (N_9489,N_6890,N_7215);
nand U9490 (N_9490,N_6584,N_6321);
or U9491 (N_9491,N_5157,N_6924);
and U9492 (N_9492,N_6941,N_6055);
nor U9493 (N_9493,N_5107,N_5941);
and U9494 (N_9494,N_6783,N_5535);
or U9495 (N_9495,N_5125,N_7495);
or U9496 (N_9496,N_6368,N_5211);
or U9497 (N_9497,N_6100,N_6930);
and U9498 (N_9498,N_6453,N_6801);
and U9499 (N_9499,N_6666,N_6173);
or U9500 (N_9500,N_5665,N_5212);
nand U9501 (N_9501,N_6484,N_5185);
and U9502 (N_9502,N_7007,N_6292);
nor U9503 (N_9503,N_5779,N_7035);
or U9504 (N_9504,N_5108,N_6342);
nor U9505 (N_9505,N_5803,N_6611);
nand U9506 (N_9506,N_5054,N_6345);
nand U9507 (N_9507,N_7177,N_5939);
nor U9508 (N_9508,N_5999,N_7274);
nor U9509 (N_9509,N_5700,N_5895);
nand U9510 (N_9510,N_5211,N_6060);
nor U9511 (N_9511,N_7382,N_6862);
nand U9512 (N_9512,N_7369,N_5957);
nor U9513 (N_9513,N_6399,N_6592);
xnor U9514 (N_9514,N_5063,N_5765);
or U9515 (N_9515,N_7275,N_6474);
and U9516 (N_9516,N_7028,N_5429);
and U9517 (N_9517,N_7223,N_5997);
and U9518 (N_9518,N_6369,N_5384);
nor U9519 (N_9519,N_5829,N_6454);
nand U9520 (N_9520,N_6809,N_5878);
and U9521 (N_9521,N_6769,N_7122);
or U9522 (N_9522,N_7452,N_7427);
nor U9523 (N_9523,N_6368,N_5609);
and U9524 (N_9524,N_6496,N_6505);
xnor U9525 (N_9525,N_6374,N_6675);
nor U9526 (N_9526,N_6474,N_6851);
nand U9527 (N_9527,N_7442,N_5312);
or U9528 (N_9528,N_5432,N_5615);
and U9529 (N_9529,N_6520,N_5180);
or U9530 (N_9530,N_5131,N_6213);
nor U9531 (N_9531,N_6871,N_6815);
nand U9532 (N_9532,N_7430,N_7132);
nand U9533 (N_9533,N_6697,N_6825);
nor U9534 (N_9534,N_6803,N_5618);
and U9535 (N_9535,N_5500,N_7259);
nor U9536 (N_9536,N_5389,N_6273);
and U9537 (N_9537,N_7393,N_5813);
and U9538 (N_9538,N_7249,N_6065);
nor U9539 (N_9539,N_7060,N_6367);
nor U9540 (N_9540,N_7025,N_6052);
or U9541 (N_9541,N_5441,N_6138);
or U9542 (N_9542,N_5768,N_7023);
nor U9543 (N_9543,N_7379,N_5056);
nor U9544 (N_9544,N_6780,N_6605);
nand U9545 (N_9545,N_7090,N_6237);
nand U9546 (N_9546,N_5099,N_5989);
nand U9547 (N_9547,N_5487,N_7462);
and U9548 (N_9548,N_5707,N_6895);
xor U9549 (N_9549,N_5044,N_5571);
nor U9550 (N_9550,N_7452,N_6088);
nand U9551 (N_9551,N_5385,N_7191);
nor U9552 (N_9552,N_5161,N_5755);
nor U9553 (N_9553,N_6657,N_6186);
or U9554 (N_9554,N_7414,N_5069);
nand U9555 (N_9555,N_6971,N_6851);
and U9556 (N_9556,N_5674,N_6344);
nor U9557 (N_9557,N_6313,N_5471);
nor U9558 (N_9558,N_6742,N_7246);
or U9559 (N_9559,N_6960,N_5436);
nand U9560 (N_9560,N_5710,N_5246);
or U9561 (N_9561,N_7458,N_6200);
nor U9562 (N_9562,N_6669,N_5145);
nor U9563 (N_9563,N_7080,N_5812);
or U9564 (N_9564,N_6648,N_6877);
or U9565 (N_9565,N_6452,N_5446);
or U9566 (N_9566,N_6782,N_5874);
or U9567 (N_9567,N_7024,N_5109);
nor U9568 (N_9568,N_5239,N_6894);
and U9569 (N_9569,N_6826,N_7188);
or U9570 (N_9570,N_6003,N_7079);
and U9571 (N_9571,N_6485,N_5130);
nor U9572 (N_9572,N_5716,N_6229);
nor U9573 (N_9573,N_5436,N_5471);
nor U9574 (N_9574,N_6554,N_5577);
nor U9575 (N_9575,N_6622,N_7408);
or U9576 (N_9576,N_5626,N_7330);
and U9577 (N_9577,N_6453,N_7325);
nand U9578 (N_9578,N_5677,N_5736);
nor U9579 (N_9579,N_5700,N_6336);
or U9580 (N_9580,N_6814,N_5538);
and U9581 (N_9581,N_6117,N_5013);
and U9582 (N_9582,N_6353,N_7378);
nand U9583 (N_9583,N_6463,N_7400);
and U9584 (N_9584,N_6601,N_5176);
or U9585 (N_9585,N_6250,N_5995);
and U9586 (N_9586,N_6799,N_5752);
and U9587 (N_9587,N_6306,N_6140);
nand U9588 (N_9588,N_6192,N_5518);
nand U9589 (N_9589,N_7003,N_6297);
nand U9590 (N_9590,N_5525,N_5770);
nor U9591 (N_9591,N_5414,N_5188);
nor U9592 (N_9592,N_6189,N_5181);
nand U9593 (N_9593,N_5517,N_6653);
and U9594 (N_9594,N_6899,N_6559);
nor U9595 (N_9595,N_7113,N_6586);
nand U9596 (N_9596,N_6657,N_6633);
and U9597 (N_9597,N_6703,N_5111);
or U9598 (N_9598,N_6791,N_5821);
and U9599 (N_9599,N_5266,N_6953);
nand U9600 (N_9600,N_5909,N_6920);
nand U9601 (N_9601,N_5720,N_7120);
and U9602 (N_9602,N_6253,N_6962);
nor U9603 (N_9603,N_6266,N_7289);
xnor U9604 (N_9604,N_7473,N_5077);
nand U9605 (N_9605,N_7498,N_5463);
and U9606 (N_9606,N_7263,N_5205);
and U9607 (N_9607,N_7420,N_6246);
nand U9608 (N_9608,N_7082,N_5573);
or U9609 (N_9609,N_6851,N_5302);
and U9610 (N_9610,N_6685,N_5705);
and U9611 (N_9611,N_5146,N_6959);
nor U9612 (N_9612,N_7089,N_5055);
xnor U9613 (N_9613,N_6291,N_6166);
nor U9614 (N_9614,N_5903,N_5672);
or U9615 (N_9615,N_7469,N_5527);
nor U9616 (N_9616,N_6617,N_6633);
nor U9617 (N_9617,N_6441,N_5571);
nor U9618 (N_9618,N_5415,N_7094);
nor U9619 (N_9619,N_7058,N_6267);
and U9620 (N_9620,N_6741,N_5397);
and U9621 (N_9621,N_5224,N_6935);
nor U9622 (N_9622,N_5418,N_6648);
or U9623 (N_9623,N_5186,N_7112);
or U9624 (N_9624,N_7499,N_6190);
and U9625 (N_9625,N_5278,N_6457);
nand U9626 (N_9626,N_6070,N_7383);
nor U9627 (N_9627,N_6360,N_7424);
and U9628 (N_9628,N_6617,N_7245);
or U9629 (N_9629,N_5591,N_5695);
nor U9630 (N_9630,N_6699,N_7180);
xnor U9631 (N_9631,N_6549,N_5611);
nor U9632 (N_9632,N_5014,N_5819);
nand U9633 (N_9633,N_7315,N_7491);
nor U9634 (N_9634,N_5550,N_6639);
nor U9635 (N_9635,N_7262,N_6010);
nand U9636 (N_9636,N_5591,N_5658);
nor U9637 (N_9637,N_5006,N_7313);
nand U9638 (N_9638,N_5828,N_5298);
and U9639 (N_9639,N_5301,N_7471);
nand U9640 (N_9640,N_6674,N_6518);
or U9641 (N_9641,N_6128,N_5609);
and U9642 (N_9642,N_6150,N_6990);
and U9643 (N_9643,N_6735,N_7149);
nand U9644 (N_9644,N_6364,N_6736);
nand U9645 (N_9645,N_6089,N_6085);
or U9646 (N_9646,N_6071,N_5178);
and U9647 (N_9647,N_6310,N_5937);
nand U9648 (N_9648,N_6911,N_5841);
xnor U9649 (N_9649,N_7299,N_5257);
nand U9650 (N_9650,N_6650,N_5202);
nand U9651 (N_9651,N_6148,N_6447);
xor U9652 (N_9652,N_5800,N_6517);
or U9653 (N_9653,N_6971,N_6378);
nor U9654 (N_9654,N_6930,N_6385);
nand U9655 (N_9655,N_7491,N_6683);
and U9656 (N_9656,N_6037,N_7386);
nor U9657 (N_9657,N_7421,N_6750);
nor U9658 (N_9658,N_6440,N_5601);
nand U9659 (N_9659,N_6334,N_5445);
nor U9660 (N_9660,N_5415,N_6887);
or U9661 (N_9661,N_7256,N_6952);
nor U9662 (N_9662,N_5759,N_6248);
nor U9663 (N_9663,N_6799,N_6791);
or U9664 (N_9664,N_7297,N_6507);
or U9665 (N_9665,N_5770,N_7095);
or U9666 (N_9666,N_6378,N_6500);
and U9667 (N_9667,N_5328,N_6615);
and U9668 (N_9668,N_6729,N_6365);
nand U9669 (N_9669,N_5693,N_6150);
or U9670 (N_9670,N_6017,N_6150);
and U9671 (N_9671,N_5054,N_6470);
and U9672 (N_9672,N_6861,N_6364);
and U9673 (N_9673,N_5874,N_5374);
and U9674 (N_9674,N_6748,N_6096);
or U9675 (N_9675,N_7465,N_5540);
nand U9676 (N_9676,N_5645,N_6501);
and U9677 (N_9677,N_6966,N_5812);
nor U9678 (N_9678,N_7204,N_5178);
and U9679 (N_9679,N_7187,N_5063);
nand U9680 (N_9680,N_6472,N_5931);
nand U9681 (N_9681,N_6976,N_6317);
and U9682 (N_9682,N_5686,N_5454);
nand U9683 (N_9683,N_5055,N_5464);
and U9684 (N_9684,N_6408,N_6898);
nor U9685 (N_9685,N_7414,N_6770);
or U9686 (N_9686,N_6212,N_5251);
nand U9687 (N_9687,N_5440,N_6542);
and U9688 (N_9688,N_5403,N_7322);
or U9689 (N_9689,N_5774,N_5009);
and U9690 (N_9690,N_5619,N_6244);
and U9691 (N_9691,N_5797,N_5033);
nand U9692 (N_9692,N_5596,N_7486);
and U9693 (N_9693,N_5078,N_5515);
and U9694 (N_9694,N_5540,N_5388);
nand U9695 (N_9695,N_6996,N_5589);
nor U9696 (N_9696,N_6944,N_5411);
nand U9697 (N_9697,N_6133,N_6100);
nand U9698 (N_9698,N_5196,N_6529);
or U9699 (N_9699,N_5792,N_5022);
or U9700 (N_9700,N_5261,N_7324);
nor U9701 (N_9701,N_5755,N_5415);
nor U9702 (N_9702,N_5242,N_5022);
and U9703 (N_9703,N_5277,N_6615);
or U9704 (N_9704,N_5045,N_6173);
nor U9705 (N_9705,N_5501,N_5108);
nor U9706 (N_9706,N_5542,N_7394);
or U9707 (N_9707,N_7174,N_6818);
or U9708 (N_9708,N_6075,N_5042);
nand U9709 (N_9709,N_7461,N_5425);
nor U9710 (N_9710,N_7292,N_5620);
or U9711 (N_9711,N_5345,N_5997);
or U9712 (N_9712,N_6929,N_7104);
nand U9713 (N_9713,N_5725,N_6539);
nand U9714 (N_9714,N_5306,N_5334);
nand U9715 (N_9715,N_5174,N_5742);
and U9716 (N_9716,N_7055,N_5081);
or U9717 (N_9717,N_7070,N_7238);
or U9718 (N_9718,N_7190,N_6644);
and U9719 (N_9719,N_6253,N_5820);
and U9720 (N_9720,N_5648,N_6247);
or U9721 (N_9721,N_7425,N_6765);
nand U9722 (N_9722,N_5041,N_6452);
or U9723 (N_9723,N_6278,N_7248);
nor U9724 (N_9724,N_7110,N_5546);
nand U9725 (N_9725,N_5915,N_7350);
or U9726 (N_9726,N_6655,N_6081);
and U9727 (N_9727,N_5340,N_7155);
and U9728 (N_9728,N_7061,N_6223);
or U9729 (N_9729,N_7351,N_7240);
or U9730 (N_9730,N_7086,N_7380);
nor U9731 (N_9731,N_5828,N_7248);
nand U9732 (N_9732,N_7261,N_5936);
nand U9733 (N_9733,N_6125,N_5521);
nand U9734 (N_9734,N_6914,N_5174);
and U9735 (N_9735,N_5275,N_6209);
nand U9736 (N_9736,N_6955,N_6281);
and U9737 (N_9737,N_7090,N_5584);
nor U9738 (N_9738,N_6170,N_5762);
nor U9739 (N_9739,N_7298,N_6518);
nor U9740 (N_9740,N_6998,N_5562);
or U9741 (N_9741,N_5805,N_6800);
nand U9742 (N_9742,N_6672,N_6303);
nand U9743 (N_9743,N_6709,N_5625);
nand U9744 (N_9744,N_5980,N_5969);
and U9745 (N_9745,N_6081,N_6745);
nand U9746 (N_9746,N_6847,N_5988);
and U9747 (N_9747,N_7212,N_7478);
and U9748 (N_9748,N_6085,N_5013);
or U9749 (N_9749,N_6645,N_6582);
and U9750 (N_9750,N_5291,N_7102);
and U9751 (N_9751,N_6403,N_5336);
nand U9752 (N_9752,N_6234,N_6132);
or U9753 (N_9753,N_6736,N_5334);
and U9754 (N_9754,N_5054,N_5285);
nand U9755 (N_9755,N_6708,N_5110);
nand U9756 (N_9756,N_6477,N_5222);
or U9757 (N_9757,N_7018,N_6642);
nor U9758 (N_9758,N_5814,N_7442);
or U9759 (N_9759,N_5198,N_5404);
nor U9760 (N_9760,N_6823,N_7382);
or U9761 (N_9761,N_6887,N_5038);
or U9762 (N_9762,N_7355,N_6535);
nand U9763 (N_9763,N_5227,N_5953);
and U9764 (N_9764,N_7085,N_6035);
and U9765 (N_9765,N_6636,N_5859);
and U9766 (N_9766,N_6867,N_5240);
xor U9767 (N_9767,N_6969,N_5904);
or U9768 (N_9768,N_6351,N_7433);
nor U9769 (N_9769,N_6088,N_6883);
xor U9770 (N_9770,N_5583,N_6117);
nor U9771 (N_9771,N_5255,N_7130);
or U9772 (N_9772,N_7186,N_6166);
and U9773 (N_9773,N_6608,N_6917);
nor U9774 (N_9774,N_6476,N_5747);
or U9775 (N_9775,N_5771,N_5854);
nand U9776 (N_9776,N_7069,N_6558);
and U9777 (N_9777,N_7457,N_6110);
nand U9778 (N_9778,N_5405,N_6776);
and U9779 (N_9779,N_7184,N_5128);
nand U9780 (N_9780,N_5957,N_5877);
or U9781 (N_9781,N_6898,N_6825);
and U9782 (N_9782,N_5719,N_6366);
nand U9783 (N_9783,N_6124,N_6185);
or U9784 (N_9784,N_5122,N_6826);
and U9785 (N_9785,N_5136,N_7421);
nor U9786 (N_9786,N_5431,N_6283);
or U9787 (N_9787,N_6459,N_5115);
nor U9788 (N_9788,N_6352,N_5032);
nand U9789 (N_9789,N_6414,N_5436);
nor U9790 (N_9790,N_6979,N_6873);
nand U9791 (N_9791,N_6097,N_6303);
or U9792 (N_9792,N_5243,N_6482);
or U9793 (N_9793,N_6091,N_6727);
nor U9794 (N_9794,N_5515,N_6883);
nor U9795 (N_9795,N_5626,N_6223);
xnor U9796 (N_9796,N_6177,N_6796);
or U9797 (N_9797,N_5166,N_6681);
nand U9798 (N_9798,N_6922,N_7063);
nand U9799 (N_9799,N_6895,N_6875);
nand U9800 (N_9800,N_6744,N_6556);
or U9801 (N_9801,N_6103,N_5404);
or U9802 (N_9802,N_6948,N_6898);
or U9803 (N_9803,N_7366,N_5711);
nor U9804 (N_9804,N_5240,N_6685);
nand U9805 (N_9805,N_5192,N_6547);
nor U9806 (N_9806,N_6652,N_5973);
nor U9807 (N_9807,N_6073,N_7383);
or U9808 (N_9808,N_7330,N_5995);
nand U9809 (N_9809,N_5268,N_5749);
and U9810 (N_9810,N_6024,N_6387);
nor U9811 (N_9811,N_5099,N_6591);
nor U9812 (N_9812,N_5536,N_6611);
nand U9813 (N_9813,N_5214,N_6970);
or U9814 (N_9814,N_6139,N_6124);
nor U9815 (N_9815,N_6137,N_6492);
nand U9816 (N_9816,N_6088,N_7462);
nor U9817 (N_9817,N_6365,N_6141);
or U9818 (N_9818,N_6595,N_7225);
or U9819 (N_9819,N_5288,N_5301);
or U9820 (N_9820,N_5709,N_7464);
nor U9821 (N_9821,N_6209,N_7464);
nand U9822 (N_9822,N_6330,N_7226);
and U9823 (N_9823,N_5245,N_7174);
or U9824 (N_9824,N_7458,N_7321);
nor U9825 (N_9825,N_6100,N_6894);
or U9826 (N_9826,N_6319,N_5248);
and U9827 (N_9827,N_7379,N_6724);
or U9828 (N_9828,N_5053,N_6227);
nor U9829 (N_9829,N_7350,N_6561);
nand U9830 (N_9830,N_6256,N_7382);
or U9831 (N_9831,N_6126,N_5693);
and U9832 (N_9832,N_5427,N_6173);
or U9833 (N_9833,N_6962,N_7354);
nor U9834 (N_9834,N_5734,N_5301);
nand U9835 (N_9835,N_6134,N_6374);
and U9836 (N_9836,N_7190,N_7272);
or U9837 (N_9837,N_7065,N_7123);
and U9838 (N_9838,N_5422,N_6231);
nand U9839 (N_9839,N_6036,N_5494);
nand U9840 (N_9840,N_5184,N_6793);
nand U9841 (N_9841,N_7408,N_7444);
and U9842 (N_9842,N_7386,N_7192);
and U9843 (N_9843,N_6010,N_6671);
nand U9844 (N_9844,N_5644,N_5210);
and U9845 (N_9845,N_6277,N_6815);
nand U9846 (N_9846,N_6110,N_6331);
nor U9847 (N_9847,N_5334,N_6628);
or U9848 (N_9848,N_6566,N_6547);
or U9849 (N_9849,N_6657,N_6742);
and U9850 (N_9850,N_5827,N_5521);
nand U9851 (N_9851,N_5663,N_5763);
or U9852 (N_9852,N_6638,N_7349);
and U9853 (N_9853,N_6519,N_7351);
and U9854 (N_9854,N_5205,N_5349);
and U9855 (N_9855,N_5402,N_5053);
or U9856 (N_9856,N_6608,N_6928);
and U9857 (N_9857,N_6079,N_7466);
or U9858 (N_9858,N_5945,N_6820);
nand U9859 (N_9859,N_7253,N_5182);
nor U9860 (N_9860,N_5049,N_5391);
nand U9861 (N_9861,N_6617,N_6029);
or U9862 (N_9862,N_7277,N_5378);
xnor U9863 (N_9863,N_5636,N_5233);
or U9864 (N_9864,N_6456,N_6013);
nor U9865 (N_9865,N_5375,N_6713);
and U9866 (N_9866,N_5779,N_7250);
and U9867 (N_9867,N_7247,N_5663);
or U9868 (N_9868,N_6722,N_5411);
nor U9869 (N_9869,N_6680,N_7122);
nor U9870 (N_9870,N_7435,N_7418);
and U9871 (N_9871,N_5977,N_6356);
nand U9872 (N_9872,N_5623,N_5077);
and U9873 (N_9873,N_7003,N_7322);
nand U9874 (N_9874,N_6437,N_5293);
xnor U9875 (N_9875,N_5793,N_5263);
nor U9876 (N_9876,N_6018,N_6338);
nand U9877 (N_9877,N_6045,N_5120);
and U9878 (N_9878,N_6383,N_6560);
xor U9879 (N_9879,N_6246,N_7332);
nand U9880 (N_9880,N_5849,N_6854);
and U9881 (N_9881,N_5169,N_7066);
or U9882 (N_9882,N_5040,N_6033);
and U9883 (N_9883,N_6458,N_6337);
and U9884 (N_9884,N_6308,N_5805);
or U9885 (N_9885,N_6950,N_5716);
nand U9886 (N_9886,N_6993,N_6227);
and U9887 (N_9887,N_5440,N_6518);
xor U9888 (N_9888,N_6352,N_6312);
and U9889 (N_9889,N_5027,N_5588);
nor U9890 (N_9890,N_5558,N_7414);
or U9891 (N_9891,N_7048,N_6026);
xor U9892 (N_9892,N_5504,N_6353);
or U9893 (N_9893,N_6273,N_5437);
nand U9894 (N_9894,N_5137,N_6707);
nor U9895 (N_9895,N_6278,N_6250);
nand U9896 (N_9896,N_7231,N_6419);
nand U9897 (N_9897,N_6929,N_6184);
or U9898 (N_9898,N_5853,N_6474);
nand U9899 (N_9899,N_6230,N_6038);
nand U9900 (N_9900,N_6828,N_7255);
nor U9901 (N_9901,N_6908,N_6563);
nand U9902 (N_9902,N_7144,N_7014);
nand U9903 (N_9903,N_6542,N_6129);
and U9904 (N_9904,N_7399,N_6519);
xnor U9905 (N_9905,N_5640,N_5309);
and U9906 (N_9906,N_7121,N_5952);
or U9907 (N_9907,N_7469,N_5621);
and U9908 (N_9908,N_6232,N_7147);
nand U9909 (N_9909,N_5448,N_7044);
nor U9910 (N_9910,N_7022,N_6088);
nor U9911 (N_9911,N_5008,N_6233);
and U9912 (N_9912,N_6638,N_6204);
and U9913 (N_9913,N_6438,N_5009);
nor U9914 (N_9914,N_6116,N_6992);
nand U9915 (N_9915,N_5310,N_5619);
and U9916 (N_9916,N_6038,N_6233);
or U9917 (N_9917,N_6156,N_6478);
nand U9918 (N_9918,N_5787,N_5087);
nand U9919 (N_9919,N_5052,N_6041);
and U9920 (N_9920,N_6641,N_6915);
or U9921 (N_9921,N_5605,N_6987);
or U9922 (N_9922,N_5736,N_5088);
and U9923 (N_9923,N_7301,N_7228);
and U9924 (N_9924,N_5533,N_6155);
and U9925 (N_9925,N_5715,N_5763);
and U9926 (N_9926,N_6182,N_5746);
nor U9927 (N_9927,N_7457,N_7275);
or U9928 (N_9928,N_6307,N_6327);
nor U9929 (N_9929,N_7134,N_7081);
or U9930 (N_9930,N_7149,N_7110);
and U9931 (N_9931,N_6373,N_6902);
nor U9932 (N_9932,N_5927,N_7421);
nand U9933 (N_9933,N_7463,N_6199);
nand U9934 (N_9934,N_5038,N_7117);
and U9935 (N_9935,N_6996,N_6465);
nor U9936 (N_9936,N_7167,N_7014);
or U9937 (N_9937,N_6560,N_6275);
nor U9938 (N_9938,N_7436,N_5504);
nor U9939 (N_9939,N_6809,N_5191);
nor U9940 (N_9940,N_6898,N_5403);
or U9941 (N_9941,N_5649,N_6258);
nand U9942 (N_9942,N_5692,N_7494);
nor U9943 (N_9943,N_6163,N_5451);
nand U9944 (N_9944,N_6835,N_7120);
or U9945 (N_9945,N_5418,N_6614);
or U9946 (N_9946,N_5232,N_6855);
nand U9947 (N_9947,N_6095,N_7419);
nor U9948 (N_9948,N_6720,N_7173);
or U9949 (N_9949,N_5088,N_6684);
nor U9950 (N_9950,N_5639,N_6649);
nand U9951 (N_9951,N_6042,N_6085);
and U9952 (N_9952,N_5877,N_5502);
nand U9953 (N_9953,N_6303,N_5062);
and U9954 (N_9954,N_5934,N_6521);
or U9955 (N_9955,N_5392,N_5689);
or U9956 (N_9956,N_7025,N_6209);
nand U9957 (N_9957,N_6359,N_5603);
or U9958 (N_9958,N_7221,N_5405);
nand U9959 (N_9959,N_5405,N_6952);
and U9960 (N_9960,N_5046,N_6715);
nand U9961 (N_9961,N_6138,N_7458);
or U9962 (N_9962,N_6240,N_5881);
nand U9963 (N_9963,N_7141,N_5590);
or U9964 (N_9964,N_7440,N_7030);
and U9965 (N_9965,N_6686,N_5364);
nor U9966 (N_9966,N_5917,N_7200);
and U9967 (N_9967,N_5733,N_6901);
nand U9968 (N_9968,N_7351,N_6032);
nor U9969 (N_9969,N_7273,N_5281);
and U9970 (N_9970,N_5545,N_6504);
and U9971 (N_9971,N_6353,N_6249);
or U9972 (N_9972,N_5597,N_5288);
and U9973 (N_9973,N_5796,N_6655);
nand U9974 (N_9974,N_7002,N_6089);
or U9975 (N_9975,N_7496,N_6327);
nor U9976 (N_9976,N_6862,N_5782);
nor U9977 (N_9977,N_5060,N_6470);
or U9978 (N_9978,N_5008,N_6677);
nor U9979 (N_9979,N_5118,N_5399);
or U9980 (N_9980,N_5806,N_6539);
nand U9981 (N_9981,N_7156,N_5116);
or U9982 (N_9982,N_6631,N_5704);
nand U9983 (N_9983,N_6828,N_6565);
nand U9984 (N_9984,N_6852,N_5550);
nand U9985 (N_9985,N_5961,N_6711);
and U9986 (N_9986,N_6490,N_6214);
xnor U9987 (N_9987,N_6463,N_7209);
and U9988 (N_9988,N_6364,N_5361);
nand U9989 (N_9989,N_5366,N_5209);
nand U9990 (N_9990,N_5816,N_6304);
nor U9991 (N_9991,N_5942,N_5406);
or U9992 (N_9992,N_6687,N_6133);
and U9993 (N_9993,N_5732,N_6340);
or U9994 (N_9994,N_6358,N_7373);
nand U9995 (N_9995,N_6505,N_7499);
nand U9996 (N_9996,N_6301,N_5403);
nor U9997 (N_9997,N_7326,N_6463);
or U9998 (N_9998,N_6263,N_5870);
nor U9999 (N_9999,N_5010,N_5827);
nor U10000 (N_10000,N_7899,N_8873);
and U10001 (N_10001,N_9369,N_8905);
nor U10002 (N_10002,N_9256,N_9961);
nand U10003 (N_10003,N_8060,N_8070);
and U10004 (N_10004,N_7807,N_8842);
or U10005 (N_10005,N_8569,N_9592);
nor U10006 (N_10006,N_9910,N_8939);
and U10007 (N_10007,N_8925,N_7783);
and U10008 (N_10008,N_9167,N_8544);
and U10009 (N_10009,N_9549,N_8081);
nor U10010 (N_10010,N_9835,N_9866);
xor U10011 (N_10011,N_9041,N_7794);
and U10012 (N_10012,N_8692,N_8056);
nor U10013 (N_10013,N_8590,N_9242);
nand U10014 (N_10014,N_9813,N_8642);
and U10015 (N_10015,N_9519,N_8741);
or U10016 (N_10016,N_9590,N_8045);
and U10017 (N_10017,N_9679,N_7881);
nand U10018 (N_10018,N_8047,N_8990);
nand U10019 (N_10019,N_7940,N_8687);
or U10020 (N_10020,N_8461,N_7671);
or U10021 (N_10021,N_9080,N_9082);
or U10022 (N_10022,N_9110,N_9526);
nor U10023 (N_10023,N_7878,N_9896);
nand U10024 (N_10024,N_9716,N_7958);
nand U10025 (N_10025,N_9875,N_8287);
xnor U10026 (N_10026,N_7667,N_7957);
or U10027 (N_10027,N_8062,N_8727);
xor U10028 (N_10028,N_8352,N_9950);
and U10029 (N_10029,N_9120,N_8637);
or U10030 (N_10030,N_8885,N_8566);
or U10031 (N_10031,N_7799,N_8484);
or U10032 (N_10032,N_7630,N_8903);
nand U10033 (N_10033,N_8582,N_7866);
and U10034 (N_10034,N_9331,N_9400);
or U10035 (N_10035,N_7681,N_9426);
nand U10036 (N_10036,N_8988,N_8949);
nand U10037 (N_10037,N_7557,N_9686);
nor U10038 (N_10038,N_8516,N_7810);
nand U10039 (N_10039,N_8184,N_8333);
or U10040 (N_10040,N_8346,N_9695);
nor U10041 (N_10041,N_7653,N_7571);
and U10042 (N_10042,N_7622,N_9604);
nand U10043 (N_10043,N_9431,N_8263);
or U10044 (N_10044,N_7549,N_8820);
nand U10045 (N_10045,N_8296,N_8746);
nor U10046 (N_10046,N_9743,N_7923);
or U10047 (N_10047,N_9446,N_9535);
and U10048 (N_10048,N_9539,N_9037);
nor U10049 (N_10049,N_9219,N_8376);
or U10050 (N_10050,N_8470,N_7656);
nor U10051 (N_10051,N_8783,N_8069);
and U10052 (N_10052,N_9885,N_8803);
and U10053 (N_10053,N_8479,N_9720);
or U10054 (N_10054,N_9580,N_9467);
nor U10055 (N_10055,N_9430,N_9291);
or U10056 (N_10056,N_9021,N_8289);
or U10057 (N_10057,N_9261,N_8183);
and U10058 (N_10058,N_8200,N_8380);
nand U10059 (N_10059,N_9315,N_7675);
and U10060 (N_10060,N_7636,N_8799);
nand U10061 (N_10061,N_8193,N_8708);
xor U10062 (N_10062,N_7516,N_8133);
nand U10063 (N_10063,N_9058,N_9469);
nand U10064 (N_10064,N_7813,N_9436);
or U10065 (N_10065,N_8092,N_8171);
nor U10066 (N_10066,N_8162,N_9480);
or U10067 (N_10067,N_8995,N_8365);
and U10068 (N_10068,N_8471,N_9477);
and U10069 (N_10069,N_8866,N_8419);
and U10070 (N_10070,N_8477,N_9935);
nor U10071 (N_10071,N_8954,N_8476);
and U10072 (N_10072,N_8485,N_7949);
and U10073 (N_10073,N_8157,N_9654);
or U10074 (N_10074,N_7598,N_9570);
nor U10075 (N_10075,N_9281,N_8316);
xnor U10076 (N_10076,N_8649,N_8797);
and U10077 (N_10077,N_9218,N_9531);
nor U10078 (N_10078,N_8015,N_8623);
nand U10079 (N_10079,N_8865,N_8153);
nor U10080 (N_10080,N_9673,N_9252);
nand U10081 (N_10081,N_9965,N_9227);
or U10082 (N_10082,N_7779,N_8384);
or U10083 (N_10083,N_8324,N_8176);
and U10084 (N_10084,N_8001,N_8144);
and U10085 (N_10085,N_9664,N_9601);
or U10086 (N_10086,N_7661,N_8932);
and U10087 (N_10087,N_8433,N_9948);
nor U10088 (N_10088,N_8268,N_8007);
or U10089 (N_10089,N_8745,N_8979);
or U10090 (N_10090,N_9070,N_9054);
xor U10091 (N_10091,N_8972,N_9949);
nand U10092 (N_10092,N_7613,N_9192);
nor U10093 (N_10093,N_9957,N_8042);
nor U10094 (N_10094,N_8115,N_7893);
and U10095 (N_10095,N_8055,N_9954);
nand U10096 (N_10096,N_7998,N_8474);
nor U10097 (N_10097,N_9048,N_9378);
xor U10098 (N_10098,N_9404,N_9484);
or U10099 (N_10099,N_8702,N_9370);
and U10100 (N_10100,N_9723,N_9072);
nand U10101 (N_10101,N_8574,N_9698);
and U10102 (N_10102,N_7904,N_9402);
nand U10103 (N_10103,N_8186,N_9650);
or U10104 (N_10104,N_8562,N_9197);
and U10105 (N_10105,N_8864,N_8618);
nand U10106 (N_10106,N_8591,N_9609);
nor U10107 (N_10107,N_8624,N_7619);
or U10108 (N_10108,N_9359,N_7537);
nand U10109 (N_10109,N_7708,N_8772);
or U10110 (N_10110,N_7758,N_8116);
nand U10111 (N_10111,N_8321,N_9019);
nand U10112 (N_10112,N_8858,N_8691);
or U10113 (N_10113,N_7967,N_7637);
nor U10114 (N_10114,N_7872,N_9794);
or U10115 (N_10115,N_7829,N_9657);
nand U10116 (N_10116,N_8067,N_9703);
or U10117 (N_10117,N_8389,N_7574);
nor U10118 (N_10118,N_9619,N_7514);
or U10119 (N_10119,N_8914,N_8585);
or U10120 (N_10120,N_8683,N_8394);
and U10121 (N_10121,N_8499,N_7827);
and U10122 (N_10122,N_7657,N_9976);
nand U10123 (N_10123,N_9702,N_8090);
or U10124 (N_10124,N_9180,N_9500);
and U10125 (N_10125,N_7736,N_9921);
or U10126 (N_10126,N_7662,N_9567);
and U10127 (N_10127,N_7624,N_8284);
and U10128 (N_10128,N_8732,N_9658);
xnor U10129 (N_10129,N_8019,N_7548);
nor U10130 (N_10130,N_7812,N_8840);
or U10131 (N_10131,N_8787,N_9968);
and U10132 (N_10132,N_9809,N_9615);
and U10133 (N_10133,N_7684,N_9052);
nor U10134 (N_10134,N_9128,N_9753);
and U10135 (N_10135,N_8426,N_9827);
and U10136 (N_10136,N_7720,N_7592);
or U10137 (N_10137,N_9582,N_9438);
nand U10138 (N_10138,N_8862,N_9762);
nor U10139 (N_10139,N_9345,N_8944);
xnor U10140 (N_10140,N_7568,N_7570);
or U10141 (N_10141,N_8785,N_9637);
or U10142 (N_10142,N_7788,N_9509);
nor U10143 (N_10143,N_8026,N_9565);
nand U10144 (N_10144,N_8434,N_9283);
nor U10145 (N_10145,N_7566,N_9955);
and U10146 (N_10146,N_8407,N_7601);
or U10147 (N_10147,N_9704,N_9731);
nor U10148 (N_10148,N_9584,N_8868);
nand U10149 (N_10149,N_9280,N_9050);
and U10150 (N_10150,N_7545,N_8826);
or U10151 (N_10151,N_9100,N_8759);
nand U10152 (N_10152,N_7861,N_7824);
nand U10153 (N_10153,N_7884,N_8031);
nor U10154 (N_10154,N_9410,N_8307);
nand U10155 (N_10155,N_8936,N_7976);
and U10156 (N_10156,N_8528,N_9861);
nor U10157 (N_10157,N_8383,N_7818);
nand U10158 (N_10158,N_9394,N_7610);
nand U10159 (N_10159,N_7654,N_8293);
nand U10160 (N_10160,N_7941,N_9734);
or U10161 (N_10161,N_9818,N_9841);
nand U10162 (N_10162,N_9895,N_9848);
and U10163 (N_10163,N_7693,N_8758);
or U10164 (N_10164,N_8613,N_9456);
or U10165 (N_10165,N_9216,N_7769);
xnor U10166 (N_10166,N_9005,N_9936);
or U10167 (N_10167,N_8898,N_8603);
and U10168 (N_10168,N_7859,N_9953);
and U10169 (N_10169,N_7980,N_8039);
or U10170 (N_10170,N_7843,N_9674);
or U10171 (N_10171,N_9867,N_9511);
or U10172 (N_10172,N_9947,N_8472);
or U10173 (N_10173,N_8464,N_9992);
nor U10174 (N_10174,N_8230,N_8154);
nor U10175 (N_10175,N_9544,N_9352);
or U10176 (N_10176,N_9661,N_7648);
and U10177 (N_10177,N_9900,N_7502);
and U10178 (N_10178,N_9271,N_7802);
or U10179 (N_10179,N_9899,N_9836);
nor U10180 (N_10180,N_8754,N_9416);
or U10181 (N_10181,N_8351,N_9497);
or U10182 (N_10182,N_8644,N_8899);
nand U10183 (N_10183,N_9353,N_9297);
nand U10184 (N_10184,N_8549,N_7734);
or U10185 (N_10185,N_8146,N_9783);
and U10186 (N_10186,N_7862,N_8347);
nand U10187 (N_10187,N_9317,N_9304);
nand U10188 (N_10188,N_9611,N_9361);
nand U10189 (N_10189,N_8685,N_7692);
nor U10190 (N_10190,N_9024,N_9721);
nor U10191 (N_10191,N_8705,N_9104);
nand U10192 (N_10192,N_8054,N_8641);
nor U10193 (N_10193,N_9379,N_8238);
and U10194 (N_10194,N_7902,N_7896);
and U10195 (N_10195,N_8833,N_7747);
nor U10196 (N_10196,N_7740,N_8431);
xor U10197 (N_10197,N_7642,N_9202);
or U10198 (N_10198,N_8933,N_9321);
and U10199 (N_10199,N_7558,N_8597);
nand U10200 (N_10200,N_9878,N_7646);
and U10201 (N_10201,N_9824,N_9164);
nand U10202 (N_10202,N_8445,N_7730);
nor U10203 (N_10203,N_9886,N_9845);
nor U10204 (N_10204,N_7728,N_9089);
nand U10205 (N_10205,N_8877,N_8423);
and U10206 (N_10206,N_8052,N_9106);
nand U10207 (N_10207,N_9069,N_7710);
and U10208 (N_10208,N_7678,N_8769);
or U10209 (N_10209,N_8500,N_8298);
nand U10210 (N_10210,N_7915,N_8610);
nand U10211 (N_10211,N_9541,N_8831);
and U10212 (N_10212,N_9022,N_9795);
nand U10213 (N_10213,N_9109,N_8437);
or U10214 (N_10214,N_8232,N_8504);
and U10215 (N_10215,N_9891,N_8374);
or U10216 (N_10216,N_9111,N_8277);
and U10217 (N_10217,N_7525,N_8595);
nor U10218 (N_10218,N_8716,N_7774);
nor U10219 (N_10219,N_7583,N_9183);
or U10220 (N_10220,N_9907,N_8128);
and U10221 (N_10221,N_8968,N_7805);
and U10222 (N_10222,N_8695,N_8598);
nor U10223 (N_10223,N_9691,N_8722);
nand U10224 (N_10224,N_9884,N_7909);
nand U10225 (N_10225,N_8740,N_9985);
nor U10226 (N_10226,N_7889,N_7856);
nand U10227 (N_10227,N_9445,N_7600);
or U10228 (N_10228,N_8962,N_8725);
nor U10229 (N_10229,N_8935,N_9201);
nand U10230 (N_10230,N_9966,N_9578);
nand U10231 (N_10231,N_9632,N_8611);
or U10232 (N_10232,N_9656,N_7739);
nor U10233 (N_10233,N_8486,N_8630);
nor U10234 (N_10234,N_8863,N_7775);
or U10235 (N_10235,N_8207,N_8029);
nand U10236 (N_10236,N_9334,N_8812);
or U10237 (N_10237,N_8571,N_9828);
nor U10238 (N_10238,N_8843,N_8229);
nor U10239 (N_10239,N_8175,N_8838);
nor U10240 (N_10240,N_8095,N_8119);
or U10241 (N_10241,N_8231,N_9787);
and U10242 (N_10242,N_7962,N_8237);
nor U10243 (N_10243,N_9136,N_8032);
xor U10244 (N_10244,N_9335,N_9903);
nand U10245 (N_10245,N_7688,N_8125);
nor U10246 (N_10246,N_8554,N_9406);
and U10247 (N_10247,N_8023,N_9710);
or U10248 (N_10248,N_8660,N_8182);
and U10249 (N_10249,N_8483,N_8650);
nand U10250 (N_10250,N_8264,N_7977);
and U10251 (N_10251,N_8282,N_8557);
nand U10252 (N_10252,N_8847,N_8841);
and U10253 (N_10253,N_7663,N_8635);
and U10254 (N_10254,N_9333,N_8672);
and U10255 (N_10255,N_9168,N_7891);
nand U10256 (N_10256,N_9343,N_9959);
and U10257 (N_10257,N_7596,N_8076);
or U10258 (N_10258,N_7741,N_9066);
nand U10259 (N_10259,N_9020,N_7582);
nor U10260 (N_10260,N_8100,N_8252);
or U10261 (N_10261,N_9407,N_8002);
or U10262 (N_10262,N_9483,N_8892);
nand U10263 (N_10263,N_9159,N_7853);
and U10264 (N_10264,N_9843,N_9073);
xnor U10265 (N_10265,N_7536,N_7551);
nor U10266 (N_10266,N_8460,N_8654);
and U10267 (N_10267,N_8615,N_8663);
nand U10268 (N_10268,N_8037,N_8927);
or U10269 (N_10269,N_9032,N_7969);
or U10270 (N_10270,N_9092,N_7863);
and U10271 (N_10271,N_7978,N_8592);
nor U10272 (N_10272,N_9203,N_9717);
or U10273 (N_10273,N_9858,N_7868);
nor U10274 (N_10274,N_8998,N_9942);
nor U10275 (N_10275,N_9941,N_8542);
nor U10276 (N_10276,N_7695,N_9278);
nor U10277 (N_10277,N_9659,N_9174);
nand U10278 (N_10278,N_9874,N_7763);
nor U10279 (N_10279,N_8911,N_8576);
nor U10280 (N_10280,N_9712,N_8216);
or U10281 (N_10281,N_8290,N_9645);
xor U10282 (N_10282,N_9478,N_8806);
nor U10283 (N_10283,N_8501,N_8401);
and U10284 (N_10284,N_9785,N_8498);
nand U10285 (N_10285,N_7660,N_9629);
or U10286 (N_10286,N_9504,N_9408);
nor U10287 (N_10287,N_8310,N_8294);
nor U10288 (N_10288,N_8386,N_8250);
nor U10289 (N_10289,N_9428,N_8168);
nand U10290 (N_10290,N_9798,N_9696);
or U10291 (N_10291,N_7946,N_8219);
nor U10292 (N_10292,N_9272,N_8077);
nand U10293 (N_10293,N_9690,N_8779);
or U10294 (N_10294,N_8412,N_9806);
or U10295 (N_10295,N_8288,N_9623);
nand U10296 (N_10296,N_7901,N_9228);
and U10297 (N_10297,N_9887,N_7554);
or U10298 (N_10298,N_8607,N_9380);
nand U10299 (N_10299,N_9765,N_9178);
nand U10300 (N_10300,N_8370,N_9507);
nor U10301 (N_10301,N_8675,N_9638);
or U10302 (N_10302,N_9460,N_7761);
nand U10303 (N_10303,N_9241,N_9444);
nor U10304 (N_10304,N_8751,N_8832);
xor U10305 (N_10305,N_9387,N_8867);
and U10306 (N_10306,N_8506,N_7870);
and U10307 (N_10307,N_7576,N_9829);
xnor U10308 (N_10308,N_9781,N_9595);
nor U10309 (N_10309,N_8786,N_8671);
and U10310 (N_10310,N_8940,N_8065);
nor U10311 (N_10311,N_8744,N_9802);
nor U10312 (N_10312,N_7777,N_8837);
nor U10313 (N_10313,N_8427,N_8358);
nor U10314 (N_10314,N_8825,N_8648);
or U10315 (N_10315,N_8969,N_9902);
nand U10316 (N_10316,N_8502,N_8537);
or U10317 (N_10317,N_8142,N_7835);
xor U10318 (N_10318,N_8855,N_8400);
and U10319 (N_10319,N_8548,N_9839);
or U10320 (N_10320,N_8191,N_8391);
xor U10321 (N_10321,N_9700,N_7883);
nor U10322 (N_10322,N_7578,N_7522);
or U10323 (N_10323,N_8947,N_9711);
or U10324 (N_10324,N_8588,N_9501);
nand U10325 (N_10325,N_9103,N_9811);
nand U10326 (N_10326,N_9084,N_9115);
or U10327 (N_10327,N_9047,N_9236);
and U10328 (N_10328,N_7632,N_7874);
nor U10329 (N_10329,N_9646,N_8964);
and U10330 (N_10330,N_8665,N_8093);
and U10331 (N_10331,N_7887,N_9474);
and U10332 (N_10332,N_8539,N_7833);
and U10333 (N_10333,N_7501,N_9760);
nor U10334 (N_10334,N_9685,N_9411);
nand U10335 (N_10335,N_8048,N_9038);
and U10336 (N_10336,N_8719,N_9277);
nand U10337 (N_10337,N_8150,N_8280);
and U10338 (N_10338,N_9926,N_8436);
or U10339 (N_10339,N_8736,N_7756);
nor U10340 (N_10340,N_8586,N_8824);
nand U10341 (N_10341,N_8341,N_7697);
nor U10342 (N_10342,N_8605,N_9081);
or U10343 (N_10343,N_9496,N_9917);
or U10344 (N_10344,N_8469,N_7711);
nor U10345 (N_10345,N_9113,N_7842);
and U10346 (N_10346,N_8385,N_9868);
or U10347 (N_10347,N_9951,N_7793);
or U10348 (N_10348,N_8659,N_8088);
nor U10349 (N_10349,N_9633,N_9791);
nand U10350 (N_10350,N_9130,N_9977);
and U10351 (N_10351,N_8633,N_9425);
nor U10352 (N_10352,N_8078,N_8177);
nor U10353 (N_10353,N_9122,N_8329);
and U10354 (N_10354,N_7649,N_9983);
or U10355 (N_10355,N_8860,N_8983);
nand U10356 (N_10356,N_8733,N_8455);
or U10357 (N_10357,N_8794,N_8068);
nor U10358 (N_10358,N_9090,N_8272);
nand U10359 (N_10359,N_9270,N_9225);
or U10360 (N_10360,N_9099,N_8697);
or U10361 (N_10361,N_7919,N_9736);
or U10362 (N_10362,N_9506,N_7507);
nand U10363 (N_10363,N_9377,N_8169);
nand U10364 (N_10364,N_9616,N_8213);
or U10365 (N_10365,N_9001,N_8894);
nor U10366 (N_10366,N_9076,N_9707);
nand U10367 (N_10367,N_8369,N_9831);
nor U10368 (N_10368,N_8614,N_9775);
or U10369 (N_10369,N_9742,N_7954);
nand U10370 (N_10370,N_7635,N_8050);
or U10371 (N_10371,N_8978,N_9964);
nand U10372 (N_10372,N_9558,N_8814);
and U10373 (N_10373,N_7933,N_9268);
nor U10374 (N_10374,N_9522,N_8756);
or U10375 (N_10375,N_7528,N_8421);
and U10376 (N_10376,N_8451,N_9979);
nand U10377 (N_10377,N_7612,N_8481);
or U10378 (N_10378,N_8710,N_9892);
and U10379 (N_10379,N_7563,N_7994);
nand U10380 (N_10380,N_9316,N_9482);
nand U10381 (N_10381,N_9078,N_7806);
nor U10382 (N_10382,N_7864,N_8425);
nor U10383 (N_10383,N_8625,N_8217);
or U10384 (N_10384,N_8226,N_7744);
and U10385 (N_10385,N_9310,N_8997);
nand U10386 (N_10386,N_9290,N_9341);
or U10387 (N_10387,N_8798,N_7982);
or U10388 (N_10388,N_9919,N_7771);
nand U10389 (N_10389,N_9642,N_7819);
and U10390 (N_10390,N_8538,N_9265);
nand U10391 (N_10391,N_8869,N_9127);
nand U10392 (N_10392,N_9026,N_8127);
nor U10393 (N_10393,N_7615,N_7956);
or U10394 (N_10394,N_8399,N_9034);
nor U10395 (N_10395,N_7588,N_9554);
nor U10396 (N_10396,N_7981,N_8893);
nand U10397 (N_10397,N_9443,N_8490);
nor U10398 (N_10398,N_8339,N_9799);
nor U10399 (N_10399,N_8244,N_8475);
nor U10400 (N_10400,N_9761,N_9059);
and U10401 (N_10401,N_9688,N_8027);
or U10402 (N_10402,N_9018,N_9759);
xor U10403 (N_10403,N_9117,N_9143);
nand U10404 (N_10404,N_8510,N_8694);
nand U10405 (N_10405,N_8243,N_9952);
nor U10406 (N_10406,N_9626,N_9978);
nor U10407 (N_10407,N_8887,N_9160);
nand U10408 (N_10408,N_9330,N_7753);
and U10409 (N_10409,N_8465,N_9651);
and U10410 (N_10410,N_8517,N_9533);
and U10411 (N_10411,N_9245,N_7840);
and U10412 (N_10412,N_7979,N_8724);
nand U10413 (N_10413,N_9226,N_8163);
xnor U10414 (N_10414,N_9705,N_9973);
or U10415 (N_10415,N_8006,N_8105);
or U10416 (N_10416,N_8491,N_7703);
or U10417 (N_10417,N_9514,N_8846);
and U10418 (N_10418,N_7992,N_9249);
or U10419 (N_10419,N_8546,N_9060);
and U10420 (N_10420,N_7855,N_8790);
nand U10421 (N_10421,N_9748,N_9000);
and U10422 (N_10422,N_9741,N_8640);
or U10423 (N_10423,N_7702,N_8955);
nor U10424 (N_10424,N_8676,N_9767);
nand U10425 (N_10425,N_8355,N_7569);
and U10426 (N_10426,N_8752,N_8203);
nor U10427 (N_10427,N_9889,N_9187);
or U10428 (N_10428,N_8620,N_8442);
and U10429 (N_10429,N_8340,N_9630);
nand U10430 (N_10430,N_7729,N_7832);
and U10431 (N_10431,N_9105,N_8432);
nor U10432 (N_10432,N_8197,N_9293);
and U10433 (N_10433,N_9063,N_8878);
nor U10434 (N_10434,N_9348,N_9146);
nor U10435 (N_10435,N_8921,N_8514);
and U10436 (N_10436,N_9162,N_8261);
nor U10437 (N_10437,N_7808,N_7903);
nand U10438 (N_10438,N_8405,N_7964);
or U10439 (N_10439,N_7745,N_9871);
nor U10440 (N_10440,N_7953,N_7694);
and U10441 (N_10441,N_8766,N_8720);
nand U10442 (N_10442,N_7689,N_9096);
and U10443 (N_10443,N_7850,N_9683);
nor U10444 (N_10444,N_7561,N_8767);
nor U10445 (N_10445,N_8242,N_8342);
nor U10446 (N_10446,N_9230,N_9777);
nand U10447 (N_10447,N_8233,N_7605);
xor U10448 (N_10448,N_7625,N_9543);
nor U10449 (N_10449,N_9028,N_8604);
or U10450 (N_10450,N_7531,N_8482);
nand U10451 (N_10451,N_9273,N_9972);
or U10452 (N_10452,N_7905,N_7676);
xnor U10453 (N_10453,N_8503,N_7722);
and U10454 (N_10454,N_8550,N_9569);
or U10455 (N_10455,N_9856,N_8072);
and U10456 (N_10456,N_9184,N_9880);
xor U10457 (N_10457,N_7918,N_9857);
nand U10458 (N_10458,N_8199,N_8526);
and U10459 (N_10459,N_8616,N_8706);
nand U10460 (N_10460,N_8690,N_8136);
nor U10461 (N_10461,N_8570,N_7886);
nor U10462 (N_10462,N_9893,N_9993);
and U10463 (N_10463,N_9385,N_8647);
nand U10464 (N_10464,N_8408,N_9513);
nand U10465 (N_10465,N_7860,N_9374);
or U10466 (N_10466,N_7597,N_9913);
nand U10467 (N_10467,N_9844,N_8757);
and U10468 (N_10468,N_9733,N_7816);
or U10469 (N_10469,N_8025,N_8249);
nand U10470 (N_10470,N_9083,N_8073);
nor U10471 (N_10471,N_9752,N_9098);
nor U10472 (N_10472,N_8034,N_9863);
and U10473 (N_10473,N_8379,N_9327);
or U10474 (N_10474,N_9088,N_8926);
nor U10475 (N_10475,N_8765,N_8446);
or U10476 (N_10476,N_9666,N_8596);
nor U10477 (N_10477,N_9206,N_8403);
or U10478 (N_10478,N_7559,N_9097);
and U10479 (N_10479,N_9172,N_9356);
and U10480 (N_10480,N_8906,N_7926);
nand U10481 (N_10481,N_9873,N_8051);
nor U10482 (N_10482,N_9571,N_9439);
nand U10483 (N_10483,N_9012,N_8278);
or U10484 (N_10484,N_9419,N_9521);
and U10485 (N_10485,N_9986,N_8326);
nor U10486 (N_10486,N_7837,N_8033);
and U10487 (N_10487,N_9555,N_7679);
and U10488 (N_10488,N_9461,N_8300);
nor U10489 (N_10489,N_8132,N_9667);
and U10490 (N_10490,N_8367,N_8668);
or U10491 (N_10491,N_7934,N_9663);
or U10492 (N_10492,N_7611,N_9613);
xor U10493 (N_10493,N_9589,N_9928);
nand U10494 (N_10494,N_7882,N_8495);
nor U10495 (N_10495,N_8830,N_9943);
nand U10496 (N_10496,N_9435,N_8565);
or U10497 (N_10497,N_7963,N_9820);
nor U10498 (N_10498,N_9373,N_7686);
or U10499 (N_10499,N_8581,N_8061);
and U10500 (N_10500,N_9217,N_7527);
and U10501 (N_10501,N_7931,N_9625);
nand U10502 (N_10502,N_8017,N_8084);
or U10503 (N_10503,N_8021,N_9056);
nor U10504 (N_10504,N_9750,N_9170);
nand U10505 (N_10505,N_9568,N_8053);
and U10506 (N_10506,N_8916,N_8958);
or U10507 (N_10507,N_7770,N_9306);
nor U10508 (N_10508,N_7603,N_7606);
and U10509 (N_10509,N_8976,N_8525);
and U10510 (N_10510,N_9129,N_8628);
or U10511 (N_10511,N_8880,N_8821);
nand U10512 (N_10512,N_7985,N_9489);
nand U10513 (N_10513,N_9150,N_9728);
nand U10514 (N_10514,N_9007,N_9528);
or U10515 (N_10515,N_7673,N_7897);
nor U10516 (N_10516,N_8579,N_8147);
and U10517 (N_10517,N_7725,N_7928);
or U10518 (N_10518,N_8188,N_8303);
nand U10519 (N_10519,N_7509,N_9969);
or U10520 (N_10520,N_9468,N_7973);
and U10521 (N_10521,N_7849,N_9823);
nor U10522 (N_10522,N_9602,N_7997);
nor U10523 (N_10523,N_9877,N_8013);
or U10524 (N_10524,N_7555,N_8742);
nand U10525 (N_10525,N_7888,N_8137);
or U10526 (N_10526,N_9518,N_9551);
nand U10527 (N_10527,N_9956,N_7553);
nand U10528 (N_10528,N_7922,N_8908);
or U10529 (N_10529,N_7647,N_9422);
nand U10530 (N_10530,N_9593,N_7965);
or U10531 (N_10531,N_8602,N_7521);
nand U10532 (N_10532,N_7988,N_9847);
nand U10533 (N_10533,N_9939,N_9744);
or U10534 (N_10534,N_7920,N_8228);
or U10535 (N_10535,N_8443,N_8992);
nor U10536 (N_10536,N_8283,N_7595);
nor U10537 (N_10537,N_8802,N_8871);
nand U10538 (N_10538,N_8192,N_9163);
nor U10539 (N_10539,N_9805,N_8975);
nor U10540 (N_10540,N_8295,N_8378);
nand U10541 (N_10541,N_9065,N_9808);
nor U10542 (N_10542,N_7540,N_9881);
nor U10543 (N_10543,N_9437,N_8255);
xnor U10544 (N_10544,N_8493,N_7727);
or U10545 (N_10545,N_9472,N_7532);
nor U10546 (N_10546,N_8234,N_7968);
or U10547 (N_10547,N_9937,N_8223);
or U10548 (N_10548,N_8808,N_7925);
or U10549 (N_10549,N_7674,N_8533);
nor U10550 (N_10550,N_9133,N_8265);
or U10551 (N_10551,N_9235,N_7641);
and U10552 (N_10552,N_8599,N_7572);
and U10553 (N_10553,N_7867,N_8509);
or U10554 (N_10554,N_7672,N_9409);
or U10555 (N_10555,N_9678,N_8559);
nand U10556 (N_10556,N_7724,N_9770);
or U10557 (N_10557,N_8123,N_7974);
or U10558 (N_10558,N_9131,N_9675);
nand U10559 (N_10559,N_7776,N_8478);
or U10560 (N_10560,N_9429,N_8104);
and U10561 (N_10561,N_9279,N_8928);
or U10562 (N_10562,N_7986,N_7828);
or U10563 (N_10563,N_8028,N_8856);
xor U10564 (N_10564,N_9627,N_7587);
and U10565 (N_10565,N_9289,N_9576);
and U10566 (N_10566,N_9605,N_7682);
and U10567 (N_10567,N_8267,N_9427);
nor U10568 (N_10568,N_7508,N_9205);
nand U10569 (N_10569,N_9890,N_9171);
and U10570 (N_10570,N_9655,N_7633);
or U10571 (N_10571,N_8488,N_9358);
nand U10572 (N_10572,N_9464,N_8547);
and U10573 (N_10573,N_9243,N_8308);
or U10574 (N_10574,N_8999,N_9768);
nor U10575 (N_10575,N_9479,N_8913);
nor U10576 (N_10576,N_9137,N_8317);
and U10577 (N_10577,N_9145,N_9516);
and U10578 (N_10578,N_8156,N_9780);
or U10579 (N_10579,N_9036,N_8415);
and U10580 (N_10580,N_7533,N_9448);
or U10581 (N_10581,N_8082,N_9132);
or U10582 (N_10582,N_9883,N_8991);
nand U10583 (N_10583,N_7547,N_8883);
or U10584 (N_10584,N_9152,N_9908);
or U10585 (N_10585,N_8160,N_7778);
xnor U10586 (N_10586,N_9967,N_9864);
nor U10587 (N_10587,N_9124,N_8564);
nor U10588 (N_10588,N_9624,N_8103);
and U10589 (N_10589,N_9190,N_9284);
and U10590 (N_10590,N_9349,N_9534);
or U10591 (N_10591,N_9577,N_7944);
nor U10592 (N_10592,N_8984,N_7942);
and U10593 (N_10593,N_9223,N_7629);
or U10594 (N_10594,N_9390,N_9699);
nand U10595 (N_10595,N_8206,N_8190);
or U10596 (N_10596,N_8518,N_9600);
or U10597 (N_10597,N_8653,N_9126);
and U10598 (N_10598,N_7701,N_9505);
or U10599 (N_10599,N_7950,N_9323);
nand U10600 (N_10600,N_9075,N_8083);
and U10601 (N_10601,N_7580,N_8239);
and U10602 (N_10602,N_8114,N_8235);
or U10603 (N_10603,N_9579,N_9295);
and U10604 (N_10604,N_8696,N_8459);
nand U10605 (N_10605,N_9552,N_9322);
and U10606 (N_10606,N_9442,N_7738);
nand U10607 (N_10607,N_8035,N_8276);
nor U10608 (N_10608,N_9308,N_9094);
and U10609 (N_10609,N_9833,N_9560);
nor U10610 (N_10610,N_8334,N_9267);
nand U10611 (N_10611,N_8536,N_8113);
or U10612 (N_10612,N_9344,N_8730);
or U10613 (N_10613,N_9930,N_8313);
or U10614 (N_10614,N_9713,N_8522);
and U10615 (N_10615,N_8922,N_7766);
nor U10616 (N_10616,N_8381,N_9998);
or U10617 (N_10617,N_8011,N_8977);
or U10618 (N_10618,N_8981,N_8845);
and U10619 (N_10619,N_9988,N_7815);
nand U10620 (N_10620,N_8849,N_8807);
or U10621 (N_10621,N_7809,N_9852);
nand U10622 (N_10622,N_9239,N_8430);
nor U10623 (N_10623,N_7817,N_9294);
nand U10624 (N_10624,N_9726,N_9586);
and U10625 (N_10625,N_9925,N_8049);
nand U10626 (N_10626,N_9876,N_9405);
or U10627 (N_10627,N_8247,N_8145);
nor U10628 (N_10628,N_8452,N_9550);
nand U10629 (N_10629,N_8809,N_8946);
nor U10630 (N_10630,N_8891,N_9357);
nor U10631 (N_10631,N_9347,N_9193);
nand U10632 (N_10632,N_7520,N_8689);
nand U10633 (N_10633,N_9452,N_7911);
nand U10634 (N_10634,N_7538,N_8319);
nand U10635 (N_10635,N_7721,N_8994);
xor U10636 (N_10636,N_7534,N_8768);
and U10637 (N_10637,N_8800,N_9599);
and U10638 (N_10638,N_9566,N_8181);
nand U10639 (N_10639,N_7782,N_9617);
nand U10640 (N_10640,N_8541,N_7898);
or U10641 (N_10641,N_7644,N_9997);
nand U10642 (N_10642,N_8360,N_8884);
and U10643 (N_10643,N_9423,N_8888);
and U10644 (N_10644,N_9398,N_9355);
nand U10645 (N_10645,N_9093,N_7543);
or U10646 (N_10646,N_9292,N_8669);
nand U10647 (N_10647,N_7907,N_8411);
and U10648 (N_10648,N_9285,N_8784);
nand U10649 (N_10649,N_8982,N_9842);
nand U10650 (N_10650,N_9594,N_9234);
and U10651 (N_10651,N_8189,N_7952);
nor U10652 (N_10652,N_7733,N_8652);
nand U10653 (N_10653,N_9363,N_8285);
nand U10654 (N_10654,N_9142,N_9838);
nand U10655 (N_10655,N_8621,N_7759);
or U10656 (N_10656,N_7945,N_8971);
xnor U10657 (N_10657,N_9463,N_9772);
nor U10658 (N_10658,N_9213,N_9782);
and U10659 (N_10659,N_8185,N_8556);
and U10660 (N_10660,N_7614,N_8583);
and U10661 (N_10661,N_7541,N_7983);
xnor U10662 (N_10662,N_7841,N_7519);
and U10663 (N_10663,N_9125,N_9288);
nor U10664 (N_10664,N_8792,N_7785);
and U10665 (N_10665,N_9635,N_8575);
nand U10666 (N_10666,N_8343,N_9662);
nor U10667 (N_10667,N_9821,N_7628);
nor U10668 (N_10668,N_9621,N_8178);
or U10669 (N_10669,N_9804,N_8256);
nor U10670 (N_10670,N_9545,N_8286);
nor U10671 (N_10671,N_9718,N_8980);
nand U10672 (N_10672,N_8662,N_8989);
or U10673 (N_10673,N_7767,N_8704);
nand U10674 (N_10674,N_9102,N_8466);
or U10675 (N_10675,N_9177,N_8224);
nor U10676 (N_10676,N_9682,N_8551);
and U10677 (N_10677,N_8122,N_9546);
or U10678 (N_10678,N_9631,N_8396);
and U10679 (N_10679,N_9392,N_9149);
and U10680 (N_10680,N_7752,N_7512);
nor U10681 (N_10681,N_8532,N_9287);
xnor U10682 (N_10682,N_7894,N_8907);
nand U10683 (N_10683,N_7960,N_8895);
nand U10684 (N_10684,N_8404,N_9557);
nand U10685 (N_10685,N_7652,N_8606);
nand U10686 (N_10686,N_8764,N_8828);
nor U10687 (N_10687,N_9364,N_8422);
or U10688 (N_10688,N_8889,N_9810);
or U10689 (N_10689,N_9714,N_8096);
or U10690 (N_10690,N_9332,N_8251);
or U10691 (N_10691,N_9865,N_9371);
nand U10692 (N_10692,N_9186,N_9139);
or U10693 (N_10693,N_8701,N_8651);
nor U10694 (N_10694,N_7797,N_8441);
or U10695 (N_10695,N_7677,N_7871);
or U10696 (N_10696,N_7826,N_9017);
nor U10697 (N_10697,N_9247,N_8008);
nor U10698 (N_10698,N_8626,N_9027);
xnor U10699 (N_10699,N_8245,N_9040);
nand U10700 (N_10700,N_8473,N_8489);
nor U10701 (N_10701,N_8534,N_8368);
or U10702 (N_10702,N_8910,N_9148);
nand U10703 (N_10703,N_8345,N_8259);
nand U10704 (N_10704,N_9276,N_9975);
or U10705 (N_10705,N_8195,N_8945);
or U10706 (N_10706,N_9540,N_9397);
or U10707 (N_10707,N_9309,N_8805);
nand U10708 (N_10708,N_7659,N_9556);
and U10709 (N_10709,N_7579,N_9553);
and U10710 (N_10710,N_8357,N_9547);
and U10711 (N_10711,N_8129,N_9990);
xor U10712 (N_10712,N_9719,N_9311);
and U10713 (N_10713,N_7550,N_7801);
nor U10714 (N_10714,N_9724,N_9801);
or U10715 (N_10715,N_9157,N_9035);
nor U10716 (N_10716,N_9123,N_8686);
nand U10717 (N_10717,N_9676,N_8515);
nor U10718 (N_10718,N_9612,N_9644);
and U10719 (N_10719,N_7599,N_8253);
and U10720 (N_10720,N_9224,N_8362);
nand U10721 (N_10721,N_9396,N_9850);
nand U10722 (N_10722,N_8492,N_9025);
or U10723 (N_10723,N_9498,N_9086);
nand U10724 (N_10724,N_9807,N_8829);
or U10725 (N_10725,N_8986,N_9194);
nand U10726 (N_10726,N_7971,N_8041);
and U10727 (N_10727,N_8819,N_7552);
and U10728 (N_10728,N_9338,N_9587);
nor U10729 (N_10729,N_8450,N_8822);
and U10730 (N_10730,N_7822,N_8839);
or U10731 (N_10731,N_8463,N_8707);
and U10732 (N_10732,N_8439,N_7539);
nand U10733 (N_10733,N_9610,N_9255);
nor U10734 (N_10734,N_7895,N_8140);
nand U10735 (N_10735,N_8619,N_9421);
nor U10736 (N_10736,N_8130,N_9510);
and U10737 (N_10737,N_8087,N_8688);
or U10738 (N_10738,N_9882,N_7620);
nor U10739 (N_10739,N_9671,N_8760);
nand U10740 (N_10740,N_9179,N_8292);
or U10741 (N_10741,N_8920,N_7865);
or U10742 (N_10742,N_8167,N_8568);
xor U10743 (N_10743,N_7687,N_7921);
nor U10744 (N_10744,N_9314,N_7798);
nor U10745 (N_10745,N_7731,N_8270);
nand U10746 (N_10746,N_8214,N_8134);
and U10747 (N_10747,N_9434,N_9351);
nor U10748 (N_10748,N_9692,N_9495);
or U10749 (N_10749,N_9238,N_7577);
nor U10750 (N_10750,N_8782,N_8117);
or U10751 (N_10751,N_9653,N_8165);
or U10752 (N_10752,N_9068,N_7513);
and U10753 (N_10753,N_8851,N_9825);
nand U10754 (N_10754,N_8101,N_9471);
or U10755 (N_10755,N_8844,N_7890);
nor U10756 (N_10756,N_9771,N_8749);
or U10757 (N_10757,N_7972,N_7995);
xor U10758 (N_10758,N_8257,N_9470);
or U10759 (N_10759,N_9339,N_7726);
or U10760 (N_10760,N_9774,N_9248);
nor U10761 (N_10761,N_9862,N_7831);
nand U10762 (N_10762,N_9044,N_8987);
and U10763 (N_10763,N_9932,N_7504);
and U10764 (N_10764,N_8363,N_8414);
nand U10765 (N_10765,N_7626,N_8447);
or U10766 (N_10766,N_9135,N_9016);
or U10767 (N_10767,N_9386,N_8004);
nand U10768 (N_10768,N_9451,N_9870);
and U10769 (N_10769,N_8311,N_9365);
nand U10770 (N_10770,N_8854,N_9298);
nand U10771 (N_10771,N_7535,N_9963);
nand U10772 (N_10772,N_7664,N_9958);
nand U10773 (N_10773,N_7691,N_8520);
or U10774 (N_10774,N_9286,N_8306);
nand U10775 (N_10775,N_9996,N_7556);
and U10776 (N_10776,N_8770,N_7500);
and U10777 (N_10777,N_8179,N_9971);
and U10778 (N_10778,N_9372,N_7627);
nor U10779 (N_10779,N_8258,N_8859);
or U10780 (N_10780,N_8638,N_8149);
xor U10781 (N_10781,N_7914,N_9901);
nand U10782 (N_10782,N_7631,N_8519);
xnor U10783 (N_10783,N_7735,N_9709);
nand U10784 (N_10784,N_9738,N_9207);
nor U10785 (N_10785,N_9381,N_9313);
nand U10786 (N_10786,N_9927,N_8996);
or U10787 (N_10787,N_9681,N_9181);
nor U10788 (N_10788,N_8438,N_8210);
nand U10789 (N_10789,N_8508,N_8018);
and U10790 (N_10790,N_7515,N_8254);
nor U10791 (N_10791,N_8763,N_8353);
nand U10792 (N_10792,N_8320,N_9250);
nand U10793 (N_10793,N_7839,N_9776);
xnor U10794 (N_10794,N_9934,N_7955);
nand U10795 (N_10795,N_9574,N_8679);
nor U10796 (N_10796,N_8016,N_8553);
nor U10797 (N_10797,N_7526,N_8375);
and U10798 (N_10798,N_9215,N_9008);
and U10799 (N_10799,N_9822,N_9764);
nor U10800 (N_10800,N_8299,N_9134);
nor U10801 (N_10801,N_7939,N_8918);
and U10802 (N_10802,N_7836,N_8139);
nand U10803 (N_10803,N_9237,N_9300);
nand U10804 (N_10804,N_9628,N_8225);
nor U10805 (N_10805,N_7716,N_8950);
and U10806 (N_10806,N_8218,N_9220);
or U10807 (N_10807,N_9779,N_8291);
and U10808 (N_10808,N_8666,N_7795);
nand U10809 (N_10809,N_9354,N_7590);
or U10810 (N_10810,N_8667,N_9537);
nor U10811 (N_10811,N_9529,N_9640);
nor U10812 (N_10812,N_7959,N_7932);
and U10813 (N_10813,N_8952,N_9485);
nand U10814 (N_10814,N_8861,N_8124);
and U10815 (N_10815,N_7709,N_9154);
and U10816 (N_10816,N_9923,N_8071);
nand U10817 (N_10817,N_7706,N_7906);
or U10818 (N_10818,N_8330,N_8205);
and U10819 (N_10819,N_7670,N_8507);
nor U10820 (N_10820,N_9746,N_9984);
nor U10821 (N_10821,N_9729,N_7742);
and U10822 (N_10822,N_8074,N_9391);
nor U10823 (N_10823,N_7573,N_9756);
nand U10824 (N_10824,N_8750,N_9817);
and U10825 (N_10825,N_7792,N_9303);
and U10826 (N_10826,N_8337,N_8513);
or U10827 (N_10827,N_8963,N_7749);
nand U10828 (N_10828,N_8923,N_8970);
nor U10829 (N_10829,N_8236,N_9453);
nand U10830 (N_10830,N_8406,N_8815);
or U10831 (N_10831,N_9418,N_8409);
nor U10832 (N_10832,N_7666,N_9403);
nor U10833 (N_10833,N_8738,N_8540);
or U10834 (N_10834,N_8875,N_9199);
xor U10835 (N_10835,N_8589,N_9591);
nor U10836 (N_10836,N_8726,N_8938);
and U10837 (N_10837,N_9458,N_7908);
nand U10838 (N_10838,N_9503,N_9095);
or U10839 (N_10839,N_8155,N_8572);
nor U10840 (N_10840,N_8126,N_9694);
nand U10841 (N_10841,N_9583,N_7991);
nor U10842 (N_10842,N_9003,N_9014);
nand U10843 (N_10843,N_9433,N_8304);
nor U10844 (N_10844,N_8684,N_9240);
nor U10845 (N_10845,N_8634,N_8530);
or U10846 (N_10846,N_9636,N_8793);
nor U10847 (N_10847,N_8496,N_9981);
xnor U10848 (N_10848,N_9087,N_9140);
nand U10849 (N_10849,N_7690,N_9269);
or U10850 (N_10850,N_7517,N_9166);
nor U10851 (N_10851,N_9641,N_8497);
or U10852 (N_10852,N_8801,N_8646);
nand U10853 (N_10853,N_8366,N_9299);
and U10854 (N_10854,N_8063,N_9257);
nand U10855 (N_10855,N_8917,N_8428);
nor U10856 (N_10856,N_9195,N_9830);
and U10857 (N_10857,N_8747,N_9530);
and U10858 (N_10858,N_7658,N_7854);
or U10859 (N_10859,N_8099,N_9816);
nor U10860 (N_10860,N_9301,N_8731);
and U10861 (N_10861,N_9015,N_9751);
or U10862 (N_10862,N_9597,N_8609);
or U10863 (N_10863,N_9198,N_9318);
nor U10864 (N_10864,N_7943,N_9517);
nor U10865 (N_10865,N_9812,N_9062);
nand U10866 (N_10866,N_9898,N_9608);
and U10867 (N_10867,N_8993,N_8612);
nand U10868 (N_10868,N_9581,N_8656);
nand U10869 (N_10869,N_9011,N_7773);
nand U10870 (N_10870,N_8909,N_9253);
or U10871 (N_10871,N_9417,N_9473);
nor U10872 (N_10872,N_7929,N_8985);
or U10873 (N_10873,N_9039,N_8246);
nand U10874 (N_10874,N_7594,N_9897);
and U10875 (N_10875,N_9840,N_8170);
xnor U10876 (N_10876,N_8166,N_8057);
nor U10877 (N_10877,N_9158,N_8377);
nand U10878 (N_10878,N_9940,N_9745);
nor U10879 (N_10879,N_7562,N_8468);
or U10880 (N_10880,N_8912,N_9031);
or U10881 (N_10881,N_8778,N_8636);
nor U10882 (N_10882,N_8161,N_7790);
nor U10883 (N_10883,N_7609,N_8402);
nand U10884 (N_10884,N_7780,N_9815);
nand U10885 (N_10885,N_8275,N_9010);
nor U10886 (N_10886,N_8965,N_8555);
or U10887 (N_10887,N_9647,N_8135);
and U10888 (N_10888,N_8834,N_8194);
nand U10889 (N_10889,N_9697,N_9176);
nand U10890 (N_10890,N_7645,N_7951);
and U10891 (N_10891,N_8836,N_9793);
or U10892 (N_10892,N_7869,N_8879);
nand U10893 (N_10893,N_9727,N_9212);
and U10894 (N_10894,N_9832,N_7760);
nor U10895 (N_10895,N_8336,N_9415);
xor U10896 (N_10896,N_8020,N_9307);
and U10897 (N_10897,N_8118,N_8111);
nand U10898 (N_10898,N_7746,N_9209);
nand U10899 (N_10899,N_8850,N_9462);
or U10900 (N_10900,N_8444,N_9962);
or U10901 (N_10901,N_8902,N_7544);
or U10902 (N_10902,N_8558,N_7719);
and U10903 (N_10903,N_8674,N_7857);
or U10904 (N_10904,N_7707,N_9114);
nand U10905 (N_10905,N_7947,N_7715);
and U10906 (N_10906,N_7700,N_7751);
xor U10907 (N_10907,N_9715,N_8097);
or U10908 (N_10908,N_7567,N_9693);
nor U10909 (N_10909,N_9320,N_9155);
and U10910 (N_10910,N_8951,N_7873);
nor U10911 (N_10911,N_7602,N_9486);
and U10912 (N_10912,N_9735,N_7565);
or U10913 (N_10913,N_8241,N_8788);
and U10914 (N_10914,N_9393,N_9042);
or U10915 (N_10915,N_7847,N_9607);
or U10916 (N_10916,N_9251,N_8356);
or U10917 (N_10917,N_8372,N_8775);
and U10918 (N_10918,N_9944,N_9057);
nor U10919 (N_10919,N_8222,N_8915);
or U10920 (N_10920,N_8957,N_7772);
nor U10921 (N_10921,N_7916,N_8529);
and U10922 (N_10922,N_7781,N_8545);
and U10923 (N_10923,N_9931,N_7650);
nor U10924 (N_10924,N_9792,N_8721);
nor U10925 (N_10925,N_9222,N_9493);
nor U10926 (N_10926,N_8680,N_9232);
nand U10927 (N_10927,N_9722,N_9029);
nand U10928 (N_10928,N_8457,N_8382);
and U10929 (N_10929,N_9030,N_8804);
or U10930 (N_10930,N_7803,N_7655);
nor U10931 (N_10931,N_8332,N_7912);
nor U10932 (N_10932,N_7564,N_7938);
and U10933 (N_10933,N_8931,N_7917);
nor U10934 (N_10934,N_9689,N_7851);
nand U10935 (N_10935,N_8335,N_8393);
xor U10936 (N_10936,N_7634,N_9946);
and U10937 (N_10937,N_8699,N_7800);
nor U10938 (N_10938,N_8064,N_9382);
nand U10939 (N_10939,N_8453,N_8388);
and U10940 (N_10940,N_9116,N_8973);
nand U10941 (N_10941,N_7984,N_9077);
and U10942 (N_10942,N_9412,N_8323);
nand U10943 (N_10943,N_8302,N_9564);
nand U10944 (N_10944,N_7768,N_8248);
or U10945 (N_10945,N_8577,N_8761);
nor U10946 (N_10946,N_9575,N_9933);
nor U10947 (N_10947,N_9786,N_8813);
or U10948 (N_10948,N_9502,N_8148);
or U10949 (N_10949,N_9614,N_9494);
or U10950 (N_10950,N_9888,N_8870);
nor U10951 (N_10951,N_9573,N_7669);
nor U10952 (N_10952,N_9169,N_8670);
or U10953 (N_10953,N_7989,N_7910);
nor U10954 (N_10954,N_8937,N_9296);
nor U10955 (N_10955,N_7546,N_9185);
or U10956 (N_10956,N_8266,N_9173);
nor U10957 (N_10957,N_8567,N_8003);
nor U10958 (N_10958,N_8771,N_7823);
or U10959 (N_10959,N_9326,N_8458);
and U10960 (N_10960,N_7765,N_9399);
nand U10961 (N_10961,N_9328,N_8348);
nand U10962 (N_10962,N_9523,N_8755);
nand U10963 (N_10963,N_9264,N_9814);
nor U10964 (N_10964,N_8066,N_9912);
and U10965 (N_10965,N_9916,N_7834);
nor U10966 (N_10966,N_8424,N_9362);
nand U10967 (N_10967,N_8657,N_7529);
and U10968 (N_10968,N_7591,N_8312);
and U10969 (N_10969,N_9778,N_8896);
or U10970 (N_10970,N_8271,N_8713);
and U10971 (N_10971,N_8967,N_9049);
nand U10972 (N_10972,N_9023,N_8681);
and U10973 (N_10973,N_8874,N_9055);
nor U10974 (N_10974,N_8344,N_8012);
and U10975 (N_10975,N_9855,N_9071);
or U10976 (N_10976,N_7585,N_9384);
or U10977 (N_10977,N_9046,N_8417);
nand U10978 (N_10978,N_9559,N_7848);
xor U10979 (N_10979,N_8934,N_9366);
nand U10980 (N_10980,N_7970,N_8531);
and U10981 (N_10981,N_8852,N_9383);
or U10982 (N_10982,N_8075,N_9266);
nor U10983 (N_10983,N_9244,N_9639);
nand U10984 (N_10984,N_9989,N_9879);
or U10985 (N_10985,N_7821,N_9603);
and U10986 (N_10986,N_8180,N_8700);
or U10987 (N_10987,N_8505,N_8373);
or U10988 (N_10988,N_8005,N_7743);
or U10989 (N_10989,N_8331,N_8221);
xor U10990 (N_10990,N_7586,N_9784);
and U10991 (N_10991,N_9282,N_8627);
nand U10992 (N_10992,N_8315,N_9708);
and U10993 (N_10993,N_8187,N_9758);
nand U10994 (N_10994,N_8058,N_8024);
nor U10995 (N_10995,N_8857,N_8729);
xor U10996 (N_10996,N_8943,N_9151);
xnor U10997 (N_10997,N_9441,N_8350);
nand U10998 (N_10998,N_7885,N_8527);
nand U10999 (N_10999,N_8279,N_8511);
nand U11000 (N_11000,N_8622,N_8102);
nor U11001 (N_11001,N_8617,N_8735);
nand U11002 (N_11002,N_9665,N_9196);
nor U11003 (N_11003,N_9319,N_7796);
nor U11004 (N_11004,N_8734,N_9945);
nand U11005 (N_11005,N_7503,N_8094);
nand U11006 (N_11006,N_9144,N_8682);
nand U11007 (N_11007,N_9987,N_9914);
nor U11008 (N_11008,N_7523,N_8349);
and U11009 (N_11009,N_7717,N_8274);
and U11010 (N_11010,N_8086,N_9994);
nand U11011 (N_11011,N_7804,N_8448);
nor U11012 (N_11012,N_9620,N_9672);
and U11013 (N_11013,N_9064,N_9211);
nand U11014 (N_11014,N_8924,N_7846);
and U11015 (N_11015,N_7683,N_8948);
and U11016 (N_11016,N_7784,N_7948);
or U11017 (N_11017,N_8748,N_7924);
and U11018 (N_11018,N_8322,N_9074);
xor U11019 (N_11019,N_9466,N_9970);
nor U11020 (N_11020,N_7789,N_8698);
nand U11021 (N_11021,N_7764,N_9789);
and U11022 (N_11022,N_7975,N_9924);
or U11023 (N_11023,N_9853,N_7966);
nand U11024 (N_11024,N_7879,N_8318);
nand U11025 (N_11025,N_9796,N_8410);
nand U11026 (N_11026,N_9210,N_9457);
or U11027 (N_11027,N_9302,N_9803);
nand U11028 (N_11028,N_7999,N_7593);
or U11029 (N_11029,N_7638,N_8776);
or U11030 (N_11030,N_7685,N_9200);
nand U11031 (N_11031,N_9045,N_9091);
nor U11032 (N_11032,N_9138,N_9481);
nor U11033 (N_11033,N_8711,N_8354);
and U11034 (N_11034,N_7900,N_7607);
and U11035 (N_11035,N_8215,N_8301);
or U11036 (N_11036,N_9175,N_8823);
nor U11037 (N_11037,N_9542,N_8131);
and U11038 (N_11038,N_8159,N_8853);
or U11039 (N_11039,N_8314,N_8494);
nor U11040 (N_11040,N_9561,N_8584);
or U11041 (N_11041,N_9401,N_8632);
or U11042 (N_11042,N_7732,N_9067);
or U11043 (N_11043,N_9312,N_8059);
and U11044 (N_11044,N_8942,N_8608);
and U11045 (N_11045,N_9112,N_9108);
and U11046 (N_11046,N_9233,N_8600);
nor U11047 (N_11047,N_9121,N_8795);
nor U11048 (N_11048,N_7542,N_8897);
or U11049 (N_11049,N_8269,N_9490);
or U11050 (N_11050,N_9755,N_8305);
and U11051 (N_11051,N_7518,N_9668);
nor U11052 (N_11052,N_9851,N_9980);
and U11053 (N_11053,N_9450,N_8328);
and U11054 (N_11054,N_9367,N_9596);
or U11055 (N_11055,N_8715,N_7589);
nor U11056 (N_11056,N_9701,N_7787);
nor U11057 (N_11057,N_8196,N_9938);
nor U11058 (N_11058,N_7604,N_9263);
or U11059 (N_11059,N_9447,N_8777);
nand U11060 (N_11060,N_8739,N_8440);
nor U11061 (N_11061,N_8420,N_8643);
nand U11062 (N_11062,N_9182,N_8085);
nand U11063 (N_11063,N_8561,N_9769);
or U11064 (N_11064,N_8462,N_8974);
nand U11065 (N_11065,N_9563,N_8714);
and U11066 (N_11066,N_9797,N_8467);
nand U11067 (N_11067,N_9368,N_8172);
or U11068 (N_11068,N_9634,N_9929);
nor U11069 (N_11069,N_8098,N_8728);
and U11070 (N_11070,N_7621,N_8121);
nor U11071 (N_11071,N_7639,N_8677);
and U11072 (N_11072,N_9849,N_8240);
and U11073 (N_11073,N_9846,N_9455);
nor U11074 (N_11074,N_9432,N_9061);
or U11075 (N_11075,N_8941,N_8881);
or U11076 (N_11076,N_9757,N_7560);
or U11077 (N_11077,N_7930,N_7913);
or U11078 (N_11078,N_9414,N_9660);
nor U11079 (N_11079,N_7880,N_8543);
and U11080 (N_11080,N_9043,N_7640);
or U11081 (N_11081,N_9706,N_9643);
nand U11082 (N_11082,N_7623,N_8789);
nor U11083 (N_11083,N_8361,N_8435);
and U11084 (N_11084,N_8202,N_9395);
nand U11085 (N_11085,N_9459,N_7651);
nor U11086 (N_11086,N_9515,N_9800);
or U11087 (N_11087,N_8281,N_9834);
and U11088 (N_11088,N_9598,N_9336);
nor U11089 (N_11089,N_9922,N_8036);
nand U11090 (N_11090,N_9562,N_8629);
and U11091 (N_11091,N_8212,N_8022);
and U11092 (N_11092,N_9449,N_7786);
and U11093 (N_11093,N_7704,N_9161);
nand U11094 (N_11094,N_7616,N_9476);
nand U11095 (N_11095,N_8297,N_8835);
or U11096 (N_11096,N_8723,N_7643);
nand U11097 (N_11097,N_8587,N_9260);
nor U11098 (N_11098,N_8010,N_8712);
or U11099 (N_11099,N_8593,N_8578);
or U11100 (N_11100,N_9342,N_9652);
nor U11101 (N_11101,N_8521,N_7713);
and U11102 (N_11102,N_9002,N_9773);
nor U11103 (N_11103,N_9413,N_9191);
and U11104 (N_11104,N_8780,N_8208);
nand U11105 (N_11105,N_9982,N_8693);
or U11106 (N_11106,N_9585,N_8774);
nand U11107 (N_11107,N_9325,N_7510);
and U11108 (N_11108,N_9618,N_9229);
nand U11109 (N_11109,N_8174,N_8890);
nand U11110 (N_11110,N_8106,N_8661);
or U11111 (N_11111,N_9754,N_9009);
nand U11112 (N_11112,N_7791,N_9340);
or U11113 (N_11113,N_7877,N_8655);
or U11114 (N_11114,N_9360,N_9826);
xnor U11115 (N_11115,N_8364,N_9763);
nor U11116 (N_11116,N_7838,N_7811);
and U11117 (N_11117,N_9013,N_9004);
nor U11118 (N_11118,N_7844,N_9388);
and U11119 (N_11119,N_8418,N_8956);
nand U11120 (N_11120,N_9214,N_9725);
nor U11121 (N_11121,N_7699,N_8535);
nand U11122 (N_11122,N_8811,N_8594);
nor U11123 (N_11123,N_7755,N_9684);
and U11124 (N_11124,N_8960,N_7825);
nor U11125 (N_11125,N_8152,N_7845);
nand U11126 (N_11126,N_7696,N_8000);
and U11127 (N_11127,N_8392,N_8512);
and U11128 (N_11128,N_8273,N_9491);
nor U11129 (N_11129,N_9337,N_8091);
or U11130 (N_11130,N_8524,N_8211);
and U11131 (N_11131,N_8930,N_8966);
nand U11132 (N_11132,N_9305,N_9420);
nand U11133 (N_11133,N_9749,N_8110);
and U11134 (N_11134,N_7617,N_9141);
and U11135 (N_11135,N_9747,N_8817);
or U11136 (N_11136,N_7506,N_7680);
nor U11137 (N_11137,N_8796,N_7748);
nand U11138 (N_11138,N_8773,N_9991);
nand U11139 (N_11139,N_8848,N_8107);
and U11140 (N_11140,N_8227,N_9730);
or U11141 (N_11141,N_8673,N_7858);
and U11142 (N_11142,N_7737,N_9905);
and U11143 (N_11143,N_9465,N_7927);
nand U11144 (N_11144,N_8718,N_8781);
nand U11145 (N_11145,N_9153,N_8014);
nand U11146 (N_11146,N_9974,N_9147);
or U11147 (N_11147,N_7718,N_9766);
and U11148 (N_11148,N_8818,N_8664);
or U11149 (N_11149,N_8112,N_8709);
nor U11150 (N_11150,N_8413,N_8449);
nor U11151 (N_11151,N_7993,N_8454);
nand U11152 (N_11152,N_8639,N_8743);
nor U11153 (N_11153,N_8044,N_8929);
nand U11154 (N_11154,N_8143,N_9085);
nand U11155 (N_11155,N_9732,N_9538);
and U11156 (N_11156,N_7936,N_7996);
nor U11157 (N_11157,N_8158,N_8038);
or U11158 (N_11158,N_9536,N_9492);
nand U11159 (N_11159,N_9739,N_8080);
nor U11160 (N_11160,N_8390,N_8580);
or U11161 (N_11161,N_9904,N_7668);
and U11162 (N_11162,N_8325,N_7705);
and U11163 (N_11163,N_8262,N_8919);
or U11164 (N_11164,N_9995,N_9532);
and U11165 (N_11165,N_9906,N_9860);
and U11166 (N_11166,N_7575,N_9524);
nand U11167 (N_11167,N_8552,N_8398);
nand U11168 (N_11168,N_9274,N_9006);
or U11169 (N_11169,N_7875,N_9740);
nand U11170 (N_11170,N_9869,N_8030);
or U11171 (N_11171,N_8560,N_8209);
nor U11172 (N_11172,N_9208,N_8961);
or U11173 (N_11173,N_9527,N_8395);
nand U11174 (N_11174,N_8327,N_8737);
nand U11175 (N_11175,N_7530,N_8753);
or U11176 (N_11176,N_8703,N_8810);
nand U11177 (N_11177,N_8631,N_9488);
and U11178 (N_11178,N_9737,N_8886);
or U11179 (N_11179,N_7581,N_9508);
or U11180 (N_11180,N_7714,N_8876);
or U11181 (N_11181,N_9440,N_8173);
nand U11182 (N_11182,N_8220,N_9254);
nand U11183 (N_11183,N_9329,N_9246);
nand U11184 (N_11184,N_8563,N_9350);
and U11185 (N_11185,N_8901,N_8204);
or U11186 (N_11186,N_8151,N_8198);
nor U11187 (N_11187,N_9819,N_8371);
and U11188 (N_11188,N_7876,N_9677);
nand U11189 (N_11189,N_9156,N_9512);
nor U11190 (N_11190,N_8480,N_9118);
and U11191 (N_11191,N_9680,N_7524);
nand U11192 (N_11192,N_7723,N_9687);
and U11193 (N_11193,N_8827,N_7830);
xnor U11194 (N_11194,N_9520,N_8900);
xnor U11195 (N_11195,N_9424,N_8959);
nand U11196 (N_11196,N_7584,N_8164);
and U11197 (N_11197,N_8601,N_9189);
nor U11198 (N_11198,N_9670,N_9918);
nor U11199 (N_11199,N_8872,N_9788);
nand U11200 (N_11200,N_9454,N_9231);
and U11201 (N_11201,N_8046,N_8120);
xor U11202 (N_11202,N_8645,N_9790);
nand U11203 (N_11203,N_9051,N_7852);
and U11204 (N_11204,N_9911,N_8040);
nor U11205 (N_11205,N_9262,N_9204);
or U11206 (N_11206,N_7987,N_7665);
and U11207 (N_11207,N_8487,N_8717);
and U11208 (N_11208,N_9606,N_7762);
nor U11209 (N_11209,N_8953,N_8009);
nand U11210 (N_11210,N_8456,N_9053);
and U11211 (N_11211,N_9622,N_7990);
nand U11212 (N_11212,N_8141,N_8309);
or U11213 (N_11213,N_8573,N_8678);
nor U11214 (N_11214,N_9275,N_9669);
or U11215 (N_11215,N_7618,N_9033);
nor U11216 (N_11216,N_9259,N_9346);
or U11217 (N_11217,N_7820,N_9572);
nor U11218 (N_11218,N_8904,N_9872);
nor U11219 (N_11219,N_7892,N_9475);
nand U11220 (N_11220,N_9119,N_9324);
or U11221 (N_11221,N_9648,N_8523);
nor U11222 (N_11222,N_9258,N_8108);
or U11223 (N_11223,N_8816,N_8882);
or U11224 (N_11224,N_7698,N_9837);
nor U11225 (N_11225,N_8260,N_7511);
or U11226 (N_11226,N_8658,N_8387);
or U11227 (N_11227,N_9487,N_8043);
and U11228 (N_11228,N_8138,N_7754);
and U11229 (N_11229,N_9854,N_8338);
nor U11230 (N_11230,N_7757,N_7505);
or U11231 (N_11231,N_7961,N_9960);
nand U11232 (N_11232,N_9915,N_9375);
or U11233 (N_11233,N_9859,N_7750);
nand U11234 (N_11234,N_8429,N_9499);
and U11235 (N_11235,N_9525,N_9079);
nand U11236 (N_11236,N_8089,N_7937);
nor U11237 (N_11237,N_9165,N_8079);
nand U11238 (N_11238,N_9894,N_9107);
or U11239 (N_11239,N_7608,N_8109);
or U11240 (N_11240,N_9909,N_8359);
nand U11241 (N_11241,N_9548,N_9999);
nand U11242 (N_11242,N_9649,N_9389);
or U11243 (N_11243,N_9188,N_8762);
and U11244 (N_11244,N_8791,N_8201);
or U11245 (N_11245,N_8397,N_9376);
nor U11246 (N_11246,N_7712,N_9221);
nor U11247 (N_11247,N_9588,N_9101);
and U11248 (N_11248,N_7935,N_8416);
nand U11249 (N_11249,N_9920,N_7814);
nand U11250 (N_11250,N_8172,N_8586);
or U11251 (N_11251,N_8517,N_9278);
nand U11252 (N_11252,N_9972,N_8483);
or U11253 (N_11253,N_8391,N_9204);
or U11254 (N_11254,N_9331,N_8597);
nand U11255 (N_11255,N_8783,N_8532);
nor U11256 (N_11256,N_8042,N_8577);
or U11257 (N_11257,N_7612,N_8157);
or U11258 (N_11258,N_7955,N_9343);
or U11259 (N_11259,N_7707,N_7534);
and U11260 (N_11260,N_8984,N_9266);
xnor U11261 (N_11261,N_7923,N_8238);
nor U11262 (N_11262,N_7802,N_9434);
and U11263 (N_11263,N_9396,N_8660);
nand U11264 (N_11264,N_7749,N_9136);
and U11265 (N_11265,N_9619,N_8749);
and U11266 (N_11266,N_9947,N_8950);
xnor U11267 (N_11267,N_9637,N_7980);
nor U11268 (N_11268,N_9376,N_9767);
or U11269 (N_11269,N_8646,N_7503);
nor U11270 (N_11270,N_8292,N_7514);
nand U11271 (N_11271,N_8420,N_7508);
or U11272 (N_11272,N_9900,N_9236);
nand U11273 (N_11273,N_9611,N_8960);
nor U11274 (N_11274,N_8750,N_8115);
nand U11275 (N_11275,N_9145,N_7988);
or U11276 (N_11276,N_8076,N_9333);
nor U11277 (N_11277,N_7742,N_9740);
and U11278 (N_11278,N_7897,N_7555);
or U11279 (N_11279,N_7592,N_8987);
and U11280 (N_11280,N_8098,N_9283);
nand U11281 (N_11281,N_9260,N_9277);
and U11282 (N_11282,N_9722,N_9630);
or U11283 (N_11283,N_9274,N_8817);
nor U11284 (N_11284,N_9859,N_8401);
or U11285 (N_11285,N_8243,N_9056);
and U11286 (N_11286,N_9166,N_7892);
nor U11287 (N_11287,N_8840,N_9449);
nor U11288 (N_11288,N_8510,N_7589);
xor U11289 (N_11289,N_9830,N_9464);
nand U11290 (N_11290,N_7626,N_7876);
and U11291 (N_11291,N_9577,N_9347);
and U11292 (N_11292,N_8744,N_8134);
or U11293 (N_11293,N_9438,N_7987);
or U11294 (N_11294,N_8932,N_9702);
and U11295 (N_11295,N_9537,N_8943);
nand U11296 (N_11296,N_9248,N_7943);
and U11297 (N_11297,N_8891,N_9889);
or U11298 (N_11298,N_7674,N_7734);
and U11299 (N_11299,N_7704,N_7721);
nor U11300 (N_11300,N_9653,N_8793);
nor U11301 (N_11301,N_8012,N_8279);
or U11302 (N_11302,N_8399,N_7668);
or U11303 (N_11303,N_8643,N_8116);
and U11304 (N_11304,N_7960,N_7653);
or U11305 (N_11305,N_7862,N_7796);
and U11306 (N_11306,N_9981,N_7803);
and U11307 (N_11307,N_8336,N_9753);
nor U11308 (N_11308,N_9456,N_8416);
and U11309 (N_11309,N_8936,N_8894);
nor U11310 (N_11310,N_8493,N_8485);
nand U11311 (N_11311,N_8489,N_9719);
nor U11312 (N_11312,N_9418,N_7553);
nor U11313 (N_11313,N_9855,N_9413);
and U11314 (N_11314,N_7910,N_7809);
nor U11315 (N_11315,N_9087,N_8408);
and U11316 (N_11316,N_9061,N_7560);
or U11317 (N_11317,N_7635,N_8887);
nand U11318 (N_11318,N_7930,N_8984);
and U11319 (N_11319,N_8494,N_7784);
or U11320 (N_11320,N_9233,N_7770);
or U11321 (N_11321,N_7889,N_9520);
and U11322 (N_11322,N_8543,N_8330);
and U11323 (N_11323,N_7671,N_7765);
nand U11324 (N_11324,N_8247,N_7962);
and U11325 (N_11325,N_7721,N_9513);
or U11326 (N_11326,N_8110,N_8338);
nor U11327 (N_11327,N_8283,N_7793);
and U11328 (N_11328,N_8451,N_9799);
nand U11329 (N_11329,N_8325,N_9227);
and U11330 (N_11330,N_7946,N_7931);
nor U11331 (N_11331,N_9310,N_8370);
and U11332 (N_11332,N_8585,N_8510);
or U11333 (N_11333,N_7965,N_7663);
and U11334 (N_11334,N_7801,N_8531);
nand U11335 (N_11335,N_9634,N_9500);
nand U11336 (N_11336,N_9162,N_9312);
or U11337 (N_11337,N_9357,N_9666);
nor U11338 (N_11338,N_9213,N_7893);
and U11339 (N_11339,N_9740,N_9535);
nor U11340 (N_11340,N_8249,N_7525);
nand U11341 (N_11341,N_8445,N_7515);
xor U11342 (N_11342,N_7731,N_9008);
nand U11343 (N_11343,N_9167,N_8215);
nand U11344 (N_11344,N_9756,N_9975);
xor U11345 (N_11345,N_8446,N_9641);
nand U11346 (N_11346,N_8560,N_9329);
nor U11347 (N_11347,N_8465,N_9358);
or U11348 (N_11348,N_8472,N_7769);
nor U11349 (N_11349,N_8300,N_8886);
and U11350 (N_11350,N_9885,N_7742);
and U11351 (N_11351,N_9213,N_9941);
nor U11352 (N_11352,N_9864,N_8207);
nand U11353 (N_11353,N_9824,N_7653);
or U11354 (N_11354,N_9780,N_8417);
nor U11355 (N_11355,N_8850,N_8220);
and U11356 (N_11356,N_8739,N_9641);
and U11357 (N_11357,N_7586,N_8680);
or U11358 (N_11358,N_9887,N_7900);
nand U11359 (N_11359,N_9943,N_8013);
or U11360 (N_11360,N_9540,N_9642);
nor U11361 (N_11361,N_7632,N_8571);
and U11362 (N_11362,N_9408,N_8672);
or U11363 (N_11363,N_9933,N_8201);
nand U11364 (N_11364,N_9845,N_8510);
and U11365 (N_11365,N_9639,N_9189);
or U11366 (N_11366,N_8428,N_8574);
and U11367 (N_11367,N_9352,N_9095);
nor U11368 (N_11368,N_9928,N_8498);
nand U11369 (N_11369,N_8463,N_9056);
nand U11370 (N_11370,N_9899,N_8146);
nand U11371 (N_11371,N_9850,N_8466);
or U11372 (N_11372,N_9330,N_8043);
nor U11373 (N_11373,N_8361,N_8487);
nand U11374 (N_11374,N_7501,N_8422);
and U11375 (N_11375,N_7510,N_9684);
nor U11376 (N_11376,N_8731,N_9288);
nand U11377 (N_11377,N_9177,N_9419);
and U11378 (N_11378,N_9473,N_8016);
and U11379 (N_11379,N_9742,N_9819);
nor U11380 (N_11380,N_9064,N_9794);
and U11381 (N_11381,N_9130,N_8850);
nand U11382 (N_11382,N_7515,N_8319);
nand U11383 (N_11383,N_9076,N_9560);
or U11384 (N_11384,N_9158,N_8846);
nor U11385 (N_11385,N_8118,N_9800);
nor U11386 (N_11386,N_8486,N_8316);
or U11387 (N_11387,N_8817,N_8876);
and U11388 (N_11388,N_9318,N_9091);
nor U11389 (N_11389,N_9919,N_9432);
nand U11390 (N_11390,N_7943,N_9127);
and U11391 (N_11391,N_8722,N_8093);
nand U11392 (N_11392,N_7746,N_7558);
or U11393 (N_11393,N_8764,N_9023);
nand U11394 (N_11394,N_9190,N_8753);
or U11395 (N_11395,N_9080,N_9432);
or U11396 (N_11396,N_9727,N_7955);
nor U11397 (N_11397,N_8487,N_7599);
nand U11398 (N_11398,N_7764,N_9394);
nor U11399 (N_11399,N_8384,N_7644);
and U11400 (N_11400,N_8986,N_7900);
nor U11401 (N_11401,N_8010,N_7667);
and U11402 (N_11402,N_8347,N_8668);
nand U11403 (N_11403,N_7722,N_8100);
nand U11404 (N_11404,N_8912,N_8249);
and U11405 (N_11405,N_9933,N_9261);
nand U11406 (N_11406,N_9804,N_9443);
nor U11407 (N_11407,N_8315,N_8284);
nand U11408 (N_11408,N_9305,N_7902);
or U11409 (N_11409,N_9837,N_9613);
nor U11410 (N_11410,N_8830,N_8314);
xnor U11411 (N_11411,N_8028,N_7908);
nand U11412 (N_11412,N_8310,N_9536);
and U11413 (N_11413,N_9609,N_9541);
and U11414 (N_11414,N_8432,N_7888);
nor U11415 (N_11415,N_8406,N_8923);
nor U11416 (N_11416,N_9935,N_7818);
nor U11417 (N_11417,N_8493,N_8981);
and U11418 (N_11418,N_8541,N_8487);
nor U11419 (N_11419,N_9354,N_9184);
or U11420 (N_11420,N_7874,N_8010);
nand U11421 (N_11421,N_8660,N_8786);
nand U11422 (N_11422,N_7573,N_9510);
and U11423 (N_11423,N_9555,N_8133);
and U11424 (N_11424,N_9867,N_9418);
nand U11425 (N_11425,N_8546,N_8216);
nand U11426 (N_11426,N_9919,N_9841);
nor U11427 (N_11427,N_7902,N_8825);
nor U11428 (N_11428,N_9571,N_8231);
and U11429 (N_11429,N_9970,N_9552);
nor U11430 (N_11430,N_8372,N_8362);
nand U11431 (N_11431,N_7805,N_9346);
nor U11432 (N_11432,N_8539,N_9507);
and U11433 (N_11433,N_8026,N_9529);
or U11434 (N_11434,N_7565,N_8458);
nand U11435 (N_11435,N_9327,N_9620);
nor U11436 (N_11436,N_7923,N_9061);
nand U11437 (N_11437,N_7683,N_9487);
and U11438 (N_11438,N_8169,N_8796);
or U11439 (N_11439,N_9892,N_9359);
nor U11440 (N_11440,N_9064,N_7998);
and U11441 (N_11441,N_8270,N_9043);
or U11442 (N_11442,N_8530,N_8237);
and U11443 (N_11443,N_7583,N_9786);
and U11444 (N_11444,N_9599,N_9916);
nand U11445 (N_11445,N_8736,N_8696);
nor U11446 (N_11446,N_9287,N_9554);
nor U11447 (N_11447,N_8439,N_9397);
and U11448 (N_11448,N_7877,N_8797);
nor U11449 (N_11449,N_9847,N_7598);
nor U11450 (N_11450,N_9310,N_9368);
nor U11451 (N_11451,N_7915,N_7626);
nor U11452 (N_11452,N_7935,N_9172);
or U11453 (N_11453,N_7997,N_9518);
or U11454 (N_11454,N_7570,N_9272);
nand U11455 (N_11455,N_9013,N_8376);
or U11456 (N_11456,N_8289,N_7751);
and U11457 (N_11457,N_7629,N_8794);
and U11458 (N_11458,N_8215,N_8261);
or U11459 (N_11459,N_9922,N_7580);
nand U11460 (N_11460,N_8605,N_9272);
nand U11461 (N_11461,N_8876,N_8773);
or U11462 (N_11462,N_8044,N_8527);
or U11463 (N_11463,N_8146,N_7745);
or U11464 (N_11464,N_8896,N_9899);
nor U11465 (N_11465,N_9504,N_9618);
nand U11466 (N_11466,N_7701,N_9139);
xor U11467 (N_11467,N_9201,N_9297);
and U11468 (N_11468,N_8402,N_9409);
or U11469 (N_11469,N_7838,N_7846);
nand U11470 (N_11470,N_9193,N_8192);
nor U11471 (N_11471,N_9721,N_9217);
nand U11472 (N_11472,N_8239,N_8676);
and U11473 (N_11473,N_8368,N_9679);
and U11474 (N_11474,N_9835,N_8516);
and U11475 (N_11475,N_8143,N_9576);
and U11476 (N_11476,N_8157,N_7599);
nand U11477 (N_11477,N_7802,N_9041);
and U11478 (N_11478,N_7744,N_9751);
and U11479 (N_11479,N_9736,N_8653);
nor U11480 (N_11480,N_8211,N_8944);
nor U11481 (N_11481,N_8661,N_8406);
nand U11482 (N_11482,N_9451,N_8082);
nor U11483 (N_11483,N_8372,N_8907);
nand U11484 (N_11484,N_9793,N_9890);
or U11485 (N_11485,N_9819,N_9726);
or U11486 (N_11486,N_9671,N_9290);
or U11487 (N_11487,N_9556,N_8607);
or U11488 (N_11488,N_8944,N_8698);
xnor U11489 (N_11489,N_8340,N_8030);
nand U11490 (N_11490,N_7538,N_8497);
or U11491 (N_11491,N_9416,N_7997);
nand U11492 (N_11492,N_9852,N_8435);
nand U11493 (N_11493,N_8751,N_9331);
nor U11494 (N_11494,N_9402,N_9157);
and U11495 (N_11495,N_8663,N_9875);
nand U11496 (N_11496,N_7551,N_9168);
and U11497 (N_11497,N_8780,N_9786);
nor U11498 (N_11498,N_8367,N_8995);
nand U11499 (N_11499,N_9449,N_9483);
nor U11500 (N_11500,N_9366,N_9569);
and U11501 (N_11501,N_9653,N_9771);
nand U11502 (N_11502,N_8658,N_8032);
nand U11503 (N_11503,N_7679,N_9848);
nor U11504 (N_11504,N_7855,N_9645);
nor U11505 (N_11505,N_7692,N_8612);
or U11506 (N_11506,N_9309,N_8373);
nand U11507 (N_11507,N_8835,N_8325);
or U11508 (N_11508,N_8701,N_7543);
or U11509 (N_11509,N_8496,N_9601);
nand U11510 (N_11510,N_9936,N_9120);
nand U11511 (N_11511,N_7914,N_8501);
or U11512 (N_11512,N_9042,N_9213);
nand U11513 (N_11513,N_8909,N_8621);
nand U11514 (N_11514,N_9733,N_9136);
or U11515 (N_11515,N_9303,N_9594);
and U11516 (N_11516,N_8199,N_9617);
nand U11517 (N_11517,N_8189,N_9492);
nor U11518 (N_11518,N_7654,N_8583);
nand U11519 (N_11519,N_7804,N_8712);
xor U11520 (N_11520,N_9679,N_8933);
or U11521 (N_11521,N_9186,N_9358);
nand U11522 (N_11522,N_7984,N_7648);
nor U11523 (N_11523,N_9658,N_8429);
nand U11524 (N_11524,N_8243,N_8944);
or U11525 (N_11525,N_8617,N_9975);
xnor U11526 (N_11526,N_8696,N_8145);
or U11527 (N_11527,N_7975,N_9149);
and U11528 (N_11528,N_9099,N_9374);
nand U11529 (N_11529,N_9712,N_9154);
nor U11530 (N_11530,N_8085,N_8068);
nor U11531 (N_11531,N_8752,N_9420);
nand U11532 (N_11532,N_9556,N_7712);
nand U11533 (N_11533,N_7650,N_7789);
or U11534 (N_11534,N_8978,N_9142);
or U11535 (N_11535,N_9988,N_7977);
nor U11536 (N_11536,N_7585,N_9571);
nor U11537 (N_11537,N_8470,N_9497);
and U11538 (N_11538,N_9073,N_9472);
and U11539 (N_11539,N_8365,N_7533);
and U11540 (N_11540,N_7745,N_8006);
nor U11541 (N_11541,N_8264,N_7790);
and U11542 (N_11542,N_9217,N_8856);
and U11543 (N_11543,N_8279,N_7629);
nand U11544 (N_11544,N_8866,N_9242);
nor U11545 (N_11545,N_7595,N_8808);
xnor U11546 (N_11546,N_7943,N_7923);
or U11547 (N_11547,N_7945,N_7712);
or U11548 (N_11548,N_7825,N_7561);
xnor U11549 (N_11549,N_9183,N_7808);
nor U11550 (N_11550,N_8862,N_8147);
or U11551 (N_11551,N_9504,N_8934);
nand U11552 (N_11552,N_7829,N_9847);
and U11553 (N_11553,N_7747,N_9961);
nand U11554 (N_11554,N_9864,N_8990);
or U11555 (N_11555,N_8888,N_9415);
nand U11556 (N_11556,N_8275,N_8904);
nand U11557 (N_11557,N_8800,N_9024);
or U11558 (N_11558,N_8611,N_8236);
or U11559 (N_11559,N_8666,N_9851);
or U11560 (N_11560,N_8938,N_7891);
and U11561 (N_11561,N_7742,N_7763);
or U11562 (N_11562,N_8203,N_7762);
and U11563 (N_11563,N_7556,N_8018);
nand U11564 (N_11564,N_7636,N_9891);
nor U11565 (N_11565,N_8505,N_8898);
or U11566 (N_11566,N_8682,N_7853);
and U11567 (N_11567,N_9606,N_9424);
or U11568 (N_11568,N_9020,N_9952);
and U11569 (N_11569,N_8955,N_9774);
nor U11570 (N_11570,N_9283,N_8411);
nor U11571 (N_11571,N_9408,N_9188);
or U11572 (N_11572,N_9059,N_8192);
and U11573 (N_11573,N_9914,N_9216);
nand U11574 (N_11574,N_9422,N_9061);
and U11575 (N_11575,N_9920,N_9316);
or U11576 (N_11576,N_7526,N_7972);
xor U11577 (N_11577,N_9023,N_9460);
or U11578 (N_11578,N_9344,N_9141);
nand U11579 (N_11579,N_8583,N_9883);
nand U11580 (N_11580,N_9477,N_7713);
nor U11581 (N_11581,N_9556,N_8403);
nand U11582 (N_11582,N_8643,N_7683);
or U11583 (N_11583,N_9203,N_7818);
xor U11584 (N_11584,N_8680,N_9718);
nor U11585 (N_11585,N_9680,N_8179);
and U11586 (N_11586,N_8483,N_9787);
and U11587 (N_11587,N_9350,N_9214);
and U11588 (N_11588,N_8566,N_9188);
and U11589 (N_11589,N_8995,N_9137);
or U11590 (N_11590,N_9387,N_7686);
nor U11591 (N_11591,N_8448,N_9506);
or U11592 (N_11592,N_8277,N_9677);
nor U11593 (N_11593,N_8952,N_9683);
or U11594 (N_11594,N_8236,N_9993);
and U11595 (N_11595,N_9477,N_7870);
nor U11596 (N_11596,N_7772,N_8920);
or U11597 (N_11597,N_8225,N_9923);
or U11598 (N_11598,N_7962,N_8866);
or U11599 (N_11599,N_7910,N_9144);
and U11600 (N_11600,N_8656,N_7876);
or U11601 (N_11601,N_7577,N_9126);
or U11602 (N_11602,N_8956,N_8842);
nor U11603 (N_11603,N_7527,N_9434);
and U11604 (N_11604,N_9346,N_8585);
nand U11605 (N_11605,N_9845,N_9288);
nand U11606 (N_11606,N_9728,N_8968);
and U11607 (N_11607,N_7612,N_8066);
and U11608 (N_11608,N_8800,N_7804);
and U11609 (N_11609,N_9122,N_9257);
or U11610 (N_11610,N_8340,N_9871);
and U11611 (N_11611,N_7677,N_8509);
nand U11612 (N_11612,N_8840,N_8047);
nor U11613 (N_11613,N_9988,N_8530);
and U11614 (N_11614,N_9652,N_7725);
and U11615 (N_11615,N_7654,N_8093);
nand U11616 (N_11616,N_7862,N_9366);
or U11617 (N_11617,N_9064,N_8711);
nand U11618 (N_11618,N_8471,N_8912);
nor U11619 (N_11619,N_9406,N_9364);
or U11620 (N_11620,N_8815,N_9125);
nand U11621 (N_11621,N_9353,N_7750);
or U11622 (N_11622,N_9331,N_8839);
nand U11623 (N_11623,N_8932,N_8584);
nand U11624 (N_11624,N_7995,N_9864);
and U11625 (N_11625,N_7792,N_8883);
and U11626 (N_11626,N_9384,N_9723);
nand U11627 (N_11627,N_9971,N_8824);
and U11628 (N_11628,N_8199,N_9162);
nor U11629 (N_11629,N_9151,N_9980);
and U11630 (N_11630,N_9650,N_9534);
nor U11631 (N_11631,N_7569,N_8318);
or U11632 (N_11632,N_9215,N_9944);
or U11633 (N_11633,N_9248,N_7774);
or U11634 (N_11634,N_8697,N_8148);
and U11635 (N_11635,N_7510,N_8974);
nor U11636 (N_11636,N_8899,N_8695);
or U11637 (N_11637,N_9571,N_9236);
nor U11638 (N_11638,N_9491,N_7949);
nor U11639 (N_11639,N_7935,N_8474);
nor U11640 (N_11640,N_8733,N_8997);
and U11641 (N_11641,N_7550,N_9244);
and U11642 (N_11642,N_9429,N_9368);
or U11643 (N_11643,N_8277,N_7867);
nor U11644 (N_11644,N_8113,N_9965);
or U11645 (N_11645,N_8797,N_7847);
and U11646 (N_11646,N_8117,N_8889);
nor U11647 (N_11647,N_8665,N_8460);
and U11648 (N_11648,N_8564,N_9369);
nand U11649 (N_11649,N_9730,N_8765);
or U11650 (N_11650,N_9858,N_8423);
nor U11651 (N_11651,N_8782,N_9920);
or U11652 (N_11652,N_9695,N_8408);
or U11653 (N_11653,N_8693,N_9220);
nor U11654 (N_11654,N_9815,N_8396);
or U11655 (N_11655,N_8454,N_7714);
and U11656 (N_11656,N_9643,N_7679);
nor U11657 (N_11657,N_8728,N_7860);
and U11658 (N_11658,N_7569,N_9458);
nor U11659 (N_11659,N_7808,N_7891);
nor U11660 (N_11660,N_9446,N_8206);
nor U11661 (N_11661,N_7799,N_9083);
nor U11662 (N_11662,N_8847,N_9593);
xor U11663 (N_11663,N_7784,N_9578);
or U11664 (N_11664,N_9378,N_9644);
and U11665 (N_11665,N_7899,N_9869);
or U11666 (N_11666,N_8823,N_7769);
nor U11667 (N_11667,N_9644,N_9182);
and U11668 (N_11668,N_9181,N_7795);
nand U11669 (N_11669,N_8258,N_8983);
nand U11670 (N_11670,N_9765,N_8019);
nand U11671 (N_11671,N_8511,N_9089);
nand U11672 (N_11672,N_9316,N_7533);
nand U11673 (N_11673,N_7961,N_9745);
xnor U11674 (N_11674,N_9502,N_9963);
nand U11675 (N_11675,N_9224,N_8462);
nor U11676 (N_11676,N_9063,N_8598);
nand U11677 (N_11677,N_8468,N_7710);
or U11678 (N_11678,N_8724,N_9975);
nor U11679 (N_11679,N_8931,N_8993);
nand U11680 (N_11680,N_9836,N_7957);
nand U11681 (N_11681,N_8646,N_9015);
and U11682 (N_11682,N_8038,N_9086);
nand U11683 (N_11683,N_8854,N_8190);
and U11684 (N_11684,N_9862,N_9359);
or U11685 (N_11685,N_9013,N_9490);
nand U11686 (N_11686,N_9451,N_7625);
nand U11687 (N_11687,N_8343,N_9035);
nand U11688 (N_11688,N_7973,N_7690);
nand U11689 (N_11689,N_8333,N_7773);
nor U11690 (N_11690,N_8299,N_9375);
and U11691 (N_11691,N_9037,N_9599);
or U11692 (N_11692,N_7528,N_8609);
or U11693 (N_11693,N_9730,N_8519);
nand U11694 (N_11694,N_9574,N_8380);
nor U11695 (N_11695,N_8244,N_9289);
or U11696 (N_11696,N_8740,N_7671);
nand U11697 (N_11697,N_9979,N_9225);
nor U11698 (N_11698,N_9430,N_7906);
and U11699 (N_11699,N_9338,N_7852);
nand U11700 (N_11700,N_9227,N_9187);
or U11701 (N_11701,N_7521,N_7693);
nand U11702 (N_11702,N_8743,N_8415);
nand U11703 (N_11703,N_7842,N_8279);
and U11704 (N_11704,N_7884,N_9371);
or U11705 (N_11705,N_8004,N_8983);
nor U11706 (N_11706,N_9160,N_9754);
and U11707 (N_11707,N_9503,N_8029);
or U11708 (N_11708,N_8284,N_8120);
nor U11709 (N_11709,N_7509,N_8766);
and U11710 (N_11710,N_8544,N_8077);
nor U11711 (N_11711,N_8105,N_7547);
nand U11712 (N_11712,N_8533,N_8050);
or U11713 (N_11713,N_7948,N_9289);
nor U11714 (N_11714,N_8170,N_8231);
nor U11715 (N_11715,N_9824,N_7933);
nand U11716 (N_11716,N_8565,N_9208);
or U11717 (N_11717,N_9757,N_7967);
and U11718 (N_11718,N_8519,N_8999);
or U11719 (N_11719,N_7863,N_8542);
or U11720 (N_11720,N_7631,N_9706);
nand U11721 (N_11721,N_8808,N_9314);
nand U11722 (N_11722,N_7639,N_8158);
nor U11723 (N_11723,N_9099,N_8889);
nor U11724 (N_11724,N_9304,N_7555);
or U11725 (N_11725,N_7712,N_7921);
xor U11726 (N_11726,N_8358,N_7631);
nand U11727 (N_11727,N_7549,N_7893);
or U11728 (N_11728,N_8173,N_8027);
or U11729 (N_11729,N_9646,N_7616);
nand U11730 (N_11730,N_7765,N_9689);
or U11731 (N_11731,N_8778,N_7954);
and U11732 (N_11732,N_8903,N_9225);
or U11733 (N_11733,N_8480,N_7900);
or U11734 (N_11734,N_7587,N_9659);
or U11735 (N_11735,N_9917,N_9557);
nor U11736 (N_11736,N_8208,N_7697);
or U11737 (N_11737,N_9221,N_9564);
or U11738 (N_11738,N_8091,N_7919);
nor U11739 (N_11739,N_8403,N_8645);
or U11740 (N_11740,N_8557,N_8244);
or U11741 (N_11741,N_7709,N_8171);
nor U11742 (N_11742,N_7861,N_7571);
nor U11743 (N_11743,N_9275,N_9926);
nor U11744 (N_11744,N_8158,N_9717);
nor U11745 (N_11745,N_8527,N_9824);
or U11746 (N_11746,N_8416,N_8966);
and U11747 (N_11747,N_7526,N_8672);
and U11748 (N_11748,N_8332,N_9591);
nor U11749 (N_11749,N_8648,N_8197);
nor U11750 (N_11750,N_8720,N_8667);
and U11751 (N_11751,N_8392,N_7993);
and U11752 (N_11752,N_9781,N_8227);
and U11753 (N_11753,N_9892,N_9607);
xnor U11754 (N_11754,N_8241,N_8626);
or U11755 (N_11755,N_7951,N_8231);
nand U11756 (N_11756,N_7843,N_8948);
nor U11757 (N_11757,N_9901,N_8897);
and U11758 (N_11758,N_7693,N_7502);
nand U11759 (N_11759,N_9271,N_8593);
nor U11760 (N_11760,N_8112,N_9024);
nor U11761 (N_11761,N_7510,N_9329);
nor U11762 (N_11762,N_9492,N_8881);
and U11763 (N_11763,N_7521,N_8843);
nor U11764 (N_11764,N_8493,N_8950);
nand U11765 (N_11765,N_8907,N_7667);
and U11766 (N_11766,N_8335,N_8492);
and U11767 (N_11767,N_9150,N_8065);
or U11768 (N_11768,N_8145,N_8566);
nand U11769 (N_11769,N_7510,N_9675);
or U11770 (N_11770,N_9644,N_9353);
and U11771 (N_11771,N_8228,N_9468);
nand U11772 (N_11772,N_8128,N_8390);
nand U11773 (N_11773,N_7678,N_9312);
nor U11774 (N_11774,N_9968,N_7982);
or U11775 (N_11775,N_9915,N_8498);
nor U11776 (N_11776,N_9971,N_9293);
nor U11777 (N_11777,N_7946,N_9442);
or U11778 (N_11778,N_9952,N_9763);
nand U11779 (N_11779,N_7981,N_9351);
and U11780 (N_11780,N_7990,N_7587);
nor U11781 (N_11781,N_9626,N_8738);
nor U11782 (N_11782,N_8375,N_8282);
or U11783 (N_11783,N_9071,N_9216);
or U11784 (N_11784,N_7861,N_7988);
and U11785 (N_11785,N_7763,N_7594);
or U11786 (N_11786,N_8179,N_9014);
nor U11787 (N_11787,N_9733,N_7725);
nand U11788 (N_11788,N_9790,N_9954);
nand U11789 (N_11789,N_8527,N_9601);
and U11790 (N_11790,N_8790,N_9081);
nor U11791 (N_11791,N_7777,N_8928);
nor U11792 (N_11792,N_9122,N_9003);
or U11793 (N_11793,N_7983,N_8789);
nand U11794 (N_11794,N_9819,N_8780);
and U11795 (N_11795,N_8072,N_9308);
nand U11796 (N_11796,N_7761,N_9450);
and U11797 (N_11797,N_9180,N_9847);
or U11798 (N_11798,N_9515,N_7893);
and U11799 (N_11799,N_8664,N_9522);
or U11800 (N_11800,N_8957,N_9519);
nor U11801 (N_11801,N_7562,N_9628);
or U11802 (N_11802,N_7892,N_9428);
or U11803 (N_11803,N_8269,N_9058);
nor U11804 (N_11804,N_8565,N_8789);
or U11805 (N_11805,N_8834,N_7959);
and U11806 (N_11806,N_9132,N_8999);
and U11807 (N_11807,N_8068,N_7957);
nor U11808 (N_11808,N_8632,N_8721);
nand U11809 (N_11809,N_9832,N_9238);
or U11810 (N_11810,N_9314,N_7782);
or U11811 (N_11811,N_9734,N_8156);
nor U11812 (N_11812,N_8015,N_8257);
nor U11813 (N_11813,N_7508,N_9113);
or U11814 (N_11814,N_7989,N_9501);
or U11815 (N_11815,N_9564,N_8920);
nand U11816 (N_11816,N_9560,N_9910);
nand U11817 (N_11817,N_9551,N_8554);
nor U11818 (N_11818,N_8207,N_9598);
nor U11819 (N_11819,N_7678,N_9623);
or U11820 (N_11820,N_7934,N_7607);
or U11821 (N_11821,N_8625,N_9379);
or U11822 (N_11822,N_8803,N_9107);
and U11823 (N_11823,N_8506,N_8023);
and U11824 (N_11824,N_8179,N_9814);
nor U11825 (N_11825,N_8699,N_7582);
nor U11826 (N_11826,N_8264,N_9089);
nor U11827 (N_11827,N_9780,N_7936);
or U11828 (N_11828,N_9532,N_9992);
nand U11829 (N_11829,N_8413,N_7980);
nor U11830 (N_11830,N_9448,N_9490);
and U11831 (N_11831,N_9831,N_7857);
nor U11832 (N_11832,N_8652,N_8547);
or U11833 (N_11833,N_8720,N_8698);
nor U11834 (N_11834,N_7863,N_8116);
or U11835 (N_11835,N_8522,N_7569);
or U11836 (N_11836,N_7996,N_9711);
nor U11837 (N_11837,N_9469,N_9959);
nor U11838 (N_11838,N_8178,N_8133);
nand U11839 (N_11839,N_9652,N_7963);
xor U11840 (N_11840,N_9755,N_8575);
nand U11841 (N_11841,N_9382,N_9100);
and U11842 (N_11842,N_8473,N_8293);
nand U11843 (N_11843,N_9357,N_8970);
nand U11844 (N_11844,N_8198,N_7775);
nor U11845 (N_11845,N_9223,N_9377);
or U11846 (N_11846,N_8118,N_8596);
nand U11847 (N_11847,N_9617,N_9466);
and U11848 (N_11848,N_9011,N_7631);
or U11849 (N_11849,N_9423,N_9610);
nor U11850 (N_11850,N_9787,N_7930);
nand U11851 (N_11851,N_7981,N_8555);
xnor U11852 (N_11852,N_8597,N_9229);
or U11853 (N_11853,N_7568,N_9846);
or U11854 (N_11854,N_7809,N_8315);
nand U11855 (N_11855,N_7910,N_9787);
or U11856 (N_11856,N_7903,N_9803);
nand U11857 (N_11857,N_9420,N_9727);
nor U11858 (N_11858,N_9527,N_7517);
and U11859 (N_11859,N_8762,N_8389);
nand U11860 (N_11860,N_9970,N_8429);
nor U11861 (N_11861,N_8267,N_9908);
nand U11862 (N_11862,N_9673,N_8890);
or U11863 (N_11863,N_8047,N_7641);
nor U11864 (N_11864,N_8601,N_8198);
nand U11865 (N_11865,N_9675,N_9008);
or U11866 (N_11866,N_7866,N_8176);
nor U11867 (N_11867,N_9510,N_8861);
nor U11868 (N_11868,N_7607,N_9083);
or U11869 (N_11869,N_7609,N_7955);
nand U11870 (N_11870,N_8772,N_8792);
or U11871 (N_11871,N_7590,N_8934);
and U11872 (N_11872,N_8511,N_8207);
nor U11873 (N_11873,N_9539,N_8239);
nor U11874 (N_11874,N_9815,N_7772);
nor U11875 (N_11875,N_9345,N_7518);
or U11876 (N_11876,N_7639,N_7675);
nor U11877 (N_11877,N_8228,N_8594);
nor U11878 (N_11878,N_7917,N_8092);
nor U11879 (N_11879,N_9518,N_8267);
nand U11880 (N_11880,N_9898,N_8803);
and U11881 (N_11881,N_7816,N_9106);
or U11882 (N_11882,N_7819,N_8999);
nand U11883 (N_11883,N_8526,N_7655);
nor U11884 (N_11884,N_9324,N_9368);
nor U11885 (N_11885,N_8584,N_7726);
nand U11886 (N_11886,N_8731,N_9380);
or U11887 (N_11887,N_7603,N_8036);
nand U11888 (N_11888,N_8810,N_9602);
and U11889 (N_11889,N_9608,N_8722);
and U11890 (N_11890,N_9523,N_9091);
or U11891 (N_11891,N_7539,N_9146);
nand U11892 (N_11892,N_8422,N_7603);
nor U11893 (N_11893,N_9793,N_8518);
and U11894 (N_11894,N_8481,N_9262);
nand U11895 (N_11895,N_8748,N_9807);
xor U11896 (N_11896,N_8439,N_9721);
and U11897 (N_11897,N_9888,N_7951);
nand U11898 (N_11898,N_9891,N_8707);
nand U11899 (N_11899,N_8291,N_8723);
and U11900 (N_11900,N_8486,N_9182);
nand U11901 (N_11901,N_7944,N_7979);
nor U11902 (N_11902,N_8721,N_9611);
nand U11903 (N_11903,N_9774,N_9239);
or U11904 (N_11904,N_9243,N_9058);
nor U11905 (N_11905,N_7515,N_8021);
nand U11906 (N_11906,N_9481,N_9587);
nand U11907 (N_11907,N_8185,N_8736);
nand U11908 (N_11908,N_7538,N_9367);
nor U11909 (N_11909,N_8232,N_8322);
nand U11910 (N_11910,N_8332,N_8113);
nand U11911 (N_11911,N_8334,N_9553);
nor U11912 (N_11912,N_7881,N_9673);
and U11913 (N_11913,N_7852,N_7534);
or U11914 (N_11914,N_7517,N_9308);
and U11915 (N_11915,N_9818,N_8705);
or U11916 (N_11916,N_7988,N_8715);
or U11917 (N_11917,N_8391,N_7836);
or U11918 (N_11918,N_9338,N_7747);
nand U11919 (N_11919,N_8470,N_7505);
and U11920 (N_11920,N_7714,N_9788);
nor U11921 (N_11921,N_8591,N_9848);
and U11922 (N_11922,N_8741,N_7614);
nor U11923 (N_11923,N_8215,N_9357);
or U11924 (N_11924,N_8159,N_8001);
nand U11925 (N_11925,N_9488,N_9302);
nand U11926 (N_11926,N_9966,N_7977);
nand U11927 (N_11927,N_8959,N_7913);
nand U11928 (N_11928,N_9868,N_8860);
nand U11929 (N_11929,N_7542,N_9760);
nor U11930 (N_11930,N_8599,N_8219);
nor U11931 (N_11931,N_9766,N_9711);
nor U11932 (N_11932,N_7640,N_8244);
nor U11933 (N_11933,N_8748,N_8124);
and U11934 (N_11934,N_9785,N_7553);
nor U11935 (N_11935,N_9964,N_9075);
and U11936 (N_11936,N_7714,N_8198);
nor U11937 (N_11937,N_9536,N_8811);
or U11938 (N_11938,N_9376,N_8007);
nor U11939 (N_11939,N_9740,N_9936);
nor U11940 (N_11940,N_9896,N_8259);
and U11941 (N_11941,N_7579,N_9666);
and U11942 (N_11942,N_8628,N_8954);
nand U11943 (N_11943,N_8859,N_9296);
or U11944 (N_11944,N_9536,N_7731);
and U11945 (N_11945,N_7937,N_9782);
nor U11946 (N_11946,N_8381,N_9107);
nor U11947 (N_11947,N_7606,N_7613);
nand U11948 (N_11948,N_8384,N_9578);
nor U11949 (N_11949,N_7552,N_8127);
nor U11950 (N_11950,N_7519,N_8543);
xnor U11951 (N_11951,N_8291,N_9469);
or U11952 (N_11952,N_7513,N_8369);
or U11953 (N_11953,N_8018,N_8354);
and U11954 (N_11954,N_8202,N_9308);
or U11955 (N_11955,N_7628,N_7784);
xor U11956 (N_11956,N_8249,N_8394);
nor U11957 (N_11957,N_8769,N_8905);
or U11958 (N_11958,N_9292,N_8820);
nor U11959 (N_11959,N_9208,N_8700);
nor U11960 (N_11960,N_8960,N_8261);
nand U11961 (N_11961,N_9790,N_9305);
and U11962 (N_11962,N_8767,N_9826);
or U11963 (N_11963,N_7991,N_8704);
nand U11964 (N_11964,N_9457,N_9190);
nor U11965 (N_11965,N_8356,N_9389);
or U11966 (N_11966,N_9886,N_8541);
and U11967 (N_11967,N_9603,N_7947);
or U11968 (N_11968,N_8599,N_8415);
nor U11969 (N_11969,N_7602,N_8776);
nor U11970 (N_11970,N_9866,N_9989);
nor U11971 (N_11971,N_9382,N_9806);
nor U11972 (N_11972,N_8634,N_7516);
and U11973 (N_11973,N_7942,N_9818);
nand U11974 (N_11974,N_8679,N_9289);
nor U11975 (N_11975,N_7798,N_8746);
xnor U11976 (N_11976,N_8675,N_8747);
or U11977 (N_11977,N_9402,N_7736);
nand U11978 (N_11978,N_8998,N_9099);
nor U11979 (N_11979,N_7672,N_8953);
or U11980 (N_11980,N_9861,N_9748);
nand U11981 (N_11981,N_8544,N_8403);
or U11982 (N_11982,N_9801,N_9508);
or U11983 (N_11983,N_9088,N_9818);
nor U11984 (N_11984,N_8194,N_9357);
or U11985 (N_11985,N_8486,N_9377);
nand U11986 (N_11986,N_8337,N_9600);
or U11987 (N_11987,N_9425,N_8118);
or U11988 (N_11988,N_7537,N_9268);
or U11989 (N_11989,N_8830,N_9014);
nor U11990 (N_11990,N_7652,N_8517);
nand U11991 (N_11991,N_8102,N_7767);
and U11992 (N_11992,N_8780,N_8299);
nand U11993 (N_11993,N_8749,N_8353);
nand U11994 (N_11994,N_9486,N_7964);
and U11995 (N_11995,N_8750,N_8652);
or U11996 (N_11996,N_8898,N_9773);
nor U11997 (N_11997,N_7677,N_8669);
and U11998 (N_11998,N_9522,N_9742);
or U11999 (N_11999,N_7647,N_8629);
or U12000 (N_12000,N_8772,N_8737);
and U12001 (N_12001,N_9319,N_7900);
nand U12002 (N_12002,N_8570,N_8052);
or U12003 (N_12003,N_9981,N_9454);
and U12004 (N_12004,N_8825,N_8582);
nand U12005 (N_12005,N_7692,N_8036);
or U12006 (N_12006,N_8695,N_9382);
or U12007 (N_12007,N_8681,N_7753);
or U12008 (N_12008,N_9506,N_7787);
or U12009 (N_12009,N_7831,N_9913);
and U12010 (N_12010,N_7644,N_9687);
nor U12011 (N_12011,N_8110,N_9831);
nor U12012 (N_12012,N_9217,N_8786);
nand U12013 (N_12013,N_8660,N_8548);
or U12014 (N_12014,N_7683,N_9685);
and U12015 (N_12015,N_7919,N_8179);
or U12016 (N_12016,N_8607,N_7610);
nand U12017 (N_12017,N_9966,N_8550);
nand U12018 (N_12018,N_8782,N_9572);
nor U12019 (N_12019,N_7501,N_9043);
and U12020 (N_12020,N_8720,N_8132);
nand U12021 (N_12021,N_9160,N_8795);
or U12022 (N_12022,N_9332,N_9914);
and U12023 (N_12023,N_8990,N_7520);
nand U12024 (N_12024,N_9969,N_7626);
nor U12025 (N_12025,N_9147,N_9050);
nand U12026 (N_12026,N_8249,N_9719);
nor U12027 (N_12027,N_8370,N_7545);
nor U12028 (N_12028,N_9888,N_9955);
xor U12029 (N_12029,N_7516,N_9770);
nand U12030 (N_12030,N_7649,N_8380);
nand U12031 (N_12031,N_9310,N_7786);
or U12032 (N_12032,N_9746,N_7941);
or U12033 (N_12033,N_7880,N_8504);
or U12034 (N_12034,N_8655,N_8227);
nor U12035 (N_12035,N_8083,N_8978);
nor U12036 (N_12036,N_8559,N_9235);
nand U12037 (N_12037,N_9405,N_8599);
or U12038 (N_12038,N_8294,N_8882);
or U12039 (N_12039,N_8591,N_9724);
or U12040 (N_12040,N_8254,N_7923);
nand U12041 (N_12041,N_9011,N_9473);
nand U12042 (N_12042,N_8714,N_7650);
nor U12043 (N_12043,N_8822,N_9640);
or U12044 (N_12044,N_7842,N_7586);
nor U12045 (N_12045,N_9828,N_8503);
and U12046 (N_12046,N_7613,N_8787);
nand U12047 (N_12047,N_9883,N_9406);
nand U12048 (N_12048,N_9000,N_7704);
nor U12049 (N_12049,N_9156,N_8073);
or U12050 (N_12050,N_9641,N_8275);
xor U12051 (N_12051,N_9850,N_7932);
nor U12052 (N_12052,N_7667,N_8542);
or U12053 (N_12053,N_8489,N_7699);
and U12054 (N_12054,N_9566,N_8695);
and U12055 (N_12055,N_9288,N_9951);
or U12056 (N_12056,N_7717,N_7856);
and U12057 (N_12057,N_8522,N_8707);
xnor U12058 (N_12058,N_9191,N_7750);
nand U12059 (N_12059,N_7611,N_8422);
or U12060 (N_12060,N_9268,N_9389);
xnor U12061 (N_12061,N_8007,N_8814);
or U12062 (N_12062,N_8322,N_9307);
nand U12063 (N_12063,N_7918,N_9142);
or U12064 (N_12064,N_9166,N_8698);
or U12065 (N_12065,N_8237,N_8633);
nand U12066 (N_12066,N_9552,N_9000);
and U12067 (N_12067,N_9032,N_8521);
or U12068 (N_12068,N_9000,N_9538);
or U12069 (N_12069,N_8380,N_8869);
nand U12070 (N_12070,N_8015,N_8322);
nand U12071 (N_12071,N_8727,N_8833);
and U12072 (N_12072,N_7529,N_7783);
nand U12073 (N_12073,N_9040,N_9241);
nor U12074 (N_12074,N_7511,N_8352);
and U12075 (N_12075,N_7977,N_9505);
or U12076 (N_12076,N_8472,N_7740);
nand U12077 (N_12077,N_9000,N_9314);
and U12078 (N_12078,N_8685,N_7693);
nor U12079 (N_12079,N_9988,N_8213);
nor U12080 (N_12080,N_9229,N_7656);
nor U12081 (N_12081,N_9867,N_7562);
and U12082 (N_12082,N_8286,N_8773);
nor U12083 (N_12083,N_7620,N_8569);
or U12084 (N_12084,N_9671,N_8551);
nand U12085 (N_12085,N_8811,N_9527);
and U12086 (N_12086,N_9654,N_8919);
nor U12087 (N_12087,N_9185,N_9657);
and U12088 (N_12088,N_8307,N_7578);
nor U12089 (N_12089,N_8852,N_7523);
or U12090 (N_12090,N_8005,N_8248);
nor U12091 (N_12091,N_9678,N_8276);
nor U12092 (N_12092,N_8589,N_9168);
nor U12093 (N_12093,N_7975,N_8427);
and U12094 (N_12094,N_8459,N_9355);
nor U12095 (N_12095,N_9430,N_9696);
nor U12096 (N_12096,N_8580,N_7597);
nor U12097 (N_12097,N_7523,N_9098);
nor U12098 (N_12098,N_9205,N_7717);
and U12099 (N_12099,N_9085,N_8550);
and U12100 (N_12100,N_7664,N_8991);
or U12101 (N_12101,N_8332,N_9664);
nor U12102 (N_12102,N_9662,N_8861);
nand U12103 (N_12103,N_7625,N_8102);
nand U12104 (N_12104,N_8614,N_7865);
and U12105 (N_12105,N_9125,N_7611);
nand U12106 (N_12106,N_9274,N_9832);
and U12107 (N_12107,N_9609,N_8688);
nand U12108 (N_12108,N_8915,N_9408);
nand U12109 (N_12109,N_8493,N_8540);
or U12110 (N_12110,N_7725,N_9277);
or U12111 (N_12111,N_9759,N_7697);
nand U12112 (N_12112,N_7966,N_8011);
and U12113 (N_12113,N_8321,N_9993);
nor U12114 (N_12114,N_8829,N_7565);
nand U12115 (N_12115,N_9770,N_9744);
nand U12116 (N_12116,N_8852,N_9855);
and U12117 (N_12117,N_9585,N_8168);
or U12118 (N_12118,N_8264,N_8664);
nor U12119 (N_12119,N_9200,N_8642);
nor U12120 (N_12120,N_8712,N_9358);
nor U12121 (N_12121,N_8014,N_8695);
nand U12122 (N_12122,N_7608,N_9103);
nand U12123 (N_12123,N_9627,N_9277);
nand U12124 (N_12124,N_8883,N_9686);
and U12125 (N_12125,N_7811,N_8369);
or U12126 (N_12126,N_7680,N_7801);
and U12127 (N_12127,N_7881,N_9753);
nand U12128 (N_12128,N_9818,N_8635);
and U12129 (N_12129,N_8562,N_9164);
and U12130 (N_12130,N_8100,N_9103);
nand U12131 (N_12131,N_8407,N_7780);
nand U12132 (N_12132,N_9666,N_7832);
nand U12133 (N_12133,N_8504,N_7507);
and U12134 (N_12134,N_9361,N_9373);
or U12135 (N_12135,N_9729,N_7884);
or U12136 (N_12136,N_8372,N_9496);
and U12137 (N_12137,N_8300,N_8192);
and U12138 (N_12138,N_9435,N_8727);
or U12139 (N_12139,N_8708,N_8746);
nand U12140 (N_12140,N_7574,N_9658);
and U12141 (N_12141,N_7699,N_8432);
nand U12142 (N_12142,N_9448,N_7782);
nand U12143 (N_12143,N_9649,N_7747);
or U12144 (N_12144,N_9568,N_8137);
nor U12145 (N_12145,N_7990,N_7693);
nor U12146 (N_12146,N_7945,N_9743);
nor U12147 (N_12147,N_8289,N_9188);
or U12148 (N_12148,N_7634,N_9217);
nor U12149 (N_12149,N_8987,N_7700);
and U12150 (N_12150,N_8287,N_7883);
or U12151 (N_12151,N_8408,N_8748);
nand U12152 (N_12152,N_9898,N_8970);
or U12153 (N_12153,N_9861,N_8260);
xor U12154 (N_12154,N_8387,N_8356);
nand U12155 (N_12155,N_9831,N_9570);
nand U12156 (N_12156,N_7719,N_9827);
or U12157 (N_12157,N_8490,N_8979);
and U12158 (N_12158,N_7949,N_8363);
and U12159 (N_12159,N_9761,N_9321);
nand U12160 (N_12160,N_8483,N_9382);
nand U12161 (N_12161,N_8015,N_9581);
nor U12162 (N_12162,N_9706,N_9027);
nor U12163 (N_12163,N_9768,N_8809);
nand U12164 (N_12164,N_8068,N_9392);
or U12165 (N_12165,N_8990,N_8140);
nor U12166 (N_12166,N_8257,N_8330);
and U12167 (N_12167,N_9829,N_9707);
or U12168 (N_12168,N_9117,N_8449);
nor U12169 (N_12169,N_9064,N_8880);
or U12170 (N_12170,N_8667,N_8071);
and U12171 (N_12171,N_8899,N_9229);
or U12172 (N_12172,N_8792,N_7510);
and U12173 (N_12173,N_8623,N_9492);
nand U12174 (N_12174,N_7794,N_9830);
nor U12175 (N_12175,N_9898,N_9067);
or U12176 (N_12176,N_9346,N_8922);
nand U12177 (N_12177,N_8070,N_8929);
and U12178 (N_12178,N_8162,N_7833);
nor U12179 (N_12179,N_7723,N_7852);
or U12180 (N_12180,N_9932,N_9976);
nor U12181 (N_12181,N_8732,N_9959);
xnor U12182 (N_12182,N_9091,N_7629);
nor U12183 (N_12183,N_8748,N_8950);
nand U12184 (N_12184,N_9296,N_9639);
and U12185 (N_12185,N_8494,N_8920);
or U12186 (N_12186,N_8864,N_9080);
and U12187 (N_12187,N_9868,N_8645);
and U12188 (N_12188,N_8385,N_8965);
nand U12189 (N_12189,N_9836,N_9827);
nand U12190 (N_12190,N_8341,N_9390);
nor U12191 (N_12191,N_8356,N_7969);
or U12192 (N_12192,N_9534,N_8007);
nand U12193 (N_12193,N_9946,N_7976);
or U12194 (N_12194,N_8739,N_7613);
or U12195 (N_12195,N_8477,N_9079);
nand U12196 (N_12196,N_9969,N_7687);
or U12197 (N_12197,N_9102,N_9163);
nor U12198 (N_12198,N_8515,N_8203);
and U12199 (N_12199,N_8621,N_9683);
nor U12200 (N_12200,N_9784,N_8139);
nor U12201 (N_12201,N_8143,N_9113);
and U12202 (N_12202,N_7818,N_9465);
and U12203 (N_12203,N_7900,N_9237);
nand U12204 (N_12204,N_9899,N_8244);
or U12205 (N_12205,N_8995,N_9670);
or U12206 (N_12206,N_9152,N_7715);
nand U12207 (N_12207,N_8604,N_8853);
nand U12208 (N_12208,N_8818,N_8802);
or U12209 (N_12209,N_9804,N_9175);
or U12210 (N_12210,N_9549,N_7629);
or U12211 (N_12211,N_9434,N_8177);
or U12212 (N_12212,N_7938,N_8117);
and U12213 (N_12213,N_8165,N_8343);
or U12214 (N_12214,N_7611,N_8402);
or U12215 (N_12215,N_9002,N_7666);
nand U12216 (N_12216,N_8340,N_9511);
and U12217 (N_12217,N_8592,N_8594);
nor U12218 (N_12218,N_9627,N_8417);
and U12219 (N_12219,N_8596,N_8143);
and U12220 (N_12220,N_9430,N_7961);
xnor U12221 (N_12221,N_7999,N_8479);
or U12222 (N_12222,N_7862,N_7606);
or U12223 (N_12223,N_7959,N_8495);
and U12224 (N_12224,N_9508,N_7546);
nor U12225 (N_12225,N_7917,N_9712);
or U12226 (N_12226,N_8505,N_9873);
or U12227 (N_12227,N_9109,N_7659);
and U12228 (N_12228,N_7991,N_9105);
and U12229 (N_12229,N_8475,N_7739);
or U12230 (N_12230,N_9004,N_9056);
nor U12231 (N_12231,N_9224,N_8800);
nor U12232 (N_12232,N_9002,N_9424);
and U12233 (N_12233,N_8035,N_8667);
nand U12234 (N_12234,N_8559,N_8858);
nand U12235 (N_12235,N_7941,N_9372);
nand U12236 (N_12236,N_7684,N_9274);
nand U12237 (N_12237,N_9509,N_9090);
nor U12238 (N_12238,N_9474,N_7889);
nand U12239 (N_12239,N_8384,N_7968);
or U12240 (N_12240,N_8737,N_8886);
xnor U12241 (N_12241,N_9705,N_8431);
nor U12242 (N_12242,N_8724,N_8209);
nor U12243 (N_12243,N_8753,N_9509);
or U12244 (N_12244,N_9875,N_8822);
nand U12245 (N_12245,N_9117,N_9033);
nand U12246 (N_12246,N_9259,N_9426);
and U12247 (N_12247,N_9407,N_9490);
nand U12248 (N_12248,N_7787,N_8569);
nor U12249 (N_12249,N_7835,N_8749);
and U12250 (N_12250,N_8541,N_8174);
or U12251 (N_12251,N_8299,N_8274);
nor U12252 (N_12252,N_9182,N_9406);
and U12253 (N_12253,N_8208,N_9735);
nor U12254 (N_12254,N_8430,N_7859);
nand U12255 (N_12255,N_8554,N_8726);
nor U12256 (N_12256,N_8451,N_9377);
xnor U12257 (N_12257,N_9134,N_8942);
nand U12258 (N_12258,N_9703,N_7980);
nand U12259 (N_12259,N_8240,N_8105);
or U12260 (N_12260,N_9956,N_8295);
nor U12261 (N_12261,N_8384,N_9672);
nand U12262 (N_12262,N_7697,N_9074);
nor U12263 (N_12263,N_9699,N_9716);
or U12264 (N_12264,N_7541,N_7738);
and U12265 (N_12265,N_9458,N_7945);
or U12266 (N_12266,N_8278,N_8660);
nor U12267 (N_12267,N_8736,N_9514);
and U12268 (N_12268,N_7866,N_9994);
or U12269 (N_12269,N_9173,N_8815);
or U12270 (N_12270,N_9734,N_9687);
nand U12271 (N_12271,N_9603,N_8242);
and U12272 (N_12272,N_9931,N_9639);
nand U12273 (N_12273,N_9562,N_8007);
or U12274 (N_12274,N_8292,N_9905);
or U12275 (N_12275,N_8550,N_9057);
or U12276 (N_12276,N_7532,N_8858);
or U12277 (N_12277,N_9649,N_9957);
and U12278 (N_12278,N_8215,N_9805);
or U12279 (N_12279,N_8011,N_8816);
or U12280 (N_12280,N_7978,N_9322);
nor U12281 (N_12281,N_7636,N_7952);
and U12282 (N_12282,N_9529,N_8644);
or U12283 (N_12283,N_7725,N_8637);
nand U12284 (N_12284,N_9495,N_8784);
and U12285 (N_12285,N_9427,N_9762);
or U12286 (N_12286,N_8824,N_9413);
or U12287 (N_12287,N_9271,N_9668);
or U12288 (N_12288,N_8096,N_8784);
nor U12289 (N_12289,N_8664,N_9619);
nor U12290 (N_12290,N_9733,N_7674);
or U12291 (N_12291,N_8314,N_8339);
or U12292 (N_12292,N_7733,N_9102);
nor U12293 (N_12293,N_9773,N_9592);
or U12294 (N_12294,N_9294,N_9459);
nand U12295 (N_12295,N_9738,N_8287);
and U12296 (N_12296,N_7988,N_8506);
or U12297 (N_12297,N_9989,N_8979);
nand U12298 (N_12298,N_9301,N_8937);
and U12299 (N_12299,N_9830,N_9098);
nand U12300 (N_12300,N_8748,N_9717);
nor U12301 (N_12301,N_8833,N_9296);
and U12302 (N_12302,N_8336,N_9913);
or U12303 (N_12303,N_8162,N_9593);
nand U12304 (N_12304,N_7796,N_8433);
nand U12305 (N_12305,N_8210,N_9991);
nor U12306 (N_12306,N_9466,N_9801);
or U12307 (N_12307,N_9870,N_9284);
or U12308 (N_12308,N_8206,N_8305);
nand U12309 (N_12309,N_7817,N_8999);
or U12310 (N_12310,N_7594,N_7725);
nor U12311 (N_12311,N_8198,N_8744);
nor U12312 (N_12312,N_9740,N_9239);
and U12313 (N_12313,N_7518,N_7797);
or U12314 (N_12314,N_7708,N_9035);
nand U12315 (N_12315,N_8386,N_8690);
nor U12316 (N_12316,N_7989,N_9508);
nor U12317 (N_12317,N_8120,N_7611);
or U12318 (N_12318,N_8233,N_9029);
nand U12319 (N_12319,N_8823,N_9918);
or U12320 (N_12320,N_7806,N_8592);
and U12321 (N_12321,N_8453,N_8114);
and U12322 (N_12322,N_8375,N_7616);
nand U12323 (N_12323,N_9637,N_7617);
nor U12324 (N_12324,N_9501,N_7957);
nand U12325 (N_12325,N_9190,N_8637);
or U12326 (N_12326,N_7787,N_9260);
nor U12327 (N_12327,N_8371,N_9737);
xor U12328 (N_12328,N_8758,N_8971);
nand U12329 (N_12329,N_7979,N_8262);
and U12330 (N_12330,N_8932,N_9739);
and U12331 (N_12331,N_8146,N_9460);
and U12332 (N_12332,N_9333,N_9466);
nor U12333 (N_12333,N_8085,N_8631);
and U12334 (N_12334,N_9466,N_8544);
and U12335 (N_12335,N_8430,N_9388);
or U12336 (N_12336,N_9969,N_7945);
xor U12337 (N_12337,N_8813,N_8281);
or U12338 (N_12338,N_9265,N_8529);
nand U12339 (N_12339,N_8160,N_8641);
or U12340 (N_12340,N_7686,N_9213);
nand U12341 (N_12341,N_8951,N_9882);
nand U12342 (N_12342,N_7833,N_9865);
or U12343 (N_12343,N_9343,N_9321);
nand U12344 (N_12344,N_8960,N_8410);
or U12345 (N_12345,N_9045,N_9635);
or U12346 (N_12346,N_8417,N_9369);
nor U12347 (N_12347,N_7678,N_8318);
and U12348 (N_12348,N_7948,N_8369);
nand U12349 (N_12349,N_8294,N_9183);
or U12350 (N_12350,N_9296,N_9585);
and U12351 (N_12351,N_9265,N_7933);
nor U12352 (N_12352,N_9375,N_7860);
nand U12353 (N_12353,N_9555,N_8915);
nand U12354 (N_12354,N_8362,N_8804);
or U12355 (N_12355,N_9123,N_8847);
and U12356 (N_12356,N_9050,N_8762);
or U12357 (N_12357,N_9553,N_7607);
nor U12358 (N_12358,N_9775,N_9312);
and U12359 (N_12359,N_7556,N_7833);
and U12360 (N_12360,N_8746,N_9910);
nor U12361 (N_12361,N_8735,N_7655);
and U12362 (N_12362,N_9057,N_8868);
or U12363 (N_12363,N_9104,N_9864);
and U12364 (N_12364,N_7647,N_9081);
nor U12365 (N_12365,N_8361,N_9771);
nor U12366 (N_12366,N_9920,N_8728);
and U12367 (N_12367,N_7829,N_9994);
nand U12368 (N_12368,N_8618,N_8334);
or U12369 (N_12369,N_9240,N_9641);
or U12370 (N_12370,N_8813,N_7934);
nor U12371 (N_12371,N_9237,N_8350);
nand U12372 (N_12372,N_8382,N_9942);
nand U12373 (N_12373,N_9848,N_9275);
or U12374 (N_12374,N_8967,N_9643);
or U12375 (N_12375,N_8160,N_9492);
nor U12376 (N_12376,N_8568,N_8845);
and U12377 (N_12377,N_8740,N_8598);
nand U12378 (N_12378,N_8624,N_9701);
and U12379 (N_12379,N_8531,N_7961);
nand U12380 (N_12380,N_9931,N_8791);
and U12381 (N_12381,N_8403,N_9489);
nand U12382 (N_12382,N_9060,N_8809);
xor U12383 (N_12383,N_8746,N_8884);
nor U12384 (N_12384,N_8182,N_9616);
xor U12385 (N_12385,N_9616,N_8322);
and U12386 (N_12386,N_8260,N_8058);
or U12387 (N_12387,N_7589,N_8048);
nand U12388 (N_12388,N_9424,N_9469);
nand U12389 (N_12389,N_9948,N_8567);
nand U12390 (N_12390,N_9019,N_8423);
nor U12391 (N_12391,N_9935,N_8654);
or U12392 (N_12392,N_9720,N_7924);
nand U12393 (N_12393,N_9364,N_8038);
nand U12394 (N_12394,N_8208,N_7651);
or U12395 (N_12395,N_7794,N_9263);
and U12396 (N_12396,N_7595,N_9592);
and U12397 (N_12397,N_8077,N_9000);
nor U12398 (N_12398,N_9890,N_8756);
nand U12399 (N_12399,N_9931,N_8544);
or U12400 (N_12400,N_8986,N_7720);
nor U12401 (N_12401,N_8993,N_7908);
nor U12402 (N_12402,N_9785,N_8016);
or U12403 (N_12403,N_9597,N_8996);
nand U12404 (N_12404,N_9102,N_9820);
or U12405 (N_12405,N_9557,N_8369);
nand U12406 (N_12406,N_9881,N_8060);
nand U12407 (N_12407,N_9926,N_9431);
and U12408 (N_12408,N_8180,N_9995);
or U12409 (N_12409,N_9070,N_9068);
xor U12410 (N_12410,N_9316,N_8782);
nor U12411 (N_12411,N_8810,N_9980);
or U12412 (N_12412,N_9874,N_9895);
nor U12413 (N_12413,N_7976,N_9722);
and U12414 (N_12414,N_8582,N_9587);
nor U12415 (N_12415,N_9592,N_9406);
nand U12416 (N_12416,N_7950,N_8493);
or U12417 (N_12417,N_9073,N_9572);
or U12418 (N_12418,N_8105,N_9615);
nor U12419 (N_12419,N_8864,N_9682);
and U12420 (N_12420,N_8139,N_9094);
or U12421 (N_12421,N_8092,N_8512);
or U12422 (N_12422,N_9377,N_9413);
and U12423 (N_12423,N_9370,N_9222);
and U12424 (N_12424,N_9604,N_8153);
or U12425 (N_12425,N_9191,N_9162);
nand U12426 (N_12426,N_7919,N_9495);
or U12427 (N_12427,N_9377,N_9503);
nand U12428 (N_12428,N_8228,N_9050);
nand U12429 (N_12429,N_8472,N_8208);
nand U12430 (N_12430,N_7613,N_8688);
and U12431 (N_12431,N_8845,N_8876);
nand U12432 (N_12432,N_8004,N_9118);
and U12433 (N_12433,N_8362,N_9342);
nor U12434 (N_12434,N_9360,N_9076);
and U12435 (N_12435,N_8560,N_8630);
nand U12436 (N_12436,N_8416,N_7943);
nor U12437 (N_12437,N_7716,N_9313);
nor U12438 (N_12438,N_7915,N_8854);
and U12439 (N_12439,N_8505,N_7767);
nand U12440 (N_12440,N_8734,N_9861);
nand U12441 (N_12441,N_9063,N_7901);
nand U12442 (N_12442,N_7501,N_8629);
or U12443 (N_12443,N_9981,N_8738);
and U12444 (N_12444,N_9348,N_7814);
nor U12445 (N_12445,N_7717,N_8632);
nand U12446 (N_12446,N_9521,N_8173);
nand U12447 (N_12447,N_9460,N_8522);
and U12448 (N_12448,N_8497,N_9935);
and U12449 (N_12449,N_8632,N_9712);
nand U12450 (N_12450,N_8371,N_8325);
nor U12451 (N_12451,N_8878,N_7673);
nand U12452 (N_12452,N_7541,N_9976);
or U12453 (N_12453,N_9970,N_9807);
nand U12454 (N_12454,N_9589,N_7982);
nand U12455 (N_12455,N_7545,N_9811);
and U12456 (N_12456,N_9000,N_7877);
and U12457 (N_12457,N_8807,N_9496);
nor U12458 (N_12458,N_7522,N_7677);
nor U12459 (N_12459,N_7755,N_9218);
nor U12460 (N_12460,N_8787,N_8612);
or U12461 (N_12461,N_8916,N_9890);
nand U12462 (N_12462,N_8847,N_8162);
or U12463 (N_12463,N_9747,N_7815);
nor U12464 (N_12464,N_9498,N_9462);
nand U12465 (N_12465,N_7630,N_9979);
and U12466 (N_12466,N_8986,N_8052);
or U12467 (N_12467,N_8467,N_9577);
and U12468 (N_12468,N_9395,N_8861);
xor U12469 (N_12469,N_7796,N_9633);
nand U12470 (N_12470,N_9536,N_8339);
and U12471 (N_12471,N_9867,N_8646);
and U12472 (N_12472,N_8425,N_7845);
or U12473 (N_12473,N_9153,N_8801);
or U12474 (N_12474,N_8303,N_9159);
nor U12475 (N_12475,N_9369,N_8801);
and U12476 (N_12476,N_8085,N_8755);
and U12477 (N_12477,N_9765,N_7831);
nor U12478 (N_12478,N_8059,N_7538);
and U12479 (N_12479,N_9951,N_9779);
and U12480 (N_12480,N_9504,N_8562);
nand U12481 (N_12481,N_9723,N_8974);
or U12482 (N_12482,N_8890,N_7949);
or U12483 (N_12483,N_8124,N_8477);
or U12484 (N_12484,N_8700,N_9420);
nand U12485 (N_12485,N_7893,N_8796);
nor U12486 (N_12486,N_8638,N_7840);
nor U12487 (N_12487,N_9976,N_9284);
nor U12488 (N_12488,N_8879,N_7874);
or U12489 (N_12489,N_8939,N_8888);
or U12490 (N_12490,N_9060,N_8907);
nor U12491 (N_12491,N_7761,N_8863);
nor U12492 (N_12492,N_8335,N_7909);
and U12493 (N_12493,N_8545,N_8626);
and U12494 (N_12494,N_8893,N_9966);
or U12495 (N_12495,N_9103,N_9324);
and U12496 (N_12496,N_8189,N_8724);
or U12497 (N_12497,N_8953,N_9248);
nand U12498 (N_12498,N_9557,N_8633);
nand U12499 (N_12499,N_7643,N_8652);
and U12500 (N_12500,N_12185,N_10258);
xor U12501 (N_12501,N_11298,N_11997);
or U12502 (N_12502,N_11552,N_11393);
nand U12503 (N_12503,N_12218,N_12256);
and U12504 (N_12504,N_11284,N_11472);
or U12505 (N_12505,N_12364,N_10216);
and U12506 (N_12506,N_12208,N_11300);
nor U12507 (N_12507,N_11959,N_10481);
or U12508 (N_12508,N_12342,N_11317);
nand U12509 (N_12509,N_10732,N_11275);
nor U12510 (N_12510,N_10426,N_12387);
nand U12511 (N_12511,N_12421,N_11404);
nor U12512 (N_12512,N_12009,N_10658);
nor U12513 (N_12513,N_11412,N_10846);
nor U12514 (N_12514,N_12236,N_11487);
nor U12515 (N_12515,N_10986,N_11790);
or U12516 (N_12516,N_12003,N_11615);
or U12517 (N_12517,N_11338,N_12044);
or U12518 (N_12518,N_11476,N_10757);
xnor U12519 (N_12519,N_12148,N_11316);
nand U12520 (N_12520,N_11577,N_12186);
and U12521 (N_12521,N_11813,N_11930);
and U12522 (N_12522,N_11799,N_10381);
nand U12523 (N_12523,N_12058,N_11427);
or U12524 (N_12524,N_11851,N_10447);
nand U12525 (N_12525,N_10365,N_12425);
or U12526 (N_12526,N_11217,N_10073);
nor U12527 (N_12527,N_10994,N_10434);
nor U12528 (N_12528,N_11486,N_12022);
nand U12529 (N_12529,N_10615,N_10504);
nor U12530 (N_12530,N_12118,N_12210);
nand U12531 (N_12531,N_10245,N_12238);
or U12532 (N_12532,N_10972,N_11146);
and U12533 (N_12533,N_10089,N_10514);
nand U12534 (N_12534,N_11594,N_11961);
or U12535 (N_12535,N_11802,N_11902);
and U12536 (N_12536,N_11387,N_10847);
and U12537 (N_12537,N_12362,N_10928);
nand U12538 (N_12538,N_12468,N_12294);
nand U12539 (N_12539,N_10257,N_10588);
nor U12540 (N_12540,N_11038,N_11304);
and U12541 (N_12541,N_11776,N_10040);
nand U12542 (N_12542,N_12126,N_11385);
or U12543 (N_12543,N_11163,N_10916);
nand U12544 (N_12544,N_11970,N_11682);
nand U12545 (N_12545,N_11992,N_10571);
or U12546 (N_12546,N_12403,N_12202);
and U12547 (N_12547,N_10085,N_12442);
nor U12548 (N_12548,N_11290,N_11332);
or U12549 (N_12549,N_10611,N_10801);
nand U12550 (N_12550,N_12190,N_12056);
or U12551 (N_12551,N_10389,N_10851);
nor U12552 (N_12552,N_11077,N_11863);
or U12553 (N_12553,N_10876,N_11017);
nor U12554 (N_12554,N_10348,N_11506);
or U12555 (N_12555,N_10749,N_11870);
and U12556 (N_12556,N_12462,N_10445);
and U12557 (N_12557,N_10619,N_10448);
xor U12558 (N_12558,N_11123,N_11478);
and U12559 (N_12559,N_10285,N_12015);
nor U12560 (N_12560,N_11706,N_11988);
nand U12561 (N_12561,N_11451,N_11494);
or U12562 (N_12562,N_10537,N_10711);
or U12563 (N_12563,N_10122,N_11314);
or U12564 (N_12564,N_11777,N_10050);
or U12565 (N_12565,N_10901,N_10460);
and U12566 (N_12566,N_11531,N_11360);
and U12567 (N_12567,N_11571,N_11532);
and U12568 (N_12568,N_10189,N_11648);
or U12569 (N_12569,N_12378,N_11735);
or U12570 (N_12570,N_12483,N_11783);
nor U12571 (N_12571,N_11471,N_10344);
nor U12572 (N_12572,N_12215,N_11892);
or U12573 (N_12573,N_10263,N_11117);
xor U12574 (N_12574,N_10693,N_11252);
nor U12575 (N_12575,N_12252,N_10311);
and U12576 (N_12576,N_10559,N_10246);
nor U12577 (N_12577,N_12465,N_10684);
nor U12578 (N_12578,N_11358,N_10510);
xor U12579 (N_12579,N_12078,N_12101);
or U12580 (N_12580,N_10715,N_11820);
nand U12581 (N_12581,N_11042,N_11812);
or U12582 (N_12582,N_11006,N_10854);
and U12583 (N_12583,N_11606,N_10168);
nand U12584 (N_12584,N_11946,N_11580);
nand U12585 (N_12585,N_11460,N_10133);
nand U12586 (N_12586,N_10443,N_11294);
or U12587 (N_12587,N_10024,N_10587);
and U12588 (N_12588,N_10591,N_11744);
nand U12589 (N_12589,N_11872,N_10261);
and U12590 (N_12590,N_12329,N_10479);
nand U12591 (N_12591,N_12280,N_10900);
nand U12592 (N_12592,N_12019,N_12436);
nor U12593 (N_12593,N_11227,N_10821);
xnor U12594 (N_12594,N_10070,N_11160);
and U12595 (N_12595,N_12334,N_11109);
and U12596 (N_12596,N_11050,N_10406);
and U12597 (N_12597,N_11188,N_11149);
nor U12598 (N_12598,N_11450,N_10411);
nor U12599 (N_12599,N_10149,N_10249);
nor U12600 (N_12600,N_10852,N_10238);
and U12601 (N_12601,N_11107,N_10606);
nor U12602 (N_12602,N_10673,N_11845);
or U12603 (N_12603,N_11180,N_10413);
nor U12604 (N_12604,N_12343,N_10409);
nand U12605 (N_12605,N_10712,N_11004);
nor U12606 (N_12606,N_10236,N_11839);
or U12607 (N_12607,N_11277,N_11835);
nor U12608 (N_12608,N_11549,N_10029);
and U12609 (N_12609,N_12061,N_11420);
nand U12610 (N_12610,N_11154,N_11773);
and U12611 (N_12611,N_11009,N_10474);
or U12612 (N_12612,N_10415,N_10277);
nand U12613 (N_12613,N_11446,N_11435);
nand U12614 (N_12614,N_12415,N_10456);
and U12615 (N_12615,N_11011,N_11235);
and U12616 (N_12616,N_10315,N_12040);
or U12617 (N_12617,N_11632,N_12457);
nor U12618 (N_12618,N_10408,N_11253);
nand U12619 (N_12619,N_11292,N_11785);
xor U12620 (N_12620,N_10913,N_10260);
xnor U12621 (N_12621,N_10656,N_11036);
nor U12622 (N_12622,N_11876,N_11803);
nand U12623 (N_12623,N_11825,N_10141);
nand U12624 (N_12624,N_10888,N_10763);
xnor U12625 (N_12625,N_10402,N_11543);
and U12626 (N_12626,N_11046,N_11743);
nand U12627 (N_12627,N_11014,N_11976);
nand U12628 (N_12628,N_11797,N_12197);
and U12629 (N_12629,N_11128,N_11082);
nor U12630 (N_12630,N_11546,N_11039);
xnor U12631 (N_12631,N_10817,N_12319);
or U12632 (N_12632,N_12487,N_11384);
nand U12633 (N_12633,N_10421,N_11365);
or U12634 (N_12634,N_11579,N_10929);
nor U12635 (N_12635,N_12482,N_11195);
or U12636 (N_12636,N_10581,N_11110);
xor U12637 (N_12637,N_12153,N_10403);
nand U12638 (N_12638,N_11201,N_10697);
and U12639 (N_12639,N_10692,N_12282);
nor U12640 (N_12640,N_10517,N_12121);
nor U12641 (N_12641,N_10094,N_10264);
and U12642 (N_12642,N_11762,N_10694);
nor U12643 (N_12643,N_11040,N_12149);
nor U12644 (N_12644,N_10225,N_10373);
nor U12645 (N_12645,N_10728,N_10390);
nand U12646 (N_12646,N_11264,N_10703);
or U12647 (N_12647,N_10629,N_12216);
nand U12648 (N_12648,N_10444,N_12412);
or U12649 (N_12649,N_11428,N_11608);
and U12650 (N_12650,N_10555,N_10207);
or U12651 (N_12651,N_10471,N_11525);
nor U12652 (N_12652,N_12097,N_11629);
nand U12653 (N_12653,N_10741,N_11700);
or U12654 (N_12654,N_10451,N_10708);
nand U12655 (N_12655,N_12318,N_12279);
nor U12656 (N_12656,N_11001,N_11928);
or U12657 (N_12657,N_10116,N_12350);
and U12658 (N_12658,N_11388,N_12154);
and U12659 (N_12659,N_11079,N_12313);
nor U12660 (N_12660,N_12481,N_11025);
and U12661 (N_12661,N_10494,N_11033);
or U12662 (N_12662,N_11516,N_11832);
nand U12663 (N_12663,N_10831,N_12330);
and U12664 (N_12664,N_12328,N_10774);
and U12665 (N_12665,N_12489,N_11389);
nor U12666 (N_12666,N_12339,N_12445);
and U12667 (N_12667,N_10096,N_10586);
nand U12668 (N_12668,N_10679,N_11564);
nand U12669 (N_12669,N_12390,N_11112);
or U12670 (N_12670,N_11096,N_11440);
nor U12671 (N_12671,N_11841,N_10843);
or U12672 (N_12672,N_10359,N_12332);
nand U12673 (N_12673,N_11794,N_12055);
nor U12674 (N_12674,N_10873,N_12065);
nand U12675 (N_12675,N_11438,N_10306);
and U12676 (N_12676,N_11757,N_12207);
nor U12677 (N_12677,N_11242,N_10534);
and U12678 (N_12678,N_10754,N_12127);
and U12679 (N_12679,N_11716,N_10989);
nor U12680 (N_12680,N_11890,N_12034);
nor U12681 (N_12681,N_10310,N_12361);
nor U12682 (N_12682,N_10395,N_11688);
nor U12683 (N_12683,N_11913,N_12103);
and U12684 (N_12684,N_11344,N_12373);
and U12685 (N_12685,N_10332,N_11533);
or U12686 (N_12686,N_10946,N_12308);
nor U12687 (N_12687,N_11179,N_11662);
or U12688 (N_12688,N_10633,N_10163);
or U12689 (N_12689,N_10565,N_12173);
nand U12690 (N_12690,N_11166,N_10914);
nand U12691 (N_12691,N_11519,N_10075);
nor U12692 (N_12692,N_10744,N_10020);
and U12693 (N_12693,N_11595,N_11311);
nand U12694 (N_12694,N_11823,N_11326);
nand U12695 (N_12695,N_11940,N_11944);
or U12696 (N_12696,N_11150,N_10996);
and U12697 (N_12697,N_12377,N_11470);
nor U12698 (N_12698,N_10286,N_10625);
nand U12699 (N_12699,N_10016,N_12099);
and U12700 (N_12700,N_10035,N_10064);
or U12701 (N_12701,N_10794,N_12352);
or U12702 (N_12702,N_11273,N_10809);
nor U12703 (N_12703,N_10021,N_11753);
or U12704 (N_12704,N_11709,N_10882);
nor U12705 (N_12705,N_11636,N_12400);
nor U12706 (N_12706,N_11570,N_11628);
or U12707 (N_12707,N_11086,N_11411);
or U12708 (N_12708,N_12370,N_10432);
or U12709 (N_12709,N_10111,N_11602);
or U12710 (N_12710,N_12180,N_10680);
nand U12711 (N_12711,N_10909,N_10604);
nor U12712 (N_12712,N_11220,N_10399);
nand U12713 (N_12713,N_11229,N_11198);
or U12714 (N_12714,N_10424,N_12440);
and U12715 (N_12715,N_10577,N_11867);
nor U12716 (N_12716,N_10204,N_12014);
xor U12717 (N_12717,N_11066,N_10377);
and U12718 (N_12718,N_10172,N_12499);
and U12719 (N_12719,N_12365,N_10138);
nand U12720 (N_12720,N_12455,N_11795);
nor U12721 (N_12721,N_11035,N_10214);
or U12722 (N_12722,N_11073,N_11241);
nand U12723 (N_12723,N_10276,N_10093);
and U12724 (N_12724,N_11711,N_10635);
nor U12725 (N_12725,N_12137,N_10318);
nor U12726 (N_12726,N_10525,N_12131);
nor U12727 (N_12727,N_11325,N_10423);
nand U12728 (N_12728,N_10923,N_11758);
and U12729 (N_12729,N_10626,N_10446);
or U12730 (N_12730,N_10101,N_12270);
or U12731 (N_12731,N_10681,N_12176);
nand U12732 (N_12732,N_12098,N_11436);
and U12733 (N_12733,N_12163,N_10484);
nand U12734 (N_12734,N_10793,N_11126);
or U12735 (N_12735,N_10937,N_10455);
and U12736 (N_12736,N_11346,N_10898);
or U12737 (N_12737,N_10000,N_10512);
nor U12738 (N_12738,N_10037,N_11538);
and U12739 (N_12739,N_11598,N_11676);
and U12740 (N_12740,N_10466,N_11665);
and U12741 (N_12741,N_11202,N_11781);
xor U12742 (N_12742,N_10495,N_10054);
or U12743 (N_12743,N_10156,N_11246);
or U12744 (N_12744,N_11568,N_11924);
or U12745 (N_12745,N_10642,N_10265);
and U12746 (N_12746,N_11653,N_10044);
and U12747 (N_12747,N_10045,N_10647);
nor U12748 (N_12748,N_11754,N_11251);
nor U12749 (N_12749,N_11501,N_11129);
nor U12750 (N_12750,N_11734,N_10030);
and U12751 (N_12751,N_10568,N_10397);
nand U12752 (N_12752,N_10939,N_11354);
or U12753 (N_12753,N_11349,N_11103);
and U12754 (N_12754,N_10487,N_10894);
nand U12755 (N_12755,N_12041,N_11736);
or U12756 (N_12756,N_10031,N_10095);
nand U12757 (N_12757,N_12434,N_10463);
or U12758 (N_12758,N_12276,N_10958);
and U12759 (N_12759,N_11534,N_11555);
or U12760 (N_12760,N_11994,N_10963);
nand U12761 (N_12761,N_10798,N_10883);
or U12762 (N_12762,N_11158,N_10392);
nor U12763 (N_12763,N_10691,N_12311);
nor U12764 (N_12764,N_10497,N_10335);
nand U12765 (N_12765,N_10362,N_10007);
or U12766 (N_12766,N_11798,N_11288);
or U12767 (N_12767,N_11207,N_11609);
and U12768 (N_12768,N_10239,N_10314);
and U12769 (N_12769,N_10280,N_10227);
and U12770 (N_12770,N_12454,N_10917);
nand U12771 (N_12771,N_12430,N_10722);
or U12772 (N_12772,N_11452,N_11638);
or U12773 (N_12773,N_11392,N_11614);
nor U12774 (N_12774,N_10878,N_12367);
and U12775 (N_12775,N_10319,N_10475);
or U12776 (N_12776,N_10863,N_11374);
nor U12777 (N_12777,N_12138,N_10905);
nor U12778 (N_12778,N_10788,N_11209);
or U12779 (N_12779,N_10750,N_10645);
nand U12780 (N_12780,N_10920,N_10439);
and U12781 (N_12781,N_11694,N_11511);
nor U12782 (N_12782,N_12397,N_10526);
nor U12783 (N_12783,N_12012,N_10739);
nor U12784 (N_12784,N_10235,N_10440);
and U12785 (N_12785,N_12023,N_10354);
nand U12786 (N_12786,N_10557,N_10698);
and U12787 (N_12787,N_10072,N_10848);
xor U12788 (N_12788,N_11740,N_11986);
or U12789 (N_12789,N_12174,N_10420);
nand U12790 (N_12790,N_11281,N_10709);
and U12791 (N_12791,N_11646,N_10748);
or U12792 (N_12792,N_11936,N_11548);
and U12793 (N_12793,N_11576,N_10099);
and U12794 (N_12794,N_10772,N_10576);
and U12795 (N_12795,N_11977,N_10719);
or U12796 (N_12796,N_10223,N_12073);
nor U12797 (N_12797,N_11348,N_10231);
nand U12798 (N_12798,N_10536,N_10844);
nand U12799 (N_12799,N_10792,N_11810);
and U12800 (N_12800,N_11425,N_11732);
or U12801 (N_12801,N_10993,N_11880);
and U12802 (N_12802,N_12222,N_11423);
nor U12803 (N_12803,N_10791,N_11654);
nand U12804 (N_12804,N_10761,N_12064);
nor U12805 (N_12805,N_11644,N_11691);
xor U12806 (N_12806,N_11286,N_10735);
or U12807 (N_12807,N_11067,N_10800);
nor U12808 (N_12808,N_10601,N_10705);
and U12809 (N_12809,N_11212,N_12299);
and U12810 (N_12810,N_11305,N_12428);
nand U12811 (N_12811,N_11875,N_11929);
nor U12812 (N_12812,N_10130,N_10702);
nand U12813 (N_12813,N_12356,N_10081);
or U12814 (N_12814,N_10871,N_10634);
or U12815 (N_12815,N_10818,N_11639);
nand U12816 (N_12816,N_12026,N_11020);
nor U12817 (N_12817,N_11413,N_11468);
or U12818 (N_12818,N_10780,N_10564);
and U12819 (N_12819,N_11172,N_11901);
nor U12820 (N_12820,N_10146,N_11942);
or U12821 (N_12821,N_10575,N_10025);
or U12822 (N_12822,N_11617,N_12347);
or U12823 (N_12823,N_11796,N_10603);
nor U12824 (N_12824,N_10043,N_12001);
nor U12825 (N_12825,N_11643,N_11453);
or U12826 (N_12826,N_11098,N_11467);
and U12827 (N_12827,N_10858,N_10023);
nor U12828 (N_12828,N_10032,N_12460);
nand U12829 (N_12829,N_11381,N_11505);
and U12830 (N_12830,N_12227,N_11012);
nand U12831 (N_12831,N_10067,N_11234);
nor U12832 (N_12832,N_10368,N_10124);
or U12833 (N_12833,N_10677,N_10562);
nand U12834 (N_12834,N_11927,N_11016);
nand U12835 (N_12835,N_12038,N_10435);
and U12836 (N_12836,N_11879,N_10540);
or U12837 (N_12837,N_12241,N_10273);
nand U12838 (N_12838,N_11829,N_11583);
nand U12839 (N_12839,N_10302,N_11843);
and U12840 (N_12840,N_11637,N_10425);
and U12841 (N_12841,N_10543,N_12226);
nand U12842 (N_12842,N_10272,N_12076);
nor U12843 (N_12843,N_12231,N_10499);
and U12844 (N_12844,N_11403,N_10296);
or U12845 (N_12845,N_10819,N_10004);
and U12846 (N_12846,N_12309,N_11692);
and U12847 (N_12847,N_12291,N_10622);
or U12848 (N_12848,N_10807,N_10457);
nor U12849 (N_12849,N_11604,N_11027);
nor U12850 (N_12850,N_11285,N_12030);
nand U12851 (N_12851,N_11704,N_12204);
nand U12852 (N_12852,N_10062,N_10449);
nor U12853 (N_12853,N_11912,N_11226);
and U12854 (N_12854,N_11416,N_11620);
nor U12855 (N_12855,N_12144,N_12447);
nand U12856 (N_12856,N_10166,N_11983);
nand U12857 (N_12857,N_10082,N_10074);
nor U12858 (N_12858,N_11958,N_11647);
nand U12859 (N_12859,N_11019,N_11041);
and U12860 (N_12860,N_11336,N_10976);
or U12861 (N_12861,N_10723,N_11926);
nand U12862 (N_12862,N_10103,N_11297);
and U12863 (N_12863,N_10663,N_10738);
nand U12864 (N_12864,N_10734,N_12444);
nor U12865 (N_12865,N_10891,N_10248);
and U12866 (N_12866,N_11828,N_12018);
nand U12867 (N_12867,N_12194,N_10653);
nand U12868 (N_12868,N_11811,N_10872);
and U12869 (N_12869,N_10226,N_10860);
and U12870 (N_12870,N_12090,N_11593);
or U12871 (N_12871,N_10637,N_10325);
nor U12872 (N_12872,N_12184,N_10941);
and U12873 (N_12873,N_10090,N_12128);
nor U12874 (N_12874,N_10825,N_12053);
nand U12875 (N_12875,N_11216,N_11968);
nor U12876 (N_12876,N_11415,N_11989);
and U12877 (N_12877,N_11562,N_10243);
and U12878 (N_12878,N_10853,N_10766);
and U12879 (N_12879,N_11142,N_12247);
or U12880 (N_12880,N_12045,N_10767);
or U12881 (N_12881,N_11171,N_11061);
and U12882 (N_12882,N_11771,N_10097);
or U12883 (N_12883,N_10470,N_12067);
or U12884 (N_12884,N_11274,N_11550);
or U12885 (N_12885,N_10500,N_10830);
or U12886 (N_12886,N_10112,N_10157);
nand U12887 (N_12887,N_11815,N_10519);
nor U12888 (N_12888,N_11031,N_12211);
nand U12889 (N_12889,N_12158,N_10178);
or U12890 (N_12890,N_10861,N_10340);
and U12891 (N_12891,N_11048,N_11243);
or U12892 (N_12892,N_11186,N_11111);
nand U12893 (N_12893,N_11949,N_10483);
nor U12894 (N_12894,N_12111,N_11013);
or U12895 (N_12895,N_10893,N_11535);
nand U12896 (N_12896,N_10755,N_10155);
and U12897 (N_12897,N_10822,N_11399);
nor U12898 (N_12898,N_11974,N_10592);
nor U12899 (N_12899,N_12446,N_10352);
and U12900 (N_12900,N_11029,N_11307);
and U12901 (N_12901,N_11437,N_11641);
or U12902 (N_12902,N_11417,N_10284);
nand U12903 (N_12903,N_11120,N_11244);
nor U12904 (N_12904,N_10185,N_11249);
and U12905 (N_12905,N_11104,N_11200);
and U12906 (N_12906,N_11204,N_10870);
or U12907 (N_12907,N_12476,N_11386);
nor U12908 (N_12908,N_11445,N_11520);
or U12909 (N_12909,N_12463,N_10566);
and U12910 (N_12910,N_12109,N_10944);
and U12911 (N_12911,N_12160,N_12000);
xnor U12912 (N_12912,N_11459,N_10026);
and U12913 (N_12913,N_11752,N_12404);
nor U12914 (N_12914,N_11359,N_11260);
nand U12915 (N_12915,N_12105,N_12136);
nor U12916 (N_12916,N_10867,N_11559);
nor U12917 (N_12917,N_11356,N_10193);
and U12918 (N_12918,N_10776,N_10197);
and U12919 (N_12919,N_11328,N_10419);
and U12920 (N_12920,N_12498,N_11105);
nor U12921 (N_12921,N_12341,N_10118);
nand U12922 (N_12922,N_10641,N_11056);
nand U12923 (N_12923,N_11108,N_10289);
and U12924 (N_12924,N_11655,N_10339);
nor U12925 (N_12925,N_12042,N_12418);
or U12926 (N_12926,N_10279,N_12170);
nand U12927 (N_12927,N_10777,N_11371);
or U12928 (N_12928,N_10052,N_11883);
or U12929 (N_12929,N_11613,N_10978);
and U12930 (N_12930,N_12116,N_11592);
and U12931 (N_12931,N_12199,N_12437);
nor U12932 (N_12932,N_11444,N_10632);
nand U12933 (N_12933,N_10164,N_11065);
or U12934 (N_12934,N_11355,N_12345);
nand U12935 (N_12935,N_10814,N_11540);
or U12936 (N_12936,N_10934,N_10682);
nand U12937 (N_12937,N_11370,N_10924);
nor U12938 (N_12938,N_12383,N_12235);
nor U12939 (N_12939,N_10433,N_11222);
and U12940 (N_12940,N_12312,N_10742);
and U12941 (N_12941,N_11458,N_10636);
and U12942 (N_12942,N_10610,N_12134);
or U12943 (N_12943,N_11181,N_11713);
and U12944 (N_12944,N_11556,N_10469);
nor U12945 (N_12945,N_11854,N_11707);
or U12946 (N_12946,N_11021,N_10862);
nand U12947 (N_12947,N_12301,N_11693);
and U12948 (N_12948,N_10935,N_10573);
nor U12949 (N_12949,N_11457,N_10211);
nor U12950 (N_12950,N_10579,N_11908);
nor U12951 (N_12951,N_10358,N_11464);
nand U12952 (N_12952,N_11071,N_10387);
and U12953 (N_12953,N_11199,N_10689);
xnor U12954 (N_12954,N_10417,N_11955);
nand U12955 (N_12955,N_11510,N_11139);
and U12956 (N_12956,N_10583,N_10110);
nand U12957 (N_12957,N_10879,N_10903);
nand U12958 (N_12958,N_10832,N_11218);
and U12959 (N_12959,N_11341,N_10770);
nor U12960 (N_12960,N_11504,N_10355);
and U12961 (N_12961,N_12479,N_10217);
and U12962 (N_12962,N_10756,N_10884);
and U12963 (N_12963,N_12459,N_11024);
nand U12964 (N_12964,N_11818,N_12193);
and U12965 (N_12965,N_12269,N_11884);
nand U12966 (N_12966,N_10160,N_12398);
nor U12967 (N_12967,N_11406,N_10088);
nand U12968 (N_12968,N_10585,N_11455);
and U12969 (N_12969,N_11739,N_10940);
nand U12970 (N_12970,N_11774,N_12198);
and U12971 (N_12971,N_11231,N_10816);
and U12972 (N_12972,N_11337,N_10290);
nand U12973 (N_12973,N_11342,N_11034);
nand U12974 (N_12974,N_11663,N_12477);
and U12975 (N_12975,N_11002,N_10102);
or U12976 (N_12976,N_12303,N_10136);
and U12977 (N_12977,N_10281,N_10049);
nor U12978 (N_12978,N_11184,N_10614);
and U12979 (N_12979,N_11809,N_10528);
xor U12980 (N_12980,N_12141,N_11581);
or U12981 (N_12981,N_10184,N_10541);
nand U12982 (N_12982,N_11775,N_12432);
nor U12983 (N_12983,N_10721,N_12119);
nand U12984 (N_12984,N_10380,N_12369);
nor U12985 (N_12985,N_11611,N_10762);
nand U12986 (N_12986,N_10312,N_10391);
nor U12987 (N_12987,N_12491,N_10595);
and U12988 (N_12988,N_11566,N_12069);
and U12989 (N_12989,N_11282,N_11650);
nand U12990 (N_12990,N_11652,N_11206);
or U12991 (N_12991,N_11456,N_10459);
nand U12992 (N_12992,N_11228,N_10580);
or U12993 (N_12993,N_10307,N_12317);
nor U12994 (N_12994,N_10987,N_10911);
nand U12995 (N_12995,N_11920,N_10795);
and U12996 (N_12996,N_10437,N_11574);
nor U12997 (N_12997,N_12416,N_10842);
and U12998 (N_12998,N_10502,N_10039);
or U12999 (N_12999,N_11116,N_10665);
and U13000 (N_13000,N_12413,N_10154);
or U13001 (N_13001,N_11352,N_11263);
and U13002 (N_13002,N_11745,N_10859);
nand U13003 (N_13003,N_10925,N_11267);
and U13004 (N_13004,N_10244,N_12095);
or U13005 (N_13005,N_11886,N_12027);
and U13006 (N_13006,N_11715,N_10785);
nand U13007 (N_13007,N_12348,N_10959);
or U13008 (N_13008,N_10549,N_12472);
xor U13009 (N_13009,N_12151,N_11779);
or U13010 (N_13010,N_11575,N_10334);
nor U13011 (N_13011,N_12395,N_10839);
and U13012 (N_13012,N_10804,N_10121);
and U13013 (N_13013,N_11834,N_11390);
nor U13014 (N_13014,N_12417,N_11256);
nor U13015 (N_13015,N_11463,N_11010);
and U13016 (N_13016,N_12191,N_10477);
or U13017 (N_13017,N_10438,N_12132);
or U13018 (N_13018,N_12494,N_11967);
or U13019 (N_13019,N_10203,N_11850);
or U13020 (N_13020,N_11043,N_10431);
nor U13021 (N_13021,N_11618,N_11363);
or U13022 (N_13022,N_10005,N_11076);
nor U13023 (N_13023,N_11971,N_11394);
nor U13024 (N_13024,N_11975,N_11668);
nor U13025 (N_13025,N_10998,N_10646);
or U13026 (N_13026,N_11634,N_10092);
nand U13027 (N_13027,N_10367,N_10802);
or U13028 (N_13028,N_10034,N_10919);
or U13029 (N_13029,N_11164,N_11094);
nor U13030 (N_13030,N_12033,N_10287);
and U13031 (N_13031,N_12147,N_10104);
or U13032 (N_13032,N_11481,N_10485);
nand U13033 (N_13033,N_12366,N_11053);
nor U13034 (N_13034,N_12100,N_10751);
nor U13035 (N_13035,N_10983,N_10385);
nor U13036 (N_13036,N_10511,N_10491);
or U13037 (N_13037,N_11848,N_11657);
or U13038 (N_13038,N_11888,N_11439);
and U13039 (N_13039,N_12165,N_12331);
nand U13040 (N_13040,N_12399,N_10055);
or U13041 (N_13041,N_10768,N_10400);
nor U13042 (N_13042,N_11152,N_11932);
nor U13043 (N_13043,N_10202,N_10600);
or U13044 (N_13044,N_11443,N_10200);
and U13045 (N_13045,N_11865,N_12175);
and U13046 (N_13046,N_11447,N_10324);
and U13047 (N_13047,N_12142,N_10270);
nand U13048 (N_13048,N_11907,N_11649);
and U13049 (N_13049,N_10538,N_10612);
and U13050 (N_13050,N_11860,N_12266);
or U13051 (N_13051,N_11672,N_10743);
nand U13052 (N_13052,N_10501,N_12409);
nand U13053 (N_13053,N_10980,N_11493);
nand U13054 (N_13054,N_11686,N_10304);
or U13055 (N_13055,N_11589,N_12429);
nor U13056 (N_13056,N_11768,N_10933);
nor U13057 (N_13057,N_11630,N_11407);
nor U13058 (N_13058,N_10109,N_11368);
and U13059 (N_13059,N_11635,N_11874);
nor U13060 (N_13060,N_11896,N_11426);
or U13061 (N_13061,N_11671,N_11490);
and U13062 (N_13062,N_11397,N_12050);
xnor U13063 (N_13063,N_12037,N_12245);
or U13064 (N_13064,N_10012,N_11135);
or U13065 (N_13065,N_12264,N_12351);
and U13066 (N_13066,N_10667,N_11542);
nor U13067 (N_13067,N_10889,N_11489);
and U13068 (N_13068,N_12401,N_10125);
or U13069 (N_13069,N_10569,N_10047);
nand U13070 (N_13070,N_11933,N_10773);
or U13071 (N_13071,N_11049,N_11786);
nand U13072 (N_13072,N_11787,N_11612);
nor U13073 (N_13073,N_12043,N_12046);
nand U13074 (N_13074,N_11278,N_11169);
or U13075 (N_13075,N_12240,N_12115);
and U13076 (N_13076,N_11712,N_11018);
xor U13077 (N_13077,N_11805,N_10194);
nor U13078 (N_13078,N_11963,N_11517);
and U13079 (N_13079,N_10418,N_10251);
or U13080 (N_13080,N_11118,N_11089);
and U13081 (N_13081,N_10544,N_10704);
nand U13082 (N_13082,N_11966,N_12188);
and U13083 (N_13083,N_11090,N_12357);
or U13084 (N_13084,N_10558,N_11964);
or U13085 (N_13085,N_12310,N_12305);
or U13086 (N_13086,N_10970,N_11093);
nand U13087 (N_13087,N_11871,N_10857);
nand U13088 (N_13088,N_10574,N_11760);
or U13089 (N_13089,N_10376,N_10165);
and U13090 (N_13090,N_11899,N_10119);
and U13091 (N_13091,N_11943,N_12322);
nor U13092 (N_13092,N_12057,N_11861);
nor U13093 (N_13093,N_11176,N_10910);
nor U13094 (N_13094,N_10664,N_11230);
nand U13095 (N_13095,N_12325,N_10880);
or U13096 (N_13096,N_10509,N_10589);
nand U13097 (N_13097,N_11826,N_11422);
nor U13098 (N_13098,N_10956,N_12267);
and U13099 (N_13099,N_11473,N_12152);
and U13100 (N_13100,N_11333,N_10797);
and U13101 (N_13101,N_12162,N_12451);
or U13102 (N_13102,N_12324,N_11174);
and U13103 (N_13103,N_11980,N_11315);
nand U13104 (N_13104,N_10215,N_10008);
and U13105 (N_13105,N_12051,N_11914);
xor U13106 (N_13106,N_11960,N_11723);
or U13107 (N_13107,N_11151,N_10826);
nor U13108 (N_13108,N_10532,N_10452);
and U13109 (N_13109,N_10942,N_10651);
and U13110 (N_13110,N_10660,N_11213);
or U13111 (N_13111,N_11347,N_11801);
and U13112 (N_13112,N_11466,N_10375);
nand U13113 (N_13113,N_10675,N_12333);
nand U13114 (N_13114,N_10718,N_12177);
nand U13115 (N_13115,N_10065,N_10209);
nor U13116 (N_13116,N_10322,N_11623);
nor U13117 (N_13117,N_10283,N_12326);
nor U13118 (N_13118,N_10904,N_10790);
nor U13119 (N_13119,N_10545,N_12145);
and U13120 (N_13120,N_11846,N_12284);
or U13121 (N_13121,N_10308,N_11837);
or U13122 (N_13122,N_12255,N_12493);
nand U13123 (N_13123,N_10551,N_12360);
nand U13124 (N_13124,N_12408,N_10892);
and U13125 (N_13125,N_10069,N_11847);
nor U13126 (N_13126,N_12171,N_11844);
or U13127 (N_13127,N_12020,N_11449);
xnor U13128 (N_13128,N_10700,N_10148);
and U13129 (N_13129,N_10508,N_12243);
xor U13130 (N_13130,N_10011,N_12139);
and U13131 (N_13131,N_12262,N_12209);
nand U13132 (N_13132,N_10053,N_12104);
nand U13133 (N_13133,N_11156,N_10357);
or U13134 (N_13134,N_10676,N_11895);
or U13135 (N_13135,N_11335,N_10627);
and U13136 (N_13136,N_11398,N_10764);
nand U13137 (N_13137,N_10683,N_12093);
nor U13138 (N_13138,N_10300,N_10208);
nor U13139 (N_13139,N_12380,N_11996);
or U13140 (N_13140,N_10533,N_10346);
or U13141 (N_13141,N_11391,N_10317);
or U13142 (N_13142,N_10806,N_11210);
nor U13143 (N_13143,N_11626,N_10961);
nor U13144 (N_13144,N_11357,N_12354);
or U13145 (N_13145,N_10786,N_12353);
and U13146 (N_13146,N_10087,N_11748);
or U13147 (N_13147,N_10548,N_10305);
nor U13148 (N_13148,N_10779,N_10567);
nor U13149 (N_13149,N_10829,N_10518);
or U13150 (N_13150,N_11957,N_10981);
and U13151 (N_13151,N_10962,N_11434);
and U13152 (N_13152,N_11431,N_10151);
or U13153 (N_13153,N_11334,N_12287);
and U13154 (N_13154,N_11287,N_10212);
and U13155 (N_13155,N_10927,N_12288);
nand U13156 (N_13156,N_10349,N_11500);
and U13157 (N_13157,N_11058,N_12016);
nor U13158 (N_13158,N_11295,N_12228);
nor U13159 (N_13159,N_11730,N_11194);
or U13160 (N_13160,N_10171,N_12402);
nor U13161 (N_13161,N_11350,N_11696);
nand U13162 (N_13162,N_12265,N_11448);
and U13163 (N_13163,N_10609,N_11182);
nor U13164 (N_13164,N_10918,N_10661);
and U13165 (N_13165,N_10758,N_11778);
or U13166 (N_13166,N_11462,N_10106);
nand U13167 (N_13167,N_10429,N_12306);
and U13168 (N_13168,N_11279,N_11044);
and U13169 (N_13169,N_11950,N_11143);
xor U13170 (N_13170,N_10803,N_10966);
nand U13171 (N_13171,N_10938,N_11161);
xnor U13172 (N_13172,N_11669,N_11881);
nand U13173 (N_13173,N_11954,N_12466);
and U13174 (N_13174,N_11134,N_10955);
nor U13175 (N_13175,N_11469,N_12258);
or U13176 (N_13176,N_10605,N_10115);
nor U13177 (N_13177,N_11310,N_11183);
nor U13178 (N_13178,N_12458,N_10572);
nor U13179 (N_13179,N_10177,N_10003);
nor U13180 (N_13180,N_10967,N_12075);
nand U13181 (N_13181,N_10699,N_12049);
or U13182 (N_13182,N_10740,N_11320);
or U13183 (N_13183,N_11807,N_12392);
nand U13184 (N_13184,N_11115,N_10405);
or U13185 (N_13185,N_10033,N_10256);
or U13186 (N_13186,N_11003,N_11911);
nand U13187 (N_13187,N_12143,N_10902);
or U13188 (N_13188,N_10957,N_12300);
nor U13189 (N_13189,N_10038,N_12372);
and U13190 (N_13190,N_11396,N_11838);
nor U13191 (N_13191,N_10142,N_10229);
nor U13192 (N_13192,N_12196,N_10874);
and U13193 (N_13193,N_11741,N_11343);
and U13194 (N_13194,N_11733,N_11170);
nand U13195 (N_13195,N_10372,N_12424);
or U13196 (N_13196,N_11793,N_11084);
nor U13197 (N_13197,N_11527,N_11257);
nor U13198 (N_13198,N_10999,N_10232);
nand U13199 (N_13199,N_11271,N_11529);
and U13200 (N_13200,N_11503,N_11121);
and U13201 (N_13201,N_10971,N_10162);
and U13202 (N_13202,N_12316,N_11719);
and U13203 (N_13203,N_10596,N_11681);
nor U13204 (N_13204,N_10268,N_12223);
nand U13205 (N_13205,N_10496,N_11095);
or U13206 (N_13206,N_10453,N_11658);
nor U13207 (N_13207,N_10654,N_10128);
or U13208 (N_13208,N_11283,N_11148);
or U13209 (N_13209,N_11113,N_11864);
nor U13210 (N_13210,N_11670,N_12385);
or U13211 (N_13211,N_11364,N_11679);
nand U13212 (N_13212,N_11536,N_12234);
or U13213 (N_13213,N_11897,N_10476);
or U13214 (N_13214,N_10205,N_10181);
or U13215 (N_13215,N_10326,N_10493);
nand U13216 (N_13216,N_10068,N_10180);
or U13217 (N_13217,N_10578,N_11051);
and U13218 (N_13218,N_10394,N_11763);
nand U13219 (N_13219,N_10114,N_11318);
or U13220 (N_13220,N_10602,N_10084);
nand U13221 (N_13221,N_12155,N_11645);
and U13222 (N_13222,N_10781,N_11474);
and U13223 (N_13223,N_10255,N_10973);
or U13224 (N_13224,N_10199,N_12084);
and U13225 (N_13225,N_12410,N_11780);
or U13226 (N_13226,N_11159,N_10554);
and U13227 (N_13227,N_10507,N_10131);
nand U13228 (N_13228,N_11193,N_11097);
or U13229 (N_13229,N_12275,N_11640);
nand U13230 (N_13230,N_12219,N_12277);
xnor U13231 (N_13231,N_12017,N_11313);
or U13232 (N_13232,N_10196,N_10932);
nor U13233 (N_13233,N_10472,N_10556);
nor U13234 (N_13234,N_11008,N_12349);
nand U13235 (N_13235,N_10327,N_10174);
nand U13236 (N_13236,N_11677,N_11157);
and U13237 (N_13237,N_12220,N_11258);
nand U13238 (N_13238,N_12257,N_11026);
and U13239 (N_13239,N_11380,N_12426);
nand U13240 (N_13240,N_11302,N_10765);
and U13241 (N_13241,N_11934,N_12251);
nor U13242 (N_13242,N_10465,N_10127);
or U13243 (N_13243,N_10837,N_10140);
nand U13244 (N_13244,N_11856,N_10678);
and U13245 (N_13245,N_11528,N_11175);
or U13246 (N_13246,N_11951,N_12338);
or U13247 (N_13247,N_10117,N_11978);
xnor U13248 (N_13248,N_10685,N_10984);
nor U13249 (N_13249,N_10242,N_11395);
nand U13250 (N_13250,N_10733,N_11660);
nor U13251 (N_13251,N_12140,N_11915);
and U13252 (N_13252,N_10877,N_12157);
or U13253 (N_13253,N_10907,N_11475);
nand U13254 (N_13254,N_11705,N_10191);
and U13255 (N_13255,N_10401,N_10370);
nor U13256 (N_13256,N_11678,N_10520);
or U13257 (N_13257,N_12200,N_10997);
nand U13258 (N_13258,N_11379,N_11689);
and U13259 (N_13259,N_11137,N_11189);
nand U13260 (N_13260,N_12358,N_12011);
or U13261 (N_13261,N_11521,N_10108);
nor U13262 (N_13262,N_11419,N_12407);
nor U13263 (N_13263,N_10309,N_10182);
nand U13264 (N_13264,N_10382,N_11289);
nor U13265 (N_13265,N_10710,N_12420);
or U13266 (N_13266,N_12192,N_10828);
nor U13267 (N_13267,N_12393,N_11197);
or U13268 (N_13268,N_11138,N_10169);
nor U13269 (N_13269,N_11429,N_10428);
nor U13270 (N_13270,N_10542,N_11114);
xor U13271 (N_13271,N_12248,N_11727);
nand U13272 (N_13272,N_11377,N_10059);
or U13273 (N_13273,N_10240,N_10018);
and U13274 (N_13274,N_11889,N_11599);
nor U13275 (N_13275,N_10553,N_12083);
nor U13276 (N_13276,N_11378,N_12346);
nor U13277 (N_13277,N_10823,N_10224);
nand U13278 (N_13278,N_11921,N_10303);
or U13279 (N_13279,N_12123,N_10135);
nand U13280 (N_13280,N_11430,N_10936);
nand U13281 (N_13281,N_10374,N_12382);
or U13282 (N_13282,N_11479,N_11935);
or U13283 (N_13283,N_10430,N_10875);
nor U13284 (N_13284,N_12478,N_10531);
or U13285 (N_13285,N_12133,N_11147);
nor U13286 (N_13286,N_11792,N_10515);
xor U13287 (N_13287,N_11339,N_11091);
nand U13288 (N_13288,N_12167,N_10462);
and U13289 (N_13289,N_10855,N_10631);
nand U13290 (N_13290,N_12293,N_11833);
and U13291 (N_13291,N_10356,N_11322);
or U13292 (N_13292,N_10295,N_12169);
nor U13293 (N_13293,N_10183,N_11830);
and U13294 (N_13294,N_11340,N_12389);
nand U13295 (N_13295,N_11674,N_10458);
or U13296 (N_13296,N_10473,N_11409);
nand U13297 (N_13297,N_10864,N_10648);
and U13298 (N_13298,N_10707,N_11465);
or U13299 (N_13299,N_11023,N_11656);
and U13300 (N_13300,N_10982,N_12381);
xor U13301 (N_13301,N_12427,N_10271);
nand U13302 (N_13302,N_10330,N_10027);
or U13303 (N_13303,N_11666,N_11366);
xnor U13304 (N_13304,N_12315,N_12485);
and U13305 (N_13305,N_10649,N_10233);
nor U13306 (N_13306,N_11319,N_11136);
and U13307 (N_13307,N_12117,N_10926);
nor U13308 (N_13308,N_10856,N_10274);
nor U13309 (N_13309,N_12336,N_10301);
nor U13310 (N_13310,N_11999,N_11270);
and U13311 (N_13311,N_12419,N_11627);
nor U13312 (N_13312,N_11591,N_12296);
nor U13313 (N_13313,N_10570,N_12074);
nor U13314 (N_13314,N_10173,N_10187);
or U13315 (N_13315,N_10945,N_12189);
nand U13316 (N_13316,N_10086,N_10139);
or U13317 (N_13317,N_11495,N_10666);
and U13318 (N_13318,N_11814,N_10262);
nand U13319 (N_13319,N_11032,N_12089);
nor U13320 (N_13320,N_10080,N_11502);
nor U13321 (N_13321,N_12007,N_10351);
and U13322 (N_13322,N_11028,N_10328);
nor U13323 (N_13323,N_12492,N_10985);
or U13324 (N_13324,N_11698,N_11858);
xor U13325 (N_13325,N_10383,N_11421);
xor U13326 (N_13326,N_11891,N_11873);
nand U13327 (N_13327,N_11099,N_12456);
nand U13328 (N_13328,N_10584,N_11893);
or U13329 (N_13329,N_12047,N_10977);
nor U13330 (N_13330,N_10066,N_11675);
xor U13331 (N_13331,N_11819,N_11699);
nor U13332 (N_13332,N_11987,N_12068);
nand U13333 (N_13333,N_11214,N_11165);
nor U13334 (N_13334,N_11939,N_11731);
and U13335 (N_13335,N_10639,N_10407);
nor U13336 (N_13336,N_11588,N_10992);
nor U13337 (N_13337,N_11972,N_11078);
and U13338 (N_13338,N_12281,N_10897);
nor U13339 (N_13339,N_10345,N_10498);
nor U13340 (N_13340,N_11991,N_11948);
nand U13341 (N_13341,N_11769,N_11585);
nor U13342 (N_13342,N_10726,N_10153);
nand U13343 (N_13343,N_12268,N_12087);
nand U13344 (N_13344,N_11223,N_10336);
nand U13345 (N_13345,N_12474,N_11125);
nand U13346 (N_13346,N_10617,N_10834);
or U13347 (N_13347,N_10291,N_12379);
and U13348 (N_13348,N_10787,N_12320);
and U13349 (N_13349,N_10597,N_10198);
or U13350 (N_13350,N_12448,N_11747);
nor U13351 (N_13351,N_10954,N_12232);
or U13352 (N_13352,N_11906,N_11068);
nor U13353 (N_13353,N_11498,N_12183);
nor U13354 (N_13354,N_10953,N_10079);
nor U13355 (N_13355,N_10561,N_11367);
and U13356 (N_13356,N_11080,N_12081);
and U13357 (N_13357,N_10594,N_10017);
and U13358 (N_13358,N_11100,N_10729);
nor U13359 (N_13359,N_12150,N_10845);
nand U13360 (N_13360,N_11751,N_11894);
and U13361 (N_13361,N_11192,N_11092);
nand U13362 (N_13362,N_12187,N_12327);
nand U13363 (N_13363,N_11215,N_12254);
nand U13364 (N_13364,N_10969,N_12124);
or U13365 (N_13365,N_10524,N_10850);
or U13366 (N_13366,N_11106,N_10492);
nand U13367 (N_13367,N_10599,N_12386);
nor U13368 (N_13368,N_10412,N_12464);
nand U13369 (N_13369,N_11537,N_11750);
and U13370 (N_13370,N_10922,N_10091);
nand U13371 (N_13371,N_11211,N_12253);
and U13372 (N_13372,N_11488,N_10006);
or U13373 (N_13373,N_10036,N_12441);
nand U13374 (N_13374,N_10789,N_11132);
or U13375 (N_13375,N_11101,N_10717);
xor U13376 (N_13376,N_12283,N_10671);
nor U13377 (N_13377,N_10275,N_12164);
and U13378 (N_13378,N_10638,N_10042);
nand U13379 (N_13379,N_11130,N_10058);
nor U13380 (N_13380,N_10886,N_10887);
nand U13381 (N_13381,N_12005,N_10838);
nand U13382 (N_13382,N_12102,N_12125);
nand U13383 (N_13383,N_10948,N_12070);
or U13384 (N_13384,N_11738,N_10840);
nor U13385 (N_13385,N_11631,N_11729);
nor U13386 (N_13386,N_12422,N_10906);
and U13387 (N_13387,N_11327,N_11789);
nand U13388 (N_13388,N_11610,N_11673);
nor U13389 (N_13389,N_10771,N_11772);
or U13390 (N_13390,N_11784,N_10478);
nand U13391 (N_13391,N_11254,N_12470);
nand U13392 (N_13392,N_12355,N_10696);
nor U13393 (N_13393,N_10145,N_12048);
nand U13394 (N_13394,N_11607,N_11737);
nand U13395 (N_13395,N_10760,N_10416);
and U13396 (N_13396,N_11539,N_10293);
and U13397 (N_13397,N_10737,N_12063);
nand U13398 (N_13398,N_12181,N_10076);
nor U13399 (N_13399,N_11303,N_11523);
nand U13400 (N_13400,N_10881,N_12229);
and U13401 (N_13401,N_11515,N_10294);
and U13402 (N_13402,N_10527,N_10061);
nor U13403 (N_13403,N_11563,N_11376);
or U13404 (N_13404,N_12246,N_10812);
and U13405 (N_13405,N_11714,N_11265);
xnor U13406 (N_13406,N_10057,N_11296);
and U13407 (N_13407,N_10482,N_11782);
and U13408 (N_13408,N_10254,N_11953);
and U13409 (N_13409,N_11836,N_10347);
and U13410 (N_13410,N_12391,N_10669);
and U13411 (N_13411,N_10921,N_11369);
nor U13412 (N_13412,N_12368,N_10230);
and U13413 (N_13413,N_12244,N_11221);
nand U13414 (N_13414,N_10134,N_10706);
nor U13415 (N_13415,N_11454,N_10745);
nor U13416 (N_13416,N_12221,N_12060);
and U13417 (N_13417,N_12021,N_12433);
and U13418 (N_13418,N_12004,N_11684);
nand U13419 (N_13419,N_11372,N_10775);
or U13420 (N_13420,N_11544,N_11240);
and U13421 (N_13421,N_11410,N_10379);
and U13422 (N_13422,N_10899,N_10333);
or U13423 (N_13423,N_11554,N_10176);
and U13424 (N_13424,N_12431,N_12302);
nor U13425 (N_13425,N_10009,N_10931);
nand U13426 (N_13426,N_10213,N_11905);
nand U13427 (N_13427,N_12112,N_11233);
and U13428 (N_13428,N_12488,N_10835);
and U13429 (N_13429,N_12054,N_12059);
and U13430 (N_13430,N_10461,N_10563);
or U13431 (N_13431,N_11237,N_12475);
and U13432 (N_13432,N_11590,N_11765);
and U13433 (N_13433,N_10158,N_11492);
and U13434 (N_13434,N_11993,N_11962);
nand U13435 (N_13435,N_12242,N_11821);
xnor U13436 (N_13436,N_11045,N_11909);
nand U13437 (N_13437,N_12495,N_10630);
xor U13438 (N_13438,N_11509,N_11621);
or U13439 (N_13439,N_11268,N_11400);
nand U13440 (N_13440,N_11685,N_12394);
and U13441 (N_13441,N_12206,N_12035);
nor U13442 (N_13442,N_11085,N_11259);
xor U13443 (N_13443,N_12225,N_11059);
nand U13444 (N_13444,N_11037,N_11007);
or U13445 (N_13445,N_10123,N_11822);
nand U13446 (N_13446,N_11600,N_11887);
nand U13447 (N_13447,N_12469,N_10731);
or U13448 (N_13448,N_11191,N_12224);
nand U13449 (N_13449,N_11664,N_11405);
nor U13450 (N_13450,N_10950,N_12039);
or U13451 (N_13451,N_10100,N_11276);
nand U13452 (N_13452,N_12467,N_10990);
or U13453 (N_13453,N_10598,N_11131);
nor U13454 (N_13454,N_10299,N_11746);
nand U13455 (N_13455,N_10810,N_10991);
or U13456 (N_13456,N_11402,N_10974);
or U13457 (N_13457,N_11605,N_12307);
xor U13458 (N_13458,N_11250,N_11956);
nor U13459 (N_13459,N_10778,N_10316);
nor U13460 (N_13460,N_11703,N_11418);
nor U13461 (N_13461,N_11800,N_12107);
nor U13462 (N_13462,N_10652,N_10535);
xnor U13463 (N_13463,N_10727,N_10650);
or U13464 (N_13464,N_12443,N_10002);
and U13465 (N_13465,N_10206,N_10353);
nand U13466 (N_13466,N_10386,N_11063);
or U13467 (N_13467,N_10607,N_11982);
nor U13468 (N_13468,N_11072,N_12156);
nor U13469 (N_13469,N_10404,N_12066);
and U13470 (N_13470,N_11770,N_11877);
nand U13471 (N_13471,N_10686,N_10001);
nand U13472 (N_13472,N_12490,N_10398);
nand U13473 (N_13473,N_11680,N_10546);
nand U13474 (N_13474,N_10237,N_10436);
nand U13475 (N_13475,N_11922,N_10071);
or U13476 (N_13476,N_10725,N_10159);
and U13477 (N_13477,N_12344,N_12453);
and U13478 (N_13478,N_12439,N_11224);
nor U13479 (N_13479,N_10259,N_11247);
nand U13480 (N_13480,N_11293,N_10960);
and U13481 (N_13481,N_10912,N_10730);
nand U13482 (N_13482,N_10618,N_12072);
nand U13483 (N_13483,N_10078,N_10427);
or U13484 (N_13484,N_10467,N_11756);
and U13485 (N_13485,N_10343,N_11064);
nor U13486 (N_13486,N_11070,N_10144);
nand U13487 (N_13487,N_12290,N_12086);
and U13488 (N_13488,N_12168,N_10820);
and U13489 (N_13489,N_11225,N_10366);
nand U13490 (N_13490,N_11616,N_12263);
or U13491 (N_13491,N_10608,N_11952);
nor U13492 (N_13492,N_10964,N_10690);
nand U13493 (N_13493,N_12129,N_11938);
nor U13494 (N_13494,N_10521,N_12274);
nand U13495 (N_13495,N_10252,N_10951);
nand U13496 (N_13496,N_11869,N_10396);
or U13497 (N_13497,N_12260,N_10869);
and U13498 (N_13498,N_12388,N_10468);
and U13499 (N_13499,N_11353,N_10179);
nand U13500 (N_13500,N_11695,N_11937);
and U13501 (N_13501,N_10486,N_10269);
or U13502 (N_13502,N_11255,N_11817);
and U13503 (N_13503,N_10885,N_10752);
or U13504 (N_13504,N_12113,N_11582);
and U13505 (N_13505,N_10736,N_11331);
nor U13506 (N_13506,N_10201,N_10724);
nand U13507 (N_13507,N_10975,N_12024);
nand U13508 (N_13508,N_11587,N_11432);
and U13509 (N_13509,N_11547,N_12008);
or U13510 (N_13510,N_11167,N_10371);
nand U13511 (N_13511,N_10147,N_11266);
and U13512 (N_13512,N_10805,N_11622);
nand U13513 (N_13513,N_10720,N_10783);
nor U13514 (N_13514,N_11062,N_11219);
nand U13515 (N_13515,N_11862,N_11299);
nand U13516 (N_13516,N_12271,N_12438);
and U13517 (N_13517,N_12473,N_11075);
or U13518 (N_13518,N_12080,N_11248);
and U13519 (N_13519,N_11766,N_11923);
or U13520 (N_13520,N_11262,N_11022);
nand U13521 (N_13521,N_10746,N_10836);
or U13522 (N_13522,N_10799,N_11903);
or U13523 (N_13523,N_11345,N_10046);
nor U13524 (N_13524,N_10320,N_11127);
nor U13525 (N_13525,N_11726,N_12233);
nand U13526 (N_13526,N_10930,N_10769);
nand U13527 (N_13527,N_12179,N_11973);
and U13528 (N_13528,N_12108,N_11990);
nand U13529 (N_13529,N_10051,N_11900);
nand U13530 (N_13530,N_10849,N_11272);
or U13531 (N_13531,N_10288,N_11530);
nand U13532 (N_13532,N_10266,N_11196);
and U13533 (N_13533,N_10450,N_10530);
or U13534 (N_13534,N_10915,N_11321);
nor U13535 (N_13535,N_12335,N_10414);
nor U13536 (N_13536,N_10616,N_11560);
or U13537 (N_13537,N_11624,N_11918);
and U13538 (N_13538,N_10297,N_11153);
or U13539 (N_13539,N_10186,N_10655);
nor U13540 (N_13540,N_11898,N_12036);
and U13541 (N_13541,N_10868,N_11433);
and U13542 (N_13542,N_11236,N_10513);
and U13543 (N_13543,N_11561,N_11323);
or U13544 (N_13544,N_10890,N_11140);
nand U13545 (N_13545,N_12250,N_11291);
nor U13546 (N_13546,N_11578,N_11831);
nor U13547 (N_13547,N_11382,N_10441);
nor U13548 (N_13548,N_10228,N_10895);
nor U13549 (N_13549,N_11401,N_11717);
nor U13550 (N_13550,N_10337,N_10796);
or U13551 (N_13551,N_11910,N_12374);
xnor U13552 (N_13552,N_11840,N_10247);
nor U13553 (N_13553,N_11081,N_12212);
nor U13554 (N_13554,N_11998,N_11508);
nor U13555 (N_13555,N_11947,N_11697);
nand U13556 (N_13556,N_10988,N_10167);
and U13557 (N_13557,N_10995,N_12452);
nand U13558 (N_13558,N_10350,N_12359);
or U13559 (N_13559,N_11659,N_11324);
or U13560 (N_13560,N_12298,N_10221);
or U13561 (N_13561,N_10150,N_12201);
nor U13562 (N_13562,N_11185,N_11069);
nand U13563 (N_13563,N_10620,N_12006);
or U13564 (N_13564,N_10210,N_11205);
and U13565 (N_13565,N_10688,N_10083);
or U13566 (N_13566,N_11309,N_11155);
nand U13567 (N_13567,N_10113,N_11308);
and U13568 (N_13568,N_10384,N_11755);
or U13569 (N_13569,N_11788,N_10341);
nor U13570 (N_13570,N_11312,N_12414);
or U13571 (N_13571,N_10278,N_10529);
or U13572 (N_13572,N_12032,N_11603);
xor U13573 (N_13573,N_11052,N_11373);
or U13574 (N_13574,N_10250,N_11965);
or U13575 (N_13575,N_10662,N_11005);
nor U13576 (N_13576,N_10022,N_12029);
or U13577 (N_13577,N_11524,N_11245);
nand U13578 (N_13578,N_11145,N_11514);
nor U13579 (N_13579,N_10550,N_12321);
nand U13580 (N_13580,N_10716,N_11904);
nor U13581 (N_13581,N_11702,N_12092);
nor U13582 (N_13582,N_12166,N_11804);
nand U13583 (N_13583,N_10028,N_10454);
or U13584 (N_13584,N_11742,N_11759);
and U13585 (N_13585,N_10152,N_11868);
nor U13586 (N_13586,N_10220,N_11569);
nor U13587 (N_13587,N_10218,N_11855);
nor U13588 (N_13588,N_11558,N_11513);
nand U13589 (N_13589,N_12411,N_12496);
or U13590 (N_13590,N_10410,N_11633);
nand U13591 (N_13591,N_11124,N_12071);
nand U13592 (N_13592,N_10522,N_10222);
nand U13593 (N_13593,N_12079,N_12278);
and U13594 (N_13594,N_10560,N_10015);
and U13595 (N_13595,N_12130,N_10361);
nand U13596 (N_13596,N_11480,N_10865);
nand U13597 (N_13597,N_11764,N_12375);
or U13598 (N_13598,N_10338,N_10811);
nor U13599 (N_13599,N_10292,N_12376);
or U13600 (N_13600,N_10896,N_10695);
xor U13601 (N_13601,N_12480,N_11728);
nor U13602 (N_13602,N_11441,N_10464);
and U13603 (N_13603,N_11507,N_11667);
nor U13604 (N_13604,N_10192,N_11767);
or U13605 (N_13605,N_10126,N_12195);
xor U13606 (N_13606,N_10323,N_12122);
and U13607 (N_13607,N_10701,N_10784);
and U13608 (N_13608,N_10378,N_10056);
nand U13609 (N_13609,N_11541,N_10363);
nor U13610 (N_13610,N_10490,N_10480);
and U13611 (N_13611,N_10659,N_12461);
nor U13612 (N_13612,N_11522,N_11015);
or U13613 (N_13613,N_11625,N_10388);
nor U13614 (N_13614,N_11173,N_11708);
or U13615 (N_13615,N_11725,N_10539);
nand U13616 (N_13616,N_12405,N_11408);
or U13617 (N_13617,N_11057,N_11597);
and U13618 (N_13618,N_11083,N_10552);
and U13619 (N_13619,N_11102,N_12237);
nor U13620 (N_13620,N_10048,N_12396);
nand U13621 (N_13621,N_10949,N_12249);
xor U13622 (N_13622,N_12052,N_12484);
or U13623 (N_13623,N_12295,N_10321);
nor U13624 (N_13624,N_10674,N_12182);
and U13625 (N_13625,N_10129,N_10342);
and U13626 (N_13626,N_10105,N_11925);
nor U13627 (N_13627,N_11945,N_10547);
and U13628 (N_13628,N_11477,N_12285);
or U13629 (N_13629,N_11060,N_10516);
or U13630 (N_13630,N_12096,N_10442);
and U13631 (N_13631,N_10628,N_11687);
and U13632 (N_13632,N_11512,N_11133);
nor U13633 (N_13633,N_11557,N_10590);
nor U13634 (N_13634,N_10234,N_10747);
xor U13635 (N_13635,N_11301,N_10188);
nor U13636 (N_13636,N_11827,N_10282);
and U13637 (N_13637,N_10640,N_11720);
and U13638 (N_13638,N_10190,N_11919);
nand U13639 (N_13639,N_11690,N_11375);
and U13640 (N_13640,N_11761,N_11984);
nand U13641 (N_13641,N_11824,N_10393);
and U13642 (N_13642,N_11178,N_10841);
nor U13643 (N_13643,N_11239,N_11553);
or U13644 (N_13644,N_12085,N_10170);
and U13645 (N_13645,N_10489,N_11931);
nand U13646 (N_13646,N_11190,N_11917);
and U13647 (N_13647,N_11573,N_11878);
or U13648 (N_13648,N_12146,N_12010);
and U13649 (N_13649,N_12297,N_11842);
nor U13650 (N_13650,N_11203,N_10979);
nor U13651 (N_13651,N_10360,N_12230);
and U13652 (N_13652,N_12203,N_12106);
and U13653 (N_13653,N_12135,N_11491);
nand U13654 (N_13654,N_11351,N_10593);
nor U13655 (N_13655,N_11916,N_11442);
nand U13656 (N_13656,N_12205,N_11485);
xor U13657 (N_13657,N_10670,N_12435);
and U13658 (N_13658,N_10161,N_11941);
xnor U13659 (N_13659,N_12172,N_10672);
nor U13660 (N_13660,N_12088,N_11985);
nand U13661 (N_13661,N_11596,N_11499);
nand U13662 (N_13662,N_11497,N_12077);
nand U13663 (N_13663,N_11518,N_11087);
and U13664 (N_13664,N_10668,N_10175);
and U13665 (N_13665,N_12304,N_11853);
or U13666 (N_13666,N_10824,N_10713);
and U13667 (N_13667,N_12423,N_12159);
nand U13668 (N_13668,N_11619,N_10714);
nand U13669 (N_13669,N_12337,N_10613);
nand U13670 (N_13670,N_11565,N_10968);
or U13671 (N_13671,N_10143,N_10060);
nor U13672 (N_13672,N_11808,N_12273);
nor U13673 (N_13673,N_11054,N_10943);
and U13674 (N_13674,N_12025,N_10833);
and U13675 (N_13675,N_10623,N_12363);
nand U13676 (N_13676,N_10063,N_10077);
and U13677 (N_13677,N_11208,N_11162);
nor U13678 (N_13678,N_11866,N_10808);
xor U13679 (N_13679,N_11232,N_12178);
and U13680 (N_13680,N_11238,N_11816);
nand U13681 (N_13681,N_10329,N_10488);
nand U13682 (N_13682,N_10582,N_12094);
or U13683 (N_13683,N_10503,N_10013);
nand U13684 (N_13684,N_12120,N_12314);
nor U13685 (N_13685,N_11177,N_10241);
and U13686 (N_13686,N_12289,N_12286);
or U13687 (N_13687,N_11424,N_12497);
nor U13688 (N_13688,N_11329,N_10369);
nor U13689 (N_13689,N_10621,N_10195);
or U13690 (N_13690,N_11710,N_11724);
nor U13691 (N_13691,N_10010,N_11261);
and U13692 (N_13692,N_11030,N_11141);
xnor U13693 (N_13693,N_11361,N_11414);
nand U13694 (N_13694,N_11362,N_12002);
nand U13695 (N_13695,N_10643,N_11526);
nand U13696 (N_13696,N_12471,N_11661);
xnor U13697 (N_13697,N_11981,N_10866);
nand U13698 (N_13698,N_10644,N_10908);
xor U13699 (N_13699,N_11791,N_11483);
or U13700 (N_13700,N_11601,N_10313);
xnor U13701 (N_13701,N_10253,N_11383);
nand U13702 (N_13702,N_11168,N_11269);
nand U13703 (N_13703,N_10759,N_11642);
xor U13704 (N_13704,N_10019,N_11701);
nor U13705 (N_13705,N_12239,N_10267);
nor U13706 (N_13706,N_11651,N_10815);
and U13707 (N_13707,N_10506,N_11330);
nor U13708 (N_13708,N_11144,N_12449);
nand U13709 (N_13709,N_11586,N_11683);
nand U13710 (N_13710,N_11718,N_10107);
and U13711 (N_13711,N_11885,N_11122);
and U13712 (N_13712,N_11545,N_11721);
xnor U13713 (N_13713,N_10827,N_10657);
or U13714 (N_13714,N_10331,N_11496);
xnor U13715 (N_13715,N_11806,N_10687);
nor U13716 (N_13716,N_11461,N_10098);
nor U13717 (N_13717,N_11995,N_12031);
nor U13718 (N_13718,N_11849,N_12292);
or U13719 (N_13719,N_11187,N_11055);
or U13720 (N_13720,N_12261,N_10132);
or U13721 (N_13721,N_10137,N_12082);
nand U13722 (N_13722,N_12013,N_11484);
nand U13723 (N_13723,N_12214,N_12161);
nor U13724 (N_13724,N_10965,N_10753);
nor U13725 (N_13725,N_11000,N_12323);
nand U13726 (N_13726,N_10298,N_11567);
and U13727 (N_13727,N_12217,N_11857);
nor U13728 (N_13728,N_11749,N_11088);
or U13729 (N_13729,N_10947,N_12486);
nor U13730 (N_13730,N_10364,N_12406);
or U13731 (N_13731,N_11047,N_11551);
and U13732 (N_13732,N_11584,N_11074);
or U13733 (N_13733,N_12114,N_10505);
nor U13734 (N_13734,N_11280,N_10782);
nor U13735 (N_13735,N_10422,N_10624);
or U13736 (N_13736,N_12384,N_11482);
or U13737 (N_13737,N_12272,N_11969);
nor U13738 (N_13738,N_12028,N_11882);
and U13739 (N_13739,N_12213,N_10120);
nor U13740 (N_13740,N_11859,N_10014);
and U13741 (N_13741,N_11119,N_12091);
or U13742 (N_13742,N_11306,N_12062);
nand U13743 (N_13743,N_10952,N_12371);
nand U13744 (N_13744,N_12110,N_10523);
and U13745 (N_13745,N_10041,N_11572);
and U13746 (N_13746,N_11979,N_11722);
and U13747 (N_13747,N_11852,N_12340);
nand U13748 (N_13748,N_10219,N_12259);
and U13749 (N_13749,N_12450,N_10813);
nor U13750 (N_13750,N_11039,N_10259);
nand U13751 (N_13751,N_11492,N_10046);
nor U13752 (N_13752,N_11742,N_10545);
or U13753 (N_13753,N_10561,N_11694);
nor U13754 (N_13754,N_10817,N_11515);
nand U13755 (N_13755,N_10163,N_10753);
or U13756 (N_13756,N_11778,N_11373);
or U13757 (N_13757,N_12471,N_11913);
or U13758 (N_13758,N_10118,N_11870);
nor U13759 (N_13759,N_11219,N_11086);
and U13760 (N_13760,N_11784,N_11662);
or U13761 (N_13761,N_12098,N_11150);
nand U13762 (N_13762,N_11333,N_10155);
nor U13763 (N_13763,N_10441,N_11837);
nand U13764 (N_13764,N_10184,N_10221);
nand U13765 (N_13765,N_11810,N_11708);
nor U13766 (N_13766,N_11211,N_10088);
nand U13767 (N_13767,N_12126,N_11134);
and U13768 (N_13768,N_11554,N_10435);
nor U13769 (N_13769,N_11607,N_10429);
nand U13770 (N_13770,N_10441,N_11840);
and U13771 (N_13771,N_10320,N_11906);
or U13772 (N_13772,N_11084,N_10696);
nor U13773 (N_13773,N_11100,N_12282);
nand U13774 (N_13774,N_11744,N_11053);
and U13775 (N_13775,N_10561,N_11872);
nand U13776 (N_13776,N_10286,N_10981);
or U13777 (N_13777,N_10679,N_11028);
nor U13778 (N_13778,N_11316,N_11784);
and U13779 (N_13779,N_12461,N_10620);
nand U13780 (N_13780,N_11962,N_11412);
or U13781 (N_13781,N_10856,N_10002);
or U13782 (N_13782,N_12141,N_10750);
and U13783 (N_13783,N_11333,N_10120);
nand U13784 (N_13784,N_12398,N_11066);
and U13785 (N_13785,N_11844,N_10524);
or U13786 (N_13786,N_10965,N_11438);
nand U13787 (N_13787,N_10650,N_10723);
or U13788 (N_13788,N_11151,N_11400);
or U13789 (N_13789,N_11113,N_10429);
and U13790 (N_13790,N_11979,N_10611);
or U13791 (N_13791,N_10576,N_10348);
or U13792 (N_13792,N_11064,N_11580);
xnor U13793 (N_13793,N_11320,N_10905);
or U13794 (N_13794,N_10872,N_10436);
nand U13795 (N_13795,N_11519,N_10611);
and U13796 (N_13796,N_10360,N_10308);
or U13797 (N_13797,N_12006,N_11597);
and U13798 (N_13798,N_10294,N_12249);
or U13799 (N_13799,N_11259,N_10091);
or U13800 (N_13800,N_10422,N_11989);
nor U13801 (N_13801,N_11846,N_10952);
and U13802 (N_13802,N_10080,N_11668);
nor U13803 (N_13803,N_12182,N_11487);
or U13804 (N_13804,N_12073,N_10339);
nor U13805 (N_13805,N_10473,N_12014);
nor U13806 (N_13806,N_10070,N_11738);
and U13807 (N_13807,N_12382,N_11424);
nor U13808 (N_13808,N_12198,N_10183);
or U13809 (N_13809,N_10785,N_12204);
or U13810 (N_13810,N_12071,N_11354);
xnor U13811 (N_13811,N_12313,N_10417);
nor U13812 (N_13812,N_12152,N_10378);
nand U13813 (N_13813,N_10456,N_10293);
and U13814 (N_13814,N_10116,N_12213);
and U13815 (N_13815,N_12244,N_12083);
or U13816 (N_13816,N_11842,N_12082);
and U13817 (N_13817,N_10228,N_10062);
nand U13818 (N_13818,N_12017,N_12147);
and U13819 (N_13819,N_10058,N_11960);
or U13820 (N_13820,N_10944,N_10945);
or U13821 (N_13821,N_10700,N_11581);
nor U13822 (N_13822,N_10489,N_10335);
and U13823 (N_13823,N_11741,N_10033);
and U13824 (N_13824,N_12140,N_11245);
and U13825 (N_13825,N_12402,N_11901);
and U13826 (N_13826,N_10031,N_10294);
nand U13827 (N_13827,N_12103,N_10591);
nor U13828 (N_13828,N_10556,N_10565);
nand U13829 (N_13829,N_10038,N_12313);
or U13830 (N_13830,N_12151,N_12304);
or U13831 (N_13831,N_11080,N_10585);
nor U13832 (N_13832,N_11492,N_11698);
xor U13833 (N_13833,N_10415,N_11637);
nand U13834 (N_13834,N_11651,N_11824);
nor U13835 (N_13835,N_11184,N_10946);
nor U13836 (N_13836,N_11267,N_11304);
xnor U13837 (N_13837,N_10115,N_10553);
nand U13838 (N_13838,N_11714,N_11854);
nor U13839 (N_13839,N_11045,N_10584);
nand U13840 (N_13840,N_12400,N_12056);
nor U13841 (N_13841,N_11319,N_11167);
and U13842 (N_13842,N_10721,N_10681);
nand U13843 (N_13843,N_10803,N_11766);
and U13844 (N_13844,N_12236,N_11540);
nor U13845 (N_13845,N_11385,N_10258);
and U13846 (N_13846,N_12342,N_12438);
or U13847 (N_13847,N_11316,N_10409);
xnor U13848 (N_13848,N_11815,N_11056);
and U13849 (N_13849,N_11288,N_12248);
nand U13850 (N_13850,N_11643,N_11368);
nor U13851 (N_13851,N_12491,N_12019);
nand U13852 (N_13852,N_11099,N_10911);
nor U13853 (N_13853,N_10461,N_11436);
nor U13854 (N_13854,N_10275,N_11950);
nor U13855 (N_13855,N_11939,N_11658);
or U13856 (N_13856,N_10764,N_12247);
nor U13857 (N_13857,N_11385,N_11502);
and U13858 (N_13858,N_10923,N_10548);
nor U13859 (N_13859,N_10288,N_12368);
or U13860 (N_13860,N_11089,N_10495);
nand U13861 (N_13861,N_12113,N_11942);
nor U13862 (N_13862,N_10366,N_12068);
and U13863 (N_13863,N_11706,N_10775);
nor U13864 (N_13864,N_11311,N_10831);
nand U13865 (N_13865,N_10599,N_11336);
or U13866 (N_13866,N_12308,N_10722);
and U13867 (N_13867,N_10738,N_12286);
nand U13868 (N_13868,N_11539,N_10918);
and U13869 (N_13869,N_11900,N_11200);
nand U13870 (N_13870,N_11801,N_10424);
nor U13871 (N_13871,N_11540,N_10687);
or U13872 (N_13872,N_11565,N_10383);
or U13873 (N_13873,N_12018,N_12419);
or U13874 (N_13874,N_11623,N_12492);
or U13875 (N_13875,N_12255,N_11934);
nor U13876 (N_13876,N_12119,N_10678);
and U13877 (N_13877,N_10286,N_10033);
nand U13878 (N_13878,N_10835,N_11057);
nor U13879 (N_13879,N_10776,N_10370);
and U13880 (N_13880,N_11132,N_11431);
nand U13881 (N_13881,N_10971,N_11222);
and U13882 (N_13882,N_10064,N_11124);
nand U13883 (N_13883,N_10399,N_10668);
nand U13884 (N_13884,N_11299,N_10072);
or U13885 (N_13885,N_11114,N_10760);
and U13886 (N_13886,N_11321,N_12247);
nor U13887 (N_13887,N_10309,N_10242);
nand U13888 (N_13888,N_12487,N_10749);
or U13889 (N_13889,N_12406,N_11033);
and U13890 (N_13890,N_11705,N_10448);
xor U13891 (N_13891,N_10016,N_10607);
or U13892 (N_13892,N_11186,N_12350);
nor U13893 (N_13893,N_10492,N_12208);
and U13894 (N_13894,N_11224,N_10132);
nand U13895 (N_13895,N_10876,N_12041);
and U13896 (N_13896,N_10020,N_11472);
and U13897 (N_13897,N_12298,N_10317);
nand U13898 (N_13898,N_11568,N_10086);
xnor U13899 (N_13899,N_10807,N_10988);
nand U13900 (N_13900,N_11698,N_10062);
or U13901 (N_13901,N_10449,N_11274);
nand U13902 (N_13902,N_11853,N_10994);
nor U13903 (N_13903,N_12156,N_11976);
or U13904 (N_13904,N_11300,N_10787);
or U13905 (N_13905,N_10772,N_10942);
or U13906 (N_13906,N_10665,N_10893);
nand U13907 (N_13907,N_11259,N_10265);
nor U13908 (N_13908,N_10297,N_10546);
nor U13909 (N_13909,N_12097,N_11107);
and U13910 (N_13910,N_10080,N_11860);
nor U13911 (N_13911,N_10123,N_10756);
nand U13912 (N_13912,N_11254,N_10870);
nor U13913 (N_13913,N_11485,N_10894);
nand U13914 (N_13914,N_12078,N_11130);
nor U13915 (N_13915,N_11920,N_11589);
and U13916 (N_13916,N_10265,N_11053);
or U13917 (N_13917,N_11266,N_12395);
or U13918 (N_13918,N_12205,N_11944);
or U13919 (N_13919,N_10358,N_10122);
nand U13920 (N_13920,N_11639,N_10203);
and U13921 (N_13921,N_11589,N_12489);
and U13922 (N_13922,N_10077,N_10229);
or U13923 (N_13923,N_10826,N_10721);
or U13924 (N_13924,N_11696,N_11462);
and U13925 (N_13925,N_11225,N_11687);
and U13926 (N_13926,N_12369,N_11732);
nand U13927 (N_13927,N_10907,N_10970);
and U13928 (N_13928,N_12489,N_10302);
or U13929 (N_13929,N_11838,N_11627);
and U13930 (N_13930,N_11691,N_10810);
and U13931 (N_13931,N_10735,N_10365);
nand U13932 (N_13932,N_11671,N_11628);
nand U13933 (N_13933,N_12040,N_10971);
and U13934 (N_13934,N_11244,N_12034);
and U13935 (N_13935,N_11411,N_10953);
nor U13936 (N_13936,N_11939,N_10038);
and U13937 (N_13937,N_11376,N_10597);
and U13938 (N_13938,N_10191,N_11579);
nand U13939 (N_13939,N_11152,N_11857);
or U13940 (N_13940,N_10918,N_10440);
nor U13941 (N_13941,N_12242,N_10013);
nor U13942 (N_13942,N_11123,N_11494);
and U13943 (N_13943,N_12125,N_11602);
nor U13944 (N_13944,N_11758,N_10938);
nand U13945 (N_13945,N_11260,N_12229);
nand U13946 (N_13946,N_12237,N_11391);
and U13947 (N_13947,N_12392,N_10559);
and U13948 (N_13948,N_10300,N_11884);
nor U13949 (N_13949,N_10405,N_11050);
and U13950 (N_13950,N_11052,N_11700);
and U13951 (N_13951,N_12065,N_11071);
nor U13952 (N_13952,N_11515,N_10899);
nand U13953 (N_13953,N_10692,N_12464);
or U13954 (N_13954,N_10753,N_11801);
xor U13955 (N_13955,N_10734,N_10958);
nand U13956 (N_13956,N_11815,N_12343);
nand U13957 (N_13957,N_12389,N_11838);
nor U13958 (N_13958,N_12339,N_12413);
and U13959 (N_13959,N_12247,N_11924);
nand U13960 (N_13960,N_11434,N_11338);
nand U13961 (N_13961,N_11671,N_10936);
and U13962 (N_13962,N_10346,N_10730);
or U13963 (N_13963,N_10286,N_12103);
nand U13964 (N_13964,N_11655,N_12017);
nand U13965 (N_13965,N_11834,N_10469);
nand U13966 (N_13966,N_10076,N_11346);
nor U13967 (N_13967,N_12193,N_12146);
nand U13968 (N_13968,N_11641,N_12143);
and U13969 (N_13969,N_10320,N_11522);
nand U13970 (N_13970,N_10850,N_11838);
nor U13971 (N_13971,N_10083,N_11381);
and U13972 (N_13972,N_10001,N_12060);
or U13973 (N_13973,N_12214,N_11353);
and U13974 (N_13974,N_12227,N_10824);
nor U13975 (N_13975,N_11658,N_11507);
nand U13976 (N_13976,N_11692,N_11175);
or U13977 (N_13977,N_11982,N_12193);
or U13978 (N_13978,N_11676,N_11246);
and U13979 (N_13979,N_11112,N_11442);
nand U13980 (N_13980,N_10472,N_11739);
nand U13981 (N_13981,N_11004,N_10428);
nand U13982 (N_13982,N_12160,N_11326);
xnor U13983 (N_13983,N_10773,N_10180);
nor U13984 (N_13984,N_10952,N_10424);
and U13985 (N_13985,N_12483,N_11021);
nor U13986 (N_13986,N_11719,N_11430);
and U13987 (N_13987,N_12093,N_12316);
and U13988 (N_13988,N_11269,N_10348);
or U13989 (N_13989,N_10024,N_10006);
nand U13990 (N_13990,N_11568,N_11677);
or U13991 (N_13991,N_12008,N_10995);
or U13992 (N_13992,N_12057,N_11462);
or U13993 (N_13993,N_10327,N_11352);
xnor U13994 (N_13994,N_10929,N_12055);
nor U13995 (N_13995,N_11663,N_10273);
nor U13996 (N_13996,N_10739,N_11800);
nor U13997 (N_13997,N_10428,N_11963);
or U13998 (N_13998,N_10250,N_11975);
nor U13999 (N_13999,N_11433,N_10143);
nor U14000 (N_14000,N_11971,N_10985);
nand U14001 (N_14001,N_11865,N_12464);
nand U14002 (N_14002,N_12184,N_12413);
nand U14003 (N_14003,N_10149,N_10999);
nor U14004 (N_14004,N_11860,N_10568);
nor U14005 (N_14005,N_11220,N_12492);
xor U14006 (N_14006,N_11109,N_10503);
or U14007 (N_14007,N_12102,N_11223);
nand U14008 (N_14008,N_11557,N_12332);
nand U14009 (N_14009,N_12329,N_10658);
xor U14010 (N_14010,N_11359,N_12073);
nor U14011 (N_14011,N_10764,N_12281);
nand U14012 (N_14012,N_10459,N_11184);
nand U14013 (N_14013,N_10428,N_12023);
nor U14014 (N_14014,N_11384,N_12499);
and U14015 (N_14015,N_11748,N_10340);
and U14016 (N_14016,N_11465,N_10557);
or U14017 (N_14017,N_10215,N_11306);
nand U14018 (N_14018,N_12215,N_11109);
nor U14019 (N_14019,N_11056,N_11005);
nor U14020 (N_14020,N_10750,N_10443);
nor U14021 (N_14021,N_11896,N_11639);
and U14022 (N_14022,N_10779,N_10319);
and U14023 (N_14023,N_10968,N_10810);
or U14024 (N_14024,N_10175,N_12363);
or U14025 (N_14025,N_12293,N_11007);
nor U14026 (N_14026,N_10465,N_10020);
nor U14027 (N_14027,N_11821,N_11440);
or U14028 (N_14028,N_10589,N_10220);
nor U14029 (N_14029,N_10274,N_10419);
or U14030 (N_14030,N_11405,N_11506);
nand U14031 (N_14031,N_11524,N_10277);
and U14032 (N_14032,N_12140,N_11448);
nor U14033 (N_14033,N_12264,N_11077);
or U14034 (N_14034,N_12140,N_11088);
or U14035 (N_14035,N_10388,N_11206);
nand U14036 (N_14036,N_10288,N_11246);
and U14037 (N_14037,N_12141,N_11321);
and U14038 (N_14038,N_12475,N_10290);
nand U14039 (N_14039,N_10313,N_10125);
nand U14040 (N_14040,N_10110,N_11284);
or U14041 (N_14041,N_10363,N_10366);
nor U14042 (N_14042,N_11750,N_12245);
nor U14043 (N_14043,N_12076,N_10139);
or U14044 (N_14044,N_11903,N_11126);
or U14045 (N_14045,N_12388,N_12270);
nand U14046 (N_14046,N_10178,N_10773);
and U14047 (N_14047,N_11273,N_12390);
and U14048 (N_14048,N_12063,N_10372);
nand U14049 (N_14049,N_10196,N_10505);
and U14050 (N_14050,N_10802,N_10381);
and U14051 (N_14051,N_12434,N_10262);
nor U14052 (N_14052,N_11531,N_10577);
nand U14053 (N_14053,N_10468,N_11067);
or U14054 (N_14054,N_10720,N_10658);
nor U14055 (N_14055,N_12180,N_11837);
nor U14056 (N_14056,N_12485,N_11271);
or U14057 (N_14057,N_11493,N_10043);
and U14058 (N_14058,N_12173,N_12005);
or U14059 (N_14059,N_10604,N_12415);
nor U14060 (N_14060,N_10531,N_11026);
and U14061 (N_14061,N_12194,N_11821);
nor U14062 (N_14062,N_12002,N_12149);
nor U14063 (N_14063,N_10224,N_10119);
xnor U14064 (N_14064,N_10198,N_12189);
nand U14065 (N_14065,N_10809,N_10981);
nor U14066 (N_14066,N_10956,N_11042);
nor U14067 (N_14067,N_10495,N_12385);
and U14068 (N_14068,N_11555,N_11952);
and U14069 (N_14069,N_11148,N_10851);
nor U14070 (N_14070,N_11586,N_10372);
nor U14071 (N_14071,N_10706,N_12328);
nor U14072 (N_14072,N_11620,N_10038);
and U14073 (N_14073,N_10814,N_10021);
or U14074 (N_14074,N_10455,N_10462);
nor U14075 (N_14075,N_11957,N_11765);
nor U14076 (N_14076,N_11066,N_10826);
nor U14077 (N_14077,N_12453,N_11615);
nor U14078 (N_14078,N_11729,N_11422);
and U14079 (N_14079,N_10867,N_11788);
and U14080 (N_14080,N_11623,N_12196);
xnor U14081 (N_14081,N_11488,N_10553);
nor U14082 (N_14082,N_11563,N_11420);
nor U14083 (N_14083,N_12209,N_10966);
nand U14084 (N_14084,N_11625,N_12439);
or U14085 (N_14085,N_11455,N_10558);
nand U14086 (N_14086,N_11033,N_12022);
nand U14087 (N_14087,N_12473,N_12032);
and U14088 (N_14088,N_11169,N_11870);
and U14089 (N_14089,N_11605,N_10316);
or U14090 (N_14090,N_10183,N_11689);
or U14091 (N_14091,N_11036,N_10682);
nand U14092 (N_14092,N_12176,N_10671);
nor U14093 (N_14093,N_10704,N_10849);
nor U14094 (N_14094,N_10889,N_10583);
or U14095 (N_14095,N_11846,N_11982);
nor U14096 (N_14096,N_12049,N_11625);
nor U14097 (N_14097,N_11420,N_11711);
nand U14098 (N_14098,N_12063,N_11270);
nand U14099 (N_14099,N_10654,N_11080);
and U14100 (N_14100,N_11954,N_10645);
or U14101 (N_14101,N_11970,N_11186);
nor U14102 (N_14102,N_10288,N_10226);
nand U14103 (N_14103,N_10099,N_10966);
nand U14104 (N_14104,N_11204,N_11690);
nand U14105 (N_14105,N_11683,N_11029);
or U14106 (N_14106,N_12347,N_10907);
nor U14107 (N_14107,N_11771,N_10587);
or U14108 (N_14108,N_12098,N_10091);
nor U14109 (N_14109,N_10154,N_11271);
and U14110 (N_14110,N_11112,N_12478);
nor U14111 (N_14111,N_10590,N_10711);
nor U14112 (N_14112,N_11947,N_12278);
nand U14113 (N_14113,N_11971,N_11477);
or U14114 (N_14114,N_12254,N_11887);
or U14115 (N_14115,N_11549,N_11037);
and U14116 (N_14116,N_12120,N_10454);
nand U14117 (N_14117,N_10710,N_11928);
and U14118 (N_14118,N_12445,N_11371);
nand U14119 (N_14119,N_10690,N_12394);
nand U14120 (N_14120,N_10747,N_10322);
nand U14121 (N_14121,N_10547,N_10787);
nand U14122 (N_14122,N_10476,N_10324);
nor U14123 (N_14123,N_10028,N_12495);
nand U14124 (N_14124,N_12084,N_11106);
or U14125 (N_14125,N_10032,N_12116);
nand U14126 (N_14126,N_11648,N_10080);
nand U14127 (N_14127,N_10146,N_11888);
and U14128 (N_14128,N_11107,N_10925);
or U14129 (N_14129,N_10942,N_10926);
and U14130 (N_14130,N_11810,N_11860);
and U14131 (N_14131,N_12308,N_12257);
nand U14132 (N_14132,N_11340,N_11509);
and U14133 (N_14133,N_10446,N_11234);
nand U14134 (N_14134,N_10657,N_12326);
or U14135 (N_14135,N_10102,N_11022);
nand U14136 (N_14136,N_10992,N_11526);
or U14137 (N_14137,N_11872,N_11618);
nor U14138 (N_14138,N_10523,N_11680);
nor U14139 (N_14139,N_11240,N_11986);
and U14140 (N_14140,N_10355,N_10640);
nor U14141 (N_14141,N_11350,N_12179);
nor U14142 (N_14142,N_11903,N_12287);
nor U14143 (N_14143,N_10949,N_10256);
and U14144 (N_14144,N_12098,N_12470);
and U14145 (N_14145,N_11831,N_12262);
nand U14146 (N_14146,N_11699,N_11583);
and U14147 (N_14147,N_10270,N_11364);
or U14148 (N_14148,N_10745,N_11102);
and U14149 (N_14149,N_11403,N_11989);
and U14150 (N_14150,N_10435,N_10407);
nand U14151 (N_14151,N_10928,N_11778);
nor U14152 (N_14152,N_11030,N_12336);
nand U14153 (N_14153,N_10999,N_10996);
nand U14154 (N_14154,N_11338,N_11178);
and U14155 (N_14155,N_10063,N_10601);
xor U14156 (N_14156,N_12320,N_10404);
nor U14157 (N_14157,N_12169,N_10542);
nand U14158 (N_14158,N_12464,N_10321);
nand U14159 (N_14159,N_10316,N_10769);
nand U14160 (N_14160,N_10817,N_12064);
nor U14161 (N_14161,N_11610,N_11654);
nor U14162 (N_14162,N_11363,N_10953);
and U14163 (N_14163,N_12035,N_10089);
and U14164 (N_14164,N_10157,N_11084);
or U14165 (N_14165,N_10890,N_11771);
or U14166 (N_14166,N_11599,N_11909);
nor U14167 (N_14167,N_12098,N_11838);
nand U14168 (N_14168,N_11489,N_11923);
and U14169 (N_14169,N_12288,N_12165);
xnor U14170 (N_14170,N_10060,N_11153);
nand U14171 (N_14171,N_11397,N_11169);
or U14172 (N_14172,N_11277,N_10870);
or U14173 (N_14173,N_12120,N_11668);
xnor U14174 (N_14174,N_11652,N_11225);
or U14175 (N_14175,N_12111,N_10486);
nor U14176 (N_14176,N_11731,N_11766);
nand U14177 (N_14177,N_10063,N_11246);
nor U14178 (N_14178,N_11826,N_10792);
or U14179 (N_14179,N_12033,N_10630);
or U14180 (N_14180,N_10944,N_10194);
or U14181 (N_14181,N_10535,N_10698);
and U14182 (N_14182,N_11202,N_12118);
nor U14183 (N_14183,N_12079,N_11289);
nor U14184 (N_14184,N_10381,N_10618);
nor U14185 (N_14185,N_12262,N_12316);
and U14186 (N_14186,N_11461,N_10635);
nor U14187 (N_14187,N_11925,N_11457);
nand U14188 (N_14188,N_12315,N_10008);
nor U14189 (N_14189,N_12172,N_11729);
and U14190 (N_14190,N_10396,N_11559);
xor U14191 (N_14191,N_11562,N_11035);
and U14192 (N_14192,N_11758,N_11707);
nand U14193 (N_14193,N_12049,N_11961);
and U14194 (N_14194,N_11924,N_10358);
and U14195 (N_14195,N_11461,N_11472);
nand U14196 (N_14196,N_10939,N_10710);
nand U14197 (N_14197,N_11539,N_11096);
or U14198 (N_14198,N_11525,N_10292);
nor U14199 (N_14199,N_12157,N_10603);
nand U14200 (N_14200,N_11172,N_11396);
nor U14201 (N_14201,N_12368,N_10370);
or U14202 (N_14202,N_10480,N_11980);
or U14203 (N_14203,N_11421,N_10270);
or U14204 (N_14204,N_10953,N_11274);
xnor U14205 (N_14205,N_10081,N_10508);
and U14206 (N_14206,N_10875,N_12351);
or U14207 (N_14207,N_12323,N_10037);
and U14208 (N_14208,N_11384,N_10097);
nor U14209 (N_14209,N_10303,N_12486);
or U14210 (N_14210,N_11867,N_10897);
nor U14211 (N_14211,N_12464,N_11533);
nand U14212 (N_14212,N_12093,N_11933);
or U14213 (N_14213,N_11207,N_10746);
nand U14214 (N_14214,N_12438,N_11581);
or U14215 (N_14215,N_10803,N_11778);
nand U14216 (N_14216,N_12201,N_10972);
nor U14217 (N_14217,N_12192,N_11851);
nand U14218 (N_14218,N_10605,N_10347);
nand U14219 (N_14219,N_12125,N_12189);
or U14220 (N_14220,N_11012,N_12156);
or U14221 (N_14221,N_10782,N_11298);
nand U14222 (N_14222,N_10819,N_11205);
nor U14223 (N_14223,N_11057,N_10760);
or U14224 (N_14224,N_12132,N_11065);
and U14225 (N_14225,N_10585,N_10581);
or U14226 (N_14226,N_10296,N_11861);
nor U14227 (N_14227,N_12048,N_10468);
and U14228 (N_14228,N_11710,N_11683);
and U14229 (N_14229,N_10724,N_10055);
nor U14230 (N_14230,N_11492,N_12020);
nor U14231 (N_14231,N_11842,N_12189);
and U14232 (N_14232,N_11401,N_10493);
or U14233 (N_14233,N_12154,N_11635);
or U14234 (N_14234,N_12242,N_10238);
nor U14235 (N_14235,N_10349,N_12388);
and U14236 (N_14236,N_11663,N_11015);
xor U14237 (N_14237,N_12067,N_10504);
and U14238 (N_14238,N_10084,N_11662);
nand U14239 (N_14239,N_10341,N_10165);
or U14240 (N_14240,N_11855,N_11528);
or U14241 (N_14241,N_10748,N_11046);
nand U14242 (N_14242,N_10641,N_10650);
and U14243 (N_14243,N_11828,N_12036);
and U14244 (N_14244,N_12225,N_11866);
or U14245 (N_14245,N_10203,N_10020);
or U14246 (N_14246,N_10932,N_12339);
and U14247 (N_14247,N_10160,N_12430);
nor U14248 (N_14248,N_12045,N_11994);
nor U14249 (N_14249,N_11024,N_10997);
nor U14250 (N_14250,N_10066,N_10244);
and U14251 (N_14251,N_12032,N_11052);
or U14252 (N_14252,N_10045,N_11224);
xnor U14253 (N_14253,N_12160,N_11966);
nand U14254 (N_14254,N_11575,N_11030);
and U14255 (N_14255,N_10892,N_12379);
nor U14256 (N_14256,N_12066,N_10135);
xor U14257 (N_14257,N_11631,N_12406);
nand U14258 (N_14258,N_11237,N_12291);
and U14259 (N_14259,N_10124,N_11662);
and U14260 (N_14260,N_10943,N_11857);
and U14261 (N_14261,N_10681,N_10760);
or U14262 (N_14262,N_12369,N_11562);
or U14263 (N_14263,N_12157,N_10478);
and U14264 (N_14264,N_10736,N_11926);
nor U14265 (N_14265,N_11943,N_11648);
or U14266 (N_14266,N_12088,N_10200);
nor U14267 (N_14267,N_11627,N_11517);
or U14268 (N_14268,N_11065,N_11936);
or U14269 (N_14269,N_10160,N_12296);
and U14270 (N_14270,N_11497,N_10308);
nand U14271 (N_14271,N_10056,N_10887);
or U14272 (N_14272,N_11895,N_10815);
or U14273 (N_14273,N_12110,N_11963);
or U14274 (N_14274,N_11571,N_10508);
or U14275 (N_14275,N_11667,N_11819);
or U14276 (N_14276,N_10432,N_11661);
nand U14277 (N_14277,N_11440,N_11619);
nor U14278 (N_14278,N_11576,N_11733);
or U14279 (N_14279,N_12038,N_12213);
nor U14280 (N_14280,N_10132,N_11089);
nand U14281 (N_14281,N_12148,N_11447);
nand U14282 (N_14282,N_11182,N_11185);
nand U14283 (N_14283,N_10413,N_12306);
and U14284 (N_14284,N_10646,N_10073);
nor U14285 (N_14285,N_10848,N_11794);
nand U14286 (N_14286,N_12279,N_11450);
nor U14287 (N_14287,N_10064,N_12137);
and U14288 (N_14288,N_11846,N_11377);
xor U14289 (N_14289,N_10708,N_10173);
nand U14290 (N_14290,N_10133,N_10772);
nand U14291 (N_14291,N_12454,N_10753);
and U14292 (N_14292,N_10533,N_10011);
or U14293 (N_14293,N_10697,N_12182);
nand U14294 (N_14294,N_12484,N_11396);
nor U14295 (N_14295,N_10620,N_12005);
or U14296 (N_14296,N_11991,N_11309);
and U14297 (N_14297,N_11455,N_11767);
nand U14298 (N_14298,N_11152,N_12249);
and U14299 (N_14299,N_11829,N_11130);
nor U14300 (N_14300,N_10270,N_12350);
nand U14301 (N_14301,N_11864,N_12056);
nor U14302 (N_14302,N_10480,N_11863);
nand U14303 (N_14303,N_10535,N_10196);
xor U14304 (N_14304,N_10691,N_11738);
nand U14305 (N_14305,N_10517,N_10515);
and U14306 (N_14306,N_10185,N_11677);
or U14307 (N_14307,N_12175,N_11481);
or U14308 (N_14308,N_11578,N_10459);
or U14309 (N_14309,N_12263,N_12494);
and U14310 (N_14310,N_11875,N_11024);
and U14311 (N_14311,N_11366,N_12155);
nand U14312 (N_14312,N_11672,N_10715);
nor U14313 (N_14313,N_11679,N_10886);
nand U14314 (N_14314,N_12209,N_11787);
xor U14315 (N_14315,N_12115,N_11928);
nand U14316 (N_14316,N_11030,N_10573);
nand U14317 (N_14317,N_10772,N_11775);
nor U14318 (N_14318,N_10947,N_10802);
and U14319 (N_14319,N_11797,N_12027);
or U14320 (N_14320,N_11755,N_10531);
nand U14321 (N_14321,N_11499,N_10638);
nand U14322 (N_14322,N_11934,N_11644);
nor U14323 (N_14323,N_11172,N_10775);
nor U14324 (N_14324,N_10459,N_10541);
or U14325 (N_14325,N_11127,N_11041);
nand U14326 (N_14326,N_12145,N_12206);
or U14327 (N_14327,N_11543,N_11873);
nor U14328 (N_14328,N_12429,N_11027);
nand U14329 (N_14329,N_10583,N_11948);
nor U14330 (N_14330,N_11742,N_11264);
nor U14331 (N_14331,N_10927,N_12027);
nand U14332 (N_14332,N_10127,N_10141);
nor U14333 (N_14333,N_10703,N_11348);
nand U14334 (N_14334,N_11203,N_12211);
and U14335 (N_14335,N_10046,N_11524);
nand U14336 (N_14336,N_10012,N_11312);
or U14337 (N_14337,N_10663,N_11118);
nor U14338 (N_14338,N_11914,N_11587);
and U14339 (N_14339,N_12168,N_10914);
or U14340 (N_14340,N_10271,N_10940);
nor U14341 (N_14341,N_11110,N_10214);
nand U14342 (N_14342,N_11688,N_12065);
or U14343 (N_14343,N_11563,N_12192);
nor U14344 (N_14344,N_10781,N_11127);
xnor U14345 (N_14345,N_10466,N_10405);
nand U14346 (N_14346,N_11502,N_11300);
and U14347 (N_14347,N_11292,N_10719);
xnor U14348 (N_14348,N_12088,N_11590);
nor U14349 (N_14349,N_11760,N_11875);
xor U14350 (N_14350,N_11907,N_10639);
nand U14351 (N_14351,N_10552,N_11629);
and U14352 (N_14352,N_10718,N_11823);
and U14353 (N_14353,N_10568,N_10432);
and U14354 (N_14354,N_11321,N_12163);
or U14355 (N_14355,N_10809,N_12128);
nand U14356 (N_14356,N_10600,N_11098);
nand U14357 (N_14357,N_10098,N_12082);
and U14358 (N_14358,N_11665,N_12140);
nor U14359 (N_14359,N_10781,N_10332);
nor U14360 (N_14360,N_10281,N_12356);
and U14361 (N_14361,N_11885,N_10957);
nand U14362 (N_14362,N_12030,N_11539);
nand U14363 (N_14363,N_10469,N_11932);
or U14364 (N_14364,N_11018,N_12246);
nor U14365 (N_14365,N_12320,N_11575);
or U14366 (N_14366,N_11781,N_11058);
nand U14367 (N_14367,N_11210,N_12468);
and U14368 (N_14368,N_11836,N_11391);
nor U14369 (N_14369,N_10612,N_12205);
and U14370 (N_14370,N_11911,N_12424);
nand U14371 (N_14371,N_11464,N_10741);
or U14372 (N_14372,N_10947,N_10065);
or U14373 (N_14373,N_11083,N_10953);
nor U14374 (N_14374,N_10666,N_11204);
nand U14375 (N_14375,N_11380,N_11339);
and U14376 (N_14376,N_10380,N_10407);
nor U14377 (N_14377,N_10443,N_11214);
and U14378 (N_14378,N_10982,N_11350);
and U14379 (N_14379,N_11283,N_10937);
nand U14380 (N_14380,N_11344,N_12421);
and U14381 (N_14381,N_11101,N_11104);
nor U14382 (N_14382,N_10682,N_11109);
or U14383 (N_14383,N_10982,N_12194);
nor U14384 (N_14384,N_11448,N_11090);
and U14385 (N_14385,N_10676,N_11486);
and U14386 (N_14386,N_11093,N_12035);
nand U14387 (N_14387,N_11233,N_10514);
nor U14388 (N_14388,N_10422,N_10556);
and U14389 (N_14389,N_10069,N_11041);
nand U14390 (N_14390,N_11432,N_10058);
or U14391 (N_14391,N_10636,N_12365);
or U14392 (N_14392,N_10071,N_11136);
or U14393 (N_14393,N_12041,N_12208);
nand U14394 (N_14394,N_12035,N_11574);
nor U14395 (N_14395,N_11528,N_10910);
nor U14396 (N_14396,N_12452,N_12097);
nor U14397 (N_14397,N_11605,N_12266);
or U14398 (N_14398,N_12303,N_11438);
and U14399 (N_14399,N_12382,N_11090);
nand U14400 (N_14400,N_10344,N_11966);
or U14401 (N_14401,N_11437,N_10292);
and U14402 (N_14402,N_11441,N_11611);
nor U14403 (N_14403,N_11344,N_10850);
and U14404 (N_14404,N_11350,N_10046);
or U14405 (N_14405,N_10355,N_10344);
or U14406 (N_14406,N_11491,N_10387);
and U14407 (N_14407,N_10325,N_10195);
nand U14408 (N_14408,N_12416,N_11533);
nor U14409 (N_14409,N_11954,N_11174);
nand U14410 (N_14410,N_10646,N_10265);
and U14411 (N_14411,N_12428,N_10194);
nor U14412 (N_14412,N_11223,N_10108);
and U14413 (N_14413,N_10116,N_12223);
or U14414 (N_14414,N_10598,N_12140);
nand U14415 (N_14415,N_11896,N_10993);
or U14416 (N_14416,N_10570,N_11324);
nor U14417 (N_14417,N_10415,N_10442);
and U14418 (N_14418,N_10395,N_12263);
nor U14419 (N_14419,N_10406,N_10794);
and U14420 (N_14420,N_11787,N_11774);
or U14421 (N_14421,N_10307,N_10152);
or U14422 (N_14422,N_11465,N_11287);
nand U14423 (N_14423,N_11931,N_10397);
nor U14424 (N_14424,N_12302,N_11338);
and U14425 (N_14425,N_11699,N_10269);
and U14426 (N_14426,N_10796,N_10825);
xor U14427 (N_14427,N_10190,N_12125);
and U14428 (N_14428,N_10798,N_11872);
or U14429 (N_14429,N_12489,N_10371);
or U14430 (N_14430,N_10873,N_10614);
nand U14431 (N_14431,N_11132,N_11790);
nor U14432 (N_14432,N_10272,N_10470);
and U14433 (N_14433,N_11988,N_10099);
and U14434 (N_14434,N_11733,N_10610);
and U14435 (N_14435,N_11473,N_12024);
xnor U14436 (N_14436,N_10772,N_11940);
or U14437 (N_14437,N_11068,N_10724);
nor U14438 (N_14438,N_11976,N_10469);
and U14439 (N_14439,N_11273,N_11475);
nor U14440 (N_14440,N_12160,N_10808);
nand U14441 (N_14441,N_10980,N_11841);
nor U14442 (N_14442,N_10526,N_10482);
and U14443 (N_14443,N_11163,N_10076);
nand U14444 (N_14444,N_10847,N_11603);
nor U14445 (N_14445,N_12103,N_12202);
nand U14446 (N_14446,N_12025,N_12169);
and U14447 (N_14447,N_10705,N_10237);
or U14448 (N_14448,N_11169,N_11382);
and U14449 (N_14449,N_12404,N_12286);
or U14450 (N_14450,N_11089,N_10567);
nand U14451 (N_14451,N_10686,N_10774);
nand U14452 (N_14452,N_10655,N_11372);
or U14453 (N_14453,N_10055,N_11015);
nor U14454 (N_14454,N_10043,N_10592);
nor U14455 (N_14455,N_10890,N_12382);
nor U14456 (N_14456,N_10157,N_11045);
nand U14457 (N_14457,N_10130,N_11998);
nor U14458 (N_14458,N_11940,N_11321);
nor U14459 (N_14459,N_10480,N_10622);
and U14460 (N_14460,N_10546,N_10026);
or U14461 (N_14461,N_11570,N_11093);
nand U14462 (N_14462,N_12027,N_10787);
and U14463 (N_14463,N_11249,N_12375);
nand U14464 (N_14464,N_10177,N_12269);
nor U14465 (N_14465,N_10900,N_10578);
nand U14466 (N_14466,N_11603,N_11707);
and U14467 (N_14467,N_10655,N_12460);
nand U14468 (N_14468,N_10748,N_12079);
nand U14469 (N_14469,N_12237,N_10622);
or U14470 (N_14470,N_12197,N_11989);
xor U14471 (N_14471,N_10416,N_11569);
nand U14472 (N_14472,N_11900,N_10539);
nor U14473 (N_14473,N_11040,N_11476);
nand U14474 (N_14474,N_10787,N_12423);
and U14475 (N_14475,N_10571,N_10694);
and U14476 (N_14476,N_11231,N_10952);
and U14477 (N_14477,N_11693,N_10038);
nor U14478 (N_14478,N_11211,N_11849);
and U14479 (N_14479,N_11043,N_11810);
nor U14480 (N_14480,N_11336,N_11524);
and U14481 (N_14481,N_12039,N_12060);
nand U14482 (N_14482,N_10608,N_11521);
and U14483 (N_14483,N_11795,N_12256);
or U14484 (N_14484,N_10147,N_11692);
or U14485 (N_14485,N_10416,N_12045);
or U14486 (N_14486,N_11865,N_11577);
nor U14487 (N_14487,N_10314,N_10502);
and U14488 (N_14488,N_11077,N_10507);
nor U14489 (N_14489,N_11520,N_11291);
and U14490 (N_14490,N_10913,N_11451);
nor U14491 (N_14491,N_11942,N_10255);
nor U14492 (N_14492,N_10929,N_10697);
and U14493 (N_14493,N_11229,N_10945);
xor U14494 (N_14494,N_10736,N_10254);
or U14495 (N_14495,N_11297,N_11439);
and U14496 (N_14496,N_11886,N_10240);
nor U14497 (N_14497,N_10127,N_11607);
and U14498 (N_14498,N_11145,N_10814);
or U14499 (N_14499,N_11016,N_12042);
or U14500 (N_14500,N_12301,N_11706);
xor U14501 (N_14501,N_12434,N_10266);
or U14502 (N_14502,N_12345,N_10701);
or U14503 (N_14503,N_10709,N_12037);
xor U14504 (N_14504,N_11477,N_10892);
and U14505 (N_14505,N_10892,N_11674);
or U14506 (N_14506,N_12261,N_11782);
nor U14507 (N_14507,N_11202,N_11924);
nand U14508 (N_14508,N_12157,N_10951);
and U14509 (N_14509,N_10856,N_10195);
and U14510 (N_14510,N_11146,N_10364);
nand U14511 (N_14511,N_12072,N_11483);
nor U14512 (N_14512,N_10204,N_12102);
nor U14513 (N_14513,N_10075,N_12137);
and U14514 (N_14514,N_10869,N_10139);
nand U14515 (N_14515,N_11302,N_11726);
and U14516 (N_14516,N_11000,N_11201);
nor U14517 (N_14517,N_10759,N_10213);
or U14518 (N_14518,N_12097,N_10338);
and U14519 (N_14519,N_12281,N_11906);
nand U14520 (N_14520,N_12177,N_12156);
and U14521 (N_14521,N_11557,N_11073);
or U14522 (N_14522,N_12460,N_10954);
and U14523 (N_14523,N_10711,N_10714);
nor U14524 (N_14524,N_11201,N_11422);
nand U14525 (N_14525,N_10470,N_11360);
or U14526 (N_14526,N_11560,N_12479);
nand U14527 (N_14527,N_11627,N_11585);
or U14528 (N_14528,N_10107,N_10596);
nor U14529 (N_14529,N_11172,N_10261);
and U14530 (N_14530,N_11014,N_11768);
nand U14531 (N_14531,N_10715,N_11400);
xnor U14532 (N_14532,N_11880,N_10125);
nand U14533 (N_14533,N_11789,N_10798);
and U14534 (N_14534,N_11281,N_10238);
and U14535 (N_14535,N_11005,N_10278);
nand U14536 (N_14536,N_12106,N_12034);
nor U14537 (N_14537,N_11295,N_12481);
nand U14538 (N_14538,N_11620,N_10254);
or U14539 (N_14539,N_12094,N_11143);
nor U14540 (N_14540,N_10085,N_12212);
and U14541 (N_14541,N_11182,N_10604);
nand U14542 (N_14542,N_10605,N_12335);
nor U14543 (N_14543,N_11099,N_10451);
or U14544 (N_14544,N_11628,N_12232);
or U14545 (N_14545,N_10762,N_12374);
or U14546 (N_14546,N_11401,N_10754);
or U14547 (N_14547,N_11383,N_10468);
nor U14548 (N_14548,N_11843,N_10668);
nor U14549 (N_14549,N_11866,N_11512);
nand U14550 (N_14550,N_11095,N_10541);
and U14551 (N_14551,N_11602,N_10755);
or U14552 (N_14552,N_11826,N_10287);
nand U14553 (N_14553,N_10555,N_10418);
and U14554 (N_14554,N_11211,N_11944);
and U14555 (N_14555,N_11532,N_10530);
xor U14556 (N_14556,N_11027,N_11387);
and U14557 (N_14557,N_10687,N_11529);
and U14558 (N_14558,N_11726,N_11511);
nor U14559 (N_14559,N_10933,N_10934);
and U14560 (N_14560,N_11073,N_12102);
nand U14561 (N_14561,N_10935,N_11478);
nor U14562 (N_14562,N_11007,N_12252);
nor U14563 (N_14563,N_10554,N_10973);
nand U14564 (N_14564,N_12237,N_12381);
nand U14565 (N_14565,N_10014,N_12286);
and U14566 (N_14566,N_11427,N_10252);
nor U14567 (N_14567,N_11107,N_10116);
or U14568 (N_14568,N_11482,N_10020);
or U14569 (N_14569,N_11880,N_10282);
and U14570 (N_14570,N_10813,N_11784);
nand U14571 (N_14571,N_10814,N_11383);
nand U14572 (N_14572,N_11034,N_11819);
or U14573 (N_14573,N_10803,N_11196);
nor U14574 (N_14574,N_10010,N_10983);
nor U14575 (N_14575,N_11340,N_10711);
and U14576 (N_14576,N_11555,N_10541);
xnor U14577 (N_14577,N_11762,N_10867);
nor U14578 (N_14578,N_12224,N_12034);
and U14579 (N_14579,N_10071,N_10190);
nor U14580 (N_14580,N_10213,N_11039);
nor U14581 (N_14581,N_10311,N_11126);
or U14582 (N_14582,N_12077,N_10027);
nand U14583 (N_14583,N_12460,N_11394);
nor U14584 (N_14584,N_11533,N_10156);
or U14585 (N_14585,N_10149,N_11734);
or U14586 (N_14586,N_11284,N_10264);
nand U14587 (N_14587,N_10459,N_10500);
and U14588 (N_14588,N_10482,N_10488);
or U14589 (N_14589,N_12294,N_11744);
nand U14590 (N_14590,N_12394,N_11257);
or U14591 (N_14591,N_12424,N_11010);
or U14592 (N_14592,N_10425,N_11463);
or U14593 (N_14593,N_11976,N_11874);
nor U14594 (N_14594,N_12105,N_10629);
nand U14595 (N_14595,N_10471,N_11022);
and U14596 (N_14596,N_10696,N_10903);
nand U14597 (N_14597,N_12303,N_10026);
nand U14598 (N_14598,N_11614,N_10566);
or U14599 (N_14599,N_10559,N_10751);
nand U14600 (N_14600,N_10735,N_11771);
and U14601 (N_14601,N_10326,N_11784);
nor U14602 (N_14602,N_10790,N_10859);
nand U14603 (N_14603,N_11855,N_10643);
nor U14604 (N_14604,N_11630,N_10964);
nand U14605 (N_14605,N_12001,N_11803);
xor U14606 (N_14606,N_11804,N_10910);
or U14607 (N_14607,N_11585,N_12077);
and U14608 (N_14608,N_12286,N_11759);
or U14609 (N_14609,N_10851,N_11965);
and U14610 (N_14610,N_11282,N_11711);
nor U14611 (N_14611,N_11360,N_10365);
nor U14612 (N_14612,N_11225,N_10545);
or U14613 (N_14613,N_12212,N_10300);
nor U14614 (N_14614,N_11938,N_10545);
nand U14615 (N_14615,N_11563,N_12119);
and U14616 (N_14616,N_10104,N_11382);
nand U14617 (N_14617,N_12256,N_11633);
or U14618 (N_14618,N_11933,N_12482);
or U14619 (N_14619,N_10231,N_11449);
nand U14620 (N_14620,N_11883,N_10099);
or U14621 (N_14621,N_11409,N_11515);
and U14622 (N_14622,N_10198,N_10191);
nor U14623 (N_14623,N_10293,N_12081);
and U14624 (N_14624,N_10644,N_10836);
and U14625 (N_14625,N_12185,N_11742);
or U14626 (N_14626,N_11237,N_10758);
nor U14627 (N_14627,N_11698,N_11304);
and U14628 (N_14628,N_10914,N_10052);
nand U14629 (N_14629,N_11118,N_12314);
nor U14630 (N_14630,N_10232,N_12060);
and U14631 (N_14631,N_10635,N_10446);
nand U14632 (N_14632,N_10232,N_10092);
nand U14633 (N_14633,N_10883,N_11535);
and U14634 (N_14634,N_12054,N_10843);
nand U14635 (N_14635,N_10641,N_10504);
or U14636 (N_14636,N_11826,N_11831);
or U14637 (N_14637,N_11768,N_10364);
nand U14638 (N_14638,N_10286,N_11116);
nand U14639 (N_14639,N_12089,N_11202);
nand U14640 (N_14640,N_11697,N_10212);
nor U14641 (N_14641,N_12210,N_10279);
nor U14642 (N_14642,N_10880,N_11231);
or U14643 (N_14643,N_11860,N_10645);
or U14644 (N_14644,N_12323,N_11099);
and U14645 (N_14645,N_12030,N_10058);
nor U14646 (N_14646,N_10114,N_12023);
nand U14647 (N_14647,N_11708,N_10299);
and U14648 (N_14648,N_10389,N_10437);
or U14649 (N_14649,N_11478,N_12314);
and U14650 (N_14650,N_12007,N_11160);
or U14651 (N_14651,N_10303,N_12215);
nand U14652 (N_14652,N_10777,N_10985);
or U14653 (N_14653,N_11247,N_11601);
nor U14654 (N_14654,N_11499,N_10563);
nand U14655 (N_14655,N_11306,N_12081);
or U14656 (N_14656,N_10248,N_10561);
and U14657 (N_14657,N_11930,N_10588);
nor U14658 (N_14658,N_11057,N_12169);
or U14659 (N_14659,N_12276,N_11931);
or U14660 (N_14660,N_12474,N_10019);
and U14661 (N_14661,N_10750,N_11707);
nor U14662 (N_14662,N_11718,N_10467);
nor U14663 (N_14663,N_11313,N_11221);
nor U14664 (N_14664,N_11196,N_12171);
nor U14665 (N_14665,N_10210,N_10790);
nor U14666 (N_14666,N_11171,N_12002);
nor U14667 (N_14667,N_11863,N_11255);
nand U14668 (N_14668,N_10300,N_12117);
nor U14669 (N_14669,N_12441,N_12134);
or U14670 (N_14670,N_11732,N_12381);
nor U14671 (N_14671,N_12036,N_11434);
nor U14672 (N_14672,N_12230,N_11684);
and U14673 (N_14673,N_10340,N_10712);
nor U14674 (N_14674,N_10973,N_10596);
and U14675 (N_14675,N_12064,N_11819);
and U14676 (N_14676,N_12091,N_10219);
or U14677 (N_14677,N_11616,N_12074);
or U14678 (N_14678,N_10515,N_12154);
and U14679 (N_14679,N_10272,N_11986);
and U14680 (N_14680,N_10969,N_12078);
or U14681 (N_14681,N_10024,N_10281);
nor U14682 (N_14682,N_12090,N_10041);
nand U14683 (N_14683,N_11960,N_10177);
or U14684 (N_14684,N_11467,N_11386);
and U14685 (N_14685,N_12294,N_12406);
nand U14686 (N_14686,N_10123,N_11886);
or U14687 (N_14687,N_11958,N_10148);
or U14688 (N_14688,N_10672,N_10546);
nand U14689 (N_14689,N_11432,N_11213);
nand U14690 (N_14690,N_10049,N_11767);
or U14691 (N_14691,N_10934,N_11105);
or U14692 (N_14692,N_10444,N_11547);
nor U14693 (N_14693,N_10409,N_12280);
or U14694 (N_14694,N_12395,N_12030);
nor U14695 (N_14695,N_10476,N_12195);
nand U14696 (N_14696,N_10456,N_10343);
nand U14697 (N_14697,N_12143,N_11393);
or U14698 (N_14698,N_10933,N_11518);
nor U14699 (N_14699,N_11983,N_11390);
nand U14700 (N_14700,N_10897,N_11290);
nand U14701 (N_14701,N_11718,N_12301);
xor U14702 (N_14702,N_11182,N_11560);
nor U14703 (N_14703,N_11554,N_12320);
or U14704 (N_14704,N_12284,N_11740);
and U14705 (N_14705,N_10466,N_11204);
xor U14706 (N_14706,N_11262,N_11559);
nand U14707 (N_14707,N_11632,N_10866);
nor U14708 (N_14708,N_11573,N_11060);
or U14709 (N_14709,N_11746,N_12425);
and U14710 (N_14710,N_11993,N_11742);
and U14711 (N_14711,N_11718,N_11980);
nand U14712 (N_14712,N_12380,N_12256);
or U14713 (N_14713,N_10101,N_11767);
and U14714 (N_14714,N_10754,N_11217);
nor U14715 (N_14715,N_11214,N_11036);
nand U14716 (N_14716,N_12137,N_12288);
and U14717 (N_14717,N_10464,N_12018);
nand U14718 (N_14718,N_11361,N_12296);
and U14719 (N_14719,N_12348,N_10084);
and U14720 (N_14720,N_11384,N_10538);
nor U14721 (N_14721,N_10864,N_11265);
or U14722 (N_14722,N_10614,N_11526);
or U14723 (N_14723,N_12303,N_11156);
xnor U14724 (N_14724,N_10554,N_11406);
nand U14725 (N_14725,N_12415,N_12480);
and U14726 (N_14726,N_10397,N_10401);
nand U14727 (N_14727,N_10144,N_10383);
nand U14728 (N_14728,N_10120,N_10108);
or U14729 (N_14729,N_10006,N_11325);
or U14730 (N_14730,N_12472,N_12347);
nand U14731 (N_14731,N_10341,N_11864);
nand U14732 (N_14732,N_12446,N_10782);
nand U14733 (N_14733,N_10718,N_11461);
or U14734 (N_14734,N_12197,N_10576);
and U14735 (N_14735,N_12467,N_10649);
nand U14736 (N_14736,N_10937,N_11828);
and U14737 (N_14737,N_12299,N_10668);
nand U14738 (N_14738,N_10614,N_11522);
nor U14739 (N_14739,N_10553,N_11521);
and U14740 (N_14740,N_10362,N_11873);
xnor U14741 (N_14741,N_11391,N_11555);
nor U14742 (N_14742,N_11015,N_10758);
nand U14743 (N_14743,N_10037,N_10507);
nor U14744 (N_14744,N_10926,N_10074);
or U14745 (N_14745,N_10633,N_10987);
xor U14746 (N_14746,N_11628,N_11625);
nor U14747 (N_14747,N_12457,N_12113);
and U14748 (N_14748,N_11450,N_12282);
and U14749 (N_14749,N_10481,N_11791);
nor U14750 (N_14750,N_10425,N_12079);
nor U14751 (N_14751,N_11340,N_10302);
nand U14752 (N_14752,N_12417,N_10006);
nand U14753 (N_14753,N_12150,N_12051);
or U14754 (N_14754,N_11304,N_12414);
nor U14755 (N_14755,N_10204,N_11391);
nand U14756 (N_14756,N_11329,N_11717);
and U14757 (N_14757,N_10218,N_11153);
or U14758 (N_14758,N_11211,N_11369);
nor U14759 (N_14759,N_11335,N_12194);
nor U14760 (N_14760,N_12422,N_10346);
and U14761 (N_14761,N_10111,N_10014);
and U14762 (N_14762,N_11232,N_10244);
or U14763 (N_14763,N_11104,N_12295);
nor U14764 (N_14764,N_11099,N_11262);
nand U14765 (N_14765,N_10688,N_12368);
or U14766 (N_14766,N_12428,N_11159);
nand U14767 (N_14767,N_11902,N_10169);
and U14768 (N_14768,N_11078,N_10313);
xor U14769 (N_14769,N_12351,N_12078);
nor U14770 (N_14770,N_10106,N_10982);
xnor U14771 (N_14771,N_12124,N_11707);
and U14772 (N_14772,N_10666,N_12459);
nor U14773 (N_14773,N_10527,N_11614);
and U14774 (N_14774,N_12356,N_12257);
or U14775 (N_14775,N_10208,N_12457);
nand U14776 (N_14776,N_10678,N_11065);
nor U14777 (N_14777,N_11850,N_10575);
nor U14778 (N_14778,N_12007,N_11001);
xor U14779 (N_14779,N_10477,N_11259);
and U14780 (N_14780,N_11190,N_11193);
and U14781 (N_14781,N_11403,N_10163);
nor U14782 (N_14782,N_10132,N_11146);
and U14783 (N_14783,N_11177,N_11527);
or U14784 (N_14784,N_11431,N_12109);
nor U14785 (N_14785,N_11393,N_10126);
nor U14786 (N_14786,N_10748,N_10022);
nand U14787 (N_14787,N_10034,N_12304);
and U14788 (N_14788,N_10210,N_12256);
and U14789 (N_14789,N_12009,N_11488);
or U14790 (N_14790,N_11783,N_11174);
nor U14791 (N_14791,N_10513,N_11711);
nand U14792 (N_14792,N_11252,N_10474);
or U14793 (N_14793,N_10142,N_10010);
nor U14794 (N_14794,N_11996,N_11026);
nand U14795 (N_14795,N_10654,N_12326);
nor U14796 (N_14796,N_10930,N_11446);
and U14797 (N_14797,N_10760,N_12346);
nand U14798 (N_14798,N_10966,N_11395);
nand U14799 (N_14799,N_10324,N_10915);
or U14800 (N_14800,N_10760,N_10195);
nand U14801 (N_14801,N_10437,N_11642);
nand U14802 (N_14802,N_12338,N_12227);
and U14803 (N_14803,N_11358,N_11202);
nor U14804 (N_14804,N_10028,N_11315);
nand U14805 (N_14805,N_11343,N_10081);
nor U14806 (N_14806,N_10251,N_12026);
nor U14807 (N_14807,N_10978,N_11520);
nand U14808 (N_14808,N_10661,N_11125);
and U14809 (N_14809,N_11038,N_10474);
or U14810 (N_14810,N_11600,N_11319);
and U14811 (N_14811,N_10106,N_12268);
nand U14812 (N_14812,N_11634,N_10855);
or U14813 (N_14813,N_11584,N_10567);
and U14814 (N_14814,N_11473,N_12390);
or U14815 (N_14815,N_12436,N_11533);
nor U14816 (N_14816,N_12024,N_10734);
or U14817 (N_14817,N_10254,N_11556);
or U14818 (N_14818,N_11253,N_10973);
nand U14819 (N_14819,N_11995,N_10039);
or U14820 (N_14820,N_10343,N_11666);
or U14821 (N_14821,N_11663,N_12031);
nand U14822 (N_14822,N_11965,N_11159);
and U14823 (N_14823,N_11154,N_10573);
or U14824 (N_14824,N_12131,N_11556);
or U14825 (N_14825,N_10939,N_12036);
or U14826 (N_14826,N_10417,N_12430);
nor U14827 (N_14827,N_11455,N_10820);
nand U14828 (N_14828,N_10750,N_12215);
and U14829 (N_14829,N_12450,N_11917);
or U14830 (N_14830,N_11380,N_11559);
xor U14831 (N_14831,N_12286,N_11821);
nor U14832 (N_14832,N_10581,N_10804);
nand U14833 (N_14833,N_10926,N_11796);
or U14834 (N_14834,N_10314,N_12153);
and U14835 (N_14835,N_10495,N_12417);
or U14836 (N_14836,N_10580,N_11631);
nor U14837 (N_14837,N_11137,N_11710);
and U14838 (N_14838,N_10033,N_12345);
and U14839 (N_14839,N_12377,N_12267);
nor U14840 (N_14840,N_10661,N_10240);
and U14841 (N_14841,N_10483,N_11037);
nor U14842 (N_14842,N_12395,N_10975);
or U14843 (N_14843,N_10624,N_12180);
and U14844 (N_14844,N_11744,N_10198);
nand U14845 (N_14845,N_12062,N_11352);
nor U14846 (N_14846,N_12337,N_10731);
nand U14847 (N_14847,N_11194,N_12447);
nor U14848 (N_14848,N_11772,N_10692);
or U14849 (N_14849,N_10234,N_10695);
or U14850 (N_14850,N_11248,N_11644);
or U14851 (N_14851,N_12396,N_10700);
or U14852 (N_14852,N_11873,N_10620);
nor U14853 (N_14853,N_11669,N_11707);
and U14854 (N_14854,N_11594,N_11661);
or U14855 (N_14855,N_10832,N_10531);
and U14856 (N_14856,N_10149,N_12189);
and U14857 (N_14857,N_11758,N_10222);
and U14858 (N_14858,N_12146,N_10971);
and U14859 (N_14859,N_11481,N_10371);
nor U14860 (N_14860,N_12239,N_11183);
nor U14861 (N_14861,N_10787,N_11865);
nor U14862 (N_14862,N_11216,N_10780);
nor U14863 (N_14863,N_10514,N_11224);
and U14864 (N_14864,N_12323,N_12215);
nand U14865 (N_14865,N_12402,N_10733);
nand U14866 (N_14866,N_11049,N_12168);
xnor U14867 (N_14867,N_11700,N_11061);
or U14868 (N_14868,N_12366,N_10479);
and U14869 (N_14869,N_12224,N_10610);
and U14870 (N_14870,N_12123,N_11594);
and U14871 (N_14871,N_11191,N_11181);
nand U14872 (N_14872,N_11491,N_10162);
nor U14873 (N_14873,N_12133,N_10642);
xnor U14874 (N_14874,N_12064,N_11384);
and U14875 (N_14875,N_12375,N_10197);
xor U14876 (N_14876,N_11057,N_12016);
or U14877 (N_14877,N_11613,N_10196);
and U14878 (N_14878,N_12018,N_10652);
xor U14879 (N_14879,N_10940,N_11305);
nand U14880 (N_14880,N_12190,N_12331);
nand U14881 (N_14881,N_11362,N_10701);
and U14882 (N_14882,N_11810,N_11879);
nand U14883 (N_14883,N_11086,N_11681);
nor U14884 (N_14884,N_11432,N_12373);
and U14885 (N_14885,N_10507,N_12008);
nand U14886 (N_14886,N_10011,N_11273);
or U14887 (N_14887,N_12250,N_10055);
and U14888 (N_14888,N_10117,N_10132);
nand U14889 (N_14889,N_11980,N_11567);
nand U14890 (N_14890,N_10922,N_11871);
and U14891 (N_14891,N_12304,N_10231);
xor U14892 (N_14892,N_10713,N_11974);
and U14893 (N_14893,N_10331,N_11734);
or U14894 (N_14894,N_10243,N_12460);
nand U14895 (N_14895,N_11910,N_10011);
and U14896 (N_14896,N_10013,N_11727);
nor U14897 (N_14897,N_11632,N_11166);
or U14898 (N_14898,N_10431,N_11524);
or U14899 (N_14899,N_12099,N_12464);
nand U14900 (N_14900,N_10786,N_12351);
or U14901 (N_14901,N_10521,N_12460);
or U14902 (N_14902,N_11482,N_11366);
nor U14903 (N_14903,N_10368,N_11450);
and U14904 (N_14904,N_12071,N_12007);
and U14905 (N_14905,N_12309,N_10650);
nand U14906 (N_14906,N_10599,N_10894);
nand U14907 (N_14907,N_11054,N_11618);
and U14908 (N_14908,N_10673,N_12299);
nor U14909 (N_14909,N_12240,N_10486);
nand U14910 (N_14910,N_11364,N_10833);
nand U14911 (N_14911,N_11693,N_12014);
nand U14912 (N_14912,N_10288,N_12051);
and U14913 (N_14913,N_10354,N_10769);
or U14914 (N_14914,N_11001,N_11670);
nand U14915 (N_14915,N_10579,N_11382);
and U14916 (N_14916,N_10306,N_11162);
nand U14917 (N_14917,N_11528,N_12154);
and U14918 (N_14918,N_10770,N_10978);
nand U14919 (N_14919,N_10759,N_11133);
or U14920 (N_14920,N_10837,N_10212);
or U14921 (N_14921,N_10622,N_11281);
nand U14922 (N_14922,N_11303,N_10803);
nor U14923 (N_14923,N_10717,N_10950);
xor U14924 (N_14924,N_10363,N_10518);
and U14925 (N_14925,N_11373,N_11633);
nor U14926 (N_14926,N_11266,N_10397);
or U14927 (N_14927,N_12452,N_12417);
or U14928 (N_14928,N_11059,N_12222);
and U14929 (N_14929,N_10753,N_10865);
and U14930 (N_14930,N_11657,N_11994);
nand U14931 (N_14931,N_10221,N_11901);
nand U14932 (N_14932,N_11816,N_10206);
nand U14933 (N_14933,N_12367,N_12144);
or U14934 (N_14934,N_11593,N_11662);
nand U14935 (N_14935,N_12201,N_11021);
and U14936 (N_14936,N_10466,N_11652);
and U14937 (N_14937,N_10959,N_10999);
nor U14938 (N_14938,N_10456,N_10065);
or U14939 (N_14939,N_11182,N_12451);
or U14940 (N_14940,N_10661,N_11375);
or U14941 (N_14941,N_11426,N_10182);
nor U14942 (N_14942,N_10286,N_11121);
nor U14943 (N_14943,N_12343,N_12108);
or U14944 (N_14944,N_11823,N_11310);
nand U14945 (N_14945,N_10065,N_10675);
nor U14946 (N_14946,N_10199,N_12187);
and U14947 (N_14947,N_11927,N_11293);
nor U14948 (N_14948,N_11605,N_11378);
and U14949 (N_14949,N_12363,N_12114);
and U14950 (N_14950,N_10559,N_10446);
nand U14951 (N_14951,N_10377,N_11919);
or U14952 (N_14952,N_11208,N_11052);
or U14953 (N_14953,N_11793,N_10792);
or U14954 (N_14954,N_10623,N_11271);
nand U14955 (N_14955,N_12025,N_11329);
or U14956 (N_14956,N_10482,N_10713);
nand U14957 (N_14957,N_12292,N_11767);
and U14958 (N_14958,N_10429,N_11066);
or U14959 (N_14959,N_11367,N_10126);
or U14960 (N_14960,N_10153,N_11846);
nand U14961 (N_14961,N_11064,N_11787);
nor U14962 (N_14962,N_12228,N_10674);
nor U14963 (N_14963,N_12468,N_12149);
or U14964 (N_14964,N_10901,N_10691);
nor U14965 (N_14965,N_11855,N_12241);
nor U14966 (N_14966,N_10439,N_11447);
and U14967 (N_14967,N_11305,N_12140);
and U14968 (N_14968,N_11840,N_10770);
or U14969 (N_14969,N_10958,N_10989);
and U14970 (N_14970,N_12482,N_10459);
or U14971 (N_14971,N_12375,N_10136);
and U14972 (N_14972,N_11851,N_10486);
nand U14973 (N_14973,N_11147,N_11945);
nor U14974 (N_14974,N_10229,N_10165);
nor U14975 (N_14975,N_11849,N_10711);
or U14976 (N_14976,N_10477,N_10060);
nand U14977 (N_14977,N_10507,N_10581);
nand U14978 (N_14978,N_11402,N_10495);
nor U14979 (N_14979,N_10900,N_10824);
or U14980 (N_14980,N_11700,N_11533);
nand U14981 (N_14981,N_10250,N_10427);
nand U14982 (N_14982,N_10763,N_12248);
nand U14983 (N_14983,N_10666,N_11597);
nand U14984 (N_14984,N_12079,N_12145);
and U14985 (N_14985,N_10021,N_11988);
nand U14986 (N_14986,N_10392,N_11698);
nor U14987 (N_14987,N_10639,N_12383);
or U14988 (N_14988,N_11741,N_11665);
and U14989 (N_14989,N_10264,N_11685);
nand U14990 (N_14990,N_11972,N_11344);
or U14991 (N_14991,N_10872,N_12065);
and U14992 (N_14992,N_10031,N_10246);
or U14993 (N_14993,N_12329,N_12177);
nor U14994 (N_14994,N_10500,N_10767);
and U14995 (N_14995,N_12433,N_11019);
nand U14996 (N_14996,N_10782,N_10691);
and U14997 (N_14997,N_11405,N_10402);
or U14998 (N_14998,N_11427,N_10927);
nor U14999 (N_14999,N_10849,N_11761);
nor U15000 (N_15000,N_14257,N_13065);
nand U15001 (N_15001,N_13059,N_14329);
or U15002 (N_15002,N_13528,N_14200);
xor U15003 (N_15003,N_13660,N_14083);
nor U15004 (N_15004,N_12732,N_12531);
nor U15005 (N_15005,N_12717,N_14190);
nor U15006 (N_15006,N_14781,N_14786);
and U15007 (N_15007,N_12904,N_12609);
or U15008 (N_15008,N_13147,N_12615);
xnor U15009 (N_15009,N_13689,N_13726);
nor U15010 (N_15010,N_12941,N_13252);
xor U15011 (N_15011,N_13184,N_14077);
and U15012 (N_15012,N_14220,N_14831);
and U15013 (N_15013,N_13724,N_14145);
nand U15014 (N_15014,N_14794,N_13008);
or U15015 (N_15015,N_13730,N_13535);
nor U15016 (N_15016,N_13221,N_14708);
and U15017 (N_15017,N_14446,N_12545);
and U15018 (N_15018,N_14139,N_14470);
and U15019 (N_15019,N_13069,N_13277);
or U15020 (N_15020,N_13132,N_12683);
nand U15021 (N_15021,N_14934,N_13722);
and U15022 (N_15022,N_13863,N_12963);
or U15023 (N_15023,N_14028,N_13579);
nor U15024 (N_15024,N_13245,N_14669);
nor U15025 (N_15025,N_14372,N_14944);
and U15026 (N_15026,N_13520,N_14108);
nand U15027 (N_15027,N_14624,N_14466);
and U15028 (N_15028,N_13011,N_14652);
or U15029 (N_15029,N_12928,N_13250);
nand U15030 (N_15030,N_13304,N_13156);
nand U15031 (N_15031,N_14534,N_12999);
nand U15032 (N_15032,N_13983,N_13920);
nor U15033 (N_15033,N_13495,N_13613);
xnor U15034 (N_15034,N_14898,N_12642);
and U15035 (N_15035,N_13403,N_13844);
and U15036 (N_15036,N_13461,N_14594);
and U15037 (N_15037,N_13067,N_14116);
or U15038 (N_15038,N_13977,N_14971);
or U15039 (N_15039,N_12739,N_14839);
and U15040 (N_15040,N_13299,N_14789);
nand U15041 (N_15041,N_14735,N_14032);
nor U15042 (N_15042,N_13849,N_12750);
nor U15043 (N_15043,N_14694,N_14851);
nor U15044 (N_15044,N_13661,N_12991);
nand U15045 (N_15045,N_14609,N_14818);
or U15046 (N_15046,N_14722,N_13697);
nor U15047 (N_15047,N_13950,N_12891);
and U15048 (N_15048,N_14821,N_13337);
nand U15049 (N_15049,N_13625,N_13100);
xor U15050 (N_15050,N_12653,N_14802);
and U15051 (N_15051,N_13344,N_13019);
and U15052 (N_15052,N_14129,N_14834);
nor U15053 (N_15053,N_13421,N_13936);
or U15054 (N_15054,N_13235,N_14113);
or U15055 (N_15055,N_13744,N_14175);
or U15056 (N_15056,N_13004,N_13387);
nand U15057 (N_15057,N_14399,N_14584);
nor U15058 (N_15058,N_13634,N_12586);
nor U15059 (N_15059,N_13257,N_14533);
nor U15060 (N_15060,N_13032,N_14138);
nor U15061 (N_15061,N_14302,N_13248);
and U15062 (N_15062,N_13971,N_13927);
or U15063 (N_15063,N_12743,N_14910);
and U15064 (N_15064,N_14580,N_14243);
nand U15065 (N_15065,N_13441,N_12795);
nand U15066 (N_15066,N_13511,N_12833);
or U15067 (N_15067,N_12767,N_14830);
nand U15068 (N_15068,N_13992,N_14305);
nor U15069 (N_15069,N_12898,N_13163);
nand U15070 (N_15070,N_13232,N_13972);
or U15071 (N_15071,N_14866,N_13050);
and U15072 (N_15072,N_13220,N_14073);
nor U15073 (N_15073,N_12501,N_13665);
nand U15074 (N_15074,N_13429,N_14563);
nand U15075 (N_15075,N_14306,N_14882);
nor U15076 (N_15076,N_12773,N_14878);
nand U15077 (N_15077,N_14948,N_12636);
nand U15078 (N_15078,N_14796,N_13669);
or U15079 (N_15079,N_13532,N_14330);
nor U15080 (N_15080,N_13126,N_14015);
nand U15081 (N_15081,N_14339,N_13400);
nor U15082 (N_15082,N_13855,N_13750);
and U15083 (N_15083,N_13305,N_12584);
or U15084 (N_15084,N_14435,N_13993);
and U15085 (N_15085,N_13349,N_13376);
nand U15086 (N_15086,N_14901,N_14541);
nand U15087 (N_15087,N_14750,N_13646);
or U15088 (N_15088,N_13153,N_14171);
and U15089 (N_15089,N_14319,N_14956);
and U15090 (N_15090,N_14179,N_12789);
or U15091 (N_15091,N_13213,N_14568);
and U15092 (N_15092,N_13228,N_13484);
or U15093 (N_15093,N_13773,N_14420);
and U15094 (N_15094,N_12864,N_14080);
or U15095 (N_15095,N_14498,N_13640);
nand U15096 (N_15096,N_14256,N_14785);
nand U15097 (N_15097,N_14599,N_14740);
and U15098 (N_15098,N_14096,N_14185);
nand U15099 (N_15099,N_14726,N_13631);
nor U15100 (N_15100,N_13289,N_13326);
nand U15101 (N_15101,N_14743,N_14749);
or U15102 (N_15102,N_13767,N_13058);
nor U15103 (N_15103,N_13015,N_14981);
nor U15104 (N_15104,N_12747,N_13831);
nor U15105 (N_15105,N_13771,N_14021);
and U15106 (N_15106,N_13715,N_13035);
nor U15107 (N_15107,N_14495,N_14439);
nor U15108 (N_15108,N_13406,N_12948);
or U15109 (N_15109,N_12654,N_12556);
and U15110 (N_15110,N_14227,N_14614);
and U15111 (N_15111,N_13399,N_12716);
or U15112 (N_15112,N_12665,N_12844);
and U15113 (N_15113,N_13224,N_14642);
and U15114 (N_15114,N_13414,N_14018);
and U15115 (N_15115,N_14904,N_13330);
or U15116 (N_15116,N_14564,N_13572);
nor U15117 (N_15117,N_14586,N_13791);
or U15118 (N_15118,N_13654,N_13493);
or U15119 (N_15119,N_13926,N_14776);
or U15120 (N_15120,N_14408,N_13494);
and U15121 (N_15121,N_14770,N_13786);
nor U15122 (N_15122,N_14198,N_13448);
and U15123 (N_15123,N_14641,N_14141);
nor U15124 (N_15124,N_14380,N_14999);
and U15125 (N_15125,N_12633,N_14062);
nand U15126 (N_15126,N_13449,N_12876);
nand U15127 (N_15127,N_12583,N_13693);
and U15128 (N_15128,N_13042,N_14538);
and U15129 (N_15129,N_13986,N_14556);
nor U15130 (N_15130,N_12511,N_13393);
nor U15131 (N_15131,N_14079,N_12679);
nor U15132 (N_15132,N_12765,N_14637);
and U15133 (N_15133,N_13763,N_14053);
nor U15134 (N_15134,N_14909,N_13995);
and U15135 (N_15135,N_13149,N_14350);
and U15136 (N_15136,N_13133,N_14665);
and U15137 (N_15137,N_14484,N_12605);
nand U15138 (N_15138,N_13630,N_13817);
xor U15139 (N_15139,N_13793,N_12618);
or U15140 (N_15140,N_14033,N_13548);
or U15141 (N_15141,N_14627,N_12906);
or U15142 (N_15142,N_13881,N_14687);
or U15143 (N_15143,N_14993,N_13322);
xnor U15144 (N_15144,N_13368,N_14915);
and U15145 (N_15145,N_13641,N_13988);
or U15146 (N_15146,N_14300,N_12643);
and U15147 (N_15147,N_13291,N_12672);
nor U15148 (N_15148,N_14346,N_14730);
nor U15149 (N_15149,N_13009,N_14165);
and U15150 (N_15150,N_14320,N_14589);
nor U15151 (N_15151,N_14112,N_13800);
and U15152 (N_15152,N_13128,N_14762);
nor U15153 (N_15153,N_13216,N_12984);
and U15154 (N_15154,N_12567,N_14157);
xnor U15155 (N_15155,N_14006,N_14701);
nor U15156 (N_15156,N_12554,N_12604);
nor U15157 (N_15157,N_13889,N_13488);
and U15158 (N_15158,N_14647,N_14772);
and U15159 (N_15159,N_14825,N_13016);
or U15160 (N_15160,N_13901,N_14558);
nor U15161 (N_15161,N_13138,N_14648);
nand U15162 (N_15162,N_14264,N_13599);
nand U15163 (N_15163,N_13981,N_14529);
and U15164 (N_15164,N_13570,N_14936);
or U15165 (N_15165,N_14155,N_12862);
nor U15166 (N_15166,N_13618,N_14613);
or U15167 (N_15167,N_14115,N_14386);
and U15168 (N_15168,N_13051,N_13336);
nand U15169 (N_15169,N_14656,N_14164);
nor U15170 (N_15170,N_13595,N_12582);
or U15171 (N_15171,N_12832,N_14737);
nand U15172 (N_15172,N_13876,N_14055);
or U15173 (N_15173,N_13062,N_13148);
nor U15174 (N_15174,N_13472,N_14700);
nand U15175 (N_15175,N_14448,N_14751);
or U15176 (N_15176,N_14536,N_14712);
nand U15177 (N_15177,N_14047,N_14102);
nor U15178 (N_15178,N_13467,N_13928);
xor U15179 (N_15179,N_14219,N_12623);
nand U15180 (N_15180,N_14421,N_13524);
nand U15181 (N_15181,N_14244,N_13783);
nand U15182 (N_15182,N_14392,N_14622);
nor U15183 (N_15183,N_13366,N_13859);
nor U15184 (N_15184,N_13940,N_13604);
and U15185 (N_15185,N_12825,N_14638);
nand U15186 (N_15186,N_13764,N_13556);
nor U15187 (N_15187,N_12896,N_14496);
or U15188 (N_15188,N_13670,N_12733);
nand U15189 (N_15189,N_12974,N_12921);
nand U15190 (N_15190,N_14389,N_12845);
nor U15191 (N_15191,N_14605,N_12805);
nand U15192 (N_15192,N_13395,N_14943);
or U15193 (N_15193,N_14537,N_12889);
nand U15194 (N_15194,N_13010,N_13696);
or U15195 (N_15195,N_14527,N_14229);
nor U15196 (N_15196,N_14042,N_13297);
or U15197 (N_15197,N_14795,N_12820);
and U15198 (N_15198,N_12885,N_13458);
nor U15199 (N_15199,N_12782,N_14530);
nand U15200 (N_15200,N_14501,N_13758);
nor U15201 (N_15201,N_12691,N_14953);
nor U15202 (N_15202,N_14431,N_12814);
nand U15203 (N_15203,N_12918,N_13707);
nand U15204 (N_15204,N_12504,N_14960);
and U15205 (N_15205,N_13283,N_14576);
and U15206 (N_15206,N_12634,N_13282);
nor U15207 (N_15207,N_14858,N_14382);
or U15208 (N_15208,N_13110,N_14307);
or U15209 (N_15209,N_13823,N_12638);
and U15210 (N_15210,N_14610,N_14460);
nor U15211 (N_15211,N_14616,N_13728);
nand U15212 (N_15212,N_14843,N_14274);
and U15213 (N_15213,N_14890,N_13898);
nor U15214 (N_15214,N_12897,N_14869);
nor U15215 (N_15215,N_14064,N_12725);
and U15216 (N_15216,N_13315,N_13644);
nor U15217 (N_15217,N_12523,N_13390);
nor U15218 (N_15218,N_14608,N_14591);
nor U15219 (N_15219,N_14745,N_14273);
or U15220 (N_15220,N_14177,N_14464);
nand U15221 (N_15221,N_14364,N_14979);
and U15222 (N_15222,N_12719,N_14929);
nor U15223 (N_15223,N_13002,N_12541);
or U15224 (N_15224,N_13990,N_14066);
and U15225 (N_15225,N_12827,N_14326);
nand U15226 (N_15226,N_14333,N_14810);
or U15227 (N_15227,N_12985,N_13473);
nor U15228 (N_15228,N_12621,N_13784);
nand U15229 (N_15229,N_14091,N_13704);
or U15230 (N_15230,N_12628,N_13692);
nor U15231 (N_15231,N_13266,N_12547);
nor U15232 (N_15232,N_13798,N_12571);
nor U15233 (N_15233,N_12835,N_13529);
or U15234 (N_15234,N_13027,N_14000);
nand U15235 (N_15235,N_12686,N_14838);
nand U15236 (N_15236,N_12637,N_12603);
and U15237 (N_15237,N_13775,N_13267);
or U15238 (N_15238,N_13655,N_14037);
nor U15239 (N_15239,N_13850,N_13721);
or U15240 (N_15240,N_12752,N_13956);
or U15241 (N_15241,N_13830,N_13578);
nand U15242 (N_15242,N_14754,N_13507);
nor U15243 (N_15243,N_13423,N_14925);
xor U15244 (N_15244,N_14957,N_13522);
or U15245 (N_15245,N_12534,N_14846);
nor U15246 (N_15246,N_14932,N_13593);
nor U15247 (N_15247,N_12701,N_13547);
nor U15248 (N_15248,N_13979,N_14973);
nand U15249 (N_15249,N_14426,N_13481);
or U15250 (N_15250,N_13064,N_14511);
nand U15251 (N_15251,N_14312,N_14285);
or U15252 (N_15252,N_12802,N_12979);
nor U15253 (N_15253,N_14572,N_13012);
nand U15254 (N_15254,N_13968,N_13437);
and U15255 (N_15255,N_13080,N_13006);
and U15256 (N_15256,N_14424,N_14410);
or U15257 (N_15257,N_12581,N_13580);
or U15258 (N_15258,N_12736,N_14031);
xnor U15259 (N_15259,N_14114,N_13822);
nor U15260 (N_15260,N_12798,N_12676);
nand U15261 (N_15261,N_12600,N_14896);
or U15262 (N_15262,N_13188,N_14293);
nor U15263 (N_15263,N_13517,N_13805);
nand U15264 (N_15264,N_13471,N_13882);
or U15265 (N_15265,N_12955,N_14275);
and U15266 (N_15266,N_14463,N_14436);
and U15267 (N_15267,N_13984,N_12549);
nor U15268 (N_15268,N_14531,N_12977);
nand U15269 (N_15269,N_13262,N_14590);
nor U15270 (N_15270,N_14188,N_14124);
and U15271 (N_15271,N_13111,N_13298);
nand U15272 (N_15272,N_14337,N_14653);
nor U15273 (N_15273,N_14880,N_13958);
nor U15274 (N_15274,N_14258,N_14504);
or U15275 (N_15275,N_12871,N_14539);
xnor U15276 (N_15276,N_12793,N_14506);
nor U15277 (N_15277,N_14768,N_12996);
nand U15278 (N_15278,N_13335,N_14912);
and U15279 (N_15279,N_12738,N_14048);
or U15280 (N_15280,N_13668,N_14991);
xor U15281 (N_15281,N_12699,N_14850);
nand U15282 (N_15282,N_13975,N_14695);
and U15283 (N_15283,N_14787,N_14111);
nor U15284 (N_15284,N_12758,N_12674);
nor U15285 (N_15285,N_13989,N_14341);
or U15286 (N_15286,N_13365,N_13193);
nor U15287 (N_15287,N_12645,N_14571);
and U15288 (N_15288,N_13211,N_13075);
and U15289 (N_15289,N_13118,N_13600);
nand U15290 (N_15290,N_13620,N_13029);
or U15291 (N_15291,N_12919,N_14940);
and U15292 (N_15292,N_14938,N_14874);
nor U15293 (N_15293,N_13942,N_12763);
nor U15294 (N_15294,N_13914,N_14672);
nor U15295 (N_15295,N_13957,N_13738);
nor U15296 (N_15296,N_12836,N_14902);
nor U15297 (N_15297,N_13417,N_14569);
and U15298 (N_15298,N_14814,N_12944);
nand U15299 (N_15299,N_14452,N_14607);
nor U15300 (N_15300,N_14253,N_14494);
xor U15301 (N_15301,N_14039,N_13333);
nor U15302 (N_15302,N_14468,N_14903);
and U15303 (N_15303,N_14365,N_13082);
nand U15304 (N_15304,N_13131,N_14913);
and U15305 (N_15305,N_13046,N_13512);
or U15306 (N_15306,N_14521,N_14894);
nand U15307 (N_15307,N_14867,N_14844);
or U15308 (N_15308,N_13385,N_14362);
nand U15309 (N_15309,N_13664,N_14434);
and U15310 (N_15310,N_14908,N_14668);
nor U15311 (N_15311,N_12585,N_12907);
or U15312 (N_15312,N_13648,N_13747);
nand U15313 (N_15313,N_14475,N_12587);
and U15314 (N_15314,N_13888,N_13558);
nor U15315 (N_15315,N_13279,N_14972);
nor U15316 (N_15316,N_14163,N_13053);
and U15317 (N_15317,N_13598,N_14335);
and U15318 (N_15318,N_14655,N_12535);
nand U15319 (N_15319,N_14173,N_13766);
and U15320 (N_15320,N_13576,N_13127);
nand U15321 (N_15321,N_13269,N_13171);
or U15322 (N_15322,N_13233,N_12791);
and U15323 (N_15323,N_13719,N_13531);
or U15324 (N_15324,N_14721,N_13091);
nand U15325 (N_15325,N_13434,N_12927);
and U15326 (N_15326,N_12666,N_14863);
and U15327 (N_15327,N_12935,N_13202);
nor U15328 (N_15328,N_12954,N_14309);
nand U15329 (N_15329,N_13913,N_14816);
and U15330 (N_15330,N_13391,N_14289);
and U15331 (N_15331,N_12680,N_14582);
nor U15332 (N_15332,N_12548,N_13347);
nand U15333 (N_15333,N_13659,N_13594);
and U15334 (N_15334,N_13929,N_12708);
or U15335 (N_15335,N_14292,N_13559);
and U15336 (N_15336,N_13637,N_12558);
nor U15337 (N_15337,N_14428,N_14001);
and U15338 (N_15338,N_14299,N_12599);
nand U15339 (N_15339,N_13606,N_12830);
and U15340 (N_15340,N_14405,N_13778);
nor U15341 (N_15341,N_13919,N_13797);
nor U15342 (N_15342,N_12868,N_14969);
and U15343 (N_15343,N_13412,N_13496);
nand U15344 (N_15344,N_14205,N_13663);
nand U15345 (N_15345,N_14396,N_14612);
nor U15346 (N_15346,N_13383,N_13045);
nor U15347 (N_15347,N_13687,N_12714);
nor U15348 (N_15348,N_14918,N_12959);
nor U15349 (N_15349,N_14856,N_13645);
nor U15350 (N_15350,N_12507,N_12910);
nand U15351 (N_15351,N_13842,N_14974);
nand U15352 (N_15352,N_14761,N_14359);
and U15353 (N_15353,N_12952,N_13883);
and U15354 (N_15354,N_13688,N_14931);
nand U15355 (N_15355,N_12980,N_12553);
nand U15356 (N_15356,N_14387,N_13591);
and U15357 (N_15357,N_13047,N_13794);
and U15358 (N_15358,N_14732,N_14875);
and U15359 (N_15359,N_14817,N_14548);
or U15360 (N_15360,N_13428,N_14551);
or U15361 (N_15361,N_12668,N_14954);
and U15362 (N_15362,N_14835,N_13690);
or U15363 (N_15363,N_14550,N_14499);
xnor U15364 (N_15364,N_13125,N_13691);
and U15365 (N_15365,N_14142,N_14003);
or U15366 (N_15366,N_14097,N_12741);
or U15367 (N_15367,N_12958,N_14284);
or U15368 (N_15368,N_13442,N_14279);
and U15369 (N_15369,N_14704,N_13152);
nand U15370 (N_15370,N_14065,N_13309);
nand U15371 (N_15371,N_12681,N_12784);
and U15372 (N_15372,N_14340,N_13733);
or U15373 (N_15373,N_13489,N_14767);
nand U15374 (N_15374,N_14950,N_13903);
and U15375 (N_15375,N_14842,N_14619);
nand U15376 (N_15376,N_12939,N_14598);
nor U15377 (N_15377,N_14041,N_14492);
nand U15378 (N_15378,N_12500,N_14181);
nor U15379 (N_15379,N_13456,N_14268);
nor U15380 (N_15380,N_13206,N_13014);
xor U15381 (N_15381,N_13499,N_12929);
nand U15382 (N_15382,N_13071,N_14467);
nor U15383 (N_15383,N_12788,N_14697);
and U15384 (N_15384,N_13633,N_14958);
and U15385 (N_15385,N_13555,N_14987);
nand U15386 (N_15386,N_12635,N_12577);
and U15387 (N_15387,N_12822,N_14643);
and U15388 (N_15388,N_13695,N_13485);
nand U15389 (N_15389,N_13677,N_12607);
xnor U15390 (N_15390,N_12533,N_12631);
or U15391 (N_15391,N_14965,N_12527);
and U15392 (N_15392,N_14170,N_14783);
nor U15393 (N_15393,N_13861,N_14314);
or U15394 (N_15394,N_13173,N_13227);
nand U15395 (N_15395,N_14099,N_12678);
and U15396 (N_15396,N_13443,N_12988);
nand U15397 (N_15397,N_13295,N_13562);
or U15398 (N_15398,N_12783,N_12702);
or U15399 (N_15399,N_13465,N_13415);
nand U15400 (N_15400,N_13139,N_12972);
nor U15401 (N_15401,N_14356,N_14617);
nor U15402 (N_15402,N_14226,N_14147);
nand U15403 (N_15403,N_13629,N_12630);
xnor U15404 (N_15404,N_13505,N_14250);
and U15405 (N_15405,N_13154,N_13867);
nand U15406 (N_15406,N_14117,N_13317);
nand U15407 (N_15407,N_14450,N_12532);
xnor U15408 (N_15408,N_13808,N_13683);
nor U15409 (N_15409,N_14507,N_14419);
nor U15410 (N_15410,N_14565,N_14084);
nand U15411 (N_15411,N_14059,N_14241);
nor U15412 (N_15412,N_13346,N_14632);
or U15413 (N_15413,N_13070,N_13085);
nand U15414 (N_15414,N_14961,N_13038);
and U15415 (N_15415,N_14277,N_14693);
nor U15416 (N_15416,N_14063,N_13210);
or U15417 (N_15417,N_14570,N_14100);
or U15418 (N_15418,N_14543,N_14528);
or U15419 (N_15419,N_14865,N_13343);
nand U15420 (N_15420,N_13497,N_14020);
nor U15421 (N_15421,N_14809,N_13431);
nand U15422 (N_15422,N_13162,N_14119);
nor U15423 (N_15423,N_12846,N_14805);
or U15424 (N_15424,N_12757,N_13577);
xor U15425 (N_15425,N_13675,N_13469);
nor U15426 (N_15426,N_14517,N_14136);
nand U15427 (N_15427,N_13628,N_14317);
or U15428 (N_15428,N_13729,N_13985);
or U15429 (N_15429,N_12660,N_14429);
nor U15430 (N_15430,N_13197,N_12539);
nor U15431 (N_15431,N_14461,N_12877);
nand U15432 (N_15432,N_14246,N_12561);
nor U15433 (N_15433,N_14857,N_14301);
nand U15434 (N_15434,N_12563,N_13894);
nor U15435 (N_15435,N_13183,N_13880);
and U15436 (N_15436,N_13063,N_13955);
nand U15437 (N_15437,N_13666,N_13945);
or U15438 (N_15438,N_12886,N_13436);
and U15439 (N_15439,N_14916,N_14515);
or U15440 (N_15440,N_14225,N_13948);
and U15441 (N_15441,N_14736,N_14442);
and U15442 (N_15442,N_13946,N_14295);
and U15443 (N_15443,N_14152,N_13476);
or U15444 (N_15444,N_14889,N_12772);
nor U15445 (N_15445,N_12713,N_14025);
or U15446 (N_15446,N_14252,N_13382);
and U15447 (N_15447,N_13312,N_14547);
nand U15448 (N_15448,N_13932,N_14272);
nand U15449 (N_15449,N_13419,N_14016);
nand U15450 (N_15450,N_14156,N_14516);
nand U15451 (N_15451,N_14160,N_12778);
nor U15452 (N_15452,N_12659,N_14240);
nor U15453 (N_15453,N_14169,N_14634);
nor U15454 (N_15454,N_13095,N_13737);
nor U15455 (N_15455,N_14161,N_13302);
nand U15456 (N_15456,N_14574,N_13701);
or U15457 (N_15457,N_13397,N_14286);
nand U15458 (N_15458,N_12626,N_14801);
or U15459 (N_15459,N_13261,N_14690);
nand U15460 (N_15460,N_14742,N_14623);
nor U15461 (N_15461,N_14308,N_14959);
nand U15462 (N_15462,N_13225,N_13355);
nor U15463 (N_15463,N_13352,N_13746);
and U15464 (N_15464,N_13066,N_13912);
or U15465 (N_15465,N_14189,N_13060);
and U15466 (N_15466,N_13886,N_13967);
nor U15467 (N_15467,N_14249,N_14445);
or U15468 (N_15468,N_12746,N_14741);
nand U15469 (N_15469,N_14725,N_13381);
or U15470 (N_15470,N_14411,N_13518);
and U15471 (N_15471,N_12518,N_14381);
and U15472 (N_15472,N_14942,N_13168);
nand U15473 (N_15473,N_13768,N_14544);
xnor U15474 (N_15474,N_14303,N_13404);
or U15475 (N_15475,N_14679,N_14233);
or U15476 (N_15476,N_13684,N_14128);
or U15477 (N_15477,N_13782,N_13769);
or U15478 (N_15478,N_13491,N_13662);
nor U15479 (N_15479,N_12620,N_14992);
or U15480 (N_15480,N_12705,N_14823);
nor U15481 (N_15481,N_14812,N_13040);
nand U15482 (N_15482,N_13270,N_13748);
or U15483 (N_15483,N_13567,N_14927);
or U15484 (N_15484,N_12987,N_12663);
nor U15485 (N_15485,N_14978,N_14034);
xor U15486 (N_15486,N_14472,N_13506);
or U15487 (N_15487,N_13150,N_13114);
and U15488 (N_15488,N_13103,N_12931);
nor U15489 (N_15489,N_12808,N_13107);
or U15490 (N_15490,N_14343,N_13761);
nand U15491 (N_15491,N_14674,N_13446);
and U15492 (N_15492,N_12971,N_13962);
nand U15493 (N_15493,N_14121,N_12780);
nor U15494 (N_15494,N_14573,N_14510);
nand U15495 (N_15495,N_12914,N_12682);
nor U15496 (N_15496,N_13937,N_13820);
or U15497 (N_15497,N_12917,N_12852);
nor U15498 (N_15498,N_13290,N_12745);
and U15499 (N_15499,N_12995,N_14231);
and U15500 (N_15500,N_13702,N_14853);
nor U15501 (N_15501,N_12508,N_12775);
or U15502 (N_15502,N_13627,N_13917);
or U15503 (N_15503,N_13345,N_14618);
nand U15504 (N_15504,N_13554,N_13199);
and U15505 (N_15505,N_14191,N_14469);
nand U15506 (N_15506,N_13650,N_13549);
nor U15507 (N_15507,N_13875,N_13218);
nor U15508 (N_15508,N_12800,N_14107);
and U15509 (N_15509,N_13061,N_14545);
and U15510 (N_15510,N_14769,N_12734);
nor U15511 (N_15511,N_14133,N_14654);
and U15512 (N_15512,N_14202,N_13477);
nand U15513 (N_15513,N_12616,N_14738);
nor U15514 (N_15514,N_12920,N_14788);
or U15515 (N_15515,N_14917,N_14363);
or U15516 (N_15516,N_13470,N_14456);
and U15517 (N_15517,N_14144,N_13966);
or U15518 (N_15518,N_14885,N_13265);
or U15519 (N_15519,N_14216,N_13970);
nor U15520 (N_15520,N_14955,N_12700);
nor U15521 (N_15521,N_12650,N_12869);
nor U15522 (N_15522,N_13569,N_13167);
nand U15523 (N_15523,N_14800,N_13310);
nor U15524 (N_15524,N_14195,N_13136);
and U15525 (N_15525,N_13504,N_12697);
nand U15526 (N_15526,N_12823,N_14146);
nor U15527 (N_15527,N_14224,N_13273);
nor U15528 (N_15528,N_12943,N_13328);
or U15529 (N_15529,N_13098,N_14698);
or U15530 (N_15530,N_13802,N_13909);
nand U15531 (N_15531,N_14377,N_13851);
and U15532 (N_15532,N_13026,N_12517);
and U15533 (N_15533,N_12712,N_13240);
nor U15534 (N_15534,N_13078,N_12933);
nor U15535 (N_15535,N_14891,N_14239);
or U15536 (N_15536,N_13454,N_14806);
or U15537 (N_15537,N_12913,N_14087);
nor U15538 (N_15538,N_12812,N_13712);
nor U15539 (N_15539,N_13364,N_13122);
and U15540 (N_15540,N_14597,N_14474);
or U15541 (N_15541,N_13978,N_13911);
nor U15542 (N_15542,N_13924,N_14118);
and U15543 (N_15543,N_14562,N_13754);
or U15544 (N_15544,N_13602,N_14397);
nor U15545 (N_15545,N_14321,N_14056);
nor U15546 (N_15546,N_14606,N_12528);
nor U15547 (N_15547,N_12892,N_12916);
xnor U15548 (N_15548,N_13824,N_13034);
or U15549 (N_15549,N_14103,N_14951);
nand U15550 (N_15550,N_14500,N_13899);
and U15551 (N_15551,N_13329,N_14489);
or U15552 (N_15552,N_13587,N_14393);
nand U15553 (N_15553,N_13597,N_14744);
nor U15554 (N_15554,N_13254,N_12968);
or U15555 (N_15555,N_14269,N_13698);
nor U15556 (N_15556,N_13681,N_14373);
nor U15557 (N_15557,N_13104,N_13037);
or U15558 (N_15558,N_14703,N_14581);
or U15559 (N_15559,N_12781,N_14413);
nor U15560 (N_15560,N_12569,N_14082);
xor U15561 (N_15561,N_13949,N_13840);
or U15562 (N_15562,N_14486,N_14692);
or U15563 (N_15563,N_13146,N_13204);
nand U15564 (N_15564,N_14298,N_14069);
nand U15565 (N_15565,N_13189,N_13005);
nor U15566 (N_15566,N_12670,N_14218);
nor U15567 (N_15567,N_14657,N_13185);
and U15568 (N_15568,N_13680,N_14479);
nand U15569 (N_15569,N_14774,N_14906);
nor U15570 (N_15570,N_14423,N_14604);
and U15571 (N_15571,N_13377,N_14193);
nor U15572 (N_15572,N_14023,N_13736);
xor U15573 (N_15573,N_13222,N_14967);
and U15574 (N_15574,N_14757,N_14123);
nand U15575 (N_15575,N_14313,N_14625);
or U15576 (N_15576,N_14101,N_12786);
nor U15577 (N_15577,N_12837,N_12890);
and U15578 (N_15578,N_13931,N_13891);
and U15579 (N_15579,N_13115,N_12870);
and U15580 (N_15580,N_12811,N_13293);
xor U15581 (N_15581,N_13087,N_14388);
and U15582 (N_15582,N_14449,N_13542);
nand U15583 (N_15583,N_14010,N_13307);
nor U15584 (N_15584,N_14443,N_12809);
nand U15585 (N_15585,N_13694,N_14180);
nand U15586 (N_15586,N_13848,N_13546);
and U15587 (N_15587,N_13776,N_14271);
and U15588 (N_15588,N_13271,N_14095);
nand U15589 (N_15589,N_14318,N_14540);
nor U15590 (N_15590,N_13196,N_12703);
nor U15591 (N_15591,N_14714,N_13890);
nor U15592 (N_15592,N_14688,N_12855);
or U15593 (N_15593,N_13124,N_13324);
nand U15594 (N_15594,N_14897,N_13020);
nor U15595 (N_15595,N_13482,N_12888);
and U15596 (N_15596,N_13099,N_14214);
and U15597 (N_15597,N_14132,N_13638);
nor U15598 (N_15598,N_14354,N_13203);
and U15599 (N_15599,N_14311,N_14525);
nand U15600 (N_15600,N_13523,N_13799);
nand U15601 (N_15601,N_14060,N_12740);
and U15602 (N_15602,N_14019,N_14398);
or U15603 (N_15603,N_14667,N_14975);
nor U15604 (N_15604,N_14676,N_13829);
or U15605 (N_15605,N_13963,N_14458);
and U15606 (N_15606,N_12536,N_12502);
nand U15607 (N_15607,N_13141,N_13348);
or U15608 (N_15608,N_13272,N_13964);
nor U15609 (N_15609,N_13134,N_14836);
or U15610 (N_15610,N_14705,N_13615);
and U15611 (N_15611,N_13292,N_13885);
or U15612 (N_15612,N_13818,N_13209);
and U15613 (N_15613,N_14194,N_14635);
nor U15614 (N_15614,N_12595,N_13510);
nor U15615 (N_15615,N_12926,N_14140);
nor U15616 (N_15616,N_14524,N_13285);
nor U15617 (N_15617,N_13947,N_14577);
nand U15618 (N_15618,N_12617,N_14659);
nand U15619 (N_15619,N_14278,N_13671);
nand U15620 (N_15620,N_13639,N_13242);
and U15621 (N_15621,N_13961,N_14686);
or U15622 (N_15622,N_13121,N_13450);
or U15623 (N_15623,N_12908,N_14438);
or U15624 (N_15624,N_12555,N_12875);
nand U15625 (N_15625,N_12596,N_14980);
or U15626 (N_15626,N_12644,N_13256);
or U15627 (N_15627,N_12505,N_12861);
and U15628 (N_15628,N_14148,N_14756);
or U15629 (N_15629,N_14230,N_13674);
and U15630 (N_15630,N_14323,N_14877);
or U15631 (N_15631,N_14137,N_14437);
nand U15632 (N_15632,N_13749,N_14376);
nor U15633 (N_15633,N_13907,N_13514);
or U15634 (N_15634,N_14522,N_12986);
nor U15635 (N_15635,N_13332,N_14030);
or U15636 (N_15636,N_14440,N_14143);
and U15637 (N_15637,N_14542,N_13418);
nor U15638 (N_15638,N_12639,N_13534);
and U15639 (N_15639,N_13440,N_12661);
and U15640 (N_15640,N_13858,N_14172);
and U15641 (N_15641,N_14182,N_14780);
nand U15642 (N_15642,N_12530,N_13259);
nand U15643 (N_15643,N_14855,N_13819);
nand U15644 (N_15644,N_14076,N_14184);
or U15645 (N_15645,N_13807,N_14645);
or U15646 (N_15646,N_13841,N_12729);
nand U15647 (N_15647,N_12860,N_13871);
or U15648 (N_15648,N_13921,N_14683);
nand U15649 (N_15649,N_13552,N_12510);
or U15650 (N_15650,N_12790,N_12576);
and U15651 (N_15651,N_13007,N_13780);
nand U15652 (N_15652,N_13872,N_14716);
or U15653 (N_15653,N_12872,N_14280);
and U15654 (N_15654,N_14159,N_13860);
or U15655 (N_15655,N_13425,N_13526);
or U15656 (N_15656,N_13044,N_13583);
nor U15657 (N_15657,N_14640,N_14027);
or U15658 (N_15658,N_14532,N_13508);
nand U15659 (N_15659,N_13374,N_13795);
or U15660 (N_15660,N_13652,N_12568);
or U15661 (N_15661,N_13057,N_13557);
nor U15662 (N_15662,N_13251,N_14876);
and U15663 (N_15663,N_13612,N_13130);
and U15664 (N_15664,N_12799,N_14666);
nand U15665 (N_15665,N_14920,N_14022);
or U15666 (N_15666,N_14104,N_14167);
xnor U15667 (N_15667,N_12730,N_13280);
nand U15668 (N_15668,N_13969,N_13838);
and U15669 (N_15669,N_14109,N_14728);
and U15670 (N_15670,N_14873,N_14731);
or U15671 (N_15671,N_14678,N_14208);
and U15672 (N_15672,N_13180,N_12774);
or U15673 (N_15673,N_13853,N_12557);
xnor U15674 (N_15674,N_13408,N_14924);
nor U15675 (N_15675,N_14503,N_13994);
nand U15676 (N_15676,N_14491,N_13237);
nand U15677 (N_15677,N_14592,N_13624);
nor U15678 (N_15678,N_13151,N_13498);
nand U15679 (N_15679,N_12841,N_12562);
or U15680 (N_15680,N_14135,N_14092);
or U15681 (N_15681,N_12610,N_13424);
or U15682 (N_15682,N_12656,N_14490);
xnor U15683 (N_15683,N_13642,N_13388);
nand U15684 (N_15684,N_13868,N_14093);
nor U15685 (N_15685,N_13161,N_13379);
nand U15686 (N_15686,N_13301,N_14206);
and U15687 (N_15687,N_12579,N_14122);
nor U15688 (N_15688,N_13021,N_14412);
or U15689 (N_15689,N_14658,N_13714);
nand U15690 (N_15690,N_13181,N_12669);
nand U15691 (N_15691,N_12937,N_14719);
or U15692 (N_15692,N_13447,N_12692);
nor U15693 (N_15693,N_14186,N_12909);
xor U15694 (N_15694,N_14615,N_14596);
nand U15695 (N_15695,N_13208,N_12828);
nor U15696 (N_15696,N_14078,N_14502);
and U15697 (N_15697,N_13068,N_13900);
nand U15698 (N_15698,N_14629,N_12880);
nor U15699 (N_15699,N_12606,N_12520);
nand U15700 (N_15700,N_13892,N_13959);
nor U15701 (N_15701,N_14746,N_14976);
and U15702 (N_15702,N_14427,N_14046);
nand U15703 (N_15703,N_13866,N_14223);
xor U15704 (N_15704,N_12550,N_13157);
nand U15705 (N_15705,N_13941,N_14207);
and U15706 (N_15706,N_13017,N_13592);
and U15707 (N_15707,N_14755,N_14892);
nand U15708 (N_15708,N_13239,N_13462);
nor U15709 (N_15709,N_13411,N_14270);
nor U15710 (N_15710,N_13581,N_13468);
and U15711 (N_15711,N_13828,N_13255);
nor U15712 (N_15712,N_13331,N_12640);
and U15713 (N_15713,N_12978,N_13611);
and U15714 (N_15714,N_14626,N_14328);
nand U15715 (N_15715,N_14859,N_14325);
nor U15716 (N_15716,N_13944,N_13717);
nor U15717 (N_15717,N_13616,N_14771);
nor U15718 (N_15718,N_12779,N_14849);
nand U15719 (N_15719,N_13323,N_13360);
nor U15720 (N_15720,N_13401,N_13113);
or U15721 (N_15721,N_14588,N_13803);
nand U15722 (N_15722,N_12942,N_14294);
and U15723 (N_15723,N_14348,N_12851);
nor U15724 (N_15724,N_13160,N_12721);
nand U15725 (N_15725,N_13621,N_12992);
and U15726 (N_15726,N_14554,N_13405);
and U15727 (N_15727,N_13353,N_13801);
nor U15728 (N_15728,N_14221,N_14071);
nand U15729 (N_15729,N_13635,N_13116);
and U15730 (N_15730,N_13887,N_14149);
or U15731 (N_15731,N_14602,N_12516);
nor U15732 (N_15732,N_13582,N_12894);
nand U15733 (N_15733,N_12608,N_12564);
or U15734 (N_15734,N_12976,N_14455);
or U15735 (N_15735,N_13568,N_12594);
or U15736 (N_15736,N_13041,N_12720);
and U15737 (N_15737,N_14480,N_13706);
and U15738 (N_15738,N_14310,N_13398);
or U15739 (N_15739,N_12759,N_12762);
nand U15740 (N_15740,N_13359,N_13372);
nand U15741 (N_15741,N_13960,N_14514);
nand U15742 (N_15742,N_13308,N_14418);
nand U15743 (N_15743,N_13804,N_14766);
or U15744 (N_15744,N_13158,N_14791);
nor U15745 (N_15745,N_14861,N_14990);
and U15746 (N_15746,N_12932,N_13610);
or U15747 (N_15747,N_12641,N_13682);
or U15748 (N_15748,N_14345,N_14315);
nor U15749 (N_15749,N_12529,N_12813);
and U15750 (N_15750,N_12707,N_13742);
nor U15751 (N_15751,N_14966,N_14351);
and U15752 (N_15752,N_14803,N_12546);
nand U15753 (N_15753,N_14383,N_12934);
or U15754 (N_15754,N_13515,N_14707);
and U15755 (N_15755,N_14662,N_13839);
nand U15756 (N_15756,N_12726,N_12658);
nor U15757 (N_15757,N_13386,N_12593);
or U15758 (N_15758,N_12748,N_14401);
or U15759 (N_15759,N_12969,N_12766);
or U15760 (N_15760,N_12981,N_13195);
and U15761 (N_15761,N_13288,N_13155);
nand U15762 (N_15762,N_14098,N_13521);
or U15763 (N_15763,N_14217,N_13792);
or U15764 (N_15764,N_12690,N_13939);
or U15765 (N_15765,N_13119,N_13922);
or U15766 (N_15766,N_14970,N_14222);
or U15767 (N_15767,N_13934,N_14513);
and U15768 (N_15768,N_13525,N_13023);
or U15769 (N_15769,N_12525,N_13303);
and U15770 (N_15770,N_12856,N_14248);
nand U15771 (N_15771,N_13910,N_14168);
nand U15772 (N_15772,N_14395,N_14709);
or U15773 (N_15773,N_14266,N_13815);
xnor U15774 (N_15774,N_13238,N_14840);
or U15775 (N_15775,N_13320,N_14797);
or U15776 (N_15776,N_14752,N_13334);
and U15777 (N_15777,N_13229,N_13996);
nor U15778 (N_15778,N_13392,N_14711);
nand U15779 (N_15779,N_14447,N_14453);
and U15780 (N_15780,N_14860,N_12818);
and U15781 (N_15781,N_14552,N_14887);
nand U15782 (N_15782,N_14519,N_12711);
nand U15783 (N_15783,N_13837,N_12883);
and U15784 (N_15784,N_12648,N_13362);
nor U15785 (N_15785,N_14051,N_12922);
xnor U15786 (N_15786,N_14886,N_13296);
nor U15787 (N_15787,N_14603,N_14566);
and U15788 (N_15788,N_12696,N_12840);
nor U15789 (N_15789,N_13605,N_13319);
nand U15790 (N_15790,N_12514,N_14720);
and U15791 (N_15791,N_13427,N_14921);
nand U15792 (N_15792,N_13560,N_13551);
xnor U15793 (N_15793,N_13825,N_13182);
xor U15794 (N_15794,N_13263,N_14651);
or U15795 (N_15795,N_13092,N_14043);
and U15796 (N_15796,N_12993,N_12874);
nand U15797 (N_15797,N_14487,N_13864);
nand U15798 (N_15798,N_14009,N_14922);
nand U15799 (N_15799,N_14777,N_13205);
or U15800 (N_15800,N_13884,N_14415);
or U15801 (N_15801,N_13101,N_14158);
or U15802 (N_15802,N_13699,N_13294);
nand U15803 (N_15803,N_12949,N_12771);
nand U15804 (N_15804,N_14560,N_14485);
and U15805 (N_15805,N_13835,N_14905);
or U15806 (N_15806,N_13013,N_14837);
nand U15807 (N_15807,N_13571,N_12960);
nor U15808 (N_15808,N_13847,N_13049);
nor U15809 (N_15809,N_12724,N_12826);
or U15810 (N_15810,N_12857,N_14621);
and U15811 (N_15811,N_13656,N_14481);
xor U15812 (N_15812,N_14360,N_14342);
nand U15813 (N_15813,N_14379,N_14407);
xnor U15814 (N_15814,N_13734,N_14765);
and U15815 (N_15815,N_14579,N_14994);
xor U15816 (N_15816,N_13832,N_13112);
nor U15817 (N_15817,N_13380,N_13954);
and U15818 (N_15818,N_14477,N_14105);
nor U15819 (N_15819,N_13311,N_14989);
nand U15820 (N_15820,N_13223,N_13340);
xnor U15821 (N_15821,N_12754,N_12764);
or U15822 (N_15822,N_14106,N_14935);
nand U15823 (N_15823,N_14234,N_13845);
nor U15824 (N_15824,N_12970,N_13673);
nand U15825 (N_15825,N_12744,N_12649);
or U15826 (N_15826,N_13074,N_14549);
nor U15827 (N_15827,N_13246,N_14465);
nor U15828 (N_15828,N_14004,N_14555);
and U15829 (N_15829,N_14409,N_12776);
and U15830 (N_15830,N_14807,N_14893);
or U15831 (N_15831,N_13865,N_12815);
nor U15832 (N_15832,N_12509,N_13198);
and U15833 (N_15833,N_14049,N_13930);
or U15834 (N_15834,N_13923,N_13607);
nor U15835 (N_15835,N_13877,N_14775);
nor U15836 (N_15836,N_14336,N_13230);
nor U15837 (N_15837,N_12807,N_14864);
nand U15838 (N_15838,N_14808,N_14758);
nor U15839 (N_15839,N_14162,N_14322);
nand U15840 (N_15840,N_13031,N_13762);
nand U15841 (N_15841,N_13166,N_13464);
or U15842 (N_15842,N_13389,N_13741);
nor U15843 (N_15843,N_12858,N_13895);
or U15844 (N_15844,N_13142,N_13918);
or U15845 (N_15845,N_13703,N_12824);
nor U15846 (N_15846,N_14557,N_14793);
and U15847 (N_15847,N_13933,N_13753);
or U15848 (N_15848,N_13354,N_13574);
nand U15849 (N_15849,N_12817,N_13420);
xnor U15850 (N_15850,N_13357,N_14471);
nand U15851 (N_15851,N_13874,N_14282);
nand U15852 (N_15852,N_13553,N_13253);
and U15853 (N_15853,N_13410,N_14238);
nand U15854 (N_15854,N_13079,N_12710);
and U15855 (N_15855,N_14433,N_12899);
nand U15856 (N_15856,N_13678,N_13215);
nand U15857 (N_15857,N_14677,N_14247);
and U15858 (N_15858,N_14828,N_14601);
or U15859 (N_15859,N_13219,N_13527);
or U15860 (N_15860,N_13338,N_14949);
nor U15861 (N_15861,N_14784,N_12706);
or U15862 (N_15862,N_12859,N_12792);
or U15863 (N_15863,N_14567,N_14254);
nor U15864 (N_15864,N_13755,N_13709);
and U15865 (N_15865,N_14523,N_13862);
or U15866 (N_15866,N_14215,N_13519);
nor U15867 (N_15867,N_14933,N_13653);
and U15868 (N_15868,N_13176,N_14002);
or U15869 (N_15869,N_14593,N_13973);
nor U15870 (N_15870,N_12566,N_12966);
and U15871 (N_15871,N_14324,N_13140);
and U15872 (N_15872,N_14778,N_14334);
nor U15873 (N_15873,N_12756,N_13459);
nand U15874 (N_15874,N_12589,N_13787);
nand U15875 (N_15875,N_14026,N_14068);
nor U15876 (N_15876,N_12731,N_14723);
and U15877 (N_15877,N_14520,N_12709);
nor U15878 (N_15878,N_13760,N_14267);
and U15879 (N_15879,N_14717,N_14798);
nor U15880 (N_15880,N_14984,N_12994);
and U15881 (N_15881,N_13938,N_13052);
and U15882 (N_15882,N_13509,N_14753);
or U15883 (N_15883,N_13486,N_13287);
nand U15884 (N_15884,N_12956,N_14211);
nand U15885 (N_15885,N_13276,N_12580);
nand U15886 (N_15886,N_12506,N_14845);
and U15887 (N_15887,N_13756,N_12625);
nand U15888 (N_15888,N_13278,N_13117);
nand U15889 (N_15889,N_13614,N_14639);
nor U15890 (N_15890,N_14011,N_14347);
nand U15891 (N_15891,N_14088,N_14561);
nor U15892 (N_15892,N_14488,N_14178);
nand U15893 (N_15893,N_12543,N_14262);
nand U15894 (N_15894,N_14578,N_13740);
nand U15895 (N_15895,N_14628,N_14518);
nand U15896 (N_15896,N_13474,N_14038);
nor U15897 (N_15897,N_14685,N_14331);
and U15898 (N_15898,N_13943,N_14459);
nor U15899 (N_15899,N_12853,N_14374);
or U15900 (N_15900,N_13413,N_12755);
nand U15901 (N_15901,N_13745,N_14804);
or U15902 (N_15902,N_13164,N_14259);
nand U15903 (N_15903,N_12924,N_14075);
and U15904 (N_15904,N_13976,N_14201);
and U15905 (N_15905,N_12964,N_13433);
nor U15906 (N_15906,N_12647,N_14483);
nand U15907 (N_15907,N_12715,N_14928);
xnor U15908 (N_15908,N_13537,N_14134);
nor U15909 (N_15909,N_14900,N_14045);
and U15910 (N_15910,N_14998,N_13821);
and U15911 (N_15911,N_13777,N_14126);
nand U15912 (N_15912,N_13394,N_12810);
xor U15913 (N_15913,N_13342,N_12804);
xnor U15914 (N_15914,N_13608,N_12983);
and U15915 (N_15915,N_13647,N_12893);
and U15916 (N_15916,N_14304,N_14997);
nor U15917 (N_15917,N_13543,N_13316);
and U15918 (N_15918,N_14699,N_13435);
and U15919 (N_15919,N_13980,N_13585);
nand U15920 (N_15920,N_14174,N_13739);
nor U15921 (N_15921,N_14673,N_13089);
nor U15922 (N_15922,N_13234,N_13178);
nor U15923 (N_15923,N_13953,N_14203);
nor U15924 (N_15924,N_13341,N_13609);
and U15925 (N_15925,N_13480,N_12526);
nand U15926 (N_15926,N_14430,N_14620);
nor U15927 (N_15927,N_12655,N_14013);
nand U15928 (N_15928,N_14153,N_14663);
nor U15929 (N_15929,N_13622,N_13632);
or U15930 (N_15930,N_13207,N_13077);
xnor U15931 (N_15931,N_13870,N_14526);
nand U15932 (N_15932,N_13544,N_14478);
nand U15933 (N_15933,N_14290,N_12673);
nor U15934 (N_15934,N_13565,N_13836);
nand U15935 (N_15935,N_12664,N_13094);
nand U15936 (N_15936,N_13137,N_13284);
or U15937 (N_15937,N_12973,N_14764);
nand U15938 (N_15938,N_14871,N_14713);
nand U15939 (N_15939,N_12849,N_14414);
nand U15940 (N_15940,N_14684,N_12901);
nand U15941 (N_15941,N_12975,N_13987);
xor U15942 (N_15942,N_12560,N_13925);
nor U15943 (N_15943,N_12884,N_12613);
or U15944 (N_15944,N_13076,N_12688);
nand U15945 (N_15945,N_12602,N_14176);
nor U15946 (N_15946,N_12619,N_14316);
nor U15947 (N_15947,N_13813,N_14739);
or U15948 (N_15948,N_12614,N_12761);
nand U15949 (N_15949,N_14151,N_13306);
nand U15950 (N_15950,N_13093,N_12850);
nand U15951 (N_15951,N_14402,N_12575);
and U15952 (N_15952,N_14245,N_12770);
nand U15953 (N_15953,N_12519,N_13438);
nand U15954 (N_15954,N_14212,N_14457);
nand U15955 (N_15955,N_12694,N_14291);
or U15956 (N_15956,N_13086,N_12998);
nor U15957 (N_15957,N_14977,N_12718);
nand U15958 (N_15958,N_12667,N_14081);
and U15959 (N_15959,N_14508,N_13533);
nor U15960 (N_15960,N_14281,N_13676);
nand U15961 (N_15961,N_14911,N_12950);
nand U15962 (N_15962,N_13054,N_13226);
nand U15963 (N_15963,N_12769,N_14297);
nor U15964 (N_15964,N_13500,N_13439);
nor U15965 (N_15965,N_14718,N_13247);
or U15966 (N_15966,N_12570,N_14228);
and U15967 (N_15967,N_12622,N_12524);
and U15968 (N_15968,N_13672,N_14166);
nor U15969 (N_15969,N_12801,N_13708);
and U15970 (N_15970,N_12821,N_13072);
and U15971 (N_15971,N_12834,N_13765);
nand U15972 (N_15972,N_12693,N_12542);
nor U15973 (N_15973,N_12951,N_13539);
or U15974 (N_15974,N_13563,N_14907);
nor U15975 (N_15975,N_14187,N_14664);
or U15976 (N_15976,N_13350,N_13573);
and U15977 (N_15977,N_12559,N_13187);
nor U15978 (N_15978,N_13658,N_13904);
and U15979 (N_15979,N_13492,N_14706);
and U15980 (N_15980,N_14209,N_13088);
and U15981 (N_15981,N_14127,N_13589);
nand U15982 (N_15982,N_14815,N_13339);
nor U15983 (N_15983,N_14422,N_14131);
xnor U15984 (N_15984,N_13952,N_13479);
xor U15985 (N_15985,N_14883,N_13809);
or U15986 (N_15986,N_13000,N_13358);
nand U15987 (N_15987,N_13998,N_13540);
nand U15988 (N_15988,N_13318,N_12551);
or U15989 (N_15989,N_12572,N_12902);
nor U15990 (N_15990,N_14848,N_13796);
or U15991 (N_15991,N_14983,N_12945);
nand U15992 (N_15992,N_14417,N_14824);
nand U15993 (N_15993,N_14792,N_14255);
and U15994 (N_15994,N_14425,N_14366);
nand U15995 (N_15995,N_13727,N_13725);
nor U15996 (N_15996,N_12652,N_12598);
or U15997 (N_15997,N_12512,N_14454);
and U15998 (N_15998,N_14941,N_14986);
nand U15999 (N_15999,N_13743,N_12990);
or U16000 (N_16000,N_12687,N_12967);
nand U16001 (N_16001,N_14829,N_14012);
and U16002 (N_16002,N_12588,N_12675);
and U16003 (N_16003,N_13025,N_14199);
nor U16004 (N_16004,N_13545,N_14884);
or U16005 (N_16005,N_13120,N_12521);
or U16006 (N_16006,N_14375,N_13081);
or U16007 (N_16007,N_14888,N_13897);
or U16008 (N_16008,N_14509,N_13575);
nand U16009 (N_16009,N_12513,N_13457);
nor U16010 (N_16010,N_14014,N_12796);
or U16011 (N_16011,N_14391,N_13463);
nor U16012 (N_16012,N_13143,N_14371);
nand U16013 (N_16013,N_13774,N_12803);
nand U16014 (N_16014,N_13048,N_13096);
and U16015 (N_16015,N_12578,N_14895);
and U16016 (N_16016,N_13194,N_12751);
and U16017 (N_16017,N_13321,N_14689);
and U16018 (N_16018,N_14384,N_14546);
nor U16019 (N_16019,N_12552,N_14394);
or U16020 (N_16020,N_14369,N_13172);
and U16021 (N_16021,N_13455,N_14017);
or U16022 (N_16022,N_13502,N_12684);
nor U16023 (N_16023,N_13313,N_14232);
nor U16024 (N_16024,N_14937,N_13258);
or U16025 (N_16025,N_14150,N_13236);
or U16026 (N_16026,N_13974,N_14914);
or U16027 (N_16027,N_13369,N_14204);
nand U16028 (N_16028,N_14696,N_14702);
nor U16029 (N_16029,N_14276,N_14827);
nand U16030 (N_16030,N_14482,N_13651);
nand U16031 (N_16031,N_13073,N_12930);
nor U16032 (N_16032,N_12923,N_12685);
or U16033 (N_16033,N_14085,N_12806);
nand U16034 (N_16034,N_14110,N_12867);
and U16035 (N_16035,N_12777,N_14355);
or U16036 (N_16036,N_13905,N_13371);
nand U16037 (N_16037,N_13264,N_12601);
and U16038 (N_16038,N_13030,N_13407);
nor U16039 (N_16039,N_12989,N_13816);
nand U16040 (N_16040,N_13997,N_12882);
or U16041 (N_16041,N_14899,N_13192);
and U16042 (N_16042,N_14930,N_12878);
nand U16043 (N_16043,N_12900,N_12854);
or U16044 (N_16044,N_13536,N_13603);
and U16045 (N_16045,N_13351,N_13043);
nand U16046 (N_16046,N_12938,N_13055);
nand U16047 (N_16047,N_13906,N_14236);
or U16048 (N_16048,N_13590,N_14782);
and U16049 (N_16049,N_14682,N_13300);
nor U16050 (N_16050,N_12662,N_12847);
nor U16051 (N_16051,N_13636,N_14054);
nand U16052 (N_16052,N_14263,N_13191);
nand U16053 (N_16053,N_13915,N_14476);
nor U16054 (N_16054,N_13106,N_12816);
and U16055 (N_16055,N_13444,N_13935);
and U16056 (N_16056,N_13561,N_14760);
and U16057 (N_16057,N_12522,N_14251);
or U16058 (N_16058,N_14400,N_13426);
and U16059 (N_16059,N_14473,N_12565);
and U16060 (N_16060,N_13490,N_14370);
nor U16061 (N_16061,N_14630,N_12842);
xor U16062 (N_16062,N_12997,N_14733);
nor U16063 (N_16063,N_13566,N_13723);
or U16064 (N_16064,N_12695,N_14332);
nand U16065 (N_16065,N_12592,N_14390);
and U16066 (N_16066,N_13601,N_13685);
nor U16067 (N_16067,N_13177,N_12965);
nor U16068 (N_16068,N_14353,N_14344);
nand U16069 (N_16069,N_12544,N_12947);
and U16070 (N_16070,N_14432,N_13241);
nand U16071 (N_16071,N_14368,N_12797);
nor U16072 (N_16072,N_14747,N_13982);
or U16073 (N_16073,N_14636,N_14759);
nand U16074 (N_16074,N_14061,N_13129);
and U16075 (N_16075,N_13667,N_13814);
or U16076 (N_16076,N_12540,N_14357);
and U16077 (N_16077,N_13810,N_13416);
nand U16078 (N_16078,N_14671,N_14050);
nor U16079 (N_16079,N_13367,N_14646);
or U16080 (N_16080,N_13378,N_13503);
nor U16081 (N_16081,N_14505,N_14261);
or U16082 (N_16082,N_14822,N_14367);
nor U16083 (N_16083,N_13244,N_14854);
nor U16084 (N_16084,N_14583,N_14790);
and U16085 (N_16085,N_13710,N_14183);
and U16086 (N_16086,N_14493,N_13466);
nor U16087 (N_16087,N_14946,N_14416);
nand U16088 (N_16088,N_14650,N_12946);
nor U16089 (N_16089,N_14497,N_14406);
and U16090 (N_16090,N_14067,N_13854);
or U16091 (N_16091,N_14361,N_14090);
nand U16092 (N_16092,N_13409,N_14287);
or U16093 (N_16093,N_13475,N_12704);
and U16094 (N_16094,N_13373,N_12627);
nand U16095 (N_16095,N_13902,N_13084);
nor U16096 (N_16096,N_13873,N_12632);
or U16097 (N_16097,N_12961,N_14996);
or U16098 (N_16098,N_13445,N_13806);
nor U16099 (N_16099,N_14939,N_13260);
or U16100 (N_16100,N_13018,N_14441);
nor U16101 (N_16101,N_14919,N_14192);
and U16102 (N_16102,N_13105,N_14729);
or U16103 (N_16103,N_13751,N_13790);
xnor U16104 (N_16104,N_13422,N_14024);
or U16105 (N_16105,N_14633,N_13453);
nor U16106 (N_16106,N_13713,N_13487);
nor U16107 (N_16107,N_13812,N_12957);
or U16108 (N_16108,N_12753,N_12591);
nand U16109 (N_16109,N_12911,N_13811);
nand U16110 (N_16110,N_13159,N_12819);
or U16111 (N_16111,N_13001,N_12925);
nor U16112 (N_16112,N_14035,N_13834);
nor U16113 (N_16113,N_13108,N_14963);
nand U16114 (N_16114,N_13878,N_14595);
nor U16115 (N_16115,N_13083,N_14462);
nor U16116 (N_16116,N_13483,N_14649);
nor U16117 (N_16117,N_12915,N_13200);
or U16118 (N_16118,N_13169,N_13617);
nand U16119 (N_16119,N_14349,N_13268);
or U16120 (N_16120,N_12612,N_14631);
nor U16121 (N_16121,N_13596,N_14945);
nand U16122 (N_16122,N_13174,N_14052);
nand U16123 (N_16123,N_13275,N_14535);
and U16124 (N_16124,N_13274,N_14154);
or U16125 (N_16125,N_14210,N_13951);
xor U16126 (N_16126,N_14819,N_13109);
xor U16127 (N_16127,N_12689,N_14044);
nand U16128 (N_16128,N_14799,N_14964);
and U16129 (N_16129,N_14660,N_13752);
and U16130 (N_16130,N_13460,N_13657);
xnor U16131 (N_16131,N_13686,N_14820);
nor U16132 (N_16132,N_14125,N_14962);
and U16133 (N_16133,N_13649,N_12671);
or U16134 (N_16134,N_14070,N_13896);
nand U16135 (N_16135,N_13916,N_12936);
nand U16136 (N_16136,N_13039,N_13869);
or U16137 (N_16137,N_14715,N_14040);
nand U16138 (N_16138,N_13090,N_13186);
nand U16139 (N_16139,N_13735,N_12831);
xor U16140 (N_16140,N_12735,N_12597);
nor U16141 (N_16141,N_13452,N_12760);
and U16142 (N_16142,N_14982,N_12538);
nor U16143 (N_16143,N_13879,N_12646);
nor U16144 (N_16144,N_12737,N_12677);
nor U16145 (N_16145,N_14727,N_14681);
nand U16146 (N_16146,N_14811,N_13732);
or U16147 (N_16147,N_12515,N_14995);
or U16148 (N_16148,N_14926,N_14404);
nand U16149 (N_16149,N_14868,N_13144);
and U16150 (N_16150,N_14327,N_13759);
and U16151 (N_16151,N_14378,N_13451);
nand U16152 (N_16152,N_12727,N_12839);
nand U16153 (N_16153,N_14923,N_12881);
nand U16154 (N_16154,N_13056,N_14826);
or U16155 (N_16155,N_14512,N_13361);
or U16156 (N_16156,N_13999,N_14288);
or U16157 (N_16157,N_14237,N_14265);
nor U16158 (N_16158,N_12829,N_12629);
and U16159 (N_16159,N_12787,N_13231);
or U16160 (N_16160,N_12723,N_12722);
xor U16161 (N_16161,N_13478,N_14242);
nand U16162 (N_16162,N_14086,N_14451);
or U16163 (N_16163,N_13588,N_13286);
and U16164 (N_16164,N_14870,N_12953);
nor U16165 (N_16165,N_13384,N_13846);
or U16166 (N_16166,N_14852,N_13785);
nor U16167 (N_16167,N_12843,N_13214);
nor U16168 (N_16168,N_13643,N_14235);
nand U16169 (N_16169,N_14847,N_14832);
or U16170 (N_16170,N_12573,N_13757);
xor U16171 (N_16171,N_14072,N_14120);
or U16172 (N_16172,N_14130,N_13513);
and U16173 (N_16173,N_14575,N_13550);
or U16174 (N_16174,N_13175,N_14587);
or U16175 (N_16175,N_13432,N_12865);
nand U16176 (N_16176,N_13145,N_14968);
and U16177 (N_16177,N_13003,N_12903);
nor U16178 (N_16178,N_13718,N_13619);
nand U16179 (N_16179,N_12698,N_12863);
xor U16180 (N_16180,N_12503,N_12651);
or U16181 (N_16181,N_14094,N_13516);
nor U16182 (N_16182,N_12848,N_14058);
and U16183 (N_16183,N_14358,N_14089);
or U16184 (N_16184,N_13281,N_12768);
or U16185 (N_16185,N_14005,N_13024);
or U16186 (N_16186,N_13586,N_12982);
or U16187 (N_16187,N_13123,N_13165);
and U16188 (N_16188,N_14813,N_12895);
nand U16189 (N_16189,N_13626,N_14644);
or U16190 (N_16190,N_14881,N_14763);
nor U16191 (N_16191,N_13501,N_13028);
and U16192 (N_16192,N_14057,N_14661);
nand U16193 (N_16193,N_13201,N_13852);
nand U16194 (N_16194,N_12962,N_13033);
and U16195 (N_16195,N_12749,N_14213);
nand U16196 (N_16196,N_12838,N_13212);
or U16197 (N_16197,N_14675,N_12590);
or U16198 (N_16198,N_13788,N_14947);
nor U16199 (N_16199,N_14952,N_13538);
and U16200 (N_16200,N_12912,N_14074);
and U16201 (N_16201,N_14007,N_12866);
xnor U16202 (N_16202,N_13541,N_12728);
or U16203 (N_16203,N_14444,N_12742);
nor U16204 (N_16204,N_14691,N_12657);
nor U16205 (N_16205,N_13325,N_13720);
xnor U16206 (N_16206,N_14585,N_14710);
nor U16207 (N_16207,N_13772,N_14748);
or U16208 (N_16208,N_14385,N_14036);
nor U16209 (N_16209,N_12905,N_13833);
and U16210 (N_16210,N_14985,N_14670);
nand U16211 (N_16211,N_13770,N_14833);
nand U16212 (N_16212,N_14559,N_14734);
nand U16213 (N_16213,N_13396,N_14197);
nor U16214 (N_16214,N_14008,N_13249);
nor U16215 (N_16215,N_13036,N_13179);
and U16216 (N_16216,N_13827,N_14779);
nor U16217 (N_16217,N_12940,N_13623);
and U16218 (N_16218,N_13243,N_13375);
and U16219 (N_16219,N_13102,N_12785);
nor U16220 (N_16220,N_13856,N_13779);
and U16221 (N_16221,N_12537,N_13716);
and U16222 (N_16222,N_13789,N_13022);
nand U16223 (N_16223,N_13356,N_13781);
nand U16224 (N_16224,N_13097,N_14773);
or U16225 (N_16225,N_14600,N_13370);
and U16226 (N_16226,N_14283,N_14680);
nand U16227 (N_16227,N_13584,N_13530);
nand U16228 (N_16228,N_13402,N_14879);
and U16229 (N_16229,N_14841,N_13135);
nor U16230 (N_16230,N_12879,N_12611);
nand U16231 (N_16231,N_14862,N_12624);
nand U16232 (N_16232,N_13363,N_14611);
nand U16233 (N_16233,N_13705,N_14872);
nor U16234 (N_16234,N_14260,N_12873);
nand U16235 (N_16235,N_13711,N_13731);
nor U16236 (N_16236,N_13893,N_13991);
or U16237 (N_16237,N_12887,N_13908);
nor U16238 (N_16238,N_13564,N_13843);
or U16239 (N_16239,N_13700,N_13327);
and U16240 (N_16240,N_13217,N_14724);
nand U16241 (N_16241,N_14352,N_13679);
nand U16242 (N_16242,N_13430,N_13826);
nand U16243 (N_16243,N_12574,N_14296);
xor U16244 (N_16244,N_13190,N_13965);
nand U16245 (N_16245,N_14196,N_14553);
xor U16246 (N_16246,N_13857,N_14988);
nand U16247 (N_16247,N_13170,N_12794);
nor U16248 (N_16248,N_13314,N_14338);
nand U16249 (N_16249,N_14029,N_14403);
xnor U16250 (N_16250,N_14889,N_12944);
or U16251 (N_16251,N_14399,N_13653);
and U16252 (N_16252,N_13358,N_13396);
and U16253 (N_16253,N_13478,N_14784);
nand U16254 (N_16254,N_13115,N_13901);
and U16255 (N_16255,N_14651,N_14660);
nor U16256 (N_16256,N_13239,N_13867);
nor U16257 (N_16257,N_13930,N_14318);
nand U16258 (N_16258,N_13254,N_13516);
or U16259 (N_16259,N_12862,N_13496);
nor U16260 (N_16260,N_14881,N_13592);
or U16261 (N_16261,N_14292,N_13060);
nor U16262 (N_16262,N_14401,N_14428);
or U16263 (N_16263,N_12581,N_13171);
or U16264 (N_16264,N_13572,N_14729);
nor U16265 (N_16265,N_14499,N_13869);
or U16266 (N_16266,N_14006,N_14757);
nand U16267 (N_16267,N_13709,N_12794);
nand U16268 (N_16268,N_14716,N_12757);
and U16269 (N_16269,N_13426,N_12731);
nand U16270 (N_16270,N_14749,N_13177);
or U16271 (N_16271,N_12856,N_14643);
or U16272 (N_16272,N_12545,N_13905);
nor U16273 (N_16273,N_14305,N_12747);
nor U16274 (N_16274,N_13328,N_14837);
or U16275 (N_16275,N_13351,N_13863);
nor U16276 (N_16276,N_13724,N_13484);
xor U16277 (N_16277,N_14747,N_12645);
nor U16278 (N_16278,N_12564,N_13023);
or U16279 (N_16279,N_12598,N_14061);
and U16280 (N_16280,N_13679,N_13168);
nor U16281 (N_16281,N_14675,N_14054);
or U16282 (N_16282,N_14882,N_13336);
nand U16283 (N_16283,N_14791,N_13243);
or U16284 (N_16284,N_14378,N_14520);
and U16285 (N_16285,N_13160,N_14599);
nor U16286 (N_16286,N_12660,N_14868);
nor U16287 (N_16287,N_12641,N_12680);
or U16288 (N_16288,N_14543,N_14850);
or U16289 (N_16289,N_13612,N_12941);
or U16290 (N_16290,N_12601,N_14948);
or U16291 (N_16291,N_13286,N_14487);
and U16292 (N_16292,N_13055,N_12685);
nor U16293 (N_16293,N_14342,N_12705);
nor U16294 (N_16294,N_13497,N_12920);
nor U16295 (N_16295,N_12728,N_13852);
or U16296 (N_16296,N_13668,N_14398);
nor U16297 (N_16297,N_13972,N_13448);
nor U16298 (N_16298,N_13008,N_13601);
nand U16299 (N_16299,N_13745,N_14093);
nand U16300 (N_16300,N_14764,N_14989);
nor U16301 (N_16301,N_14221,N_14537);
and U16302 (N_16302,N_13500,N_14591);
nor U16303 (N_16303,N_14526,N_14481);
or U16304 (N_16304,N_12861,N_14351);
nor U16305 (N_16305,N_14798,N_14982);
and U16306 (N_16306,N_12696,N_13439);
nor U16307 (N_16307,N_13427,N_12761);
xnor U16308 (N_16308,N_14187,N_14278);
xor U16309 (N_16309,N_13196,N_14978);
nand U16310 (N_16310,N_13932,N_14752);
or U16311 (N_16311,N_12797,N_13715);
nor U16312 (N_16312,N_12905,N_12928);
and U16313 (N_16313,N_13889,N_14666);
nand U16314 (N_16314,N_13214,N_14090);
and U16315 (N_16315,N_13130,N_13509);
nand U16316 (N_16316,N_13214,N_12776);
nor U16317 (N_16317,N_13026,N_14498);
nand U16318 (N_16318,N_12550,N_14309);
or U16319 (N_16319,N_14570,N_13714);
nand U16320 (N_16320,N_13454,N_13969);
nor U16321 (N_16321,N_12950,N_13963);
nand U16322 (N_16322,N_14737,N_13622);
or U16323 (N_16323,N_14974,N_14124);
nand U16324 (N_16324,N_12545,N_12723);
and U16325 (N_16325,N_13539,N_12642);
or U16326 (N_16326,N_14620,N_13519);
or U16327 (N_16327,N_14329,N_13010);
or U16328 (N_16328,N_14777,N_13711);
nor U16329 (N_16329,N_14661,N_13639);
and U16330 (N_16330,N_13376,N_13195);
or U16331 (N_16331,N_14275,N_14566);
xnor U16332 (N_16332,N_14479,N_14887);
nor U16333 (N_16333,N_14958,N_14802);
nor U16334 (N_16334,N_12741,N_14029);
nand U16335 (N_16335,N_13060,N_14608);
and U16336 (N_16336,N_12953,N_13141);
nand U16337 (N_16337,N_12893,N_13923);
and U16338 (N_16338,N_13848,N_12541);
nand U16339 (N_16339,N_14460,N_14314);
xor U16340 (N_16340,N_14402,N_14976);
nand U16341 (N_16341,N_13602,N_12884);
nor U16342 (N_16342,N_12856,N_14348);
or U16343 (N_16343,N_12819,N_13356);
or U16344 (N_16344,N_14264,N_14639);
nand U16345 (N_16345,N_12990,N_13073);
nand U16346 (N_16346,N_14323,N_14900);
or U16347 (N_16347,N_13575,N_14484);
nand U16348 (N_16348,N_13283,N_14869);
nor U16349 (N_16349,N_13109,N_13240);
nor U16350 (N_16350,N_14985,N_13957);
nand U16351 (N_16351,N_14742,N_13330);
nand U16352 (N_16352,N_13455,N_14115);
nor U16353 (N_16353,N_14596,N_14946);
and U16354 (N_16354,N_14121,N_13696);
nand U16355 (N_16355,N_13618,N_14207);
or U16356 (N_16356,N_12708,N_13374);
or U16357 (N_16357,N_13250,N_12947);
nor U16358 (N_16358,N_12977,N_13524);
nor U16359 (N_16359,N_13436,N_13566);
nor U16360 (N_16360,N_14221,N_14731);
nor U16361 (N_16361,N_12538,N_13294);
and U16362 (N_16362,N_13178,N_14072);
or U16363 (N_16363,N_13981,N_14982);
and U16364 (N_16364,N_13729,N_14555);
or U16365 (N_16365,N_13889,N_14285);
and U16366 (N_16366,N_13437,N_14121);
or U16367 (N_16367,N_13630,N_13747);
nor U16368 (N_16368,N_12683,N_13411);
xor U16369 (N_16369,N_12998,N_14599);
and U16370 (N_16370,N_13399,N_14590);
or U16371 (N_16371,N_12628,N_14799);
nor U16372 (N_16372,N_13789,N_13475);
nand U16373 (N_16373,N_13596,N_13114);
and U16374 (N_16374,N_14200,N_14604);
nor U16375 (N_16375,N_13300,N_12553);
nor U16376 (N_16376,N_12978,N_13087);
nand U16377 (N_16377,N_13786,N_14883);
nor U16378 (N_16378,N_13664,N_13196);
and U16379 (N_16379,N_13331,N_14690);
or U16380 (N_16380,N_13402,N_14700);
nor U16381 (N_16381,N_12609,N_12503);
and U16382 (N_16382,N_14459,N_13566);
and U16383 (N_16383,N_12878,N_12905);
and U16384 (N_16384,N_14032,N_12653);
nor U16385 (N_16385,N_13878,N_14425);
nand U16386 (N_16386,N_12540,N_12775);
and U16387 (N_16387,N_14705,N_14398);
and U16388 (N_16388,N_13911,N_14318);
and U16389 (N_16389,N_13053,N_13413);
nor U16390 (N_16390,N_14756,N_13958);
or U16391 (N_16391,N_12614,N_13302);
and U16392 (N_16392,N_12636,N_13432);
nor U16393 (N_16393,N_13188,N_13733);
nand U16394 (N_16394,N_12830,N_14943);
nor U16395 (N_16395,N_14729,N_13178);
or U16396 (N_16396,N_13714,N_13450);
and U16397 (N_16397,N_12613,N_14756);
or U16398 (N_16398,N_13345,N_13997);
and U16399 (N_16399,N_14940,N_12836);
xor U16400 (N_16400,N_14257,N_12990);
nor U16401 (N_16401,N_13402,N_13679);
nand U16402 (N_16402,N_14301,N_14958);
or U16403 (N_16403,N_14158,N_14699);
nand U16404 (N_16404,N_13695,N_14532);
nor U16405 (N_16405,N_13336,N_12785);
nor U16406 (N_16406,N_12645,N_14511);
and U16407 (N_16407,N_12928,N_13736);
or U16408 (N_16408,N_14360,N_13671);
or U16409 (N_16409,N_13235,N_14080);
or U16410 (N_16410,N_13876,N_12922);
and U16411 (N_16411,N_14871,N_12899);
or U16412 (N_16412,N_13694,N_14031);
xor U16413 (N_16413,N_14774,N_14250);
and U16414 (N_16414,N_13118,N_14849);
nor U16415 (N_16415,N_14436,N_14011);
or U16416 (N_16416,N_14447,N_14059);
and U16417 (N_16417,N_14668,N_13721);
or U16418 (N_16418,N_13441,N_12567);
or U16419 (N_16419,N_14376,N_12833);
or U16420 (N_16420,N_13851,N_14517);
and U16421 (N_16421,N_12953,N_13593);
nor U16422 (N_16422,N_13019,N_12782);
nand U16423 (N_16423,N_14820,N_12901);
nor U16424 (N_16424,N_12759,N_12738);
nor U16425 (N_16425,N_13834,N_14802);
nand U16426 (N_16426,N_13724,N_14183);
nor U16427 (N_16427,N_13428,N_14601);
and U16428 (N_16428,N_14038,N_12967);
nand U16429 (N_16429,N_12734,N_13259);
nand U16430 (N_16430,N_13855,N_12544);
or U16431 (N_16431,N_14022,N_14830);
nand U16432 (N_16432,N_13572,N_13363);
nand U16433 (N_16433,N_14619,N_13902);
nor U16434 (N_16434,N_14263,N_13800);
and U16435 (N_16435,N_14651,N_14080);
or U16436 (N_16436,N_13723,N_14852);
nand U16437 (N_16437,N_14081,N_12580);
or U16438 (N_16438,N_14139,N_14374);
or U16439 (N_16439,N_13770,N_13607);
or U16440 (N_16440,N_13566,N_14152);
or U16441 (N_16441,N_13494,N_13122);
or U16442 (N_16442,N_14710,N_14029);
nor U16443 (N_16443,N_12801,N_12737);
nor U16444 (N_16444,N_14249,N_14680);
nor U16445 (N_16445,N_12534,N_14045);
or U16446 (N_16446,N_14751,N_14283);
and U16447 (N_16447,N_13431,N_13674);
or U16448 (N_16448,N_14145,N_13842);
xnor U16449 (N_16449,N_14288,N_14999);
and U16450 (N_16450,N_14054,N_13278);
and U16451 (N_16451,N_13565,N_14803);
or U16452 (N_16452,N_14704,N_14007);
or U16453 (N_16453,N_13348,N_14946);
or U16454 (N_16454,N_14558,N_14436);
or U16455 (N_16455,N_14480,N_13414);
nor U16456 (N_16456,N_12538,N_14936);
or U16457 (N_16457,N_13199,N_12591);
nor U16458 (N_16458,N_13043,N_13327);
and U16459 (N_16459,N_13920,N_13114);
and U16460 (N_16460,N_14431,N_13593);
nor U16461 (N_16461,N_13433,N_13424);
nand U16462 (N_16462,N_13561,N_14481);
or U16463 (N_16463,N_12928,N_13945);
and U16464 (N_16464,N_13891,N_13221);
or U16465 (N_16465,N_14704,N_13537);
nor U16466 (N_16466,N_13986,N_14485);
nand U16467 (N_16467,N_14838,N_14072);
and U16468 (N_16468,N_14083,N_14499);
and U16469 (N_16469,N_13203,N_14161);
or U16470 (N_16470,N_14401,N_13398);
nor U16471 (N_16471,N_14000,N_12677);
nor U16472 (N_16472,N_14831,N_14915);
nor U16473 (N_16473,N_12625,N_13422);
xnor U16474 (N_16474,N_13758,N_14297);
or U16475 (N_16475,N_14723,N_14462);
nand U16476 (N_16476,N_12711,N_14958);
nand U16477 (N_16477,N_13437,N_12797);
and U16478 (N_16478,N_14801,N_14020);
nor U16479 (N_16479,N_14770,N_14240);
nand U16480 (N_16480,N_12784,N_13586);
and U16481 (N_16481,N_14018,N_14430);
or U16482 (N_16482,N_13921,N_14324);
or U16483 (N_16483,N_12831,N_14030);
nand U16484 (N_16484,N_12846,N_13845);
and U16485 (N_16485,N_14197,N_13777);
and U16486 (N_16486,N_13955,N_14727);
or U16487 (N_16487,N_14111,N_14027);
and U16488 (N_16488,N_14675,N_14993);
and U16489 (N_16489,N_14325,N_14526);
nand U16490 (N_16490,N_14952,N_13380);
nor U16491 (N_16491,N_14963,N_13307);
nor U16492 (N_16492,N_13911,N_14609);
and U16493 (N_16493,N_12512,N_14771);
or U16494 (N_16494,N_13763,N_13046);
xnor U16495 (N_16495,N_13777,N_13094);
and U16496 (N_16496,N_14632,N_12506);
nor U16497 (N_16497,N_14584,N_13856);
or U16498 (N_16498,N_13131,N_13274);
and U16499 (N_16499,N_13089,N_14339);
or U16500 (N_16500,N_12566,N_12755);
or U16501 (N_16501,N_14317,N_13218);
or U16502 (N_16502,N_13360,N_13927);
nand U16503 (N_16503,N_14798,N_14026);
or U16504 (N_16504,N_14850,N_14292);
nand U16505 (N_16505,N_14171,N_13620);
nand U16506 (N_16506,N_13759,N_13264);
nor U16507 (N_16507,N_12582,N_12974);
and U16508 (N_16508,N_13052,N_14043);
nand U16509 (N_16509,N_13972,N_12512);
nand U16510 (N_16510,N_13336,N_14583);
nand U16511 (N_16511,N_13920,N_14090);
or U16512 (N_16512,N_14487,N_12559);
or U16513 (N_16513,N_13370,N_13364);
nand U16514 (N_16514,N_12643,N_13955);
xor U16515 (N_16515,N_13563,N_14377);
and U16516 (N_16516,N_13878,N_12973);
or U16517 (N_16517,N_12859,N_14357);
or U16518 (N_16518,N_13294,N_13760);
nand U16519 (N_16519,N_13923,N_13209);
and U16520 (N_16520,N_14553,N_12787);
nand U16521 (N_16521,N_13929,N_14456);
nor U16522 (N_16522,N_13858,N_14684);
nor U16523 (N_16523,N_14975,N_13706);
xor U16524 (N_16524,N_14830,N_12645);
nand U16525 (N_16525,N_13114,N_14630);
or U16526 (N_16526,N_14045,N_14669);
xor U16527 (N_16527,N_13523,N_12948);
nor U16528 (N_16528,N_13452,N_14894);
nand U16529 (N_16529,N_14430,N_13604);
and U16530 (N_16530,N_13052,N_13085);
and U16531 (N_16531,N_12792,N_14528);
or U16532 (N_16532,N_13312,N_14316);
nor U16533 (N_16533,N_14543,N_14295);
nand U16534 (N_16534,N_13356,N_13766);
nor U16535 (N_16535,N_13092,N_12818);
nand U16536 (N_16536,N_13482,N_13863);
nor U16537 (N_16537,N_13500,N_14471);
and U16538 (N_16538,N_13132,N_13857);
nand U16539 (N_16539,N_13610,N_13438);
and U16540 (N_16540,N_13139,N_12726);
nor U16541 (N_16541,N_14285,N_14695);
and U16542 (N_16542,N_14402,N_14267);
and U16543 (N_16543,N_12622,N_13070);
and U16544 (N_16544,N_13031,N_13005);
nor U16545 (N_16545,N_12910,N_13659);
or U16546 (N_16546,N_12818,N_14101);
and U16547 (N_16547,N_14064,N_13174);
and U16548 (N_16548,N_12724,N_14287);
nor U16549 (N_16549,N_14114,N_12516);
or U16550 (N_16550,N_14179,N_14084);
or U16551 (N_16551,N_12746,N_14064);
nand U16552 (N_16552,N_12724,N_14899);
or U16553 (N_16553,N_14013,N_14681);
or U16554 (N_16554,N_14256,N_14976);
and U16555 (N_16555,N_14223,N_13651);
and U16556 (N_16556,N_14744,N_14422);
and U16557 (N_16557,N_13550,N_14831);
nand U16558 (N_16558,N_14731,N_12663);
nor U16559 (N_16559,N_13877,N_13509);
nand U16560 (N_16560,N_13736,N_12949);
nand U16561 (N_16561,N_14040,N_14430);
or U16562 (N_16562,N_14371,N_13268);
and U16563 (N_16563,N_12725,N_14462);
nor U16564 (N_16564,N_13024,N_14684);
nand U16565 (N_16565,N_13520,N_14691);
xor U16566 (N_16566,N_14522,N_12720);
or U16567 (N_16567,N_13363,N_13966);
or U16568 (N_16568,N_14048,N_13190);
or U16569 (N_16569,N_12852,N_14224);
nor U16570 (N_16570,N_14253,N_13989);
nor U16571 (N_16571,N_14986,N_13208);
or U16572 (N_16572,N_14128,N_13605);
or U16573 (N_16573,N_13049,N_13287);
and U16574 (N_16574,N_14744,N_12824);
nor U16575 (N_16575,N_14420,N_12965);
nor U16576 (N_16576,N_14025,N_12988);
and U16577 (N_16577,N_14144,N_13047);
nand U16578 (N_16578,N_14984,N_12937);
nor U16579 (N_16579,N_13528,N_13878);
nand U16580 (N_16580,N_14488,N_12502);
or U16581 (N_16581,N_14989,N_12824);
nor U16582 (N_16582,N_13902,N_12683);
nand U16583 (N_16583,N_14324,N_13313);
nand U16584 (N_16584,N_14297,N_14041);
or U16585 (N_16585,N_13674,N_14957);
nor U16586 (N_16586,N_13617,N_13258);
or U16587 (N_16587,N_14357,N_12935);
nand U16588 (N_16588,N_14165,N_13637);
or U16589 (N_16589,N_12953,N_13754);
nor U16590 (N_16590,N_12864,N_12735);
nand U16591 (N_16591,N_13402,N_13474);
or U16592 (N_16592,N_14301,N_12605);
nand U16593 (N_16593,N_13749,N_13698);
nor U16594 (N_16594,N_13929,N_14409);
nand U16595 (N_16595,N_13180,N_14265);
or U16596 (N_16596,N_13060,N_14103);
or U16597 (N_16597,N_13330,N_13877);
and U16598 (N_16598,N_13894,N_13980);
or U16599 (N_16599,N_13848,N_14143);
or U16600 (N_16600,N_13186,N_14280);
or U16601 (N_16601,N_13720,N_13931);
or U16602 (N_16602,N_12689,N_14877);
nor U16603 (N_16603,N_13273,N_13063);
or U16604 (N_16604,N_14388,N_13352);
and U16605 (N_16605,N_14664,N_13406);
nand U16606 (N_16606,N_12981,N_13544);
nor U16607 (N_16607,N_13737,N_13247);
or U16608 (N_16608,N_14105,N_12962);
nand U16609 (N_16609,N_12625,N_13763);
nand U16610 (N_16610,N_12539,N_13268);
or U16611 (N_16611,N_14046,N_13528);
nand U16612 (N_16612,N_13741,N_12668);
or U16613 (N_16613,N_12534,N_14845);
or U16614 (N_16614,N_13347,N_13490);
nor U16615 (N_16615,N_14381,N_13617);
and U16616 (N_16616,N_13074,N_12735);
nand U16617 (N_16617,N_13698,N_14128);
and U16618 (N_16618,N_13014,N_13450);
nor U16619 (N_16619,N_13540,N_13121);
nor U16620 (N_16620,N_13059,N_13909);
nand U16621 (N_16621,N_14096,N_12968);
and U16622 (N_16622,N_14855,N_14519);
and U16623 (N_16623,N_12521,N_14377);
or U16624 (N_16624,N_13617,N_12500);
nor U16625 (N_16625,N_14814,N_13102);
nor U16626 (N_16626,N_12824,N_12565);
and U16627 (N_16627,N_12775,N_12744);
nand U16628 (N_16628,N_14890,N_13750);
nand U16629 (N_16629,N_13977,N_14341);
and U16630 (N_16630,N_14820,N_14828);
or U16631 (N_16631,N_14822,N_13020);
and U16632 (N_16632,N_13512,N_13824);
or U16633 (N_16633,N_12664,N_14266);
and U16634 (N_16634,N_13489,N_13745);
and U16635 (N_16635,N_13300,N_14775);
nor U16636 (N_16636,N_14697,N_13494);
nor U16637 (N_16637,N_13870,N_13534);
or U16638 (N_16638,N_13934,N_14978);
or U16639 (N_16639,N_13366,N_14094);
and U16640 (N_16640,N_12934,N_13972);
and U16641 (N_16641,N_14783,N_12799);
and U16642 (N_16642,N_12808,N_14889);
nor U16643 (N_16643,N_14892,N_13813);
nand U16644 (N_16644,N_13912,N_14609);
or U16645 (N_16645,N_12640,N_14012);
or U16646 (N_16646,N_12681,N_13501);
nand U16647 (N_16647,N_13262,N_13778);
or U16648 (N_16648,N_13709,N_14955);
and U16649 (N_16649,N_13008,N_13890);
nor U16650 (N_16650,N_12719,N_14121);
xnor U16651 (N_16651,N_13692,N_13901);
nand U16652 (N_16652,N_13451,N_13876);
and U16653 (N_16653,N_14653,N_14229);
or U16654 (N_16654,N_14738,N_12734);
nor U16655 (N_16655,N_14280,N_13455);
or U16656 (N_16656,N_14421,N_13277);
or U16657 (N_16657,N_13524,N_12595);
nand U16658 (N_16658,N_13867,N_14041);
and U16659 (N_16659,N_14033,N_14878);
nand U16660 (N_16660,N_13236,N_13470);
and U16661 (N_16661,N_12983,N_13431);
or U16662 (N_16662,N_13926,N_14794);
and U16663 (N_16663,N_14225,N_12806);
nor U16664 (N_16664,N_13111,N_13950);
nor U16665 (N_16665,N_13069,N_14750);
and U16666 (N_16666,N_14608,N_13829);
xnor U16667 (N_16667,N_13502,N_14973);
nand U16668 (N_16668,N_13068,N_13999);
nand U16669 (N_16669,N_13610,N_14248);
or U16670 (N_16670,N_13350,N_14765);
nand U16671 (N_16671,N_12730,N_13976);
and U16672 (N_16672,N_12854,N_14490);
and U16673 (N_16673,N_12501,N_13460);
and U16674 (N_16674,N_13987,N_14380);
and U16675 (N_16675,N_14438,N_14485);
nor U16676 (N_16676,N_13514,N_14060);
or U16677 (N_16677,N_14216,N_14061);
nor U16678 (N_16678,N_12962,N_14132);
nand U16679 (N_16679,N_13026,N_13245);
or U16680 (N_16680,N_14619,N_13598);
nand U16681 (N_16681,N_14149,N_12946);
nand U16682 (N_16682,N_13443,N_13515);
and U16683 (N_16683,N_14188,N_14413);
and U16684 (N_16684,N_14407,N_13541);
or U16685 (N_16685,N_13434,N_13951);
or U16686 (N_16686,N_14056,N_13428);
nor U16687 (N_16687,N_13363,N_13921);
and U16688 (N_16688,N_12668,N_14642);
or U16689 (N_16689,N_14855,N_13032);
nand U16690 (N_16690,N_13495,N_13637);
and U16691 (N_16691,N_13273,N_13223);
nand U16692 (N_16692,N_14071,N_12586);
or U16693 (N_16693,N_13920,N_13217);
or U16694 (N_16694,N_13524,N_12616);
nor U16695 (N_16695,N_14940,N_13838);
or U16696 (N_16696,N_14540,N_14543);
nand U16697 (N_16697,N_12954,N_13166);
nand U16698 (N_16698,N_14033,N_13968);
or U16699 (N_16699,N_13452,N_14412);
nor U16700 (N_16700,N_13253,N_14924);
nand U16701 (N_16701,N_12586,N_13332);
nor U16702 (N_16702,N_13635,N_13170);
or U16703 (N_16703,N_14994,N_14021);
nor U16704 (N_16704,N_13837,N_13975);
or U16705 (N_16705,N_13592,N_12748);
or U16706 (N_16706,N_12710,N_14361);
and U16707 (N_16707,N_13945,N_14625);
and U16708 (N_16708,N_14925,N_13669);
nor U16709 (N_16709,N_14065,N_14194);
nor U16710 (N_16710,N_14760,N_13179);
or U16711 (N_16711,N_14959,N_13084);
nand U16712 (N_16712,N_13265,N_12726);
nand U16713 (N_16713,N_12731,N_14643);
or U16714 (N_16714,N_13775,N_14801);
nor U16715 (N_16715,N_12801,N_14206);
nor U16716 (N_16716,N_14754,N_12828);
nor U16717 (N_16717,N_12986,N_13923);
or U16718 (N_16718,N_14889,N_13674);
nor U16719 (N_16719,N_12987,N_12886);
or U16720 (N_16720,N_13879,N_12728);
and U16721 (N_16721,N_12917,N_12934);
or U16722 (N_16722,N_14228,N_13858);
and U16723 (N_16723,N_13668,N_12893);
nor U16724 (N_16724,N_13421,N_12861);
or U16725 (N_16725,N_13499,N_13734);
nor U16726 (N_16726,N_14145,N_14959);
nor U16727 (N_16727,N_13214,N_13852);
nand U16728 (N_16728,N_14762,N_12928);
nor U16729 (N_16729,N_13073,N_14915);
or U16730 (N_16730,N_14262,N_13504);
nand U16731 (N_16731,N_14071,N_14783);
and U16732 (N_16732,N_13499,N_13143);
nand U16733 (N_16733,N_13001,N_13695);
and U16734 (N_16734,N_14095,N_13993);
or U16735 (N_16735,N_13346,N_13576);
nand U16736 (N_16736,N_13935,N_13130);
and U16737 (N_16737,N_14554,N_12505);
or U16738 (N_16738,N_13633,N_14322);
nor U16739 (N_16739,N_13408,N_13201);
or U16740 (N_16740,N_13871,N_13992);
and U16741 (N_16741,N_13821,N_14567);
nand U16742 (N_16742,N_13301,N_13314);
and U16743 (N_16743,N_13330,N_13208);
and U16744 (N_16744,N_12668,N_14783);
nand U16745 (N_16745,N_13199,N_13315);
or U16746 (N_16746,N_14215,N_14804);
nor U16747 (N_16747,N_13999,N_14145);
or U16748 (N_16748,N_13423,N_12970);
nor U16749 (N_16749,N_12824,N_12542);
nor U16750 (N_16750,N_12911,N_14728);
nand U16751 (N_16751,N_12815,N_13312);
nor U16752 (N_16752,N_14162,N_14181);
nand U16753 (N_16753,N_13536,N_13176);
nor U16754 (N_16754,N_13427,N_13163);
nor U16755 (N_16755,N_13823,N_14937);
or U16756 (N_16756,N_13396,N_12550);
nor U16757 (N_16757,N_14007,N_13807);
or U16758 (N_16758,N_13491,N_14057);
nor U16759 (N_16759,N_13722,N_13784);
and U16760 (N_16760,N_13315,N_13477);
or U16761 (N_16761,N_13410,N_13817);
and U16762 (N_16762,N_13261,N_12680);
nor U16763 (N_16763,N_13137,N_13110);
nand U16764 (N_16764,N_13990,N_14755);
nor U16765 (N_16765,N_13654,N_12848);
nand U16766 (N_16766,N_13498,N_12685);
nand U16767 (N_16767,N_13313,N_12569);
or U16768 (N_16768,N_14142,N_13244);
nand U16769 (N_16769,N_13940,N_14799);
nor U16770 (N_16770,N_14820,N_13520);
or U16771 (N_16771,N_13768,N_12584);
nand U16772 (N_16772,N_13324,N_14421);
nor U16773 (N_16773,N_14141,N_14438);
nand U16774 (N_16774,N_13840,N_12928);
and U16775 (N_16775,N_13087,N_14651);
nand U16776 (N_16776,N_12887,N_14097);
and U16777 (N_16777,N_14806,N_13110);
and U16778 (N_16778,N_12740,N_14408);
xnor U16779 (N_16779,N_13665,N_13878);
and U16780 (N_16780,N_13784,N_14238);
or U16781 (N_16781,N_14738,N_14443);
or U16782 (N_16782,N_12791,N_13036);
or U16783 (N_16783,N_14536,N_14025);
and U16784 (N_16784,N_14178,N_14540);
or U16785 (N_16785,N_13868,N_14025);
nand U16786 (N_16786,N_13948,N_13123);
nor U16787 (N_16787,N_13225,N_12815);
or U16788 (N_16788,N_12765,N_12976);
nor U16789 (N_16789,N_13928,N_12989);
or U16790 (N_16790,N_14484,N_13871);
or U16791 (N_16791,N_13146,N_13481);
nor U16792 (N_16792,N_13245,N_12931);
nor U16793 (N_16793,N_13496,N_14857);
and U16794 (N_16794,N_12604,N_13174);
nand U16795 (N_16795,N_14112,N_13161);
nand U16796 (N_16796,N_13238,N_12552);
or U16797 (N_16797,N_13983,N_13048);
nor U16798 (N_16798,N_14513,N_13189);
and U16799 (N_16799,N_13346,N_12676);
nor U16800 (N_16800,N_13166,N_12525);
nor U16801 (N_16801,N_14273,N_13970);
and U16802 (N_16802,N_14937,N_14120);
or U16803 (N_16803,N_14688,N_14737);
nand U16804 (N_16804,N_13362,N_12805);
or U16805 (N_16805,N_14163,N_14585);
nand U16806 (N_16806,N_12530,N_12824);
nor U16807 (N_16807,N_12921,N_13121);
nor U16808 (N_16808,N_14361,N_14020);
nor U16809 (N_16809,N_14747,N_13845);
and U16810 (N_16810,N_14342,N_14031);
nor U16811 (N_16811,N_14855,N_12673);
or U16812 (N_16812,N_13097,N_14923);
xnor U16813 (N_16813,N_14932,N_14252);
nor U16814 (N_16814,N_13071,N_13036);
nand U16815 (N_16815,N_14327,N_14028);
nor U16816 (N_16816,N_12776,N_13090);
xor U16817 (N_16817,N_13116,N_13312);
and U16818 (N_16818,N_12571,N_14899);
and U16819 (N_16819,N_14776,N_13094);
or U16820 (N_16820,N_13101,N_12684);
nand U16821 (N_16821,N_14642,N_14216);
or U16822 (N_16822,N_13591,N_13109);
or U16823 (N_16823,N_12840,N_14779);
xnor U16824 (N_16824,N_13041,N_13124);
nor U16825 (N_16825,N_14312,N_13825);
or U16826 (N_16826,N_13906,N_14596);
nand U16827 (N_16827,N_14887,N_14111);
or U16828 (N_16828,N_14071,N_14243);
and U16829 (N_16829,N_13927,N_14227);
nand U16830 (N_16830,N_14341,N_14547);
nand U16831 (N_16831,N_13042,N_12943);
nor U16832 (N_16832,N_12967,N_12655);
nor U16833 (N_16833,N_13167,N_14598);
and U16834 (N_16834,N_12793,N_14222);
and U16835 (N_16835,N_13452,N_14842);
and U16836 (N_16836,N_13371,N_12585);
nor U16837 (N_16837,N_13213,N_12964);
nor U16838 (N_16838,N_14343,N_13728);
and U16839 (N_16839,N_14658,N_13421);
and U16840 (N_16840,N_14174,N_14398);
and U16841 (N_16841,N_12529,N_13999);
and U16842 (N_16842,N_13349,N_12951);
and U16843 (N_16843,N_13484,N_12816);
or U16844 (N_16844,N_14293,N_14616);
and U16845 (N_16845,N_12561,N_14108);
nor U16846 (N_16846,N_13762,N_12934);
nor U16847 (N_16847,N_12500,N_14728);
and U16848 (N_16848,N_14270,N_13160);
and U16849 (N_16849,N_13190,N_12658);
or U16850 (N_16850,N_13354,N_13390);
nand U16851 (N_16851,N_14502,N_12760);
and U16852 (N_16852,N_12878,N_13776);
or U16853 (N_16853,N_13192,N_14595);
or U16854 (N_16854,N_13317,N_13472);
or U16855 (N_16855,N_14511,N_14291);
nand U16856 (N_16856,N_14966,N_13703);
or U16857 (N_16857,N_12827,N_13810);
and U16858 (N_16858,N_13350,N_13359);
nor U16859 (N_16859,N_12947,N_12991);
and U16860 (N_16860,N_14066,N_14412);
and U16861 (N_16861,N_13017,N_13343);
nor U16862 (N_16862,N_14069,N_13269);
nor U16863 (N_16863,N_14046,N_13864);
nor U16864 (N_16864,N_13439,N_13261);
or U16865 (N_16865,N_13909,N_13818);
nor U16866 (N_16866,N_14365,N_13719);
nand U16867 (N_16867,N_13860,N_12540);
and U16868 (N_16868,N_13958,N_13836);
and U16869 (N_16869,N_13269,N_14437);
or U16870 (N_16870,N_13088,N_14705);
or U16871 (N_16871,N_14093,N_14663);
nand U16872 (N_16872,N_14771,N_13430);
nand U16873 (N_16873,N_12503,N_14380);
nor U16874 (N_16874,N_13018,N_14485);
and U16875 (N_16875,N_13825,N_12905);
or U16876 (N_16876,N_14642,N_14665);
nor U16877 (N_16877,N_14908,N_14222);
nor U16878 (N_16878,N_14277,N_12986);
nor U16879 (N_16879,N_14597,N_13450);
nor U16880 (N_16880,N_13081,N_14818);
and U16881 (N_16881,N_13192,N_13337);
or U16882 (N_16882,N_14709,N_13882);
nand U16883 (N_16883,N_13596,N_14207);
and U16884 (N_16884,N_14779,N_12595);
nor U16885 (N_16885,N_12700,N_13418);
xor U16886 (N_16886,N_14218,N_14736);
or U16887 (N_16887,N_13550,N_14605);
nand U16888 (N_16888,N_14647,N_13369);
nand U16889 (N_16889,N_12503,N_14332);
nor U16890 (N_16890,N_12658,N_14417);
nand U16891 (N_16891,N_13318,N_14492);
and U16892 (N_16892,N_13097,N_12803);
nor U16893 (N_16893,N_14635,N_13717);
nand U16894 (N_16894,N_13876,N_13096);
nand U16895 (N_16895,N_13568,N_13908);
or U16896 (N_16896,N_13606,N_13306);
nor U16897 (N_16897,N_13470,N_14971);
nor U16898 (N_16898,N_12516,N_13807);
nor U16899 (N_16899,N_14446,N_14813);
nand U16900 (N_16900,N_13001,N_13271);
nor U16901 (N_16901,N_14454,N_14889);
or U16902 (N_16902,N_14608,N_12669);
nor U16903 (N_16903,N_12939,N_13293);
nor U16904 (N_16904,N_13674,N_14284);
nand U16905 (N_16905,N_12860,N_14465);
nand U16906 (N_16906,N_14940,N_14010);
nand U16907 (N_16907,N_14117,N_12547);
nand U16908 (N_16908,N_12833,N_14894);
and U16909 (N_16909,N_14821,N_14961);
nor U16910 (N_16910,N_13316,N_13522);
or U16911 (N_16911,N_14062,N_13778);
and U16912 (N_16912,N_13367,N_13890);
nor U16913 (N_16913,N_14564,N_13319);
nand U16914 (N_16914,N_13993,N_14052);
nand U16915 (N_16915,N_13947,N_14710);
or U16916 (N_16916,N_14073,N_14021);
xor U16917 (N_16917,N_13740,N_14990);
nor U16918 (N_16918,N_12702,N_12619);
and U16919 (N_16919,N_13150,N_14233);
nand U16920 (N_16920,N_14509,N_14591);
nor U16921 (N_16921,N_13682,N_13477);
or U16922 (N_16922,N_14683,N_12591);
or U16923 (N_16923,N_14433,N_14049);
nor U16924 (N_16924,N_14736,N_14691);
and U16925 (N_16925,N_12626,N_13061);
nand U16926 (N_16926,N_13092,N_14482);
nor U16927 (N_16927,N_13641,N_14591);
or U16928 (N_16928,N_13216,N_14243);
and U16929 (N_16929,N_12726,N_13851);
nor U16930 (N_16930,N_13553,N_12955);
nand U16931 (N_16931,N_14793,N_13000);
or U16932 (N_16932,N_14995,N_12513);
and U16933 (N_16933,N_13264,N_13470);
nor U16934 (N_16934,N_14884,N_14264);
or U16935 (N_16935,N_13669,N_14997);
nor U16936 (N_16936,N_14108,N_12540);
nand U16937 (N_16937,N_13838,N_12797);
nor U16938 (N_16938,N_13992,N_12879);
nand U16939 (N_16939,N_14159,N_13769);
or U16940 (N_16940,N_12705,N_13252);
or U16941 (N_16941,N_12727,N_14104);
nor U16942 (N_16942,N_12541,N_12661);
nor U16943 (N_16943,N_13385,N_13501);
and U16944 (N_16944,N_13516,N_14229);
or U16945 (N_16945,N_12710,N_13393);
and U16946 (N_16946,N_13871,N_14005);
and U16947 (N_16947,N_14485,N_14439);
or U16948 (N_16948,N_12602,N_13673);
nand U16949 (N_16949,N_13854,N_14336);
nand U16950 (N_16950,N_12660,N_14246);
or U16951 (N_16951,N_12626,N_12838);
and U16952 (N_16952,N_12766,N_14566);
xnor U16953 (N_16953,N_14944,N_13739);
nand U16954 (N_16954,N_14373,N_12784);
nand U16955 (N_16955,N_13127,N_12693);
and U16956 (N_16956,N_14712,N_13470);
or U16957 (N_16957,N_13784,N_13298);
nand U16958 (N_16958,N_13891,N_14669);
nor U16959 (N_16959,N_12908,N_13540);
nand U16960 (N_16960,N_12649,N_13963);
and U16961 (N_16961,N_13496,N_12843);
and U16962 (N_16962,N_14711,N_14168);
or U16963 (N_16963,N_14275,N_13376);
nor U16964 (N_16964,N_12921,N_13149);
nand U16965 (N_16965,N_14554,N_13733);
nor U16966 (N_16966,N_12693,N_13082);
nor U16967 (N_16967,N_13725,N_14106);
and U16968 (N_16968,N_13087,N_14836);
nand U16969 (N_16969,N_14788,N_12890);
nor U16970 (N_16970,N_14336,N_13364);
or U16971 (N_16971,N_12967,N_14484);
nor U16972 (N_16972,N_14500,N_14801);
nand U16973 (N_16973,N_13786,N_14533);
or U16974 (N_16974,N_13714,N_13773);
nor U16975 (N_16975,N_13905,N_12828);
nor U16976 (N_16976,N_14100,N_13198);
nand U16977 (N_16977,N_12892,N_13927);
or U16978 (N_16978,N_13943,N_14417);
nor U16979 (N_16979,N_14719,N_13670);
nor U16980 (N_16980,N_13520,N_12634);
nor U16981 (N_16981,N_13672,N_13633);
nor U16982 (N_16982,N_12831,N_12875);
and U16983 (N_16983,N_13470,N_13219);
nor U16984 (N_16984,N_12592,N_14581);
nand U16985 (N_16985,N_13422,N_12650);
or U16986 (N_16986,N_13369,N_12725);
and U16987 (N_16987,N_12867,N_13761);
and U16988 (N_16988,N_13967,N_13779);
nor U16989 (N_16989,N_13054,N_14330);
and U16990 (N_16990,N_12757,N_13192);
and U16991 (N_16991,N_13977,N_13952);
and U16992 (N_16992,N_13768,N_14670);
xor U16993 (N_16993,N_14220,N_14827);
nor U16994 (N_16994,N_14467,N_14695);
and U16995 (N_16995,N_14119,N_12764);
or U16996 (N_16996,N_13732,N_13498);
and U16997 (N_16997,N_14452,N_13903);
and U16998 (N_16998,N_13230,N_14266);
and U16999 (N_16999,N_14018,N_14661);
or U17000 (N_17000,N_12891,N_13251);
nand U17001 (N_17001,N_14049,N_12601);
and U17002 (N_17002,N_13898,N_13627);
or U17003 (N_17003,N_13988,N_13879);
nor U17004 (N_17004,N_13068,N_14445);
or U17005 (N_17005,N_13817,N_14794);
xor U17006 (N_17006,N_13818,N_13460);
nand U17007 (N_17007,N_12949,N_14096);
nor U17008 (N_17008,N_13644,N_14533);
and U17009 (N_17009,N_13678,N_12561);
nor U17010 (N_17010,N_14541,N_12888);
nor U17011 (N_17011,N_14944,N_13535);
nor U17012 (N_17012,N_14841,N_12625);
nor U17013 (N_17013,N_13510,N_13754);
nand U17014 (N_17014,N_14027,N_13740);
and U17015 (N_17015,N_14867,N_12700);
xnor U17016 (N_17016,N_14032,N_13925);
nand U17017 (N_17017,N_14095,N_13325);
or U17018 (N_17018,N_12612,N_13183);
and U17019 (N_17019,N_14195,N_13248);
nor U17020 (N_17020,N_13841,N_13862);
nand U17021 (N_17021,N_14065,N_13401);
nand U17022 (N_17022,N_13088,N_13992);
and U17023 (N_17023,N_14781,N_14642);
or U17024 (N_17024,N_13137,N_14071);
nor U17025 (N_17025,N_14624,N_12943);
xor U17026 (N_17026,N_14666,N_14223);
or U17027 (N_17027,N_14984,N_14012);
nand U17028 (N_17028,N_14420,N_12880);
nand U17029 (N_17029,N_13169,N_13572);
and U17030 (N_17030,N_13404,N_14544);
and U17031 (N_17031,N_14932,N_13211);
nand U17032 (N_17032,N_14295,N_12944);
nand U17033 (N_17033,N_13521,N_13831);
and U17034 (N_17034,N_13024,N_13057);
or U17035 (N_17035,N_14317,N_14897);
and U17036 (N_17036,N_13935,N_13411);
or U17037 (N_17037,N_13637,N_14781);
nor U17038 (N_17038,N_14029,N_13627);
or U17039 (N_17039,N_12582,N_14390);
nand U17040 (N_17040,N_12885,N_12574);
xnor U17041 (N_17041,N_13518,N_12788);
nand U17042 (N_17042,N_13448,N_13321);
nand U17043 (N_17043,N_12520,N_14790);
nor U17044 (N_17044,N_14227,N_14325);
or U17045 (N_17045,N_13844,N_13538);
and U17046 (N_17046,N_13327,N_14865);
nor U17047 (N_17047,N_13246,N_13468);
or U17048 (N_17048,N_13343,N_13821);
nor U17049 (N_17049,N_12855,N_13219);
and U17050 (N_17050,N_14915,N_14418);
or U17051 (N_17051,N_13217,N_14677);
and U17052 (N_17052,N_13429,N_14186);
and U17053 (N_17053,N_14071,N_14797);
nor U17054 (N_17054,N_14123,N_14967);
and U17055 (N_17055,N_13610,N_14065);
nand U17056 (N_17056,N_13562,N_12671);
xor U17057 (N_17057,N_14838,N_13347);
nor U17058 (N_17058,N_14498,N_14178);
nand U17059 (N_17059,N_12970,N_13119);
nor U17060 (N_17060,N_13369,N_13584);
nor U17061 (N_17061,N_12930,N_13168);
nand U17062 (N_17062,N_14321,N_14830);
and U17063 (N_17063,N_14026,N_12829);
and U17064 (N_17064,N_14324,N_13954);
xor U17065 (N_17065,N_12702,N_14216);
nor U17066 (N_17066,N_12598,N_14687);
nor U17067 (N_17067,N_14886,N_14214);
nand U17068 (N_17068,N_14312,N_13093);
nor U17069 (N_17069,N_13298,N_14198);
nand U17070 (N_17070,N_12689,N_14395);
nand U17071 (N_17071,N_13886,N_12956);
nand U17072 (N_17072,N_13788,N_13648);
nor U17073 (N_17073,N_13280,N_13066);
nand U17074 (N_17074,N_13822,N_14260);
nand U17075 (N_17075,N_14568,N_12726);
nand U17076 (N_17076,N_12912,N_12860);
xor U17077 (N_17077,N_14046,N_13846);
or U17078 (N_17078,N_14343,N_14268);
and U17079 (N_17079,N_14259,N_14650);
nand U17080 (N_17080,N_13153,N_13348);
nand U17081 (N_17081,N_13636,N_14393);
or U17082 (N_17082,N_13378,N_12883);
or U17083 (N_17083,N_13527,N_14567);
nand U17084 (N_17084,N_13991,N_14903);
nand U17085 (N_17085,N_14086,N_12588);
and U17086 (N_17086,N_13844,N_13528);
and U17087 (N_17087,N_14740,N_14702);
or U17088 (N_17088,N_13879,N_14880);
nand U17089 (N_17089,N_14782,N_14555);
nor U17090 (N_17090,N_14571,N_14313);
or U17091 (N_17091,N_14019,N_13648);
or U17092 (N_17092,N_12513,N_14437);
nand U17093 (N_17093,N_14581,N_13958);
and U17094 (N_17094,N_14250,N_14991);
and U17095 (N_17095,N_12736,N_14343);
or U17096 (N_17096,N_14200,N_13692);
or U17097 (N_17097,N_14057,N_12940);
nor U17098 (N_17098,N_13545,N_13645);
or U17099 (N_17099,N_14301,N_13521);
nand U17100 (N_17100,N_13836,N_14659);
nand U17101 (N_17101,N_14951,N_13236);
or U17102 (N_17102,N_12590,N_12678);
nor U17103 (N_17103,N_14987,N_12822);
or U17104 (N_17104,N_14438,N_13018);
nand U17105 (N_17105,N_13071,N_14711);
xnor U17106 (N_17106,N_14752,N_13910);
nand U17107 (N_17107,N_13647,N_13197);
or U17108 (N_17108,N_14884,N_13254);
or U17109 (N_17109,N_13448,N_13033);
nor U17110 (N_17110,N_13732,N_12532);
or U17111 (N_17111,N_12608,N_14201);
and U17112 (N_17112,N_13841,N_12830);
nor U17113 (N_17113,N_12744,N_14325);
and U17114 (N_17114,N_14190,N_14564);
and U17115 (N_17115,N_14637,N_14804);
nand U17116 (N_17116,N_13954,N_13368);
or U17117 (N_17117,N_12986,N_14705);
and U17118 (N_17118,N_13266,N_13463);
nor U17119 (N_17119,N_13908,N_14894);
or U17120 (N_17120,N_14326,N_13471);
nor U17121 (N_17121,N_14975,N_14488);
nor U17122 (N_17122,N_14563,N_14502);
and U17123 (N_17123,N_14383,N_14404);
nor U17124 (N_17124,N_13669,N_13629);
or U17125 (N_17125,N_14232,N_12509);
nor U17126 (N_17126,N_12774,N_14316);
and U17127 (N_17127,N_12913,N_14111);
and U17128 (N_17128,N_12987,N_12771);
nor U17129 (N_17129,N_13434,N_13750);
and U17130 (N_17130,N_14174,N_13789);
nand U17131 (N_17131,N_13106,N_14891);
nor U17132 (N_17132,N_14276,N_14669);
nand U17133 (N_17133,N_12614,N_13360);
nor U17134 (N_17134,N_13913,N_12813);
nor U17135 (N_17135,N_14687,N_14122);
or U17136 (N_17136,N_12963,N_13198);
nor U17137 (N_17137,N_14027,N_13236);
nand U17138 (N_17138,N_13668,N_14789);
nand U17139 (N_17139,N_13603,N_12523);
and U17140 (N_17140,N_12948,N_14106);
nand U17141 (N_17141,N_14844,N_13739);
nor U17142 (N_17142,N_14906,N_13297);
nor U17143 (N_17143,N_13359,N_12633);
or U17144 (N_17144,N_12530,N_13771);
or U17145 (N_17145,N_12644,N_13313);
nor U17146 (N_17146,N_13382,N_13488);
nor U17147 (N_17147,N_12726,N_14897);
and U17148 (N_17148,N_13946,N_13497);
nand U17149 (N_17149,N_14595,N_14328);
nor U17150 (N_17150,N_14383,N_14670);
and U17151 (N_17151,N_12596,N_13179);
and U17152 (N_17152,N_13054,N_14714);
nand U17153 (N_17153,N_14653,N_14264);
nand U17154 (N_17154,N_13307,N_14766);
and U17155 (N_17155,N_12690,N_13848);
nor U17156 (N_17156,N_13622,N_12696);
nand U17157 (N_17157,N_13146,N_13883);
nand U17158 (N_17158,N_12885,N_13967);
nor U17159 (N_17159,N_14823,N_14248);
nand U17160 (N_17160,N_14451,N_14926);
and U17161 (N_17161,N_14589,N_13331);
and U17162 (N_17162,N_12604,N_13934);
or U17163 (N_17163,N_12649,N_12637);
or U17164 (N_17164,N_13744,N_13402);
xnor U17165 (N_17165,N_14836,N_13178);
nor U17166 (N_17166,N_13942,N_12787);
or U17167 (N_17167,N_13175,N_14611);
and U17168 (N_17168,N_12657,N_14684);
nand U17169 (N_17169,N_14352,N_14310);
nand U17170 (N_17170,N_12507,N_13705);
nand U17171 (N_17171,N_14219,N_13011);
and U17172 (N_17172,N_14644,N_13718);
and U17173 (N_17173,N_12855,N_13323);
and U17174 (N_17174,N_14294,N_14640);
nor U17175 (N_17175,N_14912,N_13056);
or U17176 (N_17176,N_14377,N_14052);
nand U17177 (N_17177,N_14663,N_12604);
nand U17178 (N_17178,N_13710,N_14550);
nand U17179 (N_17179,N_14701,N_14633);
nand U17180 (N_17180,N_14299,N_13725);
nor U17181 (N_17181,N_13458,N_12644);
nand U17182 (N_17182,N_14938,N_14464);
or U17183 (N_17183,N_14292,N_12620);
nand U17184 (N_17184,N_13248,N_12598);
nor U17185 (N_17185,N_14642,N_13746);
nor U17186 (N_17186,N_13315,N_12584);
nand U17187 (N_17187,N_12704,N_14757);
and U17188 (N_17188,N_13413,N_12609);
nor U17189 (N_17189,N_14909,N_12640);
nand U17190 (N_17190,N_13780,N_12746);
or U17191 (N_17191,N_14262,N_13050);
nor U17192 (N_17192,N_13909,N_14816);
and U17193 (N_17193,N_13212,N_14987);
nor U17194 (N_17194,N_12775,N_14888);
xnor U17195 (N_17195,N_14135,N_12994);
or U17196 (N_17196,N_12576,N_13233);
and U17197 (N_17197,N_12625,N_14035);
and U17198 (N_17198,N_14493,N_14158);
and U17199 (N_17199,N_14567,N_14262);
or U17200 (N_17200,N_12559,N_13374);
nor U17201 (N_17201,N_14343,N_14143);
nand U17202 (N_17202,N_12900,N_13207);
and U17203 (N_17203,N_14854,N_14030);
and U17204 (N_17204,N_14463,N_12931);
nor U17205 (N_17205,N_12817,N_12726);
xor U17206 (N_17206,N_12710,N_14723);
nand U17207 (N_17207,N_13847,N_14659);
nor U17208 (N_17208,N_12745,N_14439);
nand U17209 (N_17209,N_14911,N_14666);
nand U17210 (N_17210,N_13613,N_14166);
nor U17211 (N_17211,N_14031,N_13755);
nor U17212 (N_17212,N_13025,N_12726);
nand U17213 (N_17213,N_14144,N_12919);
or U17214 (N_17214,N_12910,N_14933);
nand U17215 (N_17215,N_14370,N_14889);
nor U17216 (N_17216,N_13359,N_12982);
nand U17217 (N_17217,N_12661,N_13962);
or U17218 (N_17218,N_12797,N_14350);
xor U17219 (N_17219,N_14356,N_13769);
or U17220 (N_17220,N_13738,N_13037);
nand U17221 (N_17221,N_13969,N_13406);
nand U17222 (N_17222,N_14827,N_13937);
or U17223 (N_17223,N_12969,N_14643);
and U17224 (N_17224,N_13144,N_14895);
or U17225 (N_17225,N_13393,N_14182);
or U17226 (N_17226,N_14539,N_14908);
and U17227 (N_17227,N_14963,N_12661);
nor U17228 (N_17228,N_12998,N_12929);
or U17229 (N_17229,N_14061,N_13265);
nor U17230 (N_17230,N_14690,N_13826);
nor U17231 (N_17231,N_14368,N_14625);
or U17232 (N_17232,N_14027,N_13881);
nor U17233 (N_17233,N_14425,N_13385);
nand U17234 (N_17234,N_13986,N_13561);
and U17235 (N_17235,N_14619,N_12714);
nand U17236 (N_17236,N_13925,N_12766);
nand U17237 (N_17237,N_12583,N_13160);
and U17238 (N_17238,N_14406,N_13600);
or U17239 (N_17239,N_13667,N_13836);
nand U17240 (N_17240,N_13382,N_13363);
nand U17241 (N_17241,N_14528,N_13739);
nand U17242 (N_17242,N_14524,N_14536);
and U17243 (N_17243,N_14515,N_14954);
or U17244 (N_17244,N_14921,N_13466);
nand U17245 (N_17245,N_12822,N_13909);
or U17246 (N_17246,N_14075,N_13605);
and U17247 (N_17247,N_12913,N_14662);
or U17248 (N_17248,N_14631,N_12617);
or U17249 (N_17249,N_13003,N_14056);
or U17250 (N_17250,N_12527,N_12605);
nand U17251 (N_17251,N_13702,N_12574);
or U17252 (N_17252,N_13566,N_13112);
nor U17253 (N_17253,N_14352,N_13542);
nand U17254 (N_17254,N_13552,N_12721);
nor U17255 (N_17255,N_13423,N_14302);
nand U17256 (N_17256,N_14865,N_13522);
nor U17257 (N_17257,N_13049,N_12780);
or U17258 (N_17258,N_13941,N_12924);
or U17259 (N_17259,N_12641,N_13434);
nand U17260 (N_17260,N_12849,N_12591);
nand U17261 (N_17261,N_14869,N_14552);
or U17262 (N_17262,N_13903,N_13564);
nand U17263 (N_17263,N_12796,N_13052);
and U17264 (N_17264,N_13790,N_12776);
and U17265 (N_17265,N_13150,N_13005);
or U17266 (N_17266,N_14422,N_13148);
or U17267 (N_17267,N_14274,N_14727);
nand U17268 (N_17268,N_12578,N_12813);
nand U17269 (N_17269,N_13391,N_14241);
or U17270 (N_17270,N_13442,N_13953);
nand U17271 (N_17271,N_13133,N_14023);
nor U17272 (N_17272,N_12656,N_14564);
nor U17273 (N_17273,N_14950,N_13526);
nand U17274 (N_17274,N_14608,N_12774);
or U17275 (N_17275,N_13822,N_13395);
nor U17276 (N_17276,N_13922,N_13364);
and U17277 (N_17277,N_14915,N_13306);
nor U17278 (N_17278,N_13214,N_13023);
and U17279 (N_17279,N_14291,N_14402);
and U17280 (N_17280,N_14752,N_14024);
nor U17281 (N_17281,N_14621,N_14595);
or U17282 (N_17282,N_13374,N_13916);
nand U17283 (N_17283,N_14768,N_13693);
nor U17284 (N_17284,N_12585,N_12911);
and U17285 (N_17285,N_14878,N_14023);
nor U17286 (N_17286,N_14579,N_14850);
and U17287 (N_17287,N_13038,N_13004);
nor U17288 (N_17288,N_13436,N_14809);
nor U17289 (N_17289,N_14976,N_14619);
and U17290 (N_17290,N_13591,N_13868);
nand U17291 (N_17291,N_14404,N_14960);
or U17292 (N_17292,N_13633,N_12530);
nand U17293 (N_17293,N_13856,N_13155);
nand U17294 (N_17294,N_12865,N_13497);
nand U17295 (N_17295,N_12530,N_13865);
nand U17296 (N_17296,N_14469,N_14478);
or U17297 (N_17297,N_13583,N_13194);
nand U17298 (N_17298,N_13337,N_14968);
nor U17299 (N_17299,N_14596,N_12851);
nor U17300 (N_17300,N_13381,N_14515);
nand U17301 (N_17301,N_12635,N_14463);
or U17302 (N_17302,N_14221,N_13827);
and U17303 (N_17303,N_12904,N_13117);
nand U17304 (N_17304,N_12825,N_14738);
nand U17305 (N_17305,N_12622,N_13512);
nor U17306 (N_17306,N_13675,N_13264);
or U17307 (N_17307,N_14453,N_14984);
and U17308 (N_17308,N_14392,N_14343);
and U17309 (N_17309,N_14115,N_13429);
nand U17310 (N_17310,N_13420,N_13458);
or U17311 (N_17311,N_14497,N_13348);
nand U17312 (N_17312,N_12587,N_14654);
nand U17313 (N_17313,N_13405,N_13822);
or U17314 (N_17314,N_13700,N_13115);
nand U17315 (N_17315,N_13852,N_13181);
or U17316 (N_17316,N_14616,N_13348);
or U17317 (N_17317,N_14977,N_13743);
nor U17318 (N_17318,N_13259,N_12989);
nand U17319 (N_17319,N_12597,N_14344);
and U17320 (N_17320,N_12687,N_14357);
or U17321 (N_17321,N_12662,N_13302);
xnor U17322 (N_17322,N_12623,N_12951);
and U17323 (N_17323,N_12502,N_14355);
nand U17324 (N_17324,N_13509,N_13784);
nand U17325 (N_17325,N_13811,N_13827);
nand U17326 (N_17326,N_14532,N_13662);
nand U17327 (N_17327,N_13837,N_12838);
or U17328 (N_17328,N_13744,N_12580);
and U17329 (N_17329,N_14442,N_14055);
nor U17330 (N_17330,N_13741,N_13135);
and U17331 (N_17331,N_13671,N_14115);
nand U17332 (N_17332,N_13851,N_14281);
or U17333 (N_17333,N_13904,N_14763);
or U17334 (N_17334,N_14204,N_14174);
nand U17335 (N_17335,N_13052,N_12543);
or U17336 (N_17336,N_12562,N_14709);
and U17337 (N_17337,N_13270,N_12613);
nand U17338 (N_17338,N_13425,N_14216);
and U17339 (N_17339,N_14859,N_13651);
and U17340 (N_17340,N_12586,N_14281);
or U17341 (N_17341,N_13717,N_14465);
and U17342 (N_17342,N_13348,N_13628);
nand U17343 (N_17343,N_14695,N_13196);
and U17344 (N_17344,N_12823,N_14948);
nor U17345 (N_17345,N_14124,N_13489);
nor U17346 (N_17346,N_13313,N_14192);
or U17347 (N_17347,N_13717,N_14042);
and U17348 (N_17348,N_13977,N_13483);
or U17349 (N_17349,N_13756,N_13781);
nand U17350 (N_17350,N_14866,N_13078);
nand U17351 (N_17351,N_14987,N_14672);
nor U17352 (N_17352,N_14552,N_12956);
nand U17353 (N_17353,N_13677,N_14541);
and U17354 (N_17354,N_13811,N_14639);
and U17355 (N_17355,N_14721,N_12795);
nand U17356 (N_17356,N_14690,N_12947);
nor U17357 (N_17357,N_12945,N_13030);
and U17358 (N_17358,N_14400,N_14029);
nand U17359 (N_17359,N_13437,N_13025);
nor U17360 (N_17360,N_14425,N_14683);
or U17361 (N_17361,N_14640,N_14001);
nor U17362 (N_17362,N_13947,N_14750);
and U17363 (N_17363,N_14433,N_13320);
xnor U17364 (N_17364,N_14217,N_13537);
nand U17365 (N_17365,N_13913,N_14669);
nor U17366 (N_17366,N_13243,N_12935);
and U17367 (N_17367,N_13368,N_13746);
nand U17368 (N_17368,N_14741,N_13961);
nor U17369 (N_17369,N_13692,N_12887);
or U17370 (N_17370,N_14161,N_14365);
or U17371 (N_17371,N_14367,N_13414);
and U17372 (N_17372,N_14929,N_13293);
nand U17373 (N_17373,N_12891,N_12527);
or U17374 (N_17374,N_13421,N_14489);
nand U17375 (N_17375,N_12875,N_14716);
nor U17376 (N_17376,N_12781,N_12520);
nand U17377 (N_17377,N_12662,N_14480);
or U17378 (N_17378,N_14721,N_13944);
and U17379 (N_17379,N_14890,N_13569);
and U17380 (N_17380,N_14547,N_12995);
or U17381 (N_17381,N_13849,N_14448);
or U17382 (N_17382,N_12645,N_14445);
or U17383 (N_17383,N_13512,N_14267);
nand U17384 (N_17384,N_12697,N_14279);
and U17385 (N_17385,N_13933,N_14132);
or U17386 (N_17386,N_13792,N_12861);
and U17387 (N_17387,N_12653,N_14123);
or U17388 (N_17388,N_13454,N_12734);
and U17389 (N_17389,N_12987,N_13734);
xnor U17390 (N_17390,N_14667,N_14804);
and U17391 (N_17391,N_14197,N_14813);
or U17392 (N_17392,N_12598,N_14789);
nand U17393 (N_17393,N_13596,N_14098);
nand U17394 (N_17394,N_12525,N_13792);
xnor U17395 (N_17395,N_12637,N_14623);
nand U17396 (N_17396,N_13462,N_14949);
xor U17397 (N_17397,N_14245,N_13487);
and U17398 (N_17398,N_14634,N_13684);
or U17399 (N_17399,N_12796,N_14876);
nand U17400 (N_17400,N_14771,N_14502);
and U17401 (N_17401,N_13287,N_13679);
nor U17402 (N_17402,N_13677,N_14287);
and U17403 (N_17403,N_13779,N_14014);
xnor U17404 (N_17404,N_13110,N_14013);
or U17405 (N_17405,N_13215,N_13742);
nand U17406 (N_17406,N_13076,N_14435);
nand U17407 (N_17407,N_13138,N_14887);
nand U17408 (N_17408,N_14192,N_13243);
or U17409 (N_17409,N_14768,N_12539);
and U17410 (N_17410,N_13341,N_13817);
nand U17411 (N_17411,N_13365,N_13110);
and U17412 (N_17412,N_13173,N_12530);
nor U17413 (N_17413,N_12842,N_12865);
nor U17414 (N_17414,N_14110,N_13927);
nor U17415 (N_17415,N_14436,N_14906);
nand U17416 (N_17416,N_12607,N_12636);
nor U17417 (N_17417,N_13791,N_13464);
or U17418 (N_17418,N_13160,N_13583);
nand U17419 (N_17419,N_14378,N_14870);
nor U17420 (N_17420,N_14423,N_14613);
nand U17421 (N_17421,N_14876,N_13047);
or U17422 (N_17422,N_13116,N_14694);
and U17423 (N_17423,N_13432,N_12867);
nand U17424 (N_17424,N_13048,N_13392);
or U17425 (N_17425,N_13220,N_13340);
or U17426 (N_17426,N_14106,N_13870);
nand U17427 (N_17427,N_13168,N_12599);
and U17428 (N_17428,N_12724,N_14424);
and U17429 (N_17429,N_13635,N_13175);
nand U17430 (N_17430,N_13685,N_14180);
xor U17431 (N_17431,N_13781,N_13583);
nor U17432 (N_17432,N_12868,N_13260);
or U17433 (N_17433,N_12570,N_13605);
or U17434 (N_17434,N_14848,N_14258);
and U17435 (N_17435,N_14333,N_13982);
nand U17436 (N_17436,N_13128,N_12604);
nand U17437 (N_17437,N_14753,N_14522);
or U17438 (N_17438,N_14398,N_14964);
xor U17439 (N_17439,N_13425,N_14007);
nor U17440 (N_17440,N_14434,N_14358);
nor U17441 (N_17441,N_14719,N_12927);
or U17442 (N_17442,N_13054,N_14411);
nor U17443 (N_17443,N_13379,N_13078);
or U17444 (N_17444,N_13631,N_13886);
and U17445 (N_17445,N_14506,N_14469);
nor U17446 (N_17446,N_13434,N_14425);
nand U17447 (N_17447,N_12973,N_14096);
and U17448 (N_17448,N_14341,N_12703);
or U17449 (N_17449,N_13041,N_13714);
nor U17450 (N_17450,N_14914,N_14919);
or U17451 (N_17451,N_12725,N_14885);
xor U17452 (N_17452,N_14936,N_14786);
nor U17453 (N_17453,N_12844,N_14714);
and U17454 (N_17454,N_14968,N_13381);
or U17455 (N_17455,N_14823,N_12889);
and U17456 (N_17456,N_13583,N_13758);
and U17457 (N_17457,N_14626,N_14873);
xnor U17458 (N_17458,N_13148,N_12990);
nor U17459 (N_17459,N_13974,N_13581);
or U17460 (N_17460,N_13418,N_12703);
and U17461 (N_17461,N_13178,N_14395);
or U17462 (N_17462,N_14498,N_12897);
nor U17463 (N_17463,N_13603,N_13543);
and U17464 (N_17464,N_13449,N_13181);
nor U17465 (N_17465,N_14002,N_13616);
or U17466 (N_17466,N_13176,N_12651);
nand U17467 (N_17467,N_14501,N_14459);
and U17468 (N_17468,N_12507,N_14552);
nor U17469 (N_17469,N_13985,N_14676);
nand U17470 (N_17470,N_13845,N_12723);
nand U17471 (N_17471,N_12921,N_13391);
or U17472 (N_17472,N_14257,N_14054);
or U17473 (N_17473,N_13047,N_13440);
nor U17474 (N_17474,N_13723,N_14529);
and U17475 (N_17475,N_14955,N_12708);
and U17476 (N_17476,N_14912,N_12646);
or U17477 (N_17477,N_14949,N_14751);
and U17478 (N_17478,N_13483,N_12994);
nor U17479 (N_17479,N_13379,N_13625);
nor U17480 (N_17480,N_14267,N_13375);
and U17481 (N_17481,N_14005,N_13417);
and U17482 (N_17482,N_14646,N_12612);
and U17483 (N_17483,N_14400,N_14678);
and U17484 (N_17484,N_14213,N_14568);
and U17485 (N_17485,N_13572,N_12741);
nand U17486 (N_17486,N_13758,N_13370);
nor U17487 (N_17487,N_12737,N_14888);
nor U17488 (N_17488,N_13771,N_14255);
or U17489 (N_17489,N_12819,N_14233);
or U17490 (N_17490,N_13092,N_14607);
nor U17491 (N_17491,N_13018,N_13828);
and U17492 (N_17492,N_14700,N_13352);
nand U17493 (N_17493,N_14581,N_13604);
nand U17494 (N_17494,N_14332,N_12546);
nand U17495 (N_17495,N_13326,N_14671);
or U17496 (N_17496,N_13155,N_12746);
or U17497 (N_17497,N_13702,N_14952);
nor U17498 (N_17498,N_13024,N_14178);
nor U17499 (N_17499,N_12680,N_14282);
or U17500 (N_17500,N_16428,N_15372);
nand U17501 (N_17501,N_16022,N_16312);
nor U17502 (N_17502,N_16043,N_16137);
or U17503 (N_17503,N_15167,N_16513);
or U17504 (N_17504,N_15219,N_15998);
nand U17505 (N_17505,N_17329,N_17025);
or U17506 (N_17506,N_16936,N_17413);
and U17507 (N_17507,N_15645,N_16891);
and U17508 (N_17508,N_15032,N_17009);
nand U17509 (N_17509,N_16817,N_17201);
nand U17510 (N_17510,N_16648,N_15412);
nand U17511 (N_17511,N_15734,N_17082);
nand U17512 (N_17512,N_16553,N_16248);
nor U17513 (N_17513,N_15449,N_16342);
and U17514 (N_17514,N_15124,N_15797);
nor U17515 (N_17515,N_16722,N_15564);
nand U17516 (N_17516,N_15519,N_16162);
and U17517 (N_17517,N_15098,N_15406);
xnor U17518 (N_17518,N_16194,N_17204);
nand U17519 (N_17519,N_16116,N_15060);
nand U17520 (N_17520,N_15244,N_15191);
nand U17521 (N_17521,N_15989,N_16354);
and U17522 (N_17522,N_16167,N_16495);
nand U17523 (N_17523,N_16296,N_17491);
and U17524 (N_17524,N_17095,N_16088);
and U17525 (N_17525,N_15194,N_16982);
nand U17526 (N_17526,N_16766,N_17272);
nor U17527 (N_17527,N_15254,N_15284);
nand U17528 (N_17528,N_17419,N_16590);
nor U17529 (N_17529,N_16527,N_16620);
xnor U17530 (N_17530,N_16662,N_17096);
nand U17531 (N_17531,N_16244,N_16986);
nor U17532 (N_17532,N_15788,N_15905);
nor U17533 (N_17533,N_17490,N_17286);
nand U17534 (N_17534,N_16881,N_16710);
nor U17535 (N_17535,N_17344,N_15500);
nor U17536 (N_17536,N_16206,N_15497);
xnor U17537 (N_17537,N_16123,N_15435);
or U17538 (N_17538,N_15728,N_15415);
nand U17539 (N_17539,N_15223,N_15149);
or U17540 (N_17540,N_15562,N_16509);
nand U17541 (N_17541,N_15466,N_17478);
and U17542 (N_17542,N_16602,N_15988);
or U17543 (N_17543,N_16843,N_16253);
nand U17544 (N_17544,N_15601,N_16687);
nand U17545 (N_17545,N_15690,N_17388);
nand U17546 (N_17546,N_17323,N_15793);
nand U17547 (N_17547,N_15557,N_16411);
nand U17548 (N_17548,N_16181,N_15874);
and U17549 (N_17549,N_15987,N_16155);
and U17550 (N_17550,N_16456,N_16347);
nand U17551 (N_17551,N_16337,N_16521);
nor U17552 (N_17552,N_16684,N_15606);
nand U17553 (N_17553,N_15746,N_17476);
and U17554 (N_17554,N_16115,N_15968);
or U17555 (N_17555,N_15518,N_15560);
xor U17556 (N_17556,N_15943,N_16295);
or U17557 (N_17557,N_16236,N_17430);
or U17558 (N_17558,N_16039,N_15232);
nand U17559 (N_17559,N_16593,N_16076);
nor U17560 (N_17560,N_15817,N_16873);
nand U17561 (N_17561,N_17168,N_17482);
nor U17562 (N_17562,N_16254,N_16726);
and U17563 (N_17563,N_15014,N_16694);
or U17564 (N_17564,N_15163,N_16566);
or U17565 (N_17565,N_17342,N_17186);
or U17566 (N_17566,N_17348,N_16671);
nand U17567 (N_17567,N_15040,N_15470);
and U17568 (N_17568,N_16497,N_16727);
nand U17569 (N_17569,N_16075,N_15525);
nor U17570 (N_17570,N_16277,N_15400);
nor U17571 (N_17571,N_15608,N_15352);
or U17572 (N_17572,N_16500,N_15786);
nand U17573 (N_17573,N_17078,N_15311);
nand U17574 (N_17574,N_15192,N_15565);
xnor U17575 (N_17575,N_15727,N_16153);
or U17576 (N_17576,N_17341,N_15450);
and U17577 (N_17577,N_17159,N_15778);
and U17578 (N_17578,N_16146,N_16420);
and U17579 (N_17579,N_16318,N_16361);
or U17580 (N_17580,N_17406,N_16056);
or U17581 (N_17581,N_17002,N_17194);
xor U17582 (N_17582,N_16796,N_16358);
or U17583 (N_17583,N_15657,N_16603);
and U17584 (N_17584,N_17031,N_15722);
nand U17585 (N_17585,N_15805,N_15973);
nand U17586 (N_17586,N_16205,N_16511);
nand U17587 (N_17587,N_16382,N_16239);
or U17588 (N_17588,N_16217,N_16528);
and U17589 (N_17589,N_17079,N_15618);
and U17590 (N_17590,N_17326,N_16831);
nand U17591 (N_17591,N_16884,N_15609);
nand U17592 (N_17592,N_17143,N_16346);
or U17593 (N_17593,N_16202,N_16467);
and U17594 (N_17594,N_15404,N_15629);
nor U17595 (N_17595,N_15656,N_15212);
and U17596 (N_17596,N_16326,N_15849);
nor U17597 (N_17597,N_16630,N_15659);
nor U17598 (N_17598,N_16689,N_15411);
and U17599 (N_17599,N_16588,N_17203);
and U17600 (N_17600,N_15646,N_17209);
xnor U17601 (N_17601,N_15469,N_15160);
and U17602 (N_17602,N_15062,N_17433);
nor U17603 (N_17603,N_16042,N_17006);
and U17604 (N_17604,N_15769,N_15001);
or U17605 (N_17605,N_16506,N_16679);
nand U17606 (N_17606,N_15049,N_17237);
nor U17607 (N_17607,N_17360,N_17205);
or U17608 (N_17608,N_15902,N_15140);
and U17609 (N_17609,N_15329,N_15332);
and U17610 (N_17610,N_17218,N_15842);
nand U17611 (N_17611,N_15426,N_16968);
and U17612 (N_17612,N_15750,N_16307);
and U17613 (N_17613,N_16867,N_17431);
or U17614 (N_17614,N_15282,N_15022);
nand U17615 (N_17615,N_16803,N_16138);
or U17616 (N_17616,N_15463,N_16265);
nand U17617 (N_17617,N_17142,N_15260);
and U17618 (N_17618,N_16947,N_16915);
or U17619 (N_17619,N_16486,N_15846);
nand U17620 (N_17620,N_17139,N_17175);
nand U17621 (N_17621,N_15290,N_16900);
and U17622 (N_17622,N_15365,N_16663);
and U17623 (N_17623,N_16844,N_17119);
or U17624 (N_17624,N_17451,N_16864);
nand U17625 (N_17625,N_15237,N_15950);
nand U17626 (N_17626,N_15908,N_17115);
nand U17627 (N_17627,N_17032,N_17065);
nor U17628 (N_17628,N_15483,N_15939);
and U17629 (N_17629,N_16201,N_16921);
xor U17630 (N_17630,N_17381,N_15165);
nand U17631 (N_17631,N_17040,N_16066);
or U17632 (N_17632,N_16267,N_15766);
nand U17633 (N_17633,N_16281,N_16322);
or U17634 (N_17634,N_16678,N_17362);
nor U17635 (N_17635,N_15579,N_15255);
or U17636 (N_17636,N_15401,N_17088);
and U17637 (N_17637,N_15993,N_15002);
or U17638 (N_17638,N_17280,N_17050);
nor U17639 (N_17639,N_16243,N_15681);
and U17640 (N_17640,N_17303,N_15221);
and U17641 (N_17641,N_15640,N_17108);
nor U17642 (N_17642,N_16414,N_16938);
nand U17643 (N_17643,N_17255,N_16857);
nor U17644 (N_17644,N_15906,N_16112);
nand U17645 (N_17645,N_16909,N_15082);
nor U17646 (N_17646,N_17244,N_15023);
or U17647 (N_17647,N_17181,N_16447);
and U17648 (N_17648,N_15847,N_15468);
or U17649 (N_17649,N_15200,N_16136);
and U17650 (N_17650,N_16345,N_16397);
nand U17651 (N_17651,N_16987,N_17214);
nand U17652 (N_17652,N_15665,N_16715);
nand U17653 (N_17653,N_15712,N_15678);
or U17654 (N_17654,N_16842,N_16174);
and U17655 (N_17655,N_16736,N_15442);
and U17656 (N_17656,N_15118,N_15588);
and U17657 (N_17657,N_15156,N_15374);
nor U17658 (N_17658,N_17407,N_15972);
nor U17659 (N_17659,N_15956,N_15831);
nand U17660 (N_17660,N_15181,N_17212);
or U17661 (N_17661,N_16238,N_16379);
or U17662 (N_17662,N_16335,N_16618);
and U17663 (N_17663,N_15835,N_16578);
nand U17664 (N_17664,N_15087,N_15702);
or U17665 (N_17665,N_16047,N_16608);
nor U17666 (N_17666,N_17120,N_16157);
or U17667 (N_17667,N_16216,N_15170);
and U17668 (N_17668,N_16330,N_16517);
and U17669 (N_17669,N_16799,N_15132);
nand U17670 (N_17670,N_15248,N_16187);
nor U17671 (N_17671,N_15355,N_17133);
and U17672 (N_17672,N_16926,N_16370);
nand U17673 (N_17673,N_16376,N_16712);
xor U17674 (N_17674,N_17441,N_15603);
nor U17675 (N_17675,N_15113,N_16872);
nand U17676 (N_17676,N_16407,N_15440);
nand U17677 (N_17677,N_16222,N_16709);
and U17678 (N_17678,N_15209,N_17158);
and U17679 (N_17679,N_17350,N_15028);
or U17680 (N_17680,N_15279,N_16573);
nor U17681 (N_17681,N_16655,N_16700);
nand U17682 (N_17682,N_15190,N_16950);
nand U17683 (N_17683,N_15335,N_16021);
and U17684 (N_17684,N_15157,N_15272);
xnor U17685 (N_17685,N_15923,N_16328);
or U17686 (N_17686,N_16834,N_17122);
nand U17687 (N_17687,N_16797,N_16443);
nand U17688 (N_17688,N_17409,N_15630);
nand U17689 (N_17689,N_15760,N_16139);
or U17690 (N_17690,N_16875,N_17202);
and U17691 (N_17691,N_15050,N_16654);
and U17692 (N_17692,N_16085,N_16096);
and U17693 (N_17693,N_16634,N_15651);
xnor U17694 (N_17694,N_17378,N_15333);
or U17695 (N_17695,N_15097,N_16256);
xor U17696 (N_17696,N_16004,N_17048);
or U17697 (N_17697,N_15294,N_15416);
nand U17698 (N_17698,N_17243,N_15578);
or U17699 (N_17699,N_17379,N_17488);
nor U17700 (N_17700,N_16778,N_16895);
and U17701 (N_17701,N_15739,N_16786);
and U17702 (N_17702,N_17034,N_17416);
and U17703 (N_17703,N_15992,N_16327);
nand U17704 (N_17704,N_15408,N_16898);
nand U17705 (N_17705,N_15674,N_16240);
nor U17706 (N_17706,N_16462,N_15017);
nor U17707 (N_17707,N_17465,N_15176);
nor U17708 (N_17708,N_17373,N_16317);
or U17709 (N_17709,N_15146,N_15822);
nor U17710 (N_17710,N_16739,N_15096);
nand U17711 (N_17711,N_16020,N_16331);
and U17712 (N_17712,N_17483,N_17367);
nand U17713 (N_17713,N_16910,N_15800);
nand U17714 (N_17714,N_16209,N_15452);
nor U17715 (N_17715,N_17462,N_16579);
or U17716 (N_17716,N_16760,N_17318);
nor U17717 (N_17717,N_15566,N_15222);
nor U17718 (N_17718,N_16083,N_15868);
or U17719 (N_17719,N_16089,N_17180);
and U17720 (N_17720,N_15692,N_16705);
nand U17721 (N_17721,N_17368,N_17298);
and U17722 (N_17722,N_16830,N_16059);
and U17723 (N_17723,N_16409,N_17366);
and U17724 (N_17724,N_15614,N_16348);
or U17725 (N_17725,N_15036,N_15257);
or U17726 (N_17726,N_15444,N_17163);
nor U17727 (N_17727,N_15013,N_17364);
or U17728 (N_17728,N_16051,N_15732);
nor U17729 (N_17729,N_15738,N_16286);
nor U17730 (N_17730,N_16393,N_15899);
xor U17731 (N_17731,N_15391,N_16384);
nand U17732 (N_17732,N_16568,N_15215);
nor U17733 (N_17733,N_17439,N_16816);
and U17734 (N_17734,N_15448,N_16621);
xor U17735 (N_17735,N_16970,N_15104);
xor U17736 (N_17736,N_16653,N_15536);
nor U17737 (N_17737,N_15065,N_16901);
and U17738 (N_17738,N_15632,N_17325);
nand U17739 (N_17739,N_15628,N_17189);
and U17740 (N_17740,N_16058,N_15175);
nand U17741 (N_17741,N_15396,N_16604);
nor U17742 (N_17742,N_15617,N_16747);
and U17743 (N_17743,N_15867,N_15513);
nand U17744 (N_17744,N_16308,N_15701);
or U17745 (N_17745,N_15460,N_16313);
or U17746 (N_17746,N_15366,N_16696);
nand U17747 (N_17747,N_15121,N_15976);
nor U17748 (N_17748,N_15383,N_15649);
nand U17749 (N_17749,N_15012,N_15595);
nand U17750 (N_17750,N_16888,N_15371);
nand U17751 (N_17751,N_15823,N_17258);
nand U17752 (N_17752,N_16349,N_17140);
nor U17753 (N_17753,N_15356,N_15409);
nand U17754 (N_17754,N_16589,N_16790);
and U17755 (N_17755,N_15653,N_17336);
nand U17756 (N_17756,N_16931,N_15101);
nor U17757 (N_17757,N_16541,N_15583);
and U17758 (N_17758,N_17238,N_15921);
and U17759 (N_17759,N_16363,N_15795);
nor U17760 (N_17760,N_15887,N_16249);
and U17761 (N_17761,N_15672,N_15109);
nand U17762 (N_17762,N_16865,N_15494);
nand U17763 (N_17763,N_17444,N_15507);
nor U17764 (N_17764,N_17259,N_16078);
nor U17765 (N_17765,N_15323,N_16109);
and U17766 (N_17766,N_17291,N_15938);
and U17767 (N_17767,N_15669,N_17386);
nor U17768 (N_17768,N_16724,N_15385);
or U17769 (N_17769,N_16673,N_17059);
nand U17770 (N_17770,N_17160,N_17343);
nand U17771 (N_17771,N_15892,N_17436);
or U17772 (N_17772,N_15775,N_15141);
nor U17773 (N_17773,N_15281,N_15227);
nor U17774 (N_17774,N_15825,N_17077);
or U17775 (N_17775,N_17447,N_16757);
nand U17776 (N_17776,N_15568,N_17374);
or U17777 (N_17777,N_15458,N_15686);
or U17778 (N_17778,N_17497,N_16341);
nand U17779 (N_17779,N_15115,N_17415);
nand U17780 (N_17780,N_16839,N_15089);
and U17781 (N_17781,N_16788,N_15986);
nand U17782 (N_17782,N_17464,N_15407);
or U17783 (N_17783,N_16007,N_16173);
or U17784 (N_17784,N_16917,N_16259);
or U17785 (N_17785,N_17297,N_15326);
and U17786 (N_17786,N_15172,N_16026);
nand U17787 (N_17787,N_15749,N_15554);
or U17788 (N_17788,N_16431,N_15671);
nor U17789 (N_17789,N_17155,N_15839);
nand U17790 (N_17790,N_16214,N_16751);
and U17791 (N_17791,N_16320,N_16964);
and U17792 (N_17792,N_15779,N_17279);
nand U17793 (N_17793,N_17049,N_17100);
nand U17794 (N_17794,N_16114,N_17277);
nor U17795 (N_17795,N_17260,N_15107);
or U17796 (N_17796,N_16071,N_17232);
nor U17797 (N_17797,N_16973,N_15962);
or U17798 (N_17798,N_16158,N_15488);
or U17799 (N_17799,N_16323,N_16924);
or U17800 (N_17800,N_17480,N_15187);
and U17801 (N_17801,N_16596,N_15855);
nor U17802 (N_17802,N_17003,N_15298);
and U17803 (N_17803,N_16961,N_16565);
or U17804 (N_17804,N_16121,N_17382);
or U17805 (N_17805,N_16591,N_17324);
nor U17806 (N_17806,N_15804,N_15826);
nand U17807 (N_17807,N_16377,N_17460);
xnor U17808 (N_17808,N_16721,N_16957);
and U17809 (N_17809,N_16092,N_15946);
and U17810 (N_17810,N_17396,N_15592);
or U17811 (N_17811,N_17250,N_16027);
nor U17812 (N_17812,N_17405,N_15954);
and U17813 (N_17813,N_16802,N_16967);
and U17814 (N_17814,N_15370,N_15465);
nand U17815 (N_17815,N_15801,N_16882);
nand U17816 (N_17816,N_16860,N_16728);
nor U17817 (N_17817,N_17421,N_15388);
nor U17818 (N_17818,N_17047,N_16470);
nor U17819 (N_17819,N_17098,N_16368);
and U17820 (N_17820,N_16478,N_16850);
nand U17821 (N_17821,N_16189,N_15252);
or U17822 (N_17822,N_16496,N_15034);
or U17823 (N_17823,N_15068,N_15381);
nand U17824 (N_17824,N_16661,N_15664);
nand U17825 (N_17825,N_17223,N_17173);
nor U17826 (N_17826,N_15710,N_15964);
nand U17827 (N_17827,N_16062,N_17372);
or U17828 (N_17828,N_17191,N_15848);
and U17829 (N_17829,N_16516,N_16398);
and U17830 (N_17830,N_15824,N_17335);
or U17831 (N_17831,N_15359,N_17440);
and U17832 (N_17832,N_15947,N_15083);
nor U17833 (N_17833,N_16301,N_15079);
or U17834 (N_17834,N_16876,N_16934);
and U17835 (N_17835,N_17333,N_15957);
or U17836 (N_17836,N_17162,N_17370);
xnor U17837 (N_17837,N_17294,N_15944);
nor U17838 (N_17838,N_15410,N_16252);
nand U17839 (N_17839,N_17487,N_16434);
or U17840 (N_17840,N_16396,N_17033);
nor U17841 (N_17841,N_16373,N_15879);
nand U17842 (N_17842,N_17179,N_16809);
and U17843 (N_17843,N_15907,N_16057);
nor U17844 (N_17844,N_16896,N_17193);
xnor U17845 (N_17845,N_16862,N_15870);
and U17846 (N_17846,N_15517,N_15492);
and U17847 (N_17847,N_16392,N_16220);
or U17848 (N_17848,N_16810,N_15431);
nand U17849 (N_17849,N_17365,N_16299);
or U17850 (N_17850,N_16635,N_15607);
and U17851 (N_17851,N_15178,N_17042);
nand U17852 (N_17852,N_15884,N_17429);
nand U17853 (N_17853,N_17475,N_15803);
nand U17854 (N_17854,N_16878,N_16182);
nor U17855 (N_17855,N_16235,N_16213);
nand U17856 (N_17856,N_17390,N_15457);
nor U17857 (N_17857,N_16557,N_16036);
nand U17858 (N_17858,N_17334,N_16783);
nand U17859 (N_17859,N_15813,N_15211);
nor U17860 (N_17860,N_16369,N_16180);
or U17861 (N_17861,N_17262,N_16087);
nand U17862 (N_17862,N_15770,N_15394);
xnor U17863 (N_17863,N_15904,N_16432);
and U17864 (N_17864,N_15891,N_15700);
and U17865 (N_17865,N_16276,N_16877);
nand U17866 (N_17866,N_15360,N_15573);
and U17867 (N_17867,N_16730,N_16124);
and U17868 (N_17868,N_16749,N_15477);
or U17869 (N_17869,N_16930,N_16685);
or U17870 (N_17870,N_15985,N_17315);
nor U17871 (N_17871,N_15981,N_15524);
nand U17872 (N_17872,N_17331,N_16807);
nand U17873 (N_17873,N_15496,N_16442);
nor U17874 (N_17874,N_16659,N_16820);
or U17875 (N_17875,N_16737,N_16505);
and U17876 (N_17876,N_15199,N_16919);
and U17877 (N_17877,N_15612,N_15445);
and U17878 (N_17878,N_16995,N_17131);
nand U17879 (N_17879,N_16670,N_16336);
or U17880 (N_17880,N_16381,N_15833);
and U17881 (N_17881,N_17242,N_16801);
nand U17882 (N_17882,N_15304,N_17225);
nor U17883 (N_17883,N_15195,N_17176);
nor U17884 (N_17884,N_16332,N_17014);
xor U17885 (N_17885,N_16417,N_16775);
or U17886 (N_17886,N_15834,N_16789);
or U17887 (N_17887,N_15309,N_16643);
nand U17888 (N_17888,N_16972,N_15696);
xnor U17889 (N_17889,N_15229,N_16503);
or U17890 (N_17890,N_15996,N_15004);
nor U17891 (N_17891,N_15478,N_15241);
or U17892 (N_17892,N_16585,N_16641);
or U17893 (N_17893,N_16567,N_15336);
nor U17894 (N_17894,N_15663,N_15814);
nor U17895 (N_17895,N_15596,N_17211);
nand U17896 (N_17896,N_16823,N_17450);
and U17897 (N_17897,N_15039,N_15295);
nand U17898 (N_17898,N_16292,N_16093);
and U17899 (N_17899,N_16003,N_17437);
and U17900 (N_17900,N_15027,N_16226);
and U17901 (N_17901,N_15090,N_15572);
or U17902 (N_17902,N_16283,N_15752);
nor U17903 (N_17903,N_16683,N_15080);
or U17904 (N_17904,N_17266,N_16615);
and U17905 (N_17905,N_16572,N_15966);
and U17906 (N_17906,N_16072,N_16808);
nand U17907 (N_17907,N_16143,N_16750);
nand U17908 (N_17908,N_16188,N_16971);
nand U17909 (N_17909,N_16508,N_15123);
nor U17910 (N_17910,N_15549,N_17001);
nor U17911 (N_17911,N_17219,N_15179);
nor U17912 (N_17912,N_16646,N_15828);
nand U17913 (N_17913,N_15726,N_16385);
nor U17914 (N_17914,N_15535,N_15895);
nor U17915 (N_17915,N_16371,N_15941);
and U17916 (N_17916,N_17461,N_15306);
and U17917 (N_17917,N_16871,N_15647);
and U17918 (N_17918,N_15911,N_15886);
nor U17919 (N_17919,N_15783,N_17197);
and U17920 (N_17920,N_17005,N_17332);
nand U17921 (N_17921,N_15216,N_17351);
nor U17922 (N_17922,N_17161,N_16492);
or U17923 (N_17923,N_16231,N_16245);
and U17924 (N_17924,N_15048,N_15790);
or U17925 (N_17925,N_16932,N_15740);
nand U17926 (N_17926,N_16441,N_15314);
or U17927 (N_17927,N_17392,N_17038);
and U17928 (N_17928,N_16129,N_17192);
nor U17929 (N_17929,N_16804,N_16151);
nand U17930 (N_17930,N_16049,N_15009);
or U17931 (N_17931,N_17221,N_15283);
or U17932 (N_17932,N_15054,N_15337);
and U17933 (N_17933,N_16120,N_16989);
nand U17934 (N_17934,N_15933,N_16438);
or U17935 (N_17935,N_17253,N_16111);
nor U17936 (N_17936,N_15375,N_17310);
nor U17937 (N_17937,N_16664,N_15755);
and U17938 (N_17938,N_16781,N_15155);
and U17939 (N_17939,N_15158,N_15934);
or U17940 (N_17940,N_17481,N_16592);
or U17941 (N_17941,N_17347,N_15242);
nor U17942 (N_17942,N_15982,N_15338);
or U17943 (N_17943,N_15138,N_15302);
and U17944 (N_17944,N_15648,N_15088);
or U17945 (N_17945,N_15979,N_15210);
nor U17946 (N_17946,N_15094,N_16474);
nor U17947 (N_17947,N_16996,N_16991);
nand U17948 (N_17948,N_15243,N_15520);
and U17949 (N_17949,N_16161,N_17445);
nand U17950 (N_17950,N_15376,N_17263);
xnor U17951 (N_17951,N_16263,N_16014);
or U17952 (N_17952,N_17314,N_15150);
or U17953 (N_17953,N_16183,N_15610);
or U17954 (N_17954,N_15182,N_16433);
xnor U17955 (N_17955,N_16748,N_16069);
or U17956 (N_17956,N_15358,N_16074);
nand U17957 (N_17957,N_16160,N_16403);
or U17958 (N_17958,N_16122,N_17467);
and U17959 (N_17959,N_16911,N_15958);
and U17960 (N_17960,N_15552,N_16128);
or U17961 (N_17961,N_15951,N_15278);
or U17962 (N_17962,N_16605,N_16983);
or U17963 (N_17963,N_16549,N_16001);
nor U17964 (N_17964,N_16282,N_15816);
and U17965 (N_17965,N_17000,N_15430);
and U17966 (N_17966,N_17313,N_15164);
nor U17967 (N_17967,N_17486,N_16445);
nor U17968 (N_17968,N_17355,N_15503);
nor U17969 (N_17969,N_16879,N_15684);
nor U17970 (N_17970,N_16487,N_16009);
nor U17971 (N_17971,N_15819,N_17199);
and U17972 (N_17972,N_15214,N_16774);
and U17973 (N_17973,N_15844,N_17187);
and U17974 (N_17974,N_15875,N_16853);
or U17975 (N_17975,N_16483,N_15591);
nor U17976 (N_17976,N_17021,N_15078);
or U17977 (N_17977,N_16204,N_16636);
or U17978 (N_17978,N_15840,N_17171);
nand U17979 (N_17979,N_15655,N_16031);
and U17980 (N_17980,N_15092,N_15186);
and U17981 (N_17981,N_16387,N_16692);
nand U17982 (N_17982,N_16838,N_16024);
nor U17983 (N_17983,N_17485,N_15574);
nand U17984 (N_17984,N_15263,N_16227);
nand U17985 (N_17985,N_16310,N_15873);
and U17986 (N_17986,N_15654,N_16787);
and U17987 (N_17987,N_15251,N_17083);
and U17988 (N_17988,N_16928,N_15707);
nor U17989 (N_17989,N_17185,N_15961);
and U17990 (N_17990,N_16548,N_15787);
and U17991 (N_17991,N_16916,N_16570);
or U17992 (N_17992,N_16477,N_16581);
nand U17993 (N_17993,N_17274,N_16571);
nor U17994 (N_17994,N_15791,N_16311);
nor U17995 (N_17995,N_17398,N_17322);
nor U17996 (N_17996,N_16945,N_15220);
nor U17997 (N_17997,N_16152,N_15724);
nand U17998 (N_17998,N_15025,N_16744);
and U17999 (N_17999,N_17438,N_16224);
and U18000 (N_18000,N_15652,N_15349);
nor U18001 (N_18001,N_16935,N_15820);
and U18002 (N_18002,N_16617,N_17454);
nor U18003 (N_18003,N_17110,N_16863);
or U18004 (N_18004,N_15051,N_15297);
nand U18005 (N_18005,N_15952,N_15510);
or U18006 (N_18006,N_16198,N_16560);
and U18007 (N_18007,N_15959,N_17276);
nor U18008 (N_18008,N_16271,N_17316);
nor U18009 (N_18009,N_17043,N_15922);
and U18010 (N_18010,N_15960,N_15730);
and U18011 (N_18011,N_16166,N_16556);
nand U18012 (N_18012,N_15949,N_16893);
nand U18013 (N_18013,N_17376,N_17357);
nor U18014 (N_18014,N_17012,N_15529);
nand U18015 (N_18015,N_16525,N_17146);
or U18016 (N_18016,N_15162,N_17044);
or U18017 (N_18017,N_17008,N_16962);
nand U18018 (N_18018,N_16899,N_16033);
and U18019 (N_18019,N_17104,N_17215);
or U18020 (N_18020,N_17076,N_15287);
nand U18021 (N_18021,N_15328,N_15117);
nor U18022 (N_18022,N_16294,N_15454);
nor U18023 (N_18023,N_17101,N_16821);
and U18024 (N_18024,N_16836,N_15300);
nor U18025 (N_18025,N_16257,N_17394);
and U18026 (N_18026,N_15125,N_17337);
and U18027 (N_18027,N_17251,N_15598);
and U18028 (N_18028,N_16639,N_15631);
and U18029 (N_18029,N_17422,N_15622);
or U18030 (N_18030,N_16488,N_16974);
nand U18031 (N_18031,N_16192,N_16458);
or U18032 (N_18032,N_15461,N_15203);
nand U18033 (N_18033,N_16268,N_17265);
nand U18034 (N_18034,N_15231,N_15234);
or U18035 (N_18035,N_17147,N_15086);
nand U18036 (N_18036,N_15876,N_16770);
nand U18037 (N_18037,N_15827,N_15308);
nor U18038 (N_18038,N_15289,N_17353);
nand U18039 (N_18039,N_16041,N_17190);
or U18040 (N_18040,N_17094,N_15235);
or U18041 (N_18041,N_17116,N_17494);
nand U18042 (N_18042,N_17208,N_16918);
nor U18043 (N_18043,N_16827,N_15481);
or U18044 (N_18044,N_16321,N_16598);
nor U18045 (N_18045,N_15240,N_16351);
or U18046 (N_18046,N_16008,N_16993);
nor U18047 (N_18047,N_15474,N_16357);
or U18048 (N_18048,N_16702,N_15318);
nor U18049 (N_18049,N_16280,N_15527);
xor U18050 (N_18050,N_15280,N_15484);
nor U18051 (N_18051,N_16761,N_16538);
nor U18052 (N_18052,N_16958,N_15126);
nand U18053 (N_18053,N_15658,N_15171);
and U18054 (N_18054,N_15832,N_16887);
nor U18055 (N_18055,N_15010,N_15354);
nand U18056 (N_18056,N_15856,N_17282);
and U18057 (N_18057,N_15590,N_15990);
and U18058 (N_18058,N_16415,N_16016);
nor U18059 (N_18059,N_16208,N_16476);
nand U18060 (N_18060,N_17412,N_17015);
and U18061 (N_18061,N_16005,N_16490);
or U18062 (N_18062,N_15522,N_17061);
nand U18063 (N_18063,N_15145,N_17144);
and U18064 (N_18064,N_17220,N_17107);
nand U18065 (N_18065,N_16401,N_17252);
nand U18066 (N_18066,N_16776,N_15540);
and U18067 (N_18067,N_15343,N_16002);
nand U18068 (N_18068,N_15871,N_17035);
and U18069 (N_18069,N_17408,N_16324);
xor U18070 (N_18070,N_15070,N_16309);
and U18071 (N_18071,N_15437,N_16388);
nor U18072 (N_18072,N_17312,N_15762);
or U18073 (N_18073,N_15858,N_15038);
or U18074 (N_18074,N_15368,N_17156);
and U18075 (N_18075,N_15353,N_16215);
and U18076 (N_18076,N_15133,N_15035);
and U18077 (N_18077,N_16147,N_15152);
or U18078 (N_18078,N_15135,N_17177);
nand U18079 (N_18079,N_16305,N_15558);
or U18080 (N_18080,N_15850,N_17113);
nor U18081 (N_18081,N_16242,N_16519);
and U18082 (N_18082,N_17188,N_17121);
and U18083 (N_18083,N_15148,N_16780);
and U18084 (N_18084,N_17183,N_17305);
nor U18085 (N_18085,N_15102,N_16077);
and U18086 (N_18086,N_15198,N_15725);
or U18087 (N_18087,N_17064,N_15286);
nand U18088 (N_18088,N_16627,N_16333);
or U18089 (N_18089,N_16402,N_16212);
nand U18090 (N_18090,N_15006,N_17228);
nand U18091 (N_18091,N_15880,N_15018);
and U18092 (N_18092,N_17330,N_15616);
and U18093 (N_18093,N_16861,N_17056);
or U18094 (N_18094,N_16645,N_15556);
or U18095 (N_18095,N_16233,N_15501);
or U18096 (N_18096,N_15605,N_16494);
and U18097 (N_18097,N_15361,N_16795);
or U18098 (N_18098,N_17136,N_15315);
and U18099 (N_18099,N_15576,N_17387);
nor U18100 (N_18100,N_16199,N_15928);
and U18101 (N_18101,N_15161,N_16569);
nor U18102 (N_18102,N_16742,N_16545);
or U18103 (N_18103,N_15782,N_15443);
and U18104 (N_18104,N_17073,N_15644);
or U18105 (N_18105,N_16638,N_15509);
and U18106 (N_18106,N_16052,N_16814);
nor U18107 (N_18107,N_15147,N_15069);
nor U18108 (N_18108,N_15305,N_15512);
xor U18109 (N_18109,N_15970,N_15111);
and U18110 (N_18110,N_17226,N_17062);
nor U18111 (N_18111,N_15660,N_16668);
or U18112 (N_18112,N_15703,N_15706);
xor U18113 (N_18113,N_15521,N_15586);
xnor U18114 (N_18114,N_16394,N_16944);
nor U18115 (N_18115,N_15324,N_17271);
nand U18116 (N_18116,N_15913,N_15030);
nor U18117 (N_18117,N_16698,N_16419);
and U18118 (N_18118,N_15153,N_16870);
and U18119 (N_18119,N_15258,N_15063);
nor U18120 (N_18120,N_15924,N_17129);
nand U18121 (N_18121,N_17052,N_16127);
nand U18122 (N_18122,N_15067,N_16164);
nand U18123 (N_18123,N_16101,N_15091);
nand U18124 (N_18124,N_16448,N_17268);
nand U18125 (N_18125,N_16258,N_15815);
nor U18126 (N_18126,N_16547,N_17459);
and U18127 (N_18127,N_16091,N_15571);
nand U18128 (N_18128,N_15742,N_15650);
nor U18129 (N_18129,N_16065,N_16793);
nand U18130 (N_18130,N_16468,N_17207);
and U18131 (N_18131,N_15889,N_16940);
nor U18132 (N_18132,N_17448,N_15759);
nor U18133 (N_18133,N_15688,N_15247);
and U18134 (N_18134,N_15346,N_16455);
nand U18135 (N_18135,N_15319,N_15967);
and U18136 (N_18136,N_15711,N_15723);
nand U18137 (N_18137,N_16352,N_17418);
nor U18138 (N_18138,N_17117,N_17363);
and U18139 (N_18139,N_17299,N_17091);
or U18140 (N_18140,N_16734,N_16107);
nor U18141 (N_18141,N_17397,N_15965);
nor U18142 (N_18142,N_15475,N_15144);
nand U18143 (N_18143,N_16852,N_16030);
nor U18144 (N_18144,N_15193,N_16412);
nor U18145 (N_18145,N_15539,N_16365);
and U18146 (N_18146,N_16105,N_16460);
nand U18147 (N_18147,N_16037,N_15322);
nand U18148 (N_18148,N_15802,N_16762);
nor U18149 (N_18149,N_16090,N_16677);
xnor U18150 (N_18150,N_16866,N_17057);
and U18151 (N_18151,N_16651,N_16006);
nand U18152 (N_18152,N_15047,N_17474);
and U18153 (N_18153,N_16159,N_16998);
nand U18154 (N_18154,N_15213,N_16472);
or U18155 (N_18155,N_17109,N_17469);
and U18156 (N_18156,N_15498,N_16134);
or U18157 (N_18157,N_17029,N_15741);
or U18158 (N_18158,N_16818,N_17097);
nand U18159 (N_18159,N_15351,N_17311);
or U18160 (N_18160,N_15619,N_17099);
xnor U18161 (N_18161,N_15455,N_16718);
or U18162 (N_18162,N_16699,N_15441);
or U18163 (N_18163,N_15136,N_15673);
nand U18164 (N_18164,N_17027,N_15735);
or U18165 (N_18165,N_15390,N_16666);
nand U18166 (N_18166,N_15120,N_17267);
nor U18167 (N_18167,N_16359,N_16640);
and U18168 (N_18168,N_16225,N_16686);
and U18169 (N_18169,N_16423,N_17361);
nor U18170 (N_18170,N_15721,N_15275);
and U18171 (N_18171,N_16672,N_16629);
nand U18172 (N_18172,N_15920,N_15392);
nand U18173 (N_18173,N_15955,N_15106);
and U18174 (N_18174,N_15130,N_16976);
and U18175 (N_18175,N_15530,N_15758);
or U18176 (N_18176,N_17442,N_16977);
nor U18177 (N_18177,N_16537,N_16145);
and U18178 (N_18178,N_17283,N_15490);
and U18179 (N_18179,N_17231,N_15119);
or U18180 (N_18180,N_15526,N_16012);
nand U18181 (N_18181,N_16185,N_17011);
nor U18182 (N_18182,N_17239,N_16097);
or U18183 (N_18183,N_16172,N_16933);
or U18184 (N_18184,N_16805,N_16413);
nand U18185 (N_18185,N_15877,N_16923);
nand U18186 (N_18186,N_15729,N_17004);
and U18187 (N_18187,N_15984,N_16927);
and U18188 (N_18188,N_16851,N_15930);
and U18189 (N_18189,N_15085,N_16555);
and U18190 (N_18190,N_15339,N_15074);
or U18191 (N_18191,N_15110,N_16806);
and U18192 (N_18192,N_15534,N_15969);
or U18193 (N_18193,N_17165,N_16289);
nand U18194 (N_18194,N_15818,N_16269);
and U18195 (N_18195,N_17164,N_16691);
and U18196 (N_18196,N_15357,N_16395);
or U18197 (N_18197,N_17067,N_16344);
and U18198 (N_18198,N_15626,N_17402);
nor U18199 (N_18199,N_17055,N_15317);
or U18200 (N_18200,N_16512,N_16045);
nor U18201 (N_18201,N_17296,N_15007);
or U18202 (N_18202,N_15024,N_17400);
and U18203 (N_18203,N_15399,N_16956);
nor U18204 (N_18204,N_15666,N_15387);
and U18205 (N_18205,N_17395,N_16284);
or U18206 (N_18206,N_15685,N_16422);
or U18207 (N_18207,N_15131,N_16459);
or U18208 (N_18208,N_15206,N_15114);
nand U18209 (N_18209,N_17264,N_15134);
nor U18210 (N_18210,N_17320,N_16587);
nor U18211 (N_18211,N_16287,N_17123);
and U18212 (N_18212,N_17358,N_16053);
nand U18213 (N_18213,N_15099,N_15419);
or U18214 (N_18214,N_16546,N_15382);
or U18215 (N_18215,N_16975,N_17019);
and U18216 (N_18216,N_15925,N_17321);
nand U18217 (N_18217,N_15862,N_15204);
nor U18218 (N_18218,N_16707,N_15405);
xnor U18219 (N_18219,N_16068,N_15621);
nor U18220 (N_18220,N_15467,N_17468);
nor U18221 (N_18221,N_16070,N_15093);
nand U18222 (N_18222,N_16196,N_15559);
nand U18223 (N_18223,N_16745,N_15634);
nor U18224 (N_18224,N_16094,N_16625);
or U18225 (N_18225,N_16632,N_16914);
nand U18226 (N_18226,N_16606,N_16642);
nor U18227 (N_18227,N_16708,N_15044);
nor U18228 (N_18228,N_16908,N_16250);
and U18229 (N_18229,N_16943,N_15202);
or U18230 (N_18230,N_16300,N_16725);
nand U18231 (N_18231,N_16210,N_16575);
and U18232 (N_18232,N_16819,N_17443);
and U18233 (N_18233,N_15901,N_17018);
and U18234 (N_18234,N_16399,N_16119);
nor U18235 (N_18235,N_16499,N_15495);
and U18236 (N_18236,N_16729,N_17182);
or U18237 (N_18237,N_16650,N_15581);
or U18238 (N_18238,N_16584,N_17290);
nor U18239 (N_18239,N_17495,N_15511);
and U18240 (N_18240,N_17227,N_15977);
or U18241 (N_18241,N_17022,N_16837);
nand U18242 (N_18242,N_15403,N_15896);
nor U18243 (N_18243,N_16753,N_16846);
nor U18244 (N_18244,N_17170,N_17317);
nor U18245 (N_18245,N_15485,N_17118);
nand U18246 (N_18246,N_15456,N_15643);
nor U18247 (N_18247,N_16260,N_16759);
nor U18248 (N_18248,N_16859,N_17452);
nor U18249 (N_18249,N_16563,N_17498);
nor U18250 (N_18250,N_16446,N_15045);
or U18251 (N_18251,N_15246,N_15472);
or U18252 (N_18252,N_15890,N_17106);
or U18253 (N_18253,N_16316,N_15299);
nor U18254 (N_18254,N_17399,N_16171);
nor U18255 (N_18255,N_16941,N_15691);
nand U18256 (N_18256,N_16046,N_16255);
nand U18257 (N_18257,N_15425,N_16532);
nand U18258 (N_18258,N_15076,N_15174);
and U18259 (N_18259,N_16965,N_16425);
and U18260 (N_18260,N_17081,N_15183);
and U18261 (N_18261,N_17470,N_16738);
or U18262 (N_18262,N_16117,N_15418);
or U18263 (N_18263,N_17411,N_17352);
and U18264 (N_18264,N_16599,N_16063);
nand U18265 (N_18265,N_16165,N_16922);
nand U18266 (N_18266,N_16849,N_16132);
nor U18267 (N_18267,N_16251,N_17275);
nand U18268 (N_18268,N_15929,N_15129);
xor U18269 (N_18269,N_16966,N_15551);
and U18270 (N_18270,N_16536,N_16404);
or U18271 (N_18271,N_16601,N_16028);
or U18272 (N_18272,N_16904,N_17301);
nor U18273 (N_18273,N_16314,N_16266);
nor U18274 (N_18274,N_15718,N_16756);
or U18275 (N_18275,N_17138,N_16055);
or U18276 (N_18276,N_15548,N_17288);
or U18277 (N_18277,N_16457,N_16905);
nand U18278 (N_18278,N_16288,N_15704);
and U18279 (N_18279,N_15434,N_15667);
nand U18280 (N_18280,N_16133,N_15751);
nor U18281 (N_18281,N_15307,N_16149);
or U18282 (N_18282,N_16652,N_15224);
nand U18283 (N_18283,N_16743,N_15716);
nand U18284 (N_18284,N_15589,N_15997);
and U18285 (N_18285,N_15081,N_16539);
nor U18286 (N_18286,N_17261,N_16868);
nor U18287 (N_18287,N_15537,N_16701);
or U18288 (N_18288,N_15033,N_15699);
or U18289 (N_18289,N_16577,N_15303);
nand U18290 (N_18290,N_15780,N_17380);
nand U18291 (N_18291,N_17472,N_15197);
and U18292 (N_18292,N_15531,N_16195);
nor U18293 (N_18293,N_15384,N_15451);
xnor U18294 (N_18294,N_15367,N_16315);
or U18295 (N_18295,N_16135,N_15789);
nand U18296 (N_18296,N_16082,N_17369);
nand U18297 (N_18297,N_15151,N_16023);
or U18298 (N_18298,N_15225,N_16847);
nand U18299 (N_18299,N_15291,N_15173);
or U18300 (N_18300,N_15865,N_15767);
nand U18301 (N_18301,N_15169,N_15516);
nor U18302 (N_18302,N_15505,N_15482);
or U18303 (N_18303,N_16785,N_15393);
or U18304 (N_18304,N_15881,N_17153);
or U18305 (N_18305,N_16515,N_17249);
and U18306 (N_18306,N_16405,N_15893);
and U18307 (N_18307,N_16466,N_15499);
nor U18308 (N_18308,N_17479,N_15914);
or U18309 (N_18309,N_16942,N_15810);
nand U18310 (N_18310,N_16741,N_17184);
and U18311 (N_18311,N_16274,N_16375);
nand U18312 (N_18312,N_16131,N_16435);
or U18313 (N_18313,N_16954,N_15625);
nand U18314 (N_18314,N_16580,N_15159);
and U18315 (N_18315,N_17423,N_15487);
nand U18316 (N_18316,N_16960,N_16291);
nor U18317 (N_18317,N_16913,N_16449);
nand U18318 (N_18318,N_17346,N_17401);
nor U18319 (N_18319,N_17089,N_15059);
or U18320 (N_18320,N_15974,N_16626);
and U18321 (N_18321,N_15344,N_15575);
and U18322 (N_18322,N_16832,N_17256);
or U18323 (N_18323,N_17273,N_15763);
nor U18324 (N_18324,N_16649,N_17245);
nand U18325 (N_18325,N_16229,N_16854);
nor U18326 (N_18326,N_15538,N_15533);
nand U18327 (N_18327,N_16491,N_17013);
nor U18328 (N_18328,N_16523,N_16211);
xnor U18329 (N_18329,N_15689,N_15184);
and U18330 (N_18330,N_16484,N_17457);
nor U18331 (N_18331,N_16125,N_16113);
nor U18332 (N_18332,N_16177,N_16372);
xnor U18333 (N_18333,N_15071,N_16461);
and U18334 (N_18334,N_15274,N_17020);
or U18335 (N_18335,N_16969,N_16029);
and U18336 (N_18336,N_16273,N_15694);
and U18337 (N_18337,N_17496,N_17217);
nand U18338 (N_18338,N_16583,N_16086);
and U18339 (N_18339,N_16768,N_15642);
nor U18340 (N_18340,N_16356,N_16949);
and U18341 (N_18341,N_15931,N_17071);
or U18342 (N_18342,N_16380,N_15116);
and U18343 (N_18343,N_15627,N_17093);
or U18344 (N_18344,N_16886,N_16777);
nor U18345 (N_18345,N_16594,N_17024);
and U18346 (N_18346,N_17198,N_17111);
or U18347 (N_18347,N_16169,N_15532);
and U18348 (N_18348,N_16367,N_15812);
nand U18349 (N_18349,N_15604,N_15489);
and U18350 (N_18350,N_15756,N_15773);
or U18351 (N_18351,N_16366,N_15108);
nor U18352 (N_18352,N_15838,N_16302);
and U18353 (N_18353,N_16481,N_15811);
nand U18354 (N_18354,N_15909,N_15453);
nor U18355 (N_18355,N_15668,N_15480);
nor U18356 (N_18356,N_17169,N_16374);
nor U18357 (N_18357,N_15679,N_15378);
nor U18358 (N_18358,N_17493,N_15423);
nor U18359 (N_18359,N_15971,N_15555);
and U18360 (N_18360,N_15347,N_17069);
nand U18361 (N_18361,N_16285,N_17172);
and U18362 (N_18362,N_16841,N_16391);
or U18363 (N_18363,N_16520,N_15687);
and U18364 (N_18364,N_16723,N_15910);
nand U18365 (N_18365,N_16564,N_17254);
nor U18366 (N_18366,N_17134,N_15471);
xor U18367 (N_18367,N_15615,N_17477);
nand U18368 (N_18368,N_17148,N_16903);
or U18369 (N_18369,N_16713,N_15325);
nand U18370 (N_18370,N_16141,N_16779);
or U18371 (N_18371,N_16791,N_17130);
nor U18372 (N_18372,N_16858,N_16953);
and U18373 (N_18373,N_15714,N_15866);
nor U18374 (N_18374,N_17028,N_15316);
or U18375 (N_18375,N_17236,N_15860);
nand U18376 (N_18376,N_15917,N_15869);
nand U18377 (N_18377,N_16480,N_16772);
nor U18378 (N_18378,N_16845,N_16176);
nor U18379 (N_18379,N_17037,N_17292);
or U18380 (N_18380,N_16184,N_16048);
or U18381 (N_18381,N_16234,N_15267);
xnor U18382 (N_18382,N_15011,N_15265);
and U18383 (N_18383,N_15003,N_15600);
nand U18384 (N_18384,N_16032,N_15369);
or U18385 (N_18385,N_15238,N_17074);
nor U18386 (N_18386,N_15582,N_16232);
nand U18387 (N_18387,N_16794,N_17384);
or U18388 (N_18388,N_15994,N_17499);
or U18389 (N_18389,N_15882,N_15021);
nor U18390 (N_18390,N_15424,N_15523);
nor U18391 (N_18391,N_16946,N_15670);
nand U18392 (N_18392,N_15784,N_16929);
and U18393 (N_18393,N_16614,N_16334);
or U18394 (N_18394,N_16920,N_15262);
nand U18395 (N_18395,N_15008,N_17248);
or U18396 (N_18396,N_15809,N_16660);
nor U18397 (N_18397,N_15765,N_15072);
nand U18398 (N_18398,N_16191,N_16990);
or U18399 (N_18399,N_15580,N_15502);
nor U18400 (N_18400,N_16813,N_17339);
and U18401 (N_18401,N_16680,N_16429);
nand U18402 (N_18402,N_16675,N_15386);
or U18403 (N_18403,N_15066,N_16767);
and U18404 (N_18404,N_17210,N_15745);
and U18405 (N_18405,N_15037,N_17135);
or U18406 (N_18406,N_15682,N_16303);
nand U18407 (N_18407,N_16688,N_16439);
and U18408 (N_18408,N_16054,N_16667);
nor U18409 (N_18409,N_17213,N_16963);
nand U18410 (N_18410,N_17359,N_15064);
and U18411 (N_18411,N_15479,N_16658);
nand U18412 (N_18412,N_15459,N_17103);
or U18413 (N_18413,N_16081,N_15277);
and U18414 (N_18414,N_16452,N_16540);
and U18415 (N_18415,N_16885,N_16084);
nand U18416 (N_18416,N_16338,N_16044);
nor U18417 (N_18417,N_17046,N_16140);
or U18418 (N_18418,N_16178,N_16464);
or U18419 (N_18419,N_15963,N_16247);
nand U18420 (N_18420,N_16410,N_16824);
or U18421 (N_18421,N_15843,N_15292);
and U18422 (N_18422,N_16631,N_17102);
xor U18423 (N_18423,N_17281,N_15841);
nor U18424 (N_18424,N_15676,N_16329);
or U18425 (N_18425,N_15462,N_16186);
or U18426 (N_18426,N_17200,N_15417);
nand U18427 (N_18427,N_16406,N_16179);
nand U18428 (N_18428,N_17016,N_15543);
and U18429 (N_18429,N_16350,N_16856);
xor U18430 (N_18430,N_16925,N_16221);
or U18431 (N_18431,N_17247,N_17007);
and U18432 (N_18432,N_17463,N_15348);
nand U18433 (N_18433,N_15402,N_16080);
or U18434 (N_18434,N_17072,N_15747);
or U18435 (N_18435,N_16437,N_17086);
nand U18436 (N_18436,N_16444,N_16711);
nand U18437 (N_18437,N_17377,N_16493);
and U18438 (N_18438,N_16612,N_15180);
nor U18439 (N_18439,N_17295,N_15041);
and U18440 (N_18440,N_16992,N_17427);
nor U18441 (N_18441,N_16514,N_15878);
nor U18442 (N_18442,N_15398,N_16800);
nand U18443 (N_18443,N_15433,N_16613);
nand U18444 (N_18444,N_15154,N_16430);
or U18445 (N_18445,N_17293,N_15888);
and U18446 (N_18446,N_15226,N_15105);
or U18447 (N_18447,N_16364,N_16471);
or U18448 (N_18448,N_15794,N_17068);
or U18449 (N_18449,N_16890,N_17030);
or U18450 (N_18450,N_16389,N_15380);
nor U18451 (N_18451,N_16826,N_16416);
and U18452 (N_18452,N_16015,N_16733);
nand U18453 (N_18453,N_16829,N_17287);
nand U18454 (N_18454,N_17039,N_15218);
or U18455 (N_18455,N_16261,N_17471);
nand U18456 (N_18456,N_17270,N_15301);
nand U18457 (N_18457,N_16714,N_15341);
nand U18458 (N_18458,N_16010,N_17492);
nor U18459 (N_18459,N_15550,N_15473);
and U18460 (N_18460,N_16771,N_16340);
nand U18461 (N_18461,N_15506,N_16290);
nand U18462 (N_18462,N_16355,N_17404);
nor U18463 (N_18463,N_15429,N_15073);
or U18464 (N_18464,N_15900,N_17428);
nand U18465 (N_18465,N_15926,N_16408);
or U18466 (N_18466,N_17141,N_16586);
nand U18467 (N_18467,N_15713,N_15446);
and U18468 (N_18468,N_17426,N_17174);
and U18469 (N_18469,N_15269,N_17114);
nand U18470 (N_18470,N_15142,N_15772);
nor U18471 (N_18471,N_15271,N_15781);
nand U18472 (N_18472,N_16978,N_17070);
and U18473 (N_18473,N_15288,N_16644);
nand U18474 (N_18474,N_15312,N_15122);
or U18475 (N_18475,N_15542,N_17222);
or U18476 (N_18476,N_16306,N_16902);
or U18477 (N_18477,N_16611,N_17453);
or U18478 (N_18478,N_16562,N_15641);
nor U18479 (N_18479,N_15799,N_17456);
and U18480 (N_18480,N_16731,N_15731);
and U18481 (N_18481,N_15995,N_16175);
nand U18482 (N_18482,N_17149,N_16897);
nand U18483 (N_18483,N_15715,N_15945);
or U18484 (N_18484,N_15026,N_15514);
nor U18485 (N_18485,N_16880,N_15594);
or U18486 (N_18486,N_15845,N_16237);
nor U18487 (N_18487,N_15708,N_15207);
and U18488 (N_18488,N_16019,N_15313);
nand U18489 (N_18489,N_15228,N_15428);
nor U18490 (N_18490,N_16469,N_15285);
nand U18491 (N_18491,N_15567,N_17466);
nor U18492 (N_18492,N_17319,N_17233);
and U18493 (N_18493,N_16624,N_15633);
nand U18494 (N_18494,N_16985,N_15000);
nand U18495 (N_18495,N_17023,N_16108);
nor U18496 (N_18496,N_15201,N_16690);
nand U18497 (N_18497,N_15635,N_17432);
nand U18498 (N_18498,N_15327,N_16479);
nor U18499 (N_18499,N_16436,N_16067);
nor U18500 (N_18500,N_17216,N_16293);
and U18501 (N_18501,N_16534,N_15743);
nor U18502 (N_18502,N_17125,N_15491);
nor U18503 (N_18503,N_15486,N_17124);
and U18504 (N_18504,N_16325,N_16498);
nor U18505 (N_18505,N_15230,N_15894);
or U18506 (N_18506,N_15296,N_16894);
or U18507 (N_18507,N_16619,N_16362);
nor U18508 (N_18508,N_16353,N_16883);
and U18509 (N_18509,N_16383,N_15342);
nand U18510 (N_18510,N_15885,N_16017);
or U18511 (N_18511,N_16531,N_15638);
or U18512 (N_18512,N_16623,N_15413);
nand U18513 (N_18513,N_17230,N_16765);
nor U18514 (N_18514,N_15250,N_17229);
nand U18515 (N_18515,N_16000,N_16752);
and U18516 (N_18516,N_15270,N_15139);
and U18517 (N_18517,N_15675,N_15414);
nor U18518 (N_18518,N_15276,N_16979);
xor U18519 (N_18519,N_17285,N_15253);
nand U18520 (N_18520,N_16740,N_17026);
and U18521 (N_18521,N_15599,N_16735);
xor U18522 (N_18522,N_16489,N_16574);
nor U18523 (N_18523,N_15602,N_16386);
or U18524 (N_18524,N_15857,N_17066);
and U18525 (N_18525,N_17128,N_15345);
or U18526 (N_18526,N_17053,N_15310);
and U18527 (N_18527,N_15861,N_17302);
or U18528 (N_18528,N_15331,N_15662);
and U18529 (N_18529,N_15587,N_17060);
and U18530 (N_18530,N_16647,N_16955);
or U18531 (N_18531,N_15077,N_15853);
or U18532 (N_18532,N_15916,N_15508);
and U18533 (N_18533,N_16102,N_16440);
or U18534 (N_18534,N_16637,N_17391);
or U18535 (N_18535,N_15942,N_15757);
or U18536 (N_18536,N_15863,N_15515);
nor U18537 (N_18537,N_15948,N_15553);
nor U18538 (N_18538,N_16544,N_15493);
and U18539 (N_18539,N_17206,N_17090);
nor U18540 (N_18540,N_17010,N_17340);
nand U18541 (N_18541,N_15771,N_16463);
and U18542 (N_18542,N_16061,N_15720);
nor U18543 (N_18543,N_15379,N_16656);
xor U18544 (N_18544,N_15239,N_16207);
or U18545 (N_18545,N_16319,N_16906);
nor U18546 (N_18546,N_16297,N_15761);
and U18547 (N_18547,N_16798,N_16339);
and U18548 (N_18548,N_15476,N_16025);
or U18549 (N_18549,N_16148,N_16018);
nor U18550 (N_18550,N_15320,N_16822);
nor U18551 (N_18551,N_16168,N_17356);
and U18552 (N_18552,N_15364,N_17166);
nand U18553 (N_18553,N_15217,N_17084);
and U18554 (N_18554,N_16219,N_17417);
or U18555 (N_18555,N_16343,N_16482);
or U18556 (N_18556,N_16040,N_15932);
or U18557 (N_18557,N_15733,N_15935);
nand U18558 (N_18558,N_16203,N_15055);
and U18559 (N_18559,N_15334,N_16600);
nor U18560 (N_18560,N_16424,N_15261);
nor U18561 (N_18561,N_17300,N_17278);
xnor U18562 (N_18562,N_16099,N_15020);
and U18563 (N_18563,N_17307,N_16892);
or U18564 (N_18564,N_17306,N_16792);
or U18565 (N_18565,N_15447,N_16815);
nor U18566 (N_18566,N_16079,N_15937);
nand U18567 (N_18567,N_15978,N_17424);
or U18568 (N_18568,N_16530,N_17425);
or U18569 (N_18569,N_16118,N_16390);
or U18570 (N_18570,N_16607,N_15103);
or U18571 (N_18571,N_15569,N_16518);
and U18572 (N_18572,N_15363,N_16746);
or U18573 (N_18573,N_15397,N_16576);
nand U18574 (N_18574,N_17075,N_15693);
or U18575 (N_18575,N_15680,N_15464);
nand U18576 (N_18576,N_15541,N_16170);
nor U18577 (N_18577,N_16811,N_16825);
nor U18578 (N_18578,N_15999,N_16223);
nor U18579 (N_18579,N_16784,N_16013);
or U18580 (N_18580,N_16064,N_16533);
and U18581 (N_18581,N_15774,N_16840);
nor U18582 (N_18582,N_17375,N_15613);
nand U18583 (N_18583,N_16674,N_16264);
or U18584 (N_18584,N_17289,N_16665);
and U18585 (N_18585,N_15785,N_17145);
and U18586 (N_18586,N_16100,N_15940);
nor U18587 (N_18587,N_16939,N_17178);
and U18588 (N_18588,N_17354,N_15777);
or U18589 (N_18589,N_15753,N_15883);
or U18590 (N_18590,N_17446,N_15829);
or U18591 (N_18591,N_16994,N_16855);
nand U18592 (N_18592,N_16011,N_15273);
and U18593 (N_18593,N_16669,N_16279);
nand U18594 (N_18594,N_16427,N_16912);
nand U18595 (N_18595,N_16937,N_15636);
and U18596 (N_18596,N_15208,N_17393);
nand U18597 (N_18597,N_15639,N_15637);
nor U18598 (N_18598,N_17137,N_15577);
and U18599 (N_18599,N_15168,N_15504);
or U18600 (N_18600,N_15915,N_17414);
nand U18601 (N_18601,N_17085,N_16703);
nand U18602 (N_18602,N_15395,N_15546);
and U18603 (N_18603,N_16504,N_16103);
nand U18604 (N_18604,N_15852,N_16421);
or U18605 (N_18605,N_16522,N_17489);
nand U18606 (N_18606,N_17345,N_15100);
and U18607 (N_18607,N_16948,N_16833);
nor U18608 (N_18608,N_16400,N_17410);
nor U18609 (N_18609,N_16719,N_17092);
nand U18610 (N_18610,N_15185,N_16558);
and U18611 (N_18611,N_15137,N_16999);
and U18612 (N_18612,N_15919,N_17338);
or U18613 (N_18613,N_16200,N_16764);
nor U18614 (N_18614,N_16812,N_17196);
nor U18615 (N_18615,N_16554,N_17304);
nand U18616 (N_18616,N_15872,N_15748);
or U18617 (N_18617,N_15340,N_17045);
and U18618 (N_18618,N_15584,N_15912);
and U18619 (N_18619,N_16874,N_15661);
and U18620 (N_18620,N_17235,N_16782);
or U18621 (N_18621,N_16716,N_17241);
and U18622 (N_18622,N_17036,N_15754);
or U18623 (N_18623,N_17058,N_15975);
or U18624 (N_18624,N_16828,N_15983);
nand U18625 (N_18625,N_15570,N_17127);
and U18626 (N_18626,N_17284,N_16526);
nand U18627 (N_18627,N_16657,N_16485);
and U18628 (N_18628,N_15927,N_16693);
or U18629 (N_18629,N_16542,N_15362);
xor U18630 (N_18630,N_16304,N_16230);
nor U18631 (N_18631,N_15717,N_16035);
nor U18632 (N_18632,N_17434,N_15015);
nor U18633 (N_18633,N_16163,N_15624);
or U18634 (N_18634,N_15806,N_15127);
nand U18635 (N_18635,N_17246,N_15436);
and U18636 (N_18636,N_16769,N_17473);
nand U18637 (N_18637,N_16193,N_16426);
nor U18638 (N_18638,N_16360,N_16501);
and U18639 (N_18639,N_15438,N_15854);
and U18640 (N_18640,N_15266,N_17449);
nor U18641 (N_18641,N_17051,N_16695);
and U18642 (N_18642,N_15836,N_15864);
xnor U18643 (N_18643,N_15256,N_15980);
or U18644 (N_18644,N_15061,N_15768);
and U18645 (N_18645,N_15389,N_16633);
nand U18646 (N_18646,N_17455,N_15046);
and U18647 (N_18647,N_17150,N_17112);
and U18648 (N_18648,N_17309,N_15189);
nand U18649 (N_18649,N_17458,N_15611);
or U18650 (N_18650,N_17389,N_15031);
and U18651 (N_18651,N_15330,N_16981);
or U18652 (N_18652,N_15851,N_17240);
or U18653 (N_18653,N_15422,N_15236);
and U18654 (N_18654,N_15837,N_17151);
xor U18655 (N_18655,N_17054,N_16582);
and U18656 (N_18656,N_17041,N_15807);
and U18657 (N_18657,N_15259,N_15821);
nor U18658 (N_18658,N_17435,N_15620);
or U18659 (N_18659,N_15953,N_16681);
nor U18660 (N_18660,N_16597,N_15736);
or U18661 (N_18661,N_16959,N_16952);
nor U18662 (N_18662,N_16475,N_15053);
and U18663 (N_18663,N_15043,N_15561);
nand U18664 (N_18664,N_15918,N_15058);
nand U18665 (N_18665,N_15719,N_15188);
nand U18666 (N_18666,N_16095,N_15798);
nor U18667 (N_18667,N_15056,N_15764);
nand U18668 (N_18668,N_17167,N_17224);
nand U18669 (N_18669,N_15623,N_15373);
or U18670 (N_18670,N_15677,N_16835);
nand U18671 (N_18671,N_16551,N_15321);
nand U18672 (N_18672,N_17234,N_16050);
or U18673 (N_18673,N_16510,N_15166);
or U18674 (N_18674,N_16453,N_15075);
nor U18675 (N_18675,N_15898,N_16073);
and U18676 (N_18676,N_16717,N_16561);
or U18677 (N_18677,N_15057,N_16524);
nor U18678 (N_18678,N_15084,N_15737);
nand U18679 (N_18679,N_16848,N_16241);
or U18680 (N_18680,N_16130,N_16755);
nor U18681 (N_18681,N_17484,N_15859);
nor U18682 (N_18682,N_16720,N_15128);
nor U18683 (N_18683,N_15268,N_16298);
or U18684 (N_18684,N_16278,N_17328);
nor U18685 (N_18685,N_16507,N_15544);
nor U18686 (N_18686,N_16197,N_17105);
and U18687 (N_18687,N_16773,N_16529);
and U18688 (N_18688,N_15019,N_15709);
xor U18689 (N_18689,N_16869,N_17420);
or U18690 (N_18690,N_15196,N_15698);
nor U18691 (N_18691,N_15177,N_15695);
nor U18692 (N_18692,N_15293,N_16106);
and U18693 (N_18693,N_15683,N_16190);
nor U18694 (N_18694,N_17017,N_15830);
or U18695 (N_18695,N_15585,N_17126);
nand U18696 (N_18696,N_16502,N_17327);
nand U18697 (N_18697,N_15903,N_15421);
and U18698 (N_18698,N_16038,N_16034);
or U18699 (N_18699,N_16543,N_15377);
or U18700 (N_18700,N_15744,N_15249);
or U18701 (N_18701,N_15427,N_16550);
and U18702 (N_18702,N_15776,N_16988);
nand U18703 (N_18703,N_16218,N_17063);
nand U18704 (N_18704,N_16262,N_15112);
and U18705 (N_18705,N_16997,N_16595);
and U18706 (N_18706,N_15936,N_16889);
and U18707 (N_18707,N_16609,N_15545);
and U18708 (N_18708,N_15528,N_16758);
or U18709 (N_18709,N_16156,N_16552);
and U18710 (N_18710,N_16616,N_15563);
nor U18711 (N_18711,N_16706,N_16228);
nor U18712 (N_18712,N_16535,N_16270);
or U18713 (N_18713,N_15205,N_16060);
nor U18714 (N_18714,N_17269,N_15005);
nor U18715 (N_18715,N_15705,N_16154);
xor U18716 (N_18716,N_15029,N_16104);
or U18717 (N_18717,N_16984,N_17132);
and U18718 (N_18718,N_16559,N_15233);
xor U18719 (N_18719,N_16628,N_16110);
xor U18720 (N_18720,N_15143,N_16246);
nor U18721 (N_18721,N_15420,N_16465);
nand U18722 (N_18722,N_16754,N_17349);
nand U18723 (N_18723,N_17152,N_16676);
and U18724 (N_18724,N_16144,N_16275);
or U18725 (N_18725,N_16451,N_15547);
nand U18726 (N_18726,N_15095,N_16378);
and U18727 (N_18727,N_16697,N_16418);
nand U18728 (N_18728,N_17157,N_15597);
and U18729 (N_18729,N_16610,N_15432);
nor U18730 (N_18730,N_16682,N_15593);
or U18731 (N_18731,N_15350,N_16763);
nor U18732 (N_18732,N_15991,N_16150);
or U18733 (N_18733,N_16450,N_16126);
nand U18734 (N_18734,N_15245,N_17195);
and U18735 (N_18735,N_17257,N_15264);
and U18736 (N_18736,N_16272,N_15808);
nand U18737 (N_18737,N_15042,N_16473);
or U18738 (N_18738,N_15897,N_16098);
nor U18739 (N_18739,N_15697,N_17385);
xor U18740 (N_18740,N_15016,N_15796);
and U18741 (N_18741,N_16951,N_16454);
nand U18742 (N_18742,N_16142,N_17154);
and U18743 (N_18743,N_16907,N_17403);
nor U18744 (N_18744,N_16980,N_15052);
nor U18745 (N_18745,N_17087,N_16704);
nand U18746 (N_18746,N_16622,N_15792);
and U18747 (N_18747,N_17371,N_17080);
nand U18748 (N_18748,N_15439,N_16732);
nand U18749 (N_18749,N_17383,N_17308);
or U18750 (N_18750,N_16810,N_15267);
nor U18751 (N_18751,N_15115,N_16874);
nor U18752 (N_18752,N_15597,N_17150);
or U18753 (N_18753,N_16918,N_16245);
or U18754 (N_18754,N_16501,N_16767);
and U18755 (N_18755,N_16021,N_17138);
nor U18756 (N_18756,N_16894,N_15437);
or U18757 (N_18757,N_15193,N_15803);
and U18758 (N_18758,N_16294,N_16960);
and U18759 (N_18759,N_15539,N_16844);
and U18760 (N_18760,N_15121,N_17018);
nor U18761 (N_18761,N_17330,N_15842);
or U18762 (N_18762,N_15461,N_15535);
nor U18763 (N_18763,N_17047,N_16291);
or U18764 (N_18764,N_17112,N_17158);
nand U18765 (N_18765,N_16520,N_15162);
and U18766 (N_18766,N_16580,N_16258);
nor U18767 (N_18767,N_16310,N_16618);
nand U18768 (N_18768,N_17156,N_15564);
nand U18769 (N_18769,N_17474,N_16228);
nor U18770 (N_18770,N_16427,N_15089);
nor U18771 (N_18771,N_15034,N_16585);
and U18772 (N_18772,N_16334,N_15811);
and U18773 (N_18773,N_16450,N_16902);
and U18774 (N_18774,N_15110,N_16241);
and U18775 (N_18775,N_15869,N_15876);
and U18776 (N_18776,N_17482,N_17475);
or U18777 (N_18777,N_17428,N_17166);
and U18778 (N_18778,N_16137,N_16172);
and U18779 (N_18779,N_16402,N_17352);
and U18780 (N_18780,N_17319,N_16714);
or U18781 (N_18781,N_16029,N_16648);
nand U18782 (N_18782,N_16145,N_16672);
nand U18783 (N_18783,N_17304,N_16931);
nor U18784 (N_18784,N_16718,N_16215);
nand U18785 (N_18785,N_15000,N_16692);
nor U18786 (N_18786,N_16226,N_16351);
or U18787 (N_18787,N_15926,N_16806);
and U18788 (N_18788,N_15393,N_16047);
nor U18789 (N_18789,N_16764,N_16235);
nor U18790 (N_18790,N_16002,N_15305);
or U18791 (N_18791,N_15477,N_16354);
and U18792 (N_18792,N_16260,N_16607);
or U18793 (N_18793,N_16527,N_16025);
xnor U18794 (N_18794,N_15552,N_17173);
and U18795 (N_18795,N_16344,N_15337);
nand U18796 (N_18796,N_17159,N_17153);
xnor U18797 (N_18797,N_16128,N_16994);
and U18798 (N_18798,N_17175,N_16609);
and U18799 (N_18799,N_15461,N_15771);
xor U18800 (N_18800,N_15683,N_15100);
nand U18801 (N_18801,N_15255,N_17085);
and U18802 (N_18802,N_17202,N_16353);
nor U18803 (N_18803,N_15020,N_16688);
nand U18804 (N_18804,N_15361,N_15124);
and U18805 (N_18805,N_17222,N_16541);
nand U18806 (N_18806,N_16764,N_15958);
or U18807 (N_18807,N_17220,N_16982);
nor U18808 (N_18808,N_16844,N_17495);
and U18809 (N_18809,N_16906,N_16848);
and U18810 (N_18810,N_15268,N_16328);
nand U18811 (N_18811,N_17241,N_16649);
or U18812 (N_18812,N_16018,N_17152);
or U18813 (N_18813,N_17218,N_16634);
nor U18814 (N_18814,N_17301,N_17416);
and U18815 (N_18815,N_15501,N_16625);
or U18816 (N_18816,N_15241,N_15651);
nand U18817 (N_18817,N_17173,N_16831);
nand U18818 (N_18818,N_16651,N_15850);
nor U18819 (N_18819,N_16588,N_15523);
or U18820 (N_18820,N_17406,N_16475);
nand U18821 (N_18821,N_17055,N_16568);
or U18822 (N_18822,N_16782,N_16738);
xor U18823 (N_18823,N_17134,N_15916);
and U18824 (N_18824,N_15496,N_15528);
or U18825 (N_18825,N_15268,N_17139);
or U18826 (N_18826,N_17310,N_15298);
and U18827 (N_18827,N_15024,N_15682);
and U18828 (N_18828,N_15649,N_17118);
or U18829 (N_18829,N_16228,N_16692);
nand U18830 (N_18830,N_15595,N_15434);
nor U18831 (N_18831,N_17352,N_15053);
nor U18832 (N_18832,N_17209,N_16123);
and U18833 (N_18833,N_17333,N_15645);
or U18834 (N_18834,N_17455,N_17460);
nor U18835 (N_18835,N_15954,N_16022);
and U18836 (N_18836,N_16757,N_16203);
and U18837 (N_18837,N_17439,N_17018);
or U18838 (N_18838,N_16246,N_16780);
nor U18839 (N_18839,N_16703,N_15906);
or U18840 (N_18840,N_16592,N_16873);
and U18841 (N_18841,N_15040,N_16873);
xnor U18842 (N_18842,N_15965,N_15863);
and U18843 (N_18843,N_15580,N_16836);
or U18844 (N_18844,N_16814,N_15551);
or U18845 (N_18845,N_17353,N_16575);
nor U18846 (N_18846,N_16545,N_15053);
nor U18847 (N_18847,N_15053,N_15469);
and U18848 (N_18848,N_16726,N_16465);
or U18849 (N_18849,N_16229,N_16411);
and U18850 (N_18850,N_15928,N_16631);
nand U18851 (N_18851,N_17105,N_16705);
nand U18852 (N_18852,N_16079,N_16209);
nor U18853 (N_18853,N_16780,N_15042);
and U18854 (N_18854,N_15574,N_16606);
nor U18855 (N_18855,N_15079,N_17142);
nor U18856 (N_18856,N_16838,N_17463);
nand U18857 (N_18857,N_15228,N_15508);
nand U18858 (N_18858,N_16435,N_17127);
nor U18859 (N_18859,N_15163,N_17446);
or U18860 (N_18860,N_16872,N_15782);
nor U18861 (N_18861,N_16021,N_17431);
nor U18862 (N_18862,N_16396,N_15145);
or U18863 (N_18863,N_16878,N_17199);
nor U18864 (N_18864,N_15304,N_16591);
nor U18865 (N_18865,N_16608,N_17435);
or U18866 (N_18866,N_15463,N_16899);
or U18867 (N_18867,N_15059,N_16949);
or U18868 (N_18868,N_16914,N_16766);
and U18869 (N_18869,N_15074,N_15947);
nor U18870 (N_18870,N_17236,N_16948);
and U18871 (N_18871,N_15653,N_16615);
xnor U18872 (N_18872,N_15431,N_16627);
and U18873 (N_18873,N_15515,N_16609);
nand U18874 (N_18874,N_17496,N_15954);
and U18875 (N_18875,N_17346,N_17132);
nand U18876 (N_18876,N_17271,N_15209);
nand U18877 (N_18877,N_16264,N_16243);
and U18878 (N_18878,N_16629,N_15030);
or U18879 (N_18879,N_15874,N_16006);
nor U18880 (N_18880,N_17101,N_16415);
and U18881 (N_18881,N_16363,N_15630);
and U18882 (N_18882,N_16363,N_15840);
nand U18883 (N_18883,N_17148,N_16063);
and U18884 (N_18884,N_15192,N_17394);
nor U18885 (N_18885,N_16605,N_16511);
and U18886 (N_18886,N_15956,N_15994);
or U18887 (N_18887,N_16789,N_16856);
nand U18888 (N_18888,N_16855,N_16847);
or U18889 (N_18889,N_15325,N_15003);
or U18890 (N_18890,N_16748,N_15422);
or U18891 (N_18891,N_15353,N_17258);
and U18892 (N_18892,N_16793,N_16738);
nor U18893 (N_18893,N_15270,N_17163);
or U18894 (N_18894,N_15235,N_15945);
and U18895 (N_18895,N_15763,N_17032);
xor U18896 (N_18896,N_16112,N_16235);
and U18897 (N_18897,N_16391,N_17296);
or U18898 (N_18898,N_17411,N_15280);
and U18899 (N_18899,N_16197,N_15846);
or U18900 (N_18900,N_17264,N_15989);
and U18901 (N_18901,N_16078,N_17113);
nand U18902 (N_18902,N_16921,N_16039);
or U18903 (N_18903,N_15179,N_15100);
nand U18904 (N_18904,N_17275,N_16567);
or U18905 (N_18905,N_15218,N_16968);
and U18906 (N_18906,N_16355,N_15212);
or U18907 (N_18907,N_16920,N_16605);
xnor U18908 (N_18908,N_15849,N_17292);
nor U18909 (N_18909,N_15358,N_15793);
nand U18910 (N_18910,N_16088,N_15672);
nor U18911 (N_18911,N_17335,N_16143);
and U18912 (N_18912,N_15496,N_15549);
xor U18913 (N_18913,N_15244,N_16799);
and U18914 (N_18914,N_16648,N_16560);
nor U18915 (N_18915,N_16518,N_15329);
nand U18916 (N_18916,N_16065,N_16105);
nand U18917 (N_18917,N_16715,N_15679);
nand U18918 (N_18918,N_15342,N_16013);
nand U18919 (N_18919,N_15616,N_15246);
or U18920 (N_18920,N_17259,N_15105);
nor U18921 (N_18921,N_16232,N_16784);
nor U18922 (N_18922,N_15804,N_16843);
nand U18923 (N_18923,N_15543,N_16995);
nor U18924 (N_18924,N_17472,N_17270);
xnor U18925 (N_18925,N_16317,N_16764);
nor U18926 (N_18926,N_15418,N_15053);
and U18927 (N_18927,N_16939,N_16830);
nor U18928 (N_18928,N_15822,N_16638);
nor U18929 (N_18929,N_17318,N_17090);
nand U18930 (N_18930,N_15047,N_17104);
nand U18931 (N_18931,N_15962,N_17325);
nor U18932 (N_18932,N_17425,N_15410);
nor U18933 (N_18933,N_15845,N_15290);
or U18934 (N_18934,N_15319,N_16062);
and U18935 (N_18935,N_16735,N_16700);
or U18936 (N_18936,N_17060,N_17348);
or U18937 (N_18937,N_15274,N_15966);
nand U18938 (N_18938,N_16855,N_16408);
nor U18939 (N_18939,N_16764,N_15087);
nand U18940 (N_18940,N_16533,N_15571);
and U18941 (N_18941,N_17150,N_16973);
or U18942 (N_18942,N_16049,N_15128);
nor U18943 (N_18943,N_16787,N_15956);
and U18944 (N_18944,N_16529,N_16652);
and U18945 (N_18945,N_17055,N_16461);
or U18946 (N_18946,N_16860,N_15451);
or U18947 (N_18947,N_16317,N_16344);
and U18948 (N_18948,N_17449,N_15308);
or U18949 (N_18949,N_16108,N_15904);
nor U18950 (N_18950,N_16702,N_16206);
and U18951 (N_18951,N_16166,N_15347);
nor U18952 (N_18952,N_15711,N_16412);
nand U18953 (N_18953,N_15671,N_15231);
nand U18954 (N_18954,N_16819,N_16069);
and U18955 (N_18955,N_15759,N_15318);
nand U18956 (N_18956,N_17149,N_17469);
xor U18957 (N_18957,N_15470,N_17224);
or U18958 (N_18958,N_15933,N_16600);
and U18959 (N_18959,N_16096,N_16763);
or U18960 (N_18960,N_15710,N_17225);
nor U18961 (N_18961,N_15929,N_15167);
or U18962 (N_18962,N_16489,N_17300);
xor U18963 (N_18963,N_15242,N_17489);
and U18964 (N_18964,N_15292,N_16421);
or U18965 (N_18965,N_17255,N_17066);
or U18966 (N_18966,N_17450,N_15853);
or U18967 (N_18967,N_16944,N_16408);
nor U18968 (N_18968,N_16836,N_17147);
and U18969 (N_18969,N_15820,N_16109);
xnor U18970 (N_18970,N_16475,N_15159);
nor U18971 (N_18971,N_17351,N_15317);
and U18972 (N_18972,N_17438,N_16621);
and U18973 (N_18973,N_16888,N_15636);
or U18974 (N_18974,N_15137,N_15222);
nor U18975 (N_18975,N_17220,N_15340);
xnor U18976 (N_18976,N_17187,N_15684);
or U18977 (N_18977,N_16691,N_16747);
nor U18978 (N_18978,N_16441,N_17051);
nor U18979 (N_18979,N_16685,N_17313);
and U18980 (N_18980,N_16442,N_16511);
or U18981 (N_18981,N_15332,N_16938);
nand U18982 (N_18982,N_16974,N_17438);
and U18983 (N_18983,N_15303,N_17002);
nor U18984 (N_18984,N_16921,N_15987);
nor U18985 (N_18985,N_15927,N_16091);
nand U18986 (N_18986,N_16880,N_16004);
and U18987 (N_18987,N_17397,N_15258);
or U18988 (N_18988,N_16039,N_17443);
xnor U18989 (N_18989,N_17182,N_16426);
and U18990 (N_18990,N_15278,N_17027);
nand U18991 (N_18991,N_17113,N_15932);
nand U18992 (N_18992,N_16949,N_15435);
nand U18993 (N_18993,N_15445,N_16106);
or U18994 (N_18994,N_16419,N_16066);
nand U18995 (N_18995,N_16698,N_15357);
or U18996 (N_18996,N_16959,N_16031);
and U18997 (N_18997,N_16673,N_16063);
or U18998 (N_18998,N_16103,N_15910);
and U18999 (N_18999,N_17199,N_15966);
nor U19000 (N_19000,N_15275,N_17159);
nor U19001 (N_19001,N_17345,N_16816);
and U19002 (N_19002,N_15249,N_15212);
and U19003 (N_19003,N_17151,N_17216);
or U19004 (N_19004,N_16400,N_15755);
nor U19005 (N_19005,N_15696,N_15935);
and U19006 (N_19006,N_16086,N_16655);
and U19007 (N_19007,N_15086,N_17237);
and U19008 (N_19008,N_15747,N_16446);
nand U19009 (N_19009,N_16035,N_16210);
and U19010 (N_19010,N_15766,N_17084);
or U19011 (N_19011,N_15847,N_17440);
nand U19012 (N_19012,N_16256,N_15539);
and U19013 (N_19013,N_15874,N_15048);
and U19014 (N_19014,N_15293,N_17138);
nand U19015 (N_19015,N_15374,N_16652);
and U19016 (N_19016,N_17309,N_15729);
and U19017 (N_19017,N_15616,N_15500);
and U19018 (N_19018,N_16218,N_17053);
xnor U19019 (N_19019,N_17404,N_15449);
and U19020 (N_19020,N_15852,N_15219);
and U19021 (N_19021,N_16511,N_15577);
nor U19022 (N_19022,N_17281,N_16749);
and U19023 (N_19023,N_15448,N_17232);
or U19024 (N_19024,N_16744,N_15931);
nor U19025 (N_19025,N_15844,N_16494);
nor U19026 (N_19026,N_17108,N_15765);
nand U19027 (N_19027,N_15512,N_16051);
or U19028 (N_19028,N_15646,N_16263);
nor U19029 (N_19029,N_15383,N_17251);
and U19030 (N_19030,N_16363,N_16405);
or U19031 (N_19031,N_15372,N_15214);
or U19032 (N_19032,N_15277,N_17367);
or U19033 (N_19033,N_17453,N_15130);
nand U19034 (N_19034,N_16168,N_17077);
and U19035 (N_19035,N_15626,N_15357);
and U19036 (N_19036,N_16154,N_15809);
or U19037 (N_19037,N_16526,N_17226);
and U19038 (N_19038,N_16717,N_16391);
or U19039 (N_19039,N_17058,N_15769);
or U19040 (N_19040,N_16701,N_15689);
nor U19041 (N_19041,N_16470,N_16316);
or U19042 (N_19042,N_16152,N_16585);
nor U19043 (N_19043,N_17170,N_15027);
nand U19044 (N_19044,N_15158,N_17437);
nor U19045 (N_19045,N_16027,N_15896);
or U19046 (N_19046,N_17479,N_15711);
nand U19047 (N_19047,N_15203,N_17105);
or U19048 (N_19048,N_16388,N_15907);
and U19049 (N_19049,N_15521,N_16723);
nand U19050 (N_19050,N_17289,N_16702);
or U19051 (N_19051,N_15724,N_16872);
or U19052 (N_19052,N_16831,N_17132);
nand U19053 (N_19053,N_15717,N_17204);
or U19054 (N_19054,N_15693,N_16076);
nand U19055 (N_19055,N_17147,N_16106);
nand U19056 (N_19056,N_16854,N_15658);
or U19057 (N_19057,N_16202,N_16885);
or U19058 (N_19058,N_16490,N_15965);
xor U19059 (N_19059,N_16407,N_15703);
and U19060 (N_19060,N_17328,N_17274);
or U19061 (N_19061,N_17089,N_16387);
and U19062 (N_19062,N_15127,N_15957);
and U19063 (N_19063,N_15340,N_16052);
and U19064 (N_19064,N_16000,N_16228);
nor U19065 (N_19065,N_15624,N_16744);
and U19066 (N_19066,N_15880,N_16043);
or U19067 (N_19067,N_15249,N_15087);
or U19068 (N_19068,N_16116,N_17081);
nor U19069 (N_19069,N_16946,N_16020);
nor U19070 (N_19070,N_15432,N_15199);
nand U19071 (N_19071,N_16996,N_16311);
nor U19072 (N_19072,N_15583,N_17018);
nand U19073 (N_19073,N_15707,N_16333);
nand U19074 (N_19074,N_17255,N_15432);
or U19075 (N_19075,N_17225,N_15977);
nand U19076 (N_19076,N_16353,N_16120);
nor U19077 (N_19077,N_17219,N_16878);
and U19078 (N_19078,N_15226,N_15465);
or U19079 (N_19079,N_16100,N_16152);
or U19080 (N_19080,N_17152,N_16374);
nand U19081 (N_19081,N_15313,N_15409);
or U19082 (N_19082,N_15536,N_16976);
nand U19083 (N_19083,N_16119,N_15591);
and U19084 (N_19084,N_16026,N_16538);
and U19085 (N_19085,N_15815,N_16155);
or U19086 (N_19086,N_16235,N_15493);
or U19087 (N_19087,N_15991,N_16188);
or U19088 (N_19088,N_16505,N_15234);
nand U19089 (N_19089,N_17296,N_15057);
or U19090 (N_19090,N_16223,N_17334);
and U19091 (N_19091,N_16338,N_16280);
and U19092 (N_19092,N_16030,N_16488);
and U19093 (N_19093,N_17341,N_17219);
nand U19094 (N_19094,N_16152,N_15747);
nand U19095 (N_19095,N_15247,N_15927);
nor U19096 (N_19096,N_17200,N_16909);
nand U19097 (N_19097,N_15082,N_15395);
nand U19098 (N_19098,N_16567,N_17349);
nor U19099 (N_19099,N_15777,N_16183);
nor U19100 (N_19100,N_15576,N_15812);
nor U19101 (N_19101,N_17184,N_16093);
nand U19102 (N_19102,N_15570,N_16068);
nand U19103 (N_19103,N_17477,N_16019);
and U19104 (N_19104,N_16994,N_16148);
nor U19105 (N_19105,N_15626,N_15462);
nand U19106 (N_19106,N_15944,N_16647);
nor U19107 (N_19107,N_16824,N_15182);
xnor U19108 (N_19108,N_17340,N_16440);
and U19109 (N_19109,N_15761,N_17472);
or U19110 (N_19110,N_15572,N_15515);
nor U19111 (N_19111,N_15326,N_17292);
or U19112 (N_19112,N_16477,N_16830);
and U19113 (N_19113,N_16887,N_16589);
nand U19114 (N_19114,N_17160,N_15660);
nor U19115 (N_19115,N_16122,N_16455);
or U19116 (N_19116,N_16405,N_15795);
and U19117 (N_19117,N_15729,N_16608);
and U19118 (N_19118,N_17389,N_15102);
nand U19119 (N_19119,N_15073,N_15925);
and U19120 (N_19120,N_16058,N_15290);
nand U19121 (N_19121,N_16833,N_15504);
or U19122 (N_19122,N_17358,N_16851);
or U19123 (N_19123,N_15347,N_15476);
and U19124 (N_19124,N_16428,N_17259);
nand U19125 (N_19125,N_16138,N_15596);
nand U19126 (N_19126,N_15462,N_17388);
xor U19127 (N_19127,N_17109,N_16615);
nor U19128 (N_19128,N_16145,N_15391);
nor U19129 (N_19129,N_16546,N_16414);
nand U19130 (N_19130,N_15825,N_16350);
xnor U19131 (N_19131,N_15034,N_15531);
nand U19132 (N_19132,N_16203,N_17021);
and U19133 (N_19133,N_17238,N_15167);
xnor U19134 (N_19134,N_15552,N_16366);
and U19135 (N_19135,N_16368,N_16703);
nor U19136 (N_19136,N_15446,N_15113);
nand U19137 (N_19137,N_17090,N_17385);
or U19138 (N_19138,N_17152,N_15808);
or U19139 (N_19139,N_15124,N_15459);
nand U19140 (N_19140,N_17348,N_15858);
or U19141 (N_19141,N_16659,N_17488);
nor U19142 (N_19142,N_16393,N_16553);
nor U19143 (N_19143,N_16801,N_16349);
and U19144 (N_19144,N_17090,N_16154);
nor U19145 (N_19145,N_15945,N_16968);
nor U19146 (N_19146,N_15151,N_17114);
nor U19147 (N_19147,N_17119,N_15453);
or U19148 (N_19148,N_15162,N_15628);
and U19149 (N_19149,N_16201,N_16482);
and U19150 (N_19150,N_15157,N_17412);
nand U19151 (N_19151,N_16335,N_16580);
and U19152 (N_19152,N_15686,N_17496);
nand U19153 (N_19153,N_16539,N_16301);
nor U19154 (N_19154,N_16361,N_17429);
or U19155 (N_19155,N_15239,N_15821);
nand U19156 (N_19156,N_17458,N_17092);
and U19157 (N_19157,N_17096,N_16390);
nor U19158 (N_19158,N_15723,N_16514);
nor U19159 (N_19159,N_15707,N_16900);
and U19160 (N_19160,N_16460,N_15458);
or U19161 (N_19161,N_16483,N_16516);
or U19162 (N_19162,N_17224,N_16095);
or U19163 (N_19163,N_17445,N_16589);
xnor U19164 (N_19164,N_16983,N_15748);
nor U19165 (N_19165,N_15283,N_15105);
and U19166 (N_19166,N_15456,N_16828);
nor U19167 (N_19167,N_15436,N_16316);
nand U19168 (N_19168,N_17092,N_16086);
or U19169 (N_19169,N_17363,N_16072);
and U19170 (N_19170,N_16384,N_17090);
and U19171 (N_19171,N_17070,N_16872);
nand U19172 (N_19172,N_16863,N_17313);
and U19173 (N_19173,N_16354,N_16938);
and U19174 (N_19174,N_16039,N_15793);
nor U19175 (N_19175,N_16000,N_16398);
nand U19176 (N_19176,N_15789,N_15116);
and U19177 (N_19177,N_15619,N_17025);
nand U19178 (N_19178,N_17033,N_15284);
nor U19179 (N_19179,N_16689,N_16682);
nor U19180 (N_19180,N_16577,N_17021);
and U19181 (N_19181,N_15030,N_16803);
and U19182 (N_19182,N_15043,N_15286);
or U19183 (N_19183,N_16759,N_16972);
and U19184 (N_19184,N_15175,N_15987);
or U19185 (N_19185,N_15125,N_17159);
and U19186 (N_19186,N_16138,N_15896);
nand U19187 (N_19187,N_16734,N_15554);
nand U19188 (N_19188,N_15601,N_16631);
nand U19189 (N_19189,N_16814,N_16699);
nor U19190 (N_19190,N_15942,N_15893);
nor U19191 (N_19191,N_17485,N_15090);
and U19192 (N_19192,N_16487,N_16554);
nor U19193 (N_19193,N_17017,N_15919);
or U19194 (N_19194,N_16104,N_16286);
nand U19195 (N_19195,N_16643,N_16422);
and U19196 (N_19196,N_16625,N_17295);
nor U19197 (N_19197,N_15405,N_16404);
and U19198 (N_19198,N_17483,N_15396);
and U19199 (N_19199,N_16013,N_17218);
nand U19200 (N_19200,N_15983,N_15992);
nor U19201 (N_19201,N_16036,N_15191);
or U19202 (N_19202,N_16186,N_16514);
and U19203 (N_19203,N_15983,N_16544);
or U19204 (N_19204,N_16186,N_17415);
and U19205 (N_19205,N_16411,N_16016);
nor U19206 (N_19206,N_17411,N_17481);
or U19207 (N_19207,N_16741,N_15810);
and U19208 (N_19208,N_16963,N_16355);
or U19209 (N_19209,N_16376,N_17229);
nor U19210 (N_19210,N_17343,N_15662);
nand U19211 (N_19211,N_15893,N_15569);
nor U19212 (N_19212,N_15115,N_16271);
nor U19213 (N_19213,N_16151,N_16577);
nor U19214 (N_19214,N_16713,N_15005);
and U19215 (N_19215,N_17204,N_15011);
and U19216 (N_19216,N_16506,N_15680);
nor U19217 (N_19217,N_15979,N_16482);
or U19218 (N_19218,N_16442,N_17177);
nor U19219 (N_19219,N_16484,N_17187);
nor U19220 (N_19220,N_16616,N_15300);
nor U19221 (N_19221,N_15143,N_16478);
or U19222 (N_19222,N_16943,N_16198);
and U19223 (N_19223,N_16682,N_15912);
nor U19224 (N_19224,N_16162,N_16570);
xnor U19225 (N_19225,N_16056,N_17368);
or U19226 (N_19226,N_16446,N_17348);
nor U19227 (N_19227,N_16690,N_16251);
nand U19228 (N_19228,N_16894,N_17233);
nand U19229 (N_19229,N_15665,N_16040);
and U19230 (N_19230,N_16393,N_15505);
nor U19231 (N_19231,N_15365,N_17226);
nand U19232 (N_19232,N_15713,N_16531);
and U19233 (N_19233,N_16899,N_17424);
or U19234 (N_19234,N_16260,N_16395);
nor U19235 (N_19235,N_17370,N_15360);
nor U19236 (N_19236,N_15447,N_17107);
nand U19237 (N_19237,N_15532,N_17272);
nor U19238 (N_19238,N_15396,N_17025);
or U19239 (N_19239,N_17381,N_15203);
nor U19240 (N_19240,N_17442,N_16489);
nand U19241 (N_19241,N_15494,N_17233);
or U19242 (N_19242,N_16787,N_17053);
nor U19243 (N_19243,N_17037,N_16634);
nor U19244 (N_19244,N_17412,N_15364);
nor U19245 (N_19245,N_16184,N_15091);
nand U19246 (N_19246,N_16211,N_15602);
and U19247 (N_19247,N_15858,N_16163);
and U19248 (N_19248,N_16520,N_17172);
and U19249 (N_19249,N_15767,N_16230);
nor U19250 (N_19250,N_16937,N_16678);
nor U19251 (N_19251,N_16816,N_16529);
xor U19252 (N_19252,N_17430,N_17010);
nor U19253 (N_19253,N_17408,N_17321);
nor U19254 (N_19254,N_15977,N_16246);
nor U19255 (N_19255,N_15731,N_17023);
or U19256 (N_19256,N_15004,N_15479);
or U19257 (N_19257,N_15973,N_15207);
nor U19258 (N_19258,N_15628,N_15724);
and U19259 (N_19259,N_16098,N_15380);
nand U19260 (N_19260,N_17378,N_16863);
nor U19261 (N_19261,N_17256,N_15535);
and U19262 (N_19262,N_16938,N_15924);
nor U19263 (N_19263,N_15646,N_16140);
or U19264 (N_19264,N_16830,N_15444);
nand U19265 (N_19265,N_15157,N_15164);
xnor U19266 (N_19266,N_15312,N_16687);
nand U19267 (N_19267,N_16206,N_16524);
nor U19268 (N_19268,N_17330,N_16791);
or U19269 (N_19269,N_16558,N_16579);
nor U19270 (N_19270,N_17317,N_16674);
nor U19271 (N_19271,N_16546,N_17023);
and U19272 (N_19272,N_17372,N_15073);
and U19273 (N_19273,N_16330,N_17222);
nor U19274 (N_19274,N_17398,N_16028);
or U19275 (N_19275,N_17182,N_16263);
or U19276 (N_19276,N_15174,N_16451);
nor U19277 (N_19277,N_15735,N_17121);
and U19278 (N_19278,N_15201,N_15662);
or U19279 (N_19279,N_15881,N_17096);
nor U19280 (N_19280,N_17126,N_17262);
and U19281 (N_19281,N_15937,N_16937);
or U19282 (N_19282,N_16353,N_15222);
nor U19283 (N_19283,N_16707,N_16986);
nand U19284 (N_19284,N_16371,N_15747);
nand U19285 (N_19285,N_17439,N_17283);
nor U19286 (N_19286,N_15366,N_15006);
and U19287 (N_19287,N_15753,N_16963);
or U19288 (N_19288,N_16568,N_15894);
or U19289 (N_19289,N_15091,N_15157);
and U19290 (N_19290,N_15734,N_17113);
and U19291 (N_19291,N_16561,N_15587);
and U19292 (N_19292,N_15302,N_15670);
or U19293 (N_19293,N_15277,N_16974);
nand U19294 (N_19294,N_15833,N_16111);
nor U19295 (N_19295,N_17107,N_16734);
nor U19296 (N_19296,N_15445,N_16434);
or U19297 (N_19297,N_17305,N_16332);
nor U19298 (N_19298,N_15977,N_16669);
nand U19299 (N_19299,N_17068,N_16210);
and U19300 (N_19300,N_16930,N_15295);
or U19301 (N_19301,N_16795,N_16408);
nand U19302 (N_19302,N_16371,N_15226);
nand U19303 (N_19303,N_16070,N_15228);
or U19304 (N_19304,N_15193,N_16598);
nand U19305 (N_19305,N_15311,N_15985);
nor U19306 (N_19306,N_16778,N_15846);
nor U19307 (N_19307,N_16747,N_16329);
and U19308 (N_19308,N_16381,N_17360);
nand U19309 (N_19309,N_15544,N_16477);
or U19310 (N_19310,N_15494,N_17133);
and U19311 (N_19311,N_16579,N_15521);
or U19312 (N_19312,N_15496,N_16362);
nand U19313 (N_19313,N_16750,N_17185);
and U19314 (N_19314,N_15798,N_16901);
nand U19315 (N_19315,N_16310,N_17046);
nand U19316 (N_19316,N_15769,N_15919);
nand U19317 (N_19317,N_16097,N_15102);
nand U19318 (N_19318,N_15647,N_16721);
or U19319 (N_19319,N_17150,N_17346);
nand U19320 (N_19320,N_16610,N_16956);
and U19321 (N_19321,N_16196,N_17157);
nor U19322 (N_19322,N_16932,N_15948);
or U19323 (N_19323,N_16486,N_15282);
nand U19324 (N_19324,N_15146,N_15045);
and U19325 (N_19325,N_15926,N_15172);
and U19326 (N_19326,N_15676,N_16799);
or U19327 (N_19327,N_16548,N_17350);
nor U19328 (N_19328,N_16553,N_16866);
or U19329 (N_19329,N_16846,N_17174);
nor U19330 (N_19330,N_15708,N_16293);
or U19331 (N_19331,N_16102,N_16904);
and U19332 (N_19332,N_15090,N_16748);
and U19333 (N_19333,N_15186,N_15285);
nor U19334 (N_19334,N_15668,N_15976);
or U19335 (N_19335,N_15822,N_15356);
nand U19336 (N_19336,N_15558,N_16602);
nor U19337 (N_19337,N_15342,N_17269);
nand U19338 (N_19338,N_15034,N_15760);
nand U19339 (N_19339,N_15156,N_15332);
nand U19340 (N_19340,N_16417,N_15823);
nand U19341 (N_19341,N_15162,N_16120);
and U19342 (N_19342,N_16779,N_15492);
and U19343 (N_19343,N_16194,N_17378);
and U19344 (N_19344,N_17107,N_17332);
or U19345 (N_19345,N_17341,N_15964);
or U19346 (N_19346,N_16848,N_17075);
nor U19347 (N_19347,N_17092,N_16886);
and U19348 (N_19348,N_15866,N_15224);
and U19349 (N_19349,N_16950,N_16922);
nor U19350 (N_19350,N_15491,N_15493);
xor U19351 (N_19351,N_16133,N_15653);
or U19352 (N_19352,N_17193,N_15927);
and U19353 (N_19353,N_16231,N_15883);
and U19354 (N_19354,N_17391,N_16129);
and U19355 (N_19355,N_16426,N_17398);
nor U19356 (N_19356,N_17163,N_15702);
nand U19357 (N_19357,N_16039,N_16853);
or U19358 (N_19358,N_15972,N_15131);
and U19359 (N_19359,N_15779,N_15609);
or U19360 (N_19360,N_16706,N_15544);
and U19361 (N_19361,N_15884,N_16676);
nor U19362 (N_19362,N_17449,N_17083);
nand U19363 (N_19363,N_16219,N_15695);
and U19364 (N_19364,N_17119,N_16902);
or U19365 (N_19365,N_15195,N_16545);
nand U19366 (N_19366,N_15427,N_15036);
nand U19367 (N_19367,N_16956,N_16262);
nand U19368 (N_19368,N_17219,N_15543);
and U19369 (N_19369,N_15402,N_15086);
nor U19370 (N_19370,N_17007,N_16661);
or U19371 (N_19371,N_15242,N_15360);
or U19372 (N_19372,N_16402,N_15612);
or U19373 (N_19373,N_15173,N_15729);
nor U19374 (N_19374,N_15297,N_15896);
or U19375 (N_19375,N_15724,N_16450);
and U19376 (N_19376,N_15612,N_16975);
or U19377 (N_19377,N_16821,N_17436);
or U19378 (N_19378,N_16619,N_15011);
and U19379 (N_19379,N_15967,N_15984);
nand U19380 (N_19380,N_15199,N_15437);
nand U19381 (N_19381,N_15222,N_15322);
and U19382 (N_19382,N_15268,N_16743);
and U19383 (N_19383,N_15675,N_16938);
nor U19384 (N_19384,N_15561,N_17036);
or U19385 (N_19385,N_15745,N_15973);
nand U19386 (N_19386,N_16452,N_16995);
or U19387 (N_19387,N_16355,N_16001);
nor U19388 (N_19388,N_16205,N_17494);
xor U19389 (N_19389,N_17173,N_17183);
and U19390 (N_19390,N_16036,N_16532);
nor U19391 (N_19391,N_16396,N_16135);
or U19392 (N_19392,N_16013,N_15291);
nor U19393 (N_19393,N_15723,N_16449);
nor U19394 (N_19394,N_16882,N_17095);
nor U19395 (N_19395,N_17188,N_17063);
nor U19396 (N_19396,N_15383,N_15744);
nand U19397 (N_19397,N_15963,N_16715);
nand U19398 (N_19398,N_15040,N_16942);
nor U19399 (N_19399,N_15056,N_16217);
or U19400 (N_19400,N_17068,N_17005);
or U19401 (N_19401,N_15496,N_15508);
nor U19402 (N_19402,N_16816,N_16430);
and U19403 (N_19403,N_17167,N_15544);
or U19404 (N_19404,N_16546,N_16617);
and U19405 (N_19405,N_16525,N_16477);
or U19406 (N_19406,N_16178,N_15262);
and U19407 (N_19407,N_16680,N_16248);
or U19408 (N_19408,N_16872,N_15101);
xnor U19409 (N_19409,N_15812,N_17433);
nand U19410 (N_19410,N_16902,N_15491);
or U19411 (N_19411,N_17232,N_15732);
or U19412 (N_19412,N_15489,N_16280);
nor U19413 (N_19413,N_16430,N_15400);
or U19414 (N_19414,N_15838,N_17024);
nor U19415 (N_19415,N_17285,N_15168);
or U19416 (N_19416,N_17149,N_17126);
nand U19417 (N_19417,N_16127,N_15634);
xor U19418 (N_19418,N_15321,N_15912);
nand U19419 (N_19419,N_15133,N_16320);
nand U19420 (N_19420,N_17353,N_16209);
and U19421 (N_19421,N_15752,N_15354);
nand U19422 (N_19422,N_15057,N_16277);
and U19423 (N_19423,N_16654,N_16512);
nand U19424 (N_19424,N_15795,N_15359);
nand U19425 (N_19425,N_15153,N_15023);
nand U19426 (N_19426,N_15311,N_15663);
or U19427 (N_19427,N_16218,N_16648);
nand U19428 (N_19428,N_15374,N_15702);
or U19429 (N_19429,N_16828,N_17218);
nand U19430 (N_19430,N_17401,N_15915);
and U19431 (N_19431,N_15018,N_17048);
or U19432 (N_19432,N_16761,N_16325);
nor U19433 (N_19433,N_15689,N_17012);
nand U19434 (N_19434,N_17230,N_16215);
and U19435 (N_19435,N_17104,N_15246);
and U19436 (N_19436,N_17071,N_16823);
nor U19437 (N_19437,N_15759,N_17477);
or U19438 (N_19438,N_15836,N_15056);
and U19439 (N_19439,N_17481,N_17198);
and U19440 (N_19440,N_17069,N_15172);
or U19441 (N_19441,N_16567,N_16353);
or U19442 (N_19442,N_16428,N_16476);
and U19443 (N_19443,N_16026,N_16182);
and U19444 (N_19444,N_17175,N_16717);
and U19445 (N_19445,N_15843,N_16689);
and U19446 (N_19446,N_16034,N_16728);
xnor U19447 (N_19447,N_16176,N_16748);
or U19448 (N_19448,N_16691,N_16139);
and U19449 (N_19449,N_15048,N_16839);
or U19450 (N_19450,N_15859,N_15437);
nand U19451 (N_19451,N_15053,N_16882);
nand U19452 (N_19452,N_16665,N_15195);
or U19453 (N_19453,N_16088,N_15500);
and U19454 (N_19454,N_15652,N_15960);
and U19455 (N_19455,N_15499,N_15011);
nand U19456 (N_19456,N_16888,N_15768);
and U19457 (N_19457,N_17053,N_17495);
xor U19458 (N_19458,N_15670,N_16473);
nor U19459 (N_19459,N_15435,N_15340);
or U19460 (N_19460,N_15650,N_15372);
nor U19461 (N_19461,N_16635,N_15974);
or U19462 (N_19462,N_15820,N_17328);
or U19463 (N_19463,N_17042,N_16891);
and U19464 (N_19464,N_16537,N_15249);
and U19465 (N_19465,N_17151,N_15622);
nand U19466 (N_19466,N_17498,N_16238);
nand U19467 (N_19467,N_15500,N_15324);
or U19468 (N_19468,N_16202,N_15429);
nand U19469 (N_19469,N_15022,N_16409);
or U19470 (N_19470,N_16141,N_15791);
nand U19471 (N_19471,N_16251,N_15026);
or U19472 (N_19472,N_17023,N_17008);
and U19473 (N_19473,N_17370,N_15461);
nand U19474 (N_19474,N_16724,N_15597);
or U19475 (N_19475,N_16823,N_15066);
or U19476 (N_19476,N_15353,N_15229);
nand U19477 (N_19477,N_15638,N_15210);
nand U19478 (N_19478,N_17342,N_16170);
and U19479 (N_19479,N_16479,N_16091);
nand U19480 (N_19480,N_15269,N_16435);
or U19481 (N_19481,N_16864,N_15328);
nand U19482 (N_19482,N_16875,N_16068);
or U19483 (N_19483,N_17429,N_16246);
and U19484 (N_19484,N_15092,N_16833);
nor U19485 (N_19485,N_17219,N_16929);
and U19486 (N_19486,N_16537,N_15585);
or U19487 (N_19487,N_16940,N_15653);
and U19488 (N_19488,N_17410,N_16022);
and U19489 (N_19489,N_15687,N_16943);
nand U19490 (N_19490,N_15599,N_16582);
and U19491 (N_19491,N_16433,N_15954);
and U19492 (N_19492,N_16329,N_16565);
nand U19493 (N_19493,N_15219,N_15523);
nor U19494 (N_19494,N_16288,N_17277);
nor U19495 (N_19495,N_15935,N_16442);
or U19496 (N_19496,N_15440,N_16615);
and U19497 (N_19497,N_15990,N_15832);
nor U19498 (N_19498,N_16631,N_16429);
nor U19499 (N_19499,N_16597,N_16801);
or U19500 (N_19500,N_16593,N_15098);
xor U19501 (N_19501,N_16943,N_17410);
nor U19502 (N_19502,N_16600,N_15372);
nor U19503 (N_19503,N_15208,N_17092);
and U19504 (N_19504,N_17417,N_15278);
nand U19505 (N_19505,N_15344,N_17182);
and U19506 (N_19506,N_15978,N_16865);
nand U19507 (N_19507,N_16700,N_15037);
nor U19508 (N_19508,N_16050,N_16154);
and U19509 (N_19509,N_15117,N_15577);
and U19510 (N_19510,N_16805,N_17164);
and U19511 (N_19511,N_17399,N_15317);
and U19512 (N_19512,N_16878,N_16556);
xnor U19513 (N_19513,N_16931,N_15091);
nor U19514 (N_19514,N_16987,N_16623);
or U19515 (N_19515,N_15200,N_17346);
or U19516 (N_19516,N_16850,N_15912);
and U19517 (N_19517,N_15379,N_17206);
nand U19518 (N_19518,N_17283,N_15071);
nor U19519 (N_19519,N_15595,N_16458);
and U19520 (N_19520,N_16165,N_17008);
xnor U19521 (N_19521,N_15286,N_16026);
and U19522 (N_19522,N_15674,N_16758);
nor U19523 (N_19523,N_16363,N_16812);
or U19524 (N_19524,N_15586,N_16907);
or U19525 (N_19525,N_16121,N_15571);
and U19526 (N_19526,N_17076,N_16995);
and U19527 (N_19527,N_16023,N_15520);
and U19528 (N_19528,N_15599,N_15980);
and U19529 (N_19529,N_16908,N_16823);
nor U19530 (N_19530,N_15504,N_15098);
and U19531 (N_19531,N_17192,N_15075);
or U19532 (N_19532,N_15466,N_15954);
nand U19533 (N_19533,N_15939,N_16917);
nand U19534 (N_19534,N_17360,N_16830);
nor U19535 (N_19535,N_17192,N_15001);
or U19536 (N_19536,N_15922,N_16232);
nor U19537 (N_19537,N_16603,N_16426);
or U19538 (N_19538,N_16713,N_16936);
or U19539 (N_19539,N_16817,N_15442);
nor U19540 (N_19540,N_16018,N_15052);
or U19541 (N_19541,N_16285,N_15398);
nand U19542 (N_19542,N_15974,N_16163);
or U19543 (N_19543,N_15225,N_15237);
or U19544 (N_19544,N_16693,N_15732);
or U19545 (N_19545,N_15796,N_15628);
and U19546 (N_19546,N_15590,N_17422);
or U19547 (N_19547,N_15264,N_15957);
nand U19548 (N_19548,N_16799,N_16826);
or U19549 (N_19549,N_16844,N_17107);
xor U19550 (N_19550,N_15072,N_15519);
nand U19551 (N_19551,N_16373,N_16395);
xnor U19552 (N_19552,N_15298,N_15080);
or U19553 (N_19553,N_15503,N_15622);
and U19554 (N_19554,N_16983,N_16781);
and U19555 (N_19555,N_15099,N_16749);
or U19556 (N_19556,N_16869,N_16330);
nand U19557 (N_19557,N_16168,N_16912);
and U19558 (N_19558,N_17356,N_17086);
nor U19559 (N_19559,N_16756,N_17306);
and U19560 (N_19560,N_15740,N_17445);
or U19561 (N_19561,N_16092,N_16417);
and U19562 (N_19562,N_16879,N_15788);
nand U19563 (N_19563,N_16096,N_16184);
nor U19564 (N_19564,N_16168,N_15502);
nand U19565 (N_19565,N_16912,N_15608);
and U19566 (N_19566,N_16066,N_15099);
nand U19567 (N_19567,N_15248,N_15771);
or U19568 (N_19568,N_16612,N_16680);
or U19569 (N_19569,N_15012,N_16126);
nor U19570 (N_19570,N_16902,N_16170);
nor U19571 (N_19571,N_17470,N_15218);
nand U19572 (N_19572,N_15061,N_16723);
and U19573 (N_19573,N_16138,N_17432);
nand U19574 (N_19574,N_15849,N_15468);
or U19575 (N_19575,N_15256,N_16596);
nor U19576 (N_19576,N_16220,N_15903);
nand U19577 (N_19577,N_16090,N_15378);
and U19578 (N_19578,N_16566,N_15047);
nand U19579 (N_19579,N_16822,N_16618);
and U19580 (N_19580,N_15401,N_15905);
and U19581 (N_19581,N_17157,N_15088);
nor U19582 (N_19582,N_16503,N_15615);
nand U19583 (N_19583,N_16752,N_17466);
nand U19584 (N_19584,N_15194,N_15169);
nand U19585 (N_19585,N_16713,N_16172);
or U19586 (N_19586,N_16288,N_16946);
and U19587 (N_19587,N_16493,N_15238);
xnor U19588 (N_19588,N_15238,N_15583);
xor U19589 (N_19589,N_17029,N_15172);
or U19590 (N_19590,N_15895,N_16382);
nor U19591 (N_19591,N_16254,N_16849);
or U19592 (N_19592,N_17251,N_17071);
or U19593 (N_19593,N_16159,N_17349);
nor U19594 (N_19594,N_15947,N_15145);
or U19595 (N_19595,N_15109,N_16771);
nand U19596 (N_19596,N_15751,N_15522);
and U19597 (N_19597,N_16401,N_15022);
nand U19598 (N_19598,N_15445,N_16715);
or U19599 (N_19599,N_15707,N_17132);
and U19600 (N_19600,N_17312,N_16413);
nand U19601 (N_19601,N_15848,N_15822);
nor U19602 (N_19602,N_17103,N_17466);
xnor U19603 (N_19603,N_15617,N_16354);
nand U19604 (N_19604,N_16090,N_16791);
and U19605 (N_19605,N_15529,N_15029);
or U19606 (N_19606,N_15648,N_15873);
nor U19607 (N_19607,N_17048,N_15329);
and U19608 (N_19608,N_16746,N_16084);
and U19609 (N_19609,N_15575,N_17207);
or U19610 (N_19610,N_17126,N_16674);
nor U19611 (N_19611,N_17348,N_16828);
or U19612 (N_19612,N_16772,N_15002);
nand U19613 (N_19613,N_16645,N_15732);
or U19614 (N_19614,N_15017,N_15725);
or U19615 (N_19615,N_16842,N_15027);
or U19616 (N_19616,N_16649,N_17008);
nor U19617 (N_19617,N_17474,N_16376);
and U19618 (N_19618,N_15174,N_17239);
nor U19619 (N_19619,N_17215,N_16397);
and U19620 (N_19620,N_17016,N_16695);
nor U19621 (N_19621,N_15735,N_17227);
nor U19622 (N_19622,N_15701,N_16382);
and U19623 (N_19623,N_15843,N_15133);
and U19624 (N_19624,N_15765,N_16053);
and U19625 (N_19625,N_17243,N_15745);
and U19626 (N_19626,N_15325,N_15504);
nand U19627 (N_19627,N_15323,N_15558);
nand U19628 (N_19628,N_16449,N_15966);
nand U19629 (N_19629,N_17483,N_16970);
and U19630 (N_19630,N_15228,N_17298);
and U19631 (N_19631,N_15375,N_15046);
xor U19632 (N_19632,N_17218,N_16436);
and U19633 (N_19633,N_15653,N_16219);
xor U19634 (N_19634,N_16294,N_16227);
nor U19635 (N_19635,N_16197,N_16750);
or U19636 (N_19636,N_16053,N_17247);
or U19637 (N_19637,N_15466,N_15732);
nand U19638 (N_19638,N_15493,N_16769);
nor U19639 (N_19639,N_17425,N_17402);
nand U19640 (N_19640,N_15969,N_15971);
and U19641 (N_19641,N_15283,N_15546);
and U19642 (N_19642,N_16738,N_15315);
nor U19643 (N_19643,N_15546,N_16314);
or U19644 (N_19644,N_17216,N_16592);
nor U19645 (N_19645,N_16905,N_15924);
or U19646 (N_19646,N_16583,N_16273);
nand U19647 (N_19647,N_17082,N_15662);
or U19648 (N_19648,N_16954,N_17140);
nand U19649 (N_19649,N_16981,N_15563);
nor U19650 (N_19650,N_15860,N_16848);
or U19651 (N_19651,N_15539,N_15738);
or U19652 (N_19652,N_16204,N_16908);
and U19653 (N_19653,N_16770,N_16463);
nor U19654 (N_19654,N_16918,N_17425);
or U19655 (N_19655,N_17040,N_16519);
and U19656 (N_19656,N_16151,N_15184);
or U19657 (N_19657,N_16733,N_15810);
nand U19658 (N_19658,N_16138,N_15060);
nor U19659 (N_19659,N_17345,N_15929);
and U19660 (N_19660,N_15722,N_16984);
nor U19661 (N_19661,N_16683,N_15320);
nand U19662 (N_19662,N_15075,N_16920);
and U19663 (N_19663,N_15755,N_16336);
nand U19664 (N_19664,N_16764,N_15534);
nor U19665 (N_19665,N_15923,N_15562);
or U19666 (N_19666,N_15255,N_16090);
nand U19667 (N_19667,N_15128,N_16953);
and U19668 (N_19668,N_15817,N_17135);
or U19669 (N_19669,N_17498,N_17410);
or U19670 (N_19670,N_16317,N_17199);
nand U19671 (N_19671,N_15901,N_17451);
nand U19672 (N_19672,N_15473,N_15529);
nor U19673 (N_19673,N_15309,N_15902);
and U19674 (N_19674,N_16617,N_16750);
nor U19675 (N_19675,N_16597,N_15030);
and U19676 (N_19676,N_16212,N_17481);
nand U19677 (N_19677,N_17096,N_15658);
and U19678 (N_19678,N_16138,N_15999);
and U19679 (N_19679,N_15975,N_17200);
or U19680 (N_19680,N_15334,N_16382);
nand U19681 (N_19681,N_16052,N_15777);
and U19682 (N_19682,N_15951,N_15314);
nor U19683 (N_19683,N_16442,N_16915);
nand U19684 (N_19684,N_15841,N_17245);
and U19685 (N_19685,N_17072,N_17031);
and U19686 (N_19686,N_17459,N_15618);
nor U19687 (N_19687,N_15417,N_15324);
nor U19688 (N_19688,N_16782,N_15751);
nor U19689 (N_19689,N_17495,N_16664);
nor U19690 (N_19690,N_17051,N_15366);
and U19691 (N_19691,N_15139,N_15870);
nor U19692 (N_19692,N_17168,N_16707);
nor U19693 (N_19693,N_17357,N_15573);
nand U19694 (N_19694,N_17151,N_15815);
and U19695 (N_19695,N_17111,N_15332);
and U19696 (N_19696,N_15281,N_16873);
or U19697 (N_19697,N_15984,N_17146);
nand U19698 (N_19698,N_17247,N_15913);
and U19699 (N_19699,N_15858,N_17291);
or U19700 (N_19700,N_16803,N_16394);
nor U19701 (N_19701,N_16240,N_16568);
nand U19702 (N_19702,N_16032,N_16460);
and U19703 (N_19703,N_15794,N_16917);
or U19704 (N_19704,N_16944,N_17307);
or U19705 (N_19705,N_15495,N_16120);
or U19706 (N_19706,N_15206,N_16534);
or U19707 (N_19707,N_17176,N_17203);
nand U19708 (N_19708,N_15774,N_16848);
and U19709 (N_19709,N_15558,N_15328);
nor U19710 (N_19710,N_17405,N_15806);
and U19711 (N_19711,N_16563,N_15411);
nor U19712 (N_19712,N_15837,N_15915);
nand U19713 (N_19713,N_15750,N_17018);
and U19714 (N_19714,N_16404,N_16011);
nor U19715 (N_19715,N_15843,N_16699);
nor U19716 (N_19716,N_15189,N_15062);
nand U19717 (N_19717,N_15717,N_15734);
nor U19718 (N_19718,N_16946,N_16947);
and U19719 (N_19719,N_16788,N_16792);
nor U19720 (N_19720,N_15367,N_16290);
or U19721 (N_19721,N_15840,N_17074);
or U19722 (N_19722,N_15478,N_15575);
nand U19723 (N_19723,N_15522,N_16733);
and U19724 (N_19724,N_16584,N_15850);
and U19725 (N_19725,N_17216,N_17167);
nand U19726 (N_19726,N_16227,N_15165);
or U19727 (N_19727,N_16183,N_15393);
nor U19728 (N_19728,N_16556,N_16809);
nor U19729 (N_19729,N_16992,N_16614);
or U19730 (N_19730,N_16661,N_17278);
xor U19731 (N_19731,N_17117,N_17455);
nand U19732 (N_19732,N_15248,N_15772);
and U19733 (N_19733,N_15008,N_15838);
nand U19734 (N_19734,N_16493,N_15637);
or U19735 (N_19735,N_16608,N_16166);
or U19736 (N_19736,N_15775,N_15205);
nand U19737 (N_19737,N_15941,N_15394);
and U19738 (N_19738,N_15281,N_17391);
nor U19739 (N_19739,N_16526,N_16922);
and U19740 (N_19740,N_15635,N_15880);
nand U19741 (N_19741,N_16178,N_15498);
nand U19742 (N_19742,N_16044,N_15066);
and U19743 (N_19743,N_15557,N_15197);
nand U19744 (N_19744,N_16075,N_15792);
nand U19745 (N_19745,N_15338,N_17164);
and U19746 (N_19746,N_16052,N_16698);
nor U19747 (N_19747,N_15383,N_15287);
or U19748 (N_19748,N_16690,N_15172);
nor U19749 (N_19749,N_16496,N_16499);
nand U19750 (N_19750,N_15703,N_15170);
nor U19751 (N_19751,N_16856,N_15001);
nor U19752 (N_19752,N_16922,N_15724);
or U19753 (N_19753,N_16571,N_17314);
nor U19754 (N_19754,N_17301,N_16727);
nor U19755 (N_19755,N_16497,N_17362);
xnor U19756 (N_19756,N_16093,N_15792);
nand U19757 (N_19757,N_16623,N_15446);
or U19758 (N_19758,N_16936,N_17347);
or U19759 (N_19759,N_15521,N_16778);
or U19760 (N_19760,N_15769,N_16082);
nor U19761 (N_19761,N_16950,N_17245);
and U19762 (N_19762,N_15646,N_15794);
nand U19763 (N_19763,N_15770,N_16984);
or U19764 (N_19764,N_15511,N_16304);
nand U19765 (N_19765,N_16022,N_16497);
and U19766 (N_19766,N_16567,N_15240);
nor U19767 (N_19767,N_15960,N_16629);
nor U19768 (N_19768,N_16837,N_15067);
or U19769 (N_19769,N_16115,N_16008);
and U19770 (N_19770,N_16819,N_16506);
nor U19771 (N_19771,N_15354,N_16381);
and U19772 (N_19772,N_16340,N_16124);
or U19773 (N_19773,N_15592,N_15148);
nand U19774 (N_19774,N_16993,N_15132);
and U19775 (N_19775,N_16175,N_15651);
or U19776 (N_19776,N_17343,N_15056);
nand U19777 (N_19777,N_15979,N_16373);
nor U19778 (N_19778,N_15665,N_15543);
and U19779 (N_19779,N_15109,N_15636);
nand U19780 (N_19780,N_15531,N_16085);
or U19781 (N_19781,N_17326,N_17314);
and U19782 (N_19782,N_15664,N_17282);
nor U19783 (N_19783,N_15935,N_17123);
and U19784 (N_19784,N_17380,N_15626);
nor U19785 (N_19785,N_15993,N_15551);
nand U19786 (N_19786,N_15587,N_16368);
xnor U19787 (N_19787,N_15132,N_15946);
xnor U19788 (N_19788,N_15844,N_15813);
and U19789 (N_19789,N_17149,N_16099);
or U19790 (N_19790,N_17043,N_17012);
or U19791 (N_19791,N_15256,N_16435);
nand U19792 (N_19792,N_15984,N_16906);
nor U19793 (N_19793,N_16347,N_15729);
nand U19794 (N_19794,N_15614,N_16979);
nand U19795 (N_19795,N_15980,N_16761);
nor U19796 (N_19796,N_15720,N_16175);
nor U19797 (N_19797,N_16282,N_15784);
and U19798 (N_19798,N_15461,N_16594);
nor U19799 (N_19799,N_16068,N_17232);
nand U19800 (N_19800,N_17453,N_16602);
nor U19801 (N_19801,N_15642,N_16197);
and U19802 (N_19802,N_17488,N_16291);
xnor U19803 (N_19803,N_17489,N_16246);
nand U19804 (N_19804,N_17361,N_15713);
nor U19805 (N_19805,N_16098,N_16371);
nor U19806 (N_19806,N_16474,N_16715);
and U19807 (N_19807,N_15750,N_15170);
and U19808 (N_19808,N_16249,N_17426);
and U19809 (N_19809,N_16951,N_16865);
or U19810 (N_19810,N_15369,N_15401);
xor U19811 (N_19811,N_16553,N_16271);
nor U19812 (N_19812,N_17118,N_16429);
xnor U19813 (N_19813,N_15661,N_15167);
nor U19814 (N_19814,N_16240,N_17431);
nand U19815 (N_19815,N_17395,N_15209);
xnor U19816 (N_19816,N_16300,N_17445);
nand U19817 (N_19817,N_17122,N_15222);
and U19818 (N_19818,N_17493,N_16474);
or U19819 (N_19819,N_16589,N_16827);
nand U19820 (N_19820,N_17168,N_15424);
nand U19821 (N_19821,N_16703,N_16633);
and U19822 (N_19822,N_17473,N_16716);
and U19823 (N_19823,N_15105,N_15684);
nor U19824 (N_19824,N_16699,N_17072);
nand U19825 (N_19825,N_15963,N_17353);
and U19826 (N_19826,N_16234,N_16310);
nor U19827 (N_19827,N_16217,N_16963);
nor U19828 (N_19828,N_16464,N_16200);
and U19829 (N_19829,N_15390,N_15200);
or U19830 (N_19830,N_15741,N_16159);
nand U19831 (N_19831,N_15707,N_15126);
nand U19832 (N_19832,N_16646,N_15151);
nand U19833 (N_19833,N_16120,N_15948);
or U19834 (N_19834,N_15346,N_15352);
or U19835 (N_19835,N_16114,N_15503);
or U19836 (N_19836,N_16595,N_16084);
and U19837 (N_19837,N_15503,N_15012);
or U19838 (N_19838,N_16793,N_16191);
and U19839 (N_19839,N_16006,N_15124);
or U19840 (N_19840,N_15117,N_16582);
nor U19841 (N_19841,N_16764,N_17252);
nor U19842 (N_19842,N_16351,N_16811);
or U19843 (N_19843,N_16203,N_17267);
nor U19844 (N_19844,N_16822,N_17085);
and U19845 (N_19845,N_15611,N_15391);
or U19846 (N_19846,N_15315,N_15376);
or U19847 (N_19847,N_16561,N_17369);
nor U19848 (N_19848,N_15733,N_16254);
nor U19849 (N_19849,N_16230,N_17118);
xor U19850 (N_19850,N_15514,N_16262);
nor U19851 (N_19851,N_16256,N_15998);
or U19852 (N_19852,N_16906,N_16887);
xnor U19853 (N_19853,N_17263,N_15007);
or U19854 (N_19854,N_16742,N_15618);
or U19855 (N_19855,N_15196,N_15010);
and U19856 (N_19856,N_16870,N_15647);
nor U19857 (N_19857,N_16363,N_15510);
or U19858 (N_19858,N_17007,N_17048);
and U19859 (N_19859,N_15931,N_16902);
and U19860 (N_19860,N_17483,N_16509);
nor U19861 (N_19861,N_16370,N_15267);
nand U19862 (N_19862,N_16064,N_16132);
xor U19863 (N_19863,N_17146,N_15617);
nand U19864 (N_19864,N_15621,N_16320);
or U19865 (N_19865,N_16138,N_15311);
nor U19866 (N_19866,N_17097,N_16383);
nor U19867 (N_19867,N_15026,N_15587);
or U19868 (N_19868,N_16693,N_15325);
nor U19869 (N_19869,N_15640,N_16613);
and U19870 (N_19870,N_15139,N_17452);
nand U19871 (N_19871,N_15758,N_16178);
nor U19872 (N_19872,N_17297,N_17105);
nand U19873 (N_19873,N_16298,N_16866);
and U19874 (N_19874,N_16991,N_15605);
nor U19875 (N_19875,N_15774,N_17415);
nand U19876 (N_19876,N_16872,N_17273);
or U19877 (N_19877,N_16682,N_15016);
and U19878 (N_19878,N_16424,N_16084);
nor U19879 (N_19879,N_16430,N_16095);
and U19880 (N_19880,N_15429,N_17487);
and U19881 (N_19881,N_15434,N_16482);
nor U19882 (N_19882,N_15581,N_17371);
nor U19883 (N_19883,N_16329,N_15323);
nor U19884 (N_19884,N_16698,N_16001);
nor U19885 (N_19885,N_15366,N_16097);
nor U19886 (N_19886,N_16131,N_16368);
or U19887 (N_19887,N_16033,N_15184);
nand U19888 (N_19888,N_16942,N_15932);
and U19889 (N_19889,N_15339,N_16309);
nand U19890 (N_19890,N_15463,N_15028);
or U19891 (N_19891,N_16754,N_16285);
nand U19892 (N_19892,N_15858,N_16522);
or U19893 (N_19893,N_15728,N_15903);
or U19894 (N_19894,N_16945,N_15302);
and U19895 (N_19895,N_15309,N_15954);
and U19896 (N_19896,N_15137,N_16253);
xor U19897 (N_19897,N_15641,N_16491);
nand U19898 (N_19898,N_16656,N_16417);
nand U19899 (N_19899,N_15435,N_17426);
and U19900 (N_19900,N_17064,N_15110);
and U19901 (N_19901,N_17093,N_16500);
nor U19902 (N_19902,N_15163,N_16774);
and U19903 (N_19903,N_17393,N_16083);
nand U19904 (N_19904,N_16645,N_15353);
nand U19905 (N_19905,N_16964,N_15815);
nand U19906 (N_19906,N_16632,N_16749);
nand U19907 (N_19907,N_16408,N_16009);
nand U19908 (N_19908,N_16868,N_17365);
nand U19909 (N_19909,N_17475,N_16291);
nand U19910 (N_19910,N_15879,N_16886);
or U19911 (N_19911,N_15881,N_16186);
and U19912 (N_19912,N_17306,N_16838);
and U19913 (N_19913,N_16905,N_17190);
nor U19914 (N_19914,N_16328,N_15739);
nand U19915 (N_19915,N_16430,N_15858);
nor U19916 (N_19916,N_16596,N_15062);
nand U19917 (N_19917,N_15204,N_15040);
or U19918 (N_19918,N_15935,N_17159);
nand U19919 (N_19919,N_17285,N_15173);
and U19920 (N_19920,N_16464,N_15538);
nand U19921 (N_19921,N_15567,N_17189);
or U19922 (N_19922,N_15146,N_15220);
nand U19923 (N_19923,N_15355,N_17286);
or U19924 (N_19924,N_17377,N_17093);
and U19925 (N_19925,N_15994,N_16439);
nor U19926 (N_19926,N_15831,N_15543);
and U19927 (N_19927,N_16196,N_16151);
nand U19928 (N_19928,N_16693,N_16745);
or U19929 (N_19929,N_15051,N_16336);
nor U19930 (N_19930,N_15630,N_15365);
nand U19931 (N_19931,N_17011,N_15905);
nor U19932 (N_19932,N_15744,N_15834);
nand U19933 (N_19933,N_16549,N_16570);
and U19934 (N_19934,N_15219,N_15565);
nand U19935 (N_19935,N_16315,N_15251);
or U19936 (N_19936,N_17086,N_17045);
nand U19937 (N_19937,N_15610,N_15047);
nand U19938 (N_19938,N_16635,N_17026);
nand U19939 (N_19939,N_16676,N_15922);
and U19940 (N_19940,N_17317,N_16205);
nand U19941 (N_19941,N_17419,N_15529);
nor U19942 (N_19942,N_16567,N_16994);
nand U19943 (N_19943,N_16832,N_16823);
or U19944 (N_19944,N_16258,N_16486);
nand U19945 (N_19945,N_16005,N_16645);
and U19946 (N_19946,N_16982,N_17229);
and U19947 (N_19947,N_16672,N_17096);
or U19948 (N_19948,N_17345,N_15090);
nand U19949 (N_19949,N_16990,N_15052);
and U19950 (N_19950,N_15454,N_15075);
nor U19951 (N_19951,N_16950,N_16925);
nand U19952 (N_19952,N_15599,N_16071);
nand U19953 (N_19953,N_17349,N_17051);
nor U19954 (N_19954,N_15871,N_15510);
nand U19955 (N_19955,N_15355,N_16786);
nor U19956 (N_19956,N_15761,N_16808);
nand U19957 (N_19957,N_15405,N_16451);
and U19958 (N_19958,N_16698,N_15489);
and U19959 (N_19959,N_17459,N_17367);
nand U19960 (N_19960,N_15993,N_16930);
nand U19961 (N_19961,N_16651,N_16928);
and U19962 (N_19962,N_17229,N_17388);
or U19963 (N_19963,N_15175,N_17405);
or U19964 (N_19964,N_15045,N_15996);
nor U19965 (N_19965,N_15305,N_16033);
nand U19966 (N_19966,N_15474,N_16003);
nor U19967 (N_19967,N_17163,N_17372);
nor U19968 (N_19968,N_15129,N_17008);
nand U19969 (N_19969,N_15941,N_15143);
nand U19970 (N_19970,N_15324,N_16917);
nand U19971 (N_19971,N_16623,N_16056);
and U19972 (N_19972,N_16145,N_16490);
and U19973 (N_19973,N_16074,N_16380);
nand U19974 (N_19974,N_16732,N_16454);
nand U19975 (N_19975,N_16163,N_15262);
and U19976 (N_19976,N_16218,N_17356);
or U19977 (N_19977,N_16430,N_15736);
and U19978 (N_19978,N_16186,N_16051);
nor U19979 (N_19979,N_16244,N_17297);
and U19980 (N_19980,N_15872,N_15885);
or U19981 (N_19981,N_17125,N_15916);
and U19982 (N_19982,N_16754,N_16011);
nand U19983 (N_19983,N_17055,N_15546);
nand U19984 (N_19984,N_15094,N_15026);
nand U19985 (N_19985,N_17377,N_16912);
or U19986 (N_19986,N_16674,N_15388);
nand U19987 (N_19987,N_15833,N_15417);
and U19988 (N_19988,N_16334,N_15321);
nor U19989 (N_19989,N_16133,N_17142);
and U19990 (N_19990,N_15422,N_16929);
or U19991 (N_19991,N_15801,N_15833);
or U19992 (N_19992,N_16506,N_16877);
or U19993 (N_19993,N_16077,N_16444);
nand U19994 (N_19994,N_16284,N_15603);
and U19995 (N_19995,N_15919,N_17142);
or U19996 (N_19996,N_17093,N_16244);
or U19997 (N_19997,N_15892,N_16396);
nand U19998 (N_19998,N_15694,N_15041);
and U19999 (N_19999,N_15069,N_15347);
and U20000 (N_20000,N_18878,N_18317);
and U20001 (N_20001,N_17526,N_19589);
or U20002 (N_20002,N_18845,N_19489);
nor U20003 (N_20003,N_18902,N_17979);
and U20004 (N_20004,N_19182,N_18788);
or U20005 (N_20005,N_19167,N_18622);
and U20006 (N_20006,N_18526,N_18442);
nor U20007 (N_20007,N_19729,N_18178);
and U20008 (N_20008,N_19906,N_17511);
nand U20009 (N_20009,N_18393,N_18823);
or U20010 (N_20010,N_19429,N_18258);
xor U20011 (N_20011,N_19632,N_18942);
or U20012 (N_20012,N_18734,N_19653);
nand U20013 (N_20013,N_18696,N_19655);
nor U20014 (N_20014,N_17648,N_19318);
nor U20015 (N_20015,N_19007,N_17569);
or U20016 (N_20016,N_19576,N_19979);
nand U20017 (N_20017,N_18299,N_18282);
or U20018 (N_20018,N_17970,N_18781);
and U20019 (N_20019,N_19369,N_17907);
nor U20020 (N_20020,N_17661,N_19480);
nor U20021 (N_20021,N_18080,N_19800);
or U20022 (N_20022,N_17995,N_17660);
and U20023 (N_20023,N_19929,N_18738);
or U20024 (N_20024,N_19944,N_18870);
nand U20025 (N_20025,N_19794,N_19766);
or U20026 (N_20026,N_17739,N_18789);
nor U20027 (N_20027,N_18721,N_19949);
or U20028 (N_20028,N_19364,N_17726);
or U20029 (N_20029,N_17712,N_19791);
nor U20030 (N_20030,N_18311,N_17597);
nand U20031 (N_20031,N_19848,N_19270);
nor U20032 (N_20032,N_18855,N_19246);
nand U20033 (N_20033,N_19282,N_17690);
and U20034 (N_20034,N_19898,N_17884);
nand U20035 (N_20035,N_19073,N_17854);
nor U20036 (N_20036,N_17744,N_18445);
or U20037 (N_20037,N_17947,N_18645);
and U20038 (N_20038,N_19710,N_18495);
and U20039 (N_20039,N_19478,N_19520);
nand U20040 (N_20040,N_19169,N_17656);
and U20041 (N_20041,N_17719,N_17701);
nor U20042 (N_20042,N_18292,N_19432);
nand U20043 (N_20043,N_17883,N_18695);
nand U20044 (N_20044,N_17674,N_18469);
nand U20045 (N_20045,N_17785,N_18024);
nor U20046 (N_20046,N_19644,N_18903);
nand U20047 (N_20047,N_18560,N_18991);
nand U20048 (N_20048,N_18961,N_19560);
nand U20049 (N_20049,N_18180,N_19572);
nand U20050 (N_20050,N_17833,N_19612);
and U20051 (N_20051,N_18033,N_18540);
or U20052 (N_20052,N_18073,N_18882);
xor U20053 (N_20053,N_19047,N_19715);
nor U20054 (N_20054,N_19970,N_19911);
and U20055 (N_20055,N_19778,N_17797);
and U20056 (N_20056,N_18853,N_19306);
nor U20057 (N_20057,N_19419,N_17959);
or U20058 (N_20058,N_18348,N_18126);
or U20059 (N_20059,N_19583,N_19947);
nand U20060 (N_20060,N_19773,N_18133);
nor U20061 (N_20061,N_18280,N_18682);
nand U20062 (N_20062,N_18819,N_18822);
or U20063 (N_20063,N_19476,N_19411);
and U20064 (N_20064,N_19095,N_17826);
xor U20065 (N_20065,N_19856,N_19918);
nor U20066 (N_20066,N_18850,N_18636);
and U20067 (N_20067,N_18036,N_17531);
nand U20068 (N_20068,N_19550,N_18437);
xnor U20069 (N_20069,N_19004,N_18303);
xnor U20070 (N_20070,N_18312,N_18538);
nor U20071 (N_20071,N_17522,N_18605);
or U20072 (N_20072,N_19969,N_19814);
and U20073 (N_20073,N_18729,N_19209);
and U20074 (N_20074,N_18104,N_17796);
or U20075 (N_20075,N_19418,N_19499);
and U20076 (N_20076,N_17784,N_19392);
nor U20077 (N_20077,N_17651,N_17916);
or U20078 (N_20078,N_18202,N_17670);
xnor U20079 (N_20079,N_19397,N_19538);
nand U20080 (N_20080,N_17617,N_19734);
nor U20081 (N_20081,N_18749,N_19953);
or U20082 (N_20082,N_17850,N_19366);
nor U20083 (N_20083,N_17929,N_18171);
or U20084 (N_20084,N_17693,N_19924);
nand U20085 (N_20085,N_19978,N_18323);
nand U20086 (N_20086,N_19163,N_18228);
xor U20087 (N_20087,N_19333,N_19664);
and U20088 (N_20088,N_19446,N_19985);
nor U20089 (N_20089,N_19821,N_18219);
or U20090 (N_20090,N_19016,N_17698);
and U20091 (N_20091,N_19342,N_19581);
or U20092 (N_20092,N_19926,N_19110);
and U20093 (N_20093,N_19391,N_19622);
nor U20094 (N_20094,N_19822,N_18619);
nor U20095 (N_20095,N_17862,N_19260);
nand U20096 (N_20096,N_17702,N_17703);
and U20097 (N_20097,N_19574,N_18483);
nand U20098 (N_20098,N_18458,N_18575);
nor U20099 (N_20099,N_19762,N_18857);
xor U20100 (N_20100,N_18044,N_18586);
or U20101 (N_20101,N_18324,N_17583);
and U20102 (N_20102,N_17587,N_18816);
and U20103 (N_20103,N_18487,N_18426);
nand U20104 (N_20104,N_19460,N_19836);
nor U20105 (N_20105,N_18994,N_18322);
or U20106 (N_20106,N_18745,N_19373);
nand U20107 (N_20107,N_19009,N_19332);
nor U20108 (N_20108,N_19740,N_18593);
or U20109 (N_20109,N_17776,N_18234);
nand U20110 (N_20110,N_17538,N_18807);
or U20111 (N_20111,N_19151,N_19337);
xnor U20112 (N_20112,N_18862,N_19890);
nand U20113 (N_20113,N_19784,N_18003);
nor U20114 (N_20114,N_18680,N_18809);
nand U20115 (N_20115,N_19871,N_19928);
nor U20116 (N_20116,N_18337,N_18446);
nor U20117 (N_20117,N_18800,N_18380);
nand U20118 (N_20118,N_19950,N_19630);
or U20119 (N_20119,N_19227,N_18955);
and U20120 (N_20120,N_19229,N_19505);
and U20121 (N_20121,N_18818,N_18772);
nand U20122 (N_20122,N_19138,N_17541);
nor U20123 (N_20123,N_18149,N_18410);
nor U20124 (N_20124,N_18517,N_18632);
nand U20125 (N_20125,N_19586,N_17876);
nand U20126 (N_20126,N_19995,N_19295);
or U20127 (N_20127,N_18563,N_18906);
nand U20128 (N_20128,N_19634,N_19936);
nand U20129 (N_20129,N_17766,N_19679);
nor U20130 (N_20130,N_18198,N_17891);
and U20131 (N_20131,N_18471,N_19485);
nor U20132 (N_20132,N_18327,N_19345);
and U20133 (N_20133,N_17954,N_18933);
nand U20134 (N_20134,N_19475,N_17681);
or U20135 (N_20135,N_18021,N_17837);
nand U20136 (N_20136,N_18924,N_17594);
and U20137 (N_20137,N_18806,N_18112);
or U20138 (N_20138,N_18093,N_19412);
nor U20139 (N_20139,N_18865,N_18753);
nand U20140 (N_20140,N_17643,N_17798);
nor U20141 (N_20141,N_19416,N_18060);
and U20142 (N_20142,N_17634,N_19566);
and U20143 (N_20143,N_18795,N_19874);
nand U20144 (N_20144,N_18515,N_18043);
nand U20145 (N_20145,N_19355,N_18839);
and U20146 (N_20146,N_18325,N_18866);
nor U20147 (N_20147,N_19241,N_18009);
nor U20148 (N_20148,N_18555,N_19087);
nand U20149 (N_20149,N_18901,N_18278);
and U20150 (N_20150,N_18764,N_19951);
and U20151 (N_20151,N_19452,N_19415);
nand U20152 (N_20152,N_18728,N_19435);
or U20153 (N_20153,N_18860,N_19931);
and U20154 (N_20154,N_18177,N_19696);
or U20155 (N_20155,N_18685,N_18836);
nor U20156 (N_20156,N_19107,N_18372);
or U20157 (N_20157,N_17586,N_19385);
xor U20158 (N_20158,N_18637,N_19608);
or U20159 (N_20159,N_18191,N_19902);
nand U20160 (N_20160,N_18627,N_19286);
and U20161 (N_20161,N_19602,N_19512);
nor U20162 (N_20162,N_18068,N_17655);
xor U20163 (N_20163,N_18107,N_18368);
nor U20164 (N_20164,N_18123,N_18136);
nand U20165 (N_20165,N_19739,N_17711);
nor U20166 (N_20166,N_19495,N_17662);
or U20167 (N_20167,N_19123,N_19968);
xor U20168 (N_20168,N_19530,N_17782);
nand U20169 (N_20169,N_19780,N_17788);
nand U20170 (N_20170,N_18001,N_19935);
nand U20171 (N_20171,N_18099,N_18079);
nor U20172 (N_20172,N_18186,N_18694);
and U20173 (N_20173,N_19401,N_17637);
or U20174 (N_20174,N_17957,N_17536);
nand U20175 (N_20175,N_18403,N_18692);
and U20176 (N_20176,N_19468,N_19775);
xnor U20177 (N_20177,N_18193,N_19940);
nor U20178 (N_20178,N_19642,N_18381);
nand U20179 (N_20179,N_18121,N_19381);
nand U20180 (N_20180,N_18306,N_17912);
nor U20181 (N_20181,N_19591,N_18333);
nand U20182 (N_20182,N_18146,N_18194);
nor U20183 (N_20183,N_18424,N_17834);
nand U20184 (N_20184,N_17967,N_17517);
xnor U20185 (N_20185,N_18584,N_19291);
and U20186 (N_20186,N_19109,N_18022);
nor U20187 (N_20187,N_19382,N_17896);
nand U20188 (N_20188,N_18506,N_17806);
nand U20189 (N_20189,N_19496,N_17956);
or U20190 (N_20190,N_18946,N_19298);
nand U20191 (N_20191,N_18720,N_19633);
and U20192 (N_20192,N_19544,N_18565);
nor U20193 (N_20193,N_17500,N_18274);
or U20194 (N_20194,N_17611,N_19129);
nand U20195 (N_20195,N_19052,N_19610);
nand U20196 (N_20196,N_18607,N_17828);
or U20197 (N_20197,N_19920,N_17989);
or U20198 (N_20198,N_18250,N_19863);
and U20199 (N_20199,N_19671,N_18926);
or U20200 (N_20200,N_19541,N_19252);
and U20201 (N_20201,N_19540,N_18940);
nor U20202 (N_20202,N_19697,N_18522);
and U20203 (N_20203,N_19135,N_19343);
or U20204 (N_20204,N_19666,N_19214);
and U20205 (N_20205,N_19470,N_19159);
nor U20206 (N_20206,N_19916,N_17734);
nand U20207 (N_20207,N_18799,N_18570);
nand U20208 (N_20208,N_18915,N_19050);
nand U20209 (N_20209,N_18630,N_17742);
nand U20210 (N_20210,N_17999,N_19623);
xor U20211 (N_20211,N_17976,N_17625);
nand U20212 (N_20212,N_19684,N_18081);
or U20213 (N_20213,N_19414,N_17938);
nand U20214 (N_20214,N_19807,N_19854);
and U20215 (N_20215,N_19508,N_17966);
or U20216 (N_20216,N_17584,N_17801);
nor U20217 (N_20217,N_17808,N_18864);
and U20218 (N_20218,N_19249,N_19267);
or U20219 (N_20219,N_19706,N_19562);
or U20220 (N_20220,N_18389,N_18392);
nor U20221 (N_20221,N_18331,N_17875);
or U20222 (N_20222,N_19243,N_18415);
and U20223 (N_20223,N_17772,N_18967);
nor U20224 (N_20224,N_17607,N_19082);
and U20225 (N_20225,N_19059,N_19744);
nor U20226 (N_20226,N_19939,N_19558);
nor U20227 (N_20227,N_17992,N_18597);
and U20228 (N_20228,N_18651,N_17764);
nand U20229 (N_20229,N_18817,N_17514);
and U20230 (N_20230,N_18263,N_18617);
or U20231 (N_20231,N_19165,N_18827);
nor U20232 (N_20232,N_18711,N_19036);
nor U20233 (N_20233,N_18837,N_18201);
nand U20234 (N_20234,N_18830,N_19510);
and U20235 (N_20235,N_18993,N_18014);
nand U20236 (N_20236,N_18660,N_19093);
or U20237 (N_20237,N_18141,N_19064);
nand U20238 (N_20238,N_18291,N_19804);
nor U20239 (N_20239,N_18652,N_18122);
nor U20240 (N_20240,N_19635,N_18908);
nor U20241 (N_20241,N_19074,N_19353);
nand U20242 (N_20242,N_19000,N_17932);
and U20243 (N_20243,N_18105,N_18737);
or U20244 (N_20244,N_19772,N_18985);
nor U20245 (N_20245,N_17921,N_17926);
and U20246 (N_20246,N_19893,N_18992);
nor U20247 (N_20247,N_19402,N_18190);
nor U20248 (N_20248,N_18616,N_18971);
xor U20249 (N_20249,N_19309,N_17578);
nor U20250 (N_20250,N_18640,N_19996);
nand U20251 (N_20251,N_17818,N_18918);
nand U20252 (N_20252,N_18321,N_18074);
and U20253 (N_20253,N_18248,N_18066);
nand U20254 (N_20254,N_18083,N_19732);
or U20255 (N_20255,N_17952,N_17839);
and U20256 (N_20256,N_19799,N_17774);
nand U20257 (N_20257,N_19359,N_18673);
or U20258 (N_20258,N_18497,N_19043);
or U20259 (N_20259,N_18042,N_19617);
and U20260 (N_20260,N_17532,N_19801);
xnor U20261 (N_20261,N_19197,N_18863);
nor U20262 (N_20262,N_19207,N_18037);
and U20263 (N_20263,N_19737,N_19975);
or U20264 (N_20264,N_18166,N_18599);
or U20265 (N_20265,N_18551,N_19676);
nand U20266 (N_20266,N_19105,N_18480);
nand U20267 (N_20267,N_19181,N_18422);
nor U20268 (N_20268,N_17773,N_18628);
nor U20269 (N_20269,N_18242,N_18513);
nand U20270 (N_20270,N_18345,N_17802);
and U20271 (N_20271,N_17778,N_19603);
nand U20272 (N_20272,N_19261,N_18384);
nand U20273 (N_20273,N_18569,N_17548);
or U20274 (N_20274,N_19824,N_18999);
nand U20275 (N_20275,N_18132,N_17853);
or U20276 (N_20276,N_19024,N_19075);
and U20277 (N_20277,N_18953,N_18527);
nor U20278 (N_20278,N_18189,N_19033);
or U20279 (N_20279,N_18731,N_19462);
nor U20280 (N_20280,N_19021,N_19280);
and U20281 (N_20281,N_18479,N_19628);
or U20282 (N_20282,N_17629,N_19500);
nor U20283 (N_20283,N_19058,N_18106);
nand U20284 (N_20284,N_17867,N_18664);
or U20285 (N_20285,N_17955,N_18834);
and U20286 (N_20286,N_19239,N_19713);
or U20287 (N_20287,N_19092,N_19730);
or U20288 (N_20288,N_19805,N_18709);
and U20289 (N_20289,N_19128,N_18048);
and U20290 (N_20290,N_17910,N_19048);
nand U20291 (N_20291,N_18979,N_19061);
nor U20292 (N_20292,N_18742,N_18061);
or U20293 (N_20293,N_18511,N_19872);
nand U20294 (N_20294,N_19113,N_19673);
nor U20295 (N_20295,N_19474,N_18168);
nand U20296 (N_20296,N_17993,N_18359);
and U20297 (N_20297,N_17664,N_19952);
or U20298 (N_20298,N_18935,N_19756);
or U20299 (N_20299,N_19810,N_19437);
nor U20300 (N_20300,N_17771,N_18440);
and U20301 (N_20301,N_17515,N_19442);
and U20302 (N_20302,N_19451,N_19857);
and U20303 (N_20303,N_18741,N_17871);
nand U20304 (N_20304,N_19494,N_18591);
and U20305 (N_20305,N_17622,N_18402);
nand U20306 (N_20306,N_19677,N_18606);
and U20307 (N_20307,N_18766,N_19904);
or U20308 (N_20308,N_18377,N_18046);
or U20309 (N_20309,N_19643,N_18580);
nor U20310 (N_20310,N_18466,N_18539);
and U20311 (N_20311,N_18172,N_18397);
and U20312 (N_20312,N_17874,N_18116);
and U20313 (N_20313,N_19425,N_18984);
or U20314 (N_20314,N_17628,N_19257);
nand U20315 (N_20315,N_18922,N_19307);
nand U20316 (N_20316,N_18065,N_18473);
and U20317 (N_20317,N_19681,N_19124);
and U20318 (N_20318,N_19652,N_19690);
nor U20319 (N_20319,N_19549,N_19972);
or U20320 (N_20320,N_19153,N_19980);
nor U20321 (N_20321,N_18269,N_19912);
and U20322 (N_20322,N_19795,N_18100);
and U20323 (N_20323,N_19830,N_18451);
nand U20324 (N_20324,N_18039,N_18018);
xor U20325 (N_20325,N_18447,N_19639);
nor U20326 (N_20326,N_17675,N_19284);
and U20327 (N_20327,N_19709,N_19482);
nand U20328 (N_20328,N_18117,N_18681);
nand U20329 (N_20329,N_17816,N_18925);
xnor U20330 (N_20330,N_19627,N_18416);
nor U20331 (N_20331,N_18686,N_18874);
nor U20332 (N_20332,N_18157,N_18297);
or U20333 (N_20333,N_18574,N_17668);
and U20334 (N_20334,N_18050,N_19090);
and U20335 (N_20335,N_19362,N_17881);
and U20336 (N_20336,N_18948,N_19176);
or U20337 (N_20337,N_19321,N_19860);
nand U20338 (N_20338,N_17756,N_19121);
or U20339 (N_20339,N_19380,N_19365);
xor U20340 (N_20340,N_19741,N_18502);
or U20341 (N_20341,N_17878,N_17699);
nor U20342 (N_20342,N_18842,N_17501);
and U20343 (N_20343,N_19759,N_18236);
nand U20344 (N_20344,N_18786,N_19704);
and U20345 (N_20345,N_19917,N_19449);
or U20346 (N_20346,N_19777,N_18778);
nor U20347 (N_20347,N_19955,N_18241);
or U20348 (N_20348,N_19198,N_17555);
nand U20349 (N_20349,N_18887,N_19273);
nand U20350 (N_20350,N_19014,N_17987);
or U20351 (N_20351,N_18740,N_18719);
nor U20352 (N_20352,N_18572,N_17786);
nand U20353 (N_20353,N_19873,N_19185);
and U20354 (N_20354,N_19316,N_18670);
or U20355 (N_20355,N_18071,N_19726);
and U20356 (N_20356,N_19934,N_18464);
nand U20357 (N_20357,N_19665,N_19897);
or U20358 (N_20358,N_17688,N_18541);
and U20359 (N_20359,N_18247,N_19290);
nor U20360 (N_20360,N_19427,N_17557);
nor U20361 (N_20361,N_19305,N_17749);
and U20362 (N_20362,N_19196,N_18406);
nand U20363 (N_20363,N_18429,N_19594);
nand U20364 (N_20364,N_19883,N_18218);
nand U20365 (N_20365,N_17812,N_19311);
and U20366 (N_20366,N_18880,N_17525);
and U20367 (N_20367,N_18152,N_17646);
or U20368 (N_20368,N_19098,N_18746);
and U20369 (N_20369,N_17975,N_19817);
or U20370 (N_20370,N_18420,N_18970);
nand U20371 (N_20371,N_17509,N_17942);
nor U20372 (N_20372,N_19650,N_19228);
nand U20373 (N_20373,N_19711,N_18943);
nand U20374 (N_20374,N_19884,N_18956);
or U20375 (N_20375,N_19636,N_18491);
or U20376 (N_20376,N_18160,N_18944);
nand U20377 (N_20377,N_18006,N_19276);
or U20378 (N_20378,N_17746,N_17879);
nand U20379 (N_20379,N_19625,N_17813);
or U20380 (N_20380,N_18910,N_19324);
xnor U20381 (N_20381,N_18715,N_18373);
nand U20382 (N_20382,N_18963,N_18108);
nor U20383 (N_20383,N_19275,N_17895);
nor U20384 (N_20384,N_19742,N_18702);
nand U20385 (N_20385,N_17996,N_19720);
or U20386 (N_20386,N_19348,N_18820);
and U20387 (N_20387,N_17520,N_17519);
and U20388 (N_20388,N_18723,N_18260);
nor U20389 (N_20389,N_18101,N_19640);
and U20390 (N_20390,N_17633,N_18978);
and U20391 (N_20391,N_19111,N_18335);
nand U20392 (N_20392,N_19503,N_19932);
nor U20393 (N_20393,N_17614,N_19188);
and U20394 (N_20394,N_19738,N_19956);
or U20395 (N_20395,N_18120,N_18400);
nand U20396 (N_20396,N_19587,N_18804);
nand U20397 (N_20397,N_19647,N_17645);
nor U20398 (N_20398,N_17750,N_18796);
and U20399 (N_20399,N_19685,N_18868);
and U20400 (N_20400,N_19907,N_19954);
nand U20401 (N_20401,N_19065,N_18275);
nand U20402 (N_20402,N_18679,N_17620);
and U20403 (N_20403,N_17504,N_18298);
nand U20404 (N_20404,N_19289,N_19667);
nand U20405 (N_20405,N_19447,N_19040);
or U20406 (N_20406,N_17965,N_17725);
and U20407 (N_20407,N_19086,N_17799);
or U20408 (N_20408,N_18129,N_19913);
xnor U20409 (N_20409,N_19915,N_19278);
and U20410 (N_20410,N_18162,N_19565);
nand U20411 (N_20411,N_18609,N_18712);
or U20412 (N_20412,N_17603,N_18932);
nand U20413 (N_20413,N_19695,N_17585);
nand U20414 (N_20414,N_19546,N_18595);
nand U20415 (N_20415,N_18928,N_19094);
nand U20416 (N_20416,N_18034,N_17575);
nand U20417 (N_20417,N_19104,N_17872);
and U20418 (N_20418,N_19259,N_18383);
or U20419 (N_20419,N_18545,N_18343);
or U20420 (N_20420,N_18618,N_17819);
nand U20421 (N_20421,N_18875,N_18936);
nor U20422 (N_20422,N_18750,N_19858);
and U20423 (N_20423,N_17728,N_19263);
or U20424 (N_20424,N_18854,N_18654);
nand U20425 (N_20425,N_19945,N_19049);
nand U20426 (N_20426,N_18078,N_19477);
and U20427 (N_20427,N_17757,N_18784);
and U20428 (N_20428,N_17971,N_19998);
or U20429 (N_20429,N_17759,N_19455);
or U20430 (N_20430,N_18253,N_18873);
nor U20431 (N_20431,N_19112,N_19967);
and U20432 (N_20432,N_18119,N_18030);
nor U20433 (N_20433,N_18604,N_19658);
nand U20434 (N_20434,N_19422,N_19702);
nor U20435 (N_20435,N_19819,N_19567);
and U20436 (N_20436,N_19548,N_19146);
or U20437 (N_20437,N_19728,N_19714);
or U20438 (N_20438,N_19517,N_19948);
xnor U20439 (N_20439,N_19247,N_18843);
nand U20440 (N_20440,N_18347,N_18156);
and U20441 (N_20441,N_19689,N_19611);
or U20442 (N_20442,N_18649,N_18205);
nor U20443 (N_20443,N_18592,N_18139);
nor U20444 (N_20444,N_17697,N_18677);
or U20445 (N_20445,N_19662,N_19601);
and U20446 (N_20446,N_18427,N_17745);
nand U20447 (N_20447,N_17880,N_19708);
and U20448 (N_20448,N_17551,N_18460);
and U20449 (N_20449,N_17753,N_18448);
or U20450 (N_20450,N_19178,N_18366);
and U20451 (N_20451,N_18722,N_19042);
or U20452 (N_20452,N_19269,N_19585);
nor U20453 (N_20453,N_19347,N_19308);
and U20454 (N_20454,N_19329,N_18828);
nor U20455 (N_20455,N_19674,N_19125);
nor U20456 (N_20456,N_17600,N_18055);
or U20457 (N_20457,N_19352,N_19896);
and U20458 (N_20458,N_17936,N_19498);
nand U20459 (N_20459,N_19903,N_18672);
and U20460 (N_20460,N_19668,N_18264);
nand U20461 (N_20461,N_17825,N_18792);
and U20462 (N_20462,N_19604,N_18354);
nor U20463 (N_20463,N_18656,N_19331);
or U20464 (N_20464,N_18304,N_19158);
nor U20465 (N_20465,N_19497,N_17723);
nand U20466 (N_20466,N_19160,N_17564);
nand U20467 (N_20467,N_18173,N_18755);
nand U20468 (N_20468,N_19879,N_18023);
and U20469 (N_20469,N_18613,N_19629);
nand U20470 (N_20470,N_19162,N_17527);
nor U20471 (N_20471,N_17811,N_17832);
and U20472 (N_20472,N_19002,N_18376);
and U20473 (N_20473,N_18035,N_19439);
and U20474 (N_20474,N_18611,N_18052);
nand U20475 (N_20475,N_18476,N_18884);
nor U20476 (N_20476,N_19106,N_19006);
or U20477 (N_20477,N_19204,N_19147);
nand U20478 (N_20478,N_18714,N_17866);
and U20479 (N_20479,N_17842,N_18077);
nor U20480 (N_20480,N_18414,N_19783);
nand U20481 (N_20481,N_19490,N_17972);
nand U20482 (N_20482,N_19578,N_19139);
nor U20483 (N_20483,N_18351,N_18891);
or U20484 (N_20484,N_17893,N_18045);
nand U20485 (N_20485,N_18493,N_19861);
nor U20486 (N_20486,N_19254,N_19592);
and U20487 (N_20487,N_18667,N_17964);
nor U20488 (N_20488,N_18535,N_18239);
or U20489 (N_20489,N_19976,N_18374);
or U20490 (N_20490,N_19618,N_17821);
nor U20491 (N_20491,N_19683,N_18998);
and U20492 (N_20492,N_17980,N_19989);
nand U20493 (N_20493,N_17596,N_17632);
or U20494 (N_20494,N_19885,N_18224);
and U20495 (N_20495,N_18000,N_19943);
nor U20496 (N_20496,N_19149,N_19410);
and U20497 (N_20497,N_18259,N_18968);
nand U20498 (N_20498,N_19234,N_17565);
or U20499 (N_20499,N_17649,N_18508);
nand U20500 (N_20500,N_18161,N_17706);
xor U20501 (N_20501,N_18548,N_19472);
nand U20502 (N_20502,N_19843,N_17793);
or U20503 (N_20503,N_19641,N_18209);
nor U20504 (N_20504,N_19459,N_18254);
xor U20505 (N_20505,N_17969,N_18113);
or U20506 (N_20506,N_19692,N_17767);
and U20507 (N_20507,N_19750,N_19045);
nor U20508 (N_20508,N_19761,N_19649);
xnor U20509 (N_20509,N_19370,N_17765);
and U20510 (N_20510,N_18520,N_18338);
or U20511 (N_20511,N_18724,N_19274);
or U20512 (N_20512,N_18898,N_17847);
nor U20513 (N_20513,N_19509,N_19637);
nand U20514 (N_20514,N_19440,N_19743);
xnor U20515 (N_20515,N_19217,N_18705);
nor U20516 (N_20516,N_19256,N_19789);
or U20517 (N_20517,N_18307,N_18642);
nand U20518 (N_20518,N_19097,N_18921);
nand U20519 (N_20519,N_17761,N_19757);
nand U20520 (N_20520,N_18096,N_18004);
nor U20521 (N_20521,N_19070,N_19765);
xor U20522 (N_20522,N_18401,N_19698);
or U20523 (N_20523,N_19573,N_18069);
or U20524 (N_20524,N_19925,N_18641);
or U20525 (N_20525,N_18124,N_17736);
or U20526 (N_20526,N_17677,N_18255);
nor U20527 (N_20527,N_18610,N_18477);
and U20528 (N_20528,N_18815,N_19582);
nand U20529 (N_20529,N_18752,N_18431);
and U20530 (N_20530,N_19463,N_19032);
and U20531 (N_20531,N_18761,N_18150);
or U20532 (N_20532,N_18929,N_19598);
and U20533 (N_20533,N_18029,N_18313);
and U20534 (N_20534,N_18683,N_18265);
nor U20535 (N_20535,N_17923,N_17868);
nor U20536 (N_20536,N_18895,N_19764);
nor U20537 (N_20537,N_18031,N_17521);
nand U20538 (N_20538,N_18273,N_18339);
nor U20539 (N_20539,N_17908,N_19233);
and U20540 (N_20540,N_18589,N_19682);
nand U20541 (N_20541,N_18067,N_18760);
nor U20542 (N_20542,N_17904,N_18399);
or U20543 (N_20543,N_17823,N_18983);
and U20544 (N_20544,N_18185,N_17567);
nor U20545 (N_20545,N_18251,N_17982);
nand U20546 (N_20546,N_19336,N_19561);
or U20547 (N_20547,N_18841,N_19892);
nand U20548 (N_20548,N_19317,N_17556);
or U20549 (N_20549,N_17542,N_18739);
nor U20550 (N_20550,N_17574,N_18960);
nor U20551 (N_20551,N_19659,N_19071);
or U20552 (N_20552,N_18756,N_18986);
or U20553 (N_20553,N_19143,N_19971);
and U20554 (N_20554,N_19068,N_19615);
nand U20555 (N_20555,N_17679,N_18110);
nand U20556 (N_20556,N_19938,N_18294);
or U20557 (N_20557,N_17704,N_18409);
nor U20558 (N_20558,N_18371,N_19326);
xor U20559 (N_20559,N_19235,N_19406);
nand U20560 (N_20560,N_17820,N_19688);
nor U20561 (N_20561,N_18892,N_17870);
xor U20562 (N_20562,N_17859,N_19213);
nor U20563 (N_20563,N_18899,N_18631);
and U20564 (N_20564,N_18614,N_18832);
or U20565 (N_20565,N_19251,N_18147);
and U20566 (N_20566,N_19304,N_18125);
nor U20567 (N_20567,N_19754,N_18690);
nor U20568 (N_20568,N_18010,N_18302);
and U20569 (N_20569,N_19686,N_17713);
or U20570 (N_20570,N_17800,N_18142);
and U20571 (N_20571,N_19579,N_19262);
nand U20572 (N_20572,N_17809,N_17845);
or U20573 (N_20573,N_17815,N_18434);
or U20574 (N_20574,N_17835,N_18310);
xor U20575 (N_20575,N_19005,N_17903);
nand U20576 (N_20576,N_19029,N_18470);
nand U20577 (N_20577,N_17619,N_19524);
nand U20578 (N_20578,N_19046,N_17692);
nand U20579 (N_20579,N_18957,N_17873);
and U20580 (N_20580,N_17732,N_18987);
or U20581 (N_20581,N_18578,N_19467);
and U20582 (N_20582,N_19088,N_18798);
nand U20583 (N_20583,N_18840,N_17570);
nand U20584 (N_20584,N_19798,N_19914);
nand U20585 (N_20585,N_18379,N_19609);
nor U20586 (N_20586,N_17846,N_19961);
nand U20587 (N_20587,N_19175,N_17777);
or U20588 (N_20588,N_17827,N_18566);
nor U20589 (N_20589,N_17865,N_19084);
nor U20590 (N_20590,N_18386,N_18883);
nor U20591 (N_20591,N_18767,N_19322);
or U20592 (N_20592,N_18015,N_17695);
nand U20593 (N_20593,N_18358,N_18296);
nand U20594 (N_20594,N_18747,N_18391);
nand U20595 (N_20595,N_19815,N_18553);
nor U20596 (N_20596,N_17986,N_18717);
nor U20597 (N_20597,N_17510,N_18430);
or U20598 (N_20598,N_18165,N_17804);
nand U20599 (N_20599,N_18408,N_19513);
nor U20600 (N_20600,N_18966,N_18188);
and U20601 (N_20601,N_19200,N_18964);
or U20602 (N_20602,N_19461,N_17707);
or U20603 (N_20603,N_19296,N_18954);
or U20604 (N_20604,N_18145,N_18047);
nand U20605 (N_20605,N_19779,N_18559);
nand U20606 (N_20606,N_19379,N_18349);
and U20607 (N_20607,N_18576,N_19923);
and U20608 (N_20608,N_19189,N_18858);
nand U20609 (N_20609,N_19648,N_18062);
nand U20610 (N_20610,N_17553,N_19448);
nand U20611 (N_20611,N_18546,N_18938);
or U20612 (N_20612,N_18320,N_18821);
or U20613 (N_20613,N_18183,N_18871);
nor U20614 (N_20614,N_19127,N_19958);
xor U20615 (N_20615,N_19657,N_18226);
or U20616 (N_20616,N_17779,N_17780);
nand U20617 (N_20617,N_18550,N_18780);
and U20618 (N_20618,N_18890,N_18759);
nand U20619 (N_20619,N_19186,N_18289);
nand U20620 (N_20620,N_18444,N_19875);
nor U20621 (N_20621,N_18962,N_18485);
nor U20622 (N_20622,N_19626,N_18256);
and U20623 (N_20623,N_17581,N_18221);
nor U20624 (N_20624,N_19137,N_18897);
nor U20625 (N_20625,N_19900,N_17807);
nand U20626 (N_20626,N_17927,N_18794);
and U20627 (N_20627,N_18465,N_17752);
or U20628 (N_20628,N_19551,N_19240);
and U20629 (N_20629,N_18245,N_17787);
nor U20630 (N_20630,N_18309,N_18653);
or U20631 (N_20631,N_19066,N_18669);
or U20632 (N_20632,N_19977,N_19941);
or U20633 (N_20633,N_18281,N_19763);
nor U20634 (N_20634,N_19526,N_17512);
nor U20635 (N_20635,N_17858,N_18529);
nor U20636 (N_20636,N_18418,N_19661);
nor U20637 (N_20637,N_19297,N_19533);
nor U20638 (N_20638,N_18571,N_19012);
and U20639 (N_20639,N_17943,N_19013);
nand U20640 (N_20640,N_19716,N_18064);
nand U20641 (N_20641,N_18284,N_19091);
nor U20642 (N_20642,N_17939,N_18852);
and U20643 (N_20643,N_19770,N_19384);
nand U20644 (N_20644,N_19041,N_19614);
nand U20645 (N_20645,N_18844,N_18230);
xnor U20646 (N_20646,N_18127,N_18644);
or U20647 (N_20647,N_19942,N_17963);
and U20648 (N_20648,N_18825,N_18730);
nor U20649 (N_20649,N_18225,N_18793);
nor U20650 (N_20650,N_18287,N_19563);
xor U20651 (N_20651,N_17940,N_18387);
nand U20652 (N_20652,N_19504,N_17691);
and U20653 (N_20653,N_19420,N_18361);
or U20654 (N_20654,N_19292,N_18494);
and U20655 (N_20655,N_17547,N_18328);
nor U20656 (N_20656,N_18646,N_19733);
and U20657 (N_20657,N_19266,N_18456);
nand U20658 (N_20658,N_18989,N_18534);
nor U20659 (N_20659,N_19215,N_19171);
nand U20660 (N_20660,N_19377,N_19067);
nand U20661 (N_20661,N_18148,N_19471);
xor U20662 (N_20662,N_19491,N_18474);
xnor U20663 (N_20663,N_19310,N_17685);
nand U20664 (N_20664,N_18097,N_19624);
nor U20665 (N_20665,N_19946,N_18638);
nand U20666 (N_20666,N_19901,N_19076);
and U20667 (N_20667,N_17922,N_17582);
nand U20668 (N_20668,N_18808,N_17897);
nand U20669 (N_20669,N_18937,N_19017);
nand U20670 (N_20670,N_19376,N_18095);
nor U20671 (N_20671,N_17981,N_17738);
or U20672 (N_20672,N_19554,N_17945);
nand U20673 (N_20673,N_18489,N_18102);
or U20674 (N_20674,N_19063,N_17941);
nor U20675 (N_20675,N_17885,N_17560);
and U20676 (N_20676,N_18557,N_17610);
nor U20677 (N_20677,N_19383,N_19027);
or U20678 (N_20678,N_19727,N_18626);
nand U20679 (N_20679,N_19010,N_17676);
and U20680 (N_20680,N_19545,N_19846);
or U20681 (N_20681,N_18463,N_18318);
or U20682 (N_20682,N_17731,N_19515);
nand U20683 (N_20683,N_18647,N_18342);
nand U20684 (N_20684,N_19523,N_18461);
nand U20685 (N_20685,N_18334,N_19431);
nor U20686 (N_20686,N_18507,N_17978);
nand U20687 (N_20687,N_19982,N_18192);
and U20688 (N_20688,N_19428,N_19096);
or U20689 (N_20689,N_19346,N_19271);
nor U20690 (N_20690,N_19521,N_18725);
and U20691 (N_20691,N_19785,N_19281);
xor U20692 (N_20692,N_17805,N_19486);
nand U20693 (N_20693,N_18057,N_19908);
and U20694 (N_20694,N_18472,N_19487);
nand U20695 (N_20695,N_18965,N_19535);
nand U20696 (N_20696,N_19192,N_18011);
xor U20697 (N_20697,N_19358,N_18509);
nand U20698 (N_20698,N_19368,N_19287);
or U20699 (N_20699,N_18777,N_18143);
and U20700 (N_20700,N_19421,N_17863);
xnor U20701 (N_20701,N_18635,N_19223);
nor U20702 (N_20702,N_17949,N_18917);
nand U20703 (N_20703,N_18814,N_18212);
nand U20704 (N_20704,N_18735,N_18811);
or U20705 (N_20705,N_18439,N_19144);
nand U20706 (N_20706,N_18633,N_17540);
nor U20707 (N_20707,N_18666,N_18662);
nor U20708 (N_20708,N_18733,N_19864);
or U20709 (N_20709,N_17506,N_19388);
or U20710 (N_20710,N_19119,N_19747);
nand U20711 (N_20711,N_18988,N_19851);
or U20712 (N_20712,N_18886,N_18305);
or U20713 (N_20713,N_19787,N_17915);
nand U20714 (N_20714,N_19011,N_17831);
and U20715 (N_20715,N_18267,N_18927);
nand U20716 (N_20716,N_19195,N_18582);
nand U20717 (N_20717,N_19319,N_18718);
nand U20718 (N_20718,N_18092,N_19580);
nor U20719 (N_20719,N_19170,N_17758);
or U20720 (N_20720,N_17624,N_19537);
nor U20721 (N_20721,N_19122,N_19020);
and U20722 (N_20722,N_18314,N_17605);
or U20723 (N_20723,N_18475,N_18027);
nand U20724 (N_20724,N_18385,N_17928);
nand U20725 (N_20725,N_19596,N_17654);
nand U20726 (N_20726,N_17869,N_19660);
nand U20727 (N_20727,N_19371,N_19760);
and U20728 (N_20728,N_19132,N_19393);
nor U20729 (N_20729,N_18982,N_18390);
nor U20730 (N_20730,N_18041,N_18486);
nand U20731 (N_20731,N_19751,N_18931);
and U20732 (N_20732,N_19719,N_17855);
and U20733 (N_20733,N_18261,N_19748);
xor U20734 (N_20734,N_19210,N_18196);
nor U20735 (N_20735,N_18249,N_17638);
nand U20736 (N_20736,N_17687,N_18791);
nor U20737 (N_20737,N_17672,N_18140);
nor U20738 (N_20738,N_18835,N_19823);
nand U20739 (N_20739,N_19080,N_19600);
or U20740 (N_20740,N_17968,N_18826);
or U20741 (N_20741,N_17546,N_19367);
or U20742 (N_20742,N_19838,N_17857);
xor U20743 (N_20743,N_19771,N_18594);
nor U20744 (N_20744,N_19378,N_19992);
or U20745 (N_20745,N_19469,N_18084);
nand U20746 (N_20746,N_19776,N_19361);
nor U20747 (N_20747,N_17639,N_19638);
or U20748 (N_20748,N_19868,N_18972);
nor U20749 (N_20749,N_19736,N_17905);
and U20750 (N_20750,N_18629,N_19363);
nand U20751 (N_20751,N_17877,N_19910);
or U20752 (N_20752,N_18634,N_19656);
nand U20753 (N_20753,N_17571,N_17573);
nand U20754 (N_20754,N_18623,N_18813);
or U20755 (N_20755,N_18697,N_18916);
nor U20756 (N_20756,N_18378,N_18639);
and U20757 (N_20757,N_19077,N_18369);
or U20758 (N_20758,N_18661,N_19960);
or U20759 (N_20759,N_17592,N_18829);
nor U20760 (N_20760,N_17890,N_18164);
nor U20761 (N_20761,N_18600,N_18977);
and U20762 (N_20762,N_18398,N_18950);
and U20763 (N_20763,N_18554,N_19831);
and U20764 (N_20764,N_19183,N_19283);
or U20765 (N_20765,N_19231,N_18181);
and U20766 (N_20766,N_19853,N_18668);
or U20767 (N_20767,N_19335,N_18271);
or U20768 (N_20768,N_19030,N_19328);
or U20769 (N_20769,N_18195,N_19180);
nand U20770 (N_20770,N_18128,N_19258);
nand U20771 (N_20771,N_19722,N_17836);
and U20772 (N_20772,N_18505,N_19115);
nand U20773 (N_20773,N_18382,N_18220);
and U20774 (N_20774,N_18558,N_19675);
nor U20775 (N_20775,N_19038,N_17899);
and U20776 (N_20776,N_17599,N_19407);
nand U20777 (N_20777,N_18433,N_17636);
and U20778 (N_20778,N_19405,N_19216);
and U20779 (N_20779,N_19882,N_19605);
or U20780 (N_20780,N_19465,N_18768);
nand U20781 (N_20781,N_18659,N_18848);
or U20782 (N_20782,N_18405,N_17843);
and U20783 (N_20783,N_17640,N_18969);
or U20784 (N_20784,N_19145,N_18785);
xnor U20785 (N_20785,N_17684,N_19404);
nand U20786 (N_20786,N_19792,N_17860);
or U20787 (N_20787,N_19268,N_18478);
nor U20788 (N_20788,N_18419,N_19037);
nand U20789 (N_20789,N_18707,N_18919);
and U20790 (N_20790,N_18501,N_19825);
xnor U20791 (N_20791,N_19226,N_19039);
nand U20792 (N_20792,N_18743,N_19360);
and U20793 (N_20793,N_19691,N_19015);
and U20794 (N_20794,N_17579,N_19616);
and U20795 (N_20795,N_18716,N_19441);
or U20796 (N_20796,N_19886,N_19990);
nand U20797 (N_20797,N_18336,N_18040);
or U20798 (N_20798,N_18163,N_17920);
nand U20799 (N_20799,N_19174,N_17563);
xor U20800 (N_20800,N_17630,N_19152);
nor U20801 (N_20801,N_17665,N_19248);
nor U20802 (N_20802,N_19678,N_18227);
or U20803 (N_20803,N_19157,N_19225);
or U20804 (N_20804,N_19288,N_18462);
or U20805 (N_20805,N_19493,N_18435);
or U20806 (N_20806,N_18939,N_17539);
and U20807 (N_20807,N_18665,N_19501);
nand U20808 (N_20808,N_18203,N_19072);
nor U20809 (N_20809,N_18547,N_19031);
nand U20810 (N_20810,N_18615,N_17516);
nand U20811 (N_20811,N_19705,N_18771);
nor U20812 (N_20812,N_17789,N_19255);
or U20813 (N_20813,N_18671,N_19481);
and U20814 (N_20814,N_18411,N_17840);
nand U20815 (N_20815,N_19054,N_18689);
nor U20816 (N_20816,N_18365,N_19502);
nand U20817 (N_20817,N_18199,N_19116);
or U20818 (N_20818,N_19909,N_18542);
nor U20819 (N_20819,N_17817,N_18240);
xnor U20820 (N_20820,N_17888,N_18360);
nand U20821 (N_20821,N_18959,N_18089);
nand U20822 (N_20822,N_18727,N_18070);
nand U20823 (N_20823,N_18776,N_19134);
and U20824 (N_20824,N_18115,N_18754);
nand U20825 (N_20825,N_18153,N_19142);
or U20826 (N_20826,N_18051,N_19542);
or U20827 (N_20827,N_17650,N_18293);
and U20828 (N_20828,N_17991,N_19140);
nand U20829 (N_20829,N_18454,N_18053);
nand U20830 (N_20830,N_18765,N_19511);
or U20831 (N_20831,N_19841,N_19398);
nor U20832 (N_20832,N_19962,N_19386);
nor U20833 (N_20833,N_17829,N_18769);
nor U20834 (N_20834,N_17741,N_18244);
nand U20835 (N_20835,N_19349,N_17958);
and U20836 (N_20836,N_18779,N_19927);
nand U20837 (N_20837,N_19236,N_19557);
and U20838 (N_20838,N_17566,N_17608);
or U20839 (N_20839,N_17626,N_18687);
or U20840 (N_20840,N_18367,N_18417);
nor U20841 (N_20841,N_17994,N_19651);
and U20842 (N_20842,N_19816,N_19456);
nor U20843 (N_20843,N_17534,N_18980);
nor U20844 (N_20844,N_17502,N_19905);
and U20845 (N_20845,N_17601,N_19774);
nor U20846 (N_20846,N_18663,N_18770);
and U20847 (N_20847,N_19786,N_19552);
nand U20848 (N_20848,N_17700,N_17984);
nand U20849 (N_20849,N_17589,N_18861);
and U20850 (N_20850,N_18757,N_19555);
or U20851 (N_20851,N_17644,N_18213);
or U20852 (N_20852,N_19937,N_19829);
nand U20853 (N_20853,N_19100,N_18658);
or U20854 (N_20854,N_18231,N_19529);
and U20855 (N_20855,N_18655,N_18118);
and U20856 (N_20856,N_19613,N_19922);
nand U20857 (N_20857,N_17591,N_19023);
nand U20858 (N_20858,N_18290,N_18496);
nand U20859 (N_20859,N_17559,N_18484);
and U20860 (N_20860,N_18974,N_17961);
or U20861 (N_20861,N_17983,N_18708);
and U20862 (N_20862,N_18889,N_19718);
and U20863 (N_20863,N_18130,N_19357);
nor U20864 (N_20864,N_19400,N_19987);
xnor U20865 (N_20865,N_18490,N_17545);
nand U20866 (N_20866,N_18790,N_18197);
or U20867 (N_20867,N_18233,N_18537);
or U20868 (N_20868,N_18976,N_19222);
and U20869 (N_20869,N_19194,N_17917);
nor U20870 (N_20870,N_18090,N_18773);
or U20871 (N_20871,N_17683,N_18453);
nor U20872 (N_20872,N_18905,N_18187);
nand U20873 (N_20873,N_18556,N_18941);
and U20874 (N_20874,N_19164,N_19325);
and U20875 (N_20875,N_19454,N_18002);
xor U20876 (N_20876,N_19444,N_19201);
nand U20877 (N_20877,N_18005,N_19434);
xor U20878 (N_20878,N_18363,N_18270);
and U20879 (N_20879,N_17769,N_18498);
nand U20880 (N_20880,N_19399,N_18344);
or U20881 (N_20881,N_19035,N_17529);
nand U20882 (N_20882,N_19458,N_19190);
xnor U20883 (N_20883,N_19735,N_18449);
or U20884 (N_20884,N_18923,N_19484);
nand U20885 (N_20885,N_19423,N_17659);
or U20886 (N_20886,N_18395,N_19809);
or U20887 (N_20887,N_18847,N_17708);
or U20888 (N_20888,N_17558,N_18025);
and U20889 (N_20889,N_17894,N_19599);
or U20890 (N_20890,N_19323,N_17990);
and U20891 (N_20891,N_18229,N_19062);
and U20892 (N_20892,N_19327,N_18549);
and U20893 (N_20893,N_19339,N_19842);
nor U20894 (N_20894,N_18235,N_18869);
nand U20895 (N_20895,N_17733,N_17621);
and U20896 (N_20896,N_18585,N_18996);
and U20897 (N_20897,N_18223,N_18518);
and U20898 (N_20898,N_18838,N_19208);
and U20899 (N_20899,N_19986,N_17814);
nor U20900 (N_20900,N_17852,N_19963);
or U20901 (N_20901,N_19506,N_18701);
or U20902 (N_20902,N_18763,N_19396);
xor U20903 (N_20903,N_17729,N_19717);
nor U20904 (N_20904,N_18020,N_18352);
nor U20905 (N_20905,N_19965,N_17618);
and U20906 (N_20906,N_18252,N_18500);
nor U20907 (N_20907,N_18579,N_19570);
nor U20908 (N_20908,N_17590,N_17948);
nand U20909 (N_20909,N_19790,N_18997);
or U20910 (N_20910,N_18608,N_19518);
nor U20911 (N_20911,N_18467,N_18438);
nand U20912 (N_20912,N_18782,N_19473);
nor U20913 (N_20913,N_17666,N_19237);
nor U20914 (N_20914,N_17730,N_18155);
nand U20915 (N_20915,N_19646,N_18407);
nand U20916 (N_20916,N_17861,N_18170);
xor U20917 (N_20917,N_19536,N_18425);
nand U20918 (N_20918,N_19085,N_18872);
nor U20919 (N_20919,N_19069,N_18017);
nand U20920 (N_20920,N_18762,N_17689);
nand U20921 (N_20921,N_18900,N_18098);
nand U20922 (N_20922,N_17606,N_18421);
or U20923 (N_20923,N_18214,N_18237);
nor U20924 (N_20924,N_18206,N_18443);
and U20925 (N_20925,N_18346,N_19746);
nor U20926 (N_20926,N_18357,N_19161);
or U20927 (N_20927,N_19507,N_19680);
nand U20928 (N_20928,N_19796,N_18488);
nand U20929 (N_20929,N_19571,N_18907);
nand U20930 (N_20930,N_19607,N_17657);
or U20931 (N_20931,N_19230,N_18920);
or U20932 (N_20932,N_19081,N_19788);
or U20933 (N_20933,N_17709,N_19001);
nand U20934 (N_20934,N_17507,N_19723);
nand U20935 (N_20935,N_17576,N_17530);
and U20936 (N_20936,N_19869,N_17505);
nand U20937 (N_20937,N_17513,N_19547);
and U20938 (N_20938,N_17663,N_19179);
and U20939 (N_20939,N_19919,N_18032);
nor U20940 (N_20940,N_19108,N_17935);
xor U20941 (N_20941,N_17886,N_18355);
or U20942 (N_20942,N_18945,N_17533);
nand U20943 (N_20943,N_18620,N_19781);
and U20944 (N_20944,N_19534,N_18810);
or U20945 (N_20945,N_19372,N_17720);
and U20946 (N_20946,N_19464,N_17783);
or U20947 (N_20947,N_18182,N_18054);
or U20948 (N_20948,N_19492,N_17844);
nand U20949 (N_20949,N_19118,N_18775);
nand U20950 (N_20950,N_18688,N_19219);
and U20951 (N_20951,N_17653,N_18262);
or U20952 (N_20952,N_19835,N_17715);
or U20953 (N_20953,N_18888,N_19301);
and U20954 (N_20954,N_19320,N_17930);
or U20955 (N_20955,N_19156,N_19584);
or U20956 (N_20956,N_18138,N_18482);
nand U20957 (N_20957,N_17792,N_18704);
nand U20958 (N_20958,N_18824,N_19862);
and U20959 (N_20959,N_18086,N_19350);
and U20960 (N_20960,N_19250,N_18362);
nor U20961 (N_20961,N_19700,N_18295);
and U20962 (N_20962,N_18643,N_17747);
nand U20963 (N_20963,N_17696,N_18896);
or U20964 (N_20964,N_18981,N_17528);
or U20965 (N_20965,N_19211,N_19876);
xnor U20966 (N_20966,N_17931,N_17951);
or U20967 (N_20967,N_17635,N_18876);
or U20968 (N_20968,N_19417,N_19619);
or U20969 (N_20969,N_18562,N_19859);
or U20970 (N_20970,N_18849,N_17748);
nor U20971 (N_20971,N_18169,N_17755);
or U20972 (N_20972,N_19394,N_19483);
nand U20973 (N_20973,N_19752,N_18200);
nor U20974 (N_20974,N_17669,N_18524);
and U20975 (N_20975,N_18912,N_17988);
or U20976 (N_20976,N_18783,N_17909);
or U20977 (N_20977,N_19528,N_18802);
nand U20978 (N_20978,N_19880,N_17568);
or U20979 (N_20979,N_19516,N_18038);
nor U20980 (N_20980,N_18436,N_18867);
nand U20981 (N_20981,N_19155,N_17751);
nand U20982 (N_20982,N_19395,N_18350);
or U20983 (N_20983,N_19212,N_19575);
or U20984 (N_20984,N_19532,N_19527);
and U20985 (N_20985,N_18603,N_18990);
or U20986 (N_20986,N_18648,N_19802);
or U20987 (N_20987,N_17544,N_17918);
nand U20988 (N_20988,N_17864,N_19811);
or U20989 (N_20989,N_18510,N_18457);
nand U20990 (N_20990,N_17641,N_18316);
or U20991 (N_20991,N_18413,N_19889);
and U20992 (N_20992,N_19855,N_18266);
nor U20993 (N_20993,N_17673,N_17727);
nand U20994 (N_20994,N_18441,N_19173);
xor U20995 (N_20995,N_19891,N_18774);
nor U20996 (N_20996,N_18450,N_19375);
and U20997 (N_20997,N_19438,N_18059);
nor U20998 (N_20998,N_17550,N_17623);
and U20999 (N_20999,N_19433,N_19564);
and U21000 (N_21000,N_17718,N_17710);
and U21001 (N_21001,N_19981,N_19930);
or U21002 (N_21002,N_19553,N_19621);
or U21003 (N_21003,N_17838,N_18913);
and U21004 (N_21004,N_18238,N_19450);
nand U21005 (N_21005,N_18693,N_18530);
nand U21006 (N_21006,N_17770,N_17856);
and U21007 (N_21007,N_18210,N_18277);
and U21008 (N_21008,N_19453,N_18216);
and U21009 (N_21009,N_18624,N_17790);
or U21010 (N_21010,N_19120,N_18134);
and U21011 (N_21011,N_17631,N_18703);
or U21012 (N_21012,N_18028,N_19356);
or U21013 (N_21013,N_17671,N_18257);
and U21014 (N_21014,N_19866,N_18222);
and U21015 (N_21015,N_19218,N_19531);
or U21016 (N_21016,N_18751,N_19539);
nand U21017 (N_21017,N_17602,N_17604);
nand U21018 (N_21018,N_18801,N_18678);
nor U21019 (N_21019,N_18019,N_19899);
nor U21020 (N_21020,N_19028,N_19199);
and U21021 (N_21021,N_19025,N_18951);
nand U21022 (N_21022,N_19895,N_19999);
nor U21023 (N_21023,N_19354,N_17760);
nor U21024 (N_21024,N_18521,N_18013);
nor U21025 (N_21025,N_18356,N_19293);
nor U21026 (N_21026,N_17775,N_18710);
and U21027 (N_21027,N_17658,N_18625);
and U21028 (N_21028,N_17503,N_17524);
nand U21029 (N_21029,N_18532,N_18388);
nand U21030 (N_21030,N_19313,N_19184);
nand U21031 (N_21031,N_19983,N_18706);
and U21032 (N_21032,N_18805,N_19403);
nor U21033 (N_21033,N_19820,N_17613);
nor U21034 (N_21034,N_18208,N_19285);
nor U21035 (N_21035,N_18833,N_19338);
nand U21036 (N_21036,N_18859,N_19136);
nand U21037 (N_21037,N_17721,N_19525);
and U21038 (N_21038,N_17810,N_19203);
nor U21039 (N_21039,N_19245,N_19154);
and U21040 (N_21040,N_19834,N_18076);
nor U21041 (N_21041,N_17882,N_19168);
and U21042 (N_21042,N_19753,N_19390);
and U21043 (N_21043,N_19008,N_19344);
nor U21044 (N_21044,N_17552,N_18300);
and U21045 (N_21045,N_18732,N_18621);
nand U21046 (N_21046,N_19221,N_19593);
nor U21047 (N_21047,N_19206,N_19959);
nand U21048 (N_21048,N_18958,N_18831);
nor U21049 (N_21049,N_17924,N_17598);
or U21050 (N_21050,N_19103,N_18058);
or U21051 (N_21051,N_18736,N_19057);
and U21052 (N_21052,N_18375,N_19731);
and U21053 (N_21053,N_19426,N_18088);
or U21054 (N_21054,N_18396,N_18340);
nand U21055 (N_21055,N_19457,N_18215);
and U21056 (N_21056,N_18650,N_18975);
and U21057 (N_21057,N_18531,N_18217);
nor U21058 (N_21058,N_18787,N_19782);
or U21059 (N_21059,N_17652,N_17518);
nor U21060 (N_21060,N_18481,N_19466);
and U21061 (N_21061,N_19849,N_19351);
or U21062 (N_21062,N_17694,N_17572);
nor U21063 (N_21063,N_19141,N_18544);
nand U21064 (N_21064,N_19424,N_18726);
nor U21065 (N_21065,N_17680,N_18154);
nand U21066 (N_21066,N_19202,N_19488);
nor U21067 (N_21067,N_18211,N_17998);
or U21068 (N_21068,N_18879,N_18846);
xor U21069 (N_21069,N_18904,N_19177);
and U21070 (N_21070,N_19663,N_18797);
nor U21071 (N_21071,N_19803,N_18455);
nor U21072 (N_21072,N_18674,N_17960);
nand U21073 (N_21073,N_19595,N_17762);
and U21074 (N_21074,N_18176,N_19837);
and U21075 (N_21075,N_17754,N_18007);
nor U21076 (N_21076,N_17580,N_19522);
nand U21077 (N_21077,N_18151,N_19590);
and U21078 (N_21078,N_17841,N_19341);
and U21079 (N_21079,N_18283,N_18063);
nor U21080 (N_21080,N_19870,N_19193);
nor U21081 (N_21081,N_18748,N_19887);
and U21082 (N_21082,N_18087,N_18561);
or U21083 (N_21083,N_18174,N_18577);
nand U21084 (N_21084,N_17950,N_18207);
or U21085 (N_21085,N_18503,N_19878);
nor U21086 (N_21086,N_19374,N_19242);
and U21087 (N_21087,N_18175,N_19303);
nor U21088 (N_21088,N_18684,N_19966);
nor U21089 (N_21089,N_18601,N_17974);
or U21090 (N_21090,N_19812,N_19264);
nand U21091 (N_21091,N_19479,N_17593);
or U21092 (N_21092,N_18934,N_17627);
and U21093 (N_21093,N_18135,N_19019);
nand U21094 (N_21094,N_17973,N_17722);
nand U21095 (N_21095,N_19974,N_17911);
nand U21096 (N_21096,N_18519,N_17791);
nor U21097 (N_21097,N_18049,N_18459);
and U21098 (N_21098,N_19408,N_18525);
nand U21099 (N_21099,N_17889,N_18523);
nand U21100 (N_21100,N_19126,N_18512);
nand U21101 (N_21101,N_19645,N_19768);
or U21102 (N_21102,N_19334,N_18812);
and U21103 (N_21103,N_18232,N_17937);
nand U21104 (N_21104,N_17919,N_17763);
or U21105 (N_21105,N_18914,N_17678);
nand U21106 (N_21106,N_18111,N_18552);
nand U21107 (N_21107,N_19133,N_19340);
or U21108 (N_21108,N_19172,N_19078);
nor U21109 (N_21109,N_18698,N_19839);
and U21110 (N_21110,N_19631,N_19445);
nand U21111 (N_21111,N_19330,N_19114);
nand U21112 (N_21112,N_19232,N_19833);
and U21113 (N_21113,N_17714,N_19166);
or U21114 (N_21114,N_19828,N_19693);
and U21115 (N_21115,N_17577,N_18995);
or U21116 (N_21116,N_19191,N_18094);
nand U21117 (N_21117,N_19933,N_19294);
or U21118 (N_21118,N_18012,N_17705);
and U21119 (N_21119,N_19724,N_18428);
nor U21120 (N_21120,N_18911,N_17737);
or U21121 (N_21121,N_18243,N_18803);
and U21122 (N_21122,N_19745,N_19597);
nand U21123 (N_21123,N_18851,N_18072);
nand U21124 (N_21124,N_19519,N_18598);
nor U21125 (N_21125,N_19712,N_19832);
nor U21126 (N_21126,N_19654,N_17554);
nor U21127 (N_21127,N_19669,N_19044);
nor U21128 (N_21128,N_19130,N_18602);
nand U21129 (N_21129,N_19721,N_19994);
xnor U21130 (N_21130,N_18657,N_19312);
and U21131 (N_21131,N_17887,N_19921);
nor U21132 (N_21132,N_17914,N_18567);
or U21133 (N_21133,N_18329,N_19888);
or U21134 (N_21134,N_18091,N_17612);
or U21135 (N_21135,N_18272,N_17849);
nand U21136 (N_21136,N_19099,N_17822);
nand U21137 (N_21137,N_19569,N_17682);
nand U21138 (N_21138,N_18699,N_19277);
and U21139 (N_21139,N_17543,N_17892);
nor U21140 (N_21140,N_18008,N_18332);
and U21141 (N_21141,N_19845,N_19083);
nor U21142 (N_21142,N_18279,N_19749);
nand U21143 (N_21143,N_17902,N_19053);
or U21144 (N_21144,N_19725,N_19413);
nor U21145 (N_21145,N_18326,N_19808);
nand U21146 (N_21146,N_17717,N_17933);
nor U21147 (N_21147,N_17549,N_19755);
nor U21148 (N_21148,N_18930,N_18691);
nor U21149 (N_21149,N_19514,N_18301);
nand U21150 (N_21150,N_17647,N_18394);
or U21151 (N_21151,N_19150,N_18330);
nor U21152 (N_21152,N_18285,N_17824);
and U21153 (N_21153,N_19022,N_17686);
and U21154 (N_21154,N_18315,N_18568);
nor U21155 (N_21155,N_19877,N_17716);
or U21156 (N_21156,N_18286,N_18947);
nor U21157 (N_21157,N_19687,N_19436);
nand U21158 (N_21158,N_19850,N_19806);
nor U21159 (N_21159,N_19148,N_19699);
or U21160 (N_21160,N_19314,N_18288);
nand U21161 (N_21161,N_18590,N_18082);
or U21162 (N_21162,N_18308,N_19707);
or U21163 (N_21163,N_17795,N_18341);
or U21164 (N_21164,N_19957,N_19224);
or U21165 (N_21165,N_19056,N_19769);
nor U21166 (N_21166,N_18583,N_18075);
or U21167 (N_21167,N_18412,N_17740);
nor U21168 (N_21168,N_19867,N_18499);
or U21169 (N_21169,N_17997,N_18573);
nand U21170 (N_21170,N_17851,N_19302);
nor U21171 (N_21171,N_19265,N_18370);
or U21172 (N_21172,N_18588,N_18885);
or U21173 (N_21173,N_17508,N_19797);
and U21174 (N_21174,N_19238,N_18893);
nand U21175 (N_21175,N_18675,N_17535);
nor U21176 (N_21176,N_18856,N_19187);
and U21177 (N_21177,N_19847,N_17616);
nor U21178 (N_21178,N_17934,N_19556);
nor U21179 (N_21179,N_18085,N_19272);
nor U21180 (N_21180,N_18909,N_17642);
and U21181 (N_21181,N_19606,N_19620);
nand U21182 (N_21182,N_19279,N_17985);
or U21183 (N_21183,N_19973,N_19964);
nand U21184 (N_21184,N_17781,N_18423);
and U21185 (N_21185,N_18103,N_19430);
or U21186 (N_21186,N_19299,N_19694);
or U21187 (N_21187,N_19767,N_17803);
nor U21188 (N_21188,N_17537,N_19079);
and U21189 (N_21189,N_18973,N_17946);
nor U21190 (N_21190,N_18612,N_18952);
or U21191 (N_21191,N_18516,N_18543);
nor U21192 (N_21192,N_18184,N_19826);
nand U21193 (N_21193,N_18533,N_19055);
or U21194 (N_21194,N_19988,N_18109);
or U21195 (N_21195,N_17953,N_18700);
and U21196 (N_21196,N_18026,N_19089);
or U21197 (N_21197,N_18364,N_19300);
or U21198 (N_21198,N_17913,N_18131);
and U21199 (N_21199,N_19102,N_18758);
or U21200 (N_21200,N_18536,N_19672);
and U21201 (N_21201,N_17830,N_19758);
nand U21202 (N_21202,N_18744,N_18144);
nand U21203 (N_21203,N_18114,N_18432);
nand U21204 (N_21204,N_19670,N_17609);
or U21205 (N_21205,N_19865,N_18179);
and U21206 (N_21206,N_17743,N_19703);
or U21207 (N_21207,N_19253,N_18204);
nor U21208 (N_21208,N_18137,N_18158);
nor U21209 (N_21209,N_17944,N_19559);
and U21210 (N_21210,N_19793,N_17768);
or U21211 (N_21211,N_19984,N_18949);
and U21212 (N_21212,N_18353,N_18276);
nor U21213 (N_21213,N_19443,N_19131);
or U21214 (N_21214,N_19051,N_18596);
nor U21215 (N_21215,N_19818,N_18246);
or U21216 (N_21216,N_18676,N_19701);
or U21217 (N_21217,N_18452,N_19389);
nor U21218 (N_21218,N_17900,N_17615);
or U21219 (N_21219,N_18016,N_19844);
nand U21220 (N_21220,N_18587,N_18504);
and U21221 (N_21221,N_17735,N_18564);
or U21222 (N_21222,N_17595,N_19991);
or U21223 (N_21223,N_17588,N_18056);
nand U21224 (N_21224,N_18514,N_18581);
nor U21225 (N_21225,N_17898,N_19588);
nand U21226 (N_21226,N_19220,N_19577);
nor U21227 (N_21227,N_19852,N_18167);
or U21228 (N_21228,N_18268,N_17925);
nand U21229 (N_21229,N_19881,N_17962);
xor U21230 (N_21230,N_18881,N_19894);
or U21231 (N_21231,N_19840,N_19813);
or U21232 (N_21232,N_19993,N_17848);
nor U21233 (N_21233,N_18404,N_17794);
or U21234 (N_21234,N_19315,N_19409);
nand U21235 (N_21235,N_19997,N_19387);
nor U21236 (N_21236,N_19060,N_18877);
and U21237 (N_21237,N_19003,N_19034);
nand U21238 (N_21238,N_17667,N_19827);
and U21239 (N_21239,N_17906,N_19018);
or U21240 (N_21240,N_17977,N_18528);
or U21241 (N_21241,N_19568,N_18492);
nor U21242 (N_21242,N_19117,N_18468);
and U21243 (N_21243,N_18319,N_19244);
and U21244 (N_21244,N_17901,N_19543);
nand U21245 (N_21245,N_19101,N_17561);
or U21246 (N_21246,N_18894,N_17724);
nand U21247 (N_21247,N_19026,N_17562);
nor U21248 (N_21248,N_18713,N_19205);
nor U21249 (N_21249,N_18159,N_17523);
nand U21250 (N_21250,N_17613,N_19460);
nor U21251 (N_21251,N_19622,N_18719);
and U21252 (N_21252,N_19629,N_17957);
nand U21253 (N_21253,N_17701,N_18297);
nor U21254 (N_21254,N_18969,N_19347);
or U21255 (N_21255,N_18356,N_17698);
and U21256 (N_21256,N_18872,N_18472);
or U21257 (N_21257,N_19340,N_18277);
nor U21258 (N_21258,N_17711,N_18657);
nor U21259 (N_21259,N_18219,N_19498);
nor U21260 (N_21260,N_19250,N_19680);
or U21261 (N_21261,N_18301,N_19275);
or U21262 (N_21262,N_19273,N_19233);
or U21263 (N_21263,N_19702,N_17873);
nor U21264 (N_21264,N_17744,N_17501);
nor U21265 (N_21265,N_18581,N_17866);
nor U21266 (N_21266,N_18156,N_19922);
nor U21267 (N_21267,N_18309,N_18227);
or U21268 (N_21268,N_18634,N_18758);
nor U21269 (N_21269,N_18450,N_19290);
and U21270 (N_21270,N_18930,N_17528);
and U21271 (N_21271,N_18252,N_19176);
or U21272 (N_21272,N_17741,N_18385);
nand U21273 (N_21273,N_19015,N_19752);
and U21274 (N_21274,N_19853,N_17934);
and U21275 (N_21275,N_19282,N_18394);
nor U21276 (N_21276,N_19534,N_18651);
nand U21277 (N_21277,N_18133,N_18548);
or U21278 (N_21278,N_18105,N_17711);
or U21279 (N_21279,N_19913,N_18770);
nand U21280 (N_21280,N_17663,N_18853);
nand U21281 (N_21281,N_18896,N_17597);
or U21282 (N_21282,N_19510,N_19597);
and U21283 (N_21283,N_17581,N_19235);
nand U21284 (N_21284,N_19654,N_18172);
nor U21285 (N_21285,N_19410,N_18381);
nor U21286 (N_21286,N_18736,N_18840);
nor U21287 (N_21287,N_19003,N_19742);
nand U21288 (N_21288,N_17598,N_18572);
xor U21289 (N_21289,N_18259,N_19950);
nand U21290 (N_21290,N_18136,N_18561);
nor U21291 (N_21291,N_18575,N_18200);
and U21292 (N_21292,N_19349,N_19021);
nor U21293 (N_21293,N_18962,N_17549);
or U21294 (N_21294,N_19861,N_19709);
and U21295 (N_21295,N_18906,N_19618);
nor U21296 (N_21296,N_18663,N_18252);
nor U21297 (N_21297,N_19821,N_17839);
and U21298 (N_21298,N_18351,N_19800);
nor U21299 (N_21299,N_18511,N_18825);
nor U21300 (N_21300,N_17526,N_18738);
or U21301 (N_21301,N_18724,N_19246);
nor U21302 (N_21302,N_18732,N_19575);
or U21303 (N_21303,N_18044,N_18037);
nor U21304 (N_21304,N_18025,N_19165);
nor U21305 (N_21305,N_19793,N_18073);
or U21306 (N_21306,N_19300,N_19270);
nor U21307 (N_21307,N_18480,N_18796);
nor U21308 (N_21308,N_18973,N_19778);
nand U21309 (N_21309,N_18286,N_18841);
and U21310 (N_21310,N_18877,N_18312);
xnor U21311 (N_21311,N_19325,N_19104);
nor U21312 (N_21312,N_19962,N_18679);
or U21313 (N_21313,N_19985,N_18806);
nand U21314 (N_21314,N_17948,N_18050);
and U21315 (N_21315,N_19336,N_17658);
nor U21316 (N_21316,N_19419,N_18170);
or U21317 (N_21317,N_18251,N_17804);
nor U21318 (N_21318,N_17617,N_18926);
nand U21319 (N_21319,N_19954,N_18418);
and U21320 (N_21320,N_18139,N_18127);
nand U21321 (N_21321,N_18987,N_18888);
and U21322 (N_21322,N_18170,N_18799);
nor U21323 (N_21323,N_18555,N_19549);
and U21324 (N_21324,N_18633,N_19604);
or U21325 (N_21325,N_17894,N_19481);
or U21326 (N_21326,N_17767,N_19004);
or U21327 (N_21327,N_18397,N_19902);
xnor U21328 (N_21328,N_17530,N_18210);
nor U21329 (N_21329,N_18865,N_18409);
or U21330 (N_21330,N_19243,N_18535);
nor U21331 (N_21331,N_19575,N_18553);
or U21332 (N_21332,N_19769,N_19808);
nor U21333 (N_21333,N_19309,N_19675);
and U21334 (N_21334,N_18209,N_18991);
or U21335 (N_21335,N_18601,N_19624);
and U21336 (N_21336,N_19724,N_17692);
or U21337 (N_21337,N_19660,N_18677);
and U21338 (N_21338,N_18119,N_19693);
and U21339 (N_21339,N_18759,N_17562);
and U21340 (N_21340,N_19017,N_18103);
nand U21341 (N_21341,N_19050,N_18674);
nor U21342 (N_21342,N_19286,N_19051);
nand U21343 (N_21343,N_19971,N_19142);
and U21344 (N_21344,N_17854,N_18321);
nor U21345 (N_21345,N_18425,N_18279);
nor U21346 (N_21346,N_19328,N_18982);
nor U21347 (N_21347,N_19338,N_18219);
or U21348 (N_21348,N_19287,N_18781);
nand U21349 (N_21349,N_18186,N_19924);
nand U21350 (N_21350,N_18850,N_19803);
nor U21351 (N_21351,N_18919,N_17832);
and U21352 (N_21352,N_19656,N_17870);
nor U21353 (N_21353,N_19633,N_18831);
or U21354 (N_21354,N_19172,N_19105);
and U21355 (N_21355,N_18803,N_19509);
or U21356 (N_21356,N_19387,N_18764);
nor U21357 (N_21357,N_18350,N_19145);
and U21358 (N_21358,N_18917,N_19716);
xor U21359 (N_21359,N_18450,N_17636);
and U21360 (N_21360,N_19003,N_18404);
nor U21361 (N_21361,N_18370,N_17853);
nand U21362 (N_21362,N_19383,N_18840);
nor U21363 (N_21363,N_18728,N_17819);
or U21364 (N_21364,N_19027,N_18944);
nand U21365 (N_21365,N_19123,N_17881);
and U21366 (N_21366,N_19421,N_18538);
nand U21367 (N_21367,N_18187,N_17505);
nand U21368 (N_21368,N_17716,N_18942);
or U21369 (N_21369,N_19078,N_19407);
or U21370 (N_21370,N_19136,N_19671);
nand U21371 (N_21371,N_18853,N_19157);
nor U21372 (N_21372,N_18152,N_18750);
and U21373 (N_21373,N_19273,N_17648);
or U21374 (N_21374,N_17676,N_19519);
xor U21375 (N_21375,N_18377,N_17695);
and U21376 (N_21376,N_19470,N_18336);
and U21377 (N_21377,N_19967,N_17964);
nand U21378 (N_21378,N_19536,N_18316);
nor U21379 (N_21379,N_17634,N_19762);
and U21380 (N_21380,N_19981,N_19571);
nor U21381 (N_21381,N_18917,N_19496);
or U21382 (N_21382,N_19518,N_19215);
nor U21383 (N_21383,N_19526,N_18242);
nor U21384 (N_21384,N_18333,N_19650);
or U21385 (N_21385,N_19195,N_17518);
or U21386 (N_21386,N_19550,N_18626);
or U21387 (N_21387,N_18315,N_19339);
nor U21388 (N_21388,N_19301,N_19595);
or U21389 (N_21389,N_19942,N_19221);
nor U21390 (N_21390,N_18160,N_18785);
and U21391 (N_21391,N_19991,N_19737);
or U21392 (N_21392,N_19034,N_19728);
nand U21393 (N_21393,N_18337,N_19049);
or U21394 (N_21394,N_19360,N_17819);
nand U21395 (N_21395,N_19333,N_17737);
or U21396 (N_21396,N_18516,N_19929);
nor U21397 (N_21397,N_18614,N_19659);
and U21398 (N_21398,N_19579,N_17653);
nor U21399 (N_21399,N_19292,N_19497);
and U21400 (N_21400,N_18370,N_17704);
and U21401 (N_21401,N_19542,N_17718);
nand U21402 (N_21402,N_17699,N_18377);
nand U21403 (N_21403,N_17971,N_19118);
nand U21404 (N_21404,N_17973,N_19179);
and U21405 (N_21405,N_19318,N_18426);
nand U21406 (N_21406,N_17605,N_19628);
nor U21407 (N_21407,N_18899,N_19661);
nand U21408 (N_21408,N_18283,N_18036);
and U21409 (N_21409,N_18443,N_18979);
or U21410 (N_21410,N_19476,N_19110);
and U21411 (N_21411,N_19408,N_17968);
nor U21412 (N_21412,N_19899,N_19059);
nand U21413 (N_21413,N_19630,N_19220);
or U21414 (N_21414,N_18729,N_18727);
nor U21415 (N_21415,N_18709,N_18788);
and U21416 (N_21416,N_18717,N_17536);
nand U21417 (N_21417,N_19765,N_17677);
nor U21418 (N_21418,N_18987,N_19576);
and U21419 (N_21419,N_18875,N_19862);
nand U21420 (N_21420,N_19778,N_17828);
nor U21421 (N_21421,N_17596,N_18405);
and U21422 (N_21422,N_17612,N_19812);
and U21423 (N_21423,N_18516,N_18773);
nor U21424 (N_21424,N_18076,N_19629);
and U21425 (N_21425,N_19849,N_18225);
or U21426 (N_21426,N_19866,N_18683);
nand U21427 (N_21427,N_17621,N_18141);
nand U21428 (N_21428,N_18185,N_18895);
nand U21429 (N_21429,N_18443,N_18182);
nand U21430 (N_21430,N_19671,N_19934);
nor U21431 (N_21431,N_19504,N_19997);
or U21432 (N_21432,N_17510,N_19386);
or U21433 (N_21433,N_17993,N_18638);
nand U21434 (N_21434,N_19239,N_19507);
nor U21435 (N_21435,N_17997,N_19714);
and U21436 (N_21436,N_18083,N_19532);
nand U21437 (N_21437,N_19157,N_19891);
nand U21438 (N_21438,N_19669,N_18969);
and U21439 (N_21439,N_19049,N_18088);
nand U21440 (N_21440,N_18008,N_18510);
and U21441 (N_21441,N_18220,N_18828);
and U21442 (N_21442,N_19276,N_19717);
xnor U21443 (N_21443,N_18608,N_18224);
nand U21444 (N_21444,N_18100,N_18150);
xnor U21445 (N_21445,N_18565,N_19437);
and U21446 (N_21446,N_19990,N_19974);
nand U21447 (N_21447,N_18571,N_17675);
or U21448 (N_21448,N_19441,N_19402);
and U21449 (N_21449,N_19139,N_17507);
or U21450 (N_21450,N_18030,N_18460);
nor U21451 (N_21451,N_17525,N_17916);
and U21452 (N_21452,N_19279,N_18825);
or U21453 (N_21453,N_19419,N_19376);
or U21454 (N_21454,N_19390,N_19355);
nand U21455 (N_21455,N_18232,N_19442);
or U21456 (N_21456,N_19182,N_17658);
nor U21457 (N_21457,N_19439,N_19334);
or U21458 (N_21458,N_19558,N_19030);
nand U21459 (N_21459,N_17702,N_18000);
nand U21460 (N_21460,N_17983,N_19861);
nor U21461 (N_21461,N_19934,N_18529);
nand U21462 (N_21462,N_19837,N_17603);
nor U21463 (N_21463,N_19808,N_17688);
nor U21464 (N_21464,N_18466,N_18310);
nor U21465 (N_21465,N_18529,N_19208);
nor U21466 (N_21466,N_19405,N_19751);
nand U21467 (N_21467,N_18249,N_18173);
or U21468 (N_21468,N_18074,N_18523);
and U21469 (N_21469,N_19538,N_19347);
nand U21470 (N_21470,N_18948,N_19873);
or U21471 (N_21471,N_18486,N_17521);
or U21472 (N_21472,N_18921,N_19360);
nand U21473 (N_21473,N_19651,N_19774);
nand U21474 (N_21474,N_18920,N_19620);
nand U21475 (N_21475,N_19839,N_19283);
nand U21476 (N_21476,N_19734,N_19794);
or U21477 (N_21477,N_19127,N_18259);
nand U21478 (N_21478,N_17639,N_19759);
nor U21479 (N_21479,N_17679,N_18058);
xor U21480 (N_21480,N_19242,N_17696);
or U21481 (N_21481,N_17878,N_19702);
and U21482 (N_21482,N_17781,N_19543);
nor U21483 (N_21483,N_17679,N_17983);
nand U21484 (N_21484,N_18559,N_18843);
and U21485 (N_21485,N_18616,N_19164);
or U21486 (N_21486,N_19867,N_17853);
and U21487 (N_21487,N_18156,N_19459);
xor U21488 (N_21488,N_19972,N_18888);
or U21489 (N_21489,N_18087,N_19145);
nor U21490 (N_21490,N_18859,N_18979);
and U21491 (N_21491,N_17559,N_18935);
nand U21492 (N_21492,N_19752,N_19985);
and U21493 (N_21493,N_18180,N_19429);
nor U21494 (N_21494,N_19094,N_17721);
nand U21495 (N_21495,N_18386,N_18565);
and U21496 (N_21496,N_19034,N_18867);
nand U21497 (N_21497,N_19829,N_17510);
or U21498 (N_21498,N_18124,N_19552);
xnor U21499 (N_21499,N_18897,N_19509);
or U21500 (N_21500,N_18811,N_18635);
nand U21501 (N_21501,N_19187,N_19016);
nor U21502 (N_21502,N_17662,N_19699);
or U21503 (N_21503,N_19069,N_19412);
nor U21504 (N_21504,N_19071,N_17911);
or U21505 (N_21505,N_18048,N_17668);
and U21506 (N_21506,N_18526,N_18276);
nor U21507 (N_21507,N_18937,N_17974);
and U21508 (N_21508,N_18981,N_18394);
nand U21509 (N_21509,N_19093,N_18603);
nor U21510 (N_21510,N_17833,N_17739);
nand U21511 (N_21511,N_18468,N_19346);
and U21512 (N_21512,N_18727,N_19871);
nand U21513 (N_21513,N_18654,N_18028);
and U21514 (N_21514,N_18501,N_19653);
nand U21515 (N_21515,N_19216,N_18649);
and U21516 (N_21516,N_18007,N_17547);
nor U21517 (N_21517,N_19791,N_18968);
nor U21518 (N_21518,N_19951,N_18606);
nand U21519 (N_21519,N_18300,N_18369);
or U21520 (N_21520,N_17809,N_18778);
xor U21521 (N_21521,N_19984,N_19445);
nand U21522 (N_21522,N_19364,N_18996);
and U21523 (N_21523,N_18059,N_17915);
or U21524 (N_21524,N_19442,N_19949);
or U21525 (N_21525,N_19574,N_18383);
nand U21526 (N_21526,N_19149,N_19854);
and U21527 (N_21527,N_18754,N_17628);
nor U21528 (N_21528,N_18708,N_17548);
or U21529 (N_21529,N_19375,N_19729);
nor U21530 (N_21530,N_17531,N_19924);
nor U21531 (N_21531,N_19149,N_17674);
and U21532 (N_21532,N_19500,N_17742);
and U21533 (N_21533,N_18585,N_19852);
or U21534 (N_21534,N_19959,N_19474);
or U21535 (N_21535,N_19308,N_17847);
nand U21536 (N_21536,N_19790,N_18899);
xnor U21537 (N_21537,N_19533,N_18679);
nor U21538 (N_21538,N_18254,N_19112);
and U21539 (N_21539,N_18181,N_17927);
or U21540 (N_21540,N_18405,N_18343);
or U21541 (N_21541,N_18191,N_17968);
nand U21542 (N_21542,N_17990,N_19480);
or U21543 (N_21543,N_19545,N_19305);
and U21544 (N_21544,N_18960,N_19598);
nor U21545 (N_21545,N_18955,N_19245);
xnor U21546 (N_21546,N_19477,N_18534);
nand U21547 (N_21547,N_19914,N_18332);
nand U21548 (N_21548,N_19473,N_19652);
nor U21549 (N_21549,N_17945,N_18074);
or U21550 (N_21550,N_17813,N_19014);
and U21551 (N_21551,N_18765,N_17770);
nand U21552 (N_21552,N_19803,N_19629);
nand U21553 (N_21553,N_19838,N_18116);
or U21554 (N_21554,N_18022,N_18804);
and U21555 (N_21555,N_19713,N_18377);
or U21556 (N_21556,N_17620,N_18203);
or U21557 (N_21557,N_19023,N_17864);
nor U21558 (N_21558,N_18635,N_19116);
nand U21559 (N_21559,N_18776,N_18582);
nor U21560 (N_21560,N_19814,N_19450);
and U21561 (N_21561,N_18148,N_18251);
or U21562 (N_21562,N_19291,N_19238);
or U21563 (N_21563,N_19076,N_19889);
or U21564 (N_21564,N_18796,N_17771);
nor U21565 (N_21565,N_18609,N_19763);
nor U21566 (N_21566,N_17967,N_17558);
and U21567 (N_21567,N_19551,N_19346);
nand U21568 (N_21568,N_18753,N_17710);
and U21569 (N_21569,N_18734,N_18825);
nor U21570 (N_21570,N_18857,N_18329);
or U21571 (N_21571,N_18990,N_18712);
or U21572 (N_21572,N_17770,N_19401);
and U21573 (N_21573,N_18440,N_18499);
nand U21574 (N_21574,N_17635,N_17758);
nand U21575 (N_21575,N_19170,N_18914);
or U21576 (N_21576,N_19404,N_17640);
nand U21577 (N_21577,N_18334,N_17712);
and U21578 (N_21578,N_19096,N_19125);
or U21579 (N_21579,N_19624,N_18048);
nor U21580 (N_21580,N_19981,N_19141);
or U21581 (N_21581,N_18516,N_18532);
nor U21582 (N_21582,N_19127,N_19435);
xor U21583 (N_21583,N_18710,N_18742);
nor U21584 (N_21584,N_18890,N_19535);
and U21585 (N_21585,N_17936,N_19576);
nand U21586 (N_21586,N_17854,N_18484);
nand U21587 (N_21587,N_18025,N_18616);
nand U21588 (N_21588,N_19858,N_17501);
and U21589 (N_21589,N_18627,N_17828);
and U21590 (N_21590,N_19898,N_17525);
nor U21591 (N_21591,N_19174,N_18918);
and U21592 (N_21592,N_19417,N_18088);
nand U21593 (N_21593,N_18290,N_18327);
or U21594 (N_21594,N_19657,N_18865);
xor U21595 (N_21595,N_19903,N_18623);
or U21596 (N_21596,N_19451,N_19373);
nand U21597 (N_21597,N_17983,N_18744);
nand U21598 (N_21598,N_17538,N_18741);
nor U21599 (N_21599,N_19604,N_17820);
or U21600 (N_21600,N_19301,N_19104);
and U21601 (N_21601,N_18810,N_19106);
and U21602 (N_21602,N_19035,N_19389);
nor U21603 (N_21603,N_18815,N_19184);
or U21604 (N_21604,N_18452,N_18988);
and U21605 (N_21605,N_19856,N_18338);
or U21606 (N_21606,N_19350,N_19638);
and U21607 (N_21607,N_17576,N_18926);
nand U21608 (N_21608,N_18744,N_18747);
nand U21609 (N_21609,N_18156,N_19773);
nand U21610 (N_21610,N_19696,N_17595);
and U21611 (N_21611,N_19861,N_18833);
or U21612 (N_21612,N_18887,N_18636);
and U21613 (N_21613,N_19935,N_17699);
nor U21614 (N_21614,N_19955,N_18524);
nor U21615 (N_21615,N_19464,N_19518);
nand U21616 (N_21616,N_18389,N_19703);
nor U21617 (N_21617,N_18068,N_18137);
nand U21618 (N_21618,N_17802,N_18509);
nor U21619 (N_21619,N_19349,N_18022);
or U21620 (N_21620,N_19653,N_18015);
and U21621 (N_21621,N_19634,N_19299);
nor U21622 (N_21622,N_18313,N_19681);
and U21623 (N_21623,N_19743,N_19746);
nand U21624 (N_21624,N_19870,N_19167);
nand U21625 (N_21625,N_19370,N_17572);
nand U21626 (N_21626,N_18407,N_18943);
and U21627 (N_21627,N_18362,N_19036);
nor U21628 (N_21628,N_19351,N_18918);
nand U21629 (N_21629,N_18003,N_18072);
or U21630 (N_21630,N_19556,N_18176);
nor U21631 (N_21631,N_19866,N_18759);
and U21632 (N_21632,N_18123,N_18126);
or U21633 (N_21633,N_19576,N_17769);
nor U21634 (N_21634,N_19570,N_19301);
and U21635 (N_21635,N_18960,N_18493);
nor U21636 (N_21636,N_19014,N_19760);
xnor U21637 (N_21637,N_19975,N_18860);
nand U21638 (N_21638,N_19330,N_18743);
and U21639 (N_21639,N_19078,N_19349);
or U21640 (N_21640,N_18550,N_18164);
nor U21641 (N_21641,N_17971,N_19824);
and U21642 (N_21642,N_17798,N_19863);
nor U21643 (N_21643,N_17893,N_18157);
or U21644 (N_21644,N_19322,N_19531);
nand U21645 (N_21645,N_18743,N_17669);
and U21646 (N_21646,N_18498,N_19533);
nand U21647 (N_21647,N_19056,N_18236);
and U21648 (N_21648,N_19183,N_19187);
and U21649 (N_21649,N_19514,N_19203);
or U21650 (N_21650,N_17823,N_18311);
nor U21651 (N_21651,N_19656,N_17880);
or U21652 (N_21652,N_19497,N_18614);
xor U21653 (N_21653,N_19745,N_18073);
nor U21654 (N_21654,N_18902,N_19992);
or U21655 (N_21655,N_18512,N_17787);
or U21656 (N_21656,N_18974,N_19758);
and U21657 (N_21657,N_19181,N_19464);
xnor U21658 (N_21658,N_18580,N_17889);
nor U21659 (N_21659,N_17918,N_19383);
or U21660 (N_21660,N_19294,N_18945);
or U21661 (N_21661,N_19311,N_17643);
nand U21662 (N_21662,N_19909,N_18831);
nor U21663 (N_21663,N_19362,N_17520);
nor U21664 (N_21664,N_18455,N_18365);
or U21665 (N_21665,N_18015,N_19659);
or U21666 (N_21666,N_17899,N_17991);
nor U21667 (N_21667,N_18827,N_19937);
and U21668 (N_21668,N_17966,N_18841);
or U21669 (N_21669,N_18534,N_18489);
nor U21670 (N_21670,N_19848,N_19092);
nor U21671 (N_21671,N_18923,N_18015);
and U21672 (N_21672,N_19445,N_18917);
and U21673 (N_21673,N_19686,N_19823);
nor U21674 (N_21674,N_18654,N_18818);
and U21675 (N_21675,N_17823,N_19865);
and U21676 (N_21676,N_17599,N_19320);
nor U21677 (N_21677,N_18748,N_17955);
nand U21678 (N_21678,N_19027,N_17900);
nand U21679 (N_21679,N_19403,N_19307);
nor U21680 (N_21680,N_18300,N_18295);
nor U21681 (N_21681,N_18738,N_19593);
and U21682 (N_21682,N_19940,N_18114);
nor U21683 (N_21683,N_18032,N_18343);
or U21684 (N_21684,N_17870,N_19798);
xnor U21685 (N_21685,N_18822,N_17947);
nor U21686 (N_21686,N_19054,N_17796);
and U21687 (N_21687,N_17907,N_17857);
and U21688 (N_21688,N_18057,N_19776);
nand U21689 (N_21689,N_17621,N_17937);
or U21690 (N_21690,N_19199,N_19535);
nor U21691 (N_21691,N_19641,N_19386);
or U21692 (N_21692,N_19117,N_19568);
and U21693 (N_21693,N_18090,N_18927);
nand U21694 (N_21694,N_17774,N_17743);
and U21695 (N_21695,N_18544,N_18027);
nand U21696 (N_21696,N_18032,N_18430);
or U21697 (N_21697,N_17597,N_18713);
or U21698 (N_21698,N_19027,N_17848);
nor U21699 (N_21699,N_19448,N_18294);
nand U21700 (N_21700,N_19374,N_18852);
nor U21701 (N_21701,N_18808,N_18703);
nor U21702 (N_21702,N_19735,N_17928);
and U21703 (N_21703,N_18016,N_18152);
and U21704 (N_21704,N_19515,N_19937);
and U21705 (N_21705,N_18953,N_18516);
or U21706 (N_21706,N_18648,N_19100);
or U21707 (N_21707,N_17522,N_18154);
or U21708 (N_21708,N_17916,N_19018);
or U21709 (N_21709,N_18515,N_18758);
or U21710 (N_21710,N_18065,N_19915);
nand U21711 (N_21711,N_19521,N_19683);
and U21712 (N_21712,N_19832,N_18933);
nor U21713 (N_21713,N_19269,N_17860);
nor U21714 (N_21714,N_19841,N_18364);
or U21715 (N_21715,N_19765,N_19406);
or U21716 (N_21716,N_18086,N_18023);
nor U21717 (N_21717,N_17809,N_18529);
and U21718 (N_21718,N_18010,N_18558);
and U21719 (N_21719,N_18628,N_19154);
nor U21720 (N_21720,N_18796,N_18099);
nor U21721 (N_21721,N_19230,N_17642);
nand U21722 (N_21722,N_19908,N_18486);
nand U21723 (N_21723,N_19738,N_19833);
nand U21724 (N_21724,N_18197,N_17906);
and U21725 (N_21725,N_17528,N_19838);
nand U21726 (N_21726,N_19523,N_17931);
and U21727 (N_21727,N_17872,N_19507);
and U21728 (N_21728,N_19760,N_18561);
and U21729 (N_21729,N_18358,N_18291);
nand U21730 (N_21730,N_19972,N_19085);
nand U21731 (N_21731,N_19819,N_19300);
and U21732 (N_21732,N_19509,N_18207);
and U21733 (N_21733,N_18279,N_17718);
nor U21734 (N_21734,N_18365,N_18749);
nand U21735 (N_21735,N_18983,N_19979);
nor U21736 (N_21736,N_18640,N_17872);
or U21737 (N_21737,N_18329,N_17817);
nor U21738 (N_21738,N_18448,N_19113);
nand U21739 (N_21739,N_19992,N_19227);
or U21740 (N_21740,N_17600,N_19178);
nand U21741 (N_21741,N_18472,N_17848);
or U21742 (N_21742,N_17994,N_19068);
nand U21743 (N_21743,N_18492,N_18459);
or U21744 (N_21744,N_17905,N_17927);
nor U21745 (N_21745,N_17565,N_18218);
nand U21746 (N_21746,N_19057,N_19339);
or U21747 (N_21747,N_19480,N_19879);
or U21748 (N_21748,N_19936,N_19278);
or U21749 (N_21749,N_18968,N_19667);
xnor U21750 (N_21750,N_18661,N_18813);
or U21751 (N_21751,N_18057,N_18849);
and U21752 (N_21752,N_19209,N_19977);
or U21753 (N_21753,N_18822,N_18211);
and U21754 (N_21754,N_19844,N_19672);
or U21755 (N_21755,N_17657,N_19400);
and U21756 (N_21756,N_19958,N_18870);
or U21757 (N_21757,N_18153,N_18288);
and U21758 (N_21758,N_18174,N_18325);
nor U21759 (N_21759,N_18015,N_18767);
nand U21760 (N_21760,N_17770,N_18992);
and U21761 (N_21761,N_17503,N_18211);
and U21762 (N_21762,N_18535,N_17814);
xnor U21763 (N_21763,N_18130,N_17667);
nor U21764 (N_21764,N_18951,N_18508);
nand U21765 (N_21765,N_17600,N_18661);
nand U21766 (N_21766,N_18860,N_18078);
or U21767 (N_21767,N_17882,N_18196);
and U21768 (N_21768,N_19775,N_18217);
nor U21769 (N_21769,N_18158,N_18287);
nand U21770 (N_21770,N_19396,N_17551);
or U21771 (N_21771,N_18374,N_18904);
and U21772 (N_21772,N_17717,N_18307);
and U21773 (N_21773,N_19698,N_19726);
nor U21774 (N_21774,N_18319,N_19541);
nor U21775 (N_21775,N_17980,N_19809);
or U21776 (N_21776,N_17930,N_17543);
and U21777 (N_21777,N_18974,N_19404);
nand U21778 (N_21778,N_17951,N_19372);
or U21779 (N_21779,N_18567,N_18741);
or U21780 (N_21780,N_19161,N_17581);
and U21781 (N_21781,N_18000,N_18492);
nor U21782 (N_21782,N_19292,N_19160);
nand U21783 (N_21783,N_19685,N_18854);
nor U21784 (N_21784,N_18558,N_18846);
or U21785 (N_21785,N_17975,N_18909);
and U21786 (N_21786,N_19668,N_19099);
nor U21787 (N_21787,N_18914,N_19069);
nor U21788 (N_21788,N_18947,N_17953);
and U21789 (N_21789,N_19619,N_17831);
and U21790 (N_21790,N_17878,N_17895);
and U21791 (N_21791,N_19047,N_18321);
and U21792 (N_21792,N_17616,N_19560);
or U21793 (N_21793,N_19034,N_17502);
and U21794 (N_21794,N_17522,N_18720);
nor U21795 (N_21795,N_19734,N_18673);
or U21796 (N_21796,N_18554,N_17642);
nand U21797 (N_21797,N_19414,N_18453);
nand U21798 (N_21798,N_18458,N_19778);
or U21799 (N_21799,N_18108,N_19920);
and U21800 (N_21800,N_18660,N_19173);
and U21801 (N_21801,N_18192,N_19957);
or U21802 (N_21802,N_17844,N_19117);
and U21803 (N_21803,N_18433,N_18812);
nor U21804 (N_21804,N_17787,N_19156);
or U21805 (N_21805,N_19027,N_18399);
nor U21806 (N_21806,N_18951,N_19769);
nand U21807 (N_21807,N_17795,N_17875);
or U21808 (N_21808,N_18253,N_18149);
nor U21809 (N_21809,N_18174,N_19070);
and U21810 (N_21810,N_19569,N_18729);
nor U21811 (N_21811,N_18905,N_18891);
or U21812 (N_21812,N_18914,N_18600);
or U21813 (N_21813,N_19580,N_18277);
or U21814 (N_21814,N_19008,N_18229);
and U21815 (N_21815,N_18511,N_18644);
nor U21816 (N_21816,N_17562,N_19927);
or U21817 (N_21817,N_18084,N_19618);
nand U21818 (N_21818,N_17721,N_19282);
nand U21819 (N_21819,N_18833,N_18564);
xor U21820 (N_21820,N_19271,N_19744);
nand U21821 (N_21821,N_17952,N_17568);
and U21822 (N_21822,N_18987,N_17826);
and U21823 (N_21823,N_19645,N_19680);
nand U21824 (N_21824,N_19960,N_19530);
nor U21825 (N_21825,N_19335,N_18073);
or U21826 (N_21826,N_18018,N_17552);
or U21827 (N_21827,N_18801,N_18040);
nor U21828 (N_21828,N_17641,N_17824);
xnor U21829 (N_21829,N_19556,N_18174);
and U21830 (N_21830,N_17811,N_19184);
or U21831 (N_21831,N_19587,N_17631);
xnor U21832 (N_21832,N_17800,N_17712);
nor U21833 (N_21833,N_17927,N_19788);
and U21834 (N_21834,N_18586,N_18229);
xor U21835 (N_21835,N_17897,N_18956);
and U21836 (N_21836,N_19689,N_19657);
nor U21837 (N_21837,N_19462,N_18443);
and U21838 (N_21838,N_18542,N_17569);
nor U21839 (N_21839,N_19818,N_17861);
and U21840 (N_21840,N_18500,N_19621);
nor U21841 (N_21841,N_17574,N_19012);
nor U21842 (N_21842,N_17541,N_18969);
nor U21843 (N_21843,N_18506,N_19574);
nor U21844 (N_21844,N_18872,N_19582);
nand U21845 (N_21845,N_18574,N_18401);
nand U21846 (N_21846,N_19268,N_18672);
or U21847 (N_21847,N_19965,N_18038);
and U21848 (N_21848,N_19215,N_17951);
nor U21849 (N_21849,N_17895,N_17581);
nor U21850 (N_21850,N_18047,N_18598);
nor U21851 (N_21851,N_18249,N_19625);
nor U21852 (N_21852,N_17802,N_19978);
nand U21853 (N_21853,N_18529,N_19816);
nor U21854 (N_21854,N_19565,N_18642);
or U21855 (N_21855,N_18686,N_19464);
or U21856 (N_21856,N_17523,N_19953);
or U21857 (N_21857,N_19589,N_17501);
nand U21858 (N_21858,N_18643,N_17646);
or U21859 (N_21859,N_18155,N_19320);
nor U21860 (N_21860,N_19745,N_18986);
nor U21861 (N_21861,N_17938,N_17722);
nand U21862 (N_21862,N_19004,N_17814);
nand U21863 (N_21863,N_18652,N_18781);
or U21864 (N_21864,N_17584,N_17916);
and U21865 (N_21865,N_19714,N_18471);
and U21866 (N_21866,N_19617,N_18229);
or U21867 (N_21867,N_17987,N_18584);
nand U21868 (N_21868,N_19967,N_19397);
nand U21869 (N_21869,N_19108,N_19143);
nand U21870 (N_21870,N_19730,N_18675);
and U21871 (N_21871,N_19931,N_18132);
nand U21872 (N_21872,N_17898,N_18334);
and U21873 (N_21873,N_18470,N_19237);
nor U21874 (N_21874,N_18960,N_18867);
nand U21875 (N_21875,N_19525,N_18577);
and U21876 (N_21876,N_19570,N_19162);
nor U21877 (N_21877,N_19779,N_19266);
or U21878 (N_21878,N_18849,N_19098);
nand U21879 (N_21879,N_18372,N_19467);
or U21880 (N_21880,N_19971,N_17815);
nand U21881 (N_21881,N_18780,N_19580);
or U21882 (N_21882,N_18494,N_17699);
or U21883 (N_21883,N_18910,N_18316);
and U21884 (N_21884,N_17714,N_17841);
and U21885 (N_21885,N_18913,N_18658);
nor U21886 (N_21886,N_18443,N_18419);
and U21887 (N_21887,N_17958,N_18313);
nand U21888 (N_21888,N_17831,N_18239);
xnor U21889 (N_21889,N_18846,N_19992);
nor U21890 (N_21890,N_18924,N_18441);
and U21891 (N_21891,N_18049,N_19405);
or U21892 (N_21892,N_19448,N_18546);
nand U21893 (N_21893,N_17722,N_19360);
nor U21894 (N_21894,N_19934,N_19541);
xor U21895 (N_21895,N_19071,N_18349);
nand U21896 (N_21896,N_18443,N_18915);
or U21897 (N_21897,N_19098,N_19096);
nand U21898 (N_21898,N_18925,N_18993);
or U21899 (N_21899,N_18275,N_17863);
nor U21900 (N_21900,N_19885,N_17752);
nand U21901 (N_21901,N_17964,N_19376);
and U21902 (N_21902,N_18777,N_18252);
or U21903 (N_21903,N_19294,N_18849);
nor U21904 (N_21904,N_18333,N_18275);
nand U21905 (N_21905,N_17825,N_19755);
and U21906 (N_21906,N_18748,N_19976);
nor U21907 (N_21907,N_18653,N_18893);
or U21908 (N_21908,N_18082,N_18665);
nor U21909 (N_21909,N_17780,N_18582);
nand U21910 (N_21910,N_18856,N_17835);
or U21911 (N_21911,N_19302,N_19523);
nor U21912 (N_21912,N_19732,N_17894);
and U21913 (N_21913,N_18362,N_18292);
nor U21914 (N_21914,N_18316,N_18328);
nand U21915 (N_21915,N_18583,N_19521);
and U21916 (N_21916,N_17711,N_18794);
nand U21917 (N_21917,N_19675,N_19018);
and U21918 (N_21918,N_18250,N_17626);
and U21919 (N_21919,N_18446,N_18353);
nand U21920 (N_21920,N_18613,N_17533);
nand U21921 (N_21921,N_18493,N_19363);
or U21922 (N_21922,N_18474,N_17948);
nor U21923 (N_21923,N_19688,N_19530);
nand U21924 (N_21924,N_18529,N_17512);
or U21925 (N_21925,N_19014,N_18373);
and U21926 (N_21926,N_18664,N_18994);
and U21927 (N_21927,N_17735,N_19402);
and U21928 (N_21928,N_17897,N_17766);
and U21929 (N_21929,N_19367,N_18861);
or U21930 (N_21930,N_19801,N_18668);
nand U21931 (N_21931,N_19002,N_18370);
nor U21932 (N_21932,N_19867,N_19960);
and U21933 (N_21933,N_17707,N_19097);
nor U21934 (N_21934,N_17756,N_18737);
nand U21935 (N_21935,N_17699,N_18928);
or U21936 (N_21936,N_18424,N_18948);
nor U21937 (N_21937,N_19398,N_18867);
or U21938 (N_21938,N_18668,N_18628);
or U21939 (N_21939,N_18465,N_18213);
nor U21940 (N_21940,N_18720,N_19875);
nor U21941 (N_21941,N_19555,N_17979);
or U21942 (N_21942,N_19994,N_18661);
and U21943 (N_21943,N_18443,N_19044);
nor U21944 (N_21944,N_17737,N_17847);
or U21945 (N_21945,N_19783,N_18661);
or U21946 (N_21946,N_19661,N_18303);
or U21947 (N_21947,N_18126,N_19156);
nor U21948 (N_21948,N_18119,N_19280);
nand U21949 (N_21949,N_19334,N_18223);
or U21950 (N_21950,N_19618,N_18690);
or U21951 (N_21951,N_18089,N_18119);
nor U21952 (N_21952,N_18787,N_19515);
nor U21953 (N_21953,N_18146,N_17617);
or U21954 (N_21954,N_18957,N_17515);
nor U21955 (N_21955,N_19510,N_18128);
nor U21956 (N_21956,N_17648,N_18471);
and U21957 (N_21957,N_18490,N_18360);
nand U21958 (N_21958,N_18685,N_19209);
nor U21959 (N_21959,N_18250,N_17530);
nand U21960 (N_21960,N_18182,N_18677);
and U21961 (N_21961,N_19276,N_18462);
and U21962 (N_21962,N_19259,N_18511);
nor U21963 (N_21963,N_17816,N_19274);
nand U21964 (N_21964,N_19978,N_18437);
nand U21965 (N_21965,N_18997,N_18570);
and U21966 (N_21966,N_17835,N_19144);
nand U21967 (N_21967,N_18029,N_19743);
nor U21968 (N_21968,N_19666,N_19170);
nand U21969 (N_21969,N_19231,N_19579);
nand U21970 (N_21970,N_17652,N_18786);
nand U21971 (N_21971,N_18088,N_18024);
nand U21972 (N_21972,N_17565,N_18329);
nor U21973 (N_21973,N_18231,N_17571);
nor U21974 (N_21974,N_19651,N_18158);
nand U21975 (N_21975,N_17937,N_18444);
or U21976 (N_21976,N_18831,N_19043);
or U21977 (N_21977,N_19174,N_19915);
or U21978 (N_21978,N_17586,N_19271);
and U21979 (N_21979,N_18684,N_18166);
or U21980 (N_21980,N_18500,N_18490);
or U21981 (N_21981,N_18063,N_18382);
and U21982 (N_21982,N_17740,N_19814);
nor U21983 (N_21983,N_17704,N_18071);
nand U21984 (N_21984,N_19882,N_19912);
nor U21985 (N_21985,N_18485,N_18017);
nor U21986 (N_21986,N_18440,N_19884);
xor U21987 (N_21987,N_17547,N_19099);
nor U21988 (N_21988,N_19964,N_19398);
nand U21989 (N_21989,N_19935,N_17934);
or U21990 (N_21990,N_17931,N_17564);
xor U21991 (N_21991,N_17868,N_18822);
or U21992 (N_21992,N_18123,N_19867);
nand U21993 (N_21993,N_17712,N_19624);
and U21994 (N_21994,N_18321,N_19120);
nor U21995 (N_21995,N_18290,N_19305);
nand U21996 (N_21996,N_17711,N_19751);
nand U21997 (N_21997,N_17627,N_19175);
nand U21998 (N_21998,N_18720,N_17947);
or U21999 (N_21999,N_19750,N_19274);
and U22000 (N_22000,N_19405,N_18275);
or U22001 (N_22001,N_17870,N_18354);
and U22002 (N_22002,N_19690,N_19250);
nand U22003 (N_22003,N_19722,N_18018);
nor U22004 (N_22004,N_19246,N_18648);
xor U22005 (N_22005,N_18673,N_18500);
and U22006 (N_22006,N_19957,N_17915);
nand U22007 (N_22007,N_19932,N_18077);
and U22008 (N_22008,N_18488,N_18344);
or U22009 (N_22009,N_17871,N_18457);
nor U22010 (N_22010,N_19910,N_19245);
nand U22011 (N_22011,N_18191,N_17789);
or U22012 (N_22012,N_18013,N_18545);
or U22013 (N_22013,N_18719,N_19184);
nor U22014 (N_22014,N_19891,N_19759);
nor U22015 (N_22015,N_18254,N_17888);
nand U22016 (N_22016,N_17515,N_18419);
or U22017 (N_22017,N_18126,N_19425);
or U22018 (N_22018,N_19630,N_18428);
and U22019 (N_22019,N_19536,N_19446);
and U22020 (N_22020,N_18318,N_19442);
or U22021 (N_22021,N_18249,N_18690);
nand U22022 (N_22022,N_17724,N_19796);
nand U22023 (N_22023,N_19886,N_18963);
nor U22024 (N_22024,N_18543,N_18288);
nand U22025 (N_22025,N_19331,N_18050);
nor U22026 (N_22026,N_17841,N_17514);
or U22027 (N_22027,N_18634,N_19286);
and U22028 (N_22028,N_19669,N_19076);
and U22029 (N_22029,N_19792,N_18499);
nand U22030 (N_22030,N_18278,N_19748);
nor U22031 (N_22031,N_18132,N_19269);
and U22032 (N_22032,N_19458,N_19321);
or U22033 (N_22033,N_17512,N_19054);
or U22034 (N_22034,N_18320,N_19118);
nor U22035 (N_22035,N_18871,N_19519);
or U22036 (N_22036,N_18236,N_19248);
or U22037 (N_22037,N_18150,N_18743);
and U22038 (N_22038,N_19100,N_18771);
nor U22039 (N_22039,N_19044,N_19043);
nor U22040 (N_22040,N_18256,N_18275);
nor U22041 (N_22041,N_18451,N_19089);
and U22042 (N_22042,N_19626,N_19080);
xor U22043 (N_22043,N_18109,N_17706);
nor U22044 (N_22044,N_19515,N_19068);
nand U22045 (N_22045,N_17875,N_19790);
nand U22046 (N_22046,N_18994,N_17800);
nand U22047 (N_22047,N_19572,N_18389);
nand U22048 (N_22048,N_18225,N_19318);
nand U22049 (N_22049,N_17534,N_17539);
and U22050 (N_22050,N_18296,N_19187);
nand U22051 (N_22051,N_17722,N_18513);
nand U22052 (N_22052,N_19913,N_17700);
and U22053 (N_22053,N_18311,N_19813);
nand U22054 (N_22054,N_19240,N_19980);
and U22055 (N_22055,N_19082,N_18519);
and U22056 (N_22056,N_17997,N_19250);
nand U22057 (N_22057,N_18284,N_19323);
or U22058 (N_22058,N_18884,N_19925);
nor U22059 (N_22059,N_18875,N_18548);
or U22060 (N_22060,N_19294,N_18338);
nor U22061 (N_22061,N_18574,N_17824);
and U22062 (N_22062,N_18529,N_19549);
or U22063 (N_22063,N_17703,N_19202);
nand U22064 (N_22064,N_17867,N_19814);
and U22065 (N_22065,N_19424,N_19882);
or U22066 (N_22066,N_18013,N_17809);
nor U22067 (N_22067,N_19216,N_18337);
nand U22068 (N_22068,N_19675,N_18118);
nor U22069 (N_22069,N_17818,N_19463);
and U22070 (N_22070,N_17940,N_18622);
or U22071 (N_22071,N_19515,N_19384);
nor U22072 (N_22072,N_18767,N_19219);
or U22073 (N_22073,N_18988,N_18217);
or U22074 (N_22074,N_19419,N_18898);
nor U22075 (N_22075,N_18605,N_19491);
nand U22076 (N_22076,N_18205,N_18664);
nand U22077 (N_22077,N_19784,N_18181);
nor U22078 (N_22078,N_19028,N_18074);
xor U22079 (N_22079,N_17594,N_19579);
and U22080 (N_22080,N_19381,N_19667);
or U22081 (N_22081,N_19944,N_19320);
or U22082 (N_22082,N_18625,N_19019);
nand U22083 (N_22083,N_18715,N_17882);
nor U22084 (N_22084,N_17857,N_18570);
nand U22085 (N_22085,N_19856,N_19193);
or U22086 (N_22086,N_19114,N_18279);
or U22087 (N_22087,N_19640,N_18682);
or U22088 (N_22088,N_17677,N_17966);
nand U22089 (N_22089,N_19116,N_17643);
or U22090 (N_22090,N_18752,N_19970);
nor U22091 (N_22091,N_17572,N_19347);
xnor U22092 (N_22092,N_19299,N_19119);
or U22093 (N_22093,N_19576,N_18545);
xnor U22094 (N_22094,N_18505,N_19143);
nand U22095 (N_22095,N_19725,N_18306);
or U22096 (N_22096,N_17543,N_17764);
and U22097 (N_22097,N_17611,N_19539);
or U22098 (N_22098,N_17742,N_18790);
and U22099 (N_22099,N_18426,N_19637);
or U22100 (N_22100,N_18361,N_18587);
or U22101 (N_22101,N_19859,N_17876);
nand U22102 (N_22102,N_17638,N_17861);
nor U22103 (N_22103,N_19700,N_18796);
nand U22104 (N_22104,N_19621,N_19034);
or U22105 (N_22105,N_19302,N_18111);
or U22106 (N_22106,N_18509,N_18922);
nand U22107 (N_22107,N_19445,N_19832);
or U22108 (N_22108,N_19638,N_18909);
nor U22109 (N_22109,N_19444,N_18128);
and U22110 (N_22110,N_18191,N_19590);
or U22111 (N_22111,N_18605,N_17564);
nand U22112 (N_22112,N_18978,N_19034);
nand U22113 (N_22113,N_19022,N_18552);
nand U22114 (N_22114,N_18128,N_19353);
nand U22115 (N_22115,N_19068,N_17727);
or U22116 (N_22116,N_18112,N_19118);
nor U22117 (N_22117,N_19688,N_19842);
or U22118 (N_22118,N_17739,N_19556);
or U22119 (N_22119,N_18603,N_18995);
or U22120 (N_22120,N_17676,N_19793);
nand U22121 (N_22121,N_19038,N_19745);
nor U22122 (N_22122,N_18591,N_18118);
nand U22123 (N_22123,N_18231,N_19604);
and U22124 (N_22124,N_19983,N_18482);
or U22125 (N_22125,N_17944,N_18859);
and U22126 (N_22126,N_18344,N_19866);
nor U22127 (N_22127,N_18843,N_18127);
or U22128 (N_22128,N_17824,N_18975);
or U22129 (N_22129,N_19296,N_19087);
nand U22130 (N_22130,N_17599,N_19102);
and U22131 (N_22131,N_17607,N_19230);
nor U22132 (N_22132,N_17893,N_19718);
nor U22133 (N_22133,N_17705,N_18779);
nor U22134 (N_22134,N_18001,N_18137);
nand U22135 (N_22135,N_18834,N_18038);
nand U22136 (N_22136,N_18376,N_18792);
nor U22137 (N_22137,N_18884,N_18033);
nand U22138 (N_22138,N_18642,N_18282);
and U22139 (N_22139,N_18550,N_19044);
or U22140 (N_22140,N_19050,N_18240);
nand U22141 (N_22141,N_18552,N_19730);
and U22142 (N_22142,N_19164,N_19218);
or U22143 (N_22143,N_19203,N_19966);
nand U22144 (N_22144,N_19371,N_18577);
or U22145 (N_22145,N_18380,N_18087);
nor U22146 (N_22146,N_19861,N_19868);
nand U22147 (N_22147,N_19946,N_18878);
nor U22148 (N_22148,N_18273,N_17852);
nor U22149 (N_22149,N_19624,N_18976);
or U22150 (N_22150,N_19571,N_18704);
and U22151 (N_22151,N_19960,N_17807);
or U22152 (N_22152,N_17843,N_19263);
nand U22153 (N_22153,N_17781,N_18556);
nand U22154 (N_22154,N_19366,N_19189);
nor U22155 (N_22155,N_18328,N_17509);
nor U22156 (N_22156,N_18884,N_19392);
nand U22157 (N_22157,N_18403,N_18614);
and U22158 (N_22158,N_18955,N_18216);
or U22159 (N_22159,N_19077,N_19067);
nand U22160 (N_22160,N_18074,N_18306);
nor U22161 (N_22161,N_18119,N_18629);
nand U22162 (N_22162,N_19757,N_18150);
and U22163 (N_22163,N_18894,N_17921);
and U22164 (N_22164,N_19929,N_19051);
or U22165 (N_22165,N_19134,N_17583);
nor U22166 (N_22166,N_19459,N_18805);
and U22167 (N_22167,N_19648,N_19292);
nand U22168 (N_22168,N_17635,N_19740);
nand U22169 (N_22169,N_18146,N_19290);
or U22170 (N_22170,N_17842,N_19100);
nand U22171 (N_22171,N_19880,N_17705);
nand U22172 (N_22172,N_19860,N_19772);
or U22173 (N_22173,N_18807,N_19892);
nor U22174 (N_22174,N_18621,N_19323);
nand U22175 (N_22175,N_19634,N_17823);
nor U22176 (N_22176,N_17806,N_17797);
nand U22177 (N_22177,N_17563,N_19294);
nand U22178 (N_22178,N_18963,N_19164);
nor U22179 (N_22179,N_18445,N_19425);
nor U22180 (N_22180,N_18071,N_18443);
nand U22181 (N_22181,N_19308,N_19302);
and U22182 (N_22182,N_18418,N_18246);
nand U22183 (N_22183,N_19257,N_17854);
or U22184 (N_22184,N_18119,N_17568);
or U22185 (N_22185,N_19615,N_18228);
or U22186 (N_22186,N_19074,N_19940);
nand U22187 (N_22187,N_18602,N_19122);
nor U22188 (N_22188,N_18697,N_18826);
nand U22189 (N_22189,N_17638,N_19999);
or U22190 (N_22190,N_17510,N_18975);
or U22191 (N_22191,N_18116,N_17749);
or U22192 (N_22192,N_18498,N_18685);
and U22193 (N_22193,N_18356,N_17814);
nand U22194 (N_22194,N_19284,N_19685);
or U22195 (N_22195,N_19156,N_18078);
or U22196 (N_22196,N_19837,N_18446);
or U22197 (N_22197,N_19196,N_18145);
nand U22198 (N_22198,N_18108,N_19357);
or U22199 (N_22199,N_18395,N_18396);
nor U22200 (N_22200,N_17915,N_18631);
nor U22201 (N_22201,N_17522,N_17748);
or U22202 (N_22202,N_18861,N_19709);
nand U22203 (N_22203,N_19815,N_18545);
and U22204 (N_22204,N_18472,N_19807);
nand U22205 (N_22205,N_19084,N_19513);
nand U22206 (N_22206,N_17998,N_17784);
or U22207 (N_22207,N_18206,N_18214);
or U22208 (N_22208,N_19336,N_18994);
or U22209 (N_22209,N_19997,N_18930);
nand U22210 (N_22210,N_18331,N_18808);
nand U22211 (N_22211,N_18208,N_19519);
or U22212 (N_22212,N_19718,N_17830);
or U22213 (N_22213,N_19826,N_18185);
nor U22214 (N_22214,N_17977,N_17937);
nor U22215 (N_22215,N_19920,N_19159);
nor U22216 (N_22216,N_19364,N_19186);
nand U22217 (N_22217,N_17727,N_19432);
or U22218 (N_22218,N_18817,N_19944);
or U22219 (N_22219,N_18902,N_18237);
or U22220 (N_22220,N_18633,N_17552);
nand U22221 (N_22221,N_19531,N_17998);
and U22222 (N_22222,N_19586,N_19881);
nand U22223 (N_22223,N_18296,N_18153);
nor U22224 (N_22224,N_18251,N_18759);
or U22225 (N_22225,N_19363,N_19792);
and U22226 (N_22226,N_18257,N_19624);
nand U22227 (N_22227,N_17639,N_17584);
nor U22228 (N_22228,N_19639,N_18110);
and U22229 (N_22229,N_18384,N_18627);
or U22230 (N_22230,N_19768,N_19025);
nand U22231 (N_22231,N_18165,N_18415);
or U22232 (N_22232,N_18301,N_18288);
or U22233 (N_22233,N_17835,N_18569);
or U22234 (N_22234,N_17978,N_17946);
and U22235 (N_22235,N_19521,N_19884);
and U22236 (N_22236,N_19334,N_18747);
nor U22237 (N_22237,N_18781,N_18775);
nor U22238 (N_22238,N_18788,N_18670);
or U22239 (N_22239,N_19616,N_18021);
or U22240 (N_22240,N_18969,N_18080);
nor U22241 (N_22241,N_18747,N_18726);
and U22242 (N_22242,N_19742,N_17665);
nor U22243 (N_22243,N_17524,N_18704);
nand U22244 (N_22244,N_19268,N_18001);
nor U22245 (N_22245,N_17841,N_17998);
or U22246 (N_22246,N_19326,N_19615);
or U22247 (N_22247,N_17857,N_18105);
xnor U22248 (N_22248,N_19536,N_19554);
nor U22249 (N_22249,N_18236,N_19297);
or U22250 (N_22250,N_17732,N_17946);
xnor U22251 (N_22251,N_18455,N_18128);
and U22252 (N_22252,N_18149,N_19761);
nand U22253 (N_22253,N_18699,N_19884);
or U22254 (N_22254,N_18682,N_18191);
nand U22255 (N_22255,N_19248,N_19619);
xnor U22256 (N_22256,N_19991,N_18993);
nand U22257 (N_22257,N_17937,N_19697);
and U22258 (N_22258,N_19324,N_17537);
or U22259 (N_22259,N_18555,N_19202);
nor U22260 (N_22260,N_19825,N_19783);
and U22261 (N_22261,N_19666,N_18365);
nor U22262 (N_22262,N_17773,N_19427);
and U22263 (N_22263,N_19251,N_18164);
or U22264 (N_22264,N_19004,N_17884);
nor U22265 (N_22265,N_18630,N_19491);
or U22266 (N_22266,N_18709,N_19412);
or U22267 (N_22267,N_18166,N_19406);
nand U22268 (N_22268,N_18272,N_18548);
nand U22269 (N_22269,N_19094,N_17854);
nor U22270 (N_22270,N_19697,N_19721);
or U22271 (N_22271,N_18968,N_19740);
and U22272 (N_22272,N_17787,N_17758);
or U22273 (N_22273,N_17946,N_19160);
or U22274 (N_22274,N_18611,N_18933);
nand U22275 (N_22275,N_18801,N_18838);
or U22276 (N_22276,N_18673,N_18137);
nand U22277 (N_22277,N_18406,N_19905);
nand U22278 (N_22278,N_17798,N_19238);
nand U22279 (N_22279,N_19825,N_17900);
nor U22280 (N_22280,N_18785,N_19402);
or U22281 (N_22281,N_17734,N_18630);
or U22282 (N_22282,N_19111,N_18545);
or U22283 (N_22283,N_19461,N_18964);
nand U22284 (N_22284,N_19508,N_17943);
or U22285 (N_22285,N_17855,N_18021);
nor U22286 (N_22286,N_17806,N_19748);
or U22287 (N_22287,N_17738,N_19043);
or U22288 (N_22288,N_18351,N_19853);
or U22289 (N_22289,N_18188,N_18819);
or U22290 (N_22290,N_18751,N_18588);
or U22291 (N_22291,N_18007,N_18369);
nand U22292 (N_22292,N_19786,N_18315);
or U22293 (N_22293,N_18924,N_17637);
nand U22294 (N_22294,N_18748,N_19790);
xor U22295 (N_22295,N_19675,N_18627);
or U22296 (N_22296,N_19040,N_19544);
nand U22297 (N_22297,N_18103,N_19796);
nor U22298 (N_22298,N_18685,N_19800);
and U22299 (N_22299,N_17759,N_17947);
nand U22300 (N_22300,N_18205,N_18970);
nor U22301 (N_22301,N_18846,N_18807);
nand U22302 (N_22302,N_17512,N_17730);
or U22303 (N_22303,N_18010,N_17815);
and U22304 (N_22304,N_18426,N_17609);
and U22305 (N_22305,N_18027,N_19341);
nand U22306 (N_22306,N_17635,N_18742);
nor U22307 (N_22307,N_19556,N_17801);
nand U22308 (N_22308,N_18024,N_19985);
and U22309 (N_22309,N_18402,N_18581);
nor U22310 (N_22310,N_17883,N_18679);
or U22311 (N_22311,N_19865,N_18499);
or U22312 (N_22312,N_19877,N_19963);
and U22313 (N_22313,N_18018,N_19415);
and U22314 (N_22314,N_17591,N_19503);
nand U22315 (N_22315,N_19555,N_19806);
or U22316 (N_22316,N_18746,N_18684);
nand U22317 (N_22317,N_19235,N_19944);
or U22318 (N_22318,N_17701,N_18470);
or U22319 (N_22319,N_18373,N_19469);
and U22320 (N_22320,N_18511,N_17638);
or U22321 (N_22321,N_19474,N_18463);
and U22322 (N_22322,N_17626,N_17543);
and U22323 (N_22323,N_18592,N_18358);
nor U22324 (N_22324,N_19570,N_18008);
and U22325 (N_22325,N_18831,N_19373);
and U22326 (N_22326,N_18322,N_18568);
or U22327 (N_22327,N_18418,N_17911);
nand U22328 (N_22328,N_18345,N_19828);
or U22329 (N_22329,N_17949,N_19470);
nand U22330 (N_22330,N_19792,N_17973);
or U22331 (N_22331,N_19705,N_18110);
nor U22332 (N_22332,N_18927,N_18276);
and U22333 (N_22333,N_18735,N_18249);
or U22334 (N_22334,N_18382,N_17503);
nand U22335 (N_22335,N_18529,N_19902);
nor U22336 (N_22336,N_18533,N_18803);
or U22337 (N_22337,N_18812,N_17979);
nand U22338 (N_22338,N_19886,N_18320);
nor U22339 (N_22339,N_18092,N_17566);
nor U22340 (N_22340,N_18078,N_18879);
xor U22341 (N_22341,N_19990,N_19941);
and U22342 (N_22342,N_18576,N_19977);
nor U22343 (N_22343,N_18267,N_18245);
or U22344 (N_22344,N_17509,N_17602);
or U22345 (N_22345,N_18288,N_18324);
nand U22346 (N_22346,N_18066,N_17935);
nor U22347 (N_22347,N_17780,N_19043);
nor U22348 (N_22348,N_18624,N_18308);
and U22349 (N_22349,N_19467,N_19393);
or U22350 (N_22350,N_18193,N_18028);
nand U22351 (N_22351,N_18197,N_19711);
nand U22352 (N_22352,N_19607,N_17961);
nor U22353 (N_22353,N_18259,N_18979);
nor U22354 (N_22354,N_19068,N_17936);
or U22355 (N_22355,N_19466,N_19341);
nor U22356 (N_22356,N_18237,N_19602);
nor U22357 (N_22357,N_19578,N_18852);
nand U22358 (N_22358,N_17761,N_18715);
or U22359 (N_22359,N_17812,N_18763);
and U22360 (N_22360,N_17512,N_17771);
xor U22361 (N_22361,N_18902,N_19226);
and U22362 (N_22362,N_19583,N_18991);
or U22363 (N_22363,N_19565,N_18388);
and U22364 (N_22364,N_19708,N_18010);
nor U22365 (N_22365,N_19915,N_18220);
and U22366 (N_22366,N_18230,N_18916);
xnor U22367 (N_22367,N_17502,N_18471);
nand U22368 (N_22368,N_19590,N_17793);
nor U22369 (N_22369,N_19742,N_17576);
or U22370 (N_22370,N_18404,N_19380);
nand U22371 (N_22371,N_19389,N_18890);
nand U22372 (N_22372,N_19776,N_17647);
nor U22373 (N_22373,N_19177,N_19391);
nor U22374 (N_22374,N_19291,N_19684);
or U22375 (N_22375,N_17716,N_17807);
and U22376 (N_22376,N_18808,N_19862);
or U22377 (N_22377,N_18783,N_19295);
nand U22378 (N_22378,N_18855,N_18286);
or U22379 (N_22379,N_19295,N_19911);
or U22380 (N_22380,N_19939,N_18581);
nand U22381 (N_22381,N_19084,N_18018);
nor U22382 (N_22382,N_17564,N_17538);
or U22383 (N_22383,N_17782,N_17568);
nand U22384 (N_22384,N_19373,N_18113);
or U22385 (N_22385,N_18389,N_19109);
or U22386 (N_22386,N_19126,N_17809);
nand U22387 (N_22387,N_19936,N_18826);
nor U22388 (N_22388,N_18561,N_19608);
and U22389 (N_22389,N_18203,N_18462);
nand U22390 (N_22390,N_18528,N_19080);
or U22391 (N_22391,N_19382,N_18693);
or U22392 (N_22392,N_17678,N_17939);
or U22393 (N_22393,N_17920,N_19286);
or U22394 (N_22394,N_19072,N_18229);
nand U22395 (N_22395,N_17693,N_18734);
or U22396 (N_22396,N_18287,N_18074);
nor U22397 (N_22397,N_18326,N_18447);
and U22398 (N_22398,N_18438,N_18178);
or U22399 (N_22399,N_19281,N_19656);
or U22400 (N_22400,N_19777,N_18316);
or U22401 (N_22401,N_18059,N_18655);
nor U22402 (N_22402,N_18640,N_18540);
and U22403 (N_22403,N_18875,N_19606);
and U22404 (N_22404,N_19382,N_18346);
or U22405 (N_22405,N_18734,N_18842);
or U22406 (N_22406,N_19409,N_18121);
and U22407 (N_22407,N_19871,N_18340);
nor U22408 (N_22408,N_18751,N_19292);
nor U22409 (N_22409,N_17952,N_18374);
and U22410 (N_22410,N_17567,N_18663);
nor U22411 (N_22411,N_17730,N_18167);
or U22412 (N_22412,N_18553,N_18470);
or U22413 (N_22413,N_18492,N_19019);
nor U22414 (N_22414,N_18626,N_18354);
nor U22415 (N_22415,N_18046,N_19718);
nor U22416 (N_22416,N_19402,N_19690);
nand U22417 (N_22417,N_18601,N_18435);
or U22418 (N_22418,N_18542,N_18255);
nand U22419 (N_22419,N_18606,N_18364);
or U22420 (N_22420,N_17810,N_18397);
and U22421 (N_22421,N_18101,N_17705);
and U22422 (N_22422,N_19072,N_19568);
nand U22423 (N_22423,N_18290,N_19963);
nand U22424 (N_22424,N_18088,N_18473);
and U22425 (N_22425,N_19602,N_19622);
and U22426 (N_22426,N_18531,N_18164);
nor U22427 (N_22427,N_19703,N_17976);
or U22428 (N_22428,N_18530,N_18371);
or U22429 (N_22429,N_18027,N_19966);
nor U22430 (N_22430,N_17581,N_19294);
nand U22431 (N_22431,N_18081,N_17894);
nor U22432 (N_22432,N_17933,N_19467);
nand U22433 (N_22433,N_19326,N_18799);
and U22434 (N_22434,N_17976,N_18659);
or U22435 (N_22435,N_17762,N_19648);
nand U22436 (N_22436,N_18474,N_19482);
or U22437 (N_22437,N_19086,N_18225);
and U22438 (N_22438,N_19191,N_19053);
or U22439 (N_22439,N_19535,N_19015);
nand U22440 (N_22440,N_18087,N_17696);
nor U22441 (N_22441,N_18463,N_18257);
nand U22442 (N_22442,N_19802,N_19026);
or U22443 (N_22443,N_18145,N_18303);
nand U22444 (N_22444,N_19255,N_19191);
nand U22445 (N_22445,N_19921,N_17675);
nor U22446 (N_22446,N_18693,N_19939);
or U22447 (N_22447,N_19769,N_18235);
nor U22448 (N_22448,N_17531,N_17621);
or U22449 (N_22449,N_18759,N_19587);
nand U22450 (N_22450,N_18761,N_18838);
or U22451 (N_22451,N_19502,N_19928);
and U22452 (N_22452,N_19970,N_19438);
and U22453 (N_22453,N_17730,N_18466);
or U22454 (N_22454,N_17629,N_18700);
and U22455 (N_22455,N_19000,N_19916);
nor U22456 (N_22456,N_18235,N_17753);
or U22457 (N_22457,N_19887,N_18050);
and U22458 (N_22458,N_19543,N_19012);
and U22459 (N_22459,N_19378,N_19233);
or U22460 (N_22460,N_18416,N_18215);
nand U22461 (N_22461,N_18339,N_17562);
or U22462 (N_22462,N_18005,N_18599);
nor U22463 (N_22463,N_19430,N_17708);
nand U22464 (N_22464,N_17770,N_18527);
nor U22465 (N_22465,N_18224,N_18028);
nor U22466 (N_22466,N_18067,N_17591);
or U22467 (N_22467,N_17626,N_19898);
xnor U22468 (N_22468,N_17790,N_19179);
nand U22469 (N_22469,N_17763,N_18677);
and U22470 (N_22470,N_19412,N_19282);
nor U22471 (N_22471,N_18940,N_18162);
or U22472 (N_22472,N_17885,N_19815);
nand U22473 (N_22473,N_18542,N_18493);
xnor U22474 (N_22474,N_19543,N_18937);
or U22475 (N_22475,N_17847,N_17694);
nor U22476 (N_22476,N_19009,N_19720);
nor U22477 (N_22477,N_18328,N_18053);
nand U22478 (N_22478,N_19878,N_18350);
or U22479 (N_22479,N_19120,N_18943);
and U22480 (N_22480,N_18293,N_18713);
and U22481 (N_22481,N_17574,N_18330);
and U22482 (N_22482,N_19957,N_19801);
nand U22483 (N_22483,N_18442,N_19295);
nand U22484 (N_22484,N_19195,N_18479);
nand U22485 (N_22485,N_18284,N_18539);
nor U22486 (N_22486,N_17585,N_18579);
and U22487 (N_22487,N_19185,N_19335);
nand U22488 (N_22488,N_19521,N_18922);
nand U22489 (N_22489,N_18580,N_18105);
xor U22490 (N_22490,N_19204,N_19186);
or U22491 (N_22491,N_19712,N_19679);
nand U22492 (N_22492,N_18974,N_18343);
nor U22493 (N_22493,N_19027,N_19802);
and U22494 (N_22494,N_18730,N_18043);
nand U22495 (N_22495,N_19159,N_19319);
nor U22496 (N_22496,N_18988,N_19670);
nor U22497 (N_22497,N_19863,N_19813);
nor U22498 (N_22498,N_19210,N_19385);
and U22499 (N_22499,N_18654,N_18176);
nand U22500 (N_22500,N_21764,N_20165);
nor U22501 (N_22501,N_21772,N_20570);
and U22502 (N_22502,N_21241,N_22326);
nand U22503 (N_22503,N_22375,N_21044);
or U22504 (N_22504,N_20206,N_20171);
and U22505 (N_22505,N_21702,N_22090);
nor U22506 (N_22506,N_22151,N_22488);
or U22507 (N_22507,N_20453,N_22355);
xnor U22508 (N_22508,N_20707,N_20512);
nand U22509 (N_22509,N_20082,N_20429);
nor U22510 (N_22510,N_21838,N_21851);
nor U22511 (N_22511,N_20781,N_20257);
or U22512 (N_22512,N_21275,N_21365);
nor U22513 (N_22513,N_22415,N_22483);
nand U22514 (N_22514,N_20534,N_21587);
nor U22515 (N_22515,N_20648,N_21204);
or U22516 (N_22516,N_20878,N_22149);
and U22517 (N_22517,N_20409,N_21954);
xor U22518 (N_22518,N_21350,N_20536);
nor U22519 (N_22519,N_20988,N_20805);
and U22520 (N_22520,N_21475,N_22263);
nand U22521 (N_22521,N_21928,N_20761);
or U22522 (N_22522,N_20637,N_20765);
nand U22523 (N_22523,N_21456,N_22078);
nor U22524 (N_22524,N_21194,N_20083);
nand U22525 (N_22525,N_20492,N_20321);
nand U22526 (N_22526,N_20775,N_21972);
or U22527 (N_22527,N_20454,N_22373);
and U22528 (N_22528,N_20150,N_20339);
and U22529 (N_22529,N_20399,N_22428);
and U22530 (N_22530,N_21745,N_22133);
nor U22531 (N_22531,N_21289,N_20127);
nor U22532 (N_22532,N_22416,N_20226);
nand U22533 (N_22533,N_20390,N_20588);
or U22534 (N_22534,N_20426,N_20859);
nand U22535 (N_22535,N_21001,N_21542);
and U22536 (N_22536,N_20476,N_21495);
nor U22537 (N_22537,N_21910,N_21812);
and U22538 (N_22538,N_21675,N_20575);
and U22539 (N_22539,N_21138,N_21509);
nor U22540 (N_22540,N_20522,N_20291);
nor U22541 (N_22541,N_21919,N_20465);
nand U22542 (N_22542,N_20269,N_21709);
nand U22543 (N_22543,N_21377,N_21717);
xnor U22544 (N_22544,N_21809,N_20527);
xor U22545 (N_22545,N_22402,N_21940);
or U22546 (N_22546,N_22104,N_21029);
and U22547 (N_22547,N_21452,N_22023);
and U22548 (N_22548,N_21014,N_20743);
and U22549 (N_22549,N_21477,N_22148);
nor U22550 (N_22550,N_21504,N_21166);
nand U22551 (N_22551,N_20351,N_21914);
nor U22552 (N_22552,N_21580,N_21575);
nor U22553 (N_22553,N_22153,N_20687);
nor U22554 (N_22554,N_21213,N_22260);
nand U22555 (N_22555,N_21917,N_21470);
and U22556 (N_22556,N_21943,N_22285);
nor U22557 (N_22557,N_20657,N_20101);
and U22558 (N_22558,N_21376,N_20865);
nor U22559 (N_22559,N_20025,N_22322);
or U22560 (N_22560,N_22164,N_21054);
and U22561 (N_22561,N_20948,N_21212);
nor U22562 (N_22562,N_20879,N_22203);
nand U22563 (N_22563,N_20639,N_21198);
nor U22564 (N_22564,N_20508,N_21546);
nand U22565 (N_22565,N_21332,N_21822);
or U22566 (N_22566,N_21183,N_21251);
or U22567 (N_22567,N_20645,N_20270);
xnor U22568 (N_22568,N_20896,N_21398);
or U22569 (N_22569,N_20461,N_20603);
xor U22570 (N_22570,N_20153,N_21045);
nand U22571 (N_22571,N_20642,N_21506);
nor U22572 (N_22572,N_22396,N_20183);
nor U22573 (N_22573,N_20006,N_20766);
or U22574 (N_22574,N_22468,N_22376);
or U22575 (N_22575,N_20649,N_20477);
nand U22576 (N_22576,N_20413,N_21413);
nand U22577 (N_22577,N_21474,N_22121);
nand U22578 (N_22578,N_22272,N_21424);
and U22579 (N_22579,N_22157,N_21963);
nor U22580 (N_22580,N_20480,N_20528);
nor U22581 (N_22581,N_20679,N_22030);
nor U22582 (N_22582,N_20152,N_22190);
or U22583 (N_22583,N_21069,N_20857);
nor U22584 (N_22584,N_20088,N_22115);
and U22585 (N_22585,N_21711,N_22082);
and U22586 (N_22586,N_20197,N_21967);
or U22587 (N_22587,N_21742,N_22442);
nor U22588 (N_22588,N_20682,N_21946);
xnor U22589 (N_22589,N_20620,N_22014);
or U22590 (N_22590,N_21344,N_21618);
nor U22591 (N_22591,N_21197,N_20013);
or U22592 (N_22592,N_22215,N_22460);
nor U22593 (N_22593,N_21561,N_21545);
nor U22594 (N_22594,N_20439,N_20516);
and U22595 (N_22595,N_21053,N_22039);
and U22596 (N_22596,N_20478,N_20365);
or U22597 (N_22597,N_21143,N_21427);
or U22598 (N_22598,N_21108,N_22245);
and U22599 (N_22599,N_21870,N_20190);
nor U22600 (N_22600,N_21794,N_22498);
nand U22601 (N_22601,N_21719,N_20181);
and U22602 (N_22602,N_22366,N_20387);
nand U22603 (N_22603,N_22231,N_21396);
and U22604 (N_22604,N_21072,N_20920);
nand U22605 (N_22605,N_22024,N_20909);
nor U22606 (N_22606,N_20354,N_20102);
or U22607 (N_22607,N_20033,N_21766);
or U22608 (N_22608,N_21106,N_21521);
and U22609 (N_22609,N_21127,N_20030);
and U22610 (N_22610,N_21923,N_21005);
or U22611 (N_22611,N_20685,N_20322);
nor U22612 (N_22612,N_20227,N_21607);
xor U22613 (N_22613,N_20926,N_20207);
nand U22614 (N_22614,N_20950,N_20959);
or U22615 (N_22615,N_20891,N_21018);
and U22616 (N_22616,N_21681,N_22019);
and U22617 (N_22617,N_22268,N_22292);
and U22618 (N_22618,N_21387,N_21132);
and U22619 (N_22619,N_20955,N_21942);
nor U22620 (N_22620,N_21543,N_21513);
and U22621 (N_22621,N_21278,N_21802);
nand U22622 (N_22622,N_22010,N_20933);
nand U22623 (N_22623,N_21416,N_20061);
and U22624 (N_22624,N_20334,N_21035);
or U22625 (N_22625,N_21592,N_20283);
or U22626 (N_22626,N_21654,N_21899);
nor U22627 (N_22627,N_21911,N_22420);
nor U22628 (N_22628,N_21755,N_20271);
nor U22629 (N_22629,N_20389,N_21983);
and U22630 (N_22630,N_20022,N_21306);
nor U22631 (N_22631,N_22298,N_20814);
nor U22632 (N_22632,N_21757,N_20521);
or U22633 (N_22633,N_20906,N_21276);
and U22634 (N_22634,N_21024,N_20502);
and U22635 (N_22635,N_21091,N_21554);
and U22636 (N_22636,N_22354,N_20046);
and U22637 (N_22637,N_20332,N_20386);
and U22638 (N_22638,N_20633,N_21095);
or U22639 (N_22639,N_20808,N_21872);
nand U22640 (N_22640,N_20259,N_20438);
nor U22641 (N_22641,N_22448,N_21388);
nor U22642 (N_22642,N_22181,N_20418);
or U22643 (N_22643,N_20792,N_22451);
and U22644 (N_22644,N_21989,N_22021);
and U22645 (N_22645,N_21081,N_21968);
or U22646 (N_22646,N_20884,N_20107);
xor U22647 (N_22647,N_21897,N_21234);
nor U22648 (N_22648,N_22032,N_21361);
nor U22649 (N_22649,N_20809,N_22241);
or U22650 (N_22650,N_21084,N_20134);
or U22651 (N_22651,N_20581,N_22387);
and U22652 (N_22652,N_20361,N_20268);
nand U22653 (N_22653,N_22484,N_20703);
or U22654 (N_22654,N_21614,N_21186);
nand U22655 (N_22655,N_22333,N_21130);
and U22656 (N_22656,N_20820,N_21360);
or U22657 (N_22657,N_21218,N_21982);
or U22658 (N_22658,N_22188,N_20932);
and U22659 (N_22659,N_20179,N_20910);
and U22660 (N_22660,N_20652,N_22301);
or U22661 (N_22661,N_21321,N_22206);
or U22662 (N_22662,N_21522,N_22443);
nand U22663 (N_22663,N_22319,N_20585);
or U22664 (N_22664,N_22401,N_20398);
and U22665 (N_22665,N_21668,N_20579);
nor U22666 (N_22666,N_20273,N_22093);
nand U22667 (N_22667,N_21271,N_21334);
nor U22668 (N_22668,N_20331,N_20290);
and U22669 (N_22669,N_21552,N_22105);
nand U22670 (N_22670,N_20989,N_22013);
or U22671 (N_22671,N_20234,N_20772);
nand U22672 (N_22672,N_20677,N_20239);
or U22673 (N_22673,N_21401,N_20155);
nor U22674 (N_22674,N_20482,N_20330);
nor U22675 (N_22675,N_21187,N_22352);
nand U22676 (N_22676,N_20618,N_20385);
nor U22677 (N_22677,N_22386,N_20424);
or U22678 (N_22678,N_21291,N_20366);
and U22679 (N_22679,N_21549,N_22110);
and U22680 (N_22680,N_21754,N_20299);
nand U22681 (N_22681,N_20274,N_21074);
or U22682 (N_22682,N_20975,N_20436);
nand U22683 (N_22683,N_20776,N_21059);
nor U22684 (N_22684,N_21179,N_20136);
nand U22685 (N_22685,N_22187,N_20559);
or U22686 (N_22686,N_21230,N_21013);
nor U22687 (N_22687,N_20256,N_21644);
nor U22688 (N_22688,N_21386,N_21853);
or U22689 (N_22689,N_20411,N_20939);
and U22690 (N_22690,N_22084,N_21655);
nand U22691 (N_22691,N_20035,N_20613);
and U22692 (N_22692,N_21583,N_22380);
and U22693 (N_22693,N_21075,N_21955);
and U22694 (N_22694,N_21400,N_21103);
and U22695 (N_22695,N_22081,N_20539);
and U22696 (N_22696,N_20196,N_20702);
nand U22697 (N_22697,N_21490,N_20786);
nand U22698 (N_22698,N_20208,N_20798);
nor U22699 (N_22699,N_21025,N_20683);
nand U22700 (N_22700,N_20759,N_20376);
xor U22701 (N_22701,N_20310,N_20659);
nand U22702 (N_22702,N_20621,N_22296);
xnor U22703 (N_22703,N_20452,N_22094);
nor U22704 (N_22704,N_22370,N_21993);
xnor U22705 (N_22705,N_20737,N_20060);
and U22706 (N_22706,N_20044,N_21002);
and U22707 (N_22707,N_20333,N_21450);
nand U22708 (N_22708,N_20494,N_21847);
nand U22709 (N_22709,N_21610,N_20565);
nand U22710 (N_22710,N_20953,N_21816);
nor U22711 (N_22711,N_21716,N_22103);
nand U22712 (N_22712,N_20119,N_21805);
nor U22713 (N_22713,N_20889,N_20356);
nand U22714 (N_22714,N_21517,N_22320);
or U22715 (N_22715,N_22139,N_20079);
nand U22716 (N_22716,N_22492,N_22213);
nand U22717 (N_22717,N_21881,N_20089);
and U22718 (N_22718,N_20726,N_22469);
nand U22719 (N_22719,N_21653,N_21038);
nand U22720 (N_22720,N_20839,N_20881);
and U22721 (N_22721,N_22464,N_20734);
xor U22722 (N_22722,N_21265,N_20954);
nand U22723 (N_22723,N_22334,N_22412);
or U22724 (N_22724,N_20610,N_20095);
and U22725 (N_22725,N_22365,N_21544);
or U22726 (N_22726,N_20812,N_22275);
nand U22727 (N_22727,N_20342,N_20294);
and U22728 (N_22728,N_20661,N_21697);
and U22729 (N_22729,N_22053,N_20860);
and U22730 (N_22730,N_21303,N_20093);
and U22731 (N_22731,N_21685,N_22142);
nor U22732 (N_22732,N_22134,N_21737);
or U22733 (N_22733,N_21926,N_21918);
nand U22734 (N_22734,N_20927,N_21227);
and U22735 (N_22735,N_20875,N_21604);
and U22736 (N_22736,N_20225,N_20253);
and U22737 (N_22737,N_20660,N_22225);
or U22738 (N_22738,N_20782,N_21357);
and U22739 (N_22739,N_21185,N_22064);
and U22740 (N_22740,N_20018,N_21161);
xor U22741 (N_22741,N_21100,N_22222);
or U22742 (N_22742,N_20731,N_21732);
nand U22743 (N_22743,N_20084,N_21735);
nor U22744 (N_22744,N_21727,N_21208);
nand U22745 (N_22745,N_20638,N_21432);
nand U22746 (N_22746,N_21393,N_20762);
nand U22747 (N_22747,N_21167,N_21286);
nor U22748 (N_22748,N_22179,N_22490);
or U22749 (N_22749,N_20254,N_20913);
nor U22750 (N_22750,N_21066,N_22284);
or U22751 (N_22751,N_20146,N_22017);
and U22752 (N_22752,N_20946,N_21602);
and U22753 (N_22753,N_20381,N_22259);
nand U22754 (N_22754,N_22098,N_21684);
nor U22755 (N_22755,N_21373,N_21970);
or U22756 (N_22756,N_20192,N_22397);
nor U22757 (N_22757,N_20545,N_22002);
nor U22758 (N_22758,N_21501,N_20251);
and U22759 (N_22759,N_20774,N_21071);
or U22760 (N_22760,N_21703,N_20890);
and U22761 (N_22761,N_21363,N_21534);
nor U22762 (N_22762,N_22199,N_22048);
nand U22763 (N_22763,N_20969,N_20552);
or U22764 (N_22764,N_21086,N_22317);
or U22765 (N_22765,N_22182,N_21219);
nand U22766 (N_22766,N_22453,N_21236);
nor U22767 (N_22767,N_20951,N_21990);
or U22768 (N_22768,N_22161,N_22339);
nor U22769 (N_22769,N_20304,N_20435);
or U22770 (N_22770,N_20573,N_22312);
nor U22771 (N_22771,N_21971,N_21557);
xor U22772 (N_22772,N_21240,N_20612);
and U22773 (N_22773,N_21499,N_20371);
and U22774 (N_22774,N_22118,N_21180);
and U22775 (N_22775,N_22494,N_21665);
and U22776 (N_22776,N_21525,N_20216);
nor U22777 (N_22777,N_22446,N_21154);
or U22778 (N_22778,N_20142,N_20191);
nor U22779 (N_22779,N_20325,N_20846);
and U22780 (N_22780,N_21630,N_21524);
and U22781 (N_22781,N_22129,N_20445);
and U22782 (N_22782,N_22340,N_21451);
and U22783 (N_22783,N_20999,N_21077);
and U22784 (N_22784,N_21886,N_22243);
nor U22785 (N_22785,N_20073,N_21455);
nor U22786 (N_22786,N_20400,N_20056);
nor U22787 (N_22787,N_20275,N_21032);
nor U22788 (N_22788,N_20279,N_20647);
or U22789 (N_22789,N_21620,N_20723);
and U22790 (N_22790,N_20554,N_22462);
nand U22791 (N_22791,N_21173,N_20708);
nand U22792 (N_22792,N_21964,N_22119);
or U22793 (N_22793,N_22455,N_21465);
and U22794 (N_22794,N_21383,N_22085);
and U22795 (N_22795,N_21410,N_21680);
or U22796 (N_22796,N_20384,N_20767);
and U22797 (N_22797,N_21062,N_22141);
or U22798 (N_22798,N_21638,N_21273);
nand U22799 (N_22799,N_22126,N_20748);
nor U22800 (N_22800,N_22324,N_20491);
nand U22801 (N_22801,N_21936,N_21632);
and U22802 (N_22802,N_21298,N_22388);
and U22803 (N_22803,N_22155,N_20962);
or U22804 (N_22804,N_21177,N_20286);
or U22805 (N_22805,N_21891,N_22162);
xor U22806 (N_22806,N_21789,N_20345);
or U22807 (N_22807,N_21245,N_21528);
or U22808 (N_22808,N_20267,N_22228);
nand U22809 (N_22809,N_22108,N_20617);
nand U22810 (N_22810,N_22012,N_20582);
and U22811 (N_22811,N_21503,N_20222);
and U22812 (N_22812,N_20729,N_20223);
or U22813 (N_22813,N_20866,N_21479);
nor U22814 (N_22814,N_20770,N_22174);
nor U22815 (N_22815,N_22414,N_21651);
and U22816 (N_22816,N_21340,N_22005);
nor U22817 (N_22817,N_20066,N_20580);
and U22818 (N_22818,N_22248,N_22276);
and U22819 (N_22819,N_21857,N_20212);
and U22820 (N_22820,N_21950,N_21908);
and U22821 (N_22821,N_20576,N_21786);
or U22822 (N_22822,N_22237,N_22261);
nor U22823 (N_22823,N_21048,N_20903);
or U22824 (N_22824,N_21078,N_21803);
nand U22825 (N_22825,N_20616,N_21027);
and U22826 (N_22826,N_20769,N_20180);
xor U22827 (N_22827,N_22309,N_20308);
nor U22828 (N_22828,N_21573,N_21055);
or U22829 (N_22829,N_22434,N_20763);
nor U22830 (N_22830,N_20777,N_20547);
or U22831 (N_22831,N_22267,N_22156);
nor U22832 (N_22832,N_21242,N_21641);
and U22833 (N_22833,N_21196,N_20824);
or U22834 (N_22834,N_21738,N_22191);
nor U22835 (N_22835,N_20867,N_20727);
or U22836 (N_22836,N_22158,N_20701);
nand U22837 (N_22837,N_20673,N_20740);
or U22838 (N_22838,N_21496,N_20757);
nand U22839 (N_22839,N_22229,N_21418);
nand U22840 (N_22840,N_20540,N_20758);
nor U22841 (N_22841,N_21122,N_21346);
or U22842 (N_22842,N_21415,N_22257);
or U22843 (N_22843,N_22106,N_21028);
or U22844 (N_22844,N_20276,N_21026);
nor U22845 (N_22845,N_22286,N_21800);
nor U22846 (N_22846,N_20650,N_22058);
nand U22847 (N_22847,N_20607,N_20432);
nor U22848 (N_22848,N_21671,N_22264);
nor U22849 (N_22849,N_20998,N_21611);
or U22850 (N_22850,N_22391,N_22424);
and U22851 (N_22851,N_20104,N_22236);
nor U22852 (N_22852,N_22196,N_21156);
nor U22853 (N_22853,N_21713,N_20029);
nor U22854 (N_22854,N_22258,N_21389);
nand U22855 (N_22855,N_20122,N_20052);
nor U22856 (N_22856,N_21486,N_21831);
and U22857 (N_22857,N_20898,N_20821);
nor U22858 (N_22858,N_20312,N_20721);
nand U22859 (N_22859,N_21258,N_21436);
and U22860 (N_22860,N_21070,N_20346);
nand U22861 (N_22861,N_21660,N_22266);
nand U22862 (N_22862,N_20041,N_20097);
nand U22863 (N_22863,N_20656,N_21850);
and U22864 (N_22864,N_20853,N_20979);
and U22865 (N_22865,N_21047,N_21994);
and U22866 (N_22866,N_21201,N_20460);
nor U22867 (N_22867,N_20714,N_20094);
nor U22868 (N_22868,N_21579,N_20086);
nor U22869 (N_22869,N_20340,N_20374);
nor U22870 (N_22870,N_21590,N_21426);
nor U22871 (N_22871,N_20861,N_21707);
nand U22872 (N_22872,N_22122,N_20965);
or U22873 (N_22873,N_21746,N_21814);
nand U22874 (N_22874,N_20362,N_21763);
and U22875 (N_22875,N_20943,N_22150);
and U22876 (N_22876,N_21445,N_21876);
and U22877 (N_22877,N_21372,N_21625);
and U22878 (N_22878,N_21462,N_21570);
or U22879 (N_22879,N_22439,N_21049);
and U22880 (N_22880,N_20530,N_21058);
nor U22881 (N_22881,N_20092,N_20796);
or U22882 (N_22882,N_22463,N_21793);
nand U22883 (N_22883,N_21532,N_22130);
nor U22884 (N_22884,N_22389,N_21003);
or U22885 (N_22885,N_20684,N_21798);
and U22886 (N_22886,N_21336,N_20912);
nor U22887 (N_22887,N_22102,N_20420);
and U22888 (N_22888,N_21297,N_21243);
nor U22889 (N_22889,N_21293,N_21852);
or U22890 (N_22890,N_21951,N_20490);
nor U22891 (N_22891,N_20944,N_22152);
nand U22892 (N_22892,N_22069,N_21898);
nor U22893 (N_22893,N_20428,N_21502);
nor U22894 (N_22894,N_21082,N_21520);
nor U22895 (N_22895,N_21778,N_22440);
or U22896 (N_22896,N_21998,N_20990);
and U22897 (N_22897,N_22087,N_20973);
nor U22898 (N_22898,N_20382,N_21237);
nand U22899 (N_22899,N_22478,N_20319);
nand U22900 (N_22900,N_20303,N_20817);
and U22901 (N_22901,N_21715,N_22088);
nor U22902 (N_22902,N_22323,N_20836);
or U22903 (N_22903,N_20693,N_21006);
nor U22904 (N_22904,N_21974,N_22390);
nor U22905 (N_22905,N_20031,N_20811);
or U22906 (N_22906,N_20591,N_22120);
or U22907 (N_22907,N_22057,N_20247);
xnor U22908 (N_22908,N_21113,N_22381);
or U22909 (N_22909,N_21818,N_20038);
or U22910 (N_22910,N_20100,N_22417);
nand U22911 (N_22911,N_21959,N_21080);
nor U22912 (N_22912,N_20916,N_20543);
or U22913 (N_22913,N_20558,N_22481);
nor U22914 (N_22914,N_21762,N_21957);
and U22915 (N_22915,N_21616,N_21174);
and U22916 (N_22916,N_21043,N_20444);
nand U22917 (N_22917,N_21435,N_21679);
nor U22918 (N_22918,N_21394,N_21839);
or U22919 (N_22919,N_22350,N_22249);
or U22920 (N_22920,N_22337,N_22230);
nand U22921 (N_22921,N_21461,N_21466);
or U22922 (N_22922,N_20634,N_22368);
nor U22923 (N_22923,N_20905,N_21861);
nand U22924 (N_22924,N_20040,N_22270);
nor U22925 (N_22925,N_21832,N_22227);
nand U22926 (N_22926,N_20689,N_22006);
and U22927 (N_22927,N_20285,N_20473);
or U22928 (N_22928,N_20474,N_21663);
nand U22929 (N_22929,N_20507,N_20574);
or U22930 (N_22930,N_22111,N_20406);
nor U22931 (N_22931,N_20895,N_20495);
nor U22932 (N_22932,N_22208,N_21041);
nand U22933 (N_22933,N_21965,N_22459);
nand U22934 (N_22934,N_20615,N_20974);
nand U22935 (N_22935,N_20221,N_22290);
nor U22936 (N_22936,N_21345,N_21257);
nand U22937 (N_22937,N_21391,N_20952);
or U22938 (N_22938,N_20200,N_21514);
or U22939 (N_22939,N_21912,N_20442);
nor U22940 (N_22940,N_20166,N_20768);
nor U22941 (N_22941,N_22144,N_21341);
nand U22942 (N_22942,N_20497,N_21781);
or U22943 (N_22943,N_21252,N_21149);
nand U22944 (N_22944,N_21145,N_22426);
nand U22945 (N_22945,N_21307,N_21981);
and U22946 (N_22946,N_20725,N_20015);
nor U22947 (N_22947,N_21266,N_21615);
nor U22948 (N_22948,N_21986,N_21817);
nand U22949 (N_22949,N_22168,N_20320);
nand U22950 (N_22950,N_21352,N_21358);
nand U22951 (N_22951,N_20967,N_21153);
nand U22952 (N_22952,N_21168,N_22033);
xnor U22953 (N_22953,N_20577,N_22167);
or U22954 (N_22954,N_21869,N_21433);
nor U22955 (N_22955,N_20280,N_21191);
nand U22956 (N_22956,N_20446,N_21808);
or U22957 (N_22957,N_20728,N_20121);
nand U22958 (N_22958,N_21566,N_21748);
nor U22959 (N_22959,N_20544,N_22177);
nor U22960 (N_22960,N_21728,N_22399);
and U22961 (N_22961,N_21217,N_20338);
and U22962 (N_22962,N_21449,N_21395);
nand U22963 (N_22963,N_21308,N_21444);
nand U22964 (N_22964,N_21639,N_21938);
nand U22965 (N_22965,N_20897,N_20976);
and U22966 (N_22966,N_20670,N_21067);
and U22967 (N_22967,N_20997,N_20441);
nor U22968 (N_22968,N_20403,N_20594);
or U22969 (N_22969,N_21210,N_21051);
and U22970 (N_22970,N_21821,N_21152);
xnor U22971 (N_22971,N_20605,N_20901);
nand U22972 (N_22972,N_20626,N_20855);
or U22973 (N_22973,N_20827,N_21841);
nand U22974 (N_22974,N_20224,N_20245);
nand U22975 (N_22975,N_22071,N_22178);
nor U22976 (N_22976,N_21550,N_21825);
nand U22977 (N_22977,N_21840,N_22445);
or U22978 (N_22978,N_21612,N_20675);
and U22979 (N_22979,N_21439,N_21696);
xnor U22980 (N_22980,N_22049,N_22479);
nor U22981 (N_22981,N_22305,N_21259);
and U22982 (N_22982,N_22099,N_20189);
or U22983 (N_22983,N_20471,N_21211);
and U22984 (N_22984,N_21087,N_21126);
nand U22985 (N_22985,N_20260,N_21313);
nand U22986 (N_22986,N_22351,N_21978);
nor U22987 (N_22987,N_22422,N_21662);
nor U22988 (N_22988,N_20489,N_20947);
or U22989 (N_22989,N_22018,N_20807);
or U22990 (N_22990,N_20793,N_22274);
nand U22991 (N_22991,N_21000,N_22100);
and U22992 (N_22992,N_21617,N_21867);
and U22993 (N_22993,N_21235,N_20087);
nor U22994 (N_22994,N_20614,N_20185);
or U22995 (N_22995,N_22255,N_21116);
or U22996 (N_22996,N_20364,N_20911);
nor U22997 (N_22997,N_21141,N_20694);
nor U22998 (N_22998,N_21699,N_21548);
nand U22999 (N_22999,N_22065,N_20862);
or U23000 (N_23000,N_20300,N_20131);
and U23001 (N_23001,N_20314,N_20210);
nor U23002 (N_23002,N_21353,N_20369);
and U23003 (N_23003,N_21609,N_21626);
and U23004 (N_23004,N_20417,N_20732);
nand U23005 (N_23005,N_22467,N_21385);
nand U23006 (N_23006,N_20627,N_21860);
nand U23007 (N_23007,N_20870,N_21979);
or U23008 (N_23008,N_21635,N_21464);
nand U23009 (N_23009,N_22450,N_21761);
nor U23010 (N_23010,N_21325,N_20204);
and U23011 (N_23011,N_21163,N_20880);
xor U23012 (N_23012,N_22477,N_20449);
xor U23013 (N_23013,N_21589,N_22154);
nor U23014 (N_23014,N_20803,N_21057);
or U23015 (N_23015,N_21354,N_20598);
nand U23016 (N_23016,N_20872,N_22097);
or U23017 (N_23017,N_20391,N_20572);
nand U23018 (N_23018,N_21232,N_21999);
nand U23019 (N_23019,N_22316,N_21581);
nand U23020 (N_23020,N_20397,N_20858);
nor U23021 (N_23021,N_20109,N_21190);
or U23022 (N_23022,N_21342,N_20281);
nand U23023 (N_23023,N_22204,N_20681);
nand U23024 (N_23024,N_20178,N_20934);
nor U23025 (N_23025,N_20347,N_21007);
and U23026 (N_23026,N_20704,N_21689);
or U23027 (N_23027,N_20986,N_20981);
nor U23028 (N_23028,N_21046,N_20835);
and U23029 (N_23029,N_20408,N_22047);
nor U23030 (N_23030,N_21958,N_20505);
nor U23031 (N_23031,N_21135,N_21249);
and U23032 (N_23032,N_21011,N_20311);
nor U23033 (N_23033,N_20549,N_20550);
and U23034 (N_23034,N_20466,N_20590);
and U23035 (N_23035,N_21323,N_22140);
nand U23036 (N_23036,N_22482,N_21019);
nand U23037 (N_23037,N_20050,N_21537);
and U23038 (N_23038,N_22089,N_20970);
nor U23039 (N_23039,N_22195,N_21442);
nand U23040 (N_23040,N_22232,N_20583);
or U23041 (N_23041,N_20678,N_20546);
nor U23042 (N_23042,N_20713,N_22233);
or U23043 (N_23043,N_20700,N_22055);
and U23044 (N_23044,N_20838,N_21843);
and U23045 (N_23045,N_21221,N_22076);
nand U23046 (N_23046,N_20506,N_21533);
nand U23047 (N_23047,N_20562,N_21902);
nor U23048 (N_23048,N_20026,N_22487);
and U23049 (N_23049,N_22393,N_20323);
nand U23050 (N_23050,N_21759,N_20057);
nor U23051 (N_23051,N_21770,N_21726);
and U23052 (N_23052,N_22454,N_21247);
nand U23053 (N_23053,N_20653,N_22136);
nand U23054 (N_23054,N_20161,N_21628);
or U23055 (N_23055,N_21417,N_21368);
nand U23056 (N_23056,N_21312,N_20915);
xnor U23057 (N_23057,N_20163,N_22080);
and U23058 (N_23058,N_20455,N_20004);
or U23059 (N_23059,N_20054,N_22475);
nor U23060 (N_23060,N_20388,N_21226);
nand U23061 (N_23061,N_22359,N_20359);
or U23062 (N_23062,N_20848,N_21233);
nand U23063 (N_23063,N_22034,N_20894);
nand U23064 (N_23064,N_21110,N_22300);
nor U23065 (N_23065,N_21686,N_20600);
xor U23066 (N_23066,N_21379,N_20813);
xnor U23067 (N_23067,N_21228,N_22205);
nand U23068 (N_23068,N_21599,N_21131);
nor U23069 (N_23069,N_21892,N_20779);
and U23070 (N_23070,N_22293,N_21050);
or U23071 (N_23071,N_20085,N_20075);
nor U23072 (N_23072,N_20199,N_21409);
nor U23073 (N_23073,N_21865,N_20914);
and U23074 (N_23074,N_22246,N_20167);
and U23075 (N_23075,N_22287,N_21578);
and U23076 (N_23076,N_21718,N_22360);
nand U23077 (N_23077,N_21795,N_20394);
nor U23078 (N_23078,N_21317,N_21371);
nor U23079 (N_23079,N_21913,N_21901);
nand U23080 (N_23080,N_21670,N_21292);
or U23081 (N_23081,N_20194,N_21536);
or U23082 (N_23082,N_21244,N_20863);
and U23083 (N_23083,N_22138,N_21915);
nand U23084 (N_23084,N_21052,N_20175);
or U23085 (N_23085,N_21034,N_20368);
nand U23086 (N_23086,N_21682,N_20416);
nor U23087 (N_23087,N_21073,N_20141);
nor U23088 (N_23088,N_22433,N_22452);
and U23089 (N_23089,N_20592,N_21176);
or U23090 (N_23090,N_20096,N_20071);
or U23091 (N_23091,N_20309,N_21255);
xnor U23092 (N_23092,N_20023,N_21125);
nand U23093 (N_23093,N_21659,N_22344);
nand U23094 (N_23094,N_21600,N_20238);
nor U23095 (N_23095,N_21281,N_20149);
or U23096 (N_23096,N_20511,N_22457);
and U23097 (N_23097,N_21160,N_21030);
and U23098 (N_23098,N_21692,N_21721);
nand U23099 (N_23099,N_20597,N_20919);
nand U23100 (N_23100,N_21678,N_20978);
or U23101 (N_23101,N_20968,N_21402);
and U23102 (N_23102,N_21667,N_20992);
nor U23103 (N_23103,N_20090,N_22137);
nor U23104 (N_23104,N_22436,N_20504);
nand U23105 (N_23105,N_21669,N_20077);
or U23106 (N_23106,N_21320,N_22371);
nand U23107 (N_23107,N_20784,N_20789);
nand U23108 (N_23108,N_21136,N_21494);
nor U23109 (N_23109,N_21791,N_22273);
nor U23110 (N_23110,N_20991,N_21586);
nand U23111 (N_23111,N_20818,N_21594);
xor U23112 (N_23112,N_21920,N_22165);
nor U23113 (N_23113,N_21905,N_21937);
or U23114 (N_23114,N_21165,N_20712);
nor U23115 (N_23115,N_20201,N_21288);
and U23116 (N_23116,N_20885,N_20644);
and U23117 (N_23117,N_20135,N_22183);
xor U23118 (N_23118,N_21128,N_22423);
nand U23119 (N_23119,N_21622,N_20377);
or U23120 (N_23120,N_21890,N_22295);
or U23121 (N_23121,N_21567,N_22435);
nand U23122 (N_23122,N_22146,N_20787);
nor U23123 (N_23123,N_21205,N_20106);
or U23124 (N_23124,N_21294,N_20569);
or U23125 (N_23125,N_21144,N_21150);
and U23126 (N_23126,N_22395,N_20401);
nor U23127 (N_23127,N_20568,N_20187);
nand U23128 (N_23128,N_20070,N_20523);
or U23129 (N_23129,N_22444,N_22353);
and U23130 (N_23130,N_22040,N_20561);
nor U23131 (N_23131,N_20663,N_21079);
nand U23132 (N_23132,N_20350,N_22114);
nor U23133 (N_23133,N_22252,N_22335);
nand U23134 (N_23134,N_21523,N_21478);
or U23135 (N_23135,N_22331,N_21756);
and U23136 (N_23136,N_21904,N_21374);
nand U23137 (N_23137,N_21500,N_21023);
and U23138 (N_23138,N_22280,N_21806);
nor U23139 (N_23139,N_21493,N_21744);
nand U23140 (N_23140,N_21343,N_21991);
or U23141 (N_23141,N_20519,N_21774);
nor U23142 (N_23142,N_21491,N_20353);
nor U23143 (N_23143,N_20414,N_22117);
and U23144 (N_23144,N_21751,N_22091);
nand U23145 (N_23145,N_21314,N_21253);
or U23146 (N_23146,N_20984,N_20336);
nand U23147 (N_23147,N_21516,N_20037);
nor U23148 (N_23148,N_21560,N_20921);
nand U23149 (N_23149,N_20963,N_20631);
nand U23150 (N_23150,N_22035,N_20722);
and U23151 (N_23151,N_20329,N_22083);
nand U23152 (N_23152,N_21568,N_20738);
xnor U23153 (N_23153,N_22250,N_20503);
nand U23154 (N_23154,N_20177,N_20904);
or U23155 (N_23155,N_21004,N_22438);
or U23156 (N_23156,N_20602,N_21220);
nor U23157 (N_23157,N_22011,N_20526);
nand U23158 (N_23158,N_21677,N_20541);
nand U23159 (N_23159,N_22224,N_21181);
and U23160 (N_23160,N_22383,N_21944);
nand U23161 (N_23161,N_20012,N_20868);
nor U23162 (N_23162,N_20448,N_21975);
or U23163 (N_23163,N_20458,N_21823);
nand U23164 (N_23164,N_21691,N_22303);
xnor U23165 (N_23165,N_21629,N_21339);
or U23166 (N_23166,N_21169,N_20484);
or U23167 (N_23167,N_20629,N_21810);
nand U23168 (N_23168,N_21296,N_20343);
or U23169 (N_23169,N_20646,N_21907);
nand U23170 (N_23170,N_20126,N_21956);
or U23171 (N_23171,N_22147,N_21420);
nor U23172 (N_23172,N_20518,N_21784);
or U23173 (N_23173,N_21118,N_21338);
nor U23174 (N_23174,N_22214,N_21083);
nand U23175 (N_23175,N_21571,N_21743);
nor U23176 (N_23176,N_20972,N_21489);
or U23177 (N_23177,N_21710,N_20427);
nand U23178 (N_23178,N_22074,N_20469);
and U23179 (N_23179,N_22473,N_20778);
or U23180 (N_23180,N_21063,N_20593);
and U23181 (N_23181,N_22029,N_20900);
or U23182 (N_23182,N_21666,N_22349);
nand U23183 (N_23183,N_21515,N_21022);
nor U23184 (N_23184,N_22302,N_21819);
nor U23185 (N_23185,N_20669,N_20829);
or U23186 (N_23186,N_20249,N_20295);
and U23187 (N_23187,N_22095,N_20118);
and U23188 (N_23188,N_20211,N_20856);
or U23189 (N_23189,N_21268,N_20542);
or U23190 (N_23190,N_21064,N_20942);
nor U23191 (N_23191,N_20983,N_22374);
xnor U23192 (N_23192,N_21894,N_21563);
xor U23193 (N_23193,N_21598,N_21422);
or U23194 (N_23194,N_21969,N_21895);
and U23195 (N_23195,N_20899,N_21932);
nor U23196 (N_23196,N_21159,N_22194);
nand U23197 (N_23197,N_21855,N_22015);
or U23198 (N_23198,N_21285,N_20114);
nor U23199 (N_23199,N_20832,N_20667);
and U23200 (N_23200,N_21790,N_22432);
nor U23201 (N_23201,N_21705,N_21142);
nand U23202 (N_23202,N_22184,N_20760);
and U23203 (N_23203,N_21572,N_22127);
or U23204 (N_23204,N_22458,N_20849);
nand U23205 (N_23205,N_20560,N_21114);
nand U23206 (N_23206,N_20993,N_21207);
or U23207 (N_23207,N_21621,N_22086);
or U23208 (N_23208,N_21508,N_20804);
and U23209 (N_23209,N_22345,N_21845);
nand U23210 (N_23210,N_22466,N_21813);
nand U23211 (N_23211,N_21785,N_20078);
and U23212 (N_23212,N_21170,N_20363);
and U23213 (N_23213,N_20019,N_21104);
or U23214 (N_23214,N_20302,N_21085);
or U23215 (N_23215,N_22346,N_20823);
nor U23216 (N_23216,N_20831,N_21484);
nor U23217 (N_23217,N_22400,N_22363);
and U23218 (N_23218,N_20780,N_22409);
nor U23219 (N_23219,N_21124,N_21076);
or U23220 (N_23220,N_21333,N_21574);
nor U23221 (N_23221,N_20372,N_21555);
nor U23222 (N_23222,N_22398,N_21985);
or U23223 (N_23223,N_21133,N_21569);
nand U23224 (N_23224,N_20241,N_20801);
and U23225 (N_23225,N_22437,N_21846);
and U23226 (N_23226,N_20869,N_20407);
nand U23227 (N_23227,N_20024,N_20799);
or U23228 (N_23228,N_20451,N_20845);
nand U23229 (N_23229,N_22170,N_20058);
nor U23230 (N_23230,N_21378,N_21779);
nor U23231 (N_23231,N_22025,N_20067);
or U23232 (N_23232,N_20883,N_21767);
nor U23233 (N_23233,N_21068,N_22211);
xor U23234 (N_23234,N_21878,N_20537);
and U23235 (N_23235,N_20488,N_22429);
and U23236 (N_23236,N_20834,N_20360);
nor U23237 (N_23237,N_20016,N_20318);
nand U23238 (N_23238,N_21200,N_20005);
nor U23239 (N_23239,N_21337,N_21434);
nor U23240 (N_23240,N_21636,N_20794);
nor U23241 (N_23241,N_21272,N_20754);
or U23242 (N_23242,N_20143,N_21708);
nand U23243 (N_23243,N_22471,N_21277);
nand U23244 (N_23244,N_22369,N_22308);
nor U23245 (N_23245,N_21105,N_20434);
nand U23246 (N_23246,N_20771,N_20719);
or U23247 (N_23247,N_20624,N_21884);
nor U23248 (N_23248,N_20720,N_21601);
xor U23249 (N_23249,N_21061,N_20138);
nor U23250 (N_23250,N_21299,N_22066);
nand U23251 (N_23251,N_22404,N_20810);
or U23252 (N_23252,N_22289,N_21408);
nor U23253 (N_23253,N_21295,N_21239);
nor U23254 (N_23254,N_20940,N_20440);
and U23255 (N_23255,N_21658,N_20463);
nor U23256 (N_23256,N_20039,N_21214);
or U23257 (N_23257,N_22031,N_20532);
nor U23258 (N_23258,N_21270,N_20011);
or U23259 (N_23259,N_21541,N_20929);
nand U23260 (N_23260,N_20316,N_21423);
nor U23261 (N_23261,N_20850,N_21164);
or U23262 (N_23262,N_21787,N_22410);
nand U23263 (N_23263,N_20217,N_20640);
nor U23264 (N_23264,N_21868,N_21929);
and U23265 (N_23265,N_20945,N_21414);
nand U23266 (N_23266,N_20065,N_21858);
nand U23267 (N_23267,N_21538,N_22343);
or U23268 (N_23268,N_20557,N_20010);
and U23269 (N_23269,N_21290,N_21556);
nor U23270 (N_23270,N_22009,N_21182);
or U23271 (N_23271,N_22051,N_22077);
or U23272 (N_23272,N_20213,N_22262);
or U23273 (N_23273,N_20628,N_21369);
nand U23274 (N_23274,N_20055,N_21010);
nand U23275 (N_23275,N_20064,N_21792);
nand U23276 (N_23276,N_20587,N_20292);
xnor U23277 (N_23277,N_20139,N_21056);
or U23278 (N_23278,N_21796,N_22406);
or U23279 (N_23279,N_20162,N_22041);
nand U23280 (N_23280,N_20844,N_21348);
or U23281 (N_23281,N_21246,N_21775);
and U23282 (N_23282,N_20699,N_20563);
nor U23283 (N_23283,N_21828,N_20147);
nand U23284 (N_23284,N_20985,N_22413);
and U23285 (N_23285,N_20802,N_21765);
nand U23286 (N_23286,N_20243,N_20184);
nand U23287 (N_23287,N_21009,N_20140);
or U23288 (N_23288,N_21603,N_21760);
or U23289 (N_23289,N_21585,N_20924);
or U23290 (N_23290,N_20000,N_20873);
nor U23291 (N_23291,N_21146,N_20806);
nand U23292 (N_23292,N_21037,N_22425);
or U23293 (N_23293,N_20971,N_21238);
nand U23294 (N_23294,N_20378,N_22008);
xor U23295 (N_23295,N_21797,N_22016);
or U23296 (N_23296,N_21987,N_20043);
and U23297 (N_23297,N_20589,N_21996);
or U23298 (N_23298,N_20373,N_20611);
or U23299 (N_23299,N_20773,N_21324);
nor U23300 (N_23300,N_20672,N_20170);
nor U23301 (N_23301,N_21656,N_20284);
nand U23302 (N_23302,N_22427,N_20326);
nand U23303 (N_23303,N_21305,N_21367);
nor U23304 (N_23304,N_20159,N_20186);
nand U23305 (N_23305,N_22221,N_21935);
nand U23306 (N_23306,N_20893,N_21948);
xor U23307 (N_23307,N_20108,N_22474);
nor U23308 (N_23308,N_22306,N_21284);
or U23309 (N_23309,N_21482,N_21750);
or U23310 (N_23310,N_21193,N_20262);
nand U23311 (N_23311,N_20529,N_22062);
nor U23312 (N_23312,N_21042,N_20742);
or U23313 (N_23313,N_22201,N_20051);
nor U23314 (N_23314,N_22038,N_22052);
and U23315 (N_23315,N_21883,N_21216);
nand U23316 (N_23316,N_21390,N_20567);
and U23317 (N_23317,N_20375,N_22456);
nand U23318 (N_23318,N_20531,N_21203);
nor U23319 (N_23319,N_20958,N_21351);
xor U23320 (N_23320,N_22159,N_21833);
nor U23321 (N_23321,N_20876,N_20132);
nand U23322 (N_23322,N_20111,N_20553);
nor U23323 (N_23323,N_21844,N_20240);
and U23324 (N_23324,N_20242,N_22271);
nor U23325 (N_23325,N_21224,N_20715);
nor U23326 (N_23326,N_20887,N_20129);
and U23327 (N_23327,N_22004,N_21137);
nor U23328 (N_23328,N_20063,N_21540);
and U23329 (N_23329,N_21526,N_20125);
nand U23330 (N_23330,N_20133,N_21776);
or U23331 (N_23331,N_21837,N_21316);
and U23332 (N_23332,N_20357,N_20961);
and U23333 (N_23333,N_20515,N_20641);
nor U23334 (N_23334,N_21468,N_20313);
or U23335 (N_23335,N_20696,N_21488);
nor U23336 (N_23336,N_21438,N_22315);
or U23337 (N_23337,N_22378,N_21673);
and U23338 (N_23338,N_21199,N_21527);
and U23339 (N_23339,N_20623,N_22046);
or U23340 (N_23340,N_21109,N_20233);
and U23341 (N_23341,N_21157,N_20795);
nor U23342 (N_23342,N_20745,N_21263);
nand U23343 (N_23343,N_20479,N_20908);
or U23344 (N_23344,N_20697,N_21657);
and U23345 (N_23345,N_21683,N_20468);
and U23346 (N_23346,N_20716,N_21896);
and U23347 (N_23347,N_22348,N_21172);
and U23348 (N_23348,N_22364,N_20520);
and U23349 (N_23349,N_21262,N_20499);
nand U23350 (N_23350,N_20741,N_21382);
nor U23351 (N_23351,N_21741,N_22001);
or U23352 (N_23352,N_22327,N_20380);
nand U23353 (N_23353,N_20724,N_21301);
nor U23354 (N_23354,N_21722,N_21094);
xor U23355 (N_23355,N_20680,N_21849);
or U23356 (N_23356,N_21827,N_20785);
xor U23357 (N_23357,N_21623,N_22042);
and U23358 (N_23358,N_20358,N_21752);
and U23359 (N_23359,N_20501,N_21873);
or U23360 (N_23360,N_20493,N_20710);
and U23361 (N_23361,N_21577,N_21953);
and U23362 (N_23362,N_22318,N_21460);
nor U23363 (N_23363,N_21997,N_21866);
and U23364 (N_23364,N_21158,N_20062);
and U23365 (N_23365,N_20324,N_22247);
nor U23366 (N_23366,N_21411,N_22028);
nand U23367 (N_23367,N_20996,N_21101);
and U23368 (N_23368,N_20533,N_21694);
nand U23369 (N_23369,N_22357,N_21147);
nor U23370 (N_23370,N_22160,N_21097);
and U23371 (N_23371,N_21425,N_20747);
nor U23372 (N_23372,N_21151,N_20852);
nor U23373 (N_23373,N_22314,N_20415);
and U23374 (N_23374,N_20500,N_20158);
or U23375 (N_23375,N_21099,N_21631);
and U23376 (N_23376,N_22283,N_22476);
or U23377 (N_23377,N_21723,N_22254);
nand U23378 (N_23378,N_20513,N_21282);
or U23379 (N_23379,N_22265,N_22499);
nand U23380 (N_23380,N_20496,N_21647);
nand U23381 (N_23381,N_20764,N_20888);
nand U23382 (N_23382,N_22311,N_21676);
nor U23383 (N_23383,N_21347,N_21753);
and U23384 (N_23384,N_20625,N_20327);
nor U23385 (N_23385,N_22486,N_21264);
nand U23386 (N_23386,N_21859,N_21310);
nor U23387 (N_23387,N_21961,N_20431);
nor U23388 (N_23388,N_21962,N_22385);
and U23389 (N_23389,N_21714,N_21498);
nand U23390 (N_23390,N_20049,N_21693);
or U23391 (N_23391,N_22125,N_21529);
or U23392 (N_23392,N_20752,N_20941);
or U23393 (N_23393,N_20666,N_20396);
or U23394 (N_23394,N_21088,N_20036);
and U23395 (N_23395,N_20105,N_21463);
nor U23396 (N_23396,N_21405,N_21331);
xor U23397 (N_23397,N_20877,N_21565);
or U23398 (N_23398,N_21931,N_21637);
xor U23399 (N_23399,N_21980,N_21909);
nand U23400 (N_23400,N_20918,N_20822);
nor U23401 (N_23401,N_20851,N_20705);
xnor U23402 (N_23402,N_21215,N_22128);
or U23403 (N_23403,N_20535,N_20596);
nor U23404 (N_23404,N_20665,N_22379);
and U23405 (N_23405,N_21017,N_20053);
nor U23406 (N_23406,N_22169,N_21349);
nand U23407 (N_23407,N_22092,N_21412);
or U23408 (N_23408,N_21421,N_21206);
nand U23409 (N_23409,N_20826,N_22176);
nor U23410 (N_23410,N_21223,N_20636);
nor U23411 (N_23411,N_21734,N_21992);
nand U23412 (N_23412,N_20551,N_20601);
and U23413 (N_23413,N_20828,N_22166);
and U23414 (N_23414,N_21815,N_20068);
nor U23415 (N_23415,N_20658,N_21469);
nor U23416 (N_23416,N_20571,N_21175);
nand U23417 (N_23417,N_21769,N_20555);
nor U23418 (N_23418,N_21329,N_22496);
nor U23419 (N_23419,N_20115,N_22328);
nand U23420 (N_23420,N_20252,N_20966);
nor U23421 (N_23421,N_21916,N_20790);
nand U23422 (N_23422,N_22362,N_20739);
and U23423 (N_23423,N_21862,N_20841);
nor U23424 (N_23424,N_21877,N_22238);
nor U23425 (N_23425,N_20457,N_20246);
nor U23426 (N_23426,N_20791,N_22491);
nand U23427 (N_23427,N_21829,N_20112);
nor U23428 (N_23428,N_21875,N_22411);
nor U23429 (N_23429,N_21446,N_21758);
nand U23430 (N_23430,N_21712,N_21039);
xnor U23431 (N_23431,N_20709,N_20176);
nor U23432 (N_23432,N_20156,N_22493);
nand U23433 (N_23433,N_22185,N_21888);
nor U23434 (N_23434,N_22253,N_21661);
nand U23435 (N_23435,N_21140,N_21749);
and U23436 (N_23436,N_20045,N_21804);
or U23437 (N_23437,N_21364,N_21531);
and U23438 (N_23438,N_21854,N_21093);
nand U23439 (N_23439,N_20218,N_21553);
and U23440 (N_23440,N_22135,N_22073);
xor U23441 (N_23441,N_21033,N_22330);
nand U23442 (N_23442,N_21129,N_22109);
nor U23443 (N_23443,N_20664,N_20265);
nand U23444 (N_23444,N_22209,N_22418);
or U23445 (N_23445,N_20137,N_20203);
or U23446 (N_23446,N_20566,N_21184);
nor U23447 (N_23447,N_20317,N_22218);
nand U23448 (N_23448,N_21924,N_20733);
nand U23449 (N_23449,N_21231,N_20706);
or U23450 (N_23450,N_20421,N_22197);
nand U23451 (N_23451,N_22112,N_21771);
nand U23452 (N_23452,N_20459,N_21864);
nor U23453 (N_23453,N_20949,N_20994);
nor U23454 (N_23454,N_21287,N_20854);
nor U23455 (N_23455,N_20691,N_21480);
and U23456 (N_23456,N_21016,N_20936);
nor U23457 (N_23457,N_21518,N_22212);
and U23458 (N_23458,N_22054,N_21384);
nand U23459 (N_23459,N_21519,N_22172);
nor U23460 (N_23460,N_21431,N_20383);
and U23461 (N_23461,N_21836,N_20982);
and U23462 (N_23462,N_20717,N_22465);
and U23463 (N_23463,N_20977,N_21123);
xor U23464 (N_23464,N_22235,N_22342);
or U23465 (N_23465,N_20074,N_22282);
nand U23466 (N_23466,N_22123,N_22361);
or U23467 (N_23467,N_20315,N_20938);
and U23468 (N_23468,N_21945,N_20027);
xor U23469 (N_23469,N_22407,N_20788);
nand U23470 (N_23470,N_20609,N_21473);
and U23471 (N_23471,N_20935,N_20980);
xnor U23472 (N_23472,N_20306,N_21788);
and U23473 (N_23473,N_21706,N_20874);
nor U23474 (N_23474,N_21593,N_20422);
nand U23475 (N_23475,N_21648,N_20718);
xor U23476 (N_23476,N_21701,N_22059);
nor U23477 (N_23477,N_21107,N_20483);
nor U23478 (N_23478,N_22079,N_21674);
nand U23479 (N_23479,N_21330,N_21799);
or U23480 (N_23480,N_20402,N_21724);
nand U23481 (N_23481,N_20917,N_22173);
nor U23482 (N_23482,N_21664,N_21649);
and U23483 (N_23483,N_21060,N_20735);
or U23484 (N_23484,N_22171,N_21879);
xor U23485 (N_23485,N_21120,N_21437);
and U23486 (N_23486,N_20586,N_20475);
or U23487 (N_23487,N_21267,N_21640);
or U23488 (N_23488,N_20209,N_21229);
nand U23489 (N_23489,N_20287,N_21428);
nand U23490 (N_23490,N_21893,N_21283);
or U23491 (N_23491,N_21856,N_20298);
or U23492 (N_23492,N_21487,N_22026);
nand U23493 (N_23493,N_20599,N_21250);
nand U23494 (N_23494,N_20498,N_20032);
nor U23495 (N_23495,N_22304,N_21882);
and U23496 (N_23496,N_21930,N_22384);
nand U23497 (N_23497,N_20173,N_21733);
nor U23498 (N_23498,N_21497,N_20205);
or U23499 (N_23499,N_20840,N_21279);
nand U23500 (N_23500,N_21801,N_20423);
or U23501 (N_23501,N_20220,N_22497);
nand U23502 (N_23502,N_22394,N_21720);
nand U23503 (N_23503,N_21736,N_21595);
or U23504 (N_23504,N_21261,N_22075);
nor U23505 (N_23505,N_20255,N_20578);
nor U23506 (N_23506,N_22043,N_21510);
and U23507 (N_23507,N_20662,N_21700);
nand U23508 (N_23508,N_21300,N_20655);
or U23509 (N_23509,N_21302,N_21842);
nor U23510 (N_23510,N_20931,N_20154);
nor U23511 (N_23511,N_22338,N_21582);
or U23512 (N_23512,N_22495,N_21672);
or U23513 (N_23513,N_20755,N_20517);
nor U23514 (N_23514,N_21731,N_20692);
nand U23515 (N_23515,N_20289,N_20103);
nor U23516 (N_23516,N_22223,N_20606);
or U23517 (N_23517,N_20172,N_20450);
nor U23518 (N_23518,N_21274,N_21162);
nor U23519 (N_23519,N_20736,N_22000);
nor U23520 (N_23520,N_21874,N_21036);
and U23521 (N_23521,N_22449,N_20116);
nand U23522 (N_23522,N_21627,N_22096);
and U23523 (N_23523,N_20236,N_21381);
nor U23524 (N_23524,N_20564,N_21889);
nor U23525 (N_23525,N_22132,N_20753);
nor U23526 (N_23526,N_22101,N_22022);
nor U23527 (N_23527,N_20014,N_22217);
nand U23528 (N_23528,N_21492,N_20297);
nand U23529 (N_23529,N_20756,N_20525);
nor U23530 (N_23530,N_22307,N_20690);
nand U23531 (N_23531,N_20608,N_20470);
nor U23532 (N_23532,N_21248,N_21311);
nand U23533 (N_23533,N_20235,N_22277);
and U23534 (N_23534,N_22403,N_20816);
or U23535 (N_23535,N_20462,N_20081);
and U23536 (N_23536,N_21403,N_21830);
nand U23537 (N_23537,N_20355,N_20072);
nand U23538 (N_23538,N_20419,N_20538);
or U23539 (N_23539,N_22489,N_21863);
and U23540 (N_23540,N_21688,N_21887);
nor U23541 (N_23541,N_20686,N_20261);
or U23542 (N_23542,N_20604,N_20202);
nor U23543 (N_23543,N_22113,N_21933);
and U23544 (N_23544,N_21021,N_21605);
nor U23545 (N_23545,N_21695,N_21457);
or U23546 (N_23546,N_21740,N_20328);
or U23547 (N_23547,N_21327,N_22060);
nor U23548 (N_23548,N_20837,N_21976);
nor U23549 (N_23549,N_20882,N_22461);
nand U23550 (N_23550,N_21483,N_22007);
nand U23551 (N_23551,N_20110,N_21280);
and U23552 (N_23552,N_21885,N_20833);
nor U23553 (N_23553,N_20825,N_21551);
and U23554 (N_23554,N_21747,N_20215);
and U23555 (N_23555,N_21613,N_22061);
or U23556 (N_23556,N_20229,N_21739);
nor U23557 (N_23557,N_20034,N_20871);
and U23558 (N_23558,N_20957,N_21952);
nand U23559 (N_23559,N_20797,N_21380);
nor U23560 (N_23560,N_21559,N_20214);
nand U23561 (N_23561,N_21269,N_22441);
nor U23562 (N_23562,N_21459,N_20630);
and U23563 (N_23563,N_22116,N_21505);
and U23564 (N_23564,N_20169,N_21558);
nand U23565 (N_23565,N_21650,N_21687);
and U23566 (N_23566,N_22239,N_21008);
nor U23567 (N_23567,N_20076,N_20151);
or U23568 (N_23568,N_21512,N_22356);
nand U23569 (N_23569,N_21065,N_22325);
nor U23570 (N_23570,N_21704,N_22050);
nor U23571 (N_23571,N_21652,N_20671);
nor U23572 (N_23572,N_20091,N_21597);
nor U23573 (N_23573,N_20800,N_20472);
or U23574 (N_23574,N_20902,N_22027);
or U23575 (N_23575,N_20193,N_22279);
nor U23576 (N_23576,N_21562,N_22244);
nand U23577 (N_23577,N_21319,N_20335);
nor U23578 (N_23578,N_20344,N_22045);
or U23579 (N_23579,N_20164,N_22256);
nor U23580 (N_23580,N_20635,N_20228);
and U23581 (N_23581,N_20002,N_20195);
nor U23582 (N_23582,N_22321,N_21941);
nand U23583 (N_23583,N_21690,N_20393);
nand U23584 (N_23584,N_21148,N_22367);
nor U23585 (N_23585,N_21871,N_21254);
nand U23586 (N_23586,N_22070,N_22044);
and U23587 (N_23587,N_20864,N_21015);
and U23588 (N_23588,N_21824,N_20028);
nor U23589 (N_23589,N_20437,N_21448);
nor U23590 (N_23590,N_20433,N_22288);
nand U23591 (N_23591,N_20632,N_20113);
and U23592 (N_23592,N_20425,N_21903);
nor U23593 (N_23593,N_21192,N_22210);
or U23594 (N_23594,N_20379,N_20486);
nand U23595 (N_23595,N_20847,N_22192);
nor U23596 (N_23596,N_21119,N_21359);
nor U23597 (N_23597,N_21591,N_20937);
and U23598 (N_23598,N_21584,N_21977);
nor U23599 (N_23599,N_21947,N_21485);
nand U23600 (N_23600,N_22037,N_20370);
nand U23601 (N_23601,N_21973,N_20524);
nor U23602 (N_23602,N_21188,N_22175);
nor U23603 (N_23603,N_20744,N_20886);
and U23604 (N_23604,N_20367,N_20923);
and U23605 (N_23605,N_20001,N_22372);
nor U23606 (N_23606,N_21441,N_22220);
or U23607 (N_23607,N_21399,N_21472);
xnor U23608 (N_23608,N_21178,N_21949);
nand U23609 (N_23609,N_21564,N_20080);
or U23610 (N_23610,N_20244,N_20009);
nor U23611 (N_23611,N_20907,N_21606);
nand U23612 (N_23612,N_21725,N_21780);
nor U23613 (N_23613,N_21547,N_21934);
nor U23614 (N_23614,N_20819,N_20248);
nand U23615 (N_23615,N_20219,N_21539);
nand U23616 (N_23616,N_21880,N_20751);
or U23617 (N_23617,N_20892,N_20467);
and U23618 (N_23618,N_21031,N_20405);
and U23619 (N_23619,N_22299,N_20017);
nor U23620 (N_23620,N_20584,N_20293);
nand U23621 (N_23621,N_20481,N_20843);
or U23622 (N_23622,N_21646,N_21115);
nor U23623 (N_23623,N_22198,N_20305);
and U23624 (N_23624,N_22447,N_21090);
nand U23625 (N_23625,N_22124,N_22207);
nand U23626 (N_23626,N_20047,N_20277);
nor U23627 (N_23627,N_20020,N_20188);
or U23628 (N_23628,N_22036,N_22131);
and U23629 (N_23629,N_21315,N_21356);
and U23630 (N_23630,N_22067,N_21430);
nor U23631 (N_23631,N_21820,N_22408);
and U23632 (N_23632,N_21939,N_20430);
nand U23633 (N_23633,N_20750,N_20230);
nor U23634 (N_23634,N_22405,N_21447);
nor U23635 (N_23635,N_20688,N_21260);
or U23636 (N_23636,N_22063,N_20464);
nand U23637 (N_23637,N_21089,N_22068);
and U23638 (N_23638,N_20059,N_22020);
nand U23639 (N_23639,N_21335,N_20266);
or U23640 (N_23640,N_20925,N_20341);
or U23641 (N_23641,N_21098,N_21040);
and U23642 (N_23642,N_22242,N_21111);
or U23643 (N_23643,N_21782,N_21225);
or U23644 (N_23644,N_20676,N_22347);
nand U23645 (N_23645,N_22180,N_20960);
and U23646 (N_23646,N_20168,N_21020);
nor U23647 (N_23647,N_20509,N_21811);
and U23648 (N_23648,N_21633,N_21096);
and U23649 (N_23649,N_22107,N_22421);
or U23650 (N_23650,N_21419,N_20124);
nor U23651 (N_23651,N_22145,N_20148);
nor U23652 (N_23652,N_21984,N_21453);
or U23653 (N_23653,N_21922,N_20548);
or U23654 (N_23654,N_20622,N_21467);
and U23655 (N_23655,N_20232,N_20117);
or U23656 (N_23656,N_21634,N_20069);
nor U23657 (N_23657,N_21322,N_20008);
or U23658 (N_23658,N_20643,N_20711);
and U23659 (N_23659,N_21012,N_21530);
nor U23660 (N_23660,N_22219,N_20746);
and U23661 (N_23661,N_21443,N_21729);
or U23662 (N_23662,N_21624,N_20272);
and U23663 (N_23663,N_20160,N_20174);
nor U23664 (N_23664,N_20250,N_22341);
nor U23665 (N_23665,N_22358,N_21643);
nand U23666 (N_23666,N_20301,N_21835);
and U23667 (N_23667,N_21134,N_22056);
or U23668 (N_23668,N_20447,N_21576);
xor U23669 (N_23669,N_21906,N_22313);
and U23670 (N_23670,N_22234,N_21995);
xor U23671 (N_23671,N_21454,N_20352);
nor U23672 (N_23672,N_20288,N_21588);
nor U23673 (N_23673,N_20120,N_22226);
nand U23674 (N_23674,N_21171,N_20337);
or U23675 (N_23675,N_22072,N_21777);
and U23676 (N_23676,N_21209,N_22485);
or U23677 (N_23677,N_22003,N_20237);
nand U23678 (N_23678,N_20595,N_21927);
or U23679 (N_23679,N_21121,N_21507);
or U23680 (N_23680,N_21596,N_21826);
nand U23681 (N_23681,N_22278,N_20730);
and U23682 (N_23682,N_21195,N_20654);
and U23683 (N_23683,N_22143,N_21397);
and U23684 (N_23684,N_21102,N_22269);
nand U23685 (N_23685,N_22189,N_20698);
and U23686 (N_23686,N_20231,N_20007);
nor U23687 (N_23687,N_20278,N_20296);
nor U23688 (N_23688,N_21730,N_20695);
nor U23689 (N_23689,N_20964,N_21966);
or U23690 (N_23690,N_21112,N_21256);
and U23691 (N_23691,N_20263,N_20349);
or U23692 (N_23692,N_21925,N_21481);
and U23693 (N_23693,N_20651,N_20182);
nor U23694 (N_23694,N_20348,N_21619);
or U23695 (N_23695,N_20485,N_22193);
nor U23696 (N_23696,N_20510,N_21476);
nor U23697 (N_23697,N_20123,N_22419);
nor U23698 (N_23698,N_20130,N_20021);
or U23699 (N_23699,N_21511,N_21642);
nor U23700 (N_23700,N_22310,N_20404);
nand U23701 (N_23701,N_22163,N_20668);
or U23702 (N_23702,N_21222,N_20456);
or U23703 (N_23703,N_22392,N_20556);
or U23704 (N_23704,N_21309,N_20956);
or U23705 (N_23705,N_21471,N_20815);
nand U23706 (N_23706,N_21362,N_20144);
nand U23707 (N_23707,N_20145,N_20258);
and U23708 (N_23708,N_21698,N_20264);
nand U23709 (N_23709,N_21440,N_21328);
nor U23710 (N_23710,N_21458,N_21117);
and U23711 (N_23711,N_20307,N_20048);
nor U23712 (N_23712,N_21318,N_20674);
nand U23713 (N_23713,N_21392,N_21404);
nand U23714 (N_23714,N_21429,N_20099);
xnor U23715 (N_23715,N_21304,N_20842);
nand U23716 (N_23716,N_20412,N_21848);
and U23717 (N_23717,N_22470,N_22240);
nor U23718 (N_23718,N_21366,N_20282);
or U23719 (N_23719,N_21326,N_21783);
or U23720 (N_23720,N_20922,N_20830);
nor U23721 (N_23721,N_22200,N_20003);
nor U23722 (N_23722,N_21139,N_21900);
and U23723 (N_23723,N_22332,N_21807);
nor U23724 (N_23724,N_22480,N_21155);
nor U23725 (N_23725,N_21370,N_20198);
or U23726 (N_23726,N_22291,N_20042);
or U23727 (N_23727,N_20514,N_21355);
nand U23728 (N_23728,N_22431,N_21921);
nor U23729 (N_23729,N_21960,N_22294);
nor U23730 (N_23730,N_21768,N_21092);
nand U23731 (N_23731,N_22216,N_20395);
nand U23732 (N_23732,N_21773,N_21202);
or U23733 (N_23733,N_21834,N_21645);
nor U23734 (N_23734,N_22186,N_21189);
nand U23735 (N_23735,N_20995,N_21375);
and U23736 (N_23736,N_20930,N_20783);
or U23737 (N_23737,N_20157,N_22202);
or U23738 (N_23738,N_21406,N_21608);
and U23739 (N_23739,N_20619,N_20098);
nor U23740 (N_23740,N_22336,N_20410);
or U23741 (N_23741,N_20128,N_22251);
or U23742 (N_23742,N_21988,N_22382);
or U23743 (N_23743,N_21407,N_20443);
nand U23744 (N_23744,N_22281,N_22377);
nand U23745 (N_23745,N_20487,N_22297);
and U23746 (N_23746,N_22430,N_22329);
or U23747 (N_23747,N_22472,N_20392);
nand U23748 (N_23748,N_20987,N_20928);
nor U23749 (N_23749,N_21535,N_20749);
nand U23750 (N_23750,N_20985,N_22423);
and U23751 (N_23751,N_22159,N_21212);
or U23752 (N_23752,N_22324,N_21046);
or U23753 (N_23753,N_21354,N_20251);
or U23754 (N_23754,N_21679,N_20141);
nand U23755 (N_23755,N_20168,N_21824);
or U23756 (N_23756,N_21194,N_22446);
or U23757 (N_23757,N_20355,N_22219);
nand U23758 (N_23758,N_21246,N_22068);
or U23759 (N_23759,N_22376,N_22142);
nor U23760 (N_23760,N_21516,N_21011);
nor U23761 (N_23761,N_22264,N_21385);
and U23762 (N_23762,N_21039,N_20382);
nor U23763 (N_23763,N_21360,N_21221);
and U23764 (N_23764,N_21103,N_20200);
nand U23765 (N_23765,N_20181,N_21687);
nor U23766 (N_23766,N_20737,N_21548);
and U23767 (N_23767,N_21868,N_21677);
nor U23768 (N_23768,N_20591,N_21741);
and U23769 (N_23769,N_20711,N_21703);
or U23770 (N_23770,N_21501,N_21353);
and U23771 (N_23771,N_20345,N_21246);
xnor U23772 (N_23772,N_22109,N_20585);
nand U23773 (N_23773,N_20941,N_21178);
and U23774 (N_23774,N_21098,N_20627);
xor U23775 (N_23775,N_22087,N_21083);
and U23776 (N_23776,N_20342,N_20510);
nand U23777 (N_23777,N_22132,N_22410);
and U23778 (N_23778,N_20208,N_22333);
and U23779 (N_23779,N_21580,N_21623);
nand U23780 (N_23780,N_22179,N_21867);
and U23781 (N_23781,N_21913,N_20475);
or U23782 (N_23782,N_20155,N_21234);
nor U23783 (N_23783,N_21960,N_20659);
nand U23784 (N_23784,N_21053,N_21633);
nor U23785 (N_23785,N_21630,N_22463);
nand U23786 (N_23786,N_22251,N_21571);
nor U23787 (N_23787,N_20445,N_22105);
and U23788 (N_23788,N_20653,N_22161);
or U23789 (N_23789,N_21032,N_20344);
nand U23790 (N_23790,N_21314,N_20200);
nand U23791 (N_23791,N_21648,N_20558);
nand U23792 (N_23792,N_21762,N_20530);
or U23793 (N_23793,N_20522,N_21781);
nor U23794 (N_23794,N_21937,N_21139);
or U23795 (N_23795,N_20215,N_21676);
and U23796 (N_23796,N_21478,N_20552);
nand U23797 (N_23797,N_21035,N_20977);
or U23798 (N_23798,N_21663,N_21919);
and U23799 (N_23799,N_20692,N_20325);
and U23800 (N_23800,N_21382,N_21300);
nand U23801 (N_23801,N_20004,N_20193);
or U23802 (N_23802,N_21437,N_20918);
nor U23803 (N_23803,N_22469,N_20464);
or U23804 (N_23804,N_20569,N_22323);
or U23805 (N_23805,N_21481,N_22327);
and U23806 (N_23806,N_22064,N_20129);
or U23807 (N_23807,N_22447,N_20178);
nor U23808 (N_23808,N_22351,N_21449);
nor U23809 (N_23809,N_21442,N_21405);
xor U23810 (N_23810,N_20051,N_22316);
nor U23811 (N_23811,N_21755,N_21562);
nand U23812 (N_23812,N_22432,N_21255);
and U23813 (N_23813,N_20731,N_20336);
and U23814 (N_23814,N_22105,N_21908);
or U23815 (N_23815,N_20365,N_21799);
or U23816 (N_23816,N_20559,N_21600);
nor U23817 (N_23817,N_21274,N_21210);
or U23818 (N_23818,N_21830,N_22026);
and U23819 (N_23819,N_21994,N_21613);
and U23820 (N_23820,N_22422,N_20956);
and U23821 (N_23821,N_20589,N_21949);
nand U23822 (N_23822,N_20837,N_22153);
or U23823 (N_23823,N_21135,N_22065);
and U23824 (N_23824,N_20711,N_20793);
nand U23825 (N_23825,N_21892,N_20543);
nor U23826 (N_23826,N_20171,N_20000);
or U23827 (N_23827,N_20143,N_21981);
nor U23828 (N_23828,N_22187,N_22099);
and U23829 (N_23829,N_21341,N_21961);
or U23830 (N_23830,N_20164,N_20944);
and U23831 (N_23831,N_21858,N_22121);
nor U23832 (N_23832,N_20356,N_21644);
nor U23833 (N_23833,N_20049,N_22304);
or U23834 (N_23834,N_20284,N_20303);
or U23835 (N_23835,N_21370,N_21121);
nand U23836 (N_23836,N_21704,N_22182);
and U23837 (N_23837,N_20102,N_20804);
nor U23838 (N_23838,N_20359,N_20450);
nand U23839 (N_23839,N_20398,N_21762);
nand U23840 (N_23840,N_20731,N_22112);
and U23841 (N_23841,N_20312,N_22103);
nor U23842 (N_23842,N_20571,N_21288);
nor U23843 (N_23843,N_20099,N_20337);
and U23844 (N_23844,N_20457,N_21340);
nand U23845 (N_23845,N_22450,N_21772);
nor U23846 (N_23846,N_20844,N_21272);
nor U23847 (N_23847,N_21460,N_21117);
and U23848 (N_23848,N_20568,N_21887);
or U23849 (N_23849,N_21331,N_22360);
or U23850 (N_23850,N_21224,N_22486);
nand U23851 (N_23851,N_20408,N_20808);
nand U23852 (N_23852,N_20175,N_20513);
nand U23853 (N_23853,N_22206,N_21394);
nor U23854 (N_23854,N_21869,N_20240);
or U23855 (N_23855,N_21629,N_20369);
nand U23856 (N_23856,N_21638,N_22460);
nor U23857 (N_23857,N_21257,N_21063);
nand U23858 (N_23858,N_20468,N_22113);
or U23859 (N_23859,N_20301,N_22347);
nor U23860 (N_23860,N_20142,N_20898);
and U23861 (N_23861,N_21714,N_21626);
nor U23862 (N_23862,N_20977,N_21197);
or U23863 (N_23863,N_20824,N_22300);
nor U23864 (N_23864,N_20255,N_21483);
or U23865 (N_23865,N_20793,N_20632);
and U23866 (N_23866,N_21623,N_20616);
or U23867 (N_23867,N_21751,N_21653);
xor U23868 (N_23868,N_21592,N_22128);
and U23869 (N_23869,N_21577,N_21579);
nor U23870 (N_23870,N_20680,N_21541);
and U23871 (N_23871,N_20972,N_20582);
nor U23872 (N_23872,N_21196,N_22033);
nor U23873 (N_23873,N_20260,N_21927);
nand U23874 (N_23874,N_22427,N_20805);
or U23875 (N_23875,N_22212,N_20602);
and U23876 (N_23876,N_21167,N_21330);
or U23877 (N_23877,N_21062,N_22128);
and U23878 (N_23878,N_20989,N_20541);
and U23879 (N_23879,N_20493,N_21229);
nand U23880 (N_23880,N_21540,N_22396);
nand U23881 (N_23881,N_20675,N_22100);
nor U23882 (N_23882,N_21365,N_20951);
nor U23883 (N_23883,N_21940,N_20535);
nand U23884 (N_23884,N_22062,N_21193);
or U23885 (N_23885,N_20605,N_21554);
and U23886 (N_23886,N_22108,N_21550);
and U23887 (N_23887,N_21318,N_21276);
and U23888 (N_23888,N_21302,N_20047);
and U23889 (N_23889,N_21924,N_20015);
and U23890 (N_23890,N_22096,N_21194);
nor U23891 (N_23891,N_20058,N_20294);
or U23892 (N_23892,N_22055,N_20148);
nand U23893 (N_23893,N_21554,N_20340);
nor U23894 (N_23894,N_21939,N_20608);
nand U23895 (N_23895,N_22123,N_20070);
nand U23896 (N_23896,N_21712,N_20243);
or U23897 (N_23897,N_20633,N_21488);
nor U23898 (N_23898,N_21386,N_20625);
nor U23899 (N_23899,N_21783,N_20968);
xor U23900 (N_23900,N_20502,N_20966);
nand U23901 (N_23901,N_20732,N_22116);
and U23902 (N_23902,N_21665,N_21764);
nand U23903 (N_23903,N_21485,N_22351);
nand U23904 (N_23904,N_20204,N_20068);
and U23905 (N_23905,N_21066,N_21258);
nor U23906 (N_23906,N_21928,N_22149);
and U23907 (N_23907,N_21586,N_20158);
or U23908 (N_23908,N_21416,N_21137);
or U23909 (N_23909,N_20531,N_21113);
nor U23910 (N_23910,N_21354,N_20883);
nand U23911 (N_23911,N_21173,N_21214);
or U23912 (N_23912,N_21745,N_21037);
nor U23913 (N_23913,N_20968,N_20974);
nand U23914 (N_23914,N_20459,N_20576);
and U23915 (N_23915,N_21248,N_22179);
nand U23916 (N_23916,N_21742,N_20996);
nor U23917 (N_23917,N_20633,N_21196);
or U23918 (N_23918,N_21415,N_20800);
nand U23919 (N_23919,N_20620,N_21429);
and U23920 (N_23920,N_22377,N_21367);
nand U23921 (N_23921,N_20686,N_21491);
nand U23922 (N_23922,N_21436,N_20468);
nand U23923 (N_23923,N_22025,N_20356);
nor U23924 (N_23924,N_20473,N_21582);
and U23925 (N_23925,N_21330,N_21955);
nor U23926 (N_23926,N_20250,N_22468);
or U23927 (N_23927,N_22142,N_20041);
and U23928 (N_23928,N_20710,N_21790);
nand U23929 (N_23929,N_20434,N_21474);
or U23930 (N_23930,N_21298,N_21314);
and U23931 (N_23931,N_21896,N_20928);
and U23932 (N_23932,N_20207,N_21303);
or U23933 (N_23933,N_20772,N_21419);
nand U23934 (N_23934,N_21405,N_20240);
and U23935 (N_23935,N_21158,N_20497);
nand U23936 (N_23936,N_20956,N_20163);
or U23937 (N_23937,N_21853,N_20141);
nor U23938 (N_23938,N_20785,N_21943);
or U23939 (N_23939,N_20466,N_21047);
nor U23940 (N_23940,N_21449,N_20686);
nand U23941 (N_23941,N_22480,N_22143);
or U23942 (N_23942,N_20723,N_22415);
nor U23943 (N_23943,N_21912,N_22116);
and U23944 (N_23944,N_21526,N_20790);
and U23945 (N_23945,N_20337,N_20267);
or U23946 (N_23946,N_21472,N_22144);
or U23947 (N_23947,N_22213,N_20070);
nand U23948 (N_23948,N_20181,N_21324);
or U23949 (N_23949,N_20628,N_21368);
or U23950 (N_23950,N_21719,N_22422);
nor U23951 (N_23951,N_21134,N_22127);
nand U23952 (N_23952,N_20513,N_22484);
nand U23953 (N_23953,N_22477,N_20212);
nand U23954 (N_23954,N_20777,N_21073);
nor U23955 (N_23955,N_20809,N_21407);
and U23956 (N_23956,N_20299,N_21696);
or U23957 (N_23957,N_21807,N_20949);
nand U23958 (N_23958,N_20029,N_22308);
nor U23959 (N_23959,N_22364,N_20440);
or U23960 (N_23960,N_22357,N_22235);
xor U23961 (N_23961,N_20647,N_20876);
or U23962 (N_23962,N_20111,N_22246);
nand U23963 (N_23963,N_21046,N_20484);
nor U23964 (N_23964,N_20235,N_21876);
nor U23965 (N_23965,N_22377,N_22428);
nor U23966 (N_23966,N_21010,N_21108);
xor U23967 (N_23967,N_21126,N_21374);
nor U23968 (N_23968,N_20165,N_20004);
nand U23969 (N_23969,N_21705,N_21611);
and U23970 (N_23970,N_20789,N_21904);
and U23971 (N_23971,N_20685,N_20350);
or U23972 (N_23972,N_22082,N_21481);
nand U23973 (N_23973,N_20473,N_20486);
or U23974 (N_23974,N_20627,N_22188);
and U23975 (N_23975,N_20384,N_20295);
nand U23976 (N_23976,N_21713,N_21766);
nand U23977 (N_23977,N_21775,N_20523);
nand U23978 (N_23978,N_22431,N_21071);
or U23979 (N_23979,N_20095,N_20719);
or U23980 (N_23980,N_21256,N_22481);
nand U23981 (N_23981,N_21628,N_21940);
nand U23982 (N_23982,N_21022,N_21711);
nand U23983 (N_23983,N_22166,N_21579);
and U23984 (N_23984,N_21094,N_21363);
and U23985 (N_23985,N_20825,N_22448);
and U23986 (N_23986,N_20555,N_20334);
nor U23987 (N_23987,N_20721,N_22225);
nand U23988 (N_23988,N_20550,N_20827);
and U23989 (N_23989,N_21666,N_20273);
nand U23990 (N_23990,N_21838,N_20967);
xnor U23991 (N_23991,N_20577,N_21326);
and U23992 (N_23992,N_20827,N_21946);
nand U23993 (N_23993,N_20556,N_22484);
and U23994 (N_23994,N_21714,N_20227);
nor U23995 (N_23995,N_22131,N_22434);
and U23996 (N_23996,N_21955,N_21281);
nor U23997 (N_23997,N_21760,N_21933);
and U23998 (N_23998,N_20530,N_21060);
and U23999 (N_23999,N_21086,N_20715);
or U24000 (N_24000,N_20718,N_21885);
nor U24001 (N_24001,N_21448,N_22218);
or U24002 (N_24002,N_21956,N_21190);
or U24003 (N_24003,N_20127,N_22394);
nor U24004 (N_24004,N_20952,N_20445);
and U24005 (N_24005,N_21262,N_21677);
nand U24006 (N_24006,N_20997,N_20230);
nor U24007 (N_24007,N_20961,N_20364);
nand U24008 (N_24008,N_20685,N_20162);
nand U24009 (N_24009,N_20001,N_20643);
nor U24010 (N_24010,N_22407,N_21902);
nor U24011 (N_24011,N_22446,N_21707);
nor U24012 (N_24012,N_21300,N_20099);
nor U24013 (N_24013,N_21206,N_20226);
nor U24014 (N_24014,N_21931,N_20772);
or U24015 (N_24015,N_21749,N_21625);
and U24016 (N_24016,N_22475,N_22058);
or U24017 (N_24017,N_21819,N_21103);
or U24018 (N_24018,N_20583,N_21020);
nor U24019 (N_24019,N_22098,N_20034);
nand U24020 (N_24020,N_22002,N_21358);
or U24021 (N_24021,N_22225,N_22168);
nor U24022 (N_24022,N_20956,N_21360);
and U24023 (N_24023,N_20836,N_21630);
and U24024 (N_24024,N_21459,N_21494);
or U24025 (N_24025,N_20541,N_22416);
and U24026 (N_24026,N_20143,N_22178);
nand U24027 (N_24027,N_21282,N_21137);
and U24028 (N_24028,N_21301,N_21890);
or U24029 (N_24029,N_20914,N_20498);
nor U24030 (N_24030,N_21879,N_20493);
and U24031 (N_24031,N_20678,N_22376);
or U24032 (N_24032,N_20705,N_21871);
xnor U24033 (N_24033,N_22134,N_20157);
nor U24034 (N_24034,N_21594,N_22355);
and U24035 (N_24035,N_20158,N_21915);
or U24036 (N_24036,N_22434,N_22296);
nor U24037 (N_24037,N_21210,N_20552);
nor U24038 (N_24038,N_20271,N_20876);
and U24039 (N_24039,N_20346,N_20829);
nor U24040 (N_24040,N_22466,N_20082);
or U24041 (N_24041,N_20635,N_20647);
xor U24042 (N_24042,N_21583,N_20766);
nand U24043 (N_24043,N_20246,N_21720);
nand U24044 (N_24044,N_22003,N_20403);
or U24045 (N_24045,N_22015,N_20518);
xnor U24046 (N_24046,N_20348,N_20259);
and U24047 (N_24047,N_20663,N_20635);
nand U24048 (N_24048,N_22346,N_20370);
or U24049 (N_24049,N_21286,N_22059);
nand U24050 (N_24050,N_20308,N_21679);
or U24051 (N_24051,N_20797,N_21868);
nand U24052 (N_24052,N_20358,N_21479);
nand U24053 (N_24053,N_20453,N_22081);
and U24054 (N_24054,N_20050,N_20260);
nand U24055 (N_24055,N_22430,N_22473);
and U24056 (N_24056,N_21416,N_20708);
and U24057 (N_24057,N_20236,N_20263);
or U24058 (N_24058,N_21180,N_20303);
nor U24059 (N_24059,N_22449,N_22455);
nand U24060 (N_24060,N_22485,N_21968);
and U24061 (N_24061,N_21356,N_20980);
or U24062 (N_24062,N_20331,N_20349);
nand U24063 (N_24063,N_20246,N_22048);
nor U24064 (N_24064,N_20064,N_20017);
nand U24065 (N_24065,N_20760,N_20015);
nand U24066 (N_24066,N_20221,N_21671);
and U24067 (N_24067,N_21586,N_21300);
nand U24068 (N_24068,N_21904,N_21710);
xor U24069 (N_24069,N_21514,N_20430);
nand U24070 (N_24070,N_20548,N_22262);
and U24071 (N_24071,N_22088,N_21098);
nand U24072 (N_24072,N_20304,N_20929);
nand U24073 (N_24073,N_22399,N_22046);
nand U24074 (N_24074,N_21442,N_20669);
nor U24075 (N_24075,N_20454,N_21278);
or U24076 (N_24076,N_22170,N_20268);
or U24077 (N_24077,N_21339,N_20725);
nor U24078 (N_24078,N_21497,N_21870);
nor U24079 (N_24079,N_22385,N_20729);
or U24080 (N_24080,N_20506,N_20706);
or U24081 (N_24081,N_21415,N_22127);
and U24082 (N_24082,N_20158,N_20908);
nand U24083 (N_24083,N_21432,N_21714);
and U24084 (N_24084,N_21998,N_21662);
nand U24085 (N_24085,N_20164,N_21354);
nand U24086 (N_24086,N_22437,N_20379);
nor U24087 (N_24087,N_21933,N_20966);
xor U24088 (N_24088,N_20348,N_21887);
or U24089 (N_24089,N_20888,N_21462);
or U24090 (N_24090,N_21084,N_20631);
or U24091 (N_24091,N_21359,N_20755);
nor U24092 (N_24092,N_22415,N_22239);
and U24093 (N_24093,N_21095,N_20471);
nor U24094 (N_24094,N_20312,N_22165);
nor U24095 (N_24095,N_20195,N_20740);
nand U24096 (N_24096,N_21276,N_21643);
or U24097 (N_24097,N_21660,N_22466);
nand U24098 (N_24098,N_21372,N_20245);
or U24099 (N_24099,N_20480,N_21974);
nor U24100 (N_24100,N_21620,N_20030);
nand U24101 (N_24101,N_21659,N_22491);
and U24102 (N_24102,N_21608,N_20259);
or U24103 (N_24103,N_21699,N_20597);
and U24104 (N_24104,N_21971,N_20374);
nand U24105 (N_24105,N_21363,N_20565);
nor U24106 (N_24106,N_20743,N_21831);
nand U24107 (N_24107,N_21116,N_21657);
nand U24108 (N_24108,N_21989,N_20605);
nor U24109 (N_24109,N_22235,N_20271);
nor U24110 (N_24110,N_20209,N_20126);
nor U24111 (N_24111,N_22440,N_21999);
nor U24112 (N_24112,N_20238,N_22104);
or U24113 (N_24113,N_21742,N_21457);
nand U24114 (N_24114,N_21864,N_21295);
and U24115 (N_24115,N_20289,N_21032);
or U24116 (N_24116,N_21459,N_22332);
nor U24117 (N_24117,N_21400,N_20835);
or U24118 (N_24118,N_21334,N_21267);
and U24119 (N_24119,N_21302,N_21319);
nor U24120 (N_24120,N_20993,N_21433);
nand U24121 (N_24121,N_20506,N_21975);
nor U24122 (N_24122,N_20955,N_20537);
nand U24123 (N_24123,N_20062,N_21413);
and U24124 (N_24124,N_20933,N_21285);
nand U24125 (N_24125,N_20723,N_22119);
and U24126 (N_24126,N_22326,N_21049);
and U24127 (N_24127,N_20606,N_22037);
and U24128 (N_24128,N_21629,N_20906);
nor U24129 (N_24129,N_22307,N_21318);
nand U24130 (N_24130,N_20906,N_22136);
nand U24131 (N_24131,N_20647,N_22281);
and U24132 (N_24132,N_21997,N_20908);
or U24133 (N_24133,N_21905,N_20786);
and U24134 (N_24134,N_21000,N_22456);
nor U24135 (N_24135,N_20735,N_20427);
and U24136 (N_24136,N_21893,N_20494);
nand U24137 (N_24137,N_22483,N_22058);
xor U24138 (N_24138,N_20023,N_22435);
and U24139 (N_24139,N_22262,N_22114);
nand U24140 (N_24140,N_20285,N_20742);
and U24141 (N_24141,N_21114,N_21762);
or U24142 (N_24142,N_21093,N_21987);
nand U24143 (N_24143,N_21593,N_20529);
nand U24144 (N_24144,N_22325,N_21691);
nand U24145 (N_24145,N_21184,N_21245);
nor U24146 (N_24146,N_21226,N_20565);
and U24147 (N_24147,N_21191,N_21041);
nand U24148 (N_24148,N_20341,N_21256);
nor U24149 (N_24149,N_21689,N_20964);
or U24150 (N_24150,N_20183,N_20827);
and U24151 (N_24151,N_21152,N_21140);
or U24152 (N_24152,N_21068,N_22099);
and U24153 (N_24153,N_22416,N_20663);
or U24154 (N_24154,N_22294,N_20022);
or U24155 (N_24155,N_22050,N_20549);
or U24156 (N_24156,N_21025,N_20385);
and U24157 (N_24157,N_21669,N_20614);
nand U24158 (N_24158,N_22024,N_21001);
and U24159 (N_24159,N_21428,N_21805);
or U24160 (N_24160,N_22105,N_22323);
and U24161 (N_24161,N_20591,N_21565);
or U24162 (N_24162,N_20750,N_21821);
nor U24163 (N_24163,N_22071,N_21784);
and U24164 (N_24164,N_22100,N_21643);
nor U24165 (N_24165,N_21680,N_21083);
and U24166 (N_24166,N_21023,N_20196);
xnor U24167 (N_24167,N_22435,N_22195);
and U24168 (N_24168,N_21507,N_20074);
xnor U24169 (N_24169,N_21158,N_21000);
or U24170 (N_24170,N_21004,N_20786);
nand U24171 (N_24171,N_20119,N_22263);
and U24172 (N_24172,N_22203,N_20755);
nand U24173 (N_24173,N_21605,N_20214);
and U24174 (N_24174,N_20402,N_20412);
nand U24175 (N_24175,N_20796,N_22226);
and U24176 (N_24176,N_20279,N_22077);
and U24177 (N_24177,N_20668,N_21343);
nor U24178 (N_24178,N_22477,N_20518);
nand U24179 (N_24179,N_21169,N_22205);
nand U24180 (N_24180,N_21742,N_22415);
or U24181 (N_24181,N_20481,N_20518);
nor U24182 (N_24182,N_21393,N_22328);
nand U24183 (N_24183,N_21600,N_20479);
or U24184 (N_24184,N_21192,N_20803);
or U24185 (N_24185,N_20262,N_20575);
and U24186 (N_24186,N_22188,N_20037);
nor U24187 (N_24187,N_21316,N_20175);
nor U24188 (N_24188,N_22314,N_22021);
nand U24189 (N_24189,N_20809,N_21473);
or U24190 (N_24190,N_20844,N_21766);
and U24191 (N_24191,N_21774,N_22292);
nand U24192 (N_24192,N_21713,N_21205);
nor U24193 (N_24193,N_21884,N_22082);
nand U24194 (N_24194,N_21205,N_20666);
nor U24195 (N_24195,N_20108,N_21382);
nand U24196 (N_24196,N_20736,N_21215);
or U24197 (N_24197,N_21140,N_20871);
or U24198 (N_24198,N_20286,N_21834);
and U24199 (N_24199,N_20081,N_22455);
nand U24200 (N_24200,N_20357,N_20083);
nand U24201 (N_24201,N_20722,N_20533);
nand U24202 (N_24202,N_21762,N_22091);
and U24203 (N_24203,N_21450,N_21779);
nand U24204 (N_24204,N_22404,N_21456);
or U24205 (N_24205,N_21857,N_20168);
nand U24206 (N_24206,N_21040,N_20745);
and U24207 (N_24207,N_20818,N_20858);
nor U24208 (N_24208,N_20424,N_20203);
nand U24209 (N_24209,N_20056,N_20499);
nor U24210 (N_24210,N_21570,N_22256);
nor U24211 (N_24211,N_20365,N_22309);
and U24212 (N_24212,N_22366,N_20622);
and U24213 (N_24213,N_21785,N_20447);
and U24214 (N_24214,N_21305,N_20105);
nor U24215 (N_24215,N_22451,N_21417);
nor U24216 (N_24216,N_22218,N_20407);
nor U24217 (N_24217,N_22229,N_21948);
nor U24218 (N_24218,N_20616,N_20697);
or U24219 (N_24219,N_21894,N_20939);
and U24220 (N_24220,N_22059,N_20830);
or U24221 (N_24221,N_22407,N_20757);
and U24222 (N_24222,N_20983,N_20298);
nor U24223 (N_24223,N_22444,N_20880);
or U24224 (N_24224,N_20281,N_20645);
nor U24225 (N_24225,N_22056,N_20207);
nor U24226 (N_24226,N_20057,N_21358);
and U24227 (N_24227,N_21409,N_20038);
and U24228 (N_24228,N_20757,N_20100);
nor U24229 (N_24229,N_20883,N_21458);
nor U24230 (N_24230,N_21867,N_20034);
nand U24231 (N_24231,N_21972,N_20267);
nand U24232 (N_24232,N_21573,N_21959);
or U24233 (N_24233,N_22354,N_20102);
or U24234 (N_24234,N_20658,N_22242);
nor U24235 (N_24235,N_22161,N_20420);
nand U24236 (N_24236,N_21491,N_21215);
and U24237 (N_24237,N_20486,N_21725);
nor U24238 (N_24238,N_20400,N_21341);
nand U24239 (N_24239,N_20839,N_21960);
or U24240 (N_24240,N_20656,N_21963);
and U24241 (N_24241,N_20324,N_21643);
nor U24242 (N_24242,N_20893,N_21668);
nor U24243 (N_24243,N_21625,N_20427);
nand U24244 (N_24244,N_20230,N_21416);
nor U24245 (N_24245,N_20483,N_20688);
nor U24246 (N_24246,N_20408,N_21723);
and U24247 (N_24247,N_21558,N_21159);
nand U24248 (N_24248,N_21219,N_22340);
xnor U24249 (N_24249,N_21766,N_22429);
or U24250 (N_24250,N_21994,N_22132);
and U24251 (N_24251,N_20136,N_20830);
and U24252 (N_24252,N_20513,N_21916);
nor U24253 (N_24253,N_22301,N_21405);
nor U24254 (N_24254,N_20264,N_20751);
nor U24255 (N_24255,N_20630,N_20405);
or U24256 (N_24256,N_21228,N_21242);
nand U24257 (N_24257,N_20689,N_21518);
nand U24258 (N_24258,N_20671,N_20005);
or U24259 (N_24259,N_21046,N_21224);
nor U24260 (N_24260,N_21387,N_21322);
or U24261 (N_24261,N_20792,N_20555);
and U24262 (N_24262,N_20955,N_21731);
nor U24263 (N_24263,N_21289,N_21012);
nor U24264 (N_24264,N_21110,N_20251);
and U24265 (N_24265,N_20253,N_21503);
or U24266 (N_24266,N_20992,N_20815);
nor U24267 (N_24267,N_20713,N_20847);
nor U24268 (N_24268,N_20384,N_20194);
and U24269 (N_24269,N_21070,N_20288);
or U24270 (N_24270,N_21525,N_21734);
and U24271 (N_24271,N_20541,N_21198);
nand U24272 (N_24272,N_21410,N_20776);
xor U24273 (N_24273,N_20292,N_20837);
and U24274 (N_24274,N_20360,N_20444);
or U24275 (N_24275,N_21613,N_20913);
or U24276 (N_24276,N_21190,N_20692);
and U24277 (N_24277,N_21687,N_21087);
and U24278 (N_24278,N_20213,N_21480);
and U24279 (N_24279,N_21879,N_20521);
or U24280 (N_24280,N_21610,N_21132);
and U24281 (N_24281,N_21816,N_20017);
nor U24282 (N_24282,N_21006,N_22379);
nand U24283 (N_24283,N_22078,N_20512);
nor U24284 (N_24284,N_20635,N_20341);
nor U24285 (N_24285,N_21864,N_20656);
or U24286 (N_24286,N_21482,N_20585);
and U24287 (N_24287,N_22276,N_21500);
nand U24288 (N_24288,N_21780,N_21593);
nor U24289 (N_24289,N_21855,N_22069);
nand U24290 (N_24290,N_22353,N_22457);
and U24291 (N_24291,N_21472,N_21237);
and U24292 (N_24292,N_21351,N_20537);
nand U24293 (N_24293,N_22151,N_20490);
nor U24294 (N_24294,N_20433,N_20584);
and U24295 (N_24295,N_20080,N_21625);
and U24296 (N_24296,N_20405,N_20286);
nand U24297 (N_24297,N_21818,N_20940);
nand U24298 (N_24298,N_20671,N_20292);
and U24299 (N_24299,N_22005,N_20879);
or U24300 (N_24300,N_21861,N_21815);
nand U24301 (N_24301,N_21295,N_21468);
nand U24302 (N_24302,N_20814,N_20440);
or U24303 (N_24303,N_21906,N_20662);
nor U24304 (N_24304,N_20808,N_21224);
nand U24305 (N_24305,N_20222,N_21771);
nor U24306 (N_24306,N_20674,N_21521);
nand U24307 (N_24307,N_20342,N_22193);
or U24308 (N_24308,N_20829,N_20194);
nor U24309 (N_24309,N_21449,N_20298);
nor U24310 (N_24310,N_21422,N_21152);
nor U24311 (N_24311,N_22293,N_20544);
or U24312 (N_24312,N_21213,N_21022);
nand U24313 (N_24313,N_20240,N_22458);
or U24314 (N_24314,N_20316,N_22353);
nand U24315 (N_24315,N_22295,N_22430);
nand U24316 (N_24316,N_21633,N_21258);
and U24317 (N_24317,N_20609,N_21337);
or U24318 (N_24318,N_21510,N_21682);
nor U24319 (N_24319,N_22055,N_22082);
or U24320 (N_24320,N_20111,N_20569);
and U24321 (N_24321,N_21730,N_20967);
nor U24322 (N_24322,N_20751,N_20954);
nor U24323 (N_24323,N_21767,N_21722);
nand U24324 (N_24324,N_20638,N_22353);
nor U24325 (N_24325,N_22166,N_21423);
nor U24326 (N_24326,N_20019,N_22156);
and U24327 (N_24327,N_20158,N_20567);
nand U24328 (N_24328,N_20076,N_22385);
or U24329 (N_24329,N_21201,N_20337);
nand U24330 (N_24330,N_21801,N_20033);
nor U24331 (N_24331,N_20495,N_20327);
nand U24332 (N_24332,N_21713,N_22330);
nand U24333 (N_24333,N_21019,N_21898);
or U24334 (N_24334,N_22253,N_20190);
or U24335 (N_24335,N_21373,N_22444);
xnor U24336 (N_24336,N_20988,N_20303);
nor U24337 (N_24337,N_21617,N_20882);
nand U24338 (N_24338,N_21570,N_20863);
or U24339 (N_24339,N_20959,N_20919);
and U24340 (N_24340,N_21219,N_20032);
nand U24341 (N_24341,N_20464,N_20513);
and U24342 (N_24342,N_20643,N_22026);
nand U24343 (N_24343,N_20654,N_22106);
and U24344 (N_24344,N_20818,N_21123);
nor U24345 (N_24345,N_20231,N_21466);
or U24346 (N_24346,N_20976,N_20305);
nor U24347 (N_24347,N_22151,N_20432);
nor U24348 (N_24348,N_20795,N_20154);
xor U24349 (N_24349,N_21749,N_21724);
or U24350 (N_24350,N_20699,N_21985);
nand U24351 (N_24351,N_21813,N_21604);
nand U24352 (N_24352,N_20271,N_21861);
or U24353 (N_24353,N_22303,N_20695);
and U24354 (N_24354,N_20835,N_21331);
nand U24355 (N_24355,N_20488,N_20208);
and U24356 (N_24356,N_20476,N_20638);
or U24357 (N_24357,N_21188,N_22064);
nand U24358 (N_24358,N_21179,N_20664);
and U24359 (N_24359,N_20207,N_20763);
nand U24360 (N_24360,N_21208,N_22375);
nor U24361 (N_24361,N_20542,N_21071);
nor U24362 (N_24362,N_20750,N_21385);
or U24363 (N_24363,N_21460,N_21378);
or U24364 (N_24364,N_21786,N_20903);
nand U24365 (N_24365,N_21985,N_21301);
nor U24366 (N_24366,N_21686,N_21565);
or U24367 (N_24367,N_20292,N_21001);
and U24368 (N_24368,N_20066,N_20134);
or U24369 (N_24369,N_22479,N_21052);
nand U24370 (N_24370,N_21914,N_22106);
and U24371 (N_24371,N_22428,N_20510);
and U24372 (N_24372,N_22047,N_20360);
and U24373 (N_24373,N_21355,N_21557);
nor U24374 (N_24374,N_21635,N_21606);
nor U24375 (N_24375,N_20085,N_20484);
or U24376 (N_24376,N_20228,N_20277);
nand U24377 (N_24377,N_22275,N_22041);
or U24378 (N_24378,N_21784,N_20183);
xnor U24379 (N_24379,N_21344,N_21984);
and U24380 (N_24380,N_21686,N_20864);
nand U24381 (N_24381,N_21444,N_20907);
and U24382 (N_24382,N_20198,N_20407);
nor U24383 (N_24383,N_20330,N_21414);
or U24384 (N_24384,N_20100,N_20906);
nor U24385 (N_24385,N_21186,N_22064);
nor U24386 (N_24386,N_21327,N_21544);
nor U24387 (N_24387,N_21683,N_22219);
or U24388 (N_24388,N_21126,N_20275);
nor U24389 (N_24389,N_21783,N_20989);
or U24390 (N_24390,N_21651,N_20936);
and U24391 (N_24391,N_20549,N_22317);
or U24392 (N_24392,N_22196,N_21116);
nand U24393 (N_24393,N_22060,N_20974);
or U24394 (N_24394,N_20698,N_22052);
or U24395 (N_24395,N_21574,N_22230);
nand U24396 (N_24396,N_20029,N_21486);
nor U24397 (N_24397,N_20424,N_21194);
and U24398 (N_24398,N_21610,N_22282);
nor U24399 (N_24399,N_22395,N_21590);
nor U24400 (N_24400,N_22363,N_22145);
or U24401 (N_24401,N_20268,N_21734);
or U24402 (N_24402,N_21359,N_21759);
or U24403 (N_24403,N_22258,N_22143);
nand U24404 (N_24404,N_21154,N_20618);
or U24405 (N_24405,N_21454,N_21583);
nand U24406 (N_24406,N_21039,N_21497);
nor U24407 (N_24407,N_22158,N_22423);
or U24408 (N_24408,N_21665,N_20077);
xnor U24409 (N_24409,N_22460,N_21356);
nor U24410 (N_24410,N_20252,N_22493);
nor U24411 (N_24411,N_20853,N_21631);
xor U24412 (N_24412,N_21335,N_20610);
nor U24413 (N_24413,N_22461,N_22310);
nand U24414 (N_24414,N_20923,N_21515);
nand U24415 (N_24415,N_20910,N_21892);
and U24416 (N_24416,N_22421,N_21941);
nand U24417 (N_24417,N_20896,N_20181);
nand U24418 (N_24418,N_20315,N_20144);
and U24419 (N_24419,N_22470,N_20534);
or U24420 (N_24420,N_20056,N_22353);
nand U24421 (N_24421,N_20069,N_21811);
or U24422 (N_24422,N_21056,N_20742);
nand U24423 (N_24423,N_21324,N_20331);
or U24424 (N_24424,N_21089,N_20782);
and U24425 (N_24425,N_22037,N_21644);
and U24426 (N_24426,N_21798,N_22018);
or U24427 (N_24427,N_21055,N_22146);
nor U24428 (N_24428,N_20595,N_22136);
or U24429 (N_24429,N_21706,N_22323);
nor U24430 (N_24430,N_20361,N_21587);
nand U24431 (N_24431,N_20407,N_20277);
nor U24432 (N_24432,N_20442,N_20440);
or U24433 (N_24433,N_21099,N_22247);
or U24434 (N_24434,N_21578,N_22291);
xor U24435 (N_24435,N_21157,N_20171);
and U24436 (N_24436,N_20560,N_21150);
or U24437 (N_24437,N_21936,N_21201);
xor U24438 (N_24438,N_21444,N_21197);
and U24439 (N_24439,N_22405,N_21321);
nand U24440 (N_24440,N_20652,N_22062);
or U24441 (N_24441,N_21742,N_20127);
and U24442 (N_24442,N_22119,N_21523);
nand U24443 (N_24443,N_22229,N_22391);
nor U24444 (N_24444,N_20535,N_20690);
nand U24445 (N_24445,N_21096,N_22196);
nand U24446 (N_24446,N_20501,N_21829);
nand U24447 (N_24447,N_20877,N_22005);
nand U24448 (N_24448,N_21093,N_21271);
nor U24449 (N_24449,N_20864,N_20528);
nor U24450 (N_24450,N_21145,N_20989);
or U24451 (N_24451,N_21739,N_20128);
nor U24452 (N_24452,N_20600,N_20199);
nand U24453 (N_24453,N_21906,N_21813);
and U24454 (N_24454,N_22385,N_20934);
or U24455 (N_24455,N_22128,N_21418);
nor U24456 (N_24456,N_20924,N_21916);
nand U24457 (N_24457,N_21745,N_20307);
or U24458 (N_24458,N_20194,N_20587);
or U24459 (N_24459,N_20177,N_22417);
nor U24460 (N_24460,N_22329,N_20380);
or U24461 (N_24461,N_21452,N_21386);
nand U24462 (N_24462,N_21125,N_21151);
and U24463 (N_24463,N_22442,N_21414);
or U24464 (N_24464,N_21189,N_21152);
nand U24465 (N_24465,N_21154,N_20430);
xnor U24466 (N_24466,N_21715,N_21466);
nor U24467 (N_24467,N_20167,N_22219);
or U24468 (N_24468,N_20823,N_20382);
nand U24469 (N_24469,N_20665,N_21727);
or U24470 (N_24470,N_22491,N_20218);
nor U24471 (N_24471,N_21780,N_21230);
nand U24472 (N_24472,N_21999,N_20610);
and U24473 (N_24473,N_20839,N_21716);
and U24474 (N_24474,N_21135,N_20732);
nor U24475 (N_24475,N_22387,N_22004);
nor U24476 (N_24476,N_20174,N_21920);
and U24477 (N_24477,N_21080,N_20593);
nor U24478 (N_24478,N_22431,N_20076);
nor U24479 (N_24479,N_21647,N_22162);
nand U24480 (N_24480,N_21433,N_20097);
nor U24481 (N_24481,N_20144,N_20542);
nor U24482 (N_24482,N_21921,N_21299);
nor U24483 (N_24483,N_20290,N_21889);
or U24484 (N_24484,N_20783,N_20494);
and U24485 (N_24485,N_21510,N_20854);
or U24486 (N_24486,N_20730,N_20521);
or U24487 (N_24487,N_21207,N_22451);
nor U24488 (N_24488,N_22273,N_20968);
nor U24489 (N_24489,N_22392,N_21655);
nor U24490 (N_24490,N_22334,N_21270);
or U24491 (N_24491,N_20867,N_21245);
nor U24492 (N_24492,N_21181,N_20415);
or U24493 (N_24493,N_21832,N_22033);
and U24494 (N_24494,N_21267,N_21014);
or U24495 (N_24495,N_21094,N_22208);
nand U24496 (N_24496,N_20206,N_22239);
nand U24497 (N_24497,N_20671,N_21348);
nor U24498 (N_24498,N_20371,N_21683);
nor U24499 (N_24499,N_21097,N_22125);
nor U24500 (N_24500,N_22322,N_20187);
xor U24501 (N_24501,N_21013,N_21783);
or U24502 (N_24502,N_21129,N_21648);
or U24503 (N_24503,N_21303,N_22320);
and U24504 (N_24504,N_21407,N_21296);
xor U24505 (N_24505,N_20362,N_21493);
or U24506 (N_24506,N_21261,N_20444);
and U24507 (N_24507,N_20526,N_21930);
and U24508 (N_24508,N_20434,N_21730);
or U24509 (N_24509,N_20619,N_21233);
nor U24510 (N_24510,N_21314,N_21190);
or U24511 (N_24511,N_21867,N_22077);
or U24512 (N_24512,N_20337,N_20560);
and U24513 (N_24513,N_22210,N_21823);
nand U24514 (N_24514,N_20931,N_20842);
or U24515 (N_24515,N_20439,N_22058);
nor U24516 (N_24516,N_20481,N_21956);
or U24517 (N_24517,N_20079,N_20798);
nand U24518 (N_24518,N_20420,N_22090);
nor U24519 (N_24519,N_20993,N_21909);
nor U24520 (N_24520,N_21614,N_20598);
nand U24521 (N_24521,N_21868,N_22404);
or U24522 (N_24522,N_21881,N_21925);
or U24523 (N_24523,N_22171,N_22492);
nand U24524 (N_24524,N_21911,N_20602);
and U24525 (N_24525,N_20328,N_21275);
and U24526 (N_24526,N_22232,N_21957);
nand U24527 (N_24527,N_21487,N_21107);
and U24528 (N_24528,N_22281,N_21824);
nor U24529 (N_24529,N_21440,N_21053);
or U24530 (N_24530,N_21991,N_20453);
or U24531 (N_24531,N_20988,N_22269);
and U24532 (N_24532,N_21846,N_21769);
or U24533 (N_24533,N_21550,N_21729);
or U24534 (N_24534,N_22248,N_21248);
and U24535 (N_24535,N_22288,N_20723);
and U24536 (N_24536,N_20913,N_20140);
nand U24537 (N_24537,N_21354,N_21548);
or U24538 (N_24538,N_21525,N_21284);
nor U24539 (N_24539,N_21660,N_20270);
or U24540 (N_24540,N_22334,N_20023);
and U24541 (N_24541,N_22274,N_20220);
or U24542 (N_24542,N_20460,N_20170);
or U24543 (N_24543,N_21942,N_21643);
or U24544 (N_24544,N_20952,N_21628);
nand U24545 (N_24545,N_21083,N_21097);
and U24546 (N_24546,N_21518,N_20282);
nand U24547 (N_24547,N_20567,N_22395);
nand U24548 (N_24548,N_21776,N_21721);
or U24549 (N_24549,N_21119,N_21787);
nor U24550 (N_24550,N_21584,N_21258);
or U24551 (N_24551,N_22119,N_21826);
xnor U24552 (N_24552,N_21365,N_20174);
or U24553 (N_24553,N_21774,N_20135);
and U24554 (N_24554,N_21266,N_21510);
nand U24555 (N_24555,N_20679,N_21646);
nand U24556 (N_24556,N_21343,N_20308);
nand U24557 (N_24557,N_22344,N_21557);
nor U24558 (N_24558,N_22287,N_22038);
or U24559 (N_24559,N_22178,N_20758);
and U24560 (N_24560,N_20650,N_20762);
or U24561 (N_24561,N_22390,N_20458);
nand U24562 (N_24562,N_21102,N_21161);
or U24563 (N_24563,N_20838,N_21786);
nor U24564 (N_24564,N_21844,N_20146);
nor U24565 (N_24565,N_20547,N_20149);
nor U24566 (N_24566,N_20960,N_21286);
and U24567 (N_24567,N_22351,N_22157);
or U24568 (N_24568,N_22070,N_20760);
and U24569 (N_24569,N_21328,N_21386);
or U24570 (N_24570,N_20637,N_21962);
and U24571 (N_24571,N_21974,N_22352);
or U24572 (N_24572,N_21067,N_21120);
nand U24573 (N_24573,N_21544,N_20280);
or U24574 (N_24574,N_20106,N_21534);
and U24575 (N_24575,N_21308,N_20401);
nor U24576 (N_24576,N_20036,N_22188);
or U24577 (N_24577,N_21091,N_21537);
or U24578 (N_24578,N_21534,N_21438);
and U24579 (N_24579,N_20377,N_20873);
or U24580 (N_24580,N_21444,N_21011);
nor U24581 (N_24581,N_21022,N_21616);
nor U24582 (N_24582,N_20277,N_20737);
nand U24583 (N_24583,N_20252,N_22062);
or U24584 (N_24584,N_21711,N_22243);
or U24585 (N_24585,N_20629,N_20732);
or U24586 (N_24586,N_21854,N_22497);
nor U24587 (N_24587,N_21246,N_21801);
or U24588 (N_24588,N_21606,N_22473);
nor U24589 (N_24589,N_22332,N_21561);
nor U24590 (N_24590,N_22373,N_21288);
or U24591 (N_24591,N_21743,N_21187);
and U24592 (N_24592,N_22485,N_20903);
nor U24593 (N_24593,N_21804,N_21590);
and U24594 (N_24594,N_20239,N_20414);
nor U24595 (N_24595,N_20147,N_21108);
nand U24596 (N_24596,N_20748,N_21533);
nand U24597 (N_24597,N_22328,N_20846);
nor U24598 (N_24598,N_21178,N_21247);
nor U24599 (N_24599,N_20449,N_20404);
nor U24600 (N_24600,N_20590,N_21545);
and U24601 (N_24601,N_20682,N_20960);
or U24602 (N_24602,N_20193,N_21229);
and U24603 (N_24603,N_22349,N_20489);
and U24604 (N_24604,N_20698,N_21838);
and U24605 (N_24605,N_21100,N_21309);
or U24606 (N_24606,N_20823,N_20663);
xor U24607 (N_24607,N_21525,N_21714);
nand U24608 (N_24608,N_20123,N_20772);
nand U24609 (N_24609,N_20783,N_20841);
nand U24610 (N_24610,N_22385,N_22137);
nor U24611 (N_24611,N_20254,N_20429);
nor U24612 (N_24612,N_20773,N_21647);
or U24613 (N_24613,N_22381,N_20314);
nor U24614 (N_24614,N_21193,N_20678);
nor U24615 (N_24615,N_21224,N_21352);
or U24616 (N_24616,N_20630,N_22042);
and U24617 (N_24617,N_22061,N_21798);
and U24618 (N_24618,N_20492,N_22422);
nor U24619 (N_24619,N_22397,N_22163);
nand U24620 (N_24620,N_20455,N_20296);
nor U24621 (N_24621,N_21284,N_20465);
nor U24622 (N_24622,N_20412,N_22363);
nor U24623 (N_24623,N_20506,N_20361);
and U24624 (N_24624,N_22153,N_21543);
nor U24625 (N_24625,N_21916,N_21945);
nand U24626 (N_24626,N_21147,N_21535);
nand U24627 (N_24627,N_20314,N_20426);
and U24628 (N_24628,N_20774,N_20418);
nand U24629 (N_24629,N_21731,N_22155);
or U24630 (N_24630,N_21335,N_21269);
nand U24631 (N_24631,N_20784,N_20377);
and U24632 (N_24632,N_21209,N_20754);
nor U24633 (N_24633,N_21408,N_20757);
xor U24634 (N_24634,N_21232,N_22300);
or U24635 (N_24635,N_20492,N_21308);
and U24636 (N_24636,N_21425,N_20565);
nor U24637 (N_24637,N_20479,N_20815);
and U24638 (N_24638,N_20144,N_20183);
nor U24639 (N_24639,N_20710,N_21879);
nor U24640 (N_24640,N_21872,N_20028);
nand U24641 (N_24641,N_20446,N_21303);
and U24642 (N_24642,N_21686,N_21782);
xor U24643 (N_24643,N_21256,N_22157);
and U24644 (N_24644,N_20967,N_20086);
or U24645 (N_24645,N_21590,N_20965);
nand U24646 (N_24646,N_21463,N_22364);
nor U24647 (N_24647,N_21418,N_21651);
nor U24648 (N_24648,N_21728,N_20016);
nand U24649 (N_24649,N_20988,N_21596);
nand U24650 (N_24650,N_20557,N_21439);
or U24651 (N_24651,N_20476,N_21098);
and U24652 (N_24652,N_20373,N_20567);
nor U24653 (N_24653,N_22439,N_20099);
nand U24654 (N_24654,N_20992,N_22306);
xor U24655 (N_24655,N_21223,N_21281);
nor U24656 (N_24656,N_21549,N_22412);
nand U24657 (N_24657,N_21837,N_21577);
or U24658 (N_24658,N_20735,N_21454);
or U24659 (N_24659,N_20641,N_22279);
nor U24660 (N_24660,N_21454,N_20806);
and U24661 (N_24661,N_22417,N_22250);
or U24662 (N_24662,N_20397,N_22471);
nand U24663 (N_24663,N_22287,N_21684);
and U24664 (N_24664,N_22479,N_20389);
nor U24665 (N_24665,N_20152,N_21131);
or U24666 (N_24666,N_22261,N_20952);
nor U24667 (N_24667,N_20873,N_21188);
or U24668 (N_24668,N_20197,N_21870);
nor U24669 (N_24669,N_20263,N_20489);
nand U24670 (N_24670,N_21970,N_20580);
and U24671 (N_24671,N_20619,N_20099);
or U24672 (N_24672,N_20033,N_22211);
nor U24673 (N_24673,N_20804,N_20957);
and U24674 (N_24674,N_20015,N_22193);
nor U24675 (N_24675,N_20786,N_20389);
nand U24676 (N_24676,N_20014,N_20708);
nor U24677 (N_24677,N_20674,N_21807);
and U24678 (N_24678,N_20185,N_21151);
nor U24679 (N_24679,N_21099,N_20033);
nor U24680 (N_24680,N_21074,N_20084);
and U24681 (N_24681,N_21962,N_20126);
or U24682 (N_24682,N_20304,N_20531);
or U24683 (N_24683,N_21872,N_20136);
nor U24684 (N_24684,N_21071,N_21615);
nand U24685 (N_24685,N_20466,N_20334);
or U24686 (N_24686,N_20811,N_20189);
nand U24687 (N_24687,N_21072,N_20836);
and U24688 (N_24688,N_22254,N_20431);
and U24689 (N_24689,N_21849,N_20554);
or U24690 (N_24690,N_22200,N_21722);
and U24691 (N_24691,N_20208,N_21075);
nand U24692 (N_24692,N_21037,N_21146);
or U24693 (N_24693,N_20842,N_20152);
and U24694 (N_24694,N_21538,N_21359);
nor U24695 (N_24695,N_21935,N_21289);
or U24696 (N_24696,N_22417,N_20479);
or U24697 (N_24697,N_21188,N_21156);
nor U24698 (N_24698,N_20868,N_22379);
and U24699 (N_24699,N_22293,N_20011);
or U24700 (N_24700,N_20559,N_21112);
nand U24701 (N_24701,N_20794,N_21549);
or U24702 (N_24702,N_21916,N_21587);
and U24703 (N_24703,N_20789,N_21445);
or U24704 (N_24704,N_20653,N_20713);
nor U24705 (N_24705,N_21070,N_22162);
xnor U24706 (N_24706,N_21336,N_22365);
or U24707 (N_24707,N_21525,N_20437);
nand U24708 (N_24708,N_21519,N_20371);
nor U24709 (N_24709,N_21085,N_20498);
and U24710 (N_24710,N_21642,N_22372);
and U24711 (N_24711,N_21811,N_21491);
nor U24712 (N_24712,N_22080,N_21579);
nand U24713 (N_24713,N_21475,N_22343);
nor U24714 (N_24714,N_22340,N_20724);
nor U24715 (N_24715,N_21523,N_21683);
or U24716 (N_24716,N_20527,N_21503);
and U24717 (N_24717,N_22367,N_21264);
or U24718 (N_24718,N_20060,N_21120);
nand U24719 (N_24719,N_20825,N_21325);
or U24720 (N_24720,N_21377,N_22209);
nor U24721 (N_24721,N_21241,N_20821);
xnor U24722 (N_24722,N_20867,N_21930);
nand U24723 (N_24723,N_20464,N_22102);
or U24724 (N_24724,N_21813,N_21043);
nor U24725 (N_24725,N_20287,N_21383);
and U24726 (N_24726,N_21352,N_20360);
or U24727 (N_24727,N_20625,N_21075);
nor U24728 (N_24728,N_21067,N_20054);
nand U24729 (N_24729,N_20627,N_20994);
nand U24730 (N_24730,N_21644,N_21112);
nand U24731 (N_24731,N_21534,N_20973);
nor U24732 (N_24732,N_20506,N_21310);
and U24733 (N_24733,N_20523,N_21945);
nor U24734 (N_24734,N_22457,N_21212);
or U24735 (N_24735,N_21653,N_20427);
and U24736 (N_24736,N_20528,N_21870);
nor U24737 (N_24737,N_20249,N_22354);
nor U24738 (N_24738,N_20545,N_22267);
nor U24739 (N_24739,N_21038,N_22450);
nand U24740 (N_24740,N_22020,N_21715);
nand U24741 (N_24741,N_21466,N_20344);
xor U24742 (N_24742,N_22159,N_21070);
or U24743 (N_24743,N_22160,N_20534);
nor U24744 (N_24744,N_21188,N_21393);
nand U24745 (N_24745,N_20604,N_20807);
xor U24746 (N_24746,N_21658,N_20727);
and U24747 (N_24747,N_21909,N_21199);
or U24748 (N_24748,N_22162,N_20429);
and U24749 (N_24749,N_21388,N_20164);
nor U24750 (N_24750,N_22051,N_20529);
and U24751 (N_24751,N_20599,N_22137);
or U24752 (N_24752,N_20180,N_21404);
and U24753 (N_24753,N_21917,N_21292);
nor U24754 (N_24754,N_21782,N_22170);
and U24755 (N_24755,N_21291,N_21247);
or U24756 (N_24756,N_20692,N_21531);
nand U24757 (N_24757,N_20247,N_22042);
or U24758 (N_24758,N_22174,N_21699);
nor U24759 (N_24759,N_21764,N_20405);
or U24760 (N_24760,N_21378,N_21486);
or U24761 (N_24761,N_21460,N_21736);
nor U24762 (N_24762,N_20773,N_21552);
nor U24763 (N_24763,N_20024,N_21153);
or U24764 (N_24764,N_21694,N_20687);
nor U24765 (N_24765,N_21628,N_22385);
and U24766 (N_24766,N_22484,N_22353);
nand U24767 (N_24767,N_21635,N_20142);
and U24768 (N_24768,N_20415,N_21115);
and U24769 (N_24769,N_20290,N_22084);
nand U24770 (N_24770,N_21887,N_21450);
or U24771 (N_24771,N_22017,N_22492);
or U24772 (N_24772,N_21990,N_21687);
and U24773 (N_24773,N_21026,N_21016);
and U24774 (N_24774,N_20378,N_20260);
and U24775 (N_24775,N_21468,N_20704);
nand U24776 (N_24776,N_21356,N_21879);
or U24777 (N_24777,N_20330,N_20918);
or U24778 (N_24778,N_20790,N_22417);
or U24779 (N_24779,N_20610,N_22239);
and U24780 (N_24780,N_21084,N_21717);
nand U24781 (N_24781,N_22245,N_22463);
nand U24782 (N_24782,N_20826,N_20725);
and U24783 (N_24783,N_20673,N_21069);
nand U24784 (N_24784,N_20566,N_20729);
or U24785 (N_24785,N_21593,N_21994);
or U24786 (N_24786,N_20509,N_20214);
or U24787 (N_24787,N_20575,N_21713);
or U24788 (N_24788,N_22252,N_20179);
nor U24789 (N_24789,N_21687,N_21750);
and U24790 (N_24790,N_21914,N_20176);
and U24791 (N_24791,N_20880,N_22355);
xnor U24792 (N_24792,N_20060,N_21260);
and U24793 (N_24793,N_20684,N_20501);
and U24794 (N_24794,N_20327,N_21572);
nand U24795 (N_24795,N_21441,N_21149);
nand U24796 (N_24796,N_21381,N_20120);
and U24797 (N_24797,N_22039,N_21164);
nor U24798 (N_24798,N_21185,N_21036);
and U24799 (N_24799,N_22431,N_20827);
nor U24800 (N_24800,N_21175,N_21304);
nand U24801 (N_24801,N_22339,N_21768);
and U24802 (N_24802,N_21112,N_22166);
or U24803 (N_24803,N_20316,N_20105);
and U24804 (N_24804,N_22288,N_21688);
nand U24805 (N_24805,N_20899,N_21180);
nor U24806 (N_24806,N_21029,N_20797);
nor U24807 (N_24807,N_21991,N_22133);
nand U24808 (N_24808,N_22176,N_21673);
nor U24809 (N_24809,N_22357,N_21160);
or U24810 (N_24810,N_21932,N_21848);
nand U24811 (N_24811,N_20372,N_21618);
nor U24812 (N_24812,N_21446,N_21023);
nor U24813 (N_24813,N_20471,N_20697);
and U24814 (N_24814,N_20375,N_21786);
nand U24815 (N_24815,N_21534,N_21329);
nor U24816 (N_24816,N_20405,N_20869);
or U24817 (N_24817,N_21676,N_21373);
and U24818 (N_24818,N_20635,N_22491);
nor U24819 (N_24819,N_20716,N_20678);
and U24820 (N_24820,N_20558,N_20862);
and U24821 (N_24821,N_22230,N_22498);
or U24822 (N_24822,N_21030,N_20601);
nand U24823 (N_24823,N_21874,N_20298);
nor U24824 (N_24824,N_22437,N_20288);
nand U24825 (N_24825,N_21944,N_22464);
nor U24826 (N_24826,N_20471,N_21348);
and U24827 (N_24827,N_20977,N_22464);
nor U24828 (N_24828,N_20843,N_22028);
and U24829 (N_24829,N_20891,N_20903);
and U24830 (N_24830,N_21379,N_21017);
nand U24831 (N_24831,N_20114,N_20106);
or U24832 (N_24832,N_21984,N_20786);
and U24833 (N_24833,N_22278,N_21360);
nand U24834 (N_24834,N_21457,N_20654);
nand U24835 (N_24835,N_21073,N_21233);
nand U24836 (N_24836,N_22059,N_20918);
nand U24837 (N_24837,N_21644,N_21238);
or U24838 (N_24838,N_20154,N_20850);
and U24839 (N_24839,N_21833,N_20795);
and U24840 (N_24840,N_20372,N_21125);
nor U24841 (N_24841,N_20207,N_21826);
nor U24842 (N_24842,N_20258,N_20896);
nor U24843 (N_24843,N_20517,N_21181);
and U24844 (N_24844,N_20012,N_20793);
nor U24845 (N_24845,N_21588,N_21087);
nand U24846 (N_24846,N_20742,N_21386);
nand U24847 (N_24847,N_20184,N_22370);
nand U24848 (N_24848,N_20791,N_21313);
nor U24849 (N_24849,N_20477,N_21159);
nand U24850 (N_24850,N_21020,N_20587);
and U24851 (N_24851,N_20626,N_21797);
nand U24852 (N_24852,N_20338,N_21181);
nand U24853 (N_24853,N_21681,N_22079);
xnor U24854 (N_24854,N_21613,N_21568);
nand U24855 (N_24855,N_20674,N_22210);
and U24856 (N_24856,N_21990,N_22436);
and U24857 (N_24857,N_22337,N_21868);
nand U24858 (N_24858,N_21620,N_20322);
nand U24859 (N_24859,N_21811,N_21779);
nand U24860 (N_24860,N_20426,N_20895);
nand U24861 (N_24861,N_20600,N_21574);
nor U24862 (N_24862,N_20615,N_22485);
and U24863 (N_24863,N_21935,N_21946);
nand U24864 (N_24864,N_22485,N_20431);
or U24865 (N_24865,N_20843,N_22433);
nor U24866 (N_24866,N_21551,N_20288);
nor U24867 (N_24867,N_22376,N_22364);
nor U24868 (N_24868,N_20623,N_22353);
nor U24869 (N_24869,N_21600,N_21916);
nor U24870 (N_24870,N_20465,N_22456);
nand U24871 (N_24871,N_20828,N_20479);
nor U24872 (N_24872,N_20943,N_21202);
nor U24873 (N_24873,N_21729,N_20853);
nor U24874 (N_24874,N_22273,N_21308);
nand U24875 (N_24875,N_21235,N_22453);
or U24876 (N_24876,N_20495,N_20811);
nor U24877 (N_24877,N_21009,N_21100);
and U24878 (N_24878,N_21562,N_21071);
and U24879 (N_24879,N_21391,N_20526);
nand U24880 (N_24880,N_20165,N_22344);
nor U24881 (N_24881,N_20190,N_21359);
and U24882 (N_24882,N_22472,N_20656);
or U24883 (N_24883,N_20220,N_21723);
or U24884 (N_24884,N_22373,N_20555);
nand U24885 (N_24885,N_21500,N_21530);
nor U24886 (N_24886,N_22020,N_20321);
nand U24887 (N_24887,N_20920,N_21376);
nand U24888 (N_24888,N_22336,N_21819);
and U24889 (N_24889,N_21790,N_21480);
nor U24890 (N_24890,N_20905,N_20312);
or U24891 (N_24891,N_20116,N_20459);
and U24892 (N_24892,N_20543,N_21438);
and U24893 (N_24893,N_20906,N_20936);
or U24894 (N_24894,N_21659,N_20709);
or U24895 (N_24895,N_22187,N_21431);
nor U24896 (N_24896,N_21509,N_21965);
or U24897 (N_24897,N_22318,N_21089);
or U24898 (N_24898,N_20678,N_21551);
nor U24899 (N_24899,N_22208,N_21383);
and U24900 (N_24900,N_21841,N_20065);
and U24901 (N_24901,N_21862,N_22101);
or U24902 (N_24902,N_21708,N_22373);
or U24903 (N_24903,N_20195,N_21682);
nor U24904 (N_24904,N_20073,N_21681);
nor U24905 (N_24905,N_21777,N_21568);
nand U24906 (N_24906,N_20847,N_21168);
or U24907 (N_24907,N_22266,N_20194);
and U24908 (N_24908,N_20699,N_20888);
nor U24909 (N_24909,N_20112,N_20072);
and U24910 (N_24910,N_21880,N_21215);
nor U24911 (N_24911,N_20369,N_20007);
nand U24912 (N_24912,N_20556,N_20208);
and U24913 (N_24913,N_22021,N_21710);
xnor U24914 (N_24914,N_21762,N_21494);
and U24915 (N_24915,N_20926,N_20918);
nor U24916 (N_24916,N_21505,N_20715);
or U24917 (N_24917,N_22241,N_20160);
nor U24918 (N_24918,N_21261,N_21630);
nor U24919 (N_24919,N_20126,N_21414);
nand U24920 (N_24920,N_20182,N_22324);
nand U24921 (N_24921,N_20630,N_21521);
or U24922 (N_24922,N_22387,N_21687);
and U24923 (N_24923,N_20437,N_22345);
and U24924 (N_24924,N_22197,N_22022);
and U24925 (N_24925,N_20449,N_21434);
or U24926 (N_24926,N_20562,N_21263);
nand U24927 (N_24927,N_21145,N_22226);
and U24928 (N_24928,N_20957,N_21022);
nor U24929 (N_24929,N_20342,N_21035);
and U24930 (N_24930,N_21344,N_21193);
or U24931 (N_24931,N_22064,N_21168);
xor U24932 (N_24932,N_20849,N_21577);
nand U24933 (N_24933,N_22384,N_21817);
nor U24934 (N_24934,N_21841,N_22019);
nand U24935 (N_24935,N_20647,N_20111);
nor U24936 (N_24936,N_22202,N_20503);
or U24937 (N_24937,N_21827,N_21595);
and U24938 (N_24938,N_20742,N_21023);
or U24939 (N_24939,N_20508,N_21325);
nand U24940 (N_24940,N_20812,N_20461);
or U24941 (N_24941,N_20739,N_20730);
nor U24942 (N_24942,N_20185,N_21712);
nor U24943 (N_24943,N_22349,N_20482);
nand U24944 (N_24944,N_21487,N_20666);
or U24945 (N_24945,N_21038,N_21689);
or U24946 (N_24946,N_22115,N_20378);
nor U24947 (N_24947,N_20033,N_20841);
nor U24948 (N_24948,N_21331,N_21118);
or U24949 (N_24949,N_20704,N_20889);
nand U24950 (N_24950,N_21820,N_20155);
nor U24951 (N_24951,N_20999,N_22417);
and U24952 (N_24952,N_21034,N_20439);
nor U24953 (N_24953,N_22253,N_21297);
nor U24954 (N_24954,N_21585,N_20053);
xor U24955 (N_24955,N_20288,N_21881);
or U24956 (N_24956,N_21755,N_21773);
nand U24957 (N_24957,N_22168,N_21737);
nor U24958 (N_24958,N_20725,N_20434);
nor U24959 (N_24959,N_22185,N_21729);
and U24960 (N_24960,N_20999,N_22434);
and U24961 (N_24961,N_21644,N_20761);
or U24962 (N_24962,N_20388,N_20020);
nand U24963 (N_24963,N_22249,N_21648);
and U24964 (N_24964,N_22142,N_21280);
and U24965 (N_24965,N_20140,N_21626);
nand U24966 (N_24966,N_22415,N_21617);
and U24967 (N_24967,N_21827,N_21082);
nand U24968 (N_24968,N_20044,N_21266);
or U24969 (N_24969,N_20903,N_22036);
and U24970 (N_24970,N_20162,N_22376);
nor U24971 (N_24971,N_20671,N_21856);
nand U24972 (N_24972,N_20732,N_21212);
and U24973 (N_24973,N_22469,N_21004);
nor U24974 (N_24974,N_21319,N_21132);
or U24975 (N_24975,N_20852,N_21649);
and U24976 (N_24976,N_21443,N_20589);
and U24977 (N_24977,N_20613,N_21888);
and U24978 (N_24978,N_22004,N_22256);
nand U24979 (N_24979,N_21197,N_20983);
or U24980 (N_24980,N_20203,N_21354);
and U24981 (N_24981,N_20709,N_21656);
nand U24982 (N_24982,N_20383,N_20769);
and U24983 (N_24983,N_20038,N_22436);
nor U24984 (N_24984,N_20470,N_22284);
nor U24985 (N_24985,N_21190,N_21491);
nor U24986 (N_24986,N_22295,N_22406);
and U24987 (N_24987,N_21681,N_21450);
and U24988 (N_24988,N_21313,N_22386);
and U24989 (N_24989,N_20488,N_22336);
nor U24990 (N_24990,N_20332,N_21039);
and U24991 (N_24991,N_21391,N_20946);
nand U24992 (N_24992,N_21450,N_22099);
nor U24993 (N_24993,N_20356,N_21319);
or U24994 (N_24994,N_20487,N_21553);
or U24995 (N_24995,N_20271,N_21796);
and U24996 (N_24996,N_21708,N_20577);
and U24997 (N_24997,N_22368,N_22186);
nor U24998 (N_24998,N_22328,N_21534);
nand U24999 (N_24999,N_21503,N_22367);
nor UO_0 (O_0,N_24444,N_23401);
or UO_1 (O_1,N_24325,N_23833);
and UO_2 (O_2,N_24974,N_23439);
or UO_3 (O_3,N_24052,N_23483);
or UO_4 (O_4,N_24122,N_23074);
xnor UO_5 (O_5,N_23493,N_24097);
nand UO_6 (O_6,N_24482,N_23886);
or UO_7 (O_7,N_23955,N_22611);
or UO_8 (O_8,N_22773,N_22823);
nor UO_9 (O_9,N_23871,N_24723);
or UO_10 (O_10,N_24508,N_22624);
or UO_11 (O_11,N_23432,N_22574);
nor UO_12 (O_12,N_24707,N_23595);
nand UO_13 (O_13,N_22691,N_23038);
xnor UO_14 (O_14,N_22808,N_23400);
nand UO_15 (O_15,N_23636,N_24000);
nand UO_16 (O_16,N_23316,N_23692);
and UO_17 (O_17,N_23120,N_24445);
nor UO_18 (O_18,N_23617,N_23371);
and UO_19 (O_19,N_24350,N_24581);
or UO_20 (O_20,N_24388,N_24254);
nand UO_21 (O_21,N_23440,N_22983);
or UO_22 (O_22,N_23296,N_23431);
and UO_23 (O_23,N_23682,N_23999);
xnor UO_24 (O_24,N_24976,N_23157);
and UO_25 (O_25,N_23399,N_23445);
and UO_26 (O_26,N_24830,N_24366);
nor UO_27 (O_27,N_22519,N_24661);
and UO_28 (O_28,N_24179,N_23675);
or UO_29 (O_29,N_24697,N_23072);
or UO_30 (O_30,N_24213,N_23453);
and UO_31 (O_31,N_24685,N_24170);
xnor UO_32 (O_32,N_22671,N_23248);
and UO_33 (O_33,N_24869,N_24935);
or UO_34 (O_34,N_23312,N_23963);
or UO_35 (O_35,N_22863,N_22657);
nor UO_36 (O_36,N_22775,N_24314);
and UO_37 (O_37,N_24136,N_24424);
nor UO_38 (O_38,N_22670,N_23530);
nor UO_39 (O_39,N_24165,N_24562);
and UO_40 (O_40,N_23986,N_24251);
nor UO_41 (O_41,N_24308,N_23897);
or UO_42 (O_42,N_24531,N_23497);
or UO_43 (O_43,N_23482,N_23424);
or UO_44 (O_44,N_22964,N_22552);
nor UO_45 (O_45,N_23556,N_24250);
nor UO_46 (O_46,N_23931,N_24733);
and UO_47 (O_47,N_23511,N_24345);
or UO_48 (O_48,N_23954,N_23385);
and UO_49 (O_49,N_24691,N_23063);
nand UO_50 (O_50,N_23328,N_24855);
xnor UO_51 (O_51,N_24135,N_23116);
or UO_52 (O_52,N_23438,N_23405);
nor UO_53 (O_53,N_23021,N_22750);
and UO_54 (O_54,N_22674,N_24474);
nor UO_55 (O_55,N_23374,N_23767);
nor UO_56 (O_56,N_23885,N_23714);
nand UO_57 (O_57,N_22778,N_23980);
and UO_58 (O_58,N_22570,N_23087);
and UO_59 (O_59,N_23646,N_24241);
or UO_60 (O_60,N_23997,N_24867);
and UO_61 (O_61,N_24601,N_22876);
and UO_62 (O_62,N_24646,N_24450);
xnor UO_63 (O_63,N_22903,N_23149);
and UO_64 (O_64,N_24972,N_23029);
or UO_65 (O_65,N_23967,N_22697);
and UO_66 (O_66,N_22625,N_24014);
and UO_67 (O_67,N_23232,N_23119);
and UO_68 (O_68,N_24954,N_24281);
and UO_69 (O_69,N_23152,N_23547);
nand UO_70 (O_70,N_22963,N_23478);
or UO_71 (O_71,N_24434,N_24049);
and UO_72 (O_72,N_22613,N_22988);
and UO_73 (O_73,N_23787,N_23929);
or UO_74 (O_74,N_24473,N_24083);
nor UO_75 (O_75,N_24307,N_22937);
nand UO_76 (O_76,N_24740,N_23076);
nor UO_77 (O_77,N_24619,N_22515);
or UO_78 (O_78,N_24909,N_23867);
and UO_79 (O_79,N_23621,N_23114);
nand UO_80 (O_80,N_22616,N_24469);
nand UO_81 (O_81,N_22965,N_23446);
or UO_82 (O_82,N_24537,N_24632);
or UO_83 (O_83,N_22796,N_23088);
or UO_84 (O_84,N_24893,N_24876);
xnor UO_85 (O_85,N_23090,N_24868);
nand UO_86 (O_86,N_23139,N_24512);
nor UO_87 (O_87,N_24595,N_24713);
or UO_88 (O_88,N_23529,N_24523);
nor UO_89 (O_89,N_22998,N_22545);
and UO_90 (O_90,N_23196,N_24328);
nor UO_91 (O_91,N_23056,N_22844);
nand UO_92 (O_92,N_24212,N_23190);
nand UO_93 (O_93,N_22803,N_24572);
or UO_94 (O_94,N_23026,N_23960);
nand UO_95 (O_95,N_22850,N_24813);
and UO_96 (O_96,N_23080,N_24229);
nand UO_97 (O_97,N_23845,N_23396);
or UO_98 (O_98,N_24702,N_23049);
nor UO_99 (O_99,N_24695,N_24468);
nand UO_100 (O_100,N_24311,N_24421);
and UO_101 (O_101,N_24189,N_23988);
nor UO_102 (O_102,N_22733,N_22580);
or UO_103 (O_103,N_22842,N_23659);
or UO_104 (O_104,N_23020,N_23605);
nor UO_105 (O_105,N_24109,N_24019);
nand UO_106 (O_106,N_24912,N_22522);
nand UO_107 (O_107,N_24988,N_23002);
and UO_108 (O_108,N_23790,N_23422);
or UO_109 (O_109,N_24783,N_24475);
and UO_110 (O_110,N_23594,N_22690);
and UO_111 (O_111,N_23541,N_23552);
nor UO_112 (O_112,N_23805,N_24573);
nor UO_113 (O_113,N_23146,N_24276);
or UO_114 (O_114,N_24406,N_23883);
or UO_115 (O_115,N_23343,N_24860);
and UO_116 (O_116,N_23227,N_23408);
and UO_117 (O_117,N_23661,N_24653);
nand UO_118 (O_118,N_23749,N_24509);
nand UO_119 (O_119,N_22914,N_23943);
nor UO_120 (O_120,N_23472,N_23142);
or UO_121 (O_121,N_24665,N_23054);
nor UO_122 (O_122,N_24181,N_23461);
or UO_123 (O_123,N_23180,N_22753);
and UO_124 (O_124,N_22781,N_23950);
nor UO_125 (O_125,N_22684,N_24105);
or UO_126 (O_126,N_24304,N_23794);
nor UO_127 (O_127,N_24794,N_24211);
nand UO_128 (O_128,N_22834,N_23429);
nand UO_129 (O_129,N_23225,N_22540);
and UO_130 (O_130,N_23939,N_23702);
or UO_131 (O_131,N_24614,N_22752);
or UO_132 (O_132,N_24177,N_24678);
nor UO_133 (O_133,N_24022,N_24957);
or UO_134 (O_134,N_22512,N_23420);
nor UO_135 (O_135,N_22831,N_24732);
or UO_136 (O_136,N_22547,N_24992);
nand UO_137 (O_137,N_24409,N_22524);
nor UO_138 (O_138,N_23349,N_22841);
or UO_139 (O_139,N_23220,N_24761);
nand UO_140 (O_140,N_24645,N_22666);
and UO_141 (O_141,N_24031,N_24643);
nand UO_142 (O_142,N_22770,N_23938);
nand UO_143 (O_143,N_24076,N_23647);
or UO_144 (O_144,N_23736,N_23508);
and UO_145 (O_145,N_22683,N_23103);
or UO_146 (O_146,N_23630,N_24127);
and UO_147 (O_147,N_22804,N_23747);
or UO_148 (O_148,N_23923,N_22664);
or UO_149 (O_149,N_23224,N_23753);
nor UO_150 (O_150,N_22979,N_23481);
nor UO_151 (O_151,N_23856,N_23912);
nor UO_152 (O_152,N_22676,N_24730);
nor UO_153 (O_153,N_22571,N_24817);
and UO_154 (O_154,N_23847,N_23154);
nor UO_155 (O_155,N_24499,N_24367);
nand UO_156 (O_156,N_24102,N_24519);
or UO_157 (O_157,N_24438,N_23032);
or UO_158 (O_158,N_22838,N_22660);
nor UO_159 (O_159,N_22723,N_24005);
nor UO_160 (O_160,N_24045,N_23584);
and UO_161 (O_161,N_22543,N_24630);
nor UO_162 (O_162,N_24377,N_24575);
nor UO_163 (O_163,N_23018,N_24979);
nand UO_164 (O_164,N_22650,N_23195);
nand UO_165 (O_165,N_23607,N_23359);
nand UO_166 (O_166,N_22853,N_24620);
and UO_167 (O_167,N_22910,N_24582);
nor UO_168 (O_168,N_23430,N_24717);
nor UO_169 (O_169,N_23106,N_23470);
nand UO_170 (O_170,N_23047,N_24080);
or UO_171 (O_171,N_24806,N_23690);
nor UO_172 (O_172,N_24309,N_22899);
or UO_173 (O_173,N_24948,N_23459);
nor UO_174 (O_174,N_24965,N_23167);
nor UO_175 (O_175,N_23616,N_22786);
and UO_176 (O_176,N_24820,N_24809);
nor UO_177 (O_177,N_24811,N_24106);
and UO_178 (O_178,N_24655,N_24905);
nor UO_179 (O_179,N_23598,N_22952);
nor UO_180 (O_180,N_24718,N_22587);
and UO_181 (O_181,N_24557,N_23522);
nor UO_182 (O_182,N_23689,N_22934);
nor UO_183 (O_183,N_24639,N_24313);
and UO_184 (O_184,N_24461,N_22620);
nor UO_185 (O_185,N_22962,N_24348);
and UO_186 (O_186,N_23231,N_23066);
and UO_187 (O_187,N_24664,N_24034);
and UO_188 (O_188,N_23992,N_23411);
nand UO_189 (O_189,N_23192,N_24126);
nor UO_190 (O_190,N_24810,N_24611);
and UO_191 (O_191,N_22901,N_22658);
nor UO_192 (O_192,N_22956,N_24880);
nand UO_193 (O_193,N_22761,N_23544);
and UO_194 (O_194,N_24082,N_24477);
nor UO_195 (O_195,N_23267,N_24541);
nand UO_196 (O_196,N_24962,N_22704);
or UO_197 (O_197,N_24403,N_24318);
nor UO_198 (O_198,N_24413,N_23243);
nor UO_199 (O_199,N_22629,N_23022);
and UO_200 (O_200,N_22523,N_24946);
and UO_201 (O_201,N_24815,N_24795);
nor UO_202 (O_202,N_24949,N_22961);
nand UO_203 (O_203,N_24143,N_22572);
nand UO_204 (O_204,N_23699,N_23314);
xnor UO_205 (O_205,N_23618,N_23928);
and UO_206 (O_206,N_24654,N_23474);
or UO_207 (O_207,N_24771,N_23981);
nor UO_208 (O_208,N_24090,N_22981);
and UO_209 (O_209,N_24627,N_22550);
nor UO_210 (O_210,N_23290,N_23532);
nand UO_211 (O_211,N_23683,N_23669);
nor UO_212 (O_212,N_23247,N_23573);
nand UO_213 (O_213,N_24779,N_24487);
nand UO_214 (O_214,N_24963,N_22929);
and UO_215 (O_215,N_23651,N_23202);
nand UO_216 (O_216,N_24226,N_24570);
or UO_217 (O_217,N_22977,N_22928);
nor UO_218 (O_218,N_24566,N_24004);
or UO_219 (O_219,N_23093,N_23578);
nand UO_220 (O_220,N_23326,N_24807);
nand UO_221 (O_221,N_23574,N_23306);
and UO_222 (O_222,N_24383,N_24968);
or UO_223 (O_223,N_24818,N_22996);
or UO_224 (O_224,N_23304,N_23271);
and UO_225 (O_225,N_22513,N_24452);
and UO_226 (O_226,N_22782,N_24621);
and UO_227 (O_227,N_23170,N_23638);
or UO_228 (O_228,N_22677,N_22717);
nor UO_229 (O_229,N_23887,N_23746);
and UO_230 (O_230,N_23131,N_24650);
or UO_231 (O_231,N_24491,N_22746);
nand UO_232 (O_232,N_24535,N_22588);
nand UO_233 (O_233,N_23412,N_24699);
and UO_234 (O_234,N_24134,N_23866);
and UO_235 (O_235,N_24618,N_24920);
nand UO_236 (O_236,N_22971,N_23339);
xor UO_237 (O_237,N_24094,N_24742);
and UO_238 (O_238,N_24245,N_23277);
nor UO_239 (O_239,N_24638,N_24900);
or UO_240 (O_240,N_24055,N_23193);
and UO_241 (O_241,N_24574,N_23857);
and UO_242 (O_242,N_23609,N_24986);
nor UO_243 (O_243,N_23217,N_23336);
and UO_244 (O_244,N_23899,N_23589);
nor UO_245 (O_245,N_23942,N_23759);
or UO_246 (O_246,N_24773,N_24069);
nand UO_247 (O_247,N_24703,N_24323);
nor UO_248 (O_248,N_23294,N_22789);
nor UO_249 (O_249,N_24628,N_23261);
and UO_250 (O_250,N_24032,N_23754);
and UO_251 (O_251,N_24040,N_22685);
nand UO_252 (O_252,N_23084,N_24224);
nand UO_253 (O_253,N_24694,N_23040);
or UO_254 (O_254,N_22626,N_22551);
nand UO_255 (O_255,N_22654,N_24238);
or UO_256 (O_256,N_24151,N_23330);
and UO_257 (O_257,N_23397,N_23308);
nand UO_258 (O_258,N_24684,N_23665);
or UO_259 (O_259,N_23023,N_24145);
and UO_260 (O_260,N_23017,N_24405);
and UO_261 (O_261,N_23571,N_23373);
nor UO_262 (O_262,N_24158,N_23388);
nor UO_263 (O_263,N_23460,N_24997);
and UO_264 (O_264,N_24327,N_23783);
and UO_265 (O_265,N_24175,N_24884);
nor UO_266 (O_266,N_22800,N_23464);
nand UO_267 (O_267,N_23859,N_24751);
or UO_268 (O_268,N_23164,N_22711);
xor UO_269 (O_269,N_24039,N_24285);
and UO_270 (O_270,N_22505,N_22749);
nand UO_271 (O_271,N_22906,N_22787);
and UO_272 (O_272,N_23724,N_22825);
nor UO_273 (O_273,N_24495,N_24511);
or UO_274 (O_274,N_24176,N_23537);
and UO_275 (O_275,N_23278,N_23414);
nor UO_276 (O_276,N_22887,N_23379);
nand UO_277 (O_277,N_24010,N_24816);
nor UO_278 (O_278,N_23097,N_24008);
and UO_279 (O_279,N_23198,N_24980);
nor UO_280 (O_280,N_23518,N_23569);
nor UO_281 (O_281,N_24470,N_24200);
nand UO_282 (O_282,N_23035,N_23624);
nor UO_283 (O_283,N_24674,N_23488);
nor UO_284 (O_284,N_23145,N_22900);
nand UO_285 (O_285,N_22663,N_24890);
nor UO_286 (O_286,N_24927,N_23540);
or UO_287 (O_287,N_23713,N_23698);
nand UO_288 (O_288,N_24871,N_23300);
or UO_289 (O_289,N_22705,N_23315);
and UO_290 (O_290,N_24658,N_24462);
nand UO_291 (O_291,N_24141,N_24784);
or UO_292 (O_292,N_22701,N_23737);
and UO_293 (O_293,N_22919,N_24183);
or UO_294 (O_294,N_23704,N_24063);
and UO_295 (O_295,N_23042,N_24746);
nand UO_296 (O_296,N_23117,N_24422);
and UO_297 (O_297,N_24825,N_24494);
and UO_298 (O_298,N_23810,N_24446);
and UO_299 (O_299,N_23194,N_22764);
nor UO_300 (O_300,N_24289,N_22954);
nand UO_301 (O_301,N_22542,N_23784);
and UO_302 (O_302,N_23990,N_24896);
nand UO_303 (O_303,N_22958,N_22508);
or UO_304 (O_304,N_24944,N_23345);
nor UO_305 (O_305,N_24607,N_22741);
nand UO_306 (O_306,N_24522,N_23269);
or UO_307 (O_307,N_24199,N_23521);
nor UO_308 (O_308,N_23548,N_23138);
nand UO_309 (O_309,N_23982,N_22659);
nor UO_310 (O_310,N_23283,N_23101);
or UO_311 (O_311,N_23118,N_24184);
nand UO_312 (O_312,N_24246,N_23706);
and UO_313 (O_313,N_24260,N_24616);
nor UO_314 (O_314,N_24924,N_23477);
nand UO_315 (O_315,N_23109,N_23756);
and UO_316 (O_316,N_24196,N_23615);
nand UO_317 (O_317,N_24271,N_23681);
nand UO_318 (O_318,N_24440,N_22826);
and UO_319 (O_319,N_22699,N_22763);
nor UO_320 (O_320,N_23352,N_24851);
nor UO_321 (O_321,N_24764,N_23380);
and UO_322 (O_322,N_22879,N_22707);
nand UO_323 (O_323,N_23168,N_24330);
or UO_324 (O_324,N_24776,N_23869);
or UO_325 (O_325,N_23978,N_23825);
and UO_326 (O_326,N_23898,N_24305);
nand UO_327 (O_327,N_23046,N_24803);
nand UO_328 (O_328,N_24514,N_23358);
or UO_329 (O_329,N_24819,N_23081);
and UO_330 (O_330,N_23865,N_23827);
nand UO_331 (O_331,N_23095,N_23586);
nor UO_332 (O_332,N_22722,N_23009);
nand UO_333 (O_333,N_23191,N_22639);
and UO_334 (O_334,N_24875,N_24945);
nor UO_335 (O_335,N_23357,N_24326);
and UO_336 (O_336,N_23826,N_24385);
nor UO_337 (O_337,N_23741,N_23171);
nor UO_338 (O_338,N_24534,N_22567);
and UO_339 (O_339,N_24775,N_24078);
and UO_340 (O_340,N_22589,N_23610);
or UO_341 (O_341,N_24041,N_23134);
or UO_342 (O_342,N_23496,N_23822);
and UO_343 (O_343,N_22991,N_23421);
or UO_344 (O_344,N_22821,N_24496);
nand UO_345 (O_345,N_24597,N_24364);
and UO_346 (O_346,N_23701,N_23775);
or UO_347 (O_347,N_23075,N_24966);
nor UO_348 (O_348,N_24858,N_22970);
nand UO_349 (O_349,N_23821,N_24024);
nand UO_350 (O_350,N_24692,N_24579);
or UO_351 (O_351,N_24964,N_22633);
or UO_352 (O_352,N_24365,N_24451);
nor UO_353 (O_353,N_24210,N_22669);
nor UO_354 (O_354,N_23757,N_22682);
and UO_355 (O_355,N_23674,N_23717);
nor UO_356 (O_356,N_22672,N_24417);
nor UO_357 (O_357,N_24216,N_23874);
xnor UO_358 (O_358,N_23454,N_23050);
and UO_359 (O_359,N_24370,N_24969);
or UO_360 (O_360,N_23498,N_23776);
nor UO_361 (O_361,N_23815,N_23016);
nor UO_362 (O_362,N_22916,N_23423);
or UO_363 (O_363,N_23937,N_24297);
or UO_364 (O_364,N_23773,N_22514);
or UO_365 (O_365,N_23655,N_23900);
xnor UO_366 (O_366,N_24524,N_23705);
and UO_367 (O_367,N_24208,N_23480);
nand UO_368 (O_368,N_23207,N_23280);
nor UO_369 (O_369,N_22893,N_23218);
nand UO_370 (O_370,N_23203,N_23910);
or UO_371 (O_371,N_24398,N_24735);
or UO_372 (O_372,N_24635,N_24433);
and UO_373 (O_373,N_24058,N_22873);
and UO_374 (O_374,N_24724,N_24263);
nand UO_375 (O_375,N_22725,N_24625);
nor UO_376 (O_376,N_24373,N_22767);
and UO_377 (O_377,N_22696,N_23200);
or UO_378 (O_378,N_23443,N_23186);
and UO_379 (O_379,N_22840,N_23415);
nand UO_380 (O_380,N_24361,N_23475);
and UO_381 (O_381,N_22501,N_23351);
and UO_382 (O_382,N_24124,N_23214);
nor UO_383 (O_383,N_23786,N_23677);
and UO_384 (O_384,N_22835,N_23144);
xor UO_385 (O_385,N_23069,N_22836);
and UO_386 (O_386,N_23000,N_23025);
nor UO_387 (O_387,N_23739,N_23209);
or UO_388 (O_388,N_24259,N_23505);
xor UO_389 (O_389,N_24696,N_24299);
nand UO_390 (O_390,N_23848,N_22640);
or UO_391 (O_391,N_24885,N_24479);
and UO_392 (O_392,N_23175,N_23156);
nand UO_393 (O_393,N_23284,N_23804);
xnor UO_394 (O_394,N_23995,N_23356);
nand UO_395 (O_395,N_23012,N_23223);
nand UO_396 (O_396,N_24353,N_23951);
or UO_397 (O_397,N_23004,N_23915);
or UO_398 (O_398,N_23637,N_23324);
and UO_399 (O_399,N_22875,N_24756);
or UO_400 (O_400,N_24682,N_22646);
nand UO_401 (O_401,N_24894,N_23500);
and UO_402 (O_402,N_22862,N_23542);
nor UO_403 (O_403,N_23515,N_24546);
nand UO_404 (O_404,N_22990,N_22905);
or UO_405 (O_405,N_24693,N_24140);
or UO_406 (O_406,N_24286,N_22813);
xor UO_407 (O_407,N_24466,N_24476);
and UO_408 (O_408,N_23876,N_23348);
or UO_409 (O_409,N_23592,N_24392);
or UO_410 (O_410,N_23872,N_24605);
nor UO_411 (O_411,N_24174,N_24907);
and UO_412 (O_412,N_23837,N_23758);
nand UO_413 (O_413,N_24782,N_22651);
or UO_414 (O_414,N_22637,N_24500);
nor UO_415 (O_415,N_24252,N_23612);
nand UO_416 (O_416,N_22932,N_24991);
and UO_417 (O_417,N_24240,N_23479);
nand UO_418 (O_418,N_23476,N_24018);
nor UO_419 (O_419,N_22742,N_24217);
and UO_420 (O_420,N_24780,N_24981);
and UO_421 (O_421,N_22861,N_24347);
nand UO_422 (O_422,N_22527,N_24550);
or UO_423 (O_423,N_23639,N_23591);
and UO_424 (O_424,N_23407,N_22535);
and UO_425 (O_425,N_22721,N_22632);
xor UO_426 (O_426,N_23642,N_23410);
or UO_427 (O_427,N_23961,N_22634);
nand UO_428 (O_428,N_22561,N_23516);
nand UO_429 (O_429,N_23078,N_22908);
nor UO_430 (O_430,N_22762,N_23260);
nand UO_431 (O_431,N_24928,N_22602);
nor UO_432 (O_432,N_24798,N_22621);
nor UO_433 (O_433,N_23671,N_23398);
nor UO_434 (O_434,N_23132,N_23792);
nand UO_435 (O_435,N_23831,N_22822);
or UO_436 (O_436,N_23588,N_23111);
or UO_437 (O_437,N_24651,N_24704);
xor UO_438 (O_438,N_24598,N_24973);
nand UO_439 (O_439,N_23623,N_23858);
and UO_440 (O_440,N_24493,N_23112);
nor UO_441 (O_441,N_23566,N_23484);
or UO_442 (O_442,N_23229,N_23907);
nand UO_443 (O_443,N_24796,N_23693);
and UO_444 (O_444,N_22868,N_24231);
or UO_445 (O_445,N_24624,N_24108);
and UO_446 (O_446,N_23353,N_24391);
and UO_447 (O_447,N_22993,N_24227);
nor UO_448 (O_448,N_23581,N_24037);
or UO_449 (O_449,N_23160,N_24738);
nor UO_450 (O_450,N_23246,N_24362);
or UO_451 (O_451,N_24288,N_22885);
and UO_452 (O_452,N_23127,N_23319);
nand UO_453 (O_453,N_23182,N_22516);
nor UO_454 (O_454,N_24683,N_23013);
or UO_455 (O_455,N_23129,N_23565);
nand UO_456 (O_456,N_22700,N_23881);
and UO_457 (O_457,N_24802,N_24585);
and UO_458 (O_458,N_22926,N_23830);
and UO_459 (O_459,N_23510,N_24089);
nor UO_460 (O_460,N_24025,N_24159);
and UO_461 (O_461,N_23972,N_23921);
nor UO_462 (O_462,N_24736,N_23512);
or UO_463 (O_463,N_24354,N_23770);
nand UO_464 (O_464,N_22967,N_22795);
xnor UO_465 (O_465,N_23779,N_24001);
nor UO_466 (O_466,N_23158,N_24960);
or UO_467 (O_467,N_23403,N_22801);
nand UO_468 (O_468,N_24933,N_24827);
and UO_469 (O_469,N_23732,N_22747);
or UO_470 (O_470,N_23862,N_23718);
xor UO_471 (O_471,N_24929,N_24505);
or UO_472 (O_472,N_24273,N_24119);
or UO_473 (O_473,N_24270,N_24407);
nor UO_474 (O_474,N_24480,N_24637);
nor UO_475 (O_475,N_22978,N_24322);
nand UO_476 (O_476,N_23376,N_24744);
nand UO_477 (O_477,N_23437,N_24021);
and UO_478 (O_478,N_23709,N_23204);
nor UO_479 (O_479,N_24879,N_23650);
and UO_480 (O_480,N_22600,N_24253);
or UO_481 (O_481,N_24062,N_24148);
and UO_482 (O_482,N_22756,N_23491);
nand UO_483 (O_483,N_22554,N_24551);
nand UO_484 (O_484,N_24113,N_24363);
xor UO_485 (O_485,N_23888,N_23680);
or UO_486 (O_486,N_24035,N_23884);
nand UO_487 (O_487,N_24142,N_24416);
nand UO_488 (O_488,N_22628,N_24600);
nand UO_489 (O_489,N_22755,N_24225);
nand UO_490 (O_490,N_24054,N_23846);
and UO_491 (O_491,N_24236,N_23652);
or UO_492 (O_492,N_24647,N_22779);
or UO_493 (O_493,N_23622,N_24727);
or UO_494 (O_494,N_23788,N_24087);
nand UO_495 (O_495,N_24689,N_24272);
or UO_496 (O_496,N_23909,N_24070);
nor UO_497 (O_497,N_24139,N_23514);
and UO_498 (O_498,N_24705,N_24977);
nand UO_499 (O_499,N_22673,N_24648);
nand UO_500 (O_500,N_24118,N_23729);
or UO_501 (O_501,N_24316,N_24125);
nand UO_502 (O_502,N_24914,N_24956);
nand UO_503 (O_503,N_23219,N_23849);
or UO_504 (O_504,N_22833,N_23649);
nand UO_505 (O_505,N_24836,N_24545);
or UO_506 (O_506,N_22647,N_24329);
nor UO_507 (O_507,N_24592,N_22921);
or UO_508 (O_508,N_24838,N_24571);
xnor UO_509 (O_509,N_23137,N_24721);
and UO_510 (O_510,N_24762,N_22902);
nor UO_511 (O_511,N_23176,N_24842);
nor UO_512 (O_512,N_22976,N_22563);
nand UO_513 (O_513,N_23458,N_23911);
or UO_514 (O_514,N_22615,N_22577);
nor UO_515 (O_515,N_22794,N_24056);
nor UO_516 (O_516,N_23104,N_23991);
nor UO_517 (O_517,N_23162,N_23563);
nand UO_518 (O_518,N_23242,N_24349);
nor UO_519 (O_519,N_22802,N_23307);
or UO_520 (O_520,N_24408,N_23628);
nor UO_521 (O_521,N_22718,N_22748);
nor UO_522 (O_522,N_22860,N_24553);
or UO_523 (O_523,N_23679,N_24484);
and UO_524 (O_524,N_24023,N_22935);
and UO_525 (O_525,N_23905,N_23748);
and UO_526 (O_526,N_23613,N_23686);
nand UO_527 (O_527,N_22911,N_22713);
or UO_528 (O_528,N_23672,N_24478);
or UO_529 (O_529,N_23027,N_24594);
nand UO_530 (O_530,N_24230,N_22812);
or UO_531 (O_531,N_24081,N_24679);
or UO_532 (O_532,N_23611,N_23802);
nand UO_533 (O_533,N_23620,N_24591);
nand UO_534 (O_534,N_22511,N_23383);
and UO_535 (O_535,N_23031,N_24337);
nor UO_536 (O_536,N_23199,N_24431);
or UO_537 (O_537,N_24833,N_24007);
and UO_538 (O_538,N_24269,N_23122);
nand UO_539 (O_539,N_23350,N_24629);
or UO_540 (O_540,N_23370,N_24447);
nand UO_541 (O_541,N_23561,N_23564);
nor UO_542 (O_542,N_23189,N_23258);
nand UO_543 (O_543,N_24228,N_24146);
and UO_544 (O_544,N_22549,N_24121);
or UO_545 (O_545,N_24808,N_23946);
nor UO_546 (O_546,N_23451,N_24235);
nand UO_547 (O_547,N_24642,N_22578);
nand UO_548 (O_548,N_24659,N_24321);
and UO_549 (O_549,N_24947,N_24610);
nor UO_550 (O_550,N_24352,N_23590);
nor UO_551 (O_551,N_24902,N_24050);
or UO_552 (O_552,N_22653,N_24190);
or UO_553 (O_553,N_23793,N_22506);
nand UO_554 (O_554,N_22716,N_22807);
nand UO_555 (O_555,N_24916,N_24153);
or UO_556 (O_556,N_23896,N_23098);
and UO_557 (O_557,N_23654,N_24456);
or UO_558 (O_558,N_23024,N_23015);
nor UO_559 (O_559,N_24745,N_24162);
nand UO_560 (O_560,N_22951,N_22774);
or UO_561 (O_561,N_23406,N_24411);
or UO_562 (O_562,N_23543,N_24084);
and UO_563 (O_563,N_24166,N_24777);
or UO_564 (O_564,N_24788,N_24626);
nand UO_565 (O_565,N_23091,N_23254);
nor UO_566 (O_566,N_23030,N_23712);
and UO_567 (O_567,N_22708,N_23927);
and UO_568 (O_568,N_23382,N_23235);
nand UO_569 (O_569,N_23752,N_24002);
nand UO_570 (O_570,N_24848,N_24093);
and UO_571 (O_571,N_22502,N_24925);
or UO_572 (O_572,N_23726,N_24355);
or UO_573 (O_573,N_23419,N_23455);
nand UO_574 (O_574,N_24711,N_24862);
and UO_575 (O_575,N_22788,N_24502);
or UO_576 (O_576,N_24525,N_22533);
nor UO_577 (O_577,N_22975,N_23174);
nand UO_578 (O_578,N_24837,N_22754);
nand UO_579 (O_579,N_24922,N_24955);
or UO_580 (O_580,N_24760,N_23751);
or UO_581 (O_581,N_23237,N_24994);
and UO_582 (O_582,N_23873,N_23486);
nor UO_583 (O_583,N_24953,N_24028);
nand UO_584 (O_584,N_23517,N_22957);
or UO_585 (O_585,N_23576,N_24882);
and UO_586 (O_586,N_22622,N_23436);
and UO_587 (O_587,N_22585,N_24719);
nor UO_588 (O_588,N_22909,N_22736);
nand UO_589 (O_589,N_23836,N_24111);
nand UO_590 (O_590,N_23092,N_24544);
nand UO_591 (O_591,N_24198,N_24983);
nor UO_592 (O_592,N_24921,N_23908);
nor UO_593 (O_593,N_22940,N_22559);
or UO_594 (O_594,N_23444,N_23501);
or UO_595 (O_595,N_23780,N_24749);
nand UO_596 (O_596,N_23362,N_23996);
nor UO_597 (O_597,N_22881,N_24556);
nand UO_598 (O_598,N_23173,N_23234);
nand UO_599 (O_599,N_23487,N_23377);
nor UO_600 (O_600,N_22793,N_22790);
and UO_601 (O_601,N_22744,N_24767);
nor UO_602 (O_602,N_23179,N_24284);
or UO_603 (O_603,N_24256,N_22867);
and UO_604 (O_604,N_23940,N_23393);
and UO_605 (O_605,N_22719,N_24029);
and UO_606 (O_606,N_23465,N_24906);
or UO_607 (O_607,N_24423,N_24430);
nand UO_608 (O_608,N_24060,N_24859);
nand UO_609 (O_609,N_24064,N_24086);
nor UO_610 (O_610,N_24681,N_24486);
nand UO_611 (O_611,N_23367,N_24931);
nor UO_612 (O_612,N_23567,N_24631);
nand UO_613 (O_613,N_23449,N_24507);
or UO_614 (O_614,N_24662,N_23188);
nor UO_615 (O_615,N_23723,N_24510);
and UO_616 (O_616,N_23635,N_24067);
or UO_617 (O_617,N_23390,N_22897);
nor UO_618 (O_618,N_22586,N_23948);
nand UO_619 (O_619,N_24676,N_23975);
xnor UO_620 (O_620,N_24881,N_24772);
or UO_621 (O_621,N_24913,N_24987);
nand UO_622 (O_622,N_23809,N_24940);
nor UO_623 (O_623,N_24888,N_22777);
nor UO_624 (O_624,N_24395,N_23700);
or UO_625 (O_625,N_22949,N_24099);
nand UO_626 (O_626,N_22880,N_23697);
nor UO_627 (O_627,N_22745,N_23150);
and UO_628 (O_628,N_23375,N_24396);
nor UO_629 (O_629,N_22635,N_23660);
nand UO_630 (O_630,N_22536,N_24218);
nor UO_631 (O_631,N_22837,N_24382);
nand UO_632 (O_632,N_24926,N_24743);
or UO_633 (O_633,N_22849,N_24012);
nand UO_634 (O_634,N_22884,N_23161);
and UO_635 (O_635,N_23036,N_23274);
nand UO_636 (O_636,N_23740,N_24374);
nor UO_637 (O_637,N_22738,N_22598);
nor UO_638 (O_638,N_22715,N_24492);
nand UO_639 (O_639,N_23044,N_22530);
and UO_640 (O_640,N_22771,N_23580);
and UO_641 (O_641,N_23695,N_24559);
nor UO_642 (O_642,N_24937,N_23829);
or UO_643 (O_643,N_23222,N_23100);
nor UO_644 (O_644,N_23251,N_24393);
or UO_645 (O_645,N_23877,N_24077);
nand UO_646 (O_646,N_23256,N_22941);
or UO_647 (O_647,N_23427,N_23197);
and UO_648 (O_648,N_23875,N_22558);
nor UO_649 (O_649,N_24338,N_22995);
and UO_650 (O_650,N_22847,N_24117);
or UO_651 (O_651,N_23894,N_24378);
nand UO_652 (O_652,N_23811,N_23177);
nand UO_653 (O_653,N_24441,N_24201);
or UO_654 (O_654,N_22959,N_24649);
nand UO_655 (O_655,N_24549,N_23147);
xor UO_656 (O_656,N_22854,N_22619);
and UO_657 (O_657,N_24527,N_23760);
and UO_658 (O_658,N_24978,N_23262);
and UO_659 (O_659,N_23266,N_22510);
or UO_660 (O_660,N_24340,N_23298);
and UO_661 (O_661,N_24812,N_24068);
and UO_662 (O_662,N_22799,N_24248);
and UO_663 (O_663,N_23159,N_23958);
nor UO_664 (O_664,N_23727,N_22687);
nor UO_665 (O_665,N_23614,N_24870);
and UO_666 (O_666,N_23600,N_23966);
or UO_667 (O_667,N_24220,N_23291);
nand UO_668 (O_668,N_22599,N_24157);
or UO_669 (O_669,N_24290,N_23817);
xnor UO_670 (O_670,N_22617,N_23575);
or UO_671 (O_671,N_24516,N_23070);
nand UO_672 (O_672,N_22815,N_23903);
nand UO_673 (O_673,N_24951,N_24453);
or UO_674 (O_674,N_23766,N_22851);
or UO_675 (O_675,N_24359,N_23949);
nand UO_676 (O_676,N_24520,N_23302);
or UO_677 (O_677,N_24518,N_24669);
nor UO_678 (O_678,N_24092,N_23850);
nor UO_679 (O_679,N_23233,N_23925);
and UO_680 (O_680,N_24786,N_22720);
nor UO_681 (O_681,N_23037,N_23703);
or UO_682 (O_682,N_23657,N_24791);
and UO_683 (O_683,N_23920,N_24465);
or UO_684 (O_684,N_23771,N_24454);
nor UO_685 (O_685,N_22686,N_23902);
and UO_686 (O_686,N_22569,N_22811);
nand UO_687 (O_687,N_23602,N_24203);
and UO_688 (O_688,N_22531,N_22520);
xnor UO_689 (O_689,N_23255,N_24427);
nand UO_690 (O_690,N_24415,N_24302);
nand UO_691 (O_691,N_23211,N_22517);
and UO_692 (O_692,N_23494,N_23835);
nand UO_693 (O_693,N_22818,N_23178);
nor UO_694 (O_694,N_24013,N_24532);
nand UO_695 (O_695,N_23355,N_23003);
nor UO_696 (O_696,N_22618,N_22896);
xor UO_697 (O_697,N_24932,N_24488);
nor UO_698 (O_698,N_23545,N_23524);
nor UO_699 (O_699,N_24768,N_24843);
or UO_700 (O_700,N_23730,N_24458);
nand UO_701 (O_701,N_22798,N_24797);
nor UO_702 (O_702,N_22553,N_24672);
nor UO_703 (O_703,N_23539,N_23750);
nor UO_704 (O_704,N_24129,N_24644);
or UO_705 (O_705,N_24778,N_23077);
or UO_706 (O_706,N_23808,N_22734);
or UO_707 (O_707,N_24589,N_22595);
nor UO_708 (O_708,N_22562,N_23799);
and UO_709 (O_709,N_24593,N_23124);
nand UO_710 (O_710,N_24943,N_24971);
nand UO_711 (O_711,N_22846,N_23970);
nand UO_712 (O_712,N_24372,N_23914);
or UO_713 (O_713,N_24785,N_23523);
nor UO_714 (O_714,N_24123,N_24521);
nor UO_715 (O_715,N_23386,N_24282);
or UO_716 (O_716,N_24668,N_22989);
nor UO_717 (O_717,N_23918,N_22766);
nor UO_718 (O_718,N_23534,N_22630);
nor UO_719 (O_719,N_24641,N_24279);
and UO_720 (O_720,N_23520,N_22866);
nand UO_721 (O_721,N_22714,N_23053);
nor UO_722 (O_722,N_23378,N_24789);
or UO_723 (O_723,N_23073,N_24739);
xor UO_724 (O_724,N_23932,N_24243);
or UO_725 (O_725,N_24995,N_23492);
and UO_726 (O_726,N_23987,N_22904);
or UO_727 (O_727,N_23311,N_23332);
nand UO_728 (O_728,N_24110,N_23329);
and UO_729 (O_729,N_23557,N_23851);
and UO_730 (O_730,N_22895,N_24429);
or UO_731 (O_731,N_24265,N_22609);
nand UO_732 (O_732,N_22726,N_24336);
nand UO_733 (O_733,N_24171,N_24850);
nand UO_734 (O_734,N_24435,N_24660);
and UO_735 (O_735,N_23007,N_23490);
nor UO_736 (O_736,N_24115,N_24306);
and UO_737 (O_737,N_23434,N_24538);
nor UO_738 (O_738,N_23295,N_24755);
or UO_739 (O_739,N_24801,N_22605);
nor UO_740 (O_740,N_23854,N_24847);
nand UO_741 (O_741,N_23418,N_24904);
or UO_742 (O_742,N_24242,N_23633);
or UO_743 (O_743,N_23965,N_23126);
and UO_744 (O_744,N_23670,N_24399);
nand UO_745 (O_745,N_22987,N_24237);
xor UO_746 (O_746,N_23216,N_22590);
and UO_747 (O_747,N_23001,N_23656);
or UO_748 (O_748,N_23275,N_24195);
nand UO_749 (O_749,N_22724,N_24604);
and UO_750 (O_750,N_24634,N_24009);
xor UO_751 (O_751,N_23947,N_23181);
or UO_752 (O_752,N_23263,N_23632);
nor UO_753 (O_753,N_22945,N_23366);
nor UO_754 (O_754,N_24769,N_24414);
nand UO_755 (O_755,N_22636,N_23882);
xor UO_756 (O_756,N_23064,N_23710);
and UO_757 (O_757,N_23215,N_23587);
or UO_758 (O_758,N_22883,N_23839);
and UO_759 (O_759,N_23059,N_24266);
and UO_760 (O_760,N_23525,N_22608);
or UO_761 (O_761,N_23538,N_23550);
nand UO_762 (O_762,N_23645,N_24886);
nor UO_763 (O_763,N_23806,N_23627);
nor UO_764 (O_764,N_22582,N_23664);
or UO_765 (O_765,N_24613,N_22645);
or UO_766 (O_766,N_23781,N_23519);
or UO_767 (O_767,N_24889,N_22874);
and UO_768 (O_768,N_23777,N_22973);
or UO_769 (O_769,N_23798,N_23327);
or UO_770 (O_770,N_23384,N_23507);
nand UO_771 (O_771,N_22984,N_22662);
or UO_772 (O_772,N_24319,N_23782);
or UO_773 (O_773,N_24194,N_22968);
nor UO_774 (O_774,N_23317,N_23619);
nand UO_775 (O_775,N_23226,N_24857);
nand UO_776 (O_776,N_23279,N_22592);
or UO_777 (O_777,N_24958,N_24608);
nand UO_778 (O_778,N_24178,N_24017);
xor UO_779 (O_779,N_24622,N_22675);
xnor UO_780 (O_780,N_24221,N_22792);
and UO_781 (O_781,N_24301,N_24540);
nand UO_782 (O_782,N_23082,N_23456);
or UO_783 (O_783,N_24599,N_24866);
nor UO_784 (O_784,N_23800,N_22566);
and UO_785 (O_785,N_23303,N_24787);
or UO_786 (O_786,N_24481,N_24673);
or UO_787 (O_787,N_23102,N_24670);
or UO_788 (O_788,N_22784,N_23108);
and UO_789 (O_789,N_24996,N_24163);
nand UO_790 (O_790,N_22972,N_23442);
xor UO_791 (O_791,N_24079,N_24274);
or UO_792 (O_792,N_24897,N_24188);
nand UO_793 (O_793,N_24967,N_23409);
or UO_794 (O_794,N_22912,N_23068);
nand UO_795 (O_795,N_22729,N_24580);
and UO_796 (O_796,N_23010,N_23285);
nor UO_797 (O_797,N_22565,N_23720);
nor UO_798 (O_798,N_23048,N_23466);
or UO_799 (O_799,N_22557,N_23014);
or UO_800 (O_800,N_24425,N_24845);
nand UO_801 (O_801,N_23363,N_22532);
and UO_802 (O_802,N_24419,N_24805);
and UO_803 (O_803,N_22737,N_24192);
and UO_804 (O_804,N_24294,N_24839);
and UO_805 (O_805,N_23062,N_23028);
nor UO_806 (O_806,N_22982,N_23785);
or UO_807 (O_807,N_22730,N_24455);
and UO_808 (O_808,N_23213,N_23310);
nand UO_809 (O_809,N_24332,N_24919);
or UO_810 (O_810,N_24278,N_23944);
xor UO_811 (O_811,N_23321,N_24173);
nand UO_812 (O_812,N_24877,N_24915);
or UO_813 (O_813,N_23971,N_24467);
and UO_814 (O_814,N_22688,N_24402);
and UO_815 (O_815,N_24548,N_24576);
xnor UO_816 (O_816,N_24003,N_22772);
or UO_817 (O_817,N_23998,N_24863);
nand UO_818 (O_818,N_23526,N_24268);
and UO_819 (O_819,N_22758,N_24970);
nand UO_820 (O_820,N_23506,N_23509);
and UO_821 (O_821,N_24849,N_24835);
and UO_822 (O_822,N_22638,N_24583);
nor UO_823 (O_823,N_24360,N_23011);
nand UO_824 (O_824,N_24766,N_22655);
and UO_825 (O_825,N_24376,N_24680);
and UO_826 (O_826,N_24471,N_22827);
and UO_827 (O_827,N_22848,N_24918);
or UO_828 (O_828,N_24596,N_24821);
and UO_829 (O_829,N_22791,N_24333);
or UO_830 (O_830,N_23471,N_22817);
or UO_831 (O_831,N_23957,N_24043);
nand UO_832 (O_832,N_24722,N_23206);
and UO_833 (O_833,N_22503,N_24061);
nand UO_834 (O_834,N_24726,N_24517);
or UO_835 (O_835,N_22830,N_24715);
or UO_836 (O_836,N_24185,N_24154);
nand UO_837 (O_837,N_23879,N_23772);
nand UO_838 (O_838,N_24666,N_24204);
nor UO_839 (O_839,N_23956,N_23892);
or UO_840 (O_840,N_24167,N_22689);
nand UO_841 (O_841,N_24223,N_22560);
and UO_842 (O_842,N_24844,N_23128);
nand UO_843 (O_843,N_23913,N_24464);
nor UO_844 (O_844,N_24688,N_22528);
nor UO_845 (O_845,N_23435,N_23528);
and UO_846 (O_846,N_24044,N_24144);
nor UO_847 (O_847,N_24878,N_23448);
nor UO_848 (O_848,N_24854,N_23067);
nand UO_849 (O_849,N_24765,N_22757);
nand UO_850 (O_850,N_23136,N_24156);
nor UO_851 (O_851,N_24389,N_24774);
nor UO_852 (O_852,N_24394,N_23006);
nor UO_853 (O_853,N_22856,N_23536);
or UO_854 (O_854,N_24503,N_24006);
nand UO_855 (O_855,N_24027,N_22544);
nor UO_856 (O_856,N_24369,N_24262);
nand UO_857 (O_857,N_24358,N_24103);
nor UO_858 (O_858,N_23259,N_24386);
and UO_859 (O_859,N_23606,N_22805);
nand UO_860 (O_860,N_23722,N_23250);
or UO_861 (O_861,N_24701,N_23205);
nor UO_862 (O_862,N_22927,N_23305);
and UO_863 (O_863,N_23061,N_24590);
and UO_864 (O_864,N_22814,N_24310);
nand UO_865 (O_865,N_24539,N_22614);
nand UO_866 (O_866,N_24277,N_22521);
or UO_867 (O_867,N_23135,N_23864);
nor UO_868 (O_868,N_22939,N_24042);
and UO_869 (O_869,N_24612,N_24737);
nand UO_870 (O_870,N_22816,N_22555);
and UO_871 (O_871,N_23169,N_22819);
and UO_872 (O_872,N_22918,N_24504);
nor UO_873 (O_873,N_24617,N_23105);
nor UO_874 (O_874,N_22942,N_24799);
nand UO_875 (O_875,N_23631,N_23725);
nor UO_876 (O_876,N_22785,N_24515);
nand UO_877 (O_877,N_23089,N_22541);
xnor UO_878 (O_878,N_23473,N_24128);
and UO_879 (O_879,N_24942,N_22584);
or UO_880 (O_880,N_22534,N_23416);
and UO_881 (O_881,N_22960,N_22643);
and UO_882 (O_882,N_22886,N_24215);
nand UO_883 (O_883,N_22712,N_23387);
and UO_884 (O_884,N_22606,N_23551);
nand UO_885 (O_885,N_24147,N_24436);
and UO_886 (O_886,N_24112,N_24790);
nor UO_887 (O_887,N_24899,N_24057);
nor UO_888 (O_888,N_24840,N_23281);
nand UO_889 (O_889,N_24368,N_24748);
nor UO_890 (O_890,N_22985,N_22820);
nand UO_891 (O_891,N_24232,N_23270);
nand UO_892 (O_892,N_24387,N_22692);
nor UO_893 (O_893,N_22576,N_22889);
or UO_894 (O_894,N_24356,N_23094);
or UO_895 (O_895,N_24026,N_24344);
nor UO_896 (O_896,N_23245,N_22969);
nand UO_897 (O_897,N_23450,N_23086);
nand UO_898 (O_898,N_23844,N_24244);
nor UO_899 (O_899,N_24698,N_23333);
or UO_900 (O_900,N_23323,N_24320);
or UO_901 (O_901,N_22518,N_22760);
nor UO_902 (O_902,N_24342,N_23133);
nand UO_903 (O_903,N_23583,N_22948);
nand UO_904 (O_904,N_24543,N_23763);
nor UO_905 (O_905,N_23334,N_23891);
nand UO_906 (O_906,N_24051,N_24930);
and UO_907 (O_907,N_23572,N_24187);
or UO_908 (O_908,N_23502,N_23604);
or UO_909 (O_909,N_24072,N_22936);
or UO_910 (O_910,N_24160,N_22986);
nand UO_911 (O_911,N_22933,N_23841);
and UO_912 (O_912,N_22500,N_24706);
and UO_913 (O_913,N_23462,N_23755);
or UO_914 (O_914,N_23761,N_23457);
or UO_915 (O_915,N_22955,N_24206);
nor UO_916 (O_916,N_22783,N_24312);
xor UO_917 (O_917,N_22871,N_23404);
and UO_918 (O_918,N_23360,N_23212);
nor UO_919 (O_919,N_23601,N_22627);
nand UO_920 (O_920,N_24283,N_24114);
nor UO_921 (O_921,N_22864,N_24834);
and UO_922 (O_922,N_22980,N_24233);
nor UO_923 (O_923,N_24133,N_23340);
or UO_924 (O_924,N_24137,N_24757);
and UO_925 (O_925,N_22966,N_24048);
nor UO_926 (O_926,N_24296,N_23293);
or UO_927 (O_927,N_24824,N_24687);
nor UO_928 (O_928,N_24567,N_24908);
and UO_929 (O_929,N_23789,N_24379);
or UO_930 (O_930,N_23441,N_22698);
and UO_931 (O_931,N_24011,N_24497);
nand UO_932 (O_932,N_22504,N_23533);
nand UO_933 (O_933,N_23579,N_24883);
and UO_934 (O_934,N_24874,N_23079);
nand UO_935 (O_935,N_24085,N_24759);
nand UO_936 (O_936,N_23666,N_24990);
nand UO_937 (O_937,N_24753,N_22776);
xnor UO_938 (O_938,N_24623,N_22732);
or UO_939 (O_939,N_23570,N_24712);
nand UO_940 (O_940,N_24400,N_23535);
nand UO_941 (O_941,N_22857,N_22548);
nand UO_942 (O_942,N_24763,N_24959);
nand UO_943 (O_943,N_23813,N_23870);
and UO_944 (O_944,N_23503,N_24075);
nand UO_945 (O_945,N_24603,N_24501);
nand UO_946 (O_946,N_23005,N_23582);
and UO_947 (O_947,N_24720,N_23318);
or UO_948 (O_948,N_24989,N_22865);
nand UO_949 (O_949,N_22944,N_24287);
nand UO_950 (O_950,N_22693,N_22999);
nor UO_951 (O_951,N_23236,N_24432);
nand UO_952 (O_952,N_24420,N_24747);
or UO_953 (O_953,N_23364,N_22525);
or UO_954 (O_954,N_23447,N_23240);
and UO_955 (O_955,N_23708,N_23853);
nor UO_956 (O_956,N_23742,N_24255);
and UO_957 (O_957,N_24547,N_22556);
nor UO_958 (O_958,N_23428,N_24291);
nand UO_959 (O_959,N_22706,N_23852);
and UO_960 (O_960,N_24657,N_24161);
nor UO_961 (O_961,N_23641,N_23208);
and UO_962 (O_962,N_22573,N_23979);
nand UO_963 (O_963,N_24169,N_24709);
nor UO_964 (O_964,N_22665,N_23716);
nor UO_965 (O_965,N_23369,N_22810);
nor UO_966 (O_966,N_22898,N_23941);
nor UO_967 (O_967,N_24091,N_23426);
and UO_968 (O_968,N_22649,N_23803);
nor UO_969 (O_969,N_22728,N_24459);
and UO_970 (O_970,N_23394,N_23562);
nand UO_971 (O_971,N_24088,N_24371);
and UO_972 (O_972,N_23337,N_24150);
or UO_973 (O_973,N_23019,N_23916);
nand UO_974 (O_974,N_24036,N_23549);
and UO_975 (O_975,N_23163,N_24671);
nor UO_976 (O_976,N_23959,N_23365);
nand UO_977 (O_977,N_23719,N_22894);
xnor UO_978 (O_978,N_23791,N_24261);
or UO_979 (O_979,N_23744,N_22648);
nand UO_980 (O_980,N_24384,N_24633);
and UO_981 (O_981,N_22526,N_24098);
or UO_982 (O_982,N_24901,N_24826);
or UO_983 (O_983,N_22681,N_23110);
nor UO_984 (O_984,N_22751,N_22931);
or UO_985 (O_985,N_23555,N_24485);
or UO_986 (O_986,N_23696,N_23468);
nor UO_987 (O_987,N_23843,N_23895);
nand UO_988 (O_988,N_23185,N_24191);
or UO_989 (O_989,N_24533,N_22568);
nor UO_990 (O_990,N_24472,N_22923);
nand UO_991 (O_991,N_23626,N_24741);
or UO_992 (O_992,N_23187,N_22877);
nor UO_993 (O_993,N_22644,N_24331);
nor UO_994 (O_994,N_22641,N_24380);
or UO_995 (O_995,N_24758,N_24792);
and UO_996 (O_996,N_23041,N_24952);
or UO_997 (O_997,N_23685,N_24852);
nand UO_998 (O_998,N_23264,N_24731);
and UO_999 (O_999,N_23814,N_24950);
or UO_1000 (O_1000,N_23121,N_24437);
nand UO_1001 (O_1001,N_24071,N_24390);
and UO_1002 (O_1002,N_22661,N_23301);
and UO_1003 (O_1003,N_24910,N_22872);
nor UO_1004 (O_1004,N_24636,N_23728);
nand UO_1005 (O_1005,N_23743,N_23085);
nor UO_1006 (O_1006,N_22679,N_24249);
nand UO_1007 (O_1007,N_23953,N_23863);
nand UO_1008 (O_1008,N_22538,N_23774);
or UO_1009 (O_1009,N_24038,N_22890);
or UO_1010 (O_1010,N_24381,N_23976);
nand UO_1011 (O_1011,N_22739,N_23974);
nand UO_1012 (O_1012,N_23244,N_22652);
and UO_1013 (O_1013,N_23842,N_24898);
nor UO_1014 (O_1014,N_22740,N_24754);
or UO_1015 (O_1015,N_22806,N_24853);
or UO_1016 (O_1016,N_24998,N_24448);
nand UO_1017 (O_1017,N_24341,N_24149);
and UO_1018 (O_1018,N_24555,N_24047);
or UO_1019 (O_1019,N_24734,N_23691);
and UO_1020 (O_1020,N_24205,N_23381);
or UO_1021 (O_1021,N_23257,N_23096);
or UO_1022 (O_1022,N_24700,N_22529);
and UO_1023 (O_1023,N_22564,N_24343);
nor UO_1024 (O_1024,N_24073,N_22575);
or UO_1025 (O_1025,N_24530,N_22843);
nor UO_1026 (O_1026,N_23115,N_22593);
and UO_1027 (O_1027,N_23812,N_24528);
xor UO_1028 (O_1028,N_23299,N_23559);
nor UO_1029 (O_1029,N_24410,N_23796);
nand UO_1030 (O_1030,N_24563,N_23239);
nand UO_1031 (O_1031,N_24999,N_23546);
nand UO_1032 (O_1032,N_23230,N_22888);
and UO_1033 (O_1033,N_23107,N_22537);
nand UO_1034 (O_1034,N_23893,N_23292);
or UO_1035 (O_1035,N_22925,N_24939);
nand UO_1036 (O_1036,N_23603,N_23889);
nand UO_1037 (O_1037,N_23372,N_24542);
nor UO_1038 (O_1038,N_23183,N_23985);
or UO_1039 (O_1039,N_24568,N_23391);
nand UO_1040 (O_1040,N_23878,N_24982);
and UO_1041 (O_1041,N_22878,N_24941);
nand UO_1042 (O_1042,N_24708,N_23989);
nand UO_1043 (O_1043,N_24993,N_23433);
or UO_1044 (O_1044,N_23099,N_24814);
nor UO_1045 (O_1045,N_22828,N_23662);
or UO_1046 (O_1046,N_22597,N_24923);
nand UO_1047 (O_1047,N_22727,N_23335);
and UO_1048 (O_1048,N_22695,N_24101);
nand UO_1049 (O_1049,N_22604,N_23341);
nor UO_1050 (O_1050,N_22953,N_23684);
nor UO_1051 (O_1051,N_24059,N_22974);
nand UO_1052 (O_1052,N_23663,N_23678);
nand UO_1053 (O_1053,N_22768,N_24690);
nor UO_1054 (O_1054,N_24714,N_22694);
nor UO_1055 (O_1055,N_24846,N_24588);
and UO_1056 (O_1056,N_23648,N_22709);
nor UO_1057 (O_1057,N_24822,N_24120);
nand UO_1058 (O_1058,N_22710,N_23832);
nor UO_1059 (O_1059,N_24033,N_22509);
and UO_1060 (O_1060,N_23597,N_23644);
or UO_1061 (O_1061,N_24015,N_23452);
and UO_1062 (O_1062,N_23917,N_23155);
and UO_1063 (O_1063,N_24298,N_24895);
and UO_1064 (O_1064,N_23819,N_23745);
nor UO_1065 (O_1065,N_24529,N_24984);
nor UO_1066 (O_1066,N_24275,N_23930);
nand UO_1067 (O_1067,N_24975,N_24675);
nor UO_1068 (O_1068,N_23764,N_24172);
nand UO_1069 (O_1069,N_22678,N_22869);
nand UO_1070 (O_1070,N_24770,N_22642);
and UO_1071 (O_1071,N_23765,N_23890);
or UO_1072 (O_1072,N_23253,N_24587);
nor UO_1073 (O_1073,N_23249,N_22612);
nand UO_1074 (O_1074,N_23489,N_24155);
or UO_1075 (O_1075,N_24891,N_24096);
nand UO_1076 (O_1076,N_23531,N_23934);
nand UO_1077 (O_1077,N_23969,N_23395);
nor UO_1078 (O_1078,N_23034,N_23901);
or UO_1079 (O_1079,N_24292,N_24554);
nand UO_1080 (O_1080,N_23043,N_24016);
or UO_1081 (O_1081,N_23834,N_24449);
or UO_1082 (O_1082,N_22623,N_24856);
or UO_1083 (O_1083,N_22943,N_23389);
nor UO_1084 (O_1084,N_24463,N_22915);
or UO_1085 (O_1085,N_24506,N_24065);
nand UO_1086 (O_1086,N_24903,N_22870);
xor UO_1087 (O_1087,N_22668,N_23554);
nor UO_1088 (O_1088,N_23201,N_22852);
and UO_1089 (O_1089,N_23634,N_24375);
and UO_1090 (O_1090,N_23289,N_23057);
nand UO_1091 (O_1091,N_24489,N_24729);
xor UO_1092 (O_1092,N_24652,N_23184);
nand UO_1093 (O_1093,N_24442,N_24104);
xor UO_1094 (O_1094,N_23402,N_23880);
and UO_1095 (O_1095,N_23769,N_24872);
and UO_1096 (O_1096,N_22832,N_24397);
nand UO_1097 (O_1097,N_23676,N_23731);
nor UO_1098 (O_1098,N_23060,N_24258);
nor UO_1099 (O_1099,N_24800,N_23558);
and UO_1100 (O_1100,N_23762,N_23286);
nand UO_1101 (O_1101,N_23467,N_22858);
nand UO_1102 (O_1102,N_24677,N_22845);
and UO_1103 (O_1103,N_24295,N_24443);
nand UO_1104 (O_1104,N_23964,N_23861);
or UO_1105 (O_1105,N_23828,N_24728);
nor UO_1106 (O_1106,N_24606,N_24074);
nor UO_1107 (O_1107,N_23711,N_24207);
nor UO_1108 (O_1108,N_23322,N_24303);
nor UO_1109 (O_1109,N_24640,N_23140);
and UO_1110 (O_1110,N_24752,N_24526);
or UO_1111 (O_1111,N_23855,N_23585);
nand UO_1112 (O_1112,N_22667,N_24202);
and UO_1113 (O_1113,N_22610,N_24861);
nand UO_1114 (O_1114,N_24257,N_23058);
or UO_1115 (O_1115,N_23945,N_23694);
nor UO_1116 (O_1116,N_24565,N_22769);
or UO_1117 (O_1117,N_24339,N_22997);
nor UO_1118 (O_1118,N_23868,N_23287);
nor UO_1119 (O_1119,N_22759,N_23673);
nand UO_1120 (O_1120,N_22930,N_22950);
nor UO_1121 (O_1121,N_23051,N_24936);
or UO_1122 (O_1122,N_23148,N_23413);
and UO_1123 (O_1123,N_23361,N_23824);
nand UO_1124 (O_1124,N_23983,N_22765);
nor UO_1125 (O_1125,N_23904,N_24095);
and UO_1126 (O_1126,N_24460,N_23039);
nor UO_1127 (O_1127,N_24513,N_22703);
or UO_1128 (O_1128,N_24564,N_23417);
nand UO_1129 (O_1129,N_23707,N_24214);
nand UO_1130 (O_1130,N_24280,N_24404);
xor UO_1131 (O_1131,N_22591,N_23008);
and UO_1132 (O_1132,N_22731,N_23667);
nor UO_1133 (O_1133,N_22839,N_24961);
nor UO_1134 (O_1134,N_24985,N_24219);
or UO_1135 (O_1135,N_24887,N_24030);
or UO_1136 (O_1136,N_24116,N_24351);
or UO_1137 (O_1137,N_23608,N_23936);
nand UO_1138 (O_1138,N_23313,N_24346);
nand UO_1139 (O_1139,N_22656,N_23640);
and UO_1140 (O_1140,N_23272,N_23919);
nor UO_1141 (O_1141,N_24418,N_24324);
nor UO_1142 (O_1142,N_23860,N_22583);
nand UO_1143 (O_1143,N_23935,N_24439);
or UO_1144 (O_1144,N_24804,N_23962);
nand UO_1145 (O_1145,N_24609,N_23738);
nand UO_1146 (O_1146,N_24865,N_24823);
or UO_1147 (O_1147,N_23553,N_23952);
nand UO_1148 (O_1148,N_23143,N_23141);
or UO_1149 (O_1149,N_23052,N_24046);
xnor UO_1150 (O_1150,N_23153,N_22947);
nor UO_1151 (O_1151,N_23560,N_23055);
and UO_1152 (O_1152,N_22892,N_24725);
xnor UO_1153 (O_1153,N_24300,N_22735);
and UO_1154 (O_1154,N_23653,N_24892);
nor UO_1155 (O_1155,N_22603,N_23504);
and UO_1156 (O_1156,N_23485,N_24132);
and UO_1157 (O_1157,N_23658,N_24107);
nand UO_1158 (O_1158,N_24100,N_23668);
or UO_1159 (O_1159,N_22829,N_24667);
or UO_1160 (O_1160,N_22946,N_24315);
and UO_1161 (O_1161,N_24873,N_23297);
nor UO_1162 (O_1162,N_23924,N_24066);
nor UO_1163 (O_1163,N_24193,N_24239);
nor UO_1164 (O_1164,N_22809,N_22938);
xor UO_1165 (O_1165,N_24293,N_24864);
and UO_1166 (O_1166,N_24560,N_23596);
or UO_1167 (O_1167,N_23065,N_23309);
nand UO_1168 (O_1168,N_23499,N_23113);
and UO_1169 (O_1169,N_24334,N_22882);
nor UO_1170 (O_1170,N_22920,N_24401);
and UO_1171 (O_1171,N_23282,N_24490);
nand UO_1172 (O_1172,N_24247,N_24686);
and UO_1173 (O_1173,N_24222,N_22539);
or UO_1174 (O_1174,N_23495,N_24426);
or UO_1175 (O_1175,N_23252,N_24130);
xnor UO_1176 (O_1176,N_24428,N_24558);
and UO_1177 (O_1177,N_22507,N_24020);
nor UO_1178 (O_1178,N_24578,N_24498);
nand UO_1179 (O_1179,N_23265,N_24552);
and UO_1180 (O_1180,N_24412,N_24168);
nand UO_1181 (O_1181,N_22913,N_23820);
and UO_1182 (O_1182,N_24357,N_22922);
nand UO_1183 (O_1183,N_23342,N_24577);
or UO_1184 (O_1184,N_23734,N_23733);
nand UO_1185 (O_1185,N_23984,N_22581);
nand UO_1186 (O_1186,N_24911,N_24615);
nand UO_1187 (O_1187,N_23778,N_23083);
and UO_1188 (O_1188,N_23993,N_24457);
nor UO_1189 (O_1189,N_22579,N_23273);
nor UO_1190 (O_1190,N_22596,N_22594);
nor UO_1191 (O_1191,N_23625,N_24197);
or UO_1192 (O_1192,N_23392,N_23425);
and UO_1193 (O_1193,N_23994,N_23354);
and UO_1194 (O_1194,N_23687,N_24317);
or UO_1195 (O_1195,N_22702,N_24829);
and UO_1196 (O_1196,N_22992,N_23768);
and UO_1197 (O_1197,N_23933,N_23513);
nor UO_1198 (O_1198,N_23033,N_23331);
and UO_1199 (O_1199,N_22607,N_23721);
nand UO_1200 (O_1200,N_24793,N_23123);
nand UO_1201 (O_1201,N_22601,N_24209);
or UO_1202 (O_1202,N_24152,N_24750);
nand UO_1203 (O_1203,N_23795,N_23268);
and UO_1204 (O_1204,N_23071,N_23568);
nor UO_1205 (O_1205,N_23165,N_24656);
nand UO_1206 (O_1206,N_23977,N_23688);
nand UO_1207 (O_1207,N_24828,N_24561);
nand UO_1208 (O_1208,N_23228,N_23818);
nor UO_1209 (O_1209,N_24586,N_23643);
or UO_1210 (O_1210,N_24164,N_23577);
and UO_1211 (O_1211,N_22855,N_23276);
and UO_1212 (O_1212,N_23906,N_23172);
nor UO_1213 (O_1213,N_24781,N_24335);
and UO_1214 (O_1214,N_24264,N_23320);
or UO_1215 (O_1215,N_24832,N_23045);
or UO_1216 (O_1216,N_23715,N_23125);
or UO_1217 (O_1217,N_24710,N_24716);
and UO_1218 (O_1218,N_23801,N_23368);
nand UO_1219 (O_1219,N_23166,N_23816);
and UO_1220 (O_1220,N_24186,N_23325);
and UO_1221 (O_1221,N_23344,N_23338);
nand UO_1222 (O_1222,N_23527,N_23593);
nor UO_1223 (O_1223,N_22859,N_23463);
and UO_1224 (O_1224,N_23238,N_23221);
nand UO_1225 (O_1225,N_24267,N_22631);
and UO_1226 (O_1226,N_23241,N_24831);
nor UO_1227 (O_1227,N_24569,N_23807);
or UO_1228 (O_1228,N_22743,N_23823);
nand UO_1229 (O_1229,N_23926,N_23151);
and UO_1230 (O_1230,N_24182,N_22797);
nor UO_1231 (O_1231,N_24053,N_24938);
xnor UO_1232 (O_1232,N_23968,N_22824);
nand UO_1233 (O_1233,N_24483,N_24663);
nand UO_1234 (O_1234,N_23469,N_23210);
and UO_1235 (O_1235,N_23840,N_23599);
or UO_1236 (O_1236,N_22780,N_24180);
and UO_1237 (O_1237,N_24584,N_23838);
or UO_1238 (O_1238,N_24234,N_24841);
nand UO_1239 (O_1239,N_22680,N_23346);
or UO_1240 (O_1240,N_22994,N_24536);
nor UO_1241 (O_1241,N_23347,N_23130);
or UO_1242 (O_1242,N_23288,N_22924);
nor UO_1243 (O_1243,N_23922,N_23797);
nand UO_1244 (O_1244,N_24934,N_24602);
and UO_1245 (O_1245,N_24917,N_23629);
nand UO_1246 (O_1246,N_22891,N_22907);
nand UO_1247 (O_1247,N_24138,N_22917);
nor UO_1248 (O_1248,N_22546,N_24131);
and UO_1249 (O_1249,N_23973,N_23735);
nor UO_1250 (O_1250,N_22624,N_23509);
or UO_1251 (O_1251,N_24346,N_23287);
nand UO_1252 (O_1252,N_22764,N_23483);
nor UO_1253 (O_1253,N_24468,N_23632);
nand UO_1254 (O_1254,N_22730,N_23568);
or UO_1255 (O_1255,N_24061,N_23602);
and UO_1256 (O_1256,N_23601,N_22751);
and UO_1257 (O_1257,N_22949,N_22880);
nand UO_1258 (O_1258,N_24176,N_24146);
nor UO_1259 (O_1259,N_23415,N_24755);
nor UO_1260 (O_1260,N_22820,N_22855);
nor UO_1261 (O_1261,N_24575,N_23532);
nor UO_1262 (O_1262,N_24697,N_24504);
nand UO_1263 (O_1263,N_24771,N_24593);
nor UO_1264 (O_1264,N_22934,N_24916);
and UO_1265 (O_1265,N_23856,N_23378);
and UO_1266 (O_1266,N_24438,N_23194);
and UO_1267 (O_1267,N_24959,N_23846);
or UO_1268 (O_1268,N_23084,N_24525);
and UO_1269 (O_1269,N_24721,N_24474);
nand UO_1270 (O_1270,N_23583,N_22867);
and UO_1271 (O_1271,N_22665,N_24338);
or UO_1272 (O_1272,N_23147,N_24042);
and UO_1273 (O_1273,N_23905,N_24607);
or UO_1274 (O_1274,N_24230,N_24016);
nor UO_1275 (O_1275,N_23939,N_24409);
or UO_1276 (O_1276,N_22692,N_23660);
and UO_1277 (O_1277,N_23768,N_23224);
and UO_1278 (O_1278,N_23435,N_23887);
and UO_1279 (O_1279,N_22628,N_23370);
or UO_1280 (O_1280,N_23224,N_23200);
nand UO_1281 (O_1281,N_24255,N_24059);
and UO_1282 (O_1282,N_24986,N_24708);
and UO_1283 (O_1283,N_24546,N_24524);
nand UO_1284 (O_1284,N_23052,N_24452);
or UO_1285 (O_1285,N_22562,N_24233);
or UO_1286 (O_1286,N_24260,N_22733);
or UO_1287 (O_1287,N_24913,N_23032);
nor UO_1288 (O_1288,N_24545,N_22565);
and UO_1289 (O_1289,N_23572,N_23626);
and UO_1290 (O_1290,N_23414,N_23446);
nand UO_1291 (O_1291,N_22700,N_23376);
nand UO_1292 (O_1292,N_23848,N_23455);
or UO_1293 (O_1293,N_23481,N_23310);
nand UO_1294 (O_1294,N_23389,N_23313);
nand UO_1295 (O_1295,N_23786,N_24773);
xor UO_1296 (O_1296,N_22660,N_23346);
nor UO_1297 (O_1297,N_24199,N_23322);
nand UO_1298 (O_1298,N_24563,N_23771);
nor UO_1299 (O_1299,N_24603,N_23490);
or UO_1300 (O_1300,N_22790,N_23025);
nor UO_1301 (O_1301,N_22792,N_24490);
nor UO_1302 (O_1302,N_24492,N_23565);
or UO_1303 (O_1303,N_22846,N_23698);
nor UO_1304 (O_1304,N_24511,N_24611);
and UO_1305 (O_1305,N_24200,N_24952);
nand UO_1306 (O_1306,N_23615,N_24758);
and UO_1307 (O_1307,N_22940,N_22757);
nor UO_1308 (O_1308,N_24860,N_24938);
nor UO_1309 (O_1309,N_23747,N_24460);
nor UO_1310 (O_1310,N_24278,N_24127);
or UO_1311 (O_1311,N_23180,N_24237);
nand UO_1312 (O_1312,N_24685,N_22565);
nand UO_1313 (O_1313,N_24555,N_23702);
nand UO_1314 (O_1314,N_23536,N_23184);
nor UO_1315 (O_1315,N_24624,N_24748);
and UO_1316 (O_1316,N_24231,N_24874);
and UO_1317 (O_1317,N_22934,N_23373);
and UO_1318 (O_1318,N_24080,N_24518);
nand UO_1319 (O_1319,N_22865,N_22843);
or UO_1320 (O_1320,N_24900,N_24105);
xnor UO_1321 (O_1321,N_23598,N_24553);
and UO_1322 (O_1322,N_24704,N_22795);
nand UO_1323 (O_1323,N_24535,N_24159);
or UO_1324 (O_1324,N_22582,N_23632);
nand UO_1325 (O_1325,N_23171,N_22891);
and UO_1326 (O_1326,N_24117,N_22632);
nand UO_1327 (O_1327,N_24661,N_23457);
and UO_1328 (O_1328,N_24773,N_24464);
nor UO_1329 (O_1329,N_24800,N_24974);
nand UO_1330 (O_1330,N_23206,N_24805);
or UO_1331 (O_1331,N_22884,N_22953);
or UO_1332 (O_1332,N_24346,N_24997);
and UO_1333 (O_1333,N_22656,N_22761);
and UO_1334 (O_1334,N_22956,N_22771);
or UO_1335 (O_1335,N_23498,N_23399);
nand UO_1336 (O_1336,N_22654,N_22746);
or UO_1337 (O_1337,N_24120,N_23886);
and UO_1338 (O_1338,N_22872,N_22930);
and UO_1339 (O_1339,N_23117,N_23828);
or UO_1340 (O_1340,N_23431,N_22930);
and UO_1341 (O_1341,N_24359,N_23219);
or UO_1342 (O_1342,N_23168,N_24416);
and UO_1343 (O_1343,N_23386,N_22835);
and UO_1344 (O_1344,N_24644,N_23639);
or UO_1345 (O_1345,N_23605,N_23498);
and UO_1346 (O_1346,N_22897,N_23258);
and UO_1347 (O_1347,N_23592,N_24278);
xor UO_1348 (O_1348,N_23037,N_23356);
or UO_1349 (O_1349,N_23731,N_24742);
nand UO_1350 (O_1350,N_24927,N_24262);
or UO_1351 (O_1351,N_24395,N_24209);
and UO_1352 (O_1352,N_24102,N_24485);
or UO_1353 (O_1353,N_24835,N_24497);
nor UO_1354 (O_1354,N_23178,N_22774);
nand UO_1355 (O_1355,N_22637,N_23443);
or UO_1356 (O_1356,N_24502,N_22861);
nand UO_1357 (O_1357,N_22539,N_22571);
and UO_1358 (O_1358,N_23275,N_23010);
nand UO_1359 (O_1359,N_23829,N_23217);
nor UO_1360 (O_1360,N_23636,N_23198);
nor UO_1361 (O_1361,N_24348,N_23331);
nor UO_1362 (O_1362,N_23615,N_24591);
nand UO_1363 (O_1363,N_22954,N_23726);
xor UO_1364 (O_1364,N_24863,N_24790);
and UO_1365 (O_1365,N_24983,N_24820);
nand UO_1366 (O_1366,N_23756,N_22653);
or UO_1367 (O_1367,N_23235,N_22942);
or UO_1368 (O_1368,N_23350,N_23039);
nor UO_1369 (O_1369,N_24518,N_24593);
nor UO_1370 (O_1370,N_24667,N_23952);
and UO_1371 (O_1371,N_22839,N_24540);
nand UO_1372 (O_1372,N_23650,N_22727);
nor UO_1373 (O_1373,N_24327,N_23420);
nor UO_1374 (O_1374,N_23977,N_23112);
nor UO_1375 (O_1375,N_22631,N_24200);
nor UO_1376 (O_1376,N_23926,N_24017);
nor UO_1377 (O_1377,N_24626,N_24226);
and UO_1378 (O_1378,N_22814,N_24095);
or UO_1379 (O_1379,N_22988,N_24603);
nand UO_1380 (O_1380,N_23565,N_22741);
nor UO_1381 (O_1381,N_24234,N_24133);
nor UO_1382 (O_1382,N_24550,N_22513);
and UO_1383 (O_1383,N_23494,N_23764);
nand UO_1384 (O_1384,N_24236,N_22997);
nand UO_1385 (O_1385,N_24204,N_24501);
and UO_1386 (O_1386,N_24141,N_24618);
nor UO_1387 (O_1387,N_23607,N_23426);
nand UO_1388 (O_1388,N_24371,N_24108);
or UO_1389 (O_1389,N_24846,N_23924);
or UO_1390 (O_1390,N_23433,N_24985);
and UO_1391 (O_1391,N_22835,N_22575);
xnor UO_1392 (O_1392,N_23624,N_23886);
nand UO_1393 (O_1393,N_22850,N_22713);
or UO_1394 (O_1394,N_24166,N_23779);
nor UO_1395 (O_1395,N_23644,N_24543);
or UO_1396 (O_1396,N_24815,N_23385);
and UO_1397 (O_1397,N_23943,N_23554);
and UO_1398 (O_1398,N_23461,N_23194);
nand UO_1399 (O_1399,N_22860,N_22734);
nand UO_1400 (O_1400,N_23518,N_24608);
nand UO_1401 (O_1401,N_23973,N_24484);
and UO_1402 (O_1402,N_24253,N_22653);
and UO_1403 (O_1403,N_23127,N_24274);
xor UO_1404 (O_1404,N_24553,N_23832);
nand UO_1405 (O_1405,N_24091,N_23398);
or UO_1406 (O_1406,N_23493,N_24121);
or UO_1407 (O_1407,N_23049,N_23497);
and UO_1408 (O_1408,N_23660,N_22814);
nand UO_1409 (O_1409,N_24026,N_24417);
and UO_1410 (O_1410,N_23791,N_23560);
and UO_1411 (O_1411,N_24768,N_24881);
nand UO_1412 (O_1412,N_24774,N_23116);
nand UO_1413 (O_1413,N_24216,N_24297);
and UO_1414 (O_1414,N_24571,N_23959);
or UO_1415 (O_1415,N_23108,N_22820);
nand UO_1416 (O_1416,N_23461,N_23925);
or UO_1417 (O_1417,N_24420,N_23549);
or UO_1418 (O_1418,N_23952,N_22638);
nand UO_1419 (O_1419,N_24879,N_23025);
nand UO_1420 (O_1420,N_23284,N_24534);
nor UO_1421 (O_1421,N_23213,N_24920);
or UO_1422 (O_1422,N_23935,N_24480);
nor UO_1423 (O_1423,N_24350,N_24166);
nor UO_1424 (O_1424,N_22670,N_23522);
or UO_1425 (O_1425,N_23665,N_22659);
nor UO_1426 (O_1426,N_24197,N_23883);
nor UO_1427 (O_1427,N_24637,N_22779);
nand UO_1428 (O_1428,N_24570,N_23440);
xnor UO_1429 (O_1429,N_24346,N_24743);
nor UO_1430 (O_1430,N_22882,N_22737);
nor UO_1431 (O_1431,N_23792,N_24837);
nand UO_1432 (O_1432,N_22584,N_24897);
nand UO_1433 (O_1433,N_23681,N_24932);
or UO_1434 (O_1434,N_24082,N_24923);
nand UO_1435 (O_1435,N_23764,N_24717);
and UO_1436 (O_1436,N_24511,N_24499);
and UO_1437 (O_1437,N_24704,N_24939);
or UO_1438 (O_1438,N_22676,N_22685);
nand UO_1439 (O_1439,N_23863,N_23033);
and UO_1440 (O_1440,N_24438,N_23874);
and UO_1441 (O_1441,N_22723,N_24900);
and UO_1442 (O_1442,N_24048,N_23797);
or UO_1443 (O_1443,N_22937,N_22568);
nor UO_1444 (O_1444,N_22699,N_23660);
and UO_1445 (O_1445,N_23456,N_22754);
and UO_1446 (O_1446,N_22709,N_24177);
nand UO_1447 (O_1447,N_23460,N_22902);
or UO_1448 (O_1448,N_24263,N_23767);
or UO_1449 (O_1449,N_24689,N_23521);
nand UO_1450 (O_1450,N_24695,N_23343);
nor UO_1451 (O_1451,N_24178,N_22648);
nor UO_1452 (O_1452,N_24707,N_22708);
nand UO_1453 (O_1453,N_24821,N_22788);
or UO_1454 (O_1454,N_22504,N_24204);
or UO_1455 (O_1455,N_22580,N_22773);
xnor UO_1456 (O_1456,N_23897,N_24393);
nor UO_1457 (O_1457,N_24867,N_23051);
and UO_1458 (O_1458,N_23436,N_24229);
or UO_1459 (O_1459,N_23154,N_24563);
nor UO_1460 (O_1460,N_22740,N_24102);
nor UO_1461 (O_1461,N_22725,N_23776);
nand UO_1462 (O_1462,N_23218,N_24919);
and UO_1463 (O_1463,N_23853,N_23576);
or UO_1464 (O_1464,N_24357,N_24554);
or UO_1465 (O_1465,N_24120,N_24312);
and UO_1466 (O_1466,N_22928,N_24239);
nor UO_1467 (O_1467,N_24194,N_24191);
or UO_1468 (O_1468,N_24726,N_22872);
nor UO_1469 (O_1469,N_23096,N_22504);
nor UO_1470 (O_1470,N_24998,N_22853);
and UO_1471 (O_1471,N_24907,N_23724);
nand UO_1472 (O_1472,N_24359,N_22802);
or UO_1473 (O_1473,N_23458,N_24155);
and UO_1474 (O_1474,N_24757,N_22559);
nand UO_1475 (O_1475,N_23269,N_24550);
or UO_1476 (O_1476,N_24649,N_24088);
and UO_1477 (O_1477,N_24802,N_23681);
and UO_1478 (O_1478,N_22923,N_23006);
or UO_1479 (O_1479,N_23114,N_23075);
or UO_1480 (O_1480,N_23405,N_24092);
and UO_1481 (O_1481,N_24538,N_24422);
nand UO_1482 (O_1482,N_24771,N_23651);
nor UO_1483 (O_1483,N_23891,N_24282);
nand UO_1484 (O_1484,N_24844,N_22700);
or UO_1485 (O_1485,N_23098,N_24534);
nor UO_1486 (O_1486,N_23897,N_24142);
and UO_1487 (O_1487,N_23697,N_24229);
or UO_1488 (O_1488,N_23163,N_23589);
and UO_1489 (O_1489,N_22812,N_23098);
or UO_1490 (O_1490,N_23219,N_24139);
and UO_1491 (O_1491,N_24422,N_23083);
or UO_1492 (O_1492,N_24563,N_23545);
and UO_1493 (O_1493,N_24722,N_24913);
nand UO_1494 (O_1494,N_23074,N_23259);
and UO_1495 (O_1495,N_24959,N_23121);
or UO_1496 (O_1496,N_24947,N_24965);
nand UO_1497 (O_1497,N_23103,N_23089);
nor UO_1498 (O_1498,N_24582,N_22981);
nor UO_1499 (O_1499,N_22992,N_23634);
nand UO_1500 (O_1500,N_24672,N_24770);
and UO_1501 (O_1501,N_23435,N_22878);
or UO_1502 (O_1502,N_23504,N_23133);
nand UO_1503 (O_1503,N_23704,N_22602);
and UO_1504 (O_1504,N_24260,N_23695);
nor UO_1505 (O_1505,N_24120,N_23420);
nand UO_1506 (O_1506,N_24341,N_23082);
nand UO_1507 (O_1507,N_22731,N_24286);
or UO_1508 (O_1508,N_22809,N_22510);
nand UO_1509 (O_1509,N_24094,N_23351);
nand UO_1510 (O_1510,N_24654,N_24074);
nand UO_1511 (O_1511,N_24257,N_23745);
nand UO_1512 (O_1512,N_22622,N_24685);
nand UO_1513 (O_1513,N_23597,N_23900);
nor UO_1514 (O_1514,N_22818,N_24773);
nor UO_1515 (O_1515,N_23322,N_24360);
and UO_1516 (O_1516,N_23700,N_23423);
and UO_1517 (O_1517,N_23654,N_24156);
or UO_1518 (O_1518,N_22525,N_23823);
or UO_1519 (O_1519,N_22529,N_23231);
nor UO_1520 (O_1520,N_22897,N_22732);
and UO_1521 (O_1521,N_23017,N_24879);
nand UO_1522 (O_1522,N_23403,N_23662);
or UO_1523 (O_1523,N_22827,N_24152);
or UO_1524 (O_1524,N_24650,N_24330);
or UO_1525 (O_1525,N_23834,N_22554);
xnor UO_1526 (O_1526,N_22774,N_23923);
nor UO_1527 (O_1527,N_22810,N_23346);
or UO_1528 (O_1528,N_22882,N_23858);
or UO_1529 (O_1529,N_24774,N_24193);
and UO_1530 (O_1530,N_24246,N_24276);
and UO_1531 (O_1531,N_24058,N_24866);
or UO_1532 (O_1532,N_23339,N_24923);
or UO_1533 (O_1533,N_23193,N_24993);
nor UO_1534 (O_1534,N_22503,N_24179);
nor UO_1535 (O_1535,N_24959,N_23774);
or UO_1536 (O_1536,N_24312,N_24809);
or UO_1537 (O_1537,N_24361,N_24532);
nor UO_1538 (O_1538,N_24778,N_24801);
nor UO_1539 (O_1539,N_23381,N_22818);
nor UO_1540 (O_1540,N_22714,N_23705);
or UO_1541 (O_1541,N_23741,N_23753);
nor UO_1542 (O_1542,N_23627,N_23367);
nor UO_1543 (O_1543,N_23785,N_24113);
and UO_1544 (O_1544,N_23837,N_23909);
xor UO_1545 (O_1545,N_23418,N_23394);
and UO_1546 (O_1546,N_24568,N_24889);
and UO_1547 (O_1547,N_24454,N_22849);
or UO_1548 (O_1548,N_23295,N_24986);
nor UO_1549 (O_1549,N_23987,N_23674);
or UO_1550 (O_1550,N_22727,N_24697);
and UO_1551 (O_1551,N_24681,N_24556);
nand UO_1552 (O_1552,N_23803,N_23985);
or UO_1553 (O_1553,N_24569,N_24228);
and UO_1554 (O_1554,N_24794,N_22917);
or UO_1555 (O_1555,N_24214,N_23772);
or UO_1556 (O_1556,N_23356,N_22762);
or UO_1557 (O_1557,N_23913,N_24217);
or UO_1558 (O_1558,N_23377,N_22797);
or UO_1559 (O_1559,N_23570,N_23160);
nor UO_1560 (O_1560,N_24795,N_22652);
or UO_1561 (O_1561,N_24637,N_23748);
nor UO_1562 (O_1562,N_24725,N_23686);
nor UO_1563 (O_1563,N_23101,N_23264);
and UO_1564 (O_1564,N_24921,N_22983);
nor UO_1565 (O_1565,N_22696,N_24576);
and UO_1566 (O_1566,N_23401,N_24996);
nand UO_1567 (O_1567,N_24370,N_22674);
or UO_1568 (O_1568,N_24289,N_23207);
nor UO_1569 (O_1569,N_24191,N_22643);
and UO_1570 (O_1570,N_24475,N_23270);
and UO_1571 (O_1571,N_22965,N_24841);
nor UO_1572 (O_1572,N_23031,N_24108);
nor UO_1573 (O_1573,N_23650,N_22724);
nand UO_1574 (O_1574,N_23732,N_22875);
or UO_1575 (O_1575,N_23950,N_22879);
nor UO_1576 (O_1576,N_24748,N_24283);
nand UO_1577 (O_1577,N_23930,N_22941);
nor UO_1578 (O_1578,N_24923,N_23303);
nor UO_1579 (O_1579,N_23333,N_24482);
and UO_1580 (O_1580,N_23596,N_23963);
nand UO_1581 (O_1581,N_22538,N_24392);
nor UO_1582 (O_1582,N_23108,N_22773);
or UO_1583 (O_1583,N_23180,N_23767);
nor UO_1584 (O_1584,N_24261,N_23995);
nand UO_1585 (O_1585,N_24332,N_23094);
nand UO_1586 (O_1586,N_24638,N_23806);
and UO_1587 (O_1587,N_23882,N_24159);
nand UO_1588 (O_1588,N_23154,N_23900);
nand UO_1589 (O_1589,N_23572,N_23488);
and UO_1590 (O_1590,N_24506,N_23769);
or UO_1591 (O_1591,N_23860,N_24852);
nand UO_1592 (O_1592,N_24313,N_24162);
or UO_1593 (O_1593,N_24076,N_23456);
or UO_1594 (O_1594,N_23003,N_23398);
or UO_1595 (O_1595,N_22660,N_24237);
nor UO_1596 (O_1596,N_22588,N_22966);
nor UO_1597 (O_1597,N_24361,N_23469);
nor UO_1598 (O_1598,N_22643,N_24674);
nand UO_1599 (O_1599,N_22835,N_24039);
nor UO_1600 (O_1600,N_22976,N_23951);
nor UO_1601 (O_1601,N_22763,N_24683);
nor UO_1602 (O_1602,N_23907,N_23904);
and UO_1603 (O_1603,N_24263,N_22679);
and UO_1604 (O_1604,N_24316,N_24177);
nand UO_1605 (O_1605,N_23149,N_24794);
or UO_1606 (O_1606,N_23702,N_24227);
xor UO_1607 (O_1607,N_23970,N_24789);
nand UO_1608 (O_1608,N_22503,N_23679);
nor UO_1609 (O_1609,N_23063,N_24361);
or UO_1610 (O_1610,N_24288,N_24352);
nand UO_1611 (O_1611,N_23159,N_24890);
nor UO_1612 (O_1612,N_24033,N_23050);
nand UO_1613 (O_1613,N_23261,N_24038);
and UO_1614 (O_1614,N_24123,N_23244);
or UO_1615 (O_1615,N_24040,N_24396);
and UO_1616 (O_1616,N_23251,N_24007);
nand UO_1617 (O_1617,N_24464,N_24850);
or UO_1618 (O_1618,N_24483,N_23851);
and UO_1619 (O_1619,N_22680,N_24205);
and UO_1620 (O_1620,N_22728,N_24907);
or UO_1621 (O_1621,N_23220,N_23169);
and UO_1622 (O_1622,N_24037,N_23863);
and UO_1623 (O_1623,N_22824,N_23284);
or UO_1624 (O_1624,N_24752,N_24251);
nand UO_1625 (O_1625,N_23868,N_23837);
nand UO_1626 (O_1626,N_24546,N_24587);
and UO_1627 (O_1627,N_22890,N_24380);
or UO_1628 (O_1628,N_22893,N_23650);
and UO_1629 (O_1629,N_23987,N_22586);
nor UO_1630 (O_1630,N_22540,N_23812);
xor UO_1631 (O_1631,N_23832,N_24959);
nor UO_1632 (O_1632,N_24627,N_24734);
nor UO_1633 (O_1633,N_24147,N_22689);
and UO_1634 (O_1634,N_22981,N_23841);
or UO_1635 (O_1635,N_22618,N_24990);
nor UO_1636 (O_1636,N_23573,N_24671);
and UO_1637 (O_1637,N_22761,N_23483);
or UO_1638 (O_1638,N_24369,N_24746);
nor UO_1639 (O_1639,N_24798,N_24234);
xor UO_1640 (O_1640,N_24097,N_23496);
xnor UO_1641 (O_1641,N_23280,N_24355);
nand UO_1642 (O_1642,N_23723,N_22731);
nand UO_1643 (O_1643,N_24805,N_23364);
or UO_1644 (O_1644,N_23921,N_23900);
nand UO_1645 (O_1645,N_23218,N_24525);
xnor UO_1646 (O_1646,N_23785,N_22799);
nand UO_1647 (O_1647,N_24547,N_23868);
or UO_1648 (O_1648,N_22636,N_22521);
nor UO_1649 (O_1649,N_22790,N_23268);
xnor UO_1650 (O_1650,N_24507,N_23374);
nand UO_1651 (O_1651,N_23278,N_23119);
or UO_1652 (O_1652,N_22881,N_23461);
nor UO_1653 (O_1653,N_23511,N_22908);
and UO_1654 (O_1654,N_24678,N_23037);
and UO_1655 (O_1655,N_23495,N_24408);
and UO_1656 (O_1656,N_24046,N_24313);
and UO_1657 (O_1657,N_22905,N_23669);
nand UO_1658 (O_1658,N_23823,N_22718);
or UO_1659 (O_1659,N_24986,N_23537);
or UO_1660 (O_1660,N_24063,N_24148);
nand UO_1661 (O_1661,N_23309,N_23622);
nor UO_1662 (O_1662,N_23586,N_23852);
and UO_1663 (O_1663,N_24989,N_23280);
nor UO_1664 (O_1664,N_23845,N_24562);
nand UO_1665 (O_1665,N_24551,N_23850);
nand UO_1666 (O_1666,N_22801,N_24939);
nand UO_1667 (O_1667,N_24875,N_24428);
and UO_1668 (O_1668,N_24450,N_23869);
nand UO_1669 (O_1669,N_23607,N_24918);
and UO_1670 (O_1670,N_22995,N_23043);
or UO_1671 (O_1671,N_24922,N_24312);
or UO_1672 (O_1672,N_24678,N_22666);
nand UO_1673 (O_1673,N_24506,N_23374);
and UO_1674 (O_1674,N_23444,N_22701);
nor UO_1675 (O_1675,N_24254,N_24077);
nor UO_1676 (O_1676,N_24033,N_24091);
or UO_1677 (O_1677,N_23338,N_23145);
and UO_1678 (O_1678,N_24149,N_23155);
nand UO_1679 (O_1679,N_24028,N_23278);
nand UO_1680 (O_1680,N_23223,N_24984);
or UO_1681 (O_1681,N_24727,N_23815);
or UO_1682 (O_1682,N_23225,N_22889);
nor UO_1683 (O_1683,N_23149,N_24382);
nor UO_1684 (O_1684,N_24878,N_23189);
or UO_1685 (O_1685,N_24040,N_24259);
nand UO_1686 (O_1686,N_22558,N_24730);
and UO_1687 (O_1687,N_24983,N_23147);
and UO_1688 (O_1688,N_24479,N_24189);
nor UO_1689 (O_1689,N_24793,N_23143);
nor UO_1690 (O_1690,N_24941,N_22851);
and UO_1691 (O_1691,N_24380,N_22715);
nand UO_1692 (O_1692,N_24773,N_23853);
or UO_1693 (O_1693,N_24037,N_22561);
and UO_1694 (O_1694,N_23479,N_23996);
and UO_1695 (O_1695,N_24697,N_22514);
and UO_1696 (O_1696,N_24402,N_22918);
nor UO_1697 (O_1697,N_22737,N_23318);
nand UO_1698 (O_1698,N_23590,N_23159);
or UO_1699 (O_1699,N_22673,N_24397);
nor UO_1700 (O_1700,N_23779,N_22627);
nand UO_1701 (O_1701,N_24364,N_22505);
and UO_1702 (O_1702,N_22815,N_22570);
or UO_1703 (O_1703,N_23035,N_24761);
or UO_1704 (O_1704,N_23706,N_24932);
or UO_1705 (O_1705,N_22608,N_23270);
or UO_1706 (O_1706,N_23524,N_23724);
xor UO_1707 (O_1707,N_24903,N_24539);
nand UO_1708 (O_1708,N_22690,N_23259);
nor UO_1709 (O_1709,N_24646,N_23221);
xor UO_1710 (O_1710,N_22742,N_24187);
or UO_1711 (O_1711,N_24483,N_23234);
nor UO_1712 (O_1712,N_22988,N_24462);
nor UO_1713 (O_1713,N_23184,N_23892);
and UO_1714 (O_1714,N_22553,N_24855);
or UO_1715 (O_1715,N_23148,N_23869);
xor UO_1716 (O_1716,N_24355,N_23325);
nand UO_1717 (O_1717,N_23516,N_22955);
nand UO_1718 (O_1718,N_24576,N_22918);
and UO_1719 (O_1719,N_22668,N_24060);
and UO_1720 (O_1720,N_24939,N_24440);
and UO_1721 (O_1721,N_23989,N_22900);
and UO_1722 (O_1722,N_24639,N_23123);
or UO_1723 (O_1723,N_23607,N_23353);
or UO_1724 (O_1724,N_23177,N_24920);
nand UO_1725 (O_1725,N_24164,N_22921);
and UO_1726 (O_1726,N_24430,N_23764);
or UO_1727 (O_1727,N_24069,N_23665);
xnor UO_1728 (O_1728,N_24124,N_22629);
or UO_1729 (O_1729,N_24409,N_23766);
and UO_1730 (O_1730,N_24301,N_23401);
or UO_1731 (O_1731,N_24993,N_24889);
nor UO_1732 (O_1732,N_22697,N_22869);
xor UO_1733 (O_1733,N_24495,N_23163);
nand UO_1734 (O_1734,N_23291,N_22854);
or UO_1735 (O_1735,N_23840,N_23990);
nand UO_1736 (O_1736,N_23036,N_23438);
nor UO_1737 (O_1737,N_24982,N_23226);
nand UO_1738 (O_1738,N_23447,N_24399);
or UO_1739 (O_1739,N_24121,N_24053);
or UO_1740 (O_1740,N_22914,N_24079);
xor UO_1741 (O_1741,N_24748,N_22995);
or UO_1742 (O_1742,N_24672,N_22853);
nand UO_1743 (O_1743,N_24298,N_23896);
or UO_1744 (O_1744,N_23861,N_23148);
or UO_1745 (O_1745,N_23483,N_24016);
nand UO_1746 (O_1746,N_23122,N_22598);
and UO_1747 (O_1747,N_24136,N_22620);
or UO_1748 (O_1748,N_24394,N_24396);
and UO_1749 (O_1749,N_23298,N_23882);
and UO_1750 (O_1750,N_23363,N_24231);
and UO_1751 (O_1751,N_24487,N_22760);
nor UO_1752 (O_1752,N_23868,N_24666);
and UO_1753 (O_1753,N_24866,N_23624);
and UO_1754 (O_1754,N_23238,N_24055);
nand UO_1755 (O_1755,N_23600,N_22971);
or UO_1756 (O_1756,N_24960,N_24912);
and UO_1757 (O_1757,N_24034,N_24410);
or UO_1758 (O_1758,N_23205,N_23244);
or UO_1759 (O_1759,N_24992,N_23748);
nand UO_1760 (O_1760,N_24833,N_22703);
nor UO_1761 (O_1761,N_23371,N_23455);
nand UO_1762 (O_1762,N_22747,N_23600);
nor UO_1763 (O_1763,N_23311,N_24845);
nor UO_1764 (O_1764,N_22964,N_23877);
and UO_1765 (O_1765,N_22961,N_23443);
xor UO_1766 (O_1766,N_22814,N_24435);
and UO_1767 (O_1767,N_22855,N_23625);
nor UO_1768 (O_1768,N_23319,N_22511);
or UO_1769 (O_1769,N_24239,N_22516);
nor UO_1770 (O_1770,N_23859,N_22501);
xor UO_1771 (O_1771,N_23077,N_23313);
or UO_1772 (O_1772,N_22658,N_24340);
nor UO_1773 (O_1773,N_22809,N_23696);
nor UO_1774 (O_1774,N_24739,N_23314);
or UO_1775 (O_1775,N_22975,N_22728);
or UO_1776 (O_1776,N_24077,N_24784);
nand UO_1777 (O_1777,N_22875,N_23779);
xor UO_1778 (O_1778,N_23331,N_22739);
nand UO_1779 (O_1779,N_22953,N_23657);
nand UO_1780 (O_1780,N_24962,N_24975);
nand UO_1781 (O_1781,N_22770,N_23259);
nor UO_1782 (O_1782,N_22651,N_23046);
nand UO_1783 (O_1783,N_23991,N_24522);
nor UO_1784 (O_1784,N_24865,N_22990);
or UO_1785 (O_1785,N_24906,N_23628);
or UO_1786 (O_1786,N_24855,N_23154);
nor UO_1787 (O_1787,N_24521,N_24483);
nand UO_1788 (O_1788,N_23722,N_24746);
or UO_1789 (O_1789,N_24507,N_24870);
and UO_1790 (O_1790,N_24902,N_24453);
nand UO_1791 (O_1791,N_24793,N_23151);
and UO_1792 (O_1792,N_23065,N_23836);
and UO_1793 (O_1793,N_23824,N_24267);
nand UO_1794 (O_1794,N_24879,N_22625);
and UO_1795 (O_1795,N_24356,N_23987);
nand UO_1796 (O_1796,N_24728,N_24403);
nand UO_1797 (O_1797,N_22858,N_23665);
nand UO_1798 (O_1798,N_22856,N_24146);
nor UO_1799 (O_1799,N_24769,N_23744);
and UO_1800 (O_1800,N_23110,N_23571);
or UO_1801 (O_1801,N_24603,N_22637);
nor UO_1802 (O_1802,N_23388,N_22543);
nor UO_1803 (O_1803,N_23161,N_22635);
nand UO_1804 (O_1804,N_23313,N_22711);
or UO_1805 (O_1805,N_23705,N_23400);
nor UO_1806 (O_1806,N_22760,N_23351);
and UO_1807 (O_1807,N_23660,N_24527);
nand UO_1808 (O_1808,N_24630,N_22701);
and UO_1809 (O_1809,N_22706,N_22932);
and UO_1810 (O_1810,N_24517,N_23631);
and UO_1811 (O_1811,N_24468,N_23821);
nor UO_1812 (O_1812,N_22734,N_24745);
nor UO_1813 (O_1813,N_23419,N_24723);
nand UO_1814 (O_1814,N_23391,N_23594);
or UO_1815 (O_1815,N_22585,N_22941);
or UO_1816 (O_1816,N_23745,N_23343);
or UO_1817 (O_1817,N_23182,N_23086);
or UO_1818 (O_1818,N_24729,N_23752);
nor UO_1819 (O_1819,N_24661,N_23009);
and UO_1820 (O_1820,N_24356,N_23587);
and UO_1821 (O_1821,N_23378,N_24546);
and UO_1822 (O_1822,N_24005,N_23922);
and UO_1823 (O_1823,N_24521,N_24759);
and UO_1824 (O_1824,N_23982,N_23378);
xnor UO_1825 (O_1825,N_22903,N_24370);
xor UO_1826 (O_1826,N_23499,N_23349);
nand UO_1827 (O_1827,N_23416,N_23866);
and UO_1828 (O_1828,N_24676,N_22591);
or UO_1829 (O_1829,N_23503,N_23054);
and UO_1830 (O_1830,N_22863,N_24458);
nor UO_1831 (O_1831,N_22900,N_22545);
nor UO_1832 (O_1832,N_23378,N_22532);
and UO_1833 (O_1833,N_24351,N_22978);
nor UO_1834 (O_1834,N_23205,N_23050);
nor UO_1835 (O_1835,N_23240,N_23074);
or UO_1836 (O_1836,N_24061,N_22563);
or UO_1837 (O_1837,N_22606,N_23408);
nand UO_1838 (O_1838,N_23991,N_24577);
nand UO_1839 (O_1839,N_24160,N_24147);
nor UO_1840 (O_1840,N_24194,N_22542);
nand UO_1841 (O_1841,N_23766,N_24931);
and UO_1842 (O_1842,N_22915,N_22661);
and UO_1843 (O_1843,N_24470,N_23305);
nor UO_1844 (O_1844,N_23008,N_23171);
nand UO_1845 (O_1845,N_24782,N_23251);
nand UO_1846 (O_1846,N_24163,N_22602);
or UO_1847 (O_1847,N_23737,N_24084);
nor UO_1848 (O_1848,N_23842,N_24856);
xor UO_1849 (O_1849,N_23102,N_24473);
nor UO_1850 (O_1850,N_23856,N_23577);
and UO_1851 (O_1851,N_23428,N_22582);
nor UO_1852 (O_1852,N_24644,N_24492);
xnor UO_1853 (O_1853,N_24260,N_24715);
nor UO_1854 (O_1854,N_24881,N_23114);
nor UO_1855 (O_1855,N_23851,N_24017);
or UO_1856 (O_1856,N_23488,N_23061);
nand UO_1857 (O_1857,N_22944,N_22837);
and UO_1858 (O_1858,N_24748,N_23960);
nor UO_1859 (O_1859,N_22761,N_23410);
and UO_1860 (O_1860,N_24712,N_22697);
nor UO_1861 (O_1861,N_24306,N_22944);
nand UO_1862 (O_1862,N_22553,N_22526);
or UO_1863 (O_1863,N_24073,N_24253);
nor UO_1864 (O_1864,N_22509,N_24377);
nand UO_1865 (O_1865,N_22518,N_23285);
nand UO_1866 (O_1866,N_23197,N_22920);
and UO_1867 (O_1867,N_23364,N_24660);
or UO_1868 (O_1868,N_22802,N_24740);
nor UO_1869 (O_1869,N_23865,N_23823);
and UO_1870 (O_1870,N_22991,N_23365);
nand UO_1871 (O_1871,N_24980,N_23247);
and UO_1872 (O_1872,N_23986,N_24707);
and UO_1873 (O_1873,N_24816,N_23701);
and UO_1874 (O_1874,N_23953,N_24133);
and UO_1875 (O_1875,N_23397,N_23114);
nor UO_1876 (O_1876,N_23348,N_24623);
nand UO_1877 (O_1877,N_24097,N_23170);
or UO_1878 (O_1878,N_22557,N_22793);
nor UO_1879 (O_1879,N_24832,N_22966);
nor UO_1880 (O_1880,N_23349,N_22987);
nand UO_1881 (O_1881,N_24256,N_23561);
and UO_1882 (O_1882,N_24341,N_24904);
or UO_1883 (O_1883,N_22860,N_23663);
nand UO_1884 (O_1884,N_24670,N_23507);
nand UO_1885 (O_1885,N_24484,N_22689);
nor UO_1886 (O_1886,N_22754,N_23904);
or UO_1887 (O_1887,N_22965,N_23722);
or UO_1888 (O_1888,N_24219,N_22538);
or UO_1889 (O_1889,N_24213,N_24863);
or UO_1890 (O_1890,N_24785,N_22615);
and UO_1891 (O_1891,N_24610,N_23522);
nor UO_1892 (O_1892,N_24042,N_23123);
nand UO_1893 (O_1893,N_22658,N_22798);
or UO_1894 (O_1894,N_23533,N_23320);
nor UO_1895 (O_1895,N_23560,N_24618);
or UO_1896 (O_1896,N_23734,N_22638);
xor UO_1897 (O_1897,N_23342,N_24227);
and UO_1898 (O_1898,N_23103,N_22837);
or UO_1899 (O_1899,N_23658,N_24297);
nor UO_1900 (O_1900,N_23278,N_24759);
nor UO_1901 (O_1901,N_22907,N_24161);
nor UO_1902 (O_1902,N_23203,N_23360);
and UO_1903 (O_1903,N_22751,N_23508);
nand UO_1904 (O_1904,N_24284,N_24306);
or UO_1905 (O_1905,N_23604,N_23617);
or UO_1906 (O_1906,N_22648,N_24188);
nand UO_1907 (O_1907,N_23846,N_24410);
xnor UO_1908 (O_1908,N_24776,N_23071);
xor UO_1909 (O_1909,N_23881,N_23902);
nor UO_1910 (O_1910,N_22595,N_24840);
or UO_1911 (O_1911,N_24282,N_23215);
nand UO_1912 (O_1912,N_23878,N_23768);
or UO_1913 (O_1913,N_24569,N_23781);
and UO_1914 (O_1914,N_23966,N_22722);
and UO_1915 (O_1915,N_23677,N_23162);
or UO_1916 (O_1916,N_23893,N_24202);
and UO_1917 (O_1917,N_23544,N_24526);
or UO_1918 (O_1918,N_24938,N_23443);
or UO_1919 (O_1919,N_24463,N_23178);
or UO_1920 (O_1920,N_23394,N_23763);
or UO_1921 (O_1921,N_24258,N_23376);
nor UO_1922 (O_1922,N_24251,N_24294);
and UO_1923 (O_1923,N_23885,N_22815);
nor UO_1924 (O_1924,N_24971,N_22701);
xor UO_1925 (O_1925,N_24626,N_24135);
and UO_1926 (O_1926,N_23344,N_23419);
nand UO_1927 (O_1927,N_22995,N_22604);
nand UO_1928 (O_1928,N_23306,N_23190);
nand UO_1929 (O_1929,N_23544,N_24916);
or UO_1930 (O_1930,N_23111,N_24493);
nand UO_1931 (O_1931,N_23929,N_24179);
xor UO_1932 (O_1932,N_23455,N_24323);
nor UO_1933 (O_1933,N_23348,N_24357);
and UO_1934 (O_1934,N_23512,N_23389);
nor UO_1935 (O_1935,N_23426,N_24136);
nand UO_1936 (O_1936,N_24322,N_23062);
xnor UO_1937 (O_1937,N_24568,N_23539);
and UO_1938 (O_1938,N_24120,N_23460);
and UO_1939 (O_1939,N_24796,N_24931);
or UO_1940 (O_1940,N_23928,N_22568);
nor UO_1941 (O_1941,N_23408,N_24432);
xor UO_1942 (O_1942,N_22536,N_23154);
or UO_1943 (O_1943,N_23498,N_24005);
nor UO_1944 (O_1944,N_22546,N_24156);
nand UO_1945 (O_1945,N_23996,N_24872);
nand UO_1946 (O_1946,N_23833,N_23145);
or UO_1947 (O_1947,N_23718,N_22880);
or UO_1948 (O_1948,N_24334,N_24750);
and UO_1949 (O_1949,N_22565,N_23115);
nand UO_1950 (O_1950,N_23580,N_24362);
nand UO_1951 (O_1951,N_24431,N_24029);
nand UO_1952 (O_1952,N_22837,N_22930);
nor UO_1953 (O_1953,N_24384,N_23239);
and UO_1954 (O_1954,N_24310,N_24598);
xnor UO_1955 (O_1955,N_24451,N_23729);
nand UO_1956 (O_1956,N_24928,N_23382);
or UO_1957 (O_1957,N_22785,N_23531);
nand UO_1958 (O_1958,N_24153,N_23178);
or UO_1959 (O_1959,N_23043,N_24130);
nand UO_1960 (O_1960,N_24431,N_24957);
nor UO_1961 (O_1961,N_22953,N_23384);
nand UO_1962 (O_1962,N_24670,N_22800);
nor UO_1963 (O_1963,N_22924,N_24671);
and UO_1964 (O_1964,N_22616,N_23064);
and UO_1965 (O_1965,N_24409,N_23541);
nand UO_1966 (O_1966,N_22662,N_24653);
and UO_1967 (O_1967,N_23177,N_24419);
nor UO_1968 (O_1968,N_23918,N_23308);
or UO_1969 (O_1969,N_22659,N_22676);
and UO_1970 (O_1970,N_24132,N_23517);
or UO_1971 (O_1971,N_24062,N_24803);
xor UO_1972 (O_1972,N_24519,N_24976);
nor UO_1973 (O_1973,N_23677,N_24662);
nor UO_1974 (O_1974,N_24911,N_24927);
nand UO_1975 (O_1975,N_22952,N_23789);
nand UO_1976 (O_1976,N_23960,N_22849);
or UO_1977 (O_1977,N_24059,N_23816);
nand UO_1978 (O_1978,N_22640,N_23237);
nand UO_1979 (O_1979,N_24241,N_24298);
or UO_1980 (O_1980,N_24985,N_24794);
and UO_1981 (O_1981,N_24359,N_24174);
nand UO_1982 (O_1982,N_23935,N_23552);
or UO_1983 (O_1983,N_24089,N_22879);
nand UO_1984 (O_1984,N_23739,N_23603);
or UO_1985 (O_1985,N_24093,N_23280);
nor UO_1986 (O_1986,N_24988,N_24940);
and UO_1987 (O_1987,N_23346,N_24325);
nand UO_1988 (O_1988,N_23659,N_23809);
nor UO_1989 (O_1989,N_23493,N_22892);
nor UO_1990 (O_1990,N_23208,N_24263);
nand UO_1991 (O_1991,N_24913,N_24773);
or UO_1992 (O_1992,N_24857,N_23317);
nor UO_1993 (O_1993,N_22558,N_23201);
xor UO_1994 (O_1994,N_24126,N_24862);
nand UO_1995 (O_1995,N_23280,N_23208);
nand UO_1996 (O_1996,N_22972,N_23294);
and UO_1997 (O_1997,N_22964,N_22712);
or UO_1998 (O_1998,N_24017,N_23128);
nor UO_1999 (O_1999,N_22961,N_24547);
or UO_2000 (O_2000,N_22828,N_23332);
nand UO_2001 (O_2001,N_22771,N_24340);
nor UO_2002 (O_2002,N_22769,N_24702);
nor UO_2003 (O_2003,N_23337,N_23483);
or UO_2004 (O_2004,N_23674,N_22741);
and UO_2005 (O_2005,N_24286,N_23609);
or UO_2006 (O_2006,N_22835,N_24844);
nor UO_2007 (O_2007,N_24399,N_23183);
or UO_2008 (O_2008,N_22753,N_24027);
nand UO_2009 (O_2009,N_23727,N_22532);
and UO_2010 (O_2010,N_24326,N_24533);
or UO_2011 (O_2011,N_23351,N_22933);
or UO_2012 (O_2012,N_22673,N_24871);
nor UO_2013 (O_2013,N_24243,N_23624);
nor UO_2014 (O_2014,N_22892,N_23136);
or UO_2015 (O_2015,N_23260,N_24661);
nor UO_2016 (O_2016,N_23662,N_24131);
nand UO_2017 (O_2017,N_24222,N_22533);
nand UO_2018 (O_2018,N_24741,N_24122);
and UO_2019 (O_2019,N_22603,N_22763);
and UO_2020 (O_2020,N_24934,N_23588);
or UO_2021 (O_2021,N_23367,N_24777);
xnor UO_2022 (O_2022,N_23384,N_22675);
nor UO_2023 (O_2023,N_23820,N_23387);
nand UO_2024 (O_2024,N_24501,N_23004);
nor UO_2025 (O_2025,N_24604,N_23572);
nand UO_2026 (O_2026,N_24902,N_23169);
nor UO_2027 (O_2027,N_24109,N_22976);
nand UO_2028 (O_2028,N_22805,N_23262);
nor UO_2029 (O_2029,N_23833,N_24775);
nand UO_2030 (O_2030,N_23211,N_23732);
nor UO_2031 (O_2031,N_23022,N_23775);
or UO_2032 (O_2032,N_23187,N_22530);
nor UO_2033 (O_2033,N_24333,N_24209);
nand UO_2034 (O_2034,N_24467,N_23182);
nand UO_2035 (O_2035,N_22523,N_24993);
xor UO_2036 (O_2036,N_23415,N_23054);
or UO_2037 (O_2037,N_23568,N_24402);
nor UO_2038 (O_2038,N_23779,N_24998);
or UO_2039 (O_2039,N_22553,N_23321);
nand UO_2040 (O_2040,N_23674,N_24453);
or UO_2041 (O_2041,N_24882,N_22518);
and UO_2042 (O_2042,N_23169,N_24724);
nor UO_2043 (O_2043,N_24138,N_24491);
or UO_2044 (O_2044,N_24035,N_24299);
or UO_2045 (O_2045,N_23289,N_24980);
and UO_2046 (O_2046,N_22557,N_23067);
or UO_2047 (O_2047,N_24393,N_22621);
nand UO_2048 (O_2048,N_22756,N_24579);
and UO_2049 (O_2049,N_24310,N_23880);
nor UO_2050 (O_2050,N_24089,N_24847);
or UO_2051 (O_2051,N_24860,N_22855);
nor UO_2052 (O_2052,N_24879,N_24066);
and UO_2053 (O_2053,N_24566,N_23338);
nand UO_2054 (O_2054,N_23097,N_22626);
or UO_2055 (O_2055,N_23593,N_24074);
or UO_2056 (O_2056,N_23342,N_23468);
nand UO_2057 (O_2057,N_23189,N_23760);
and UO_2058 (O_2058,N_24990,N_23564);
and UO_2059 (O_2059,N_23775,N_23163);
nand UO_2060 (O_2060,N_23161,N_23287);
nand UO_2061 (O_2061,N_23858,N_23635);
and UO_2062 (O_2062,N_23323,N_23340);
xnor UO_2063 (O_2063,N_24257,N_23199);
nand UO_2064 (O_2064,N_24430,N_23974);
nor UO_2065 (O_2065,N_24965,N_24287);
nor UO_2066 (O_2066,N_23585,N_23684);
nor UO_2067 (O_2067,N_23634,N_23739);
nor UO_2068 (O_2068,N_22687,N_24753);
or UO_2069 (O_2069,N_24435,N_24682);
nand UO_2070 (O_2070,N_23232,N_24365);
and UO_2071 (O_2071,N_24257,N_23728);
nor UO_2072 (O_2072,N_23218,N_24748);
nor UO_2073 (O_2073,N_24863,N_22533);
nand UO_2074 (O_2074,N_24023,N_24827);
nor UO_2075 (O_2075,N_23240,N_24805);
or UO_2076 (O_2076,N_22687,N_23251);
or UO_2077 (O_2077,N_23490,N_24129);
and UO_2078 (O_2078,N_23059,N_24814);
nor UO_2079 (O_2079,N_23780,N_24459);
nor UO_2080 (O_2080,N_24269,N_23303);
or UO_2081 (O_2081,N_24742,N_24061);
nand UO_2082 (O_2082,N_23187,N_24304);
and UO_2083 (O_2083,N_23338,N_22618);
nand UO_2084 (O_2084,N_23063,N_24056);
nor UO_2085 (O_2085,N_24963,N_22547);
nand UO_2086 (O_2086,N_22832,N_23722);
nor UO_2087 (O_2087,N_23526,N_23236);
nor UO_2088 (O_2088,N_22786,N_23318);
nand UO_2089 (O_2089,N_24282,N_22872);
nand UO_2090 (O_2090,N_24057,N_24859);
nand UO_2091 (O_2091,N_24373,N_22635);
and UO_2092 (O_2092,N_23456,N_23292);
nor UO_2093 (O_2093,N_22869,N_24679);
or UO_2094 (O_2094,N_24962,N_22582);
nor UO_2095 (O_2095,N_23679,N_23122);
nor UO_2096 (O_2096,N_23011,N_23979);
nand UO_2097 (O_2097,N_23996,N_22739);
and UO_2098 (O_2098,N_24263,N_22831);
nand UO_2099 (O_2099,N_24676,N_23509);
or UO_2100 (O_2100,N_23168,N_24815);
nand UO_2101 (O_2101,N_23897,N_24056);
nand UO_2102 (O_2102,N_22778,N_23033);
nor UO_2103 (O_2103,N_23867,N_24013);
and UO_2104 (O_2104,N_24504,N_23576);
nand UO_2105 (O_2105,N_23541,N_23971);
nor UO_2106 (O_2106,N_22652,N_23883);
nand UO_2107 (O_2107,N_23477,N_24823);
nand UO_2108 (O_2108,N_24417,N_22754);
or UO_2109 (O_2109,N_24313,N_23539);
or UO_2110 (O_2110,N_24498,N_24135);
nand UO_2111 (O_2111,N_24959,N_22553);
nand UO_2112 (O_2112,N_24980,N_23610);
nand UO_2113 (O_2113,N_23161,N_23926);
or UO_2114 (O_2114,N_23997,N_23141);
or UO_2115 (O_2115,N_24025,N_22891);
nor UO_2116 (O_2116,N_24146,N_24579);
nand UO_2117 (O_2117,N_23159,N_23922);
and UO_2118 (O_2118,N_24971,N_23872);
nand UO_2119 (O_2119,N_24202,N_24939);
and UO_2120 (O_2120,N_23911,N_24627);
nor UO_2121 (O_2121,N_24838,N_23210);
nand UO_2122 (O_2122,N_22854,N_24160);
or UO_2123 (O_2123,N_24501,N_24919);
nand UO_2124 (O_2124,N_23623,N_24801);
nand UO_2125 (O_2125,N_23292,N_23076);
nand UO_2126 (O_2126,N_23425,N_23258);
nor UO_2127 (O_2127,N_24281,N_24553);
or UO_2128 (O_2128,N_24133,N_24761);
nand UO_2129 (O_2129,N_23970,N_24661);
nor UO_2130 (O_2130,N_22599,N_23640);
or UO_2131 (O_2131,N_23555,N_24700);
and UO_2132 (O_2132,N_24619,N_24221);
xnor UO_2133 (O_2133,N_22720,N_23026);
nor UO_2134 (O_2134,N_24530,N_22869);
and UO_2135 (O_2135,N_23054,N_24882);
or UO_2136 (O_2136,N_22624,N_24310);
or UO_2137 (O_2137,N_24843,N_24838);
or UO_2138 (O_2138,N_23105,N_22699);
xnor UO_2139 (O_2139,N_23140,N_23375);
or UO_2140 (O_2140,N_24295,N_24980);
or UO_2141 (O_2141,N_24251,N_23521);
or UO_2142 (O_2142,N_24495,N_23939);
or UO_2143 (O_2143,N_23233,N_23960);
and UO_2144 (O_2144,N_22903,N_24033);
or UO_2145 (O_2145,N_24183,N_22701);
nand UO_2146 (O_2146,N_23635,N_24924);
nand UO_2147 (O_2147,N_24454,N_23155);
or UO_2148 (O_2148,N_23664,N_22670);
and UO_2149 (O_2149,N_24380,N_24215);
or UO_2150 (O_2150,N_23406,N_24979);
and UO_2151 (O_2151,N_22731,N_22522);
nor UO_2152 (O_2152,N_23720,N_24218);
nor UO_2153 (O_2153,N_24011,N_24964);
nor UO_2154 (O_2154,N_24611,N_23208);
or UO_2155 (O_2155,N_23108,N_23807);
nand UO_2156 (O_2156,N_23357,N_24354);
or UO_2157 (O_2157,N_23750,N_22606);
nor UO_2158 (O_2158,N_23138,N_23944);
or UO_2159 (O_2159,N_24167,N_23770);
nor UO_2160 (O_2160,N_23380,N_22652);
or UO_2161 (O_2161,N_24582,N_23522);
nand UO_2162 (O_2162,N_23291,N_24599);
and UO_2163 (O_2163,N_24218,N_24406);
and UO_2164 (O_2164,N_23473,N_22595);
nor UO_2165 (O_2165,N_24433,N_23249);
nand UO_2166 (O_2166,N_22536,N_24958);
or UO_2167 (O_2167,N_24362,N_23277);
nand UO_2168 (O_2168,N_22543,N_24628);
nor UO_2169 (O_2169,N_23311,N_22622);
or UO_2170 (O_2170,N_24327,N_23437);
and UO_2171 (O_2171,N_24162,N_22587);
and UO_2172 (O_2172,N_24908,N_22806);
nand UO_2173 (O_2173,N_23183,N_23195);
or UO_2174 (O_2174,N_24212,N_24321);
nor UO_2175 (O_2175,N_22665,N_24091);
and UO_2176 (O_2176,N_24948,N_23759);
nor UO_2177 (O_2177,N_23989,N_24079);
and UO_2178 (O_2178,N_24934,N_23149);
nor UO_2179 (O_2179,N_24993,N_24554);
or UO_2180 (O_2180,N_22908,N_23703);
or UO_2181 (O_2181,N_23450,N_24441);
nor UO_2182 (O_2182,N_23264,N_24261);
or UO_2183 (O_2183,N_23585,N_22632);
and UO_2184 (O_2184,N_24241,N_24685);
and UO_2185 (O_2185,N_24905,N_24319);
nand UO_2186 (O_2186,N_22624,N_24290);
or UO_2187 (O_2187,N_24493,N_24551);
or UO_2188 (O_2188,N_24310,N_22705);
nor UO_2189 (O_2189,N_23338,N_23387);
nor UO_2190 (O_2190,N_24337,N_23503);
or UO_2191 (O_2191,N_23308,N_22998);
nand UO_2192 (O_2192,N_23425,N_23237);
nand UO_2193 (O_2193,N_24485,N_23380);
nor UO_2194 (O_2194,N_22792,N_23657);
nor UO_2195 (O_2195,N_24495,N_24518);
nand UO_2196 (O_2196,N_23392,N_24318);
nor UO_2197 (O_2197,N_23728,N_23408);
nor UO_2198 (O_2198,N_24187,N_22733);
or UO_2199 (O_2199,N_22760,N_24869);
and UO_2200 (O_2200,N_23643,N_24581);
nor UO_2201 (O_2201,N_23146,N_24243);
xnor UO_2202 (O_2202,N_24773,N_23968);
nor UO_2203 (O_2203,N_23781,N_23060);
nor UO_2204 (O_2204,N_24997,N_22911);
or UO_2205 (O_2205,N_24395,N_23543);
nor UO_2206 (O_2206,N_23554,N_23340);
or UO_2207 (O_2207,N_22908,N_23824);
and UO_2208 (O_2208,N_23018,N_24038);
nor UO_2209 (O_2209,N_22857,N_23472);
nor UO_2210 (O_2210,N_24935,N_24216);
or UO_2211 (O_2211,N_24710,N_23084);
and UO_2212 (O_2212,N_23580,N_23340);
nor UO_2213 (O_2213,N_24113,N_22789);
and UO_2214 (O_2214,N_23786,N_24672);
nor UO_2215 (O_2215,N_23289,N_24689);
nand UO_2216 (O_2216,N_23936,N_23021);
or UO_2217 (O_2217,N_23103,N_23691);
and UO_2218 (O_2218,N_24971,N_23244);
nand UO_2219 (O_2219,N_23660,N_23326);
nand UO_2220 (O_2220,N_23236,N_23504);
and UO_2221 (O_2221,N_24020,N_23523);
or UO_2222 (O_2222,N_23725,N_24822);
nor UO_2223 (O_2223,N_24905,N_24240);
nor UO_2224 (O_2224,N_23949,N_24530);
nand UO_2225 (O_2225,N_22724,N_23443);
or UO_2226 (O_2226,N_23242,N_24051);
or UO_2227 (O_2227,N_23516,N_24284);
or UO_2228 (O_2228,N_23006,N_23554);
or UO_2229 (O_2229,N_24204,N_24001);
or UO_2230 (O_2230,N_24478,N_24793);
and UO_2231 (O_2231,N_22810,N_22835);
nor UO_2232 (O_2232,N_23014,N_24748);
or UO_2233 (O_2233,N_24221,N_24313);
nor UO_2234 (O_2234,N_23169,N_23665);
or UO_2235 (O_2235,N_24642,N_24610);
or UO_2236 (O_2236,N_23660,N_24262);
or UO_2237 (O_2237,N_23736,N_23476);
nor UO_2238 (O_2238,N_23314,N_23497);
and UO_2239 (O_2239,N_23080,N_24754);
nor UO_2240 (O_2240,N_24669,N_24325);
nor UO_2241 (O_2241,N_24927,N_22673);
and UO_2242 (O_2242,N_24348,N_23923);
and UO_2243 (O_2243,N_22517,N_22819);
or UO_2244 (O_2244,N_24526,N_24912);
or UO_2245 (O_2245,N_24220,N_23825);
and UO_2246 (O_2246,N_24341,N_23801);
or UO_2247 (O_2247,N_24848,N_24539);
nand UO_2248 (O_2248,N_23157,N_23814);
nand UO_2249 (O_2249,N_22538,N_23079);
nand UO_2250 (O_2250,N_22779,N_23394);
nor UO_2251 (O_2251,N_24627,N_22565);
nor UO_2252 (O_2252,N_22767,N_23467);
or UO_2253 (O_2253,N_24380,N_24260);
nand UO_2254 (O_2254,N_24203,N_24516);
nand UO_2255 (O_2255,N_23282,N_23709);
nor UO_2256 (O_2256,N_24451,N_22932);
nor UO_2257 (O_2257,N_23206,N_23091);
nand UO_2258 (O_2258,N_22675,N_24832);
nor UO_2259 (O_2259,N_24394,N_24387);
and UO_2260 (O_2260,N_24723,N_22840);
nand UO_2261 (O_2261,N_22677,N_23325);
and UO_2262 (O_2262,N_23985,N_23843);
or UO_2263 (O_2263,N_22769,N_23525);
nand UO_2264 (O_2264,N_22876,N_24807);
or UO_2265 (O_2265,N_24724,N_23032);
nand UO_2266 (O_2266,N_24497,N_22965);
and UO_2267 (O_2267,N_22643,N_23985);
nand UO_2268 (O_2268,N_23711,N_23931);
nand UO_2269 (O_2269,N_22830,N_23214);
and UO_2270 (O_2270,N_23122,N_23725);
nor UO_2271 (O_2271,N_22710,N_23777);
nand UO_2272 (O_2272,N_23425,N_22559);
xor UO_2273 (O_2273,N_23299,N_23903);
or UO_2274 (O_2274,N_23476,N_23426);
and UO_2275 (O_2275,N_22929,N_24044);
nand UO_2276 (O_2276,N_23826,N_23577);
nor UO_2277 (O_2277,N_23834,N_24790);
nor UO_2278 (O_2278,N_24643,N_23337);
nand UO_2279 (O_2279,N_23027,N_22960);
and UO_2280 (O_2280,N_23729,N_24396);
nor UO_2281 (O_2281,N_23712,N_23516);
or UO_2282 (O_2282,N_24944,N_24746);
and UO_2283 (O_2283,N_23145,N_24054);
or UO_2284 (O_2284,N_23807,N_24877);
nor UO_2285 (O_2285,N_23707,N_23426);
and UO_2286 (O_2286,N_23609,N_22517);
nor UO_2287 (O_2287,N_24020,N_23992);
nor UO_2288 (O_2288,N_23038,N_23070);
nand UO_2289 (O_2289,N_24846,N_24025);
and UO_2290 (O_2290,N_22744,N_24950);
nand UO_2291 (O_2291,N_24879,N_23529);
and UO_2292 (O_2292,N_22982,N_23348);
nand UO_2293 (O_2293,N_22962,N_23005);
nor UO_2294 (O_2294,N_24808,N_23205);
and UO_2295 (O_2295,N_23772,N_23137);
nor UO_2296 (O_2296,N_23875,N_24265);
nor UO_2297 (O_2297,N_22721,N_24080);
nor UO_2298 (O_2298,N_23841,N_23236);
and UO_2299 (O_2299,N_24532,N_24277);
and UO_2300 (O_2300,N_23843,N_24834);
or UO_2301 (O_2301,N_22989,N_24974);
and UO_2302 (O_2302,N_23859,N_24736);
nand UO_2303 (O_2303,N_24852,N_23025);
and UO_2304 (O_2304,N_23397,N_23115);
or UO_2305 (O_2305,N_23294,N_23289);
and UO_2306 (O_2306,N_24844,N_24703);
nand UO_2307 (O_2307,N_23045,N_23329);
or UO_2308 (O_2308,N_24559,N_24482);
or UO_2309 (O_2309,N_23940,N_24952);
and UO_2310 (O_2310,N_22706,N_22860);
nor UO_2311 (O_2311,N_23783,N_22517);
and UO_2312 (O_2312,N_24597,N_22854);
and UO_2313 (O_2313,N_24931,N_24855);
nor UO_2314 (O_2314,N_23671,N_22654);
and UO_2315 (O_2315,N_23689,N_24480);
nor UO_2316 (O_2316,N_22634,N_24107);
or UO_2317 (O_2317,N_24085,N_23186);
or UO_2318 (O_2318,N_23620,N_22700);
nand UO_2319 (O_2319,N_22860,N_23933);
or UO_2320 (O_2320,N_24785,N_22583);
nor UO_2321 (O_2321,N_24221,N_24886);
and UO_2322 (O_2322,N_24738,N_23174);
and UO_2323 (O_2323,N_23897,N_23255);
or UO_2324 (O_2324,N_22930,N_24172);
nor UO_2325 (O_2325,N_23124,N_23301);
or UO_2326 (O_2326,N_24369,N_22656);
nor UO_2327 (O_2327,N_23709,N_22693);
or UO_2328 (O_2328,N_22638,N_22923);
and UO_2329 (O_2329,N_22899,N_23663);
nor UO_2330 (O_2330,N_22718,N_24900);
nand UO_2331 (O_2331,N_24750,N_23667);
or UO_2332 (O_2332,N_23900,N_23839);
or UO_2333 (O_2333,N_24893,N_22602);
and UO_2334 (O_2334,N_23377,N_24721);
nor UO_2335 (O_2335,N_23416,N_24189);
nand UO_2336 (O_2336,N_24024,N_22979);
nor UO_2337 (O_2337,N_24706,N_24708);
nand UO_2338 (O_2338,N_22759,N_23664);
nor UO_2339 (O_2339,N_22750,N_23420);
or UO_2340 (O_2340,N_23171,N_24134);
nand UO_2341 (O_2341,N_23012,N_24227);
nand UO_2342 (O_2342,N_23727,N_24744);
or UO_2343 (O_2343,N_23543,N_23510);
nor UO_2344 (O_2344,N_24348,N_23980);
or UO_2345 (O_2345,N_23048,N_23725);
or UO_2346 (O_2346,N_22692,N_24917);
nor UO_2347 (O_2347,N_24328,N_23161);
nor UO_2348 (O_2348,N_23830,N_23986);
and UO_2349 (O_2349,N_23013,N_22995);
nand UO_2350 (O_2350,N_23906,N_23032);
nor UO_2351 (O_2351,N_23795,N_24303);
and UO_2352 (O_2352,N_23885,N_24604);
or UO_2353 (O_2353,N_23068,N_23257);
and UO_2354 (O_2354,N_24887,N_24763);
or UO_2355 (O_2355,N_23502,N_23087);
nand UO_2356 (O_2356,N_24720,N_24385);
and UO_2357 (O_2357,N_24239,N_24799);
or UO_2358 (O_2358,N_22803,N_23601);
nand UO_2359 (O_2359,N_22777,N_22961);
nor UO_2360 (O_2360,N_22732,N_22974);
and UO_2361 (O_2361,N_24334,N_22989);
and UO_2362 (O_2362,N_24764,N_23912);
nand UO_2363 (O_2363,N_23712,N_23938);
and UO_2364 (O_2364,N_24085,N_22780);
and UO_2365 (O_2365,N_23497,N_24085);
and UO_2366 (O_2366,N_22947,N_23886);
nor UO_2367 (O_2367,N_24258,N_22833);
nand UO_2368 (O_2368,N_23747,N_24150);
or UO_2369 (O_2369,N_23354,N_23008);
or UO_2370 (O_2370,N_24388,N_24351);
or UO_2371 (O_2371,N_24950,N_24374);
and UO_2372 (O_2372,N_22674,N_23981);
or UO_2373 (O_2373,N_24743,N_22577);
nand UO_2374 (O_2374,N_24430,N_23461);
and UO_2375 (O_2375,N_23767,N_24214);
or UO_2376 (O_2376,N_24794,N_24763);
xnor UO_2377 (O_2377,N_24485,N_22715);
and UO_2378 (O_2378,N_24413,N_24686);
or UO_2379 (O_2379,N_23958,N_24951);
and UO_2380 (O_2380,N_24798,N_23298);
nor UO_2381 (O_2381,N_23299,N_23555);
and UO_2382 (O_2382,N_23084,N_23500);
nor UO_2383 (O_2383,N_24906,N_22793);
nor UO_2384 (O_2384,N_23539,N_23000);
nor UO_2385 (O_2385,N_22689,N_23596);
nor UO_2386 (O_2386,N_22706,N_24156);
nand UO_2387 (O_2387,N_22994,N_24903);
nor UO_2388 (O_2388,N_22527,N_24548);
nand UO_2389 (O_2389,N_22565,N_22959);
and UO_2390 (O_2390,N_22511,N_23875);
xnor UO_2391 (O_2391,N_24937,N_24307);
nor UO_2392 (O_2392,N_24139,N_23978);
or UO_2393 (O_2393,N_24804,N_24490);
and UO_2394 (O_2394,N_24624,N_24251);
and UO_2395 (O_2395,N_23199,N_24381);
and UO_2396 (O_2396,N_24299,N_22998);
nor UO_2397 (O_2397,N_24569,N_24045);
nand UO_2398 (O_2398,N_23618,N_24678);
nor UO_2399 (O_2399,N_22907,N_22720);
and UO_2400 (O_2400,N_22783,N_24134);
nor UO_2401 (O_2401,N_24876,N_23112);
nor UO_2402 (O_2402,N_24307,N_22531);
or UO_2403 (O_2403,N_24858,N_24193);
and UO_2404 (O_2404,N_24816,N_23208);
nor UO_2405 (O_2405,N_23825,N_24959);
and UO_2406 (O_2406,N_22697,N_23579);
or UO_2407 (O_2407,N_24105,N_23871);
or UO_2408 (O_2408,N_22657,N_23145);
nor UO_2409 (O_2409,N_24579,N_23993);
or UO_2410 (O_2410,N_23057,N_23525);
or UO_2411 (O_2411,N_22933,N_22977);
nor UO_2412 (O_2412,N_24368,N_24067);
and UO_2413 (O_2413,N_22992,N_24487);
and UO_2414 (O_2414,N_24442,N_24743);
and UO_2415 (O_2415,N_23556,N_24167);
nor UO_2416 (O_2416,N_24932,N_22581);
or UO_2417 (O_2417,N_23114,N_22501);
xnor UO_2418 (O_2418,N_23773,N_23519);
nand UO_2419 (O_2419,N_23926,N_24049);
nor UO_2420 (O_2420,N_22623,N_23360);
xor UO_2421 (O_2421,N_23871,N_23701);
nor UO_2422 (O_2422,N_24709,N_22778);
and UO_2423 (O_2423,N_24678,N_23718);
nor UO_2424 (O_2424,N_23168,N_24900);
and UO_2425 (O_2425,N_23414,N_22864);
nor UO_2426 (O_2426,N_24493,N_23462);
and UO_2427 (O_2427,N_23413,N_23027);
and UO_2428 (O_2428,N_23434,N_23428);
nor UO_2429 (O_2429,N_23277,N_22645);
nor UO_2430 (O_2430,N_23551,N_24216);
nand UO_2431 (O_2431,N_22844,N_22606);
nor UO_2432 (O_2432,N_23303,N_22927);
nor UO_2433 (O_2433,N_24911,N_24703);
nor UO_2434 (O_2434,N_24447,N_24330);
or UO_2435 (O_2435,N_22936,N_22977);
xnor UO_2436 (O_2436,N_23717,N_23401);
nor UO_2437 (O_2437,N_24513,N_24729);
nor UO_2438 (O_2438,N_24511,N_24491);
or UO_2439 (O_2439,N_23655,N_22748);
nand UO_2440 (O_2440,N_23857,N_24581);
nand UO_2441 (O_2441,N_23342,N_24477);
nor UO_2442 (O_2442,N_23550,N_23349);
nand UO_2443 (O_2443,N_24023,N_23233);
nor UO_2444 (O_2444,N_23220,N_23256);
and UO_2445 (O_2445,N_23841,N_23938);
and UO_2446 (O_2446,N_23123,N_24770);
nor UO_2447 (O_2447,N_24958,N_24125);
nand UO_2448 (O_2448,N_23069,N_22795);
nand UO_2449 (O_2449,N_23529,N_24671);
nor UO_2450 (O_2450,N_23974,N_24422);
xor UO_2451 (O_2451,N_22882,N_23695);
nor UO_2452 (O_2452,N_24540,N_22621);
or UO_2453 (O_2453,N_24049,N_22981);
and UO_2454 (O_2454,N_23586,N_23981);
nand UO_2455 (O_2455,N_24451,N_24436);
nor UO_2456 (O_2456,N_23987,N_23020);
nand UO_2457 (O_2457,N_23999,N_24469);
nand UO_2458 (O_2458,N_22965,N_22712);
or UO_2459 (O_2459,N_24554,N_23615);
and UO_2460 (O_2460,N_24843,N_22656);
or UO_2461 (O_2461,N_24906,N_22570);
nand UO_2462 (O_2462,N_23438,N_24172);
nand UO_2463 (O_2463,N_22886,N_24084);
nor UO_2464 (O_2464,N_24583,N_24783);
or UO_2465 (O_2465,N_22993,N_24511);
and UO_2466 (O_2466,N_24274,N_22508);
nand UO_2467 (O_2467,N_24450,N_23987);
nand UO_2468 (O_2468,N_24286,N_24266);
or UO_2469 (O_2469,N_23459,N_22574);
nor UO_2470 (O_2470,N_24089,N_24321);
nand UO_2471 (O_2471,N_24511,N_24972);
or UO_2472 (O_2472,N_22965,N_23882);
and UO_2473 (O_2473,N_24855,N_23850);
and UO_2474 (O_2474,N_24334,N_23763);
and UO_2475 (O_2475,N_23002,N_22531);
nor UO_2476 (O_2476,N_23457,N_23715);
or UO_2477 (O_2477,N_23693,N_23373);
and UO_2478 (O_2478,N_23725,N_23313);
xor UO_2479 (O_2479,N_22771,N_22638);
nor UO_2480 (O_2480,N_24825,N_24811);
or UO_2481 (O_2481,N_22876,N_24247);
and UO_2482 (O_2482,N_24628,N_24916);
and UO_2483 (O_2483,N_23713,N_24675);
or UO_2484 (O_2484,N_23716,N_23158);
or UO_2485 (O_2485,N_23192,N_24441);
nand UO_2486 (O_2486,N_22677,N_23418);
nor UO_2487 (O_2487,N_23521,N_23792);
nor UO_2488 (O_2488,N_24340,N_23247);
nor UO_2489 (O_2489,N_22925,N_24873);
nand UO_2490 (O_2490,N_22685,N_22729);
or UO_2491 (O_2491,N_24309,N_24719);
and UO_2492 (O_2492,N_24599,N_22889);
or UO_2493 (O_2493,N_22552,N_24787);
nand UO_2494 (O_2494,N_23730,N_22994);
and UO_2495 (O_2495,N_22921,N_23968);
nor UO_2496 (O_2496,N_24327,N_24139);
or UO_2497 (O_2497,N_24892,N_24694);
and UO_2498 (O_2498,N_23203,N_24119);
and UO_2499 (O_2499,N_22512,N_23804);
nor UO_2500 (O_2500,N_23668,N_23679);
nand UO_2501 (O_2501,N_24666,N_22541);
or UO_2502 (O_2502,N_23342,N_24369);
and UO_2503 (O_2503,N_23638,N_23485);
and UO_2504 (O_2504,N_24070,N_23926);
nor UO_2505 (O_2505,N_24683,N_24463);
nand UO_2506 (O_2506,N_22940,N_24380);
nor UO_2507 (O_2507,N_23600,N_23210);
nor UO_2508 (O_2508,N_23521,N_23574);
nor UO_2509 (O_2509,N_24129,N_23444);
nand UO_2510 (O_2510,N_23873,N_22942);
nor UO_2511 (O_2511,N_24909,N_22793);
nor UO_2512 (O_2512,N_24601,N_23371);
or UO_2513 (O_2513,N_24450,N_24088);
nand UO_2514 (O_2514,N_23094,N_24396);
nor UO_2515 (O_2515,N_23770,N_24042);
or UO_2516 (O_2516,N_23363,N_23880);
xnor UO_2517 (O_2517,N_24744,N_24592);
or UO_2518 (O_2518,N_23028,N_24985);
or UO_2519 (O_2519,N_23401,N_22717);
or UO_2520 (O_2520,N_23039,N_24648);
or UO_2521 (O_2521,N_22962,N_24350);
nor UO_2522 (O_2522,N_23304,N_24264);
nand UO_2523 (O_2523,N_23136,N_24719);
or UO_2524 (O_2524,N_23018,N_24127);
or UO_2525 (O_2525,N_24505,N_24045);
and UO_2526 (O_2526,N_24764,N_23306);
nand UO_2527 (O_2527,N_23276,N_22676);
and UO_2528 (O_2528,N_24562,N_23866);
xor UO_2529 (O_2529,N_24492,N_22687);
xnor UO_2530 (O_2530,N_23166,N_24989);
nand UO_2531 (O_2531,N_23245,N_24295);
xnor UO_2532 (O_2532,N_24729,N_22707);
xnor UO_2533 (O_2533,N_23125,N_22517);
or UO_2534 (O_2534,N_24096,N_23108);
nand UO_2535 (O_2535,N_23106,N_24389);
or UO_2536 (O_2536,N_22924,N_24839);
nand UO_2537 (O_2537,N_24959,N_24687);
or UO_2538 (O_2538,N_24872,N_23796);
and UO_2539 (O_2539,N_24485,N_22548);
or UO_2540 (O_2540,N_22628,N_22610);
or UO_2541 (O_2541,N_23313,N_24807);
or UO_2542 (O_2542,N_23733,N_22780);
and UO_2543 (O_2543,N_24497,N_24396);
and UO_2544 (O_2544,N_22806,N_23403);
and UO_2545 (O_2545,N_22865,N_22779);
nor UO_2546 (O_2546,N_24451,N_23692);
nand UO_2547 (O_2547,N_24967,N_24762);
xnor UO_2548 (O_2548,N_24736,N_22546);
nor UO_2549 (O_2549,N_23012,N_24428);
nand UO_2550 (O_2550,N_23413,N_22879);
or UO_2551 (O_2551,N_23319,N_23052);
or UO_2552 (O_2552,N_23678,N_22533);
or UO_2553 (O_2553,N_23273,N_22564);
or UO_2554 (O_2554,N_23279,N_24557);
or UO_2555 (O_2555,N_24304,N_22776);
nand UO_2556 (O_2556,N_22882,N_22915);
nand UO_2557 (O_2557,N_23102,N_24985);
nor UO_2558 (O_2558,N_23647,N_23264);
nor UO_2559 (O_2559,N_24816,N_22810);
and UO_2560 (O_2560,N_23867,N_24610);
or UO_2561 (O_2561,N_24991,N_24156);
or UO_2562 (O_2562,N_24716,N_22933);
or UO_2563 (O_2563,N_22798,N_22893);
nor UO_2564 (O_2564,N_23707,N_23350);
and UO_2565 (O_2565,N_22768,N_23718);
nand UO_2566 (O_2566,N_24467,N_22946);
and UO_2567 (O_2567,N_22523,N_22970);
nor UO_2568 (O_2568,N_24566,N_23701);
nor UO_2569 (O_2569,N_24550,N_22671);
nand UO_2570 (O_2570,N_24385,N_23915);
or UO_2571 (O_2571,N_23586,N_23144);
or UO_2572 (O_2572,N_23480,N_23388);
or UO_2573 (O_2573,N_23127,N_22930);
nor UO_2574 (O_2574,N_24065,N_23096);
nand UO_2575 (O_2575,N_23824,N_24625);
nand UO_2576 (O_2576,N_23209,N_24706);
nor UO_2577 (O_2577,N_24788,N_23786);
or UO_2578 (O_2578,N_22939,N_24256);
and UO_2579 (O_2579,N_24125,N_22884);
nand UO_2580 (O_2580,N_23057,N_24728);
nand UO_2581 (O_2581,N_22637,N_24664);
xnor UO_2582 (O_2582,N_23970,N_24199);
nor UO_2583 (O_2583,N_23625,N_23181);
nand UO_2584 (O_2584,N_22825,N_23575);
or UO_2585 (O_2585,N_24107,N_23004);
or UO_2586 (O_2586,N_24205,N_24041);
nor UO_2587 (O_2587,N_23589,N_23230);
nor UO_2588 (O_2588,N_22908,N_24839);
nor UO_2589 (O_2589,N_24540,N_24378);
and UO_2590 (O_2590,N_22576,N_23376);
nand UO_2591 (O_2591,N_23615,N_23293);
and UO_2592 (O_2592,N_23310,N_24240);
nand UO_2593 (O_2593,N_23765,N_23803);
or UO_2594 (O_2594,N_23921,N_23245);
or UO_2595 (O_2595,N_22860,N_23655);
and UO_2596 (O_2596,N_24903,N_24472);
nand UO_2597 (O_2597,N_22548,N_23375);
nor UO_2598 (O_2598,N_24279,N_24302);
nand UO_2599 (O_2599,N_24470,N_23874);
nor UO_2600 (O_2600,N_22908,N_23475);
nor UO_2601 (O_2601,N_24742,N_22679);
and UO_2602 (O_2602,N_24163,N_23889);
or UO_2603 (O_2603,N_23024,N_22603);
or UO_2604 (O_2604,N_23587,N_24836);
or UO_2605 (O_2605,N_24523,N_23211);
nor UO_2606 (O_2606,N_23708,N_22599);
xnor UO_2607 (O_2607,N_24821,N_23508);
xnor UO_2608 (O_2608,N_24252,N_24823);
xnor UO_2609 (O_2609,N_22592,N_22524);
and UO_2610 (O_2610,N_22846,N_23032);
nand UO_2611 (O_2611,N_24854,N_23601);
and UO_2612 (O_2612,N_24437,N_23124);
or UO_2613 (O_2613,N_23281,N_24529);
and UO_2614 (O_2614,N_24529,N_24444);
nor UO_2615 (O_2615,N_23696,N_24607);
nor UO_2616 (O_2616,N_24882,N_24172);
or UO_2617 (O_2617,N_23926,N_23588);
or UO_2618 (O_2618,N_23826,N_23653);
nand UO_2619 (O_2619,N_24982,N_23767);
or UO_2620 (O_2620,N_24462,N_24452);
nor UO_2621 (O_2621,N_24850,N_24687);
nand UO_2622 (O_2622,N_24118,N_23702);
nor UO_2623 (O_2623,N_22650,N_24272);
nor UO_2624 (O_2624,N_24826,N_22626);
nor UO_2625 (O_2625,N_23083,N_24772);
nand UO_2626 (O_2626,N_23264,N_22936);
and UO_2627 (O_2627,N_23322,N_24008);
nor UO_2628 (O_2628,N_23211,N_24993);
xnor UO_2629 (O_2629,N_24401,N_23697);
nand UO_2630 (O_2630,N_23228,N_23506);
nand UO_2631 (O_2631,N_23205,N_24104);
xnor UO_2632 (O_2632,N_22850,N_24408);
and UO_2633 (O_2633,N_24587,N_23190);
and UO_2634 (O_2634,N_23160,N_22554);
or UO_2635 (O_2635,N_23576,N_24883);
nand UO_2636 (O_2636,N_23563,N_23884);
xor UO_2637 (O_2637,N_23904,N_24772);
nor UO_2638 (O_2638,N_23357,N_24278);
nand UO_2639 (O_2639,N_23582,N_24522);
nor UO_2640 (O_2640,N_23682,N_24310);
nor UO_2641 (O_2641,N_24907,N_23341);
and UO_2642 (O_2642,N_24347,N_22526);
nand UO_2643 (O_2643,N_22843,N_24784);
nor UO_2644 (O_2644,N_23562,N_24004);
or UO_2645 (O_2645,N_23318,N_24982);
xnor UO_2646 (O_2646,N_24308,N_24455);
or UO_2647 (O_2647,N_22935,N_24170);
nor UO_2648 (O_2648,N_23081,N_24958);
or UO_2649 (O_2649,N_23403,N_23317);
and UO_2650 (O_2650,N_24137,N_24579);
nor UO_2651 (O_2651,N_23264,N_23716);
or UO_2652 (O_2652,N_22587,N_23107);
nand UO_2653 (O_2653,N_22790,N_24954);
and UO_2654 (O_2654,N_23751,N_23085);
or UO_2655 (O_2655,N_22851,N_24519);
nor UO_2656 (O_2656,N_23435,N_23880);
and UO_2657 (O_2657,N_23193,N_24773);
nand UO_2658 (O_2658,N_23322,N_22571);
and UO_2659 (O_2659,N_23655,N_24273);
nand UO_2660 (O_2660,N_24047,N_23028);
nand UO_2661 (O_2661,N_24554,N_22969);
and UO_2662 (O_2662,N_24183,N_22586);
nand UO_2663 (O_2663,N_23123,N_24201);
and UO_2664 (O_2664,N_24419,N_23671);
xnor UO_2665 (O_2665,N_24306,N_23335);
nand UO_2666 (O_2666,N_23703,N_22708);
or UO_2667 (O_2667,N_24878,N_24276);
and UO_2668 (O_2668,N_23274,N_24211);
nor UO_2669 (O_2669,N_23927,N_24036);
and UO_2670 (O_2670,N_24952,N_22527);
nand UO_2671 (O_2671,N_23948,N_24771);
and UO_2672 (O_2672,N_22817,N_23131);
or UO_2673 (O_2673,N_23741,N_23928);
nand UO_2674 (O_2674,N_23230,N_23263);
nand UO_2675 (O_2675,N_23735,N_22767);
or UO_2676 (O_2676,N_22562,N_23289);
nand UO_2677 (O_2677,N_24161,N_23990);
nand UO_2678 (O_2678,N_23130,N_24765);
nand UO_2679 (O_2679,N_23082,N_24513);
or UO_2680 (O_2680,N_23058,N_23371);
nand UO_2681 (O_2681,N_23034,N_23067);
nand UO_2682 (O_2682,N_24401,N_24415);
nand UO_2683 (O_2683,N_24086,N_24006);
nor UO_2684 (O_2684,N_22591,N_22522);
and UO_2685 (O_2685,N_23515,N_24593);
nand UO_2686 (O_2686,N_24265,N_23152);
and UO_2687 (O_2687,N_24958,N_24420);
or UO_2688 (O_2688,N_24814,N_24060);
nor UO_2689 (O_2689,N_24163,N_22671);
nand UO_2690 (O_2690,N_24454,N_23280);
or UO_2691 (O_2691,N_23762,N_23918);
or UO_2692 (O_2692,N_22660,N_24907);
and UO_2693 (O_2693,N_23157,N_22539);
nand UO_2694 (O_2694,N_24789,N_23676);
nor UO_2695 (O_2695,N_24985,N_24118);
nand UO_2696 (O_2696,N_23662,N_24193);
nor UO_2697 (O_2697,N_24500,N_23610);
or UO_2698 (O_2698,N_24701,N_22686);
nand UO_2699 (O_2699,N_23266,N_24395);
or UO_2700 (O_2700,N_23822,N_22526);
nand UO_2701 (O_2701,N_23913,N_23447);
nor UO_2702 (O_2702,N_24453,N_23109);
or UO_2703 (O_2703,N_23256,N_23312);
nor UO_2704 (O_2704,N_23408,N_23763);
nor UO_2705 (O_2705,N_24191,N_24274);
and UO_2706 (O_2706,N_24040,N_24305);
and UO_2707 (O_2707,N_23725,N_23963);
or UO_2708 (O_2708,N_23338,N_24965);
nor UO_2709 (O_2709,N_24014,N_24676);
or UO_2710 (O_2710,N_23570,N_22608);
and UO_2711 (O_2711,N_24309,N_23685);
nand UO_2712 (O_2712,N_22852,N_24652);
nor UO_2713 (O_2713,N_24926,N_24952);
and UO_2714 (O_2714,N_22909,N_23455);
or UO_2715 (O_2715,N_23144,N_22765);
nand UO_2716 (O_2716,N_22944,N_22984);
or UO_2717 (O_2717,N_22765,N_23101);
nor UO_2718 (O_2718,N_22700,N_23939);
nor UO_2719 (O_2719,N_23344,N_24136);
nor UO_2720 (O_2720,N_22971,N_24900);
and UO_2721 (O_2721,N_22530,N_24497);
nor UO_2722 (O_2722,N_24779,N_22679);
or UO_2723 (O_2723,N_24640,N_22902);
or UO_2724 (O_2724,N_24462,N_23053);
nand UO_2725 (O_2725,N_24773,N_23362);
or UO_2726 (O_2726,N_24980,N_23253);
or UO_2727 (O_2727,N_24858,N_23889);
and UO_2728 (O_2728,N_22842,N_23636);
nand UO_2729 (O_2729,N_23583,N_24431);
nand UO_2730 (O_2730,N_24446,N_24884);
or UO_2731 (O_2731,N_23909,N_24273);
nor UO_2732 (O_2732,N_22832,N_23306);
nand UO_2733 (O_2733,N_23495,N_22707);
nand UO_2734 (O_2734,N_22613,N_24272);
and UO_2735 (O_2735,N_22979,N_24673);
nor UO_2736 (O_2736,N_23870,N_23440);
or UO_2737 (O_2737,N_23986,N_24686);
or UO_2738 (O_2738,N_23962,N_24805);
nand UO_2739 (O_2739,N_24887,N_23987);
nand UO_2740 (O_2740,N_24749,N_22727);
nor UO_2741 (O_2741,N_24314,N_22810);
and UO_2742 (O_2742,N_24077,N_23075);
nor UO_2743 (O_2743,N_24432,N_23317);
nor UO_2744 (O_2744,N_23915,N_23155);
and UO_2745 (O_2745,N_23712,N_23037);
nand UO_2746 (O_2746,N_24283,N_23015);
nand UO_2747 (O_2747,N_24178,N_24005);
or UO_2748 (O_2748,N_23313,N_23508);
xnor UO_2749 (O_2749,N_24498,N_23087);
or UO_2750 (O_2750,N_23301,N_24392);
nor UO_2751 (O_2751,N_22972,N_23517);
and UO_2752 (O_2752,N_24297,N_23587);
or UO_2753 (O_2753,N_23559,N_24805);
or UO_2754 (O_2754,N_23648,N_24538);
and UO_2755 (O_2755,N_22600,N_23278);
nor UO_2756 (O_2756,N_24299,N_24567);
or UO_2757 (O_2757,N_22587,N_23329);
nor UO_2758 (O_2758,N_24550,N_24583);
and UO_2759 (O_2759,N_22912,N_24361);
or UO_2760 (O_2760,N_24549,N_23724);
or UO_2761 (O_2761,N_24742,N_24261);
xor UO_2762 (O_2762,N_22783,N_22715);
nand UO_2763 (O_2763,N_23246,N_23188);
nor UO_2764 (O_2764,N_23865,N_23453);
and UO_2765 (O_2765,N_22944,N_23160);
and UO_2766 (O_2766,N_22544,N_24442);
nor UO_2767 (O_2767,N_22713,N_23243);
or UO_2768 (O_2768,N_23529,N_24964);
nor UO_2769 (O_2769,N_23899,N_23931);
nor UO_2770 (O_2770,N_24839,N_23989);
nand UO_2771 (O_2771,N_24647,N_24424);
nand UO_2772 (O_2772,N_22749,N_24750);
nand UO_2773 (O_2773,N_24410,N_23208);
nand UO_2774 (O_2774,N_24747,N_24584);
nor UO_2775 (O_2775,N_22762,N_23875);
nor UO_2776 (O_2776,N_22598,N_22967);
nor UO_2777 (O_2777,N_24442,N_23310);
and UO_2778 (O_2778,N_23100,N_24223);
and UO_2779 (O_2779,N_23213,N_24443);
or UO_2780 (O_2780,N_22979,N_23588);
xnor UO_2781 (O_2781,N_22854,N_23393);
nor UO_2782 (O_2782,N_23812,N_24844);
nand UO_2783 (O_2783,N_22989,N_23986);
or UO_2784 (O_2784,N_23767,N_24270);
and UO_2785 (O_2785,N_24049,N_22562);
nor UO_2786 (O_2786,N_24053,N_23509);
and UO_2787 (O_2787,N_22929,N_23613);
or UO_2788 (O_2788,N_24660,N_23060);
xor UO_2789 (O_2789,N_23583,N_24880);
and UO_2790 (O_2790,N_24418,N_24650);
or UO_2791 (O_2791,N_22624,N_23026);
xnor UO_2792 (O_2792,N_23745,N_22516);
and UO_2793 (O_2793,N_23946,N_23497);
or UO_2794 (O_2794,N_23349,N_24258);
or UO_2795 (O_2795,N_24245,N_23575);
or UO_2796 (O_2796,N_24368,N_24631);
and UO_2797 (O_2797,N_23641,N_23819);
and UO_2798 (O_2798,N_23185,N_24968);
nor UO_2799 (O_2799,N_24375,N_23164);
nor UO_2800 (O_2800,N_24057,N_22611);
nor UO_2801 (O_2801,N_23541,N_24633);
and UO_2802 (O_2802,N_22778,N_24579);
or UO_2803 (O_2803,N_22709,N_23018);
nor UO_2804 (O_2804,N_24950,N_24789);
nor UO_2805 (O_2805,N_23590,N_24333);
and UO_2806 (O_2806,N_22812,N_22833);
nand UO_2807 (O_2807,N_24502,N_23510);
nand UO_2808 (O_2808,N_23863,N_24938);
or UO_2809 (O_2809,N_24382,N_23171);
or UO_2810 (O_2810,N_24103,N_24833);
nor UO_2811 (O_2811,N_23198,N_22742);
nor UO_2812 (O_2812,N_24822,N_24634);
or UO_2813 (O_2813,N_22906,N_24086);
or UO_2814 (O_2814,N_22972,N_24415);
and UO_2815 (O_2815,N_23832,N_23684);
nand UO_2816 (O_2816,N_23656,N_24172);
xnor UO_2817 (O_2817,N_22955,N_22934);
and UO_2818 (O_2818,N_23667,N_23192);
or UO_2819 (O_2819,N_22889,N_24445);
nand UO_2820 (O_2820,N_24726,N_23881);
and UO_2821 (O_2821,N_23555,N_23366);
and UO_2822 (O_2822,N_24947,N_24930);
xnor UO_2823 (O_2823,N_24479,N_23416);
and UO_2824 (O_2824,N_23622,N_24811);
nand UO_2825 (O_2825,N_22543,N_23195);
nor UO_2826 (O_2826,N_22877,N_24362);
nand UO_2827 (O_2827,N_23604,N_23520);
nand UO_2828 (O_2828,N_24128,N_23555);
nand UO_2829 (O_2829,N_24228,N_23470);
nand UO_2830 (O_2830,N_24928,N_23331);
and UO_2831 (O_2831,N_23766,N_22705);
nand UO_2832 (O_2832,N_24378,N_23827);
nand UO_2833 (O_2833,N_23131,N_23361);
nor UO_2834 (O_2834,N_22602,N_24548);
or UO_2835 (O_2835,N_23689,N_23614);
nand UO_2836 (O_2836,N_23000,N_23869);
or UO_2837 (O_2837,N_24992,N_24918);
nand UO_2838 (O_2838,N_22874,N_24444);
or UO_2839 (O_2839,N_23594,N_24907);
or UO_2840 (O_2840,N_23877,N_22898);
nand UO_2841 (O_2841,N_22565,N_23408);
nor UO_2842 (O_2842,N_23738,N_23214);
nand UO_2843 (O_2843,N_23708,N_23706);
nand UO_2844 (O_2844,N_23291,N_24997);
nand UO_2845 (O_2845,N_24856,N_23069);
and UO_2846 (O_2846,N_24877,N_23062);
or UO_2847 (O_2847,N_24259,N_23842);
xor UO_2848 (O_2848,N_23854,N_24070);
or UO_2849 (O_2849,N_23411,N_22857);
nor UO_2850 (O_2850,N_23346,N_24806);
xnor UO_2851 (O_2851,N_24528,N_22610);
or UO_2852 (O_2852,N_24535,N_24850);
nor UO_2853 (O_2853,N_23192,N_22753);
nand UO_2854 (O_2854,N_24642,N_23685);
nor UO_2855 (O_2855,N_23465,N_22656);
or UO_2856 (O_2856,N_24728,N_24502);
and UO_2857 (O_2857,N_24239,N_23693);
nand UO_2858 (O_2858,N_24680,N_23704);
and UO_2859 (O_2859,N_23858,N_23630);
or UO_2860 (O_2860,N_23406,N_24063);
or UO_2861 (O_2861,N_23438,N_23215);
and UO_2862 (O_2862,N_24137,N_23539);
or UO_2863 (O_2863,N_24681,N_24240);
nor UO_2864 (O_2864,N_22537,N_23298);
or UO_2865 (O_2865,N_23006,N_24767);
xnor UO_2866 (O_2866,N_24427,N_23372);
or UO_2867 (O_2867,N_22969,N_22626);
or UO_2868 (O_2868,N_22566,N_23516);
nor UO_2869 (O_2869,N_23138,N_24904);
and UO_2870 (O_2870,N_23635,N_23533);
nor UO_2871 (O_2871,N_23296,N_24210);
and UO_2872 (O_2872,N_22929,N_24705);
nor UO_2873 (O_2873,N_24033,N_22738);
nor UO_2874 (O_2874,N_22524,N_23469);
or UO_2875 (O_2875,N_24043,N_24670);
or UO_2876 (O_2876,N_22635,N_24634);
nand UO_2877 (O_2877,N_23848,N_23306);
and UO_2878 (O_2878,N_23614,N_24335);
or UO_2879 (O_2879,N_24154,N_22636);
nand UO_2880 (O_2880,N_22938,N_24443);
xor UO_2881 (O_2881,N_24763,N_22553);
and UO_2882 (O_2882,N_23720,N_24420);
and UO_2883 (O_2883,N_24473,N_22859);
and UO_2884 (O_2884,N_22727,N_24460);
and UO_2885 (O_2885,N_22670,N_23447);
nor UO_2886 (O_2886,N_23931,N_24209);
xor UO_2887 (O_2887,N_23094,N_24184);
nand UO_2888 (O_2888,N_24556,N_23224);
and UO_2889 (O_2889,N_23296,N_22704);
nor UO_2890 (O_2890,N_24134,N_23555);
or UO_2891 (O_2891,N_22729,N_23403);
nor UO_2892 (O_2892,N_24012,N_24005);
or UO_2893 (O_2893,N_24666,N_23004);
and UO_2894 (O_2894,N_22901,N_23856);
or UO_2895 (O_2895,N_24039,N_22684);
nor UO_2896 (O_2896,N_24806,N_24653);
and UO_2897 (O_2897,N_24001,N_24576);
or UO_2898 (O_2898,N_23478,N_23196);
and UO_2899 (O_2899,N_24566,N_23770);
or UO_2900 (O_2900,N_24721,N_22632);
and UO_2901 (O_2901,N_22766,N_22602);
nor UO_2902 (O_2902,N_23504,N_23001);
and UO_2903 (O_2903,N_24771,N_23069);
nand UO_2904 (O_2904,N_22593,N_24401);
and UO_2905 (O_2905,N_23599,N_24694);
nor UO_2906 (O_2906,N_23882,N_23919);
or UO_2907 (O_2907,N_24306,N_24523);
or UO_2908 (O_2908,N_22939,N_23975);
and UO_2909 (O_2909,N_23301,N_23860);
and UO_2910 (O_2910,N_23243,N_22861);
nor UO_2911 (O_2911,N_23184,N_24995);
and UO_2912 (O_2912,N_22534,N_24974);
or UO_2913 (O_2913,N_24726,N_24587);
and UO_2914 (O_2914,N_24330,N_24671);
nor UO_2915 (O_2915,N_23239,N_23765);
and UO_2916 (O_2916,N_23431,N_23189);
or UO_2917 (O_2917,N_24286,N_24913);
nand UO_2918 (O_2918,N_22901,N_24916);
xnor UO_2919 (O_2919,N_24502,N_24553);
nand UO_2920 (O_2920,N_24496,N_24837);
and UO_2921 (O_2921,N_24633,N_22890);
and UO_2922 (O_2922,N_24306,N_23001);
or UO_2923 (O_2923,N_22510,N_23463);
nor UO_2924 (O_2924,N_24897,N_24967);
nand UO_2925 (O_2925,N_23415,N_24073);
or UO_2926 (O_2926,N_24387,N_24398);
and UO_2927 (O_2927,N_24179,N_24872);
nor UO_2928 (O_2928,N_23527,N_22501);
and UO_2929 (O_2929,N_23089,N_24165);
and UO_2930 (O_2930,N_23542,N_23168);
and UO_2931 (O_2931,N_23747,N_23494);
and UO_2932 (O_2932,N_23839,N_22864);
and UO_2933 (O_2933,N_24625,N_22527);
and UO_2934 (O_2934,N_22876,N_23875);
nor UO_2935 (O_2935,N_24542,N_23148);
nand UO_2936 (O_2936,N_24249,N_23217);
or UO_2937 (O_2937,N_23066,N_24701);
nor UO_2938 (O_2938,N_24131,N_23827);
and UO_2939 (O_2939,N_23060,N_23726);
and UO_2940 (O_2940,N_24459,N_23517);
or UO_2941 (O_2941,N_23961,N_23128);
and UO_2942 (O_2942,N_24317,N_24964);
and UO_2943 (O_2943,N_23420,N_23416);
nand UO_2944 (O_2944,N_22517,N_24048);
and UO_2945 (O_2945,N_23801,N_22509);
nand UO_2946 (O_2946,N_24053,N_24401);
nand UO_2947 (O_2947,N_24854,N_24381);
xor UO_2948 (O_2948,N_24477,N_23822);
xnor UO_2949 (O_2949,N_24157,N_23912);
nand UO_2950 (O_2950,N_24104,N_23852);
nand UO_2951 (O_2951,N_24654,N_23890);
and UO_2952 (O_2952,N_22763,N_23572);
nor UO_2953 (O_2953,N_24749,N_24575);
or UO_2954 (O_2954,N_24052,N_23819);
and UO_2955 (O_2955,N_24869,N_23833);
nand UO_2956 (O_2956,N_22933,N_24151);
or UO_2957 (O_2957,N_22949,N_22683);
nand UO_2958 (O_2958,N_24298,N_23385);
or UO_2959 (O_2959,N_22963,N_22699);
and UO_2960 (O_2960,N_22886,N_23724);
or UO_2961 (O_2961,N_22891,N_23997);
or UO_2962 (O_2962,N_23588,N_24098);
nor UO_2963 (O_2963,N_22679,N_23987);
nand UO_2964 (O_2964,N_24593,N_24523);
nor UO_2965 (O_2965,N_24942,N_24090);
nand UO_2966 (O_2966,N_22855,N_24883);
nand UO_2967 (O_2967,N_23753,N_24593);
and UO_2968 (O_2968,N_22703,N_23598);
and UO_2969 (O_2969,N_24956,N_23938);
nand UO_2970 (O_2970,N_24221,N_23207);
or UO_2971 (O_2971,N_22989,N_22904);
and UO_2972 (O_2972,N_24394,N_24306);
and UO_2973 (O_2973,N_23001,N_24246);
or UO_2974 (O_2974,N_24730,N_24561);
nand UO_2975 (O_2975,N_22936,N_23901);
nor UO_2976 (O_2976,N_24141,N_23287);
or UO_2977 (O_2977,N_24990,N_23514);
and UO_2978 (O_2978,N_24531,N_22667);
nand UO_2979 (O_2979,N_23675,N_22624);
and UO_2980 (O_2980,N_24655,N_22701);
and UO_2981 (O_2981,N_24140,N_22578);
nor UO_2982 (O_2982,N_22505,N_24279);
or UO_2983 (O_2983,N_23048,N_22781);
nand UO_2984 (O_2984,N_23486,N_24329);
nor UO_2985 (O_2985,N_22653,N_23574);
and UO_2986 (O_2986,N_23310,N_24185);
or UO_2987 (O_2987,N_24498,N_23444);
or UO_2988 (O_2988,N_24103,N_23799);
nand UO_2989 (O_2989,N_23352,N_24235);
and UO_2990 (O_2990,N_24590,N_23101);
nand UO_2991 (O_2991,N_24571,N_23816);
or UO_2992 (O_2992,N_23242,N_23112);
and UO_2993 (O_2993,N_23039,N_24378);
nand UO_2994 (O_2994,N_22676,N_23870);
nor UO_2995 (O_2995,N_23939,N_24938);
and UO_2996 (O_2996,N_22604,N_22619);
and UO_2997 (O_2997,N_22836,N_22764);
or UO_2998 (O_2998,N_23452,N_24748);
or UO_2999 (O_2999,N_24565,N_24527);
endmodule