module basic_1500_15000_2000_50_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_386,In_1293);
xor U1 (N_1,In_1269,In_1097);
nand U2 (N_2,In_667,In_1177);
nor U3 (N_3,In_709,In_1286);
or U4 (N_4,In_440,In_1290);
nand U5 (N_5,In_941,In_394);
nor U6 (N_6,In_28,In_756);
or U7 (N_7,In_335,In_1429);
and U8 (N_8,In_920,In_1197);
xnor U9 (N_9,In_1476,In_727);
or U10 (N_10,In_147,In_34);
or U11 (N_11,In_1417,In_1003);
nor U12 (N_12,In_928,In_1173);
or U13 (N_13,In_215,In_229);
xor U14 (N_14,In_745,In_927);
nand U15 (N_15,In_1015,In_644);
xnor U16 (N_16,In_155,In_411);
nand U17 (N_17,In_1115,In_647);
or U18 (N_18,In_843,In_429);
xnor U19 (N_19,In_1331,In_111);
and U20 (N_20,In_49,In_255);
nor U21 (N_21,In_555,In_8);
or U22 (N_22,In_403,In_1186);
or U23 (N_23,In_252,In_445);
nor U24 (N_24,In_1227,In_1165);
or U25 (N_25,In_878,In_1270);
and U26 (N_26,In_113,In_295);
nor U27 (N_27,In_880,In_862);
nand U28 (N_28,In_391,In_1248);
xnor U29 (N_29,In_782,In_686);
and U30 (N_30,In_580,In_72);
xor U31 (N_31,In_1253,In_17);
xnor U32 (N_32,In_636,In_1088);
and U33 (N_33,In_237,In_856);
xnor U34 (N_34,In_160,In_733);
nor U35 (N_35,In_506,In_951);
nand U36 (N_36,In_0,In_109);
and U37 (N_37,In_275,In_973);
and U38 (N_38,In_62,In_39);
and U39 (N_39,In_1171,In_785);
xor U40 (N_40,In_1163,In_765);
and U41 (N_41,In_1013,In_1355);
and U42 (N_42,In_1378,In_485);
nor U43 (N_43,In_1243,In_406);
xnor U44 (N_44,In_57,In_979);
nand U45 (N_45,In_1334,In_286);
xor U46 (N_46,In_194,In_1235);
and U47 (N_47,In_866,In_990);
or U48 (N_48,In_190,In_422);
and U49 (N_49,In_371,In_730);
xnor U50 (N_50,In_400,In_248);
nor U51 (N_51,In_1296,In_1387);
or U52 (N_52,In_899,In_1279);
or U53 (N_53,In_1313,In_211);
nand U54 (N_54,In_337,In_495);
nor U55 (N_55,In_724,In_1374);
nand U56 (N_56,In_274,In_232);
or U57 (N_57,In_1388,In_330);
nand U58 (N_58,In_1112,In_1477);
xor U59 (N_59,In_616,In_463);
or U60 (N_60,In_932,In_914);
nor U61 (N_61,In_1246,In_1300);
and U62 (N_62,In_1001,In_1025);
nor U63 (N_63,In_638,In_235);
or U64 (N_64,In_52,In_652);
or U65 (N_65,In_1095,In_283);
or U66 (N_66,In_830,In_369);
xnor U67 (N_67,In_601,In_504);
nor U68 (N_68,In_46,In_768);
nor U69 (N_69,In_379,In_1483);
xor U70 (N_70,In_717,In_712);
nor U71 (N_71,In_1148,In_1376);
and U72 (N_72,In_962,In_632);
or U73 (N_73,In_1481,In_1366);
or U74 (N_74,In_491,In_447);
and U75 (N_75,In_981,In_1326);
and U76 (N_76,In_808,In_493);
or U77 (N_77,In_1098,In_1183);
nand U78 (N_78,In_596,In_245);
xor U79 (N_79,In_895,In_929);
or U80 (N_80,In_1126,In_604);
and U81 (N_81,In_1179,In_630);
xnor U82 (N_82,In_633,In_1198);
nand U83 (N_83,In_1049,In_1256);
or U84 (N_84,In_1434,In_790);
and U85 (N_85,In_494,In_313);
and U86 (N_86,In_231,In_1441);
nor U87 (N_87,In_14,In_519);
xor U88 (N_88,In_95,In_964);
or U89 (N_89,In_413,In_1124);
nor U90 (N_90,In_615,In_547);
nor U91 (N_91,In_253,In_937);
or U92 (N_92,In_1192,In_1090);
nand U93 (N_93,In_75,In_346);
xnor U94 (N_94,In_1393,In_935);
xnor U95 (N_95,In_674,In_1223);
nor U96 (N_96,In_404,In_199);
xnor U97 (N_97,In_846,In_1005);
and U98 (N_98,In_870,In_924);
or U99 (N_99,In_1237,In_884);
nor U100 (N_100,In_1428,In_99);
nand U101 (N_101,In_366,In_639);
and U102 (N_102,In_41,In_781);
xor U103 (N_103,In_1475,In_108);
and U104 (N_104,In_287,In_254);
and U105 (N_105,In_530,In_1038);
and U106 (N_106,In_1031,In_967);
nor U107 (N_107,In_691,In_706);
nand U108 (N_108,In_634,In_1405);
or U109 (N_109,In_1278,In_668);
nand U110 (N_110,In_955,In_1101);
and U111 (N_111,In_1046,In_240);
nor U112 (N_112,In_1318,In_364);
xnor U113 (N_113,In_224,In_910);
and U114 (N_114,In_33,In_897);
nand U115 (N_115,In_961,In_261);
nor U116 (N_116,In_1356,In_418);
or U117 (N_117,In_1160,In_236);
nand U118 (N_118,In_760,In_883);
xor U119 (N_119,In_265,In_1258);
nor U120 (N_120,In_1219,In_1487);
or U121 (N_121,In_50,In_584);
or U122 (N_122,In_289,In_200);
and U123 (N_123,In_1080,In_1406);
nand U124 (N_124,In_526,In_581);
nand U125 (N_125,In_110,In_1315);
nand U126 (N_126,In_729,In_350);
nand U127 (N_127,In_693,In_1491);
nor U128 (N_128,In_954,In_621);
or U129 (N_129,In_1130,In_424);
nor U130 (N_130,In_1178,In_999);
nand U131 (N_131,In_1322,In_1480);
and U132 (N_132,In_1415,In_1139);
xor U133 (N_133,In_1207,In_150);
and U134 (N_134,In_351,In_857);
nand U135 (N_135,In_1352,In_757);
nand U136 (N_136,In_262,In_590);
and U137 (N_137,In_1104,In_1363);
nor U138 (N_138,In_1304,In_1255);
nor U139 (N_139,In_1102,In_456);
nor U140 (N_140,In_1340,In_972);
nand U141 (N_141,In_991,In_421);
nand U142 (N_142,In_1037,In_796);
and U143 (N_143,In_6,In_672);
nor U144 (N_144,In_564,In_1348);
nor U145 (N_145,In_436,In_585);
nor U146 (N_146,In_55,In_1051);
nor U147 (N_147,In_101,In_764);
and U148 (N_148,In_1087,In_1027);
or U149 (N_149,In_353,In_741);
nor U150 (N_150,In_690,In_141);
xor U151 (N_151,In_1089,In_1042);
nand U152 (N_152,In_838,In_882);
or U153 (N_153,In_1040,In_901);
nor U154 (N_154,In_356,In_692);
nor U155 (N_155,In_348,In_654);
and U156 (N_156,In_698,In_370);
nand U157 (N_157,In_1189,In_1133);
nor U158 (N_158,In_589,In_1156);
nand U159 (N_159,In_378,In_338);
nor U160 (N_160,In_73,In_334);
and U161 (N_161,In_306,In_340);
nor U162 (N_162,In_855,In_1072);
or U163 (N_163,In_569,In_1041);
and U164 (N_164,In_1064,In_292);
and U165 (N_165,In_67,In_1267);
nor U166 (N_166,In_184,In_812);
or U167 (N_167,In_412,In_1266);
nand U168 (N_168,In_1474,In_68);
and U169 (N_169,In_1377,In_174);
nand U170 (N_170,In_993,In_10);
and U171 (N_171,In_43,In_361);
nor U172 (N_172,In_836,In_169);
and U173 (N_173,In_1209,In_1389);
or U174 (N_174,In_665,In_1022);
or U175 (N_175,In_1368,In_662);
nand U176 (N_176,In_239,In_1347);
nand U177 (N_177,In_571,In_980);
and U178 (N_178,In_544,In_136);
nand U179 (N_179,In_598,In_1048);
and U180 (N_180,In_650,In_1221);
and U181 (N_181,In_688,In_680);
nor U182 (N_182,In_1199,In_343);
and U183 (N_183,In_816,In_323);
and U184 (N_184,In_1118,In_24);
xnor U185 (N_185,In_936,In_517);
xor U186 (N_186,In_1411,In_845);
or U187 (N_187,In_135,In_824);
nand U188 (N_188,In_297,In_1397);
xnor U189 (N_189,In_800,In_1438);
xnor U190 (N_190,In_1229,In_342);
or U191 (N_191,In_627,In_798);
and U192 (N_192,In_282,In_132);
xnor U193 (N_193,In_1435,In_787);
xnor U194 (N_194,In_610,In_1194);
or U195 (N_195,In_1478,In_839);
xnor U196 (N_196,In_1075,In_1402);
nand U197 (N_197,In_763,In_21);
and U198 (N_198,In_1070,In_1215);
and U199 (N_199,In_457,In_820);
xnor U200 (N_200,In_779,In_1424);
nor U201 (N_201,In_892,In_104);
or U202 (N_202,In_1086,In_1181);
and U203 (N_203,In_988,In_1365);
xor U204 (N_204,In_1020,In_202);
xor U205 (N_205,In_1386,In_276);
or U206 (N_206,In_532,In_697);
or U207 (N_207,In_965,In_778);
or U208 (N_208,In_1350,In_122);
nor U209 (N_209,In_689,In_1372);
and U210 (N_210,In_40,In_1230);
nand U211 (N_211,In_791,In_588);
xor U212 (N_212,In_835,In_432);
nor U213 (N_213,In_1360,In_1128);
nand U214 (N_214,In_175,In_1000);
nor U215 (N_215,In_268,In_960);
xnor U216 (N_216,In_1259,In_328);
and U217 (N_217,In_1107,In_1214);
xnor U218 (N_218,In_1451,In_116);
nor U219 (N_219,In_818,In_1362);
and U220 (N_220,In_1079,In_1254);
nand U221 (N_221,In_645,In_944);
xor U222 (N_222,In_79,In_1288);
nand U223 (N_223,In_1157,In_437);
nor U224 (N_224,In_1303,In_1263);
and U225 (N_225,In_948,In_885);
xor U226 (N_226,In_829,In_879);
or U227 (N_227,In_1106,In_701);
and U228 (N_228,In_721,In_933);
nand U229 (N_229,In_1314,In_619);
and U230 (N_230,In_238,In_718);
and U231 (N_231,In_1081,In_696);
nand U232 (N_232,In_625,In_148);
nor U233 (N_233,In_1470,In_687);
and U234 (N_234,In_922,In_320);
nand U235 (N_235,In_1400,In_213);
or U236 (N_236,In_212,In_85);
and U237 (N_237,In_694,In_637);
xnor U238 (N_238,In_1455,In_1419);
and U239 (N_239,In_1301,In_583);
or U240 (N_240,In_195,In_774);
or U241 (N_241,In_209,In_725);
and U242 (N_242,In_217,In_592);
xor U243 (N_243,In_264,In_32);
or U244 (N_244,In_204,In_678);
nand U245 (N_245,In_1463,In_1490);
nand U246 (N_246,In_1002,In_61);
xor U247 (N_247,In_735,In_1467);
or U248 (N_248,In_2,In_871);
xor U249 (N_249,In_290,In_640);
nand U250 (N_250,In_279,In_308);
or U251 (N_251,In_214,In_448);
and U252 (N_252,In_89,In_1358);
nand U253 (N_253,In_548,In_128);
nor U254 (N_254,In_60,In_1325);
xnor U255 (N_255,In_461,In_1203);
or U256 (N_256,In_565,In_464);
or U257 (N_257,In_1494,In_159);
xor U258 (N_258,In_316,In_499);
or U259 (N_259,In_854,In_244);
and U260 (N_260,In_179,In_1091);
nor U261 (N_261,In_620,In_606);
or U262 (N_262,In_989,In_1142);
nor U263 (N_263,In_1496,In_587);
nor U264 (N_264,In_139,In_524);
nand U265 (N_265,In_1423,In_858);
or U266 (N_266,In_522,In_481);
nand U267 (N_267,In_1265,In_918);
and U268 (N_268,In_705,In_984);
or U269 (N_269,In_1457,In_1344);
nor U270 (N_270,In_907,In_1078);
and U271 (N_271,In_30,In_1010);
nand U272 (N_272,In_489,In_1076);
xor U273 (N_273,In_700,In_188);
and U274 (N_274,In_986,In_154);
xor U275 (N_275,In_82,In_134);
and U276 (N_276,In_656,In_842);
xnor U277 (N_277,In_76,In_849);
nor U278 (N_278,In_586,In_1220);
nand U279 (N_279,In_832,In_18);
xor U280 (N_280,In_728,In_917);
nor U281 (N_281,In_266,In_1240);
and U282 (N_282,In_35,In_103);
xor U283 (N_283,In_850,In_1416);
nand U284 (N_284,In_1309,In_607);
nor U285 (N_285,In_575,In_1234);
nand U286 (N_286,In_722,In_1057);
and U287 (N_287,In_574,In_1029);
nor U288 (N_288,In_1446,In_1291);
xnor U289 (N_289,In_1151,In_669);
and U290 (N_290,In_834,In_1082);
nor U291 (N_291,In_227,In_365);
and U292 (N_292,In_864,In_1336);
nand U293 (N_293,In_243,In_1058);
nor U294 (N_294,In_53,In_626);
nand U295 (N_295,In_203,In_950);
nand U296 (N_296,In_71,In_1453);
or U297 (N_297,In_1152,In_1361);
nor U298 (N_298,In_325,In_507);
or U299 (N_299,In_556,In_848);
xnor U300 (N_300,In_1120,In_1131);
nor U301 (N_301,N_110,In_1425);
nand U302 (N_302,In_786,In_1498);
xor U303 (N_303,N_6,In_119);
or U304 (N_304,In_1295,In_172);
nor U305 (N_305,In_624,N_92);
and U306 (N_306,N_244,In_594);
xnor U307 (N_307,In_543,In_987);
nand U308 (N_308,In_515,In_710);
xnor U309 (N_309,In_367,In_1287);
nor U310 (N_310,In_372,In_91);
nand U311 (N_311,In_995,In_1073);
nand U312 (N_312,In_359,In_1052);
nor U313 (N_313,N_56,In_58);
xnor U314 (N_314,In_390,In_152);
nand U315 (N_315,In_1026,In_1384);
or U316 (N_316,In_699,In_285);
or U317 (N_317,In_671,N_72);
nor U318 (N_318,In_1277,In_1135);
nor U319 (N_319,In_431,In_1461);
and U320 (N_320,In_943,N_26);
or U321 (N_321,In_1050,In_501);
xor U322 (N_322,In_271,In_3);
nor U323 (N_323,N_194,In_1273);
nor U324 (N_324,In_868,In_1153);
and U325 (N_325,In_1018,N_0);
and U326 (N_326,N_67,N_223);
nor U327 (N_327,In_996,In_242);
and U328 (N_328,In_761,In_1310);
or U329 (N_329,In_1172,N_134);
and U330 (N_330,In_197,N_188);
and U331 (N_331,N_35,In_438);
xor U332 (N_332,In_653,In_178);
nand U333 (N_333,In_87,In_1452);
nor U334 (N_334,In_465,In_523);
nand U335 (N_335,In_1328,In_1321);
nand U336 (N_336,N_169,In_1167);
nor U337 (N_337,In_780,In_823);
nand U338 (N_338,In_1188,In_971);
nand U339 (N_339,In_566,In_222);
nor U340 (N_340,In_446,In_332);
xnor U341 (N_341,In_605,In_613);
nand U342 (N_342,In_947,In_131);
nand U343 (N_343,In_1224,N_193);
nand U344 (N_344,In_1044,In_121);
or U345 (N_345,In_428,In_807);
nor U346 (N_346,In_11,In_1132);
xnor U347 (N_347,In_1196,In_296);
or U348 (N_348,In_923,In_1395);
and U349 (N_349,N_117,In_1479);
xor U350 (N_350,In_1100,N_124);
and U351 (N_351,In_561,In_853);
nand U352 (N_352,In_1436,In_751);
or U353 (N_353,In_453,In_549);
or U354 (N_354,N_65,In_354);
nor U355 (N_355,In_873,In_97);
and U356 (N_356,In_673,N_100);
nand U357 (N_357,In_1187,In_272);
and U358 (N_358,N_201,N_136);
xnor U359 (N_359,In_1191,In_1047);
nand U360 (N_360,In_1205,In_1062);
nand U361 (N_361,In_1482,N_78);
nor U362 (N_362,N_190,N_88);
and U363 (N_363,In_591,In_939);
and U364 (N_364,In_450,N_15);
and U365 (N_365,In_1054,N_210);
and U366 (N_366,In_908,In_25);
nand U367 (N_367,N_149,N_60);
and U368 (N_368,In_528,In_1385);
and U369 (N_369,In_234,In_402);
nor U370 (N_370,In_31,N_90);
xnor U371 (N_371,In_567,In_1138);
xor U372 (N_372,In_916,In_479);
nand U373 (N_373,N_218,In_930);
nand U374 (N_374,In_734,In_142);
or U375 (N_375,In_415,N_271);
or U376 (N_376,In_23,In_550);
xnor U377 (N_377,In_416,In_488);
and U378 (N_378,In_1252,In_1176);
xnor U379 (N_379,In_389,N_144);
nand U380 (N_380,In_247,In_92);
and U381 (N_381,In_70,In_1443);
xnor U382 (N_382,In_992,In_341);
and U383 (N_383,In_525,In_600);
xnor U384 (N_384,In_913,In_959);
nor U385 (N_385,N_203,In_860);
and U386 (N_386,In_906,In_315);
and U387 (N_387,N_74,N_32);
and U388 (N_388,In_100,In_737);
and U389 (N_389,In_478,N_183);
xnor U390 (N_390,In_291,In_677);
or U391 (N_391,In_1016,In_299);
or U392 (N_392,In_1202,N_199);
nand U393 (N_393,N_3,N_7);
nor U394 (N_394,In_623,In_1113);
or U395 (N_395,In_1056,N_66);
or U396 (N_396,In_553,In_743);
xor U397 (N_397,In_475,In_631);
and U398 (N_398,In_814,In_865);
nand U399 (N_399,N_185,In_758);
nand U400 (N_400,In_1201,In_953);
nand U401 (N_401,In_1185,N_47);
nor U402 (N_402,N_299,N_236);
xor U403 (N_403,N_125,N_232);
xnor U404 (N_404,In_225,In_1364);
nand U405 (N_405,In_414,In_1009);
or U406 (N_406,In_535,In_1004);
nor U407 (N_407,N_4,In_784);
nor U408 (N_408,In_792,N_9);
or U409 (N_409,N_273,In_395);
or U410 (N_410,In_1430,In_137);
nand U411 (N_411,In_298,In_889);
nand U412 (N_412,In_1369,N_276);
or U413 (N_413,In_554,In_1413);
or U414 (N_414,In_1329,In_1489);
and U415 (N_415,In_664,In_1373);
and U416 (N_416,N_103,In_380);
or U417 (N_417,N_274,In_876);
and U418 (N_418,In_382,In_746);
xor U419 (N_419,In_1302,In_572);
xnor U420 (N_420,In_182,N_163);
xnor U421 (N_421,In_484,In_1271);
and U422 (N_422,In_357,N_79);
nand U423 (N_423,In_1085,N_182);
or U424 (N_424,In_900,In_133);
nand U425 (N_425,In_852,N_95);
xor U426 (N_426,In_1306,In_915);
nand U427 (N_427,In_384,In_26);
xnor U428 (N_428,In_1261,In_831);
nand U429 (N_429,In_997,In_711);
or U430 (N_430,N_114,In_1281);
nand U431 (N_431,In_1280,In_319);
and U432 (N_432,In_704,N_253);
nand U433 (N_433,N_251,In_1459);
nand U434 (N_434,In_1043,In_1216);
nor U435 (N_435,In_618,In_189);
nor U436 (N_436,In_1337,In_509);
nand U437 (N_437,In_1370,N_187);
or U438 (N_438,In_508,N_162);
xnor U439 (N_439,N_52,N_292);
or U440 (N_440,In_1014,In_1150);
xor U441 (N_441,In_166,In_218);
nor U442 (N_442,In_314,In_803);
or U443 (N_443,In_284,N_170);
and U444 (N_444,In_426,In_809);
and U445 (N_445,N_120,In_1061);
nand U446 (N_446,In_1067,N_280);
nor U447 (N_447,In_683,In_747);
nand U448 (N_448,In_492,In_258);
and U449 (N_449,In_1096,N_231);
xnor U450 (N_450,In_408,In_516);
and U451 (N_451,In_1083,N_84);
nand U452 (N_452,In_1351,In_1412);
nor U453 (N_453,In_42,In_173);
or U454 (N_454,In_1063,N_54);
nand U455 (N_455,In_767,N_58);
xnor U456 (N_456,N_106,N_161);
nor U457 (N_457,In_388,N_73);
or U458 (N_458,In_158,In_740);
nor U459 (N_459,In_716,In_851);
and U460 (N_460,In_1024,In_707);
or U461 (N_461,N_186,In_1059);
or U462 (N_462,In_1146,In_145);
nand U463 (N_463,In_536,In_221);
and U464 (N_464,N_171,In_230);
and U465 (N_465,N_36,N_238);
and U466 (N_466,In_383,In_1440);
nor U467 (N_467,In_1380,N_98);
or U468 (N_468,In_1212,In_303);
and U469 (N_469,In_1137,In_660);
or U470 (N_470,In_1407,In_186);
and U471 (N_471,N_43,N_22);
and U472 (N_472,In_1210,In_250);
nor U473 (N_473,N_207,In_744);
or U474 (N_474,In_301,In_793);
or U475 (N_475,In_661,In_1427);
or U476 (N_476,In_1055,N_235);
or U477 (N_477,N_25,N_255);
nor U478 (N_478,N_206,In_806);
nor U479 (N_479,In_321,N_234);
and U480 (N_480,In_1166,N_93);
xor U481 (N_481,N_38,In_776);
and U482 (N_482,In_890,In_210);
nand U483 (N_483,In_251,N_34);
xnor U484 (N_484,In_934,In_278);
xnor U485 (N_485,N_27,In_942);
nand U486 (N_486,In_451,In_861);
or U487 (N_487,In_309,In_393);
nand U488 (N_488,N_243,In_1021);
nor U489 (N_489,N_127,N_222);
or U490 (N_490,In_381,In_1383);
nand U491 (N_491,N_2,N_146);
xnor U492 (N_492,In_280,In_1422);
nor U493 (N_493,In_407,In_64);
nand U494 (N_494,N_16,In_635);
and U495 (N_495,In_373,In_603);
nor U496 (N_496,In_518,N_113);
nand U497 (N_497,In_1447,In_1053);
nand U498 (N_498,In_1335,In_966);
xor U499 (N_499,In_893,In_208);
nor U500 (N_500,In_1211,In_1488);
nand U501 (N_501,N_189,N_5);
and U502 (N_502,In_1464,In_958);
or U503 (N_503,In_124,N_21);
nor U504 (N_504,In_777,In_1282);
nand U505 (N_505,In_1460,N_263);
nand U506 (N_506,N_8,In_770);
or U507 (N_507,In_775,In_568);
and U508 (N_508,N_168,N_220);
nand U509 (N_509,In_1324,N_211);
nand U510 (N_510,N_46,N_63);
nand U511 (N_511,In_1338,In_719);
xor U512 (N_512,N_85,In_511);
or U513 (N_513,In_1257,In_1231);
nor U514 (N_514,In_458,In_1247);
nand U515 (N_515,In_540,In_527);
and U516 (N_516,In_505,In_1276);
and U517 (N_517,N_219,N_229);
xnor U518 (N_518,In_1421,N_41);
and U519 (N_519,N_115,In_467);
nand U520 (N_520,N_293,In_1071);
nand U521 (N_521,In_433,In_201);
nand U522 (N_522,In_293,In_593);
xnor U523 (N_523,In_1105,In_742);
xnor U524 (N_524,In_22,In_1442);
or U525 (N_525,In_56,In_1353);
and U526 (N_526,In_1099,N_230);
nor U527 (N_527,In_270,In_1418);
nor U528 (N_528,In_1204,In_1006);
and U529 (N_529,In_1123,In_294);
and U530 (N_530,In_891,In_196);
nor U531 (N_531,In_410,In_1284);
nor U532 (N_532,In_185,N_99);
nand U533 (N_533,In_127,In_233);
nor U534 (N_534,In_423,N_62);
xnor U535 (N_535,N_87,In_1307);
xnor U536 (N_536,In_1346,In_715);
xnor U537 (N_537,In_1359,In_663);
nor U538 (N_538,N_250,In_1206);
nor U539 (N_539,In_1484,In_602);
xnor U540 (N_540,In_1272,In_1426);
xnor U541 (N_541,In_1190,N_240);
or U542 (N_542,In_1110,In_867);
and U543 (N_543,In_1164,In_12);
nor U544 (N_544,In_1122,N_192);
and U545 (N_545,In_573,In_20);
nand U546 (N_546,In_84,N_265);
nand U547 (N_547,In_77,In_161);
nor U548 (N_548,N_283,In_1391);
nand U549 (N_549,N_143,N_17);
nor U550 (N_550,In_327,In_1045);
nor U551 (N_551,In_1065,In_643);
nand U552 (N_552,In_875,In_1226);
and U553 (N_553,In_1109,In_1381);
nand U554 (N_554,In_347,In_1330);
or U555 (N_555,In_1069,In_534);
and U556 (N_556,In_1017,N_200);
or U557 (N_557,In_685,In_1217);
nand U558 (N_558,In_802,N_44);
xor U559 (N_559,In_376,In_617);
xnor U560 (N_560,N_59,N_142);
nor U561 (N_561,In_1140,In_344);
nand U562 (N_562,In_970,In_703);
nor U563 (N_563,In_1195,In_1033);
or U564 (N_564,In_260,N_155);
or U565 (N_565,In_1129,In_360);
and U566 (N_566,In_542,In_611);
nor U567 (N_567,In_401,N_298);
or U568 (N_568,In_1074,In_546);
or U569 (N_569,In_963,N_279);
and U570 (N_570,In_191,In_1264);
nor U571 (N_571,In_810,In_487);
or U572 (N_572,In_374,In_521);
and U573 (N_573,In_397,N_141);
or U574 (N_574,In_482,N_151);
nand U575 (N_575,In_460,In_1114);
or U576 (N_576,In_1289,In_106);
xnor U577 (N_577,In_1404,N_19);
and U578 (N_578,In_66,In_1239);
nor U579 (N_579,In_249,In_307);
and U580 (N_580,N_51,N_264);
xor U581 (N_581,N_226,In_80);
xnor U582 (N_582,In_7,In_982);
xnor U583 (N_583,N_156,In_472);
nor U584 (N_584,N_277,In_1035);
xnor U585 (N_585,In_538,In_666);
nand U586 (N_586,In_682,N_20);
or U587 (N_587,N_198,In_676);
nand U588 (N_588,In_1312,In_675);
and U589 (N_589,In_363,In_1499);
nand U590 (N_590,In_1431,In_1396);
xor U591 (N_591,In_1141,In_430);
xor U592 (N_592,In_470,In_324);
nor U593 (N_593,In_1316,N_267);
nand U594 (N_594,In_1305,In_925);
or U595 (N_595,In_1174,In_1077);
xor U596 (N_596,In_739,In_1285);
nor U597 (N_597,In_541,In_45);
and U598 (N_598,In_163,In_1162);
nand U599 (N_599,N_40,In_597);
nand U600 (N_600,N_409,N_583);
nor U601 (N_601,N_425,In_529);
and U602 (N_602,In_1342,In_952);
nand U603 (N_603,In_670,N_541);
and U604 (N_604,In_983,N_262);
xnor U605 (N_605,N_550,In_288);
and U606 (N_606,In_469,N_568);
or U607 (N_607,N_112,N_282);
xor U608 (N_608,N_507,N_549);
nor U609 (N_609,N_566,In_216);
or U610 (N_610,N_439,In_1311);
or U611 (N_611,N_594,N_416);
or U612 (N_612,N_407,N_97);
or U613 (N_613,N_420,N_153);
nand U614 (N_614,In_887,N_179);
and U615 (N_615,In_888,N_131);
nand U616 (N_616,In_468,N_152);
and U617 (N_617,N_383,N_391);
nand U618 (N_618,In_648,N_332);
nor U619 (N_619,In_1472,N_348);
and U620 (N_620,In_392,N_428);
or U621 (N_621,In_1339,N_309);
or U622 (N_622,In_1297,In_51);
and U623 (N_623,N_553,In_869);
nand U624 (N_624,In_819,N_64);
and U625 (N_625,N_177,In_1094);
xor U626 (N_626,N_366,In_153);
nor U627 (N_627,N_498,N_272);
and U628 (N_628,N_522,N_509);
and U629 (N_629,N_316,In_1319);
xor U630 (N_630,N_599,In_1420);
and U631 (N_631,In_766,In_1093);
nor U632 (N_632,In_828,N_14);
xor U633 (N_633,In_1493,N_312);
nor U634 (N_634,In_1084,N_39);
nor U635 (N_635,In_769,In_614);
nand U636 (N_636,N_215,In_537);
xor U637 (N_637,In_329,In_577);
nand U638 (N_638,N_321,N_96);
nor U639 (N_639,In_1249,N_576);
and U640 (N_640,In_1327,In_998);
nand U641 (N_641,In_817,N_580);
and U642 (N_642,In_207,In_1241);
and U643 (N_643,N_29,In_300);
xnor U644 (N_644,N_486,In_443);
and U645 (N_645,N_445,N_390);
nand U646 (N_646,In_1317,In_220);
xnor U647 (N_647,N_572,In_946);
and U648 (N_648,In_442,N_429);
and U649 (N_649,N_216,In_1108);
nand U650 (N_650,N_421,In_192);
nor U651 (N_651,N_166,N_543);
and U652 (N_652,In_969,In_65);
nor U653 (N_653,N_132,N_252);
or U654 (N_654,In_78,N_441);
nand U655 (N_655,N_517,N_268);
nand U656 (N_656,In_476,In_1260);
or U657 (N_657,N_577,In_1414);
nand U658 (N_658,N_431,In_881);
and U659 (N_659,In_168,N_315);
or U660 (N_660,In_1486,N_501);
nor U661 (N_661,N_224,In_126);
nor U662 (N_662,In_474,N_465);
nor U663 (N_663,N_322,In_462);
xor U664 (N_664,N_520,N_237);
and U665 (N_665,N_320,N_487);
and U666 (N_666,N_239,N_197);
nand U667 (N_667,In_318,N_380);
xnor U668 (N_668,In_1218,In_302);
xnor U669 (N_669,In_841,In_54);
nand U670 (N_670,In_1437,N_288);
or U671 (N_671,In_919,N_562);
xnor U672 (N_672,N_83,In_1143);
or U673 (N_673,In_926,In_1394);
nand U674 (N_674,N_12,In_310);
nor U675 (N_675,In_459,N_393);
nand U676 (N_676,In_748,N_55);
xnor U677 (N_677,In_1244,In_679);
or U678 (N_678,N_172,In_1019);
and U679 (N_679,In_317,N_138);
or U680 (N_680,N_564,N_281);
xor U681 (N_681,In_844,N_514);
and U682 (N_682,In_840,In_1145);
xor U683 (N_683,In_560,In_1323);
or U684 (N_684,N_524,N_527);
nand U685 (N_685,N_77,N_505);
and U686 (N_686,N_398,N_516);
and U687 (N_687,In_187,In_612);
or U688 (N_688,N_382,In_651);
nand U689 (N_689,In_19,In_749);
or U690 (N_690,N_471,In_420);
nand U691 (N_691,In_1159,N_515);
nand U692 (N_692,N_330,In_105);
xnor U693 (N_693,In_377,N_491);
or U694 (N_694,N_266,N_444);
and U695 (N_695,In_130,In_473);
or U696 (N_696,N_427,In_655);
and U697 (N_697,In_642,In_1242);
and U698 (N_698,N_482,N_310);
and U699 (N_699,N_488,N_569);
xnor U700 (N_700,In_441,N_81);
nand U701 (N_701,N_1,N_291);
or U702 (N_702,In_165,N_404);
nor U703 (N_703,N_457,In_352);
or U704 (N_704,N_337,In_1454);
or U705 (N_705,In_1060,N_45);
or U706 (N_706,In_576,N_184);
or U707 (N_707,N_140,In_822);
xor U708 (N_708,In_773,N_49);
and U709 (N_709,N_378,N_31);
or U710 (N_710,N_408,N_176);
nand U711 (N_711,N_592,In_968);
or U712 (N_712,N_137,In_1283);
or U713 (N_713,N_37,N_414);
nand U714 (N_714,N_69,N_147);
nand U715 (N_715,N_534,In_164);
or U716 (N_716,In_502,N_470);
nand U717 (N_717,N_209,In_1299);
and U718 (N_718,N_275,N_111);
and U719 (N_719,N_508,In_38);
or U720 (N_720,N_212,N_159);
xor U721 (N_721,N_53,N_290);
nor U722 (N_722,In_622,N_402);
and U723 (N_723,In_193,N_308);
or U724 (N_724,N_356,N_443);
xnor U725 (N_725,N_563,In_1169);
and U726 (N_726,N_13,In_1401);
nand U727 (N_727,N_518,In_417);
nand U728 (N_728,In_396,In_304);
or U729 (N_729,N_94,In_1127);
nand U730 (N_730,N_573,N_537);
nand U731 (N_731,In_223,In_579);
and U732 (N_732,N_175,N_379);
and U733 (N_733,In_731,N_381);
nor U734 (N_734,N_319,In_477);
or U735 (N_735,In_156,N_389);
nor U736 (N_736,N_349,N_284);
nand U737 (N_737,N_295,N_297);
nand U738 (N_738,In_1345,N_551);
or U739 (N_739,N_546,N_476);
xor U740 (N_740,N_181,N_375);
nor U741 (N_741,In_1333,In_123);
nor U742 (N_742,N_123,In_241);
xor U743 (N_743,N_305,In_1357);
and U744 (N_744,N_475,In_1294);
nor U745 (N_745,N_289,N_302);
and U746 (N_746,In_1170,In_1462);
nand U747 (N_747,N_108,N_467);
and U748 (N_748,N_318,In_466);
and U749 (N_749,In_1012,In_783);
nand U750 (N_750,In_931,N_535);
xor U751 (N_751,In_74,N_560);
xor U752 (N_752,In_795,In_500);
or U753 (N_753,In_1228,N_68);
and U754 (N_754,In_825,In_497);
and U755 (N_755,In_595,N_242);
and U756 (N_756,N_70,N_254);
or U757 (N_757,N_430,N_437);
and U758 (N_758,In_1154,N_285);
or U759 (N_759,In_1371,N_101);
nand U760 (N_760,In_659,N_269);
nor U761 (N_761,In_486,In_1011);
nand U762 (N_762,In_759,N_529);
nor U763 (N_763,N_202,N_484);
nand U764 (N_764,N_257,In_833);
nor U765 (N_765,In_259,In_801);
or U766 (N_766,In_1445,N_403);
or U767 (N_767,In_206,N_459);
and U768 (N_768,N_278,N_582);
nand U769 (N_769,N_413,In_1182);
nor U770 (N_770,N_557,In_246);
xnor U771 (N_771,In_976,In_1250);
and U772 (N_772,In_256,In_753);
xnor U773 (N_773,In_738,N_586);
or U774 (N_774,N_48,In_641);
nand U775 (N_775,In_863,In_311);
nand U776 (N_776,N_385,N_353);
or U777 (N_777,In_1193,N_419);
nand U778 (N_778,In_562,In_170);
xnor U779 (N_779,N_424,In_874);
nand U780 (N_780,N_453,In_551);
nand U781 (N_781,N_555,In_1399);
and U782 (N_782,N_167,N_331);
nor U783 (N_783,N_545,N_584);
xnor U784 (N_784,N_208,N_513);
nor U785 (N_785,N_345,N_540);
nor U786 (N_786,N_245,In_94);
nand U787 (N_787,N_139,In_273);
xnor U788 (N_788,In_559,In_439);
nand U789 (N_789,In_578,N_227);
nand U790 (N_790,In_557,In_894);
xnor U791 (N_791,In_205,N_334);
and U792 (N_792,N_479,N_360);
nor U793 (N_793,N_89,N_359);
or U794 (N_794,N_128,In_1039);
nand U795 (N_795,N_596,In_1292);
or U796 (N_796,N_423,N_489);
nor U797 (N_797,N_347,In_877);
xnor U798 (N_798,N_493,N_104);
or U799 (N_799,In_1409,N_75);
xor U800 (N_800,In_452,In_1225);
and U801 (N_801,In_1155,N_384);
and U802 (N_802,In_435,N_300);
or U803 (N_803,N_502,In_114);
xnor U804 (N_804,N_412,In_1403);
and U805 (N_805,N_474,In_1433);
and U806 (N_806,In_496,In_608);
and U807 (N_807,N_335,In_1268);
or U808 (N_808,N_145,N_119);
or U809 (N_809,N_511,In_27);
or U810 (N_810,N_157,In_398);
and U811 (N_811,In_118,In_978);
and U812 (N_812,N_561,N_129);
nor U813 (N_813,In_385,N_248);
and U814 (N_814,In_1367,In_1275);
nor U815 (N_815,N_503,In_898);
xor U816 (N_816,In_333,In_1136);
and U817 (N_817,In_723,In_714);
nor U818 (N_818,N_461,In_514);
nor U819 (N_819,In_16,In_1298);
xnor U820 (N_820,In_1485,N_196);
nand U821 (N_821,N_542,In_322);
or U822 (N_822,In_269,In_797);
xnor U823 (N_823,In_167,In_1251);
or U824 (N_824,In_93,In_1410);
nor U825 (N_825,N_130,In_1125);
nand U826 (N_826,In_129,In_1066);
or U827 (N_827,N_354,N_458);
xor U828 (N_828,N_570,In_305);
or U829 (N_829,N_178,In_449);
nand U830 (N_830,N_61,In_994);
nand U831 (N_831,N_116,N_102);
or U832 (N_832,In_912,In_570);
nand U833 (N_833,In_684,In_1497);
nor U834 (N_834,In_1,In_940);
or U835 (N_835,In_646,N_344);
xnor U836 (N_836,In_444,In_98);
xor U837 (N_837,In_228,In_1213);
or U838 (N_838,In_859,In_1466);
nand U839 (N_839,In_140,In_171);
nor U840 (N_840,N_261,In_1161);
nor U841 (N_841,In_281,In_1117);
nand U842 (N_842,N_126,In_180);
nand U843 (N_843,N_536,N_490);
or U844 (N_844,In_512,In_47);
or U845 (N_845,In_503,In_681);
nor U846 (N_846,In_1450,N_164);
nor U847 (N_847,In_582,N_418);
nor U848 (N_848,N_247,N_221);
or U849 (N_849,N_371,N_339);
nand U850 (N_850,In_480,In_977);
and U851 (N_851,In_312,N_519);
and U852 (N_852,In_277,N_213);
and U853 (N_853,N_395,N_500);
nor U854 (N_854,In_1274,In_1208);
or U855 (N_855,In_1121,N_10);
or U856 (N_856,N_352,In_37);
xor U857 (N_857,In_533,N_422);
or U858 (N_858,In_387,In_1390);
nand U859 (N_859,In_107,In_702);
nand U860 (N_860,N_448,N_478);
or U861 (N_861,N_483,In_975);
nor U862 (N_862,In_815,N_531);
nand U863 (N_863,N_118,N_370);
nand U864 (N_864,In_1392,N_496);
nor U865 (N_865,N_228,In_510);
nand U866 (N_866,N_342,In_1473);
nand U867 (N_867,N_341,N_523);
and U868 (N_868,N_258,In_539);
and U869 (N_869,In_146,N_333);
nor U870 (N_870,In_896,In_13);
nand U871 (N_871,N_450,In_117);
or U872 (N_872,N_376,N_436);
xnor U873 (N_873,In_1245,N_91);
and U874 (N_874,In_1233,In_419);
xor U875 (N_875,In_1232,In_872);
or U876 (N_876,N_386,N_526);
nor U877 (N_877,In_805,In_83);
and U878 (N_878,In_1495,In_658);
and U879 (N_879,N_304,In_1175);
and U880 (N_880,In_789,In_811);
xnor U881 (N_881,In_1341,In_498);
nor U882 (N_882,In_1134,N_154);
nor U883 (N_883,N_174,N_548);
nand U884 (N_884,N_477,N_544);
and U885 (N_885,In_736,N_559);
nand U886 (N_886,In_176,N_241);
and U887 (N_887,N_521,N_435);
xor U888 (N_888,In_563,N_447);
nand U889 (N_889,In_1007,In_886);
and U890 (N_890,In_331,N_397);
xnor U891 (N_891,N_121,In_455);
nand U892 (N_892,In_904,In_427);
xor U893 (N_893,N_538,In_520);
or U894 (N_894,In_69,In_29);
xor U895 (N_895,N_579,N_259);
nor U896 (N_896,N_510,N_480);
or U897 (N_897,N_442,In_375);
or U898 (N_898,In_974,N_307);
nand U899 (N_899,In_1032,In_226);
xnor U900 (N_900,In_1144,N_460);
xnor U901 (N_901,N_173,N_721);
and U902 (N_902,In_799,N_369);
or U903 (N_903,N_575,N_400);
and U904 (N_904,N_672,N_636);
and U905 (N_905,N_801,In_1028);
nand U906 (N_906,N_837,In_1238);
xor U907 (N_907,N_694,N_287);
nor U908 (N_908,In_657,In_326);
nor U909 (N_909,N_367,In_115);
nand U910 (N_910,N_891,N_653);
nor U911 (N_911,N_691,In_409);
and U912 (N_912,N_667,N_711);
nor U913 (N_913,N_451,In_1468);
or U914 (N_914,N_775,N_740);
and U915 (N_915,N_757,N_314);
or U916 (N_916,N_865,N_639);
xnor U917 (N_917,N_754,N_411);
xnor U918 (N_918,N_899,N_578);
xor U919 (N_919,In_471,N_768);
nor U920 (N_920,N_606,In_257);
nor U921 (N_921,N_804,N_456);
nor U922 (N_922,N_313,In_143);
nand U923 (N_923,In_454,N_660);
nor U924 (N_924,N_363,N_699);
xor U925 (N_925,N_633,N_664);
nor U926 (N_926,In_1184,N_871);
xnor U927 (N_927,N_434,N_652);
xor U928 (N_928,In_1375,N_530);
nor U929 (N_929,N_859,In_921);
or U930 (N_930,N_631,N_848);
xnor U931 (N_931,N_759,N_782);
and U932 (N_932,N_643,N_574);
or U933 (N_933,In_1262,N_632);
nor U934 (N_934,N_685,N_687);
and U935 (N_935,N_627,N_260);
and U936 (N_936,In_88,N_387);
and U937 (N_937,N_849,N_830);
and U938 (N_938,N_670,In_183);
or U939 (N_939,In_81,In_558);
nand U940 (N_940,N_286,N_876);
and U941 (N_941,N_760,In_1103);
and U942 (N_942,N_786,N_294);
xnor U943 (N_943,N_492,N_705);
nand U944 (N_944,In_1200,In_144);
xnor U945 (N_945,N_351,N_817);
and U946 (N_946,N_713,N_788);
nor U947 (N_947,In_5,N_887);
and U948 (N_948,N_373,N_191);
xnor U949 (N_949,In_1149,In_1465);
or U950 (N_950,N_755,N_326);
and U951 (N_951,N_868,N_343);
nor U952 (N_952,In_112,N_76);
nor U953 (N_953,N_853,N_214);
xor U954 (N_954,In_911,N_884);
or U955 (N_955,N_802,N_765);
xnor U956 (N_956,N_620,In_772);
nand U957 (N_957,In_368,N_861);
nor U958 (N_958,N_256,N_787);
or U959 (N_959,N_468,In_695);
or U960 (N_960,In_1469,N_635);
or U961 (N_961,N_655,N_372);
and U962 (N_962,N_649,N_898);
xnor U963 (N_963,N_693,N_827);
xor U964 (N_964,N_640,N_807);
and U965 (N_965,N_764,N_738);
nor U966 (N_966,N_452,N_658);
or U967 (N_967,N_410,N_624);
nand U968 (N_968,N_11,N_626);
xnor U969 (N_969,N_692,In_1382);
nor U970 (N_970,N_661,N_158);
nor U971 (N_971,In_821,N_790);
and U972 (N_972,N_821,N_109);
xor U973 (N_973,N_834,In_355);
and U974 (N_974,N_824,N_616);
nand U975 (N_975,In_1168,N_350);
xor U976 (N_976,N_645,N_303);
nor U977 (N_977,In_762,In_949);
nand U978 (N_978,N_50,N_604);
nand U979 (N_979,N_225,N_438);
or U980 (N_980,N_246,N_777);
or U981 (N_981,N_602,N_862);
or U982 (N_982,In_1354,N_831);
xnor U983 (N_983,In_125,In_336);
and U984 (N_984,In_826,In_86);
or U985 (N_985,N_832,N_107);
xor U986 (N_986,N_638,In_837);
nor U987 (N_987,In_434,N_712);
nand U988 (N_988,In_198,N_682);
nand U989 (N_989,N_897,N_622);
and U990 (N_990,N_684,In_15);
nand U991 (N_991,N_761,N_499);
or U992 (N_992,N_204,In_36);
xor U993 (N_993,N_481,N_399);
nand U994 (N_994,N_895,N_892);
xor U995 (N_995,In_755,N_882);
nor U996 (N_996,N_472,N_24);
nor U997 (N_997,N_889,N_717);
nor U998 (N_998,N_135,In_804);
xor U999 (N_999,N_737,N_648);
or U1000 (N_1000,N_567,N_819);
and U1001 (N_1001,N_585,In_945);
or U1002 (N_1002,N_893,N_133);
nand U1003 (N_1003,N_615,In_102);
or U1004 (N_1004,N_742,N_763);
or U1005 (N_1005,N_748,N_57);
and U1006 (N_1006,N_440,N_883);
or U1007 (N_1007,N_735,N_838);
or U1008 (N_1008,In_1444,N_880);
xnor U1009 (N_1009,N_532,N_33);
or U1010 (N_1010,N_317,In_63);
nand U1011 (N_1011,N_866,N_329);
or U1012 (N_1012,N_847,N_533);
or U1013 (N_1013,N_785,In_1008);
nor U1014 (N_1014,N_659,N_603);
or U1015 (N_1015,N_677,N_396);
nor U1016 (N_1016,In_1439,N_811);
xor U1017 (N_1017,N_357,N_803);
and U1018 (N_1018,N_607,N_644);
nor U1019 (N_1019,N_650,In_219);
nand U1020 (N_1020,N_854,N_205);
xnor U1021 (N_1021,N_815,N_504);
xor U1022 (N_1022,N_249,N_829);
nor U1023 (N_1023,N_844,In_362);
or U1024 (N_1024,N_466,N_818);
xnor U1025 (N_1025,N_695,N_703);
or U1026 (N_1026,N_361,N_628);
xor U1027 (N_1027,N_728,In_708);
xnor U1028 (N_1028,N_417,N_752);
xor U1029 (N_1029,N_816,In_177);
and U1030 (N_1030,N_799,N_629);
and U1031 (N_1031,In_1222,N_855);
nand U1032 (N_1032,N_797,N_873);
nand U1033 (N_1033,N_610,N_870);
xor U1034 (N_1034,N_311,N_528);
or U1035 (N_1035,N_30,N_556);
nor U1036 (N_1036,N_630,N_651);
nor U1037 (N_1037,In_827,N_836);
nand U1038 (N_1038,N_724,N_619);
or U1039 (N_1039,N_497,N_462);
or U1040 (N_1040,N_825,In_732);
nor U1041 (N_1041,N_405,In_1180);
xor U1042 (N_1042,N_747,N_368);
or U1043 (N_1043,N_780,In_162);
nor U1044 (N_1044,N_751,N_726);
xor U1045 (N_1045,N_863,N_609);
nand U1046 (N_1046,N_364,N_762);
xor U1047 (N_1047,N_858,In_1111);
xor U1048 (N_1048,N_841,N_690);
nor U1049 (N_1049,N_796,In_609);
nor U1050 (N_1050,In_1349,N_750);
nor U1051 (N_1051,N_820,N_706);
xor U1052 (N_1052,N_587,N_828);
and U1053 (N_1053,N_707,N_666);
and U1054 (N_1054,N_554,N_793);
nor U1055 (N_1055,N_449,N_42);
or U1056 (N_1056,N_822,N_669);
nand U1057 (N_1057,N_617,N_657);
xor U1058 (N_1058,In_44,N_365);
nor U1059 (N_1059,N_646,N_723);
and U1060 (N_1060,N_845,N_180);
and U1061 (N_1061,N_595,N_150);
and U1062 (N_1062,N_446,In_1320);
nor U1063 (N_1063,N_700,N_769);
and U1064 (N_1064,In_425,N_784);
xor U1065 (N_1065,In_1023,In_1092);
nand U1066 (N_1066,In_1116,N_71);
xnor U1067 (N_1067,N_686,N_336);
nand U1068 (N_1068,In_48,In_1343);
nand U1069 (N_1069,In_1308,In_1492);
xnor U1070 (N_1070,N_464,N_864);
or U1071 (N_1071,N_814,N_857);
nor U1072 (N_1072,In_985,N_377);
and U1073 (N_1073,N_709,N_598);
xnor U1074 (N_1074,N_28,N_770);
xnor U1075 (N_1075,N_730,In_181);
and U1076 (N_1076,N_597,In_349);
xnor U1077 (N_1077,In_754,N_743);
xor U1078 (N_1078,N_890,N_744);
nand U1079 (N_1079,N_772,In_794);
and U1080 (N_1080,N_673,N_338);
nand U1081 (N_1081,N_697,N_346);
and U1082 (N_1082,N_774,N_601);
or U1083 (N_1083,N_731,N_839);
xnor U1084 (N_1084,N_702,N_328);
nand U1085 (N_1085,N_565,N_809);
nand U1086 (N_1086,In_531,N_374);
and U1087 (N_1087,N_794,N_856);
nor U1088 (N_1088,N_506,N_850);
nor U1089 (N_1089,N_781,N_806);
or U1090 (N_1090,N_148,In_151);
nand U1091 (N_1091,N_525,In_552);
and U1092 (N_1092,N_618,In_263);
xnor U1093 (N_1093,In_1398,N_625);
xnor U1094 (N_1094,N_415,N_881);
nand U1095 (N_1095,N_810,N_872);
nor U1096 (N_1096,N_792,N_725);
nor U1097 (N_1097,N_647,N_846);
and U1098 (N_1098,N_433,N_122);
nand U1099 (N_1099,In_96,N_18);
xnor U1100 (N_1100,N_852,N_86);
nand U1101 (N_1101,In_720,In_771);
or U1102 (N_1102,N_401,N_722);
or U1103 (N_1103,N_869,N_662);
or U1104 (N_1104,N_621,In_545);
and U1105 (N_1105,N_512,N_879);
nand U1106 (N_1106,N_296,N_874);
and U1107 (N_1107,N_195,N_270);
or U1108 (N_1108,N_432,N_813);
and U1109 (N_1109,N_591,N_698);
nand U1110 (N_1110,N_160,N_668);
or U1111 (N_1111,N_704,N_681);
nand U1112 (N_1112,N_745,N_325);
xnor U1113 (N_1113,N_495,N_732);
and U1114 (N_1114,In_267,N_323);
and U1115 (N_1115,In_649,N_355);
and U1116 (N_1116,N_588,N_720);
xor U1117 (N_1117,In_938,N_710);
xor U1118 (N_1118,N_696,N_689);
nand U1119 (N_1119,N_741,In_788);
or U1120 (N_1120,N_678,In_1147);
xor U1121 (N_1121,N_388,N_608);
xnor U1122 (N_1122,N_547,N_539);
nor U1123 (N_1123,N_105,N_485);
nand U1124 (N_1124,N_826,In_752);
or U1125 (N_1125,In_1456,In_405);
nand U1126 (N_1126,N_558,N_80);
xnor U1127 (N_1127,N_642,N_463);
and U1128 (N_1128,N_674,In_149);
nand U1129 (N_1129,In_1068,N_860);
and U1130 (N_1130,N_843,N_842);
and U1131 (N_1131,N_552,In_628);
and U1132 (N_1132,In_1034,N_823);
xor U1133 (N_1133,N_878,In_157);
nand U1134 (N_1134,N_894,In_726);
and U1135 (N_1135,N_800,N_778);
nor U1136 (N_1136,N_805,In_1119);
and U1137 (N_1137,N_885,N_634);
nor U1138 (N_1138,N_701,N_888);
nor U1139 (N_1139,N_455,N_593);
and U1140 (N_1140,In_599,N_875);
nor U1141 (N_1141,N_454,N_611);
nand U1142 (N_1142,N_473,In_1036);
or U1143 (N_1143,N_733,N_896);
nand U1144 (N_1144,N_766,N_773);
and U1145 (N_1145,N_165,N_571);
nor U1146 (N_1146,N_654,In_339);
nor U1147 (N_1147,N_362,N_756);
and U1148 (N_1148,N_749,N_739);
and U1149 (N_1149,N_729,N_718);
nor U1150 (N_1150,In_483,In_1236);
xnor U1151 (N_1151,In_713,N_808);
and U1152 (N_1152,N_688,N_771);
and U1153 (N_1153,N_840,N_589);
and U1154 (N_1154,N_758,N_394);
nand U1155 (N_1155,N_680,In_490);
nand U1156 (N_1156,N_392,N_665);
nand U1157 (N_1157,In_90,N_641);
nor U1158 (N_1158,In_345,In_399);
xnor U1159 (N_1159,N_734,In_956);
nand U1160 (N_1160,In_59,N_727);
and U1161 (N_1161,N_469,In_909);
nand U1162 (N_1162,N_791,N_358);
and U1163 (N_1163,N_306,N_776);
nand U1164 (N_1164,N_406,N_789);
nand U1165 (N_1165,N_851,N_746);
and U1166 (N_1166,In_1458,In_9);
and U1167 (N_1167,In_1379,N_877);
and U1168 (N_1168,N_327,N_426);
nand U1169 (N_1169,N_612,N_605);
nand U1170 (N_1170,N_217,In_1332);
nor U1171 (N_1171,N_716,N_812);
xor U1172 (N_1172,N_637,In_120);
xor U1173 (N_1173,In_1432,N_798);
nor U1174 (N_1174,In_629,In_847);
nand U1175 (N_1175,N_867,N_581);
nand U1176 (N_1176,N_714,N_715);
and U1177 (N_1177,In_1471,N_663);
nor U1178 (N_1178,N_795,In_1449);
or U1179 (N_1179,N_767,N_833);
xor U1180 (N_1180,N_736,In_358);
and U1181 (N_1181,In_957,N_623);
nor U1182 (N_1182,N_494,In_750);
nor U1183 (N_1183,In_1448,N_590);
nand U1184 (N_1184,N_708,N_835);
xnor U1185 (N_1185,In_1030,N_719);
and U1186 (N_1186,In_1408,N_679);
nand U1187 (N_1187,N_656,N_671);
xnor U1188 (N_1188,N_82,N_886);
nand U1189 (N_1189,In_1158,In_902);
and U1190 (N_1190,In_138,N_614);
xnor U1191 (N_1191,N_233,N_676);
nor U1192 (N_1192,In_4,N_613);
or U1193 (N_1193,N_600,N_340);
xor U1194 (N_1194,In_903,In_905);
nand U1195 (N_1195,N_753,In_813);
and U1196 (N_1196,N_779,In_513);
nand U1197 (N_1197,N_783,N_683);
nand U1198 (N_1198,N_675,N_23);
nand U1199 (N_1199,N_324,N_301);
nor U1200 (N_1200,N_1047,N_1184);
nand U1201 (N_1201,N_948,N_1060);
xor U1202 (N_1202,N_1157,N_918);
or U1203 (N_1203,N_1191,N_911);
nand U1204 (N_1204,N_1038,N_1099);
nor U1205 (N_1205,N_1061,N_1092);
nand U1206 (N_1206,N_945,N_917);
nor U1207 (N_1207,N_1050,N_1023);
or U1208 (N_1208,N_1154,N_1105);
xor U1209 (N_1209,N_927,N_951);
or U1210 (N_1210,N_1056,N_940);
and U1211 (N_1211,N_1034,N_904);
and U1212 (N_1212,N_925,N_1111);
or U1213 (N_1213,N_1027,N_961);
nor U1214 (N_1214,N_1019,N_1101);
nor U1215 (N_1215,N_983,N_1146);
xor U1216 (N_1216,N_1195,N_992);
xnor U1217 (N_1217,N_1002,N_1073);
or U1218 (N_1218,N_1076,N_1074);
nor U1219 (N_1219,N_1030,N_1045);
nor U1220 (N_1220,N_1199,N_1125);
or U1221 (N_1221,N_1057,N_1156);
or U1222 (N_1222,N_1140,N_909);
nor U1223 (N_1223,N_1014,N_1024);
nor U1224 (N_1224,N_1121,N_908);
nand U1225 (N_1225,N_965,N_907);
nor U1226 (N_1226,N_1150,N_1033);
nand U1227 (N_1227,N_1133,N_1013);
nand U1228 (N_1228,N_901,N_968);
xnor U1229 (N_1229,N_973,N_954);
or U1230 (N_1230,N_1107,N_1194);
or U1231 (N_1231,N_1127,N_929);
xnor U1232 (N_1232,N_1123,N_1085);
nand U1233 (N_1233,N_1134,N_1097);
or U1234 (N_1234,N_994,N_1011);
xor U1235 (N_1235,N_1167,N_919);
or U1236 (N_1236,N_905,N_978);
and U1237 (N_1237,N_1041,N_1058);
xnor U1238 (N_1238,N_1178,N_1122);
xnor U1239 (N_1239,N_1098,N_1071);
xnor U1240 (N_1240,N_949,N_1175);
nand U1241 (N_1241,N_963,N_1080);
nor U1242 (N_1242,N_1119,N_1020);
and U1243 (N_1243,N_970,N_1114);
or U1244 (N_1244,N_1035,N_962);
and U1245 (N_1245,N_971,N_1177);
and U1246 (N_1246,N_969,N_1006);
nor U1247 (N_1247,N_1088,N_958);
nor U1248 (N_1248,N_1001,N_935);
and U1249 (N_1249,N_947,N_1144);
and U1250 (N_1250,N_975,N_984);
nor U1251 (N_1251,N_1046,N_943);
nand U1252 (N_1252,N_1043,N_1064);
and U1253 (N_1253,N_1168,N_1093);
and U1254 (N_1254,N_1077,N_955);
nand U1255 (N_1255,N_1160,N_979);
and U1256 (N_1256,N_923,N_900);
and U1257 (N_1257,N_1100,N_1003);
nor U1258 (N_1258,N_956,N_912);
nand U1259 (N_1259,N_1120,N_1179);
nor U1260 (N_1260,N_1089,N_930);
and U1261 (N_1261,N_1075,N_1065);
or U1262 (N_1262,N_1062,N_1172);
or U1263 (N_1263,N_1174,N_1040);
or U1264 (N_1264,N_1136,N_1083);
xnor U1265 (N_1265,N_991,N_1108);
and U1266 (N_1266,N_922,N_967);
nor U1267 (N_1267,N_1182,N_1082);
or U1268 (N_1268,N_1012,N_1055);
nor U1269 (N_1269,N_1037,N_1022);
nand U1270 (N_1270,N_937,N_997);
and U1271 (N_1271,N_946,N_1192);
nand U1272 (N_1272,N_942,N_1053);
nor U1273 (N_1273,N_1059,N_1078);
nor U1274 (N_1274,N_913,N_1084);
nand U1275 (N_1275,N_1106,N_1044);
nand U1276 (N_1276,N_931,N_985);
xor U1277 (N_1277,N_1010,N_1126);
nor U1278 (N_1278,N_906,N_939);
or U1279 (N_1279,N_1096,N_974);
and U1280 (N_1280,N_1132,N_1015);
xnor U1281 (N_1281,N_1124,N_987);
nor U1282 (N_1282,N_1066,N_1070);
nor U1283 (N_1283,N_1000,N_933);
and U1284 (N_1284,N_1028,N_1161);
nand U1285 (N_1285,N_938,N_1137);
xnor U1286 (N_1286,N_1159,N_1051);
xnor U1287 (N_1287,N_1104,N_1189);
nor U1288 (N_1288,N_1063,N_1094);
nand U1289 (N_1289,N_1095,N_1118);
xnor U1290 (N_1290,N_1004,N_1026);
or U1291 (N_1291,N_1052,N_1117);
and U1292 (N_1292,N_902,N_1171);
or U1293 (N_1293,N_1102,N_950);
nand U1294 (N_1294,N_1173,N_976);
xnor U1295 (N_1295,N_1185,N_1018);
nand U1296 (N_1296,N_1016,N_1183);
or U1297 (N_1297,N_964,N_1151);
or U1298 (N_1298,N_966,N_1109);
xor U1299 (N_1299,N_1090,N_903);
and U1300 (N_1300,N_996,N_1176);
or U1301 (N_1301,N_957,N_1143);
nor U1302 (N_1302,N_988,N_1112);
nor U1303 (N_1303,N_1079,N_1032);
and U1304 (N_1304,N_993,N_1007);
or U1305 (N_1305,N_921,N_986);
nand U1306 (N_1306,N_1181,N_1153);
xor U1307 (N_1307,N_1054,N_915);
or U1308 (N_1308,N_999,N_936);
xor U1309 (N_1309,N_914,N_1113);
xnor U1310 (N_1310,N_1039,N_1067);
xnor U1311 (N_1311,N_953,N_1196);
xnor U1312 (N_1312,N_952,N_1188);
nor U1313 (N_1313,N_1009,N_1198);
nor U1314 (N_1314,N_1091,N_1029);
or U1315 (N_1315,N_916,N_1021);
nand U1316 (N_1316,N_941,N_920);
xnor U1317 (N_1317,N_1148,N_1141);
xnor U1318 (N_1318,N_926,N_998);
nand U1319 (N_1319,N_1048,N_1036);
nand U1320 (N_1320,N_910,N_981);
nand U1321 (N_1321,N_1025,N_1031);
nor U1322 (N_1322,N_980,N_972);
and U1323 (N_1323,N_1081,N_1186);
and U1324 (N_1324,N_1110,N_1138);
and U1325 (N_1325,N_1042,N_934);
and U1326 (N_1326,N_1152,N_1164);
nand U1327 (N_1327,N_1139,N_995);
or U1328 (N_1328,N_1086,N_1149);
xor U1329 (N_1329,N_928,N_1072);
or U1330 (N_1330,N_924,N_944);
nand U1331 (N_1331,N_1103,N_1163);
xor U1332 (N_1332,N_1135,N_1170);
and U1333 (N_1333,N_1008,N_1131);
and U1334 (N_1334,N_1180,N_989);
xor U1335 (N_1335,N_1128,N_1169);
nor U1336 (N_1336,N_1162,N_977);
or U1337 (N_1337,N_1087,N_1142);
or U1338 (N_1338,N_1187,N_1068);
nand U1339 (N_1339,N_1005,N_959);
xnor U1340 (N_1340,N_1193,N_1069);
nand U1341 (N_1341,N_960,N_1197);
nand U1342 (N_1342,N_1116,N_1049);
xnor U1343 (N_1343,N_1165,N_990);
nand U1344 (N_1344,N_1129,N_1115);
nand U1345 (N_1345,N_1190,N_1158);
xnor U1346 (N_1346,N_1145,N_1017);
or U1347 (N_1347,N_1166,N_932);
and U1348 (N_1348,N_1155,N_1130);
or U1349 (N_1349,N_1147,N_982);
nor U1350 (N_1350,N_918,N_1071);
xnor U1351 (N_1351,N_1014,N_1175);
xnor U1352 (N_1352,N_1063,N_1124);
nand U1353 (N_1353,N_927,N_1061);
nor U1354 (N_1354,N_1070,N_1083);
nor U1355 (N_1355,N_1091,N_1044);
nand U1356 (N_1356,N_964,N_912);
xnor U1357 (N_1357,N_911,N_960);
xor U1358 (N_1358,N_1144,N_1006);
xnor U1359 (N_1359,N_1009,N_991);
nand U1360 (N_1360,N_989,N_1126);
and U1361 (N_1361,N_997,N_900);
nand U1362 (N_1362,N_1033,N_1120);
and U1363 (N_1363,N_927,N_1069);
nand U1364 (N_1364,N_1152,N_1088);
and U1365 (N_1365,N_952,N_1085);
xor U1366 (N_1366,N_1022,N_1006);
and U1367 (N_1367,N_1097,N_1176);
or U1368 (N_1368,N_969,N_1096);
or U1369 (N_1369,N_984,N_1149);
or U1370 (N_1370,N_1033,N_919);
nand U1371 (N_1371,N_1184,N_1155);
nand U1372 (N_1372,N_1076,N_1182);
nand U1373 (N_1373,N_987,N_1175);
xnor U1374 (N_1374,N_1019,N_1023);
nor U1375 (N_1375,N_1113,N_994);
nand U1376 (N_1376,N_1093,N_925);
and U1377 (N_1377,N_946,N_1012);
nand U1378 (N_1378,N_904,N_1097);
nor U1379 (N_1379,N_1010,N_1174);
nor U1380 (N_1380,N_964,N_958);
nand U1381 (N_1381,N_1199,N_1030);
nand U1382 (N_1382,N_931,N_998);
nor U1383 (N_1383,N_1198,N_976);
nand U1384 (N_1384,N_1119,N_1127);
nand U1385 (N_1385,N_1171,N_1115);
nor U1386 (N_1386,N_1133,N_1032);
xor U1387 (N_1387,N_1197,N_964);
nor U1388 (N_1388,N_974,N_944);
xor U1389 (N_1389,N_909,N_1100);
nand U1390 (N_1390,N_1140,N_1151);
nor U1391 (N_1391,N_966,N_1102);
nor U1392 (N_1392,N_1009,N_980);
xor U1393 (N_1393,N_900,N_926);
nand U1394 (N_1394,N_1176,N_963);
nor U1395 (N_1395,N_1039,N_1192);
and U1396 (N_1396,N_1014,N_937);
nand U1397 (N_1397,N_1158,N_1053);
nor U1398 (N_1398,N_1183,N_952);
or U1399 (N_1399,N_961,N_1095);
nor U1400 (N_1400,N_940,N_1140);
xnor U1401 (N_1401,N_1079,N_962);
nor U1402 (N_1402,N_1113,N_1177);
nor U1403 (N_1403,N_1034,N_945);
nand U1404 (N_1404,N_1162,N_1054);
xor U1405 (N_1405,N_1030,N_1082);
and U1406 (N_1406,N_995,N_1186);
and U1407 (N_1407,N_1069,N_1050);
xor U1408 (N_1408,N_1175,N_1194);
nor U1409 (N_1409,N_902,N_1063);
and U1410 (N_1410,N_1033,N_945);
xor U1411 (N_1411,N_1020,N_1091);
or U1412 (N_1412,N_1166,N_1141);
and U1413 (N_1413,N_998,N_1035);
and U1414 (N_1414,N_997,N_979);
or U1415 (N_1415,N_1011,N_1147);
nand U1416 (N_1416,N_1116,N_1100);
xnor U1417 (N_1417,N_1058,N_1042);
nor U1418 (N_1418,N_977,N_946);
nand U1419 (N_1419,N_980,N_1137);
or U1420 (N_1420,N_958,N_1139);
nand U1421 (N_1421,N_1162,N_1186);
xnor U1422 (N_1422,N_1057,N_989);
nor U1423 (N_1423,N_1119,N_1038);
and U1424 (N_1424,N_943,N_975);
nor U1425 (N_1425,N_976,N_921);
or U1426 (N_1426,N_1122,N_1039);
and U1427 (N_1427,N_1038,N_1036);
and U1428 (N_1428,N_1189,N_1139);
nand U1429 (N_1429,N_975,N_1018);
or U1430 (N_1430,N_1018,N_1039);
nor U1431 (N_1431,N_1169,N_1172);
and U1432 (N_1432,N_959,N_1115);
nand U1433 (N_1433,N_1073,N_1067);
and U1434 (N_1434,N_1023,N_1082);
nand U1435 (N_1435,N_939,N_928);
nor U1436 (N_1436,N_1006,N_1111);
nor U1437 (N_1437,N_967,N_1069);
nand U1438 (N_1438,N_913,N_1169);
and U1439 (N_1439,N_988,N_1050);
or U1440 (N_1440,N_1097,N_1130);
or U1441 (N_1441,N_966,N_1196);
nand U1442 (N_1442,N_1063,N_967);
xor U1443 (N_1443,N_1088,N_1096);
xor U1444 (N_1444,N_1139,N_928);
xor U1445 (N_1445,N_1054,N_1038);
or U1446 (N_1446,N_961,N_1141);
and U1447 (N_1447,N_1056,N_1110);
nand U1448 (N_1448,N_1068,N_1005);
xor U1449 (N_1449,N_1107,N_1151);
xnor U1450 (N_1450,N_1192,N_994);
nor U1451 (N_1451,N_1121,N_1113);
and U1452 (N_1452,N_935,N_1186);
or U1453 (N_1453,N_1052,N_914);
xor U1454 (N_1454,N_1018,N_1074);
nand U1455 (N_1455,N_1109,N_1140);
and U1456 (N_1456,N_1154,N_1027);
xor U1457 (N_1457,N_1173,N_1078);
and U1458 (N_1458,N_1182,N_1117);
or U1459 (N_1459,N_943,N_935);
nand U1460 (N_1460,N_1045,N_913);
or U1461 (N_1461,N_931,N_901);
nand U1462 (N_1462,N_1074,N_1034);
xnor U1463 (N_1463,N_1157,N_1028);
nor U1464 (N_1464,N_1173,N_1183);
or U1465 (N_1465,N_1192,N_957);
and U1466 (N_1466,N_977,N_1033);
or U1467 (N_1467,N_1128,N_934);
nor U1468 (N_1468,N_1162,N_1089);
xor U1469 (N_1469,N_900,N_1159);
nand U1470 (N_1470,N_1182,N_1053);
and U1471 (N_1471,N_907,N_961);
nand U1472 (N_1472,N_963,N_1022);
nor U1473 (N_1473,N_902,N_901);
nand U1474 (N_1474,N_970,N_1084);
or U1475 (N_1475,N_1194,N_939);
and U1476 (N_1476,N_1183,N_998);
nor U1477 (N_1477,N_1051,N_992);
and U1478 (N_1478,N_1158,N_1058);
and U1479 (N_1479,N_1108,N_1063);
nor U1480 (N_1480,N_1090,N_1006);
and U1481 (N_1481,N_916,N_931);
and U1482 (N_1482,N_1007,N_1080);
or U1483 (N_1483,N_957,N_1020);
xnor U1484 (N_1484,N_1118,N_1061);
nand U1485 (N_1485,N_1048,N_1052);
nand U1486 (N_1486,N_990,N_1077);
nand U1487 (N_1487,N_1050,N_1171);
or U1488 (N_1488,N_976,N_931);
nor U1489 (N_1489,N_955,N_1199);
nand U1490 (N_1490,N_1027,N_1037);
or U1491 (N_1491,N_1034,N_1127);
nor U1492 (N_1492,N_946,N_1101);
nand U1493 (N_1493,N_993,N_1130);
or U1494 (N_1494,N_1032,N_1120);
or U1495 (N_1495,N_990,N_910);
nand U1496 (N_1496,N_999,N_1187);
or U1497 (N_1497,N_1016,N_1133);
nand U1498 (N_1498,N_954,N_936);
nand U1499 (N_1499,N_1124,N_1017);
or U1500 (N_1500,N_1379,N_1345);
nor U1501 (N_1501,N_1326,N_1392);
nand U1502 (N_1502,N_1406,N_1347);
and U1503 (N_1503,N_1352,N_1495);
xnor U1504 (N_1504,N_1258,N_1290);
xnor U1505 (N_1505,N_1436,N_1362);
nand U1506 (N_1506,N_1405,N_1282);
or U1507 (N_1507,N_1200,N_1480);
nand U1508 (N_1508,N_1264,N_1312);
xor U1509 (N_1509,N_1297,N_1434);
and U1510 (N_1510,N_1230,N_1241);
xnor U1511 (N_1511,N_1284,N_1412);
and U1512 (N_1512,N_1265,N_1250);
or U1513 (N_1513,N_1219,N_1270);
xor U1514 (N_1514,N_1422,N_1260);
and U1515 (N_1515,N_1215,N_1237);
xor U1516 (N_1516,N_1202,N_1232);
nand U1517 (N_1517,N_1280,N_1369);
or U1518 (N_1518,N_1397,N_1466);
or U1519 (N_1519,N_1387,N_1273);
nand U1520 (N_1520,N_1337,N_1207);
nand U1521 (N_1521,N_1228,N_1209);
or U1522 (N_1522,N_1233,N_1238);
and U1523 (N_1523,N_1400,N_1223);
or U1524 (N_1524,N_1229,N_1225);
nor U1525 (N_1525,N_1256,N_1363);
nor U1526 (N_1526,N_1383,N_1445);
and U1527 (N_1527,N_1309,N_1303);
and U1528 (N_1528,N_1221,N_1449);
nand U1529 (N_1529,N_1319,N_1351);
nand U1530 (N_1530,N_1361,N_1304);
nor U1531 (N_1531,N_1401,N_1353);
nor U1532 (N_1532,N_1349,N_1458);
nor U1533 (N_1533,N_1399,N_1205);
nor U1534 (N_1534,N_1269,N_1486);
xnor U1535 (N_1535,N_1492,N_1371);
and U1536 (N_1536,N_1360,N_1462);
xor U1537 (N_1537,N_1453,N_1285);
nand U1538 (N_1538,N_1451,N_1490);
or U1539 (N_1539,N_1427,N_1268);
nand U1540 (N_1540,N_1348,N_1300);
xnor U1541 (N_1541,N_1407,N_1472);
nor U1542 (N_1542,N_1204,N_1414);
nand U1543 (N_1543,N_1313,N_1263);
xnor U1544 (N_1544,N_1368,N_1343);
nor U1545 (N_1545,N_1419,N_1333);
nor U1546 (N_1546,N_1331,N_1432);
and U1547 (N_1547,N_1247,N_1289);
and U1548 (N_1548,N_1234,N_1336);
nor U1549 (N_1549,N_1306,N_1327);
and U1550 (N_1550,N_1378,N_1315);
nand U1551 (N_1551,N_1271,N_1307);
nor U1552 (N_1552,N_1267,N_1311);
xor U1553 (N_1553,N_1213,N_1310);
and U1554 (N_1554,N_1208,N_1476);
nand U1555 (N_1555,N_1496,N_1474);
nor U1556 (N_1556,N_1467,N_1291);
or U1557 (N_1557,N_1497,N_1342);
or U1558 (N_1558,N_1236,N_1418);
and U1559 (N_1559,N_1388,N_1257);
xor U1560 (N_1560,N_1464,N_1469);
and U1561 (N_1561,N_1416,N_1372);
or U1562 (N_1562,N_1424,N_1356);
or U1563 (N_1563,N_1428,N_1235);
and U1564 (N_1564,N_1296,N_1346);
and U1565 (N_1565,N_1358,N_1435);
or U1566 (N_1566,N_1266,N_1277);
nor U1567 (N_1567,N_1222,N_1354);
nor U1568 (N_1568,N_1366,N_1301);
and U1569 (N_1569,N_1377,N_1485);
and U1570 (N_1570,N_1365,N_1364);
nor U1571 (N_1571,N_1384,N_1450);
or U1572 (N_1572,N_1488,N_1394);
nor U1573 (N_1573,N_1275,N_1477);
xnor U1574 (N_1574,N_1386,N_1463);
or U1575 (N_1575,N_1456,N_1339);
nand U1576 (N_1576,N_1396,N_1433);
nor U1577 (N_1577,N_1447,N_1210);
nor U1578 (N_1578,N_1468,N_1441);
and U1579 (N_1579,N_1359,N_1431);
and U1580 (N_1580,N_1211,N_1494);
nand U1581 (N_1581,N_1295,N_1376);
nor U1582 (N_1582,N_1478,N_1212);
or U1583 (N_1583,N_1410,N_1471);
and U1584 (N_1584,N_1324,N_1465);
xnor U1585 (N_1585,N_1243,N_1214);
xor U1586 (N_1586,N_1218,N_1389);
nand U1587 (N_1587,N_1314,N_1374);
nand U1588 (N_1588,N_1201,N_1344);
and U1589 (N_1589,N_1261,N_1459);
or U1590 (N_1590,N_1370,N_1413);
or U1591 (N_1591,N_1231,N_1323);
xor U1592 (N_1592,N_1278,N_1489);
nor U1593 (N_1593,N_1240,N_1252);
nor U1594 (N_1594,N_1475,N_1398);
and U1595 (N_1595,N_1249,N_1224);
and U1596 (N_1596,N_1409,N_1251);
nand U1597 (N_1597,N_1391,N_1440);
xnor U1598 (N_1598,N_1421,N_1457);
xor U1599 (N_1599,N_1294,N_1334);
or U1600 (N_1600,N_1439,N_1382);
or U1601 (N_1601,N_1227,N_1206);
xnor U1602 (N_1602,N_1417,N_1385);
nor U1603 (N_1603,N_1322,N_1253);
and U1604 (N_1604,N_1443,N_1246);
or U1605 (N_1605,N_1481,N_1338);
nor U1606 (N_1606,N_1317,N_1293);
nand U1607 (N_1607,N_1242,N_1438);
nand U1608 (N_1608,N_1281,N_1473);
or U1609 (N_1609,N_1255,N_1444);
or U1610 (N_1610,N_1332,N_1248);
nor U1611 (N_1611,N_1454,N_1262);
and U1612 (N_1612,N_1355,N_1491);
nand U1613 (N_1613,N_1320,N_1393);
nor U1614 (N_1614,N_1493,N_1498);
nor U1615 (N_1615,N_1216,N_1272);
xnor U1616 (N_1616,N_1380,N_1461);
or U1617 (N_1617,N_1402,N_1276);
xnor U1618 (N_1618,N_1239,N_1318);
xnor U1619 (N_1619,N_1423,N_1203);
nor U1620 (N_1620,N_1429,N_1254);
xor U1621 (N_1621,N_1442,N_1437);
nor U1622 (N_1622,N_1305,N_1287);
and U1623 (N_1623,N_1302,N_1357);
or U1624 (N_1624,N_1483,N_1446);
xnor U1625 (N_1625,N_1217,N_1487);
or U1626 (N_1626,N_1482,N_1321);
nor U1627 (N_1627,N_1330,N_1340);
or U1628 (N_1628,N_1408,N_1373);
nand U1629 (N_1629,N_1430,N_1367);
nor U1630 (N_1630,N_1341,N_1415);
nand U1631 (N_1631,N_1325,N_1470);
nand U1632 (N_1632,N_1460,N_1335);
or U1633 (N_1633,N_1279,N_1420);
and U1634 (N_1634,N_1328,N_1329);
nand U1635 (N_1635,N_1274,N_1226);
or U1636 (N_1636,N_1452,N_1292);
nor U1637 (N_1637,N_1308,N_1448);
nand U1638 (N_1638,N_1390,N_1245);
and U1639 (N_1639,N_1479,N_1395);
or U1640 (N_1640,N_1244,N_1299);
nor U1641 (N_1641,N_1403,N_1425);
nand U1642 (N_1642,N_1220,N_1288);
and U1643 (N_1643,N_1404,N_1426);
and U1644 (N_1644,N_1499,N_1381);
nor U1645 (N_1645,N_1411,N_1484);
or U1646 (N_1646,N_1298,N_1350);
or U1647 (N_1647,N_1259,N_1286);
or U1648 (N_1648,N_1375,N_1316);
nand U1649 (N_1649,N_1455,N_1283);
xnor U1650 (N_1650,N_1419,N_1472);
xnor U1651 (N_1651,N_1322,N_1474);
or U1652 (N_1652,N_1300,N_1384);
nor U1653 (N_1653,N_1413,N_1493);
or U1654 (N_1654,N_1357,N_1374);
and U1655 (N_1655,N_1364,N_1371);
nor U1656 (N_1656,N_1377,N_1252);
or U1657 (N_1657,N_1269,N_1200);
and U1658 (N_1658,N_1233,N_1375);
nand U1659 (N_1659,N_1496,N_1278);
nand U1660 (N_1660,N_1215,N_1287);
xnor U1661 (N_1661,N_1272,N_1226);
nand U1662 (N_1662,N_1206,N_1288);
xnor U1663 (N_1663,N_1243,N_1211);
nor U1664 (N_1664,N_1492,N_1201);
or U1665 (N_1665,N_1380,N_1234);
nand U1666 (N_1666,N_1362,N_1300);
and U1667 (N_1667,N_1420,N_1275);
and U1668 (N_1668,N_1282,N_1380);
xor U1669 (N_1669,N_1262,N_1227);
xnor U1670 (N_1670,N_1230,N_1456);
or U1671 (N_1671,N_1375,N_1439);
xnor U1672 (N_1672,N_1392,N_1456);
or U1673 (N_1673,N_1391,N_1369);
xor U1674 (N_1674,N_1491,N_1290);
nor U1675 (N_1675,N_1225,N_1440);
and U1676 (N_1676,N_1267,N_1260);
nor U1677 (N_1677,N_1369,N_1449);
nor U1678 (N_1678,N_1379,N_1325);
or U1679 (N_1679,N_1451,N_1394);
and U1680 (N_1680,N_1478,N_1299);
or U1681 (N_1681,N_1395,N_1225);
nand U1682 (N_1682,N_1249,N_1462);
or U1683 (N_1683,N_1396,N_1430);
nand U1684 (N_1684,N_1250,N_1249);
nor U1685 (N_1685,N_1263,N_1273);
xor U1686 (N_1686,N_1372,N_1493);
xor U1687 (N_1687,N_1245,N_1483);
nor U1688 (N_1688,N_1479,N_1359);
nand U1689 (N_1689,N_1431,N_1406);
nand U1690 (N_1690,N_1288,N_1448);
xor U1691 (N_1691,N_1297,N_1320);
nand U1692 (N_1692,N_1484,N_1252);
nor U1693 (N_1693,N_1317,N_1397);
nor U1694 (N_1694,N_1257,N_1299);
nand U1695 (N_1695,N_1318,N_1365);
and U1696 (N_1696,N_1408,N_1277);
and U1697 (N_1697,N_1351,N_1303);
or U1698 (N_1698,N_1483,N_1234);
or U1699 (N_1699,N_1318,N_1379);
nand U1700 (N_1700,N_1224,N_1355);
xor U1701 (N_1701,N_1372,N_1324);
nor U1702 (N_1702,N_1490,N_1388);
nor U1703 (N_1703,N_1499,N_1361);
and U1704 (N_1704,N_1380,N_1474);
or U1705 (N_1705,N_1430,N_1230);
xnor U1706 (N_1706,N_1250,N_1372);
nand U1707 (N_1707,N_1264,N_1484);
and U1708 (N_1708,N_1444,N_1355);
xnor U1709 (N_1709,N_1208,N_1364);
and U1710 (N_1710,N_1257,N_1262);
nor U1711 (N_1711,N_1296,N_1208);
nand U1712 (N_1712,N_1359,N_1207);
xnor U1713 (N_1713,N_1232,N_1496);
xnor U1714 (N_1714,N_1417,N_1228);
and U1715 (N_1715,N_1423,N_1435);
nor U1716 (N_1716,N_1303,N_1200);
and U1717 (N_1717,N_1377,N_1433);
or U1718 (N_1718,N_1239,N_1472);
xnor U1719 (N_1719,N_1460,N_1275);
xnor U1720 (N_1720,N_1329,N_1296);
or U1721 (N_1721,N_1266,N_1445);
nand U1722 (N_1722,N_1417,N_1313);
xor U1723 (N_1723,N_1363,N_1245);
or U1724 (N_1724,N_1421,N_1272);
or U1725 (N_1725,N_1350,N_1232);
and U1726 (N_1726,N_1408,N_1321);
nor U1727 (N_1727,N_1295,N_1279);
nor U1728 (N_1728,N_1475,N_1410);
xnor U1729 (N_1729,N_1398,N_1294);
nand U1730 (N_1730,N_1314,N_1290);
or U1731 (N_1731,N_1371,N_1318);
and U1732 (N_1732,N_1334,N_1476);
and U1733 (N_1733,N_1471,N_1348);
xnor U1734 (N_1734,N_1485,N_1334);
xor U1735 (N_1735,N_1254,N_1454);
nor U1736 (N_1736,N_1208,N_1468);
or U1737 (N_1737,N_1481,N_1464);
xor U1738 (N_1738,N_1242,N_1363);
and U1739 (N_1739,N_1337,N_1335);
nand U1740 (N_1740,N_1325,N_1497);
xnor U1741 (N_1741,N_1391,N_1242);
nand U1742 (N_1742,N_1452,N_1357);
nor U1743 (N_1743,N_1483,N_1315);
nor U1744 (N_1744,N_1231,N_1295);
or U1745 (N_1745,N_1269,N_1476);
or U1746 (N_1746,N_1343,N_1249);
nor U1747 (N_1747,N_1284,N_1322);
and U1748 (N_1748,N_1358,N_1421);
nand U1749 (N_1749,N_1264,N_1433);
nand U1750 (N_1750,N_1228,N_1380);
xor U1751 (N_1751,N_1255,N_1267);
nor U1752 (N_1752,N_1319,N_1336);
or U1753 (N_1753,N_1235,N_1233);
nor U1754 (N_1754,N_1207,N_1330);
or U1755 (N_1755,N_1488,N_1389);
or U1756 (N_1756,N_1422,N_1259);
nor U1757 (N_1757,N_1425,N_1433);
xnor U1758 (N_1758,N_1480,N_1205);
nand U1759 (N_1759,N_1447,N_1253);
or U1760 (N_1760,N_1345,N_1224);
and U1761 (N_1761,N_1457,N_1477);
nand U1762 (N_1762,N_1228,N_1443);
or U1763 (N_1763,N_1391,N_1442);
and U1764 (N_1764,N_1400,N_1338);
and U1765 (N_1765,N_1234,N_1360);
or U1766 (N_1766,N_1225,N_1386);
xnor U1767 (N_1767,N_1336,N_1299);
and U1768 (N_1768,N_1470,N_1263);
nand U1769 (N_1769,N_1358,N_1426);
xor U1770 (N_1770,N_1477,N_1463);
nor U1771 (N_1771,N_1256,N_1436);
xnor U1772 (N_1772,N_1269,N_1230);
and U1773 (N_1773,N_1264,N_1396);
xor U1774 (N_1774,N_1467,N_1268);
nand U1775 (N_1775,N_1209,N_1339);
nand U1776 (N_1776,N_1201,N_1448);
and U1777 (N_1777,N_1493,N_1257);
xnor U1778 (N_1778,N_1255,N_1358);
and U1779 (N_1779,N_1326,N_1437);
nand U1780 (N_1780,N_1332,N_1235);
nand U1781 (N_1781,N_1285,N_1430);
or U1782 (N_1782,N_1478,N_1424);
or U1783 (N_1783,N_1311,N_1431);
nor U1784 (N_1784,N_1257,N_1324);
and U1785 (N_1785,N_1331,N_1216);
nor U1786 (N_1786,N_1235,N_1210);
nand U1787 (N_1787,N_1378,N_1493);
nand U1788 (N_1788,N_1425,N_1376);
and U1789 (N_1789,N_1296,N_1383);
nand U1790 (N_1790,N_1385,N_1299);
and U1791 (N_1791,N_1238,N_1456);
or U1792 (N_1792,N_1363,N_1203);
xor U1793 (N_1793,N_1294,N_1209);
and U1794 (N_1794,N_1293,N_1347);
and U1795 (N_1795,N_1252,N_1454);
nand U1796 (N_1796,N_1309,N_1377);
nand U1797 (N_1797,N_1466,N_1233);
nor U1798 (N_1798,N_1439,N_1342);
nand U1799 (N_1799,N_1454,N_1288);
and U1800 (N_1800,N_1587,N_1681);
xnor U1801 (N_1801,N_1791,N_1527);
or U1802 (N_1802,N_1513,N_1611);
and U1803 (N_1803,N_1603,N_1741);
xor U1804 (N_1804,N_1636,N_1652);
nor U1805 (N_1805,N_1761,N_1610);
xnor U1806 (N_1806,N_1789,N_1702);
xnor U1807 (N_1807,N_1774,N_1629);
xor U1808 (N_1808,N_1614,N_1539);
nor U1809 (N_1809,N_1787,N_1695);
nor U1810 (N_1810,N_1512,N_1550);
or U1811 (N_1811,N_1618,N_1536);
nand U1812 (N_1812,N_1660,N_1646);
or U1813 (N_1813,N_1534,N_1654);
and U1814 (N_1814,N_1622,N_1708);
nand U1815 (N_1815,N_1548,N_1678);
or U1816 (N_1816,N_1540,N_1692);
nand U1817 (N_1817,N_1743,N_1552);
nor U1818 (N_1818,N_1549,N_1572);
or U1819 (N_1819,N_1634,N_1713);
and U1820 (N_1820,N_1686,N_1505);
nand U1821 (N_1821,N_1580,N_1560);
xnor U1822 (N_1822,N_1746,N_1579);
nand U1823 (N_1823,N_1775,N_1597);
or U1824 (N_1824,N_1518,N_1767);
nor U1825 (N_1825,N_1737,N_1734);
and U1826 (N_1826,N_1592,N_1638);
and U1827 (N_1827,N_1709,N_1687);
nand U1828 (N_1828,N_1680,N_1724);
nand U1829 (N_1829,N_1684,N_1595);
nand U1830 (N_1830,N_1751,N_1707);
or U1831 (N_1831,N_1764,N_1798);
xnor U1832 (N_1832,N_1656,N_1703);
xor U1833 (N_1833,N_1717,N_1691);
nand U1834 (N_1834,N_1779,N_1528);
and U1835 (N_1835,N_1665,N_1671);
xnor U1836 (N_1836,N_1768,N_1542);
xnor U1837 (N_1837,N_1771,N_1613);
nor U1838 (N_1838,N_1608,N_1586);
and U1839 (N_1839,N_1716,N_1705);
nand U1840 (N_1840,N_1625,N_1555);
nand U1841 (N_1841,N_1679,N_1601);
or U1842 (N_1842,N_1753,N_1551);
and U1843 (N_1843,N_1759,N_1696);
or U1844 (N_1844,N_1710,N_1756);
or U1845 (N_1845,N_1624,N_1711);
nand U1846 (N_1846,N_1514,N_1793);
xor U1847 (N_1847,N_1644,N_1591);
nor U1848 (N_1848,N_1570,N_1720);
or U1849 (N_1849,N_1571,N_1739);
nor U1850 (N_1850,N_1783,N_1772);
nor U1851 (N_1851,N_1668,N_1784);
and U1852 (N_1852,N_1576,N_1502);
or U1853 (N_1853,N_1564,N_1547);
or U1854 (N_1854,N_1565,N_1590);
nand U1855 (N_1855,N_1732,N_1581);
nor U1856 (N_1856,N_1525,N_1790);
nor U1857 (N_1857,N_1728,N_1504);
xor U1858 (N_1858,N_1569,N_1503);
or U1859 (N_1859,N_1511,N_1657);
and U1860 (N_1860,N_1796,N_1604);
and U1861 (N_1861,N_1749,N_1606);
xor U1862 (N_1862,N_1556,N_1619);
nor U1863 (N_1863,N_1718,N_1651);
or U1864 (N_1864,N_1785,N_1582);
and U1865 (N_1865,N_1689,N_1723);
nor U1866 (N_1866,N_1721,N_1522);
xor U1867 (N_1867,N_1704,N_1637);
and U1868 (N_1868,N_1607,N_1700);
and U1869 (N_1869,N_1593,N_1635);
xnor U1870 (N_1870,N_1612,N_1596);
nand U1871 (N_1871,N_1529,N_1517);
nand U1872 (N_1872,N_1735,N_1726);
or U1873 (N_1873,N_1788,N_1698);
and U1874 (N_1874,N_1575,N_1500);
or U1875 (N_1875,N_1538,N_1760);
xor U1876 (N_1876,N_1633,N_1758);
nand U1877 (N_1877,N_1740,N_1562);
nor U1878 (N_1878,N_1567,N_1515);
or U1879 (N_1879,N_1588,N_1541);
nor U1880 (N_1880,N_1583,N_1672);
nand U1881 (N_1881,N_1545,N_1757);
nand U1882 (N_1882,N_1766,N_1674);
or U1883 (N_1883,N_1670,N_1677);
nand U1884 (N_1884,N_1714,N_1508);
or U1885 (N_1885,N_1568,N_1747);
and U1886 (N_1886,N_1778,N_1520);
or U1887 (N_1887,N_1566,N_1530);
nor U1888 (N_1888,N_1594,N_1537);
nor U1889 (N_1889,N_1647,N_1676);
nand U1890 (N_1890,N_1605,N_1682);
nand U1891 (N_1891,N_1697,N_1573);
or U1892 (N_1892,N_1762,N_1533);
nor U1893 (N_1893,N_1685,N_1577);
or U1894 (N_1894,N_1763,N_1782);
xor U1895 (N_1895,N_1627,N_1616);
nand U1896 (N_1896,N_1799,N_1706);
nand U1897 (N_1897,N_1731,N_1744);
nor U1898 (N_1898,N_1509,N_1786);
or U1899 (N_1899,N_1535,N_1725);
xor U1900 (N_1900,N_1609,N_1712);
nor U1901 (N_1901,N_1554,N_1752);
nor U1902 (N_1902,N_1795,N_1645);
nor U1903 (N_1903,N_1683,N_1715);
xor U1904 (N_1904,N_1532,N_1755);
xor U1905 (N_1905,N_1543,N_1599);
xor U1906 (N_1906,N_1623,N_1584);
nor U1907 (N_1907,N_1643,N_1516);
nor U1908 (N_1908,N_1510,N_1776);
nand U1909 (N_1909,N_1701,N_1648);
or U1910 (N_1910,N_1598,N_1585);
and U1911 (N_1911,N_1639,N_1777);
or U1912 (N_1912,N_1736,N_1770);
nor U1913 (N_1913,N_1693,N_1563);
and U1914 (N_1914,N_1673,N_1675);
nor U1915 (N_1915,N_1750,N_1773);
or U1916 (N_1916,N_1501,N_1559);
nand U1917 (N_1917,N_1655,N_1523);
nor U1918 (N_1918,N_1506,N_1658);
nor U1919 (N_1919,N_1653,N_1589);
nand U1920 (N_1920,N_1663,N_1600);
nor U1921 (N_1921,N_1729,N_1602);
or U1922 (N_1922,N_1667,N_1632);
or U1923 (N_1923,N_1621,N_1519);
nor U1924 (N_1924,N_1666,N_1558);
and U1925 (N_1925,N_1688,N_1617);
xor U1926 (N_1926,N_1662,N_1615);
xnor U1927 (N_1927,N_1631,N_1557);
and U1928 (N_1928,N_1641,N_1745);
nor U1929 (N_1929,N_1620,N_1630);
xor U1930 (N_1930,N_1578,N_1524);
nand U1931 (N_1931,N_1574,N_1733);
nor U1932 (N_1932,N_1738,N_1765);
nor U1933 (N_1933,N_1628,N_1626);
and U1934 (N_1934,N_1649,N_1669);
nor U1935 (N_1935,N_1699,N_1526);
or U1936 (N_1936,N_1780,N_1546);
nor U1937 (N_1937,N_1719,N_1659);
nand U1938 (N_1938,N_1794,N_1544);
and U1939 (N_1939,N_1664,N_1690);
xnor U1940 (N_1940,N_1642,N_1661);
nand U1941 (N_1941,N_1640,N_1769);
nand U1942 (N_1942,N_1507,N_1781);
or U1943 (N_1943,N_1797,N_1531);
nand U1944 (N_1944,N_1792,N_1748);
or U1945 (N_1945,N_1694,N_1742);
or U1946 (N_1946,N_1650,N_1561);
or U1947 (N_1947,N_1727,N_1754);
xor U1948 (N_1948,N_1722,N_1521);
xor U1949 (N_1949,N_1730,N_1553);
nand U1950 (N_1950,N_1506,N_1739);
nand U1951 (N_1951,N_1641,N_1701);
or U1952 (N_1952,N_1691,N_1708);
nand U1953 (N_1953,N_1715,N_1594);
nor U1954 (N_1954,N_1648,N_1719);
and U1955 (N_1955,N_1677,N_1779);
nor U1956 (N_1956,N_1631,N_1597);
nor U1957 (N_1957,N_1779,N_1667);
xnor U1958 (N_1958,N_1671,N_1504);
nand U1959 (N_1959,N_1670,N_1550);
and U1960 (N_1960,N_1593,N_1543);
or U1961 (N_1961,N_1554,N_1570);
nor U1962 (N_1962,N_1743,N_1624);
nor U1963 (N_1963,N_1676,N_1654);
nand U1964 (N_1964,N_1662,N_1698);
xnor U1965 (N_1965,N_1645,N_1601);
or U1966 (N_1966,N_1631,N_1532);
or U1967 (N_1967,N_1692,N_1657);
nor U1968 (N_1968,N_1686,N_1567);
nor U1969 (N_1969,N_1634,N_1594);
and U1970 (N_1970,N_1738,N_1758);
nand U1971 (N_1971,N_1609,N_1523);
nand U1972 (N_1972,N_1536,N_1592);
xor U1973 (N_1973,N_1756,N_1522);
nand U1974 (N_1974,N_1759,N_1500);
xor U1975 (N_1975,N_1534,N_1586);
nor U1976 (N_1976,N_1575,N_1593);
or U1977 (N_1977,N_1651,N_1677);
nor U1978 (N_1978,N_1584,N_1656);
nor U1979 (N_1979,N_1655,N_1756);
or U1980 (N_1980,N_1633,N_1554);
xnor U1981 (N_1981,N_1718,N_1695);
and U1982 (N_1982,N_1760,N_1727);
nand U1983 (N_1983,N_1560,N_1672);
or U1984 (N_1984,N_1617,N_1619);
or U1985 (N_1985,N_1680,N_1603);
and U1986 (N_1986,N_1700,N_1677);
xnor U1987 (N_1987,N_1635,N_1530);
nand U1988 (N_1988,N_1751,N_1673);
xor U1989 (N_1989,N_1578,N_1725);
nor U1990 (N_1990,N_1609,N_1518);
or U1991 (N_1991,N_1540,N_1506);
nand U1992 (N_1992,N_1774,N_1662);
xor U1993 (N_1993,N_1534,N_1751);
xor U1994 (N_1994,N_1562,N_1571);
nand U1995 (N_1995,N_1538,N_1579);
or U1996 (N_1996,N_1611,N_1705);
nor U1997 (N_1997,N_1568,N_1674);
nor U1998 (N_1998,N_1704,N_1646);
and U1999 (N_1999,N_1724,N_1584);
and U2000 (N_2000,N_1779,N_1605);
nor U2001 (N_2001,N_1603,N_1686);
nor U2002 (N_2002,N_1715,N_1798);
nand U2003 (N_2003,N_1735,N_1618);
xnor U2004 (N_2004,N_1567,N_1587);
nand U2005 (N_2005,N_1570,N_1580);
nand U2006 (N_2006,N_1732,N_1617);
or U2007 (N_2007,N_1699,N_1693);
xor U2008 (N_2008,N_1525,N_1532);
nor U2009 (N_2009,N_1734,N_1626);
nor U2010 (N_2010,N_1539,N_1598);
nand U2011 (N_2011,N_1538,N_1540);
or U2012 (N_2012,N_1697,N_1602);
or U2013 (N_2013,N_1771,N_1649);
and U2014 (N_2014,N_1625,N_1709);
nor U2015 (N_2015,N_1743,N_1774);
and U2016 (N_2016,N_1721,N_1673);
or U2017 (N_2017,N_1731,N_1571);
and U2018 (N_2018,N_1526,N_1593);
and U2019 (N_2019,N_1595,N_1772);
or U2020 (N_2020,N_1733,N_1572);
nor U2021 (N_2021,N_1727,N_1694);
nand U2022 (N_2022,N_1629,N_1515);
nor U2023 (N_2023,N_1692,N_1783);
nor U2024 (N_2024,N_1738,N_1577);
or U2025 (N_2025,N_1547,N_1576);
and U2026 (N_2026,N_1675,N_1719);
nor U2027 (N_2027,N_1733,N_1546);
nand U2028 (N_2028,N_1619,N_1614);
or U2029 (N_2029,N_1512,N_1567);
xor U2030 (N_2030,N_1573,N_1775);
nor U2031 (N_2031,N_1688,N_1564);
nor U2032 (N_2032,N_1611,N_1508);
xor U2033 (N_2033,N_1552,N_1687);
nor U2034 (N_2034,N_1786,N_1553);
nand U2035 (N_2035,N_1588,N_1641);
nand U2036 (N_2036,N_1782,N_1705);
nor U2037 (N_2037,N_1681,N_1682);
and U2038 (N_2038,N_1622,N_1679);
nor U2039 (N_2039,N_1589,N_1687);
or U2040 (N_2040,N_1662,N_1760);
and U2041 (N_2041,N_1671,N_1582);
or U2042 (N_2042,N_1546,N_1529);
nand U2043 (N_2043,N_1799,N_1521);
nor U2044 (N_2044,N_1646,N_1567);
and U2045 (N_2045,N_1577,N_1739);
or U2046 (N_2046,N_1509,N_1734);
and U2047 (N_2047,N_1760,N_1597);
or U2048 (N_2048,N_1696,N_1738);
nor U2049 (N_2049,N_1520,N_1515);
or U2050 (N_2050,N_1610,N_1744);
xor U2051 (N_2051,N_1612,N_1553);
nor U2052 (N_2052,N_1605,N_1644);
or U2053 (N_2053,N_1731,N_1540);
xor U2054 (N_2054,N_1759,N_1769);
xnor U2055 (N_2055,N_1781,N_1528);
xor U2056 (N_2056,N_1519,N_1513);
xor U2057 (N_2057,N_1597,N_1746);
nor U2058 (N_2058,N_1661,N_1575);
or U2059 (N_2059,N_1539,N_1798);
nand U2060 (N_2060,N_1675,N_1626);
nor U2061 (N_2061,N_1672,N_1570);
nor U2062 (N_2062,N_1744,N_1633);
nor U2063 (N_2063,N_1688,N_1700);
or U2064 (N_2064,N_1684,N_1746);
or U2065 (N_2065,N_1642,N_1741);
nand U2066 (N_2066,N_1770,N_1684);
or U2067 (N_2067,N_1512,N_1709);
nand U2068 (N_2068,N_1730,N_1776);
xor U2069 (N_2069,N_1697,N_1685);
nor U2070 (N_2070,N_1634,N_1685);
nand U2071 (N_2071,N_1506,N_1635);
and U2072 (N_2072,N_1534,N_1643);
and U2073 (N_2073,N_1586,N_1638);
nand U2074 (N_2074,N_1778,N_1588);
nor U2075 (N_2075,N_1783,N_1690);
or U2076 (N_2076,N_1682,N_1662);
and U2077 (N_2077,N_1765,N_1754);
xnor U2078 (N_2078,N_1702,N_1539);
nand U2079 (N_2079,N_1576,N_1500);
nand U2080 (N_2080,N_1566,N_1757);
and U2081 (N_2081,N_1655,N_1769);
and U2082 (N_2082,N_1623,N_1609);
xnor U2083 (N_2083,N_1779,N_1581);
or U2084 (N_2084,N_1622,N_1621);
and U2085 (N_2085,N_1685,N_1750);
nand U2086 (N_2086,N_1560,N_1582);
nand U2087 (N_2087,N_1716,N_1646);
or U2088 (N_2088,N_1626,N_1690);
xnor U2089 (N_2089,N_1598,N_1548);
xor U2090 (N_2090,N_1627,N_1648);
or U2091 (N_2091,N_1760,N_1539);
and U2092 (N_2092,N_1725,N_1669);
xor U2093 (N_2093,N_1540,N_1695);
xor U2094 (N_2094,N_1536,N_1531);
nand U2095 (N_2095,N_1534,N_1701);
and U2096 (N_2096,N_1595,N_1529);
xnor U2097 (N_2097,N_1629,N_1663);
or U2098 (N_2098,N_1756,N_1501);
xnor U2099 (N_2099,N_1508,N_1726);
nand U2100 (N_2100,N_1925,N_2049);
and U2101 (N_2101,N_1939,N_1856);
nand U2102 (N_2102,N_2083,N_1974);
nand U2103 (N_2103,N_1881,N_1801);
nor U2104 (N_2104,N_1833,N_2027);
xnor U2105 (N_2105,N_1943,N_2099);
xor U2106 (N_2106,N_1844,N_2096);
or U2107 (N_2107,N_2055,N_2064);
xor U2108 (N_2108,N_1824,N_2056);
nor U2109 (N_2109,N_1828,N_2067);
and U2110 (N_2110,N_2035,N_2072);
or U2111 (N_2111,N_1859,N_1810);
xor U2112 (N_2112,N_1924,N_2018);
and U2113 (N_2113,N_1904,N_1841);
nand U2114 (N_2114,N_2048,N_1911);
nand U2115 (N_2115,N_1890,N_2097);
and U2116 (N_2116,N_1807,N_1851);
and U2117 (N_2117,N_1854,N_1991);
nand U2118 (N_2118,N_2063,N_1944);
xor U2119 (N_2119,N_1948,N_1889);
xor U2120 (N_2120,N_1843,N_1933);
and U2121 (N_2121,N_1966,N_2006);
and U2122 (N_2122,N_1817,N_2069);
or U2123 (N_2123,N_2008,N_1831);
or U2124 (N_2124,N_1829,N_1835);
xnor U2125 (N_2125,N_1969,N_1962);
nand U2126 (N_2126,N_2038,N_1899);
nand U2127 (N_2127,N_1814,N_1901);
nor U2128 (N_2128,N_1955,N_2002);
nor U2129 (N_2129,N_2082,N_1910);
xnor U2130 (N_2130,N_2052,N_2085);
and U2131 (N_2131,N_2065,N_2098);
nand U2132 (N_2132,N_1845,N_1877);
nor U2133 (N_2133,N_1909,N_1903);
and U2134 (N_2134,N_2050,N_2060);
or U2135 (N_2135,N_2093,N_2051);
xnor U2136 (N_2136,N_1802,N_1972);
nand U2137 (N_2137,N_1968,N_1998);
nand U2138 (N_2138,N_1941,N_2005);
or U2139 (N_2139,N_2086,N_1971);
nand U2140 (N_2140,N_1945,N_2075);
nand U2141 (N_2141,N_1888,N_1914);
nor U2142 (N_2142,N_1860,N_1883);
nor U2143 (N_2143,N_1973,N_1999);
or U2144 (N_2144,N_2031,N_1842);
or U2145 (N_2145,N_1989,N_1976);
xor U2146 (N_2146,N_2009,N_2054);
and U2147 (N_2147,N_2045,N_1988);
or U2148 (N_2148,N_1997,N_2017);
xnor U2149 (N_2149,N_1876,N_1895);
nand U2150 (N_2150,N_1803,N_2020);
nor U2151 (N_2151,N_1894,N_1806);
or U2152 (N_2152,N_2077,N_1867);
or U2153 (N_2153,N_1953,N_2012);
and U2154 (N_2154,N_2028,N_1957);
or U2155 (N_2155,N_1961,N_1846);
xnor U2156 (N_2156,N_1855,N_1872);
xor U2157 (N_2157,N_1800,N_2080);
xor U2158 (N_2158,N_1849,N_1866);
xor U2159 (N_2159,N_1805,N_2090);
and U2160 (N_2160,N_1879,N_2047);
nor U2161 (N_2161,N_1908,N_2032);
and U2162 (N_2162,N_1886,N_1907);
xnor U2163 (N_2163,N_2003,N_1900);
nand U2164 (N_2164,N_1956,N_1868);
nand U2165 (N_2165,N_1946,N_2068);
nor U2166 (N_2166,N_1947,N_1898);
xnor U2167 (N_2167,N_1864,N_1874);
nand U2168 (N_2168,N_2013,N_2010);
nand U2169 (N_2169,N_1906,N_1813);
nand U2170 (N_2170,N_1830,N_1836);
and U2171 (N_2171,N_1847,N_1878);
nand U2172 (N_2172,N_1819,N_2034);
and U2173 (N_2173,N_2039,N_1981);
or U2174 (N_2174,N_1934,N_1921);
nand U2175 (N_2175,N_1954,N_1808);
nand U2176 (N_2176,N_2059,N_1926);
and U2177 (N_2177,N_1990,N_2021);
nor U2178 (N_2178,N_2016,N_2043);
nor U2179 (N_2179,N_1994,N_1858);
nand U2180 (N_2180,N_1928,N_1963);
or U2181 (N_2181,N_1865,N_1960);
xor U2182 (N_2182,N_1970,N_1861);
xnor U2183 (N_2183,N_2074,N_1893);
and U2184 (N_2184,N_2011,N_1915);
and U2185 (N_2185,N_1984,N_2041);
nor U2186 (N_2186,N_1837,N_1992);
and U2187 (N_2187,N_1822,N_1916);
nor U2188 (N_2188,N_2095,N_2029);
and U2189 (N_2189,N_2007,N_1959);
xnor U2190 (N_2190,N_2033,N_1869);
or U2191 (N_2191,N_2070,N_2084);
xor U2192 (N_2192,N_1983,N_1977);
xnor U2193 (N_2193,N_1985,N_1949);
nand U2194 (N_2194,N_2088,N_2044);
nor U2195 (N_2195,N_1982,N_2053);
nand U2196 (N_2196,N_1930,N_1832);
xor U2197 (N_2197,N_2042,N_1811);
or U2198 (N_2198,N_1812,N_2094);
nand U2199 (N_2199,N_2066,N_1825);
nor U2200 (N_2200,N_1838,N_2022);
nor U2201 (N_2201,N_2004,N_2079);
and U2202 (N_2202,N_1882,N_2071);
nor U2203 (N_2203,N_2046,N_2091);
nor U2204 (N_2204,N_1986,N_1852);
or U2205 (N_2205,N_1958,N_1885);
nor U2206 (N_2206,N_1965,N_1850);
and U2207 (N_2207,N_2089,N_2001);
or U2208 (N_2208,N_1840,N_2000);
or U2209 (N_2209,N_1905,N_1951);
xor U2210 (N_2210,N_1952,N_1938);
nand U2211 (N_2211,N_1834,N_1929);
or U2212 (N_2212,N_2023,N_1902);
nand U2213 (N_2213,N_1871,N_2036);
and U2214 (N_2214,N_2014,N_2015);
nand U2215 (N_2215,N_1919,N_1923);
and U2216 (N_2216,N_1935,N_1862);
nor U2217 (N_2217,N_1920,N_1942);
xor U2218 (N_2218,N_1912,N_2058);
and U2219 (N_2219,N_1809,N_1875);
xor U2220 (N_2220,N_1870,N_1880);
nand U2221 (N_2221,N_1827,N_2076);
nor U2222 (N_2222,N_2087,N_2024);
xor U2223 (N_2223,N_1927,N_1826);
and U2224 (N_2224,N_1884,N_1804);
or U2225 (N_2225,N_1993,N_2057);
nand U2226 (N_2226,N_1980,N_1987);
nor U2227 (N_2227,N_2030,N_1917);
or U2228 (N_2228,N_1896,N_1863);
xor U2229 (N_2229,N_1967,N_1936);
nand U2230 (N_2230,N_1887,N_2061);
nor U2231 (N_2231,N_2081,N_2025);
and U2232 (N_2232,N_1996,N_1816);
nand U2233 (N_2233,N_1853,N_1979);
nand U2234 (N_2234,N_1995,N_2078);
and U2235 (N_2235,N_1848,N_1815);
nand U2236 (N_2236,N_1897,N_1821);
and U2237 (N_2237,N_1975,N_2062);
or U2238 (N_2238,N_1922,N_2026);
nor U2239 (N_2239,N_2040,N_2037);
nand U2240 (N_2240,N_1857,N_1964);
and U2241 (N_2241,N_2019,N_1823);
or U2242 (N_2242,N_1892,N_1931);
nand U2243 (N_2243,N_1873,N_1940);
nor U2244 (N_2244,N_2092,N_2073);
and U2245 (N_2245,N_1978,N_1818);
xnor U2246 (N_2246,N_1950,N_1820);
or U2247 (N_2247,N_1918,N_1937);
nand U2248 (N_2248,N_1932,N_1839);
xnor U2249 (N_2249,N_1891,N_1913);
xnor U2250 (N_2250,N_1904,N_2069);
and U2251 (N_2251,N_1955,N_1933);
and U2252 (N_2252,N_1925,N_1815);
nand U2253 (N_2253,N_2076,N_1982);
xnor U2254 (N_2254,N_2052,N_1973);
nor U2255 (N_2255,N_2083,N_1886);
and U2256 (N_2256,N_2078,N_2056);
xnor U2257 (N_2257,N_2038,N_1964);
or U2258 (N_2258,N_1852,N_1851);
and U2259 (N_2259,N_1838,N_1919);
xor U2260 (N_2260,N_1842,N_1847);
and U2261 (N_2261,N_1896,N_1988);
or U2262 (N_2262,N_1851,N_2099);
xnor U2263 (N_2263,N_1943,N_2007);
nor U2264 (N_2264,N_1867,N_1874);
or U2265 (N_2265,N_1958,N_2013);
xnor U2266 (N_2266,N_2052,N_2030);
nor U2267 (N_2267,N_1831,N_2056);
or U2268 (N_2268,N_1896,N_1932);
xnor U2269 (N_2269,N_2050,N_1926);
or U2270 (N_2270,N_1955,N_1897);
or U2271 (N_2271,N_1963,N_1966);
xnor U2272 (N_2272,N_2013,N_1818);
xnor U2273 (N_2273,N_1963,N_2027);
and U2274 (N_2274,N_1853,N_2031);
nor U2275 (N_2275,N_1828,N_1802);
nand U2276 (N_2276,N_1849,N_2035);
and U2277 (N_2277,N_2040,N_2082);
xnor U2278 (N_2278,N_2020,N_1849);
or U2279 (N_2279,N_2098,N_1856);
xor U2280 (N_2280,N_1852,N_1944);
and U2281 (N_2281,N_1982,N_2071);
xnor U2282 (N_2282,N_1870,N_2009);
nor U2283 (N_2283,N_2079,N_1921);
or U2284 (N_2284,N_2004,N_1967);
nand U2285 (N_2285,N_2064,N_2060);
and U2286 (N_2286,N_1990,N_1871);
xnor U2287 (N_2287,N_1867,N_1937);
nor U2288 (N_2288,N_2030,N_1870);
nor U2289 (N_2289,N_2054,N_1922);
or U2290 (N_2290,N_2026,N_1894);
xnor U2291 (N_2291,N_1928,N_2075);
nor U2292 (N_2292,N_1800,N_2032);
nand U2293 (N_2293,N_1911,N_1876);
nor U2294 (N_2294,N_1876,N_1934);
xnor U2295 (N_2295,N_1955,N_2073);
and U2296 (N_2296,N_2020,N_1915);
or U2297 (N_2297,N_1921,N_1893);
and U2298 (N_2298,N_1974,N_1894);
and U2299 (N_2299,N_1827,N_1947);
xnor U2300 (N_2300,N_1877,N_1914);
nor U2301 (N_2301,N_2015,N_1962);
and U2302 (N_2302,N_1915,N_1865);
xor U2303 (N_2303,N_1973,N_1919);
nand U2304 (N_2304,N_1907,N_1817);
and U2305 (N_2305,N_1891,N_2013);
nor U2306 (N_2306,N_1807,N_2000);
and U2307 (N_2307,N_1937,N_1993);
nor U2308 (N_2308,N_1946,N_1819);
nand U2309 (N_2309,N_2099,N_1974);
nor U2310 (N_2310,N_1849,N_1932);
nand U2311 (N_2311,N_1891,N_1809);
xnor U2312 (N_2312,N_1890,N_1905);
or U2313 (N_2313,N_1973,N_1906);
nor U2314 (N_2314,N_1822,N_1805);
xor U2315 (N_2315,N_2062,N_1894);
nand U2316 (N_2316,N_1929,N_1951);
xnor U2317 (N_2317,N_1930,N_1974);
xor U2318 (N_2318,N_1878,N_1976);
or U2319 (N_2319,N_1878,N_1951);
or U2320 (N_2320,N_1836,N_1989);
xor U2321 (N_2321,N_1817,N_2053);
nand U2322 (N_2322,N_1937,N_2037);
nor U2323 (N_2323,N_1882,N_1948);
and U2324 (N_2324,N_2010,N_2044);
and U2325 (N_2325,N_2018,N_1863);
nand U2326 (N_2326,N_2026,N_1984);
or U2327 (N_2327,N_2095,N_2081);
nand U2328 (N_2328,N_2037,N_2026);
and U2329 (N_2329,N_1905,N_1909);
xnor U2330 (N_2330,N_2033,N_1934);
xnor U2331 (N_2331,N_1994,N_1914);
nor U2332 (N_2332,N_1882,N_2074);
xor U2333 (N_2333,N_2035,N_1800);
nor U2334 (N_2334,N_1820,N_1838);
or U2335 (N_2335,N_1993,N_2032);
nand U2336 (N_2336,N_1927,N_2038);
or U2337 (N_2337,N_2071,N_1986);
nor U2338 (N_2338,N_1836,N_1903);
and U2339 (N_2339,N_1852,N_1952);
and U2340 (N_2340,N_2036,N_2095);
nor U2341 (N_2341,N_1870,N_1837);
or U2342 (N_2342,N_2073,N_2077);
xor U2343 (N_2343,N_2016,N_1854);
nand U2344 (N_2344,N_2098,N_1857);
or U2345 (N_2345,N_1891,N_1894);
xnor U2346 (N_2346,N_1999,N_1931);
xor U2347 (N_2347,N_1904,N_1979);
nor U2348 (N_2348,N_1993,N_1826);
and U2349 (N_2349,N_2041,N_2009);
or U2350 (N_2350,N_1820,N_2090);
or U2351 (N_2351,N_1937,N_2061);
or U2352 (N_2352,N_1937,N_1899);
nand U2353 (N_2353,N_2052,N_1988);
xnor U2354 (N_2354,N_1907,N_2030);
nor U2355 (N_2355,N_1995,N_2041);
and U2356 (N_2356,N_1916,N_1990);
nand U2357 (N_2357,N_1929,N_2063);
or U2358 (N_2358,N_1825,N_2003);
or U2359 (N_2359,N_1948,N_1890);
xnor U2360 (N_2360,N_1948,N_1942);
or U2361 (N_2361,N_1997,N_1905);
nor U2362 (N_2362,N_2035,N_1917);
or U2363 (N_2363,N_2077,N_1954);
or U2364 (N_2364,N_1821,N_1822);
or U2365 (N_2365,N_1856,N_2047);
nor U2366 (N_2366,N_1964,N_1914);
nand U2367 (N_2367,N_1869,N_1976);
nand U2368 (N_2368,N_2008,N_1865);
nor U2369 (N_2369,N_1864,N_1883);
or U2370 (N_2370,N_2076,N_1824);
or U2371 (N_2371,N_2005,N_1853);
or U2372 (N_2372,N_1976,N_1973);
and U2373 (N_2373,N_2079,N_1929);
and U2374 (N_2374,N_2071,N_1893);
and U2375 (N_2375,N_2050,N_2061);
and U2376 (N_2376,N_1981,N_1940);
xor U2377 (N_2377,N_1800,N_1999);
nand U2378 (N_2378,N_1910,N_2058);
xnor U2379 (N_2379,N_1828,N_2099);
nor U2380 (N_2380,N_1922,N_1974);
nand U2381 (N_2381,N_1918,N_2057);
and U2382 (N_2382,N_1897,N_1861);
or U2383 (N_2383,N_1876,N_1924);
or U2384 (N_2384,N_2087,N_1910);
and U2385 (N_2385,N_1812,N_2061);
nand U2386 (N_2386,N_2009,N_1902);
xnor U2387 (N_2387,N_1840,N_2084);
and U2388 (N_2388,N_1807,N_2066);
nand U2389 (N_2389,N_2081,N_1948);
xor U2390 (N_2390,N_2097,N_1988);
xnor U2391 (N_2391,N_1859,N_1923);
or U2392 (N_2392,N_2021,N_2046);
and U2393 (N_2393,N_1886,N_1869);
nor U2394 (N_2394,N_1855,N_1915);
or U2395 (N_2395,N_1820,N_2027);
nand U2396 (N_2396,N_1878,N_1891);
and U2397 (N_2397,N_1990,N_1810);
xnor U2398 (N_2398,N_1821,N_1814);
and U2399 (N_2399,N_1840,N_2005);
nand U2400 (N_2400,N_2351,N_2101);
nand U2401 (N_2401,N_2138,N_2185);
nand U2402 (N_2402,N_2366,N_2261);
and U2403 (N_2403,N_2197,N_2106);
and U2404 (N_2404,N_2136,N_2223);
nor U2405 (N_2405,N_2196,N_2380);
and U2406 (N_2406,N_2111,N_2354);
and U2407 (N_2407,N_2158,N_2392);
xor U2408 (N_2408,N_2234,N_2239);
or U2409 (N_2409,N_2144,N_2263);
nand U2410 (N_2410,N_2266,N_2168);
nand U2411 (N_2411,N_2246,N_2332);
nor U2412 (N_2412,N_2133,N_2167);
xnor U2413 (N_2413,N_2273,N_2140);
or U2414 (N_2414,N_2375,N_2237);
nand U2415 (N_2415,N_2328,N_2200);
xnor U2416 (N_2416,N_2291,N_2290);
xor U2417 (N_2417,N_2125,N_2303);
and U2418 (N_2418,N_2206,N_2336);
xnor U2419 (N_2419,N_2177,N_2378);
and U2420 (N_2420,N_2151,N_2281);
and U2421 (N_2421,N_2107,N_2365);
and U2422 (N_2422,N_2146,N_2199);
nor U2423 (N_2423,N_2319,N_2219);
or U2424 (N_2424,N_2267,N_2343);
nor U2425 (N_2425,N_2265,N_2118);
and U2426 (N_2426,N_2306,N_2318);
xnor U2427 (N_2427,N_2211,N_2156);
and U2428 (N_2428,N_2189,N_2307);
xor U2429 (N_2429,N_2141,N_2396);
nor U2430 (N_2430,N_2322,N_2201);
and U2431 (N_2431,N_2297,N_2180);
nor U2432 (N_2432,N_2342,N_2169);
and U2433 (N_2433,N_2245,N_2347);
or U2434 (N_2434,N_2228,N_2313);
xor U2435 (N_2435,N_2293,N_2383);
xnor U2436 (N_2436,N_2345,N_2119);
xor U2437 (N_2437,N_2126,N_2262);
nor U2438 (N_2438,N_2305,N_2213);
and U2439 (N_2439,N_2357,N_2353);
or U2440 (N_2440,N_2127,N_2268);
and U2441 (N_2441,N_2372,N_2391);
xnor U2442 (N_2442,N_2230,N_2277);
and U2443 (N_2443,N_2362,N_2376);
xnor U2444 (N_2444,N_2202,N_2320);
nor U2445 (N_2445,N_2386,N_2339);
xnor U2446 (N_2446,N_2282,N_2183);
nor U2447 (N_2447,N_2166,N_2257);
nand U2448 (N_2448,N_2373,N_2165);
or U2449 (N_2449,N_2130,N_2374);
xor U2450 (N_2450,N_2109,N_2317);
nand U2451 (N_2451,N_2278,N_2143);
nor U2452 (N_2452,N_2215,N_2224);
nand U2453 (N_2453,N_2135,N_2231);
or U2454 (N_2454,N_2292,N_2232);
nor U2455 (N_2455,N_2112,N_2186);
and U2456 (N_2456,N_2218,N_2210);
or U2457 (N_2457,N_2280,N_2304);
nor U2458 (N_2458,N_2175,N_2123);
or U2459 (N_2459,N_2301,N_2134);
nand U2460 (N_2460,N_2300,N_2128);
or U2461 (N_2461,N_2371,N_2203);
xnor U2462 (N_2462,N_2236,N_2172);
nor U2463 (N_2463,N_2251,N_2275);
nand U2464 (N_2464,N_2227,N_2395);
and U2465 (N_2465,N_2338,N_2149);
and U2466 (N_2466,N_2387,N_2335);
nor U2467 (N_2467,N_2152,N_2212);
xor U2468 (N_2468,N_2367,N_2187);
nand U2469 (N_2469,N_2244,N_2360);
and U2470 (N_2470,N_2184,N_2247);
or U2471 (N_2471,N_2285,N_2220);
xnor U2472 (N_2472,N_2173,N_2270);
nand U2473 (N_2473,N_2302,N_2346);
nor U2474 (N_2474,N_2121,N_2358);
nor U2475 (N_2475,N_2364,N_2209);
or U2476 (N_2476,N_2154,N_2340);
xnor U2477 (N_2477,N_2296,N_2384);
nand U2478 (N_2478,N_2115,N_2284);
and U2479 (N_2479,N_2299,N_2221);
nand U2480 (N_2480,N_2204,N_2195);
nor U2481 (N_2481,N_2164,N_2113);
nor U2482 (N_2482,N_2238,N_2258);
xor U2483 (N_2483,N_2329,N_2207);
xnor U2484 (N_2484,N_2259,N_2192);
nor U2485 (N_2485,N_2120,N_2361);
and U2486 (N_2486,N_2235,N_2389);
xnor U2487 (N_2487,N_2170,N_2142);
nand U2488 (N_2488,N_2225,N_2311);
or U2489 (N_2489,N_2214,N_2148);
nor U2490 (N_2490,N_2162,N_2363);
nor U2491 (N_2491,N_2163,N_2161);
nand U2492 (N_2492,N_2334,N_2131);
nand U2493 (N_2493,N_2388,N_2205);
xor U2494 (N_2494,N_2287,N_2254);
or U2495 (N_2495,N_2139,N_2153);
xor U2496 (N_2496,N_2321,N_2348);
and U2497 (N_2497,N_2325,N_2255);
xnor U2498 (N_2498,N_2276,N_2355);
xor U2499 (N_2499,N_2132,N_2289);
nand U2500 (N_2500,N_2344,N_2331);
xor U2501 (N_2501,N_2264,N_2124);
nor U2502 (N_2502,N_2310,N_2381);
xor U2503 (N_2503,N_2271,N_2190);
xnor U2504 (N_2504,N_2324,N_2250);
nor U2505 (N_2505,N_2145,N_2368);
xnor U2506 (N_2506,N_2191,N_2102);
xor U2507 (N_2507,N_2178,N_2352);
xnor U2508 (N_2508,N_2316,N_2253);
nand U2509 (N_2509,N_2100,N_2286);
nand U2510 (N_2510,N_2110,N_2308);
nor U2511 (N_2511,N_2315,N_2114);
nor U2512 (N_2512,N_2176,N_2117);
xor U2513 (N_2513,N_2159,N_2382);
nand U2514 (N_2514,N_2260,N_2150);
xor U2515 (N_2515,N_2103,N_2198);
and U2516 (N_2516,N_2279,N_2229);
or U2517 (N_2517,N_2249,N_2327);
or U2518 (N_2518,N_2104,N_2397);
and U2519 (N_2519,N_2147,N_2314);
or U2520 (N_2520,N_2349,N_2194);
nand U2521 (N_2521,N_2122,N_2393);
nand U2522 (N_2522,N_2359,N_2274);
xor U2523 (N_2523,N_2193,N_2252);
nor U2524 (N_2524,N_2160,N_2269);
nor U2525 (N_2525,N_2243,N_2295);
and U2526 (N_2526,N_2226,N_2155);
nor U2527 (N_2527,N_2171,N_2216);
and U2528 (N_2528,N_2323,N_2182);
and U2529 (N_2529,N_2129,N_2174);
or U2530 (N_2530,N_2379,N_2248);
nor U2531 (N_2531,N_2242,N_2377);
xor U2532 (N_2532,N_2333,N_2385);
and U2533 (N_2533,N_2241,N_2108);
nor U2534 (N_2534,N_2233,N_2341);
nand U2535 (N_2535,N_2350,N_2116);
or U2536 (N_2536,N_2294,N_2309);
or U2537 (N_2537,N_2398,N_2188);
or U2538 (N_2538,N_2181,N_2370);
xor U2539 (N_2539,N_2356,N_2179);
and U2540 (N_2540,N_2288,N_2240);
nor U2541 (N_2541,N_2369,N_2157);
nor U2542 (N_2542,N_2330,N_2222);
nor U2543 (N_2543,N_2337,N_2394);
xnor U2544 (N_2544,N_2217,N_2272);
and U2545 (N_2545,N_2208,N_2312);
or U2546 (N_2546,N_2390,N_2256);
xor U2547 (N_2547,N_2137,N_2298);
xnor U2548 (N_2548,N_2283,N_2399);
or U2549 (N_2549,N_2326,N_2105);
xor U2550 (N_2550,N_2346,N_2106);
or U2551 (N_2551,N_2119,N_2299);
or U2552 (N_2552,N_2368,N_2385);
and U2553 (N_2553,N_2199,N_2204);
nand U2554 (N_2554,N_2294,N_2325);
xnor U2555 (N_2555,N_2189,N_2335);
xor U2556 (N_2556,N_2193,N_2200);
xor U2557 (N_2557,N_2362,N_2254);
and U2558 (N_2558,N_2110,N_2237);
nand U2559 (N_2559,N_2227,N_2350);
nand U2560 (N_2560,N_2219,N_2224);
xor U2561 (N_2561,N_2271,N_2129);
nor U2562 (N_2562,N_2397,N_2194);
and U2563 (N_2563,N_2255,N_2292);
and U2564 (N_2564,N_2129,N_2330);
xor U2565 (N_2565,N_2341,N_2180);
and U2566 (N_2566,N_2220,N_2175);
xnor U2567 (N_2567,N_2197,N_2186);
or U2568 (N_2568,N_2115,N_2136);
or U2569 (N_2569,N_2393,N_2133);
nor U2570 (N_2570,N_2262,N_2341);
and U2571 (N_2571,N_2266,N_2177);
and U2572 (N_2572,N_2288,N_2352);
nand U2573 (N_2573,N_2239,N_2198);
or U2574 (N_2574,N_2270,N_2137);
nor U2575 (N_2575,N_2310,N_2151);
xnor U2576 (N_2576,N_2231,N_2255);
nor U2577 (N_2577,N_2308,N_2318);
nor U2578 (N_2578,N_2103,N_2205);
or U2579 (N_2579,N_2324,N_2395);
or U2580 (N_2580,N_2347,N_2289);
or U2581 (N_2581,N_2153,N_2149);
and U2582 (N_2582,N_2153,N_2163);
and U2583 (N_2583,N_2271,N_2119);
nand U2584 (N_2584,N_2305,N_2210);
and U2585 (N_2585,N_2386,N_2337);
nand U2586 (N_2586,N_2156,N_2260);
or U2587 (N_2587,N_2107,N_2227);
and U2588 (N_2588,N_2263,N_2372);
or U2589 (N_2589,N_2264,N_2260);
xor U2590 (N_2590,N_2130,N_2174);
xor U2591 (N_2591,N_2117,N_2216);
nand U2592 (N_2592,N_2283,N_2208);
nor U2593 (N_2593,N_2132,N_2393);
xnor U2594 (N_2594,N_2312,N_2190);
and U2595 (N_2595,N_2348,N_2187);
or U2596 (N_2596,N_2302,N_2399);
xor U2597 (N_2597,N_2231,N_2109);
nand U2598 (N_2598,N_2388,N_2394);
nand U2599 (N_2599,N_2306,N_2158);
nand U2600 (N_2600,N_2144,N_2300);
and U2601 (N_2601,N_2394,N_2233);
or U2602 (N_2602,N_2204,N_2125);
or U2603 (N_2603,N_2324,N_2138);
nand U2604 (N_2604,N_2127,N_2303);
xnor U2605 (N_2605,N_2130,N_2206);
xor U2606 (N_2606,N_2393,N_2359);
xor U2607 (N_2607,N_2255,N_2383);
nand U2608 (N_2608,N_2248,N_2195);
nor U2609 (N_2609,N_2210,N_2362);
nor U2610 (N_2610,N_2327,N_2321);
xnor U2611 (N_2611,N_2240,N_2168);
and U2612 (N_2612,N_2388,N_2191);
xnor U2613 (N_2613,N_2396,N_2229);
nor U2614 (N_2614,N_2200,N_2353);
xnor U2615 (N_2615,N_2303,N_2193);
nand U2616 (N_2616,N_2153,N_2337);
and U2617 (N_2617,N_2194,N_2362);
xnor U2618 (N_2618,N_2101,N_2301);
nor U2619 (N_2619,N_2327,N_2132);
nand U2620 (N_2620,N_2244,N_2270);
and U2621 (N_2621,N_2363,N_2352);
xor U2622 (N_2622,N_2133,N_2125);
xor U2623 (N_2623,N_2339,N_2245);
nor U2624 (N_2624,N_2278,N_2233);
and U2625 (N_2625,N_2394,N_2308);
nand U2626 (N_2626,N_2239,N_2126);
and U2627 (N_2627,N_2333,N_2167);
or U2628 (N_2628,N_2388,N_2274);
and U2629 (N_2629,N_2195,N_2290);
and U2630 (N_2630,N_2322,N_2368);
nor U2631 (N_2631,N_2192,N_2309);
nand U2632 (N_2632,N_2187,N_2155);
nand U2633 (N_2633,N_2238,N_2151);
xnor U2634 (N_2634,N_2100,N_2157);
nand U2635 (N_2635,N_2233,N_2389);
or U2636 (N_2636,N_2391,N_2379);
nand U2637 (N_2637,N_2189,N_2331);
nor U2638 (N_2638,N_2382,N_2363);
or U2639 (N_2639,N_2203,N_2273);
or U2640 (N_2640,N_2239,N_2135);
nand U2641 (N_2641,N_2393,N_2171);
nor U2642 (N_2642,N_2318,N_2352);
nor U2643 (N_2643,N_2174,N_2182);
xnor U2644 (N_2644,N_2280,N_2179);
nand U2645 (N_2645,N_2271,N_2286);
nor U2646 (N_2646,N_2321,N_2267);
xor U2647 (N_2647,N_2130,N_2275);
nor U2648 (N_2648,N_2312,N_2211);
nor U2649 (N_2649,N_2383,N_2263);
or U2650 (N_2650,N_2315,N_2344);
xor U2651 (N_2651,N_2156,N_2107);
or U2652 (N_2652,N_2153,N_2306);
and U2653 (N_2653,N_2310,N_2317);
nand U2654 (N_2654,N_2356,N_2219);
xor U2655 (N_2655,N_2188,N_2331);
nand U2656 (N_2656,N_2155,N_2211);
nand U2657 (N_2657,N_2101,N_2299);
nand U2658 (N_2658,N_2131,N_2101);
nand U2659 (N_2659,N_2340,N_2383);
nor U2660 (N_2660,N_2202,N_2342);
xor U2661 (N_2661,N_2260,N_2396);
nor U2662 (N_2662,N_2262,N_2387);
xor U2663 (N_2663,N_2179,N_2297);
nand U2664 (N_2664,N_2275,N_2231);
xor U2665 (N_2665,N_2197,N_2385);
nor U2666 (N_2666,N_2181,N_2122);
and U2667 (N_2667,N_2383,N_2177);
nand U2668 (N_2668,N_2280,N_2282);
nand U2669 (N_2669,N_2228,N_2136);
nor U2670 (N_2670,N_2352,N_2218);
and U2671 (N_2671,N_2223,N_2227);
and U2672 (N_2672,N_2201,N_2117);
nor U2673 (N_2673,N_2220,N_2246);
nand U2674 (N_2674,N_2226,N_2216);
xnor U2675 (N_2675,N_2211,N_2202);
xnor U2676 (N_2676,N_2138,N_2104);
nor U2677 (N_2677,N_2146,N_2106);
or U2678 (N_2678,N_2372,N_2262);
and U2679 (N_2679,N_2155,N_2186);
nor U2680 (N_2680,N_2166,N_2331);
or U2681 (N_2681,N_2268,N_2273);
and U2682 (N_2682,N_2319,N_2273);
nand U2683 (N_2683,N_2370,N_2199);
xnor U2684 (N_2684,N_2152,N_2240);
xor U2685 (N_2685,N_2339,N_2338);
nor U2686 (N_2686,N_2317,N_2359);
or U2687 (N_2687,N_2128,N_2396);
nand U2688 (N_2688,N_2202,N_2253);
or U2689 (N_2689,N_2343,N_2350);
nand U2690 (N_2690,N_2295,N_2298);
and U2691 (N_2691,N_2154,N_2331);
and U2692 (N_2692,N_2280,N_2129);
or U2693 (N_2693,N_2244,N_2346);
nand U2694 (N_2694,N_2215,N_2151);
nor U2695 (N_2695,N_2307,N_2298);
or U2696 (N_2696,N_2216,N_2368);
or U2697 (N_2697,N_2299,N_2386);
nand U2698 (N_2698,N_2141,N_2372);
and U2699 (N_2699,N_2116,N_2182);
and U2700 (N_2700,N_2415,N_2662);
nand U2701 (N_2701,N_2539,N_2444);
nor U2702 (N_2702,N_2660,N_2499);
or U2703 (N_2703,N_2431,N_2677);
or U2704 (N_2704,N_2401,N_2656);
xor U2705 (N_2705,N_2652,N_2436);
xnor U2706 (N_2706,N_2519,N_2681);
or U2707 (N_2707,N_2558,N_2636);
xor U2708 (N_2708,N_2560,N_2615);
nand U2709 (N_2709,N_2628,N_2573);
xnor U2710 (N_2710,N_2638,N_2692);
nor U2711 (N_2711,N_2508,N_2459);
nor U2712 (N_2712,N_2440,N_2445);
xnor U2713 (N_2713,N_2470,N_2498);
or U2714 (N_2714,N_2654,N_2613);
nand U2715 (N_2715,N_2507,N_2490);
and U2716 (N_2716,N_2663,N_2515);
xor U2717 (N_2717,N_2512,N_2647);
nor U2718 (N_2718,N_2630,N_2481);
xor U2719 (N_2719,N_2426,N_2501);
nor U2720 (N_2720,N_2581,N_2469);
nand U2721 (N_2721,N_2411,N_2588);
and U2722 (N_2722,N_2535,N_2649);
or U2723 (N_2723,N_2443,N_2489);
nor U2724 (N_2724,N_2653,N_2509);
xnor U2725 (N_2725,N_2477,N_2658);
or U2726 (N_2726,N_2450,N_2479);
xor U2727 (N_2727,N_2424,N_2529);
xnor U2728 (N_2728,N_2453,N_2597);
xor U2729 (N_2729,N_2549,N_2641);
nor U2730 (N_2730,N_2563,N_2464);
nor U2731 (N_2731,N_2448,N_2403);
nand U2732 (N_2732,N_2593,N_2527);
or U2733 (N_2733,N_2603,N_2579);
nand U2734 (N_2734,N_2585,N_2446);
and U2735 (N_2735,N_2689,N_2428);
nor U2736 (N_2736,N_2609,N_2659);
and U2737 (N_2737,N_2602,N_2556);
nor U2738 (N_2738,N_2548,N_2550);
or U2739 (N_2739,N_2666,N_2574);
nor U2740 (N_2740,N_2472,N_2571);
xnor U2741 (N_2741,N_2665,N_2610);
nand U2742 (N_2742,N_2577,N_2427);
and U2743 (N_2743,N_2668,N_2463);
xnor U2744 (N_2744,N_2678,N_2420);
nor U2745 (N_2745,N_2644,N_2657);
nor U2746 (N_2746,N_2449,N_2456);
nor U2747 (N_2747,N_2570,N_2514);
xnor U2748 (N_2748,N_2538,N_2651);
or U2749 (N_2749,N_2698,N_2505);
nand U2750 (N_2750,N_2604,N_2475);
xor U2751 (N_2751,N_2451,N_2540);
or U2752 (N_2752,N_2695,N_2642);
nor U2753 (N_2753,N_2435,N_2575);
or U2754 (N_2754,N_2466,N_2525);
nor U2755 (N_2755,N_2438,N_2670);
and U2756 (N_2756,N_2618,N_2530);
or U2757 (N_2757,N_2608,N_2655);
nand U2758 (N_2758,N_2639,N_2410);
nor U2759 (N_2759,N_2684,N_2646);
or U2760 (N_2760,N_2640,N_2569);
xnor U2761 (N_2761,N_2605,N_2524);
nor U2762 (N_2762,N_2686,N_2416);
nor U2763 (N_2763,N_2633,N_2476);
xor U2764 (N_2764,N_2429,N_2637);
nor U2765 (N_2765,N_2617,N_2546);
or U2766 (N_2766,N_2664,N_2425);
and U2767 (N_2767,N_2598,N_2611);
xor U2768 (N_2768,N_2582,N_2408);
nand U2769 (N_2769,N_2553,N_2528);
or U2770 (N_2770,N_2567,N_2554);
xnor U2771 (N_2771,N_2502,N_2627);
and U2772 (N_2772,N_2417,N_2442);
and U2773 (N_2773,N_2612,N_2454);
and U2774 (N_2774,N_2566,N_2537);
and U2775 (N_2775,N_2418,N_2606);
and U2776 (N_2776,N_2441,N_2688);
and U2777 (N_2777,N_2500,N_2552);
nor U2778 (N_2778,N_2691,N_2675);
or U2779 (N_2779,N_2584,N_2591);
xnor U2780 (N_2780,N_2572,N_2600);
or U2781 (N_2781,N_2690,N_2685);
xnor U2782 (N_2782,N_2619,N_2473);
and U2783 (N_2783,N_2545,N_2465);
xor U2784 (N_2784,N_2496,N_2467);
and U2785 (N_2785,N_2557,N_2414);
or U2786 (N_2786,N_2580,N_2419);
xor U2787 (N_2787,N_2493,N_2457);
and U2788 (N_2788,N_2504,N_2517);
xnor U2789 (N_2789,N_2632,N_2626);
and U2790 (N_2790,N_2421,N_2541);
nand U2791 (N_2791,N_2621,N_2562);
xnor U2792 (N_2792,N_2650,N_2516);
nand U2793 (N_2793,N_2699,N_2595);
or U2794 (N_2794,N_2521,N_2596);
and U2795 (N_2795,N_2634,N_2526);
nand U2796 (N_2796,N_2543,N_2648);
or U2797 (N_2797,N_2682,N_2486);
xor U2798 (N_2798,N_2452,N_2506);
and U2799 (N_2799,N_2680,N_2511);
xor U2800 (N_2800,N_2484,N_2439);
and U2801 (N_2801,N_2536,N_2400);
and U2802 (N_2802,N_2482,N_2462);
nor U2803 (N_2803,N_2518,N_2405);
nand U2804 (N_2804,N_2643,N_2561);
or U2805 (N_2805,N_2565,N_2673);
or U2806 (N_2806,N_2513,N_2487);
and U2807 (N_2807,N_2607,N_2503);
and U2808 (N_2808,N_2474,N_2614);
nand U2809 (N_2809,N_2413,N_2460);
xnor U2810 (N_2810,N_2471,N_2461);
nor U2811 (N_2811,N_2667,N_2622);
xor U2812 (N_2812,N_2583,N_2423);
and U2813 (N_2813,N_2551,N_2693);
and U2814 (N_2814,N_2679,N_2629);
xor U2815 (N_2815,N_2576,N_2531);
xnor U2816 (N_2816,N_2491,N_2671);
and U2817 (N_2817,N_2555,N_2495);
nor U2818 (N_2818,N_2586,N_2631);
or U2819 (N_2819,N_2432,N_2404);
and U2820 (N_2820,N_2601,N_2485);
or U2821 (N_2821,N_2625,N_2589);
or U2822 (N_2822,N_2520,N_2623);
nand U2823 (N_2823,N_2587,N_2694);
and U2824 (N_2824,N_2468,N_2624);
or U2825 (N_2825,N_2409,N_2559);
nor U2826 (N_2826,N_2687,N_2455);
xor U2827 (N_2827,N_2532,N_2533);
and U2828 (N_2828,N_2433,N_2661);
or U2829 (N_2829,N_2447,N_2592);
or U2830 (N_2830,N_2497,N_2406);
and U2831 (N_2831,N_2458,N_2616);
nor U2832 (N_2832,N_2483,N_2696);
xor U2833 (N_2833,N_2645,N_2488);
and U2834 (N_2834,N_2534,N_2674);
xnor U2835 (N_2835,N_2412,N_2547);
nor U2836 (N_2836,N_2494,N_2599);
or U2837 (N_2837,N_2407,N_2542);
or U2838 (N_2838,N_2510,N_2523);
nor U2839 (N_2839,N_2568,N_2478);
xor U2840 (N_2840,N_2564,N_2683);
nor U2841 (N_2841,N_2672,N_2522);
nand U2842 (N_2842,N_2635,N_2480);
nor U2843 (N_2843,N_2594,N_2697);
nor U2844 (N_2844,N_2676,N_2590);
nand U2845 (N_2845,N_2492,N_2620);
xnor U2846 (N_2846,N_2430,N_2402);
or U2847 (N_2847,N_2544,N_2437);
and U2848 (N_2848,N_2578,N_2434);
nand U2849 (N_2849,N_2669,N_2422);
nor U2850 (N_2850,N_2621,N_2532);
nand U2851 (N_2851,N_2569,N_2570);
nor U2852 (N_2852,N_2533,N_2619);
and U2853 (N_2853,N_2567,N_2621);
nor U2854 (N_2854,N_2575,N_2592);
or U2855 (N_2855,N_2546,N_2539);
xor U2856 (N_2856,N_2683,N_2403);
xnor U2857 (N_2857,N_2510,N_2644);
xnor U2858 (N_2858,N_2656,N_2605);
nor U2859 (N_2859,N_2462,N_2467);
or U2860 (N_2860,N_2678,N_2628);
and U2861 (N_2861,N_2616,N_2499);
or U2862 (N_2862,N_2402,N_2560);
nor U2863 (N_2863,N_2635,N_2572);
xor U2864 (N_2864,N_2632,N_2404);
or U2865 (N_2865,N_2523,N_2475);
xor U2866 (N_2866,N_2649,N_2642);
nor U2867 (N_2867,N_2653,N_2446);
nor U2868 (N_2868,N_2692,N_2627);
and U2869 (N_2869,N_2656,N_2647);
nor U2870 (N_2870,N_2473,N_2439);
nand U2871 (N_2871,N_2438,N_2635);
nand U2872 (N_2872,N_2554,N_2529);
xnor U2873 (N_2873,N_2650,N_2644);
nor U2874 (N_2874,N_2692,N_2504);
or U2875 (N_2875,N_2698,N_2484);
and U2876 (N_2876,N_2589,N_2630);
xor U2877 (N_2877,N_2453,N_2443);
nand U2878 (N_2878,N_2609,N_2603);
xor U2879 (N_2879,N_2686,N_2600);
and U2880 (N_2880,N_2501,N_2676);
and U2881 (N_2881,N_2652,N_2570);
and U2882 (N_2882,N_2514,N_2530);
nand U2883 (N_2883,N_2539,N_2555);
nand U2884 (N_2884,N_2503,N_2629);
xor U2885 (N_2885,N_2489,N_2591);
xnor U2886 (N_2886,N_2536,N_2452);
xnor U2887 (N_2887,N_2626,N_2406);
and U2888 (N_2888,N_2639,N_2510);
or U2889 (N_2889,N_2617,N_2525);
xnor U2890 (N_2890,N_2587,N_2675);
nor U2891 (N_2891,N_2525,N_2689);
nor U2892 (N_2892,N_2514,N_2451);
nor U2893 (N_2893,N_2693,N_2414);
nor U2894 (N_2894,N_2554,N_2558);
nor U2895 (N_2895,N_2407,N_2527);
xnor U2896 (N_2896,N_2544,N_2418);
and U2897 (N_2897,N_2401,N_2437);
nor U2898 (N_2898,N_2452,N_2478);
nor U2899 (N_2899,N_2687,N_2546);
xnor U2900 (N_2900,N_2492,N_2630);
or U2901 (N_2901,N_2591,N_2412);
nor U2902 (N_2902,N_2630,N_2433);
nand U2903 (N_2903,N_2581,N_2570);
nor U2904 (N_2904,N_2672,N_2634);
nor U2905 (N_2905,N_2678,N_2435);
nand U2906 (N_2906,N_2651,N_2691);
xnor U2907 (N_2907,N_2612,N_2697);
nor U2908 (N_2908,N_2652,N_2596);
nor U2909 (N_2909,N_2505,N_2476);
xor U2910 (N_2910,N_2674,N_2411);
or U2911 (N_2911,N_2499,N_2575);
and U2912 (N_2912,N_2554,N_2615);
nor U2913 (N_2913,N_2690,N_2411);
nor U2914 (N_2914,N_2485,N_2407);
nor U2915 (N_2915,N_2512,N_2597);
or U2916 (N_2916,N_2416,N_2586);
nand U2917 (N_2917,N_2559,N_2600);
xor U2918 (N_2918,N_2538,N_2549);
and U2919 (N_2919,N_2444,N_2583);
nor U2920 (N_2920,N_2503,N_2417);
xnor U2921 (N_2921,N_2489,N_2604);
xnor U2922 (N_2922,N_2421,N_2609);
xor U2923 (N_2923,N_2464,N_2415);
or U2924 (N_2924,N_2470,N_2571);
nand U2925 (N_2925,N_2628,N_2597);
xor U2926 (N_2926,N_2405,N_2657);
and U2927 (N_2927,N_2547,N_2486);
nor U2928 (N_2928,N_2427,N_2559);
nand U2929 (N_2929,N_2637,N_2677);
nor U2930 (N_2930,N_2672,N_2631);
nand U2931 (N_2931,N_2668,N_2640);
or U2932 (N_2932,N_2612,N_2447);
and U2933 (N_2933,N_2665,N_2550);
nor U2934 (N_2934,N_2587,N_2595);
or U2935 (N_2935,N_2466,N_2539);
or U2936 (N_2936,N_2421,N_2439);
nor U2937 (N_2937,N_2618,N_2466);
and U2938 (N_2938,N_2454,N_2592);
nor U2939 (N_2939,N_2430,N_2445);
nand U2940 (N_2940,N_2574,N_2566);
nand U2941 (N_2941,N_2597,N_2440);
xor U2942 (N_2942,N_2569,N_2656);
xnor U2943 (N_2943,N_2663,N_2673);
xnor U2944 (N_2944,N_2623,N_2459);
or U2945 (N_2945,N_2513,N_2416);
or U2946 (N_2946,N_2694,N_2612);
nand U2947 (N_2947,N_2689,N_2698);
nand U2948 (N_2948,N_2422,N_2454);
xor U2949 (N_2949,N_2482,N_2555);
xnor U2950 (N_2950,N_2517,N_2515);
and U2951 (N_2951,N_2462,N_2589);
nand U2952 (N_2952,N_2479,N_2579);
xor U2953 (N_2953,N_2596,N_2590);
nor U2954 (N_2954,N_2446,N_2654);
nand U2955 (N_2955,N_2466,N_2547);
nand U2956 (N_2956,N_2471,N_2505);
nand U2957 (N_2957,N_2496,N_2581);
and U2958 (N_2958,N_2471,N_2500);
and U2959 (N_2959,N_2582,N_2478);
xor U2960 (N_2960,N_2618,N_2465);
xnor U2961 (N_2961,N_2500,N_2567);
xor U2962 (N_2962,N_2597,N_2621);
nor U2963 (N_2963,N_2695,N_2488);
or U2964 (N_2964,N_2690,N_2501);
or U2965 (N_2965,N_2613,N_2421);
or U2966 (N_2966,N_2556,N_2686);
nand U2967 (N_2967,N_2554,N_2638);
or U2968 (N_2968,N_2428,N_2651);
nand U2969 (N_2969,N_2543,N_2482);
and U2970 (N_2970,N_2446,N_2657);
or U2971 (N_2971,N_2619,N_2464);
xor U2972 (N_2972,N_2415,N_2677);
xor U2973 (N_2973,N_2692,N_2678);
nor U2974 (N_2974,N_2407,N_2457);
and U2975 (N_2975,N_2563,N_2594);
nand U2976 (N_2976,N_2427,N_2525);
xor U2977 (N_2977,N_2416,N_2564);
xnor U2978 (N_2978,N_2430,N_2535);
xnor U2979 (N_2979,N_2514,N_2681);
and U2980 (N_2980,N_2590,N_2607);
xnor U2981 (N_2981,N_2600,N_2555);
nor U2982 (N_2982,N_2627,N_2653);
nor U2983 (N_2983,N_2481,N_2636);
and U2984 (N_2984,N_2661,N_2482);
xnor U2985 (N_2985,N_2543,N_2468);
or U2986 (N_2986,N_2693,N_2576);
nand U2987 (N_2987,N_2484,N_2471);
nand U2988 (N_2988,N_2454,N_2581);
xnor U2989 (N_2989,N_2660,N_2592);
nand U2990 (N_2990,N_2616,N_2413);
nor U2991 (N_2991,N_2487,N_2630);
or U2992 (N_2992,N_2651,N_2673);
or U2993 (N_2993,N_2509,N_2484);
and U2994 (N_2994,N_2551,N_2419);
nor U2995 (N_2995,N_2559,N_2677);
and U2996 (N_2996,N_2683,N_2474);
xnor U2997 (N_2997,N_2614,N_2501);
or U2998 (N_2998,N_2508,N_2647);
and U2999 (N_2999,N_2460,N_2598);
nand U3000 (N_3000,N_2812,N_2874);
nand U3001 (N_3001,N_2797,N_2966);
and U3002 (N_3002,N_2886,N_2959);
and U3003 (N_3003,N_2781,N_2744);
xor U3004 (N_3004,N_2904,N_2936);
or U3005 (N_3005,N_2964,N_2819);
and U3006 (N_3006,N_2960,N_2701);
nor U3007 (N_3007,N_2953,N_2779);
nand U3008 (N_3008,N_2765,N_2832);
nor U3009 (N_3009,N_2728,N_2963);
xor U3010 (N_3010,N_2946,N_2705);
or U3011 (N_3011,N_2947,N_2853);
and U3012 (N_3012,N_2907,N_2862);
and U3013 (N_3013,N_2861,N_2961);
xor U3014 (N_3014,N_2807,N_2790);
and U3015 (N_3015,N_2784,N_2796);
or U3016 (N_3016,N_2711,N_2774);
nor U3017 (N_3017,N_2773,N_2938);
nor U3018 (N_3018,N_2937,N_2893);
or U3019 (N_3019,N_2943,N_2822);
and U3020 (N_3020,N_2756,N_2917);
nand U3021 (N_3021,N_2992,N_2923);
xor U3022 (N_3022,N_2787,N_2981);
and U3023 (N_3023,N_2973,N_2748);
or U3024 (N_3024,N_2767,N_2898);
or U3025 (N_3025,N_2914,N_2899);
xor U3026 (N_3026,N_2778,N_2795);
xnor U3027 (N_3027,N_2785,N_2809);
nor U3028 (N_3028,N_2997,N_2873);
nand U3029 (N_3029,N_2841,N_2743);
or U3030 (N_3030,N_2894,N_2855);
xnor U3031 (N_3031,N_2846,N_2872);
and U3032 (N_3032,N_2972,N_2916);
xnor U3033 (N_3033,N_2901,N_2933);
nor U3034 (N_3034,N_2956,N_2840);
nand U3035 (N_3035,N_2977,N_2830);
or U3036 (N_3036,N_2948,N_2805);
or U3037 (N_3037,N_2967,N_2726);
or U3038 (N_3038,N_2780,N_2965);
nand U3039 (N_3039,N_2794,N_2739);
xnor U3040 (N_3040,N_2706,N_2771);
nor U3041 (N_3041,N_2906,N_2751);
nand U3042 (N_3042,N_2957,N_2721);
or U3043 (N_3043,N_2772,N_2883);
and U3044 (N_3044,N_2952,N_2745);
nor U3045 (N_3045,N_2789,N_2718);
and U3046 (N_3046,N_2725,N_2754);
and U3047 (N_3047,N_2791,N_2708);
and U3048 (N_3048,N_2940,N_2740);
and U3049 (N_3049,N_2820,N_2742);
xnor U3050 (N_3050,N_2881,N_2985);
nor U3051 (N_3051,N_2835,N_2715);
nand U3052 (N_3052,N_2995,N_2803);
or U3053 (N_3053,N_2837,N_2860);
nor U3054 (N_3054,N_2935,N_2849);
xnor U3055 (N_3055,N_2833,N_2878);
xnor U3056 (N_3056,N_2991,N_2926);
and U3057 (N_3057,N_2769,N_2804);
nand U3058 (N_3058,N_2723,N_2736);
or U3059 (N_3059,N_2815,N_2752);
xor U3060 (N_3060,N_2802,N_2863);
xnor U3061 (N_3061,N_2851,N_2984);
xnor U3062 (N_3062,N_2854,N_2996);
xnor U3063 (N_3063,N_2871,N_2889);
nand U3064 (N_3064,N_2817,N_2707);
nand U3065 (N_3065,N_2896,N_2989);
nor U3066 (N_3066,N_2912,N_2888);
nand U3067 (N_3067,N_2870,N_2798);
or U3068 (N_3068,N_2836,N_2763);
or U3069 (N_3069,N_2910,N_2920);
nor U3070 (N_3070,N_2848,N_2824);
nand U3071 (N_3071,N_2806,N_2844);
nor U3072 (N_3072,N_2955,N_2958);
and U3073 (N_3073,N_2845,N_2843);
or U3074 (N_3074,N_2999,N_2944);
nand U3075 (N_3075,N_2924,N_2993);
and U3076 (N_3076,N_2818,N_2929);
nor U3077 (N_3077,N_2903,N_2786);
nor U3078 (N_3078,N_2799,N_2770);
and U3079 (N_3079,N_2868,N_2750);
or U3080 (N_3080,N_2969,N_2749);
xor U3081 (N_3081,N_2814,N_2852);
nand U3082 (N_3082,N_2962,N_2988);
nand U3083 (N_3083,N_2867,N_2792);
and U3084 (N_3084,N_2941,N_2950);
xnor U3085 (N_3085,N_2908,N_2776);
xor U3086 (N_3086,N_2753,N_2828);
or U3087 (N_3087,N_2983,N_2880);
nor U3088 (N_3088,N_2831,N_2813);
and U3089 (N_3089,N_2755,N_2827);
xor U3090 (N_3090,N_2713,N_2700);
or U3091 (N_3091,N_2925,N_2759);
nand U3092 (N_3092,N_2857,N_2890);
or U3093 (N_3093,N_2746,N_2879);
nor U3094 (N_3094,N_2724,N_2709);
nand U3095 (N_3095,N_2712,N_2704);
and U3096 (N_3096,N_2865,N_2826);
or U3097 (N_3097,N_2987,N_2877);
and U3098 (N_3098,N_2856,N_2887);
or U3099 (N_3099,N_2823,N_2945);
nor U3100 (N_3100,N_2764,N_2980);
xnor U3101 (N_3101,N_2869,N_2892);
xnor U3102 (N_3102,N_2825,N_2735);
xor U3103 (N_3103,N_2930,N_2951);
nor U3104 (N_3104,N_2733,N_2994);
and U3105 (N_3105,N_2884,N_2968);
xor U3106 (N_3106,N_2876,N_2975);
nor U3107 (N_3107,N_2954,N_2839);
xor U3108 (N_3108,N_2921,N_2990);
or U3109 (N_3109,N_2782,N_2838);
or U3110 (N_3110,N_2928,N_2834);
nand U3111 (N_3111,N_2913,N_2768);
nand U3112 (N_3112,N_2777,N_2801);
and U3113 (N_3113,N_2891,N_2760);
and U3114 (N_3114,N_2788,N_2942);
and U3115 (N_3115,N_2998,N_2730);
xor U3116 (N_3116,N_2727,N_2741);
or U3117 (N_3117,N_2927,N_2738);
and U3118 (N_3118,N_2895,N_2931);
and U3119 (N_3119,N_2847,N_2978);
and U3120 (N_3120,N_2934,N_2900);
or U3121 (N_3121,N_2783,N_2710);
nor U3122 (N_3122,N_2714,N_2829);
nor U3123 (N_3123,N_2702,N_2808);
xor U3124 (N_3124,N_2897,N_2758);
nand U3125 (N_3125,N_2717,N_2949);
and U3126 (N_3126,N_2982,N_2939);
nand U3127 (N_3127,N_2800,N_2766);
nand U3128 (N_3128,N_2793,N_2859);
nor U3129 (N_3129,N_2703,N_2732);
or U3130 (N_3130,N_2979,N_2731);
xnor U3131 (N_3131,N_2885,N_2762);
nor U3132 (N_3132,N_2974,N_2722);
and U3133 (N_3133,N_2919,N_2729);
xnor U3134 (N_3134,N_2775,N_2882);
xor U3135 (N_3135,N_2905,N_2918);
nor U3136 (N_3136,N_2911,N_2976);
nand U3137 (N_3137,N_2821,N_2761);
and U3138 (N_3138,N_2971,N_2719);
nand U3139 (N_3139,N_2737,N_2986);
nor U3140 (N_3140,N_2915,N_2734);
nand U3141 (N_3141,N_2720,N_2970);
or U3142 (N_3142,N_2902,N_2850);
and U3143 (N_3143,N_2716,N_2810);
and U3144 (N_3144,N_2747,N_2922);
nand U3145 (N_3145,N_2811,N_2757);
or U3146 (N_3146,N_2866,N_2875);
nand U3147 (N_3147,N_2932,N_2842);
xnor U3148 (N_3148,N_2816,N_2858);
and U3149 (N_3149,N_2909,N_2864);
nand U3150 (N_3150,N_2737,N_2803);
xnor U3151 (N_3151,N_2733,N_2883);
and U3152 (N_3152,N_2729,N_2779);
nand U3153 (N_3153,N_2872,N_2819);
and U3154 (N_3154,N_2956,N_2702);
or U3155 (N_3155,N_2763,N_2761);
or U3156 (N_3156,N_2784,N_2834);
or U3157 (N_3157,N_2911,N_2870);
xor U3158 (N_3158,N_2703,N_2876);
nand U3159 (N_3159,N_2756,N_2886);
nor U3160 (N_3160,N_2887,N_2749);
xnor U3161 (N_3161,N_2964,N_2742);
nor U3162 (N_3162,N_2764,N_2805);
nor U3163 (N_3163,N_2768,N_2874);
nand U3164 (N_3164,N_2756,N_2904);
or U3165 (N_3165,N_2780,N_2840);
or U3166 (N_3166,N_2768,N_2867);
and U3167 (N_3167,N_2891,N_2701);
and U3168 (N_3168,N_2973,N_2700);
xor U3169 (N_3169,N_2776,N_2767);
or U3170 (N_3170,N_2848,N_2838);
nand U3171 (N_3171,N_2971,N_2707);
or U3172 (N_3172,N_2948,N_2836);
or U3173 (N_3173,N_2901,N_2790);
nor U3174 (N_3174,N_2914,N_2741);
or U3175 (N_3175,N_2738,N_2705);
xor U3176 (N_3176,N_2918,N_2943);
nor U3177 (N_3177,N_2891,N_2783);
nand U3178 (N_3178,N_2802,N_2974);
nor U3179 (N_3179,N_2702,N_2700);
or U3180 (N_3180,N_2876,N_2937);
nor U3181 (N_3181,N_2763,N_2870);
xor U3182 (N_3182,N_2967,N_2881);
nand U3183 (N_3183,N_2916,N_2925);
xor U3184 (N_3184,N_2874,N_2927);
nand U3185 (N_3185,N_2940,N_2853);
nand U3186 (N_3186,N_2910,N_2752);
and U3187 (N_3187,N_2950,N_2885);
and U3188 (N_3188,N_2734,N_2821);
nor U3189 (N_3189,N_2925,N_2860);
nor U3190 (N_3190,N_2909,N_2878);
nor U3191 (N_3191,N_2945,N_2822);
nor U3192 (N_3192,N_2812,N_2958);
xor U3193 (N_3193,N_2958,N_2940);
xor U3194 (N_3194,N_2845,N_2965);
or U3195 (N_3195,N_2818,N_2914);
and U3196 (N_3196,N_2843,N_2993);
or U3197 (N_3197,N_2863,N_2706);
or U3198 (N_3198,N_2909,N_2720);
nand U3199 (N_3199,N_2781,N_2955);
or U3200 (N_3200,N_2866,N_2773);
nor U3201 (N_3201,N_2899,N_2719);
or U3202 (N_3202,N_2715,N_2815);
xor U3203 (N_3203,N_2745,N_2839);
and U3204 (N_3204,N_2834,N_2882);
nand U3205 (N_3205,N_2982,N_2921);
nor U3206 (N_3206,N_2999,N_2714);
xnor U3207 (N_3207,N_2760,N_2955);
nor U3208 (N_3208,N_2917,N_2848);
and U3209 (N_3209,N_2870,N_2835);
nand U3210 (N_3210,N_2791,N_2767);
xnor U3211 (N_3211,N_2924,N_2843);
or U3212 (N_3212,N_2802,N_2953);
and U3213 (N_3213,N_2704,N_2744);
xor U3214 (N_3214,N_2766,N_2820);
or U3215 (N_3215,N_2911,N_2927);
or U3216 (N_3216,N_2783,N_2933);
xnor U3217 (N_3217,N_2934,N_2983);
nor U3218 (N_3218,N_2875,N_2766);
nand U3219 (N_3219,N_2780,N_2984);
nand U3220 (N_3220,N_2842,N_2839);
xor U3221 (N_3221,N_2775,N_2754);
and U3222 (N_3222,N_2996,N_2870);
nand U3223 (N_3223,N_2983,N_2855);
xnor U3224 (N_3224,N_2774,N_2960);
nor U3225 (N_3225,N_2995,N_2814);
xnor U3226 (N_3226,N_2788,N_2836);
and U3227 (N_3227,N_2815,N_2978);
nand U3228 (N_3228,N_2847,N_2889);
nand U3229 (N_3229,N_2712,N_2859);
and U3230 (N_3230,N_2764,N_2804);
and U3231 (N_3231,N_2704,N_2988);
and U3232 (N_3232,N_2839,N_2730);
nor U3233 (N_3233,N_2785,N_2884);
and U3234 (N_3234,N_2786,N_2825);
xor U3235 (N_3235,N_2890,N_2782);
or U3236 (N_3236,N_2988,N_2782);
nand U3237 (N_3237,N_2754,N_2880);
or U3238 (N_3238,N_2988,N_2742);
nand U3239 (N_3239,N_2849,N_2974);
and U3240 (N_3240,N_2776,N_2954);
and U3241 (N_3241,N_2813,N_2844);
or U3242 (N_3242,N_2961,N_2829);
nand U3243 (N_3243,N_2827,N_2732);
nor U3244 (N_3244,N_2723,N_2970);
nand U3245 (N_3245,N_2988,N_2824);
nor U3246 (N_3246,N_2772,N_2908);
nand U3247 (N_3247,N_2884,N_2883);
xor U3248 (N_3248,N_2899,N_2802);
or U3249 (N_3249,N_2757,N_2718);
and U3250 (N_3250,N_2915,N_2727);
nor U3251 (N_3251,N_2972,N_2870);
or U3252 (N_3252,N_2711,N_2839);
and U3253 (N_3253,N_2728,N_2928);
nand U3254 (N_3254,N_2722,N_2746);
and U3255 (N_3255,N_2973,N_2908);
xor U3256 (N_3256,N_2742,N_2831);
or U3257 (N_3257,N_2767,N_2820);
or U3258 (N_3258,N_2762,N_2767);
nand U3259 (N_3259,N_2994,N_2845);
xor U3260 (N_3260,N_2742,N_2775);
nor U3261 (N_3261,N_2855,N_2734);
nand U3262 (N_3262,N_2760,N_2997);
and U3263 (N_3263,N_2997,N_2894);
xor U3264 (N_3264,N_2915,N_2818);
or U3265 (N_3265,N_2791,N_2934);
nor U3266 (N_3266,N_2871,N_2945);
or U3267 (N_3267,N_2997,N_2824);
nand U3268 (N_3268,N_2731,N_2773);
nor U3269 (N_3269,N_2936,N_2919);
xor U3270 (N_3270,N_2845,N_2998);
nand U3271 (N_3271,N_2782,N_2943);
or U3272 (N_3272,N_2822,N_2820);
nor U3273 (N_3273,N_2710,N_2997);
and U3274 (N_3274,N_2909,N_2780);
and U3275 (N_3275,N_2817,N_2908);
and U3276 (N_3276,N_2881,N_2808);
nand U3277 (N_3277,N_2882,N_2906);
nand U3278 (N_3278,N_2892,N_2724);
xnor U3279 (N_3279,N_2768,N_2901);
or U3280 (N_3280,N_2920,N_2970);
and U3281 (N_3281,N_2886,N_2924);
xor U3282 (N_3282,N_2854,N_2770);
and U3283 (N_3283,N_2814,N_2973);
xnor U3284 (N_3284,N_2953,N_2773);
or U3285 (N_3285,N_2820,N_2970);
and U3286 (N_3286,N_2848,N_2712);
and U3287 (N_3287,N_2773,N_2811);
or U3288 (N_3288,N_2988,N_2790);
xnor U3289 (N_3289,N_2905,N_2746);
and U3290 (N_3290,N_2841,N_2868);
xnor U3291 (N_3291,N_2770,N_2805);
nand U3292 (N_3292,N_2756,N_2833);
nor U3293 (N_3293,N_2700,N_2826);
xnor U3294 (N_3294,N_2870,N_2705);
xor U3295 (N_3295,N_2798,N_2790);
xnor U3296 (N_3296,N_2728,N_2770);
or U3297 (N_3297,N_2716,N_2887);
nand U3298 (N_3298,N_2777,N_2804);
nor U3299 (N_3299,N_2818,N_2937);
and U3300 (N_3300,N_3208,N_3185);
and U3301 (N_3301,N_3226,N_3148);
xnor U3302 (N_3302,N_3143,N_3243);
nand U3303 (N_3303,N_3200,N_3202);
or U3304 (N_3304,N_3132,N_3090);
and U3305 (N_3305,N_3121,N_3071);
xor U3306 (N_3306,N_3274,N_3150);
and U3307 (N_3307,N_3223,N_3125);
nand U3308 (N_3308,N_3113,N_3245);
nand U3309 (N_3309,N_3041,N_3066);
or U3310 (N_3310,N_3250,N_3221);
and U3311 (N_3311,N_3294,N_3012);
nand U3312 (N_3312,N_3198,N_3218);
nand U3313 (N_3313,N_3038,N_3118);
or U3314 (N_3314,N_3084,N_3297);
xnor U3315 (N_3315,N_3036,N_3133);
xor U3316 (N_3316,N_3107,N_3230);
nor U3317 (N_3317,N_3251,N_3023);
xor U3318 (N_3318,N_3264,N_3186);
or U3319 (N_3319,N_3089,N_3163);
or U3320 (N_3320,N_3234,N_3281);
and U3321 (N_3321,N_3085,N_3063);
or U3322 (N_3322,N_3286,N_3181);
nor U3323 (N_3323,N_3296,N_3224);
and U3324 (N_3324,N_3276,N_3057);
or U3325 (N_3325,N_3255,N_3015);
and U3326 (N_3326,N_3101,N_3029);
and U3327 (N_3327,N_3231,N_3169);
xnor U3328 (N_3328,N_3190,N_3266);
nand U3329 (N_3329,N_3065,N_3261);
and U3330 (N_3330,N_3222,N_3152);
nor U3331 (N_3331,N_3244,N_3058);
xnor U3332 (N_3332,N_3116,N_3111);
xnor U3333 (N_3333,N_3177,N_3040);
and U3334 (N_3334,N_3178,N_3265);
and U3335 (N_3335,N_3135,N_3045);
xor U3336 (N_3336,N_3158,N_3099);
nor U3337 (N_3337,N_3124,N_3034);
or U3338 (N_3338,N_3102,N_3184);
or U3339 (N_3339,N_3284,N_3044);
xnor U3340 (N_3340,N_3174,N_3262);
xnor U3341 (N_3341,N_3130,N_3056);
and U3342 (N_3342,N_3217,N_3160);
and U3343 (N_3343,N_3214,N_3215);
or U3344 (N_3344,N_3013,N_3128);
xor U3345 (N_3345,N_3093,N_3175);
and U3346 (N_3346,N_3127,N_3249);
and U3347 (N_3347,N_3061,N_3104);
or U3348 (N_3348,N_3191,N_3188);
nand U3349 (N_3349,N_3120,N_3080);
or U3350 (N_3350,N_3164,N_3009);
nand U3351 (N_3351,N_3087,N_3292);
nand U3352 (N_3352,N_3033,N_3103);
nand U3353 (N_3353,N_3176,N_3254);
or U3354 (N_3354,N_3242,N_3142);
and U3355 (N_3355,N_3094,N_3026);
nor U3356 (N_3356,N_3278,N_3024);
xnor U3357 (N_3357,N_3021,N_3110);
nor U3358 (N_3358,N_3020,N_3138);
xnor U3359 (N_3359,N_3232,N_3059);
or U3360 (N_3360,N_3027,N_3165);
xor U3361 (N_3361,N_3241,N_3210);
xnor U3362 (N_3362,N_3277,N_3194);
and U3363 (N_3363,N_3035,N_3134);
or U3364 (N_3364,N_3289,N_3207);
nor U3365 (N_3365,N_3117,N_3016);
and U3366 (N_3366,N_3098,N_3285);
xor U3367 (N_3367,N_3287,N_3227);
xnor U3368 (N_3368,N_3060,N_3204);
nand U3369 (N_3369,N_3256,N_3258);
nand U3370 (N_3370,N_3180,N_3288);
and U3371 (N_3371,N_3161,N_3273);
or U3372 (N_3372,N_3039,N_3031);
nor U3373 (N_3373,N_3229,N_3129);
nand U3374 (N_3374,N_3228,N_3046);
nand U3375 (N_3375,N_3077,N_3079);
nand U3376 (N_3376,N_3115,N_3239);
nor U3377 (N_3377,N_3270,N_3053);
and U3378 (N_3378,N_3048,N_3083);
nand U3379 (N_3379,N_3139,N_3106);
nor U3380 (N_3380,N_3193,N_3192);
and U3381 (N_3381,N_3213,N_3182);
nor U3382 (N_3382,N_3076,N_3268);
nor U3383 (N_3383,N_3141,N_3216);
nand U3384 (N_3384,N_3206,N_3153);
nor U3385 (N_3385,N_3167,N_3097);
nor U3386 (N_3386,N_3203,N_3237);
nand U3387 (N_3387,N_3002,N_3290);
nor U3388 (N_3388,N_3131,N_3280);
and U3389 (N_3389,N_3299,N_3267);
nor U3390 (N_3390,N_3095,N_3197);
nor U3391 (N_3391,N_3248,N_3259);
or U3392 (N_3392,N_3147,N_3017);
nor U3393 (N_3393,N_3233,N_3108);
and U3394 (N_3394,N_3081,N_3269);
or U3395 (N_3395,N_3211,N_3070);
xnor U3396 (N_3396,N_3008,N_3088);
xor U3397 (N_3397,N_3173,N_3253);
and U3398 (N_3398,N_3205,N_3189);
or U3399 (N_3399,N_3183,N_3054);
and U3400 (N_3400,N_3092,N_3220);
and U3401 (N_3401,N_3072,N_3159);
nand U3402 (N_3402,N_3005,N_3082);
nand U3403 (N_3403,N_3022,N_3049);
and U3404 (N_3404,N_3279,N_3050);
nor U3405 (N_3405,N_3140,N_3225);
nand U3406 (N_3406,N_3298,N_3187);
and U3407 (N_3407,N_3042,N_3260);
and U3408 (N_3408,N_3019,N_3114);
nand U3409 (N_3409,N_3007,N_3137);
nor U3410 (N_3410,N_3257,N_3100);
nor U3411 (N_3411,N_3105,N_3052);
xnor U3412 (N_3412,N_3155,N_3064);
and U3413 (N_3413,N_3025,N_3004);
and U3414 (N_3414,N_3014,N_3271);
and U3415 (N_3415,N_3078,N_3272);
nand U3416 (N_3416,N_3145,N_3295);
or U3417 (N_3417,N_3162,N_3263);
nor U3418 (N_3418,N_3126,N_3144);
and U3419 (N_3419,N_3073,N_3096);
nand U3420 (N_3420,N_3119,N_3157);
and U3421 (N_3421,N_3195,N_3011);
and U3422 (N_3422,N_3006,N_3001);
and U3423 (N_3423,N_3172,N_3283);
xnor U3424 (N_3424,N_3109,N_3043);
and U3425 (N_3425,N_3209,N_3170);
nor U3426 (N_3426,N_3136,N_3146);
and U3427 (N_3427,N_3247,N_3235);
or U3428 (N_3428,N_3246,N_3168);
and U3429 (N_3429,N_3151,N_3091);
xor U3430 (N_3430,N_3201,N_3069);
nand U3431 (N_3431,N_3028,N_3112);
nand U3432 (N_3432,N_3018,N_3219);
xnor U3433 (N_3433,N_3075,N_3055);
xor U3434 (N_3434,N_3010,N_3051);
or U3435 (N_3435,N_3238,N_3030);
or U3436 (N_3436,N_3282,N_3123);
and U3437 (N_3437,N_3212,N_3196);
nand U3438 (N_3438,N_3149,N_3240);
and U3439 (N_3439,N_3291,N_3086);
nor U3440 (N_3440,N_3074,N_3236);
and U3441 (N_3441,N_3067,N_3003);
or U3442 (N_3442,N_3171,N_3122);
nand U3443 (N_3443,N_3047,N_3275);
or U3444 (N_3444,N_3166,N_3199);
or U3445 (N_3445,N_3068,N_3179);
nor U3446 (N_3446,N_3037,N_3252);
and U3447 (N_3447,N_3062,N_3000);
nor U3448 (N_3448,N_3293,N_3156);
nor U3449 (N_3449,N_3032,N_3154);
or U3450 (N_3450,N_3025,N_3200);
nor U3451 (N_3451,N_3211,N_3256);
and U3452 (N_3452,N_3278,N_3022);
and U3453 (N_3453,N_3058,N_3205);
or U3454 (N_3454,N_3289,N_3134);
nand U3455 (N_3455,N_3271,N_3072);
nand U3456 (N_3456,N_3051,N_3044);
and U3457 (N_3457,N_3138,N_3283);
nand U3458 (N_3458,N_3057,N_3079);
or U3459 (N_3459,N_3079,N_3183);
nor U3460 (N_3460,N_3047,N_3010);
xor U3461 (N_3461,N_3220,N_3224);
nand U3462 (N_3462,N_3237,N_3170);
nor U3463 (N_3463,N_3111,N_3016);
nor U3464 (N_3464,N_3170,N_3250);
or U3465 (N_3465,N_3006,N_3105);
nor U3466 (N_3466,N_3137,N_3011);
nor U3467 (N_3467,N_3271,N_3209);
and U3468 (N_3468,N_3152,N_3129);
xor U3469 (N_3469,N_3267,N_3014);
xnor U3470 (N_3470,N_3156,N_3017);
nor U3471 (N_3471,N_3028,N_3182);
and U3472 (N_3472,N_3060,N_3001);
or U3473 (N_3473,N_3160,N_3053);
nor U3474 (N_3474,N_3094,N_3204);
or U3475 (N_3475,N_3047,N_3169);
or U3476 (N_3476,N_3267,N_3132);
and U3477 (N_3477,N_3009,N_3181);
and U3478 (N_3478,N_3224,N_3134);
nor U3479 (N_3479,N_3026,N_3056);
xor U3480 (N_3480,N_3167,N_3207);
xnor U3481 (N_3481,N_3128,N_3277);
nor U3482 (N_3482,N_3211,N_3167);
or U3483 (N_3483,N_3016,N_3193);
or U3484 (N_3484,N_3094,N_3287);
xnor U3485 (N_3485,N_3043,N_3133);
and U3486 (N_3486,N_3174,N_3037);
xnor U3487 (N_3487,N_3220,N_3080);
or U3488 (N_3488,N_3272,N_3240);
xor U3489 (N_3489,N_3247,N_3104);
xnor U3490 (N_3490,N_3248,N_3169);
xor U3491 (N_3491,N_3256,N_3177);
nand U3492 (N_3492,N_3193,N_3165);
nand U3493 (N_3493,N_3010,N_3054);
xor U3494 (N_3494,N_3064,N_3215);
xnor U3495 (N_3495,N_3074,N_3094);
nand U3496 (N_3496,N_3083,N_3227);
or U3497 (N_3497,N_3242,N_3179);
nor U3498 (N_3498,N_3014,N_3118);
and U3499 (N_3499,N_3145,N_3161);
nor U3500 (N_3500,N_3208,N_3272);
nand U3501 (N_3501,N_3226,N_3113);
or U3502 (N_3502,N_3232,N_3189);
nand U3503 (N_3503,N_3041,N_3091);
or U3504 (N_3504,N_3180,N_3104);
nor U3505 (N_3505,N_3199,N_3215);
or U3506 (N_3506,N_3049,N_3269);
or U3507 (N_3507,N_3112,N_3173);
or U3508 (N_3508,N_3013,N_3026);
and U3509 (N_3509,N_3212,N_3114);
xor U3510 (N_3510,N_3171,N_3039);
or U3511 (N_3511,N_3178,N_3269);
nand U3512 (N_3512,N_3250,N_3003);
and U3513 (N_3513,N_3138,N_3239);
or U3514 (N_3514,N_3284,N_3140);
and U3515 (N_3515,N_3213,N_3198);
nand U3516 (N_3516,N_3118,N_3255);
and U3517 (N_3517,N_3177,N_3145);
xor U3518 (N_3518,N_3227,N_3030);
and U3519 (N_3519,N_3077,N_3106);
and U3520 (N_3520,N_3062,N_3194);
or U3521 (N_3521,N_3147,N_3096);
nor U3522 (N_3522,N_3191,N_3127);
and U3523 (N_3523,N_3139,N_3148);
or U3524 (N_3524,N_3243,N_3201);
nand U3525 (N_3525,N_3273,N_3255);
xor U3526 (N_3526,N_3125,N_3217);
or U3527 (N_3527,N_3275,N_3117);
xnor U3528 (N_3528,N_3140,N_3061);
or U3529 (N_3529,N_3051,N_3212);
or U3530 (N_3530,N_3249,N_3174);
or U3531 (N_3531,N_3145,N_3252);
nor U3532 (N_3532,N_3092,N_3031);
or U3533 (N_3533,N_3089,N_3287);
nor U3534 (N_3534,N_3283,N_3043);
or U3535 (N_3535,N_3203,N_3170);
nand U3536 (N_3536,N_3256,N_3262);
nor U3537 (N_3537,N_3138,N_3145);
nor U3538 (N_3538,N_3215,N_3223);
nor U3539 (N_3539,N_3143,N_3234);
or U3540 (N_3540,N_3130,N_3109);
nand U3541 (N_3541,N_3129,N_3296);
and U3542 (N_3542,N_3068,N_3286);
and U3543 (N_3543,N_3025,N_3287);
xnor U3544 (N_3544,N_3128,N_3056);
or U3545 (N_3545,N_3131,N_3214);
xor U3546 (N_3546,N_3027,N_3083);
and U3547 (N_3547,N_3294,N_3205);
nor U3548 (N_3548,N_3081,N_3031);
and U3549 (N_3549,N_3168,N_3118);
nand U3550 (N_3550,N_3221,N_3024);
and U3551 (N_3551,N_3150,N_3207);
nor U3552 (N_3552,N_3213,N_3189);
xnor U3553 (N_3553,N_3113,N_3053);
nor U3554 (N_3554,N_3121,N_3059);
nor U3555 (N_3555,N_3159,N_3004);
nand U3556 (N_3556,N_3285,N_3293);
and U3557 (N_3557,N_3264,N_3206);
nor U3558 (N_3558,N_3117,N_3183);
or U3559 (N_3559,N_3299,N_3113);
nand U3560 (N_3560,N_3240,N_3214);
nor U3561 (N_3561,N_3181,N_3267);
and U3562 (N_3562,N_3009,N_3255);
nand U3563 (N_3563,N_3103,N_3061);
xnor U3564 (N_3564,N_3071,N_3000);
nand U3565 (N_3565,N_3271,N_3166);
nor U3566 (N_3566,N_3131,N_3162);
nor U3567 (N_3567,N_3099,N_3055);
or U3568 (N_3568,N_3013,N_3295);
nand U3569 (N_3569,N_3269,N_3036);
nor U3570 (N_3570,N_3280,N_3050);
nor U3571 (N_3571,N_3065,N_3007);
and U3572 (N_3572,N_3049,N_3078);
and U3573 (N_3573,N_3268,N_3112);
nor U3574 (N_3574,N_3267,N_3095);
nor U3575 (N_3575,N_3284,N_3016);
nand U3576 (N_3576,N_3139,N_3058);
xnor U3577 (N_3577,N_3213,N_3017);
nand U3578 (N_3578,N_3240,N_3153);
nand U3579 (N_3579,N_3018,N_3033);
or U3580 (N_3580,N_3140,N_3286);
or U3581 (N_3581,N_3292,N_3164);
or U3582 (N_3582,N_3219,N_3116);
xor U3583 (N_3583,N_3095,N_3223);
nor U3584 (N_3584,N_3196,N_3065);
nor U3585 (N_3585,N_3072,N_3077);
or U3586 (N_3586,N_3107,N_3002);
nor U3587 (N_3587,N_3190,N_3008);
nand U3588 (N_3588,N_3122,N_3189);
nand U3589 (N_3589,N_3169,N_3083);
xor U3590 (N_3590,N_3060,N_3202);
nand U3591 (N_3591,N_3221,N_3283);
nand U3592 (N_3592,N_3102,N_3172);
and U3593 (N_3593,N_3033,N_3042);
and U3594 (N_3594,N_3240,N_3223);
xnor U3595 (N_3595,N_3036,N_3200);
nand U3596 (N_3596,N_3174,N_3213);
or U3597 (N_3597,N_3084,N_3106);
xor U3598 (N_3598,N_3232,N_3176);
and U3599 (N_3599,N_3047,N_3182);
nand U3600 (N_3600,N_3497,N_3456);
nand U3601 (N_3601,N_3589,N_3541);
or U3602 (N_3602,N_3590,N_3583);
xor U3603 (N_3603,N_3436,N_3434);
nor U3604 (N_3604,N_3438,N_3479);
xor U3605 (N_3605,N_3525,N_3408);
xnor U3606 (N_3606,N_3341,N_3562);
xnor U3607 (N_3607,N_3578,N_3377);
or U3608 (N_3608,N_3474,N_3320);
or U3609 (N_3609,N_3343,N_3493);
nor U3610 (N_3610,N_3547,N_3482);
nor U3611 (N_3611,N_3512,N_3430);
or U3612 (N_3612,N_3523,N_3432);
xnor U3613 (N_3613,N_3490,N_3545);
and U3614 (N_3614,N_3591,N_3526);
nor U3615 (N_3615,N_3557,N_3404);
nand U3616 (N_3616,N_3559,N_3387);
or U3617 (N_3617,N_3385,N_3326);
nand U3618 (N_3618,N_3515,N_3459);
nand U3619 (N_3619,N_3542,N_3593);
xor U3620 (N_3620,N_3575,N_3533);
and U3621 (N_3621,N_3386,N_3349);
or U3622 (N_3622,N_3450,N_3330);
nor U3623 (N_3623,N_3571,N_3465);
nand U3624 (N_3624,N_3508,N_3527);
and U3625 (N_3625,N_3599,N_3317);
xnor U3626 (N_3626,N_3572,N_3372);
xnor U3627 (N_3627,N_3417,N_3472);
or U3628 (N_3628,N_3480,N_3457);
nor U3629 (N_3629,N_3448,N_3581);
xor U3630 (N_3630,N_3391,N_3580);
and U3631 (N_3631,N_3498,N_3302);
and U3632 (N_3632,N_3312,N_3440);
nor U3633 (N_3633,N_3588,N_3462);
or U3634 (N_3634,N_3379,N_3367);
xnor U3635 (N_3635,N_3524,N_3470);
xor U3636 (N_3636,N_3332,N_3419);
and U3637 (N_3637,N_3411,N_3370);
nor U3638 (N_3638,N_3458,N_3516);
or U3639 (N_3639,N_3431,N_3475);
or U3640 (N_3640,N_3418,N_3460);
nor U3641 (N_3641,N_3494,N_3528);
xor U3642 (N_3642,N_3439,N_3551);
xnor U3643 (N_3643,N_3483,N_3501);
nor U3644 (N_3644,N_3521,N_3577);
nand U3645 (N_3645,N_3441,N_3337);
and U3646 (N_3646,N_3374,N_3336);
and U3647 (N_3647,N_3429,N_3595);
or U3648 (N_3648,N_3442,N_3363);
nor U3649 (N_3649,N_3415,N_3504);
xor U3650 (N_3650,N_3354,N_3485);
or U3651 (N_3651,N_3300,N_3371);
and U3652 (N_3652,N_3325,N_3424);
nor U3653 (N_3653,N_3453,N_3513);
and U3654 (N_3654,N_3544,N_3303);
or U3655 (N_3655,N_3333,N_3394);
nand U3656 (N_3656,N_3369,N_3576);
xnor U3657 (N_3657,N_3530,N_3564);
nor U3658 (N_3658,N_3356,N_3335);
nor U3659 (N_3659,N_3534,N_3445);
nor U3660 (N_3660,N_3409,N_3405);
nand U3661 (N_3661,N_3433,N_3536);
and U3662 (N_3662,N_3381,N_3520);
xnor U3663 (N_3663,N_3507,N_3584);
and U3664 (N_3664,N_3410,N_3362);
nand U3665 (N_3665,N_3423,N_3582);
nor U3666 (N_3666,N_3505,N_3447);
xor U3667 (N_3667,N_3412,N_3509);
nand U3668 (N_3668,N_3471,N_3484);
nand U3669 (N_3669,N_3489,N_3383);
or U3670 (N_3670,N_3449,N_3364);
nor U3671 (N_3671,N_3594,N_3554);
xor U3672 (N_3672,N_3334,N_3368);
and U3673 (N_3673,N_3388,N_3579);
nand U3674 (N_3674,N_3307,N_3322);
nor U3675 (N_3675,N_3398,N_3309);
or U3676 (N_3676,N_3426,N_3568);
nor U3677 (N_3677,N_3455,N_3304);
xor U3678 (N_3678,N_3446,N_3306);
nor U3679 (N_3679,N_3478,N_3382);
and U3680 (N_3680,N_3339,N_3556);
or U3681 (N_3681,N_3351,N_3323);
nand U3682 (N_3682,N_3375,N_3466);
nor U3683 (N_3683,N_3558,N_3443);
or U3684 (N_3684,N_3403,N_3522);
nor U3685 (N_3685,N_3392,N_3360);
nor U3686 (N_3686,N_3384,N_3315);
xor U3687 (N_3687,N_3451,N_3597);
and U3688 (N_3688,N_3329,N_3587);
xor U3689 (N_3689,N_3517,N_3569);
nand U3690 (N_3690,N_3305,N_3477);
or U3691 (N_3691,N_3406,N_3567);
nand U3692 (N_3692,N_3301,N_3319);
nor U3693 (N_3693,N_3510,N_3346);
nand U3694 (N_3694,N_3464,N_3352);
nand U3695 (N_3695,N_3586,N_3324);
nor U3696 (N_3696,N_3425,N_3347);
and U3697 (N_3697,N_3413,N_3531);
nand U3698 (N_3698,N_3444,N_3563);
nand U3699 (N_3699,N_3555,N_3560);
xnor U3700 (N_3700,N_3401,N_3592);
and U3701 (N_3701,N_3348,N_3313);
and U3702 (N_3702,N_3344,N_3553);
nand U3703 (N_3703,N_3473,N_3511);
nor U3704 (N_3704,N_3596,N_3397);
xor U3705 (N_3705,N_3355,N_3492);
and U3706 (N_3706,N_3486,N_3598);
nand U3707 (N_3707,N_3357,N_3331);
xor U3708 (N_3708,N_3316,N_3548);
or U3709 (N_3709,N_3566,N_3506);
xnor U3710 (N_3710,N_3353,N_3543);
and U3711 (N_3711,N_3499,N_3389);
nand U3712 (N_3712,N_3538,N_3540);
xor U3713 (N_3713,N_3550,N_3414);
nor U3714 (N_3714,N_3565,N_3361);
nor U3715 (N_3715,N_3314,N_3487);
nand U3716 (N_3716,N_3365,N_3561);
nand U3717 (N_3717,N_3310,N_3463);
nor U3718 (N_3718,N_3503,N_3338);
and U3719 (N_3719,N_3476,N_3529);
xor U3720 (N_3720,N_3532,N_3342);
or U3721 (N_3721,N_3539,N_3366);
xnor U3722 (N_3722,N_3340,N_3491);
and U3723 (N_3723,N_3359,N_3574);
xor U3724 (N_3724,N_3488,N_3437);
or U3725 (N_3725,N_3350,N_3400);
nand U3726 (N_3726,N_3519,N_3549);
and U3727 (N_3727,N_3454,N_3469);
nand U3728 (N_3728,N_3496,N_3500);
or U3729 (N_3729,N_3461,N_3327);
xor U3730 (N_3730,N_3546,N_3345);
nor U3731 (N_3731,N_3502,N_3376);
nand U3732 (N_3732,N_3396,N_3570);
or U3733 (N_3733,N_3537,N_3428);
nor U3734 (N_3734,N_3318,N_3380);
or U3735 (N_3735,N_3407,N_3495);
nor U3736 (N_3736,N_3311,N_3308);
nor U3737 (N_3737,N_3467,N_3393);
nor U3738 (N_3738,N_3321,N_3518);
and U3739 (N_3739,N_3427,N_3468);
nand U3740 (N_3740,N_3585,N_3420);
or U3741 (N_3741,N_3399,N_3373);
or U3742 (N_3742,N_3358,N_3395);
nand U3743 (N_3743,N_3552,N_3573);
or U3744 (N_3744,N_3402,N_3514);
or U3745 (N_3745,N_3535,N_3481);
and U3746 (N_3746,N_3416,N_3452);
or U3747 (N_3747,N_3421,N_3328);
or U3748 (N_3748,N_3435,N_3422);
xnor U3749 (N_3749,N_3378,N_3390);
nor U3750 (N_3750,N_3300,N_3333);
nor U3751 (N_3751,N_3315,N_3485);
nand U3752 (N_3752,N_3374,N_3573);
xor U3753 (N_3753,N_3538,N_3478);
and U3754 (N_3754,N_3565,N_3582);
nand U3755 (N_3755,N_3457,N_3581);
or U3756 (N_3756,N_3535,N_3467);
nor U3757 (N_3757,N_3598,N_3592);
and U3758 (N_3758,N_3527,N_3543);
xor U3759 (N_3759,N_3400,N_3459);
and U3760 (N_3760,N_3515,N_3487);
or U3761 (N_3761,N_3366,N_3336);
nor U3762 (N_3762,N_3544,N_3584);
nor U3763 (N_3763,N_3332,N_3390);
nand U3764 (N_3764,N_3465,N_3481);
nor U3765 (N_3765,N_3561,N_3551);
or U3766 (N_3766,N_3321,N_3301);
xnor U3767 (N_3767,N_3423,N_3492);
or U3768 (N_3768,N_3493,N_3488);
or U3769 (N_3769,N_3589,N_3555);
and U3770 (N_3770,N_3303,N_3513);
or U3771 (N_3771,N_3573,N_3445);
nor U3772 (N_3772,N_3373,N_3478);
xnor U3773 (N_3773,N_3427,N_3323);
xnor U3774 (N_3774,N_3474,N_3562);
or U3775 (N_3775,N_3408,N_3481);
or U3776 (N_3776,N_3349,N_3583);
nor U3777 (N_3777,N_3549,N_3562);
nand U3778 (N_3778,N_3561,N_3503);
nand U3779 (N_3779,N_3524,N_3458);
xor U3780 (N_3780,N_3574,N_3430);
or U3781 (N_3781,N_3512,N_3532);
and U3782 (N_3782,N_3557,N_3389);
nor U3783 (N_3783,N_3430,N_3524);
nand U3784 (N_3784,N_3313,N_3351);
nand U3785 (N_3785,N_3523,N_3399);
nand U3786 (N_3786,N_3556,N_3539);
nor U3787 (N_3787,N_3531,N_3512);
xor U3788 (N_3788,N_3340,N_3571);
and U3789 (N_3789,N_3446,N_3402);
nor U3790 (N_3790,N_3386,N_3598);
and U3791 (N_3791,N_3316,N_3569);
nor U3792 (N_3792,N_3514,N_3379);
nand U3793 (N_3793,N_3349,N_3377);
and U3794 (N_3794,N_3459,N_3478);
or U3795 (N_3795,N_3356,N_3451);
and U3796 (N_3796,N_3438,N_3374);
nor U3797 (N_3797,N_3370,N_3320);
xor U3798 (N_3798,N_3536,N_3518);
xnor U3799 (N_3799,N_3523,N_3583);
nor U3800 (N_3800,N_3371,N_3379);
nor U3801 (N_3801,N_3540,N_3347);
and U3802 (N_3802,N_3388,N_3509);
nand U3803 (N_3803,N_3545,N_3355);
xnor U3804 (N_3804,N_3312,N_3365);
and U3805 (N_3805,N_3436,N_3431);
or U3806 (N_3806,N_3435,N_3443);
xor U3807 (N_3807,N_3358,N_3370);
nor U3808 (N_3808,N_3455,N_3540);
or U3809 (N_3809,N_3439,N_3530);
or U3810 (N_3810,N_3546,N_3334);
xor U3811 (N_3811,N_3439,N_3330);
nand U3812 (N_3812,N_3363,N_3538);
nor U3813 (N_3813,N_3489,N_3459);
xor U3814 (N_3814,N_3415,N_3474);
nor U3815 (N_3815,N_3350,N_3515);
nand U3816 (N_3816,N_3401,N_3322);
nand U3817 (N_3817,N_3451,N_3443);
xnor U3818 (N_3818,N_3424,N_3378);
and U3819 (N_3819,N_3373,N_3543);
xor U3820 (N_3820,N_3504,N_3572);
nor U3821 (N_3821,N_3494,N_3462);
and U3822 (N_3822,N_3549,N_3572);
nand U3823 (N_3823,N_3405,N_3388);
and U3824 (N_3824,N_3461,N_3307);
nand U3825 (N_3825,N_3398,N_3566);
nand U3826 (N_3826,N_3584,N_3521);
nor U3827 (N_3827,N_3532,N_3518);
and U3828 (N_3828,N_3342,N_3471);
or U3829 (N_3829,N_3501,N_3596);
or U3830 (N_3830,N_3368,N_3431);
or U3831 (N_3831,N_3577,N_3317);
xnor U3832 (N_3832,N_3339,N_3517);
or U3833 (N_3833,N_3455,N_3452);
and U3834 (N_3834,N_3349,N_3408);
or U3835 (N_3835,N_3584,N_3562);
and U3836 (N_3836,N_3307,N_3405);
or U3837 (N_3837,N_3456,N_3542);
nor U3838 (N_3838,N_3313,N_3481);
nor U3839 (N_3839,N_3304,N_3312);
nor U3840 (N_3840,N_3439,N_3469);
and U3841 (N_3841,N_3300,N_3440);
or U3842 (N_3842,N_3347,N_3586);
nor U3843 (N_3843,N_3510,N_3533);
nor U3844 (N_3844,N_3493,N_3535);
nor U3845 (N_3845,N_3370,N_3398);
and U3846 (N_3846,N_3435,N_3491);
or U3847 (N_3847,N_3365,N_3333);
nor U3848 (N_3848,N_3494,N_3471);
nor U3849 (N_3849,N_3406,N_3311);
or U3850 (N_3850,N_3529,N_3370);
or U3851 (N_3851,N_3520,N_3513);
nor U3852 (N_3852,N_3461,N_3518);
nand U3853 (N_3853,N_3506,N_3324);
or U3854 (N_3854,N_3341,N_3316);
or U3855 (N_3855,N_3514,N_3520);
and U3856 (N_3856,N_3308,N_3424);
and U3857 (N_3857,N_3599,N_3497);
nor U3858 (N_3858,N_3583,N_3509);
and U3859 (N_3859,N_3591,N_3563);
and U3860 (N_3860,N_3506,N_3339);
nor U3861 (N_3861,N_3492,N_3410);
or U3862 (N_3862,N_3468,N_3391);
nand U3863 (N_3863,N_3497,N_3513);
nand U3864 (N_3864,N_3590,N_3493);
nor U3865 (N_3865,N_3516,N_3576);
nor U3866 (N_3866,N_3513,N_3368);
nand U3867 (N_3867,N_3447,N_3511);
xor U3868 (N_3868,N_3485,N_3462);
nand U3869 (N_3869,N_3369,N_3586);
nor U3870 (N_3870,N_3483,N_3387);
nor U3871 (N_3871,N_3402,N_3412);
and U3872 (N_3872,N_3467,N_3434);
or U3873 (N_3873,N_3415,N_3427);
and U3874 (N_3874,N_3507,N_3524);
or U3875 (N_3875,N_3390,N_3507);
nand U3876 (N_3876,N_3489,N_3578);
xnor U3877 (N_3877,N_3572,N_3305);
or U3878 (N_3878,N_3316,N_3432);
nand U3879 (N_3879,N_3317,N_3520);
or U3880 (N_3880,N_3490,N_3466);
nor U3881 (N_3881,N_3558,N_3351);
and U3882 (N_3882,N_3328,N_3571);
xnor U3883 (N_3883,N_3360,N_3368);
or U3884 (N_3884,N_3471,N_3431);
xor U3885 (N_3885,N_3549,N_3470);
and U3886 (N_3886,N_3495,N_3470);
xor U3887 (N_3887,N_3561,N_3497);
nor U3888 (N_3888,N_3492,N_3430);
and U3889 (N_3889,N_3524,N_3555);
nand U3890 (N_3890,N_3380,N_3311);
or U3891 (N_3891,N_3395,N_3565);
nand U3892 (N_3892,N_3513,N_3543);
nor U3893 (N_3893,N_3328,N_3528);
xor U3894 (N_3894,N_3394,N_3583);
xor U3895 (N_3895,N_3537,N_3589);
xnor U3896 (N_3896,N_3447,N_3391);
or U3897 (N_3897,N_3568,N_3480);
nor U3898 (N_3898,N_3543,N_3354);
or U3899 (N_3899,N_3568,N_3436);
xor U3900 (N_3900,N_3861,N_3688);
nand U3901 (N_3901,N_3682,N_3735);
nor U3902 (N_3902,N_3674,N_3847);
nand U3903 (N_3903,N_3809,N_3814);
nor U3904 (N_3904,N_3810,N_3652);
or U3905 (N_3905,N_3668,N_3840);
xnor U3906 (N_3906,N_3705,N_3691);
and U3907 (N_3907,N_3713,N_3830);
xor U3908 (N_3908,N_3633,N_3724);
nand U3909 (N_3909,N_3807,N_3663);
nor U3910 (N_3910,N_3707,N_3669);
or U3911 (N_3911,N_3845,N_3632);
and U3912 (N_3912,N_3804,N_3865);
or U3913 (N_3913,N_3750,N_3858);
and U3914 (N_3914,N_3676,N_3784);
nand U3915 (N_3915,N_3736,N_3684);
or U3916 (N_3916,N_3681,N_3687);
nor U3917 (N_3917,N_3887,N_3811);
and U3918 (N_3918,N_3734,N_3685);
xor U3919 (N_3919,N_3829,N_3741);
and U3920 (N_3920,N_3850,N_3789);
and U3921 (N_3921,N_3667,N_3717);
nand U3922 (N_3922,N_3884,N_3631);
xor U3923 (N_3923,N_3823,N_3785);
nand U3924 (N_3924,N_3826,N_3798);
xor U3925 (N_3925,N_3604,N_3838);
nor U3926 (N_3926,N_3625,N_3739);
and U3927 (N_3927,N_3801,N_3764);
and U3928 (N_3928,N_3844,N_3656);
nor U3929 (N_3929,N_3609,N_3749);
nor U3930 (N_3930,N_3639,N_3660);
and U3931 (N_3931,N_3710,N_3647);
nand U3932 (N_3932,N_3783,N_3760);
xnor U3933 (N_3933,N_3831,N_3712);
or U3934 (N_3934,N_3730,N_3683);
or U3935 (N_3935,N_3820,N_3637);
or U3936 (N_3936,N_3792,N_3602);
nand U3937 (N_3937,N_3606,N_3839);
xnor U3938 (N_3938,N_3800,N_3716);
nand U3939 (N_3939,N_3700,N_3770);
xnor U3940 (N_3940,N_3813,N_3786);
nor U3941 (N_3941,N_3690,N_3790);
or U3942 (N_3942,N_3748,N_3697);
and U3943 (N_3943,N_3703,N_3888);
xor U3944 (N_3944,N_3653,N_3864);
nand U3945 (N_3945,N_3859,N_3781);
and U3946 (N_3946,N_3816,N_3837);
or U3947 (N_3947,N_3610,N_3648);
and U3948 (N_3948,N_3751,N_3832);
nand U3949 (N_3949,N_3628,N_3627);
or U3950 (N_3950,N_3862,N_3729);
nand U3951 (N_3951,N_3871,N_3744);
xnor U3952 (N_3952,N_3853,N_3763);
and U3953 (N_3953,N_3722,N_3646);
xor U3954 (N_3954,N_3673,N_3822);
xnor U3955 (N_3955,N_3689,N_3616);
nand U3956 (N_3956,N_3893,N_3677);
and U3957 (N_3957,N_3880,N_3793);
or U3958 (N_3958,N_3718,N_3733);
and U3959 (N_3959,N_3617,N_3852);
xor U3960 (N_3960,N_3626,N_3745);
or U3961 (N_3961,N_3740,N_3692);
nand U3962 (N_3962,N_3834,N_3777);
and U3963 (N_3963,N_3870,N_3780);
and U3964 (N_3964,N_3738,N_3726);
and U3965 (N_3965,N_3708,N_3867);
xnor U3966 (N_3966,N_3695,N_3641);
xor U3967 (N_3967,N_3879,N_3638);
nor U3968 (N_3968,N_3620,N_3696);
xnor U3969 (N_3969,N_3698,N_3630);
xor U3970 (N_3970,N_3899,N_3699);
and U3971 (N_3971,N_3782,N_3754);
xor U3972 (N_3972,N_3768,N_3753);
or U3973 (N_3973,N_3772,N_3752);
nand U3974 (N_3974,N_3773,N_3731);
nor U3975 (N_3975,N_3621,N_3650);
xor U3976 (N_3976,N_3608,N_3769);
or U3977 (N_3977,N_3874,N_3868);
nand U3978 (N_3978,N_3614,N_3894);
nand U3979 (N_3979,N_3720,N_3882);
and U3980 (N_3980,N_3841,N_3603);
or U3981 (N_3981,N_3775,N_3824);
and U3982 (N_3982,N_3743,N_3881);
nand U3983 (N_3983,N_3605,N_3624);
nand U3984 (N_3984,N_3833,N_3857);
xnor U3985 (N_3985,N_3767,N_3846);
nor U3986 (N_3986,N_3842,N_3642);
and U3987 (N_3987,N_3851,N_3611);
nor U3988 (N_3988,N_3732,N_3883);
or U3989 (N_3989,N_3849,N_3797);
nand U3990 (N_3990,N_3694,N_3788);
nand U3991 (N_3991,N_3623,N_3817);
nand U3992 (N_3992,N_3774,N_3686);
and U3993 (N_3993,N_3778,N_3892);
xor U3994 (N_3994,N_3856,N_3701);
or U3995 (N_3995,N_3728,N_3600);
and U3996 (N_3996,N_3827,N_3657);
nand U3997 (N_3997,N_3799,N_3619);
nand U3998 (N_3998,N_3765,N_3723);
or U3999 (N_3999,N_3651,N_3725);
or U4000 (N_4000,N_3742,N_3803);
and U4001 (N_4001,N_3702,N_3890);
nand U4002 (N_4002,N_3661,N_3771);
and U4003 (N_4003,N_3670,N_3891);
nand U4004 (N_4004,N_3885,N_3805);
or U4005 (N_4005,N_3643,N_3711);
or U4006 (N_4006,N_3761,N_3866);
nor U4007 (N_4007,N_3658,N_3618);
nor U4008 (N_4008,N_3693,N_3675);
xor U4009 (N_4009,N_3678,N_3812);
or U4010 (N_4010,N_3806,N_3709);
nand U4011 (N_4011,N_3818,N_3855);
or U4012 (N_4012,N_3665,N_3671);
nor U4013 (N_4013,N_3721,N_3819);
nand U4014 (N_4014,N_3755,N_3808);
nand U4015 (N_4015,N_3766,N_3848);
nand U4016 (N_4016,N_3654,N_3897);
xnor U4017 (N_4017,N_3664,N_3795);
nor U4018 (N_4018,N_3762,N_3757);
or U4019 (N_4019,N_3869,N_3791);
xnor U4020 (N_4020,N_3636,N_3727);
xnor U4021 (N_4021,N_3796,N_3672);
and U4022 (N_4022,N_3640,N_3655);
or U4023 (N_4023,N_3601,N_3613);
xor U4024 (N_4024,N_3872,N_3645);
nand U4025 (N_4025,N_3828,N_3825);
xor U4026 (N_4026,N_3714,N_3878);
and U4027 (N_4027,N_3622,N_3649);
or U4028 (N_4028,N_3875,N_3758);
xnor U4029 (N_4029,N_3863,N_3860);
xor U4030 (N_4030,N_3666,N_3896);
nor U4031 (N_4031,N_3836,N_3715);
and U4032 (N_4032,N_3843,N_3776);
and U4033 (N_4033,N_3835,N_3607);
nor U4034 (N_4034,N_3854,N_3759);
nor U4035 (N_4035,N_3889,N_3612);
nand U4036 (N_4036,N_3895,N_3706);
nand U4037 (N_4037,N_3737,N_3779);
or U4038 (N_4038,N_3719,N_3615);
or U4039 (N_4039,N_3679,N_3787);
and U4040 (N_4040,N_3802,N_3704);
and U4041 (N_4041,N_3794,N_3876);
nor U4042 (N_4042,N_3662,N_3756);
or U4043 (N_4043,N_3635,N_3821);
nor U4044 (N_4044,N_3747,N_3877);
or U4045 (N_4045,N_3898,N_3644);
xor U4046 (N_4046,N_3886,N_3629);
nand U4047 (N_4047,N_3815,N_3659);
xor U4048 (N_4048,N_3746,N_3634);
or U4049 (N_4049,N_3873,N_3680);
nand U4050 (N_4050,N_3768,N_3873);
xor U4051 (N_4051,N_3701,N_3688);
nand U4052 (N_4052,N_3684,N_3618);
and U4053 (N_4053,N_3775,N_3751);
nor U4054 (N_4054,N_3645,N_3714);
xnor U4055 (N_4055,N_3843,N_3866);
and U4056 (N_4056,N_3622,N_3783);
nor U4057 (N_4057,N_3605,N_3736);
xnor U4058 (N_4058,N_3688,N_3630);
or U4059 (N_4059,N_3724,N_3781);
and U4060 (N_4060,N_3849,N_3739);
nand U4061 (N_4061,N_3656,N_3660);
nor U4062 (N_4062,N_3691,N_3607);
xor U4063 (N_4063,N_3867,N_3680);
nor U4064 (N_4064,N_3795,N_3721);
nand U4065 (N_4065,N_3807,N_3646);
nor U4066 (N_4066,N_3693,N_3834);
xor U4067 (N_4067,N_3673,N_3798);
nand U4068 (N_4068,N_3668,N_3772);
or U4069 (N_4069,N_3749,N_3815);
nand U4070 (N_4070,N_3696,N_3836);
or U4071 (N_4071,N_3723,N_3716);
or U4072 (N_4072,N_3868,N_3622);
nand U4073 (N_4073,N_3823,N_3876);
and U4074 (N_4074,N_3882,N_3739);
nor U4075 (N_4075,N_3829,N_3679);
nor U4076 (N_4076,N_3717,N_3605);
or U4077 (N_4077,N_3893,N_3685);
nor U4078 (N_4078,N_3666,N_3851);
and U4079 (N_4079,N_3762,N_3702);
nor U4080 (N_4080,N_3707,N_3799);
nand U4081 (N_4081,N_3796,N_3828);
nand U4082 (N_4082,N_3798,N_3716);
and U4083 (N_4083,N_3662,N_3635);
xor U4084 (N_4084,N_3682,N_3830);
nand U4085 (N_4085,N_3620,N_3782);
nor U4086 (N_4086,N_3743,N_3728);
and U4087 (N_4087,N_3793,N_3711);
and U4088 (N_4088,N_3706,N_3861);
or U4089 (N_4089,N_3776,N_3675);
and U4090 (N_4090,N_3896,N_3647);
nand U4091 (N_4091,N_3702,N_3761);
xnor U4092 (N_4092,N_3737,N_3686);
xor U4093 (N_4093,N_3626,N_3819);
nand U4094 (N_4094,N_3756,N_3745);
nand U4095 (N_4095,N_3758,N_3814);
nand U4096 (N_4096,N_3636,N_3627);
or U4097 (N_4097,N_3834,N_3705);
and U4098 (N_4098,N_3827,N_3638);
nor U4099 (N_4099,N_3815,N_3820);
or U4100 (N_4100,N_3826,N_3688);
nor U4101 (N_4101,N_3833,N_3677);
xor U4102 (N_4102,N_3699,N_3665);
nand U4103 (N_4103,N_3869,N_3765);
xnor U4104 (N_4104,N_3691,N_3868);
or U4105 (N_4105,N_3716,N_3670);
and U4106 (N_4106,N_3638,N_3646);
xnor U4107 (N_4107,N_3782,N_3768);
nand U4108 (N_4108,N_3862,N_3813);
and U4109 (N_4109,N_3711,N_3691);
nor U4110 (N_4110,N_3756,N_3755);
and U4111 (N_4111,N_3611,N_3792);
or U4112 (N_4112,N_3660,N_3603);
xor U4113 (N_4113,N_3648,N_3785);
and U4114 (N_4114,N_3702,N_3716);
or U4115 (N_4115,N_3754,N_3631);
xnor U4116 (N_4116,N_3643,N_3738);
nor U4117 (N_4117,N_3790,N_3647);
or U4118 (N_4118,N_3643,N_3748);
or U4119 (N_4119,N_3694,N_3806);
xnor U4120 (N_4120,N_3723,N_3671);
nand U4121 (N_4121,N_3885,N_3740);
nor U4122 (N_4122,N_3805,N_3858);
nor U4123 (N_4123,N_3852,N_3851);
nor U4124 (N_4124,N_3665,N_3803);
or U4125 (N_4125,N_3855,N_3692);
nand U4126 (N_4126,N_3824,N_3825);
and U4127 (N_4127,N_3685,N_3871);
nand U4128 (N_4128,N_3617,N_3716);
and U4129 (N_4129,N_3823,N_3849);
and U4130 (N_4130,N_3729,N_3865);
and U4131 (N_4131,N_3887,N_3686);
xnor U4132 (N_4132,N_3791,N_3836);
nor U4133 (N_4133,N_3687,N_3755);
nand U4134 (N_4134,N_3811,N_3678);
and U4135 (N_4135,N_3709,N_3743);
nand U4136 (N_4136,N_3752,N_3753);
nor U4137 (N_4137,N_3717,N_3657);
xor U4138 (N_4138,N_3858,N_3816);
and U4139 (N_4139,N_3720,N_3788);
or U4140 (N_4140,N_3657,N_3795);
nand U4141 (N_4141,N_3881,N_3696);
nor U4142 (N_4142,N_3666,N_3752);
nor U4143 (N_4143,N_3645,N_3741);
and U4144 (N_4144,N_3645,N_3722);
and U4145 (N_4145,N_3794,N_3855);
nand U4146 (N_4146,N_3699,N_3613);
and U4147 (N_4147,N_3614,N_3656);
xnor U4148 (N_4148,N_3837,N_3784);
and U4149 (N_4149,N_3625,N_3797);
and U4150 (N_4150,N_3850,N_3681);
xnor U4151 (N_4151,N_3804,N_3864);
nand U4152 (N_4152,N_3608,N_3883);
nor U4153 (N_4153,N_3664,N_3723);
or U4154 (N_4154,N_3808,N_3868);
or U4155 (N_4155,N_3867,N_3697);
nand U4156 (N_4156,N_3600,N_3655);
or U4157 (N_4157,N_3679,N_3730);
nand U4158 (N_4158,N_3868,N_3781);
nor U4159 (N_4159,N_3763,N_3735);
nand U4160 (N_4160,N_3710,N_3753);
or U4161 (N_4161,N_3717,N_3785);
nor U4162 (N_4162,N_3843,N_3605);
xor U4163 (N_4163,N_3841,N_3834);
xnor U4164 (N_4164,N_3650,N_3807);
or U4165 (N_4165,N_3760,N_3884);
xor U4166 (N_4166,N_3661,N_3667);
or U4167 (N_4167,N_3651,N_3753);
nor U4168 (N_4168,N_3808,N_3794);
nand U4169 (N_4169,N_3839,N_3642);
nand U4170 (N_4170,N_3716,N_3792);
or U4171 (N_4171,N_3609,N_3711);
or U4172 (N_4172,N_3764,N_3672);
nor U4173 (N_4173,N_3849,N_3805);
xor U4174 (N_4174,N_3735,N_3897);
nand U4175 (N_4175,N_3627,N_3840);
xnor U4176 (N_4176,N_3807,N_3781);
and U4177 (N_4177,N_3616,N_3661);
or U4178 (N_4178,N_3600,N_3742);
and U4179 (N_4179,N_3861,N_3898);
or U4180 (N_4180,N_3868,N_3659);
nor U4181 (N_4181,N_3732,N_3684);
nor U4182 (N_4182,N_3636,N_3680);
and U4183 (N_4183,N_3713,N_3635);
or U4184 (N_4184,N_3845,N_3836);
nor U4185 (N_4185,N_3643,N_3697);
xor U4186 (N_4186,N_3696,N_3880);
nand U4187 (N_4187,N_3759,N_3685);
nor U4188 (N_4188,N_3608,N_3641);
nor U4189 (N_4189,N_3692,N_3711);
and U4190 (N_4190,N_3869,N_3838);
or U4191 (N_4191,N_3858,N_3813);
or U4192 (N_4192,N_3744,N_3666);
nand U4193 (N_4193,N_3707,N_3814);
or U4194 (N_4194,N_3784,N_3624);
or U4195 (N_4195,N_3654,N_3683);
nor U4196 (N_4196,N_3894,N_3886);
xnor U4197 (N_4197,N_3828,N_3642);
or U4198 (N_4198,N_3738,N_3673);
and U4199 (N_4199,N_3865,N_3649);
and U4200 (N_4200,N_4191,N_4184);
xnor U4201 (N_4201,N_4125,N_4085);
xor U4202 (N_4202,N_4162,N_4012);
nor U4203 (N_4203,N_4106,N_4021);
or U4204 (N_4204,N_4047,N_4152);
nor U4205 (N_4205,N_4182,N_3988);
and U4206 (N_4206,N_4010,N_4108);
or U4207 (N_4207,N_4151,N_3980);
or U4208 (N_4208,N_4006,N_3901);
nor U4209 (N_4209,N_3977,N_4019);
nand U4210 (N_4210,N_3995,N_4079);
nor U4211 (N_4211,N_4144,N_4103);
nand U4212 (N_4212,N_3904,N_3942);
or U4213 (N_4213,N_4175,N_4163);
nor U4214 (N_4214,N_3998,N_3951);
or U4215 (N_4215,N_3919,N_4008);
or U4216 (N_4216,N_3950,N_3996);
and U4217 (N_4217,N_4137,N_4114);
xnor U4218 (N_4218,N_3931,N_4068);
nor U4219 (N_4219,N_4084,N_4189);
and U4220 (N_4220,N_4029,N_4030);
nand U4221 (N_4221,N_3955,N_4015);
xnor U4222 (N_4222,N_4093,N_4009);
nor U4223 (N_4223,N_4195,N_4073);
nand U4224 (N_4224,N_4028,N_4109);
nand U4225 (N_4225,N_3908,N_3911);
nor U4226 (N_4226,N_3945,N_3935);
nand U4227 (N_4227,N_3905,N_4132);
nand U4228 (N_4228,N_4027,N_3994);
nand U4229 (N_4229,N_4198,N_4026);
xnor U4230 (N_4230,N_3913,N_4062);
nor U4231 (N_4231,N_4120,N_3915);
nand U4232 (N_4232,N_4098,N_3979);
nor U4233 (N_4233,N_4080,N_4142);
nor U4234 (N_4234,N_4083,N_4116);
xnor U4235 (N_4235,N_3933,N_4178);
xnor U4236 (N_4236,N_4075,N_3938);
xor U4237 (N_4237,N_4183,N_4122);
nand U4238 (N_4238,N_4007,N_4065);
nor U4239 (N_4239,N_3906,N_3940);
nand U4240 (N_4240,N_4131,N_4089);
or U4241 (N_4241,N_4092,N_3964);
nor U4242 (N_4242,N_4104,N_4154);
nor U4243 (N_4243,N_4034,N_4164);
xor U4244 (N_4244,N_4000,N_4158);
xnor U4245 (N_4245,N_4051,N_4173);
or U4246 (N_4246,N_4038,N_4128);
nor U4247 (N_4247,N_3963,N_4039);
xnor U4248 (N_4248,N_3927,N_3917);
or U4249 (N_4249,N_4139,N_4107);
nand U4250 (N_4250,N_3936,N_3986);
nor U4251 (N_4251,N_3972,N_4172);
xnor U4252 (N_4252,N_4035,N_4072);
or U4253 (N_4253,N_3989,N_4159);
xnor U4254 (N_4254,N_4135,N_3944);
or U4255 (N_4255,N_3999,N_3921);
nand U4256 (N_4256,N_4003,N_4196);
or U4257 (N_4257,N_4123,N_4187);
and U4258 (N_4258,N_3953,N_4001);
nor U4259 (N_4259,N_4186,N_4060);
or U4260 (N_4260,N_4024,N_4117);
and U4261 (N_4261,N_3984,N_4077);
xor U4262 (N_4262,N_4022,N_4168);
nand U4263 (N_4263,N_3907,N_3903);
nand U4264 (N_4264,N_4097,N_3914);
or U4265 (N_4265,N_3956,N_4059);
and U4266 (N_4266,N_4004,N_3966);
and U4267 (N_4267,N_4129,N_3971);
and U4268 (N_4268,N_4005,N_4160);
and U4269 (N_4269,N_3910,N_4161);
nor U4270 (N_4270,N_4181,N_4145);
and U4271 (N_4271,N_4100,N_3923);
nand U4272 (N_4272,N_3968,N_4043);
or U4273 (N_4273,N_4141,N_4091);
or U4274 (N_4274,N_4094,N_3990);
nor U4275 (N_4275,N_4112,N_3928);
and U4276 (N_4276,N_4165,N_4190);
or U4277 (N_4277,N_3946,N_3929);
nor U4278 (N_4278,N_3900,N_4121);
or U4279 (N_4279,N_3987,N_3932);
nor U4280 (N_4280,N_3974,N_3969);
and U4281 (N_4281,N_3973,N_4052);
or U4282 (N_4282,N_3912,N_3937);
xor U4283 (N_4283,N_3952,N_4110);
nand U4284 (N_4284,N_4033,N_4067);
and U4285 (N_4285,N_3902,N_4082);
or U4286 (N_4286,N_4048,N_4115);
nor U4287 (N_4287,N_3941,N_4179);
and U4288 (N_4288,N_4188,N_3967);
nor U4289 (N_4289,N_4076,N_4101);
nand U4290 (N_4290,N_4055,N_4090);
xor U4291 (N_4291,N_3959,N_4025);
or U4292 (N_4292,N_4031,N_4197);
nand U4293 (N_4293,N_4049,N_3957);
or U4294 (N_4294,N_3922,N_3965);
nand U4295 (N_4295,N_4119,N_4011);
or U4296 (N_4296,N_4053,N_4126);
nand U4297 (N_4297,N_4061,N_4037);
xnor U4298 (N_4298,N_4177,N_4199);
or U4299 (N_4299,N_4018,N_4078);
nor U4300 (N_4300,N_4113,N_3991);
and U4301 (N_4301,N_4020,N_3954);
and U4302 (N_4302,N_3983,N_3939);
nand U4303 (N_4303,N_4130,N_4124);
or U4304 (N_4304,N_3926,N_4118);
nand U4305 (N_4305,N_3943,N_4111);
and U4306 (N_4306,N_4002,N_3924);
xnor U4307 (N_4307,N_4074,N_4180);
or U4308 (N_4308,N_4134,N_3970);
and U4309 (N_4309,N_3982,N_4167);
xnor U4310 (N_4310,N_4127,N_3918);
and U4311 (N_4311,N_4157,N_3920);
or U4312 (N_4312,N_3975,N_4050);
xor U4313 (N_4313,N_4169,N_4174);
and U4314 (N_4314,N_4176,N_4042);
nand U4315 (N_4315,N_3948,N_4086);
xor U4316 (N_4316,N_4040,N_4099);
and U4317 (N_4317,N_4140,N_3992);
or U4318 (N_4318,N_4194,N_4096);
or U4319 (N_4319,N_4063,N_3949);
nand U4320 (N_4320,N_4170,N_4192);
nand U4321 (N_4321,N_4166,N_3976);
nand U4322 (N_4322,N_4155,N_4058);
nand U4323 (N_4323,N_4148,N_3930);
and U4324 (N_4324,N_4046,N_4014);
xor U4325 (N_4325,N_4044,N_4071);
nor U4326 (N_4326,N_4069,N_4066);
and U4327 (N_4327,N_4171,N_4017);
and U4328 (N_4328,N_4133,N_3962);
or U4329 (N_4329,N_4036,N_3993);
nand U4330 (N_4330,N_3925,N_4057);
xor U4331 (N_4331,N_4045,N_3985);
xnor U4332 (N_4332,N_3981,N_3934);
nor U4333 (N_4333,N_4150,N_4087);
nor U4334 (N_4334,N_4032,N_3909);
and U4335 (N_4335,N_4185,N_3916);
xor U4336 (N_4336,N_4146,N_4095);
nand U4337 (N_4337,N_4153,N_3958);
and U4338 (N_4338,N_4054,N_4070);
xor U4339 (N_4339,N_3947,N_4056);
xnor U4340 (N_4340,N_3997,N_3978);
xor U4341 (N_4341,N_4143,N_4088);
xnor U4342 (N_4342,N_3961,N_4016);
and U4343 (N_4343,N_4193,N_4102);
nor U4344 (N_4344,N_4013,N_4081);
nand U4345 (N_4345,N_4138,N_4136);
and U4346 (N_4346,N_4149,N_4023);
nand U4347 (N_4347,N_3960,N_4147);
nor U4348 (N_4348,N_4105,N_4041);
or U4349 (N_4349,N_4156,N_4064);
and U4350 (N_4350,N_3971,N_3951);
and U4351 (N_4351,N_4165,N_4184);
or U4352 (N_4352,N_4156,N_4116);
xnor U4353 (N_4353,N_4159,N_3978);
nand U4354 (N_4354,N_4017,N_3978);
xnor U4355 (N_4355,N_3924,N_4198);
nand U4356 (N_4356,N_3955,N_3974);
or U4357 (N_4357,N_4004,N_4027);
or U4358 (N_4358,N_3963,N_4095);
or U4359 (N_4359,N_4177,N_3984);
nor U4360 (N_4360,N_3991,N_3992);
or U4361 (N_4361,N_3914,N_4017);
nand U4362 (N_4362,N_4142,N_4157);
nor U4363 (N_4363,N_3963,N_4064);
nor U4364 (N_4364,N_4181,N_4059);
or U4365 (N_4365,N_4188,N_4047);
nor U4366 (N_4366,N_4145,N_4052);
nor U4367 (N_4367,N_3938,N_3940);
nand U4368 (N_4368,N_4044,N_3960);
xnor U4369 (N_4369,N_3961,N_3988);
or U4370 (N_4370,N_4107,N_4067);
xnor U4371 (N_4371,N_3987,N_4194);
or U4372 (N_4372,N_4198,N_4115);
xnor U4373 (N_4373,N_3925,N_4016);
and U4374 (N_4374,N_4086,N_4075);
xor U4375 (N_4375,N_4134,N_3974);
or U4376 (N_4376,N_3960,N_4030);
nor U4377 (N_4377,N_4127,N_4016);
and U4378 (N_4378,N_4090,N_4078);
or U4379 (N_4379,N_3905,N_4131);
xor U4380 (N_4380,N_4132,N_4009);
or U4381 (N_4381,N_3907,N_4031);
or U4382 (N_4382,N_4001,N_4155);
or U4383 (N_4383,N_4186,N_4149);
xor U4384 (N_4384,N_4003,N_3927);
and U4385 (N_4385,N_4170,N_4083);
and U4386 (N_4386,N_3917,N_4009);
nor U4387 (N_4387,N_4193,N_3976);
xnor U4388 (N_4388,N_4103,N_3942);
and U4389 (N_4389,N_4098,N_3967);
and U4390 (N_4390,N_4080,N_4070);
nand U4391 (N_4391,N_4191,N_4006);
or U4392 (N_4392,N_4149,N_4138);
nor U4393 (N_4393,N_3949,N_3919);
nand U4394 (N_4394,N_3971,N_3944);
nand U4395 (N_4395,N_4144,N_3942);
or U4396 (N_4396,N_4194,N_4078);
or U4397 (N_4397,N_4198,N_4129);
xor U4398 (N_4398,N_3989,N_4017);
xor U4399 (N_4399,N_4060,N_4108);
nor U4400 (N_4400,N_4011,N_4080);
nor U4401 (N_4401,N_4160,N_4094);
and U4402 (N_4402,N_4031,N_4018);
xnor U4403 (N_4403,N_4034,N_4057);
and U4404 (N_4404,N_3950,N_3908);
nand U4405 (N_4405,N_4174,N_4021);
and U4406 (N_4406,N_3953,N_4088);
nor U4407 (N_4407,N_3992,N_4094);
nand U4408 (N_4408,N_4067,N_4196);
nor U4409 (N_4409,N_4102,N_3968);
nor U4410 (N_4410,N_3902,N_3970);
xnor U4411 (N_4411,N_4044,N_3948);
or U4412 (N_4412,N_3904,N_4091);
xnor U4413 (N_4413,N_4072,N_3911);
and U4414 (N_4414,N_4002,N_3991);
or U4415 (N_4415,N_3921,N_4120);
nor U4416 (N_4416,N_4002,N_3973);
and U4417 (N_4417,N_4183,N_4164);
nor U4418 (N_4418,N_3950,N_3965);
nand U4419 (N_4419,N_3901,N_4013);
nand U4420 (N_4420,N_3954,N_4024);
nor U4421 (N_4421,N_4134,N_3975);
and U4422 (N_4422,N_4009,N_4163);
or U4423 (N_4423,N_4072,N_4064);
nand U4424 (N_4424,N_3986,N_4116);
and U4425 (N_4425,N_3973,N_4011);
nor U4426 (N_4426,N_4023,N_3949);
nand U4427 (N_4427,N_3918,N_4000);
and U4428 (N_4428,N_3990,N_4128);
or U4429 (N_4429,N_4157,N_3932);
nand U4430 (N_4430,N_4117,N_4033);
and U4431 (N_4431,N_4119,N_3968);
and U4432 (N_4432,N_3931,N_3916);
nand U4433 (N_4433,N_4015,N_4004);
xor U4434 (N_4434,N_4077,N_3914);
nor U4435 (N_4435,N_4112,N_3985);
nand U4436 (N_4436,N_4075,N_3941);
xor U4437 (N_4437,N_3989,N_4190);
and U4438 (N_4438,N_4005,N_4051);
nor U4439 (N_4439,N_4024,N_4186);
nor U4440 (N_4440,N_3937,N_4018);
and U4441 (N_4441,N_4092,N_4051);
and U4442 (N_4442,N_3928,N_4181);
and U4443 (N_4443,N_3936,N_4075);
or U4444 (N_4444,N_4065,N_3902);
xor U4445 (N_4445,N_3998,N_3985);
and U4446 (N_4446,N_4105,N_4160);
xnor U4447 (N_4447,N_4004,N_3905);
nor U4448 (N_4448,N_3926,N_4143);
nor U4449 (N_4449,N_3992,N_4027);
xor U4450 (N_4450,N_3966,N_3982);
xor U4451 (N_4451,N_4168,N_4057);
xor U4452 (N_4452,N_4081,N_4038);
xor U4453 (N_4453,N_3900,N_4155);
nand U4454 (N_4454,N_4026,N_3955);
nand U4455 (N_4455,N_4120,N_3968);
nor U4456 (N_4456,N_3943,N_4163);
and U4457 (N_4457,N_3947,N_3915);
nand U4458 (N_4458,N_4083,N_4010);
and U4459 (N_4459,N_3907,N_3957);
nor U4460 (N_4460,N_3935,N_3913);
nor U4461 (N_4461,N_4011,N_4041);
or U4462 (N_4462,N_3909,N_4096);
xor U4463 (N_4463,N_4077,N_3975);
nand U4464 (N_4464,N_4057,N_4037);
xor U4465 (N_4465,N_4170,N_4126);
xor U4466 (N_4466,N_4005,N_4129);
nand U4467 (N_4467,N_4105,N_4016);
or U4468 (N_4468,N_4091,N_3910);
and U4469 (N_4469,N_4112,N_4075);
xnor U4470 (N_4470,N_3971,N_4153);
nor U4471 (N_4471,N_4001,N_4176);
or U4472 (N_4472,N_4055,N_3928);
nand U4473 (N_4473,N_4095,N_3948);
xor U4474 (N_4474,N_4043,N_4073);
nand U4475 (N_4475,N_4017,N_4125);
xor U4476 (N_4476,N_3918,N_3917);
and U4477 (N_4477,N_4126,N_4166);
nand U4478 (N_4478,N_3921,N_4044);
nand U4479 (N_4479,N_3976,N_4062);
xnor U4480 (N_4480,N_4112,N_4042);
nand U4481 (N_4481,N_4158,N_3952);
and U4482 (N_4482,N_4129,N_4007);
or U4483 (N_4483,N_4104,N_4085);
or U4484 (N_4484,N_3976,N_4135);
nand U4485 (N_4485,N_4041,N_3964);
and U4486 (N_4486,N_3950,N_4023);
xor U4487 (N_4487,N_3935,N_3984);
nand U4488 (N_4488,N_4006,N_4115);
xnor U4489 (N_4489,N_3920,N_4172);
and U4490 (N_4490,N_4019,N_4172);
nor U4491 (N_4491,N_4038,N_4144);
and U4492 (N_4492,N_4047,N_4005);
nor U4493 (N_4493,N_4151,N_4126);
xor U4494 (N_4494,N_3913,N_4027);
or U4495 (N_4495,N_4009,N_3907);
nor U4496 (N_4496,N_4097,N_3995);
or U4497 (N_4497,N_4133,N_3932);
nor U4498 (N_4498,N_4069,N_4125);
xor U4499 (N_4499,N_4084,N_4079);
or U4500 (N_4500,N_4337,N_4410);
nor U4501 (N_4501,N_4288,N_4426);
and U4502 (N_4502,N_4304,N_4283);
and U4503 (N_4503,N_4313,N_4282);
nor U4504 (N_4504,N_4256,N_4390);
or U4505 (N_4505,N_4420,N_4305);
xor U4506 (N_4506,N_4472,N_4280);
nor U4507 (N_4507,N_4306,N_4269);
nor U4508 (N_4508,N_4348,N_4308);
or U4509 (N_4509,N_4315,N_4419);
or U4510 (N_4510,N_4376,N_4260);
or U4511 (N_4511,N_4486,N_4251);
nor U4512 (N_4512,N_4298,N_4445);
xnor U4513 (N_4513,N_4401,N_4201);
nand U4514 (N_4514,N_4385,N_4292);
or U4515 (N_4515,N_4415,N_4205);
and U4516 (N_4516,N_4229,N_4342);
nand U4517 (N_4517,N_4258,N_4244);
xnor U4518 (N_4518,N_4365,N_4370);
xor U4519 (N_4519,N_4466,N_4249);
or U4520 (N_4520,N_4465,N_4446);
nand U4521 (N_4521,N_4477,N_4443);
xor U4522 (N_4522,N_4338,N_4356);
and U4523 (N_4523,N_4469,N_4448);
nor U4524 (N_4524,N_4276,N_4203);
and U4525 (N_4525,N_4450,N_4422);
or U4526 (N_4526,N_4362,N_4257);
nor U4527 (N_4527,N_4470,N_4271);
xor U4528 (N_4528,N_4206,N_4263);
or U4529 (N_4529,N_4346,N_4393);
nor U4530 (N_4530,N_4418,N_4232);
and U4531 (N_4531,N_4495,N_4382);
and U4532 (N_4532,N_4303,N_4235);
nor U4533 (N_4533,N_4440,N_4319);
or U4534 (N_4534,N_4293,N_4333);
nand U4535 (N_4535,N_4241,N_4457);
xor U4536 (N_4536,N_4468,N_4312);
nor U4537 (N_4537,N_4444,N_4275);
nand U4538 (N_4538,N_4334,N_4340);
nor U4539 (N_4539,N_4279,N_4259);
and U4540 (N_4540,N_4374,N_4291);
nand U4541 (N_4541,N_4322,N_4460);
xnor U4542 (N_4542,N_4364,N_4451);
and U4543 (N_4543,N_4217,N_4476);
and U4544 (N_4544,N_4243,N_4351);
and U4545 (N_4545,N_4246,N_4408);
or U4546 (N_4546,N_4454,N_4341);
and U4547 (N_4547,N_4371,N_4361);
nor U4548 (N_4548,N_4358,N_4483);
nand U4549 (N_4549,N_4473,N_4392);
nor U4550 (N_4550,N_4383,N_4219);
and U4551 (N_4551,N_4388,N_4377);
nand U4552 (N_4552,N_4265,N_4350);
xor U4553 (N_4553,N_4368,N_4210);
or U4554 (N_4554,N_4421,N_4327);
nor U4555 (N_4555,N_4406,N_4359);
nor U4556 (N_4556,N_4387,N_4266);
nor U4557 (N_4557,N_4287,N_4498);
nand U4558 (N_4558,N_4496,N_4449);
nand U4559 (N_4559,N_4300,N_4435);
and U4560 (N_4560,N_4253,N_4238);
or U4561 (N_4561,N_4400,N_4321);
and U4562 (N_4562,N_4455,N_4428);
and U4563 (N_4563,N_4230,N_4429);
xnor U4564 (N_4564,N_4492,N_4307);
nand U4565 (N_4565,N_4297,N_4237);
and U4566 (N_4566,N_4480,N_4438);
nor U4567 (N_4567,N_4325,N_4414);
xor U4568 (N_4568,N_4336,N_4234);
nor U4569 (N_4569,N_4310,N_4441);
nand U4570 (N_4570,N_4360,N_4458);
and U4571 (N_4571,N_4270,N_4326);
and U4572 (N_4572,N_4424,N_4323);
nor U4573 (N_4573,N_4431,N_4425);
nand U4574 (N_4574,N_4459,N_4286);
xor U4575 (N_4575,N_4335,N_4309);
nor U4576 (N_4576,N_4373,N_4491);
nand U4577 (N_4577,N_4343,N_4273);
nor U4578 (N_4578,N_4233,N_4290);
nor U4579 (N_4579,N_4467,N_4225);
xnor U4580 (N_4580,N_4404,N_4231);
nand U4581 (N_4581,N_4284,N_4324);
and U4582 (N_4582,N_4433,N_4484);
and U4583 (N_4583,N_4316,N_4320);
nand U4584 (N_4584,N_4239,N_4411);
or U4585 (N_4585,N_4452,N_4281);
xnor U4586 (N_4586,N_4436,N_4499);
nor U4587 (N_4587,N_4437,N_4430);
or U4588 (N_4588,N_4240,N_4366);
nor U4589 (N_4589,N_4395,N_4353);
nor U4590 (N_4590,N_4223,N_4481);
or U4591 (N_4591,N_4255,N_4345);
nand U4592 (N_4592,N_4434,N_4349);
and U4593 (N_4593,N_4407,N_4478);
nor U4594 (N_4594,N_4453,N_4221);
nand U4595 (N_4595,N_4285,N_4427);
and U4596 (N_4596,N_4222,N_4216);
or U4597 (N_4597,N_4208,N_4236);
xor U4598 (N_4598,N_4482,N_4215);
xor U4599 (N_4599,N_4367,N_4250);
nor U4600 (N_4600,N_4295,N_4242);
nor U4601 (N_4601,N_4226,N_4254);
xnor U4602 (N_4602,N_4227,N_4369);
or U4603 (N_4603,N_4212,N_4296);
nor U4604 (N_4604,N_4299,N_4442);
xor U4605 (N_4605,N_4409,N_4248);
xor U4606 (N_4606,N_4261,N_4267);
nand U4607 (N_4607,N_4456,N_4403);
nor U4608 (N_4608,N_4294,N_4494);
xnor U4609 (N_4609,N_4352,N_4463);
and U4610 (N_4610,N_4372,N_4471);
nand U4611 (N_4611,N_4375,N_4493);
nand U4612 (N_4612,N_4489,N_4354);
nor U4613 (N_4613,N_4416,N_4397);
and U4614 (N_4614,N_4207,N_4423);
xor U4615 (N_4615,N_4490,N_4462);
and U4616 (N_4616,N_4380,N_4432);
or U4617 (N_4617,N_4417,N_4413);
nor U4618 (N_4618,N_4202,N_4487);
and U4619 (N_4619,N_4314,N_4301);
or U4620 (N_4620,N_4497,N_4330);
or U4621 (N_4621,N_4398,N_4220);
nor U4622 (N_4622,N_4347,N_4381);
or U4623 (N_4623,N_4389,N_4209);
or U4624 (N_4624,N_4268,N_4332);
xor U4625 (N_4625,N_4344,N_4379);
nand U4626 (N_4626,N_4384,N_4224);
xor U4627 (N_4627,N_4214,N_4204);
nand U4628 (N_4628,N_4399,N_4339);
or U4629 (N_4629,N_4252,N_4311);
or U4630 (N_4630,N_4474,N_4247);
or U4631 (N_4631,N_4405,N_4488);
or U4632 (N_4632,N_4302,N_4386);
xnor U4633 (N_4633,N_4363,N_4264);
nand U4634 (N_4634,N_4200,N_4213);
and U4635 (N_4635,N_4412,N_4262);
xnor U4636 (N_4636,N_4289,N_4391);
and U4637 (N_4637,N_4479,N_4447);
and U4638 (N_4638,N_4464,N_4439);
or U4639 (N_4639,N_4329,N_4475);
nand U4640 (N_4640,N_4396,N_4461);
nor U4641 (N_4641,N_4278,N_4355);
nand U4642 (N_4642,N_4318,N_4218);
nand U4643 (N_4643,N_4485,N_4394);
or U4644 (N_4644,N_4211,N_4228);
nand U4645 (N_4645,N_4317,N_4274);
xnor U4646 (N_4646,N_4357,N_4328);
or U4647 (N_4647,N_4245,N_4331);
or U4648 (N_4648,N_4378,N_4272);
xor U4649 (N_4649,N_4277,N_4402);
nand U4650 (N_4650,N_4459,N_4277);
and U4651 (N_4651,N_4240,N_4238);
nor U4652 (N_4652,N_4421,N_4312);
or U4653 (N_4653,N_4276,N_4438);
and U4654 (N_4654,N_4395,N_4374);
and U4655 (N_4655,N_4380,N_4409);
or U4656 (N_4656,N_4400,N_4402);
xnor U4657 (N_4657,N_4280,N_4411);
and U4658 (N_4658,N_4338,N_4209);
nand U4659 (N_4659,N_4326,N_4491);
nand U4660 (N_4660,N_4224,N_4336);
and U4661 (N_4661,N_4220,N_4468);
nand U4662 (N_4662,N_4379,N_4405);
nand U4663 (N_4663,N_4420,N_4408);
nor U4664 (N_4664,N_4273,N_4481);
or U4665 (N_4665,N_4203,N_4269);
nor U4666 (N_4666,N_4225,N_4344);
and U4667 (N_4667,N_4276,N_4274);
nand U4668 (N_4668,N_4366,N_4411);
xnor U4669 (N_4669,N_4484,N_4465);
xnor U4670 (N_4670,N_4202,N_4279);
or U4671 (N_4671,N_4480,N_4499);
nor U4672 (N_4672,N_4293,N_4393);
nor U4673 (N_4673,N_4379,N_4422);
nor U4674 (N_4674,N_4446,N_4250);
nor U4675 (N_4675,N_4343,N_4203);
nand U4676 (N_4676,N_4212,N_4351);
or U4677 (N_4677,N_4443,N_4372);
nand U4678 (N_4678,N_4401,N_4298);
and U4679 (N_4679,N_4294,N_4474);
nor U4680 (N_4680,N_4497,N_4365);
nand U4681 (N_4681,N_4378,N_4308);
nor U4682 (N_4682,N_4225,N_4480);
and U4683 (N_4683,N_4450,N_4485);
nand U4684 (N_4684,N_4438,N_4397);
nor U4685 (N_4685,N_4317,N_4417);
or U4686 (N_4686,N_4295,N_4200);
nor U4687 (N_4687,N_4466,N_4268);
nor U4688 (N_4688,N_4285,N_4362);
nor U4689 (N_4689,N_4313,N_4433);
xor U4690 (N_4690,N_4268,N_4272);
xnor U4691 (N_4691,N_4219,N_4346);
or U4692 (N_4692,N_4257,N_4484);
xnor U4693 (N_4693,N_4286,N_4321);
xor U4694 (N_4694,N_4296,N_4463);
xnor U4695 (N_4695,N_4337,N_4310);
and U4696 (N_4696,N_4372,N_4462);
nand U4697 (N_4697,N_4484,N_4208);
nand U4698 (N_4698,N_4476,N_4495);
xnor U4699 (N_4699,N_4440,N_4263);
or U4700 (N_4700,N_4437,N_4253);
nor U4701 (N_4701,N_4201,N_4389);
nor U4702 (N_4702,N_4288,N_4308);
nand U4703 (N_4703,N_4477,N_4411);
nand U4704 (N_4704,N_4272,N_4300);
and U4705 (N_4705,N_4432,N_4218);
xnor U4706 (N_4706,N_4239,N_4371);
nor U4707 (N_4707,N_4451,N_4443);
and U4708 (N_4708,N_4407,N_4378);
xor U4709 (N_4709,N_4491,N_4223);
and U4710 (N_4710,N_4446,N_4435);
and U4711 (N_4711,N_4205,N_4369);
nand U4712 (N_4712,N_4364,N_4312);
nor U4713 (N_4713,N_4336,N_4456);
xnor U4714 (N_4714,N_4378,N_4485);
and U4715 (N_4715,N_4480,N_4495);
nand U4716 (N_4716,N_4465,N_4480);
or U4717 (N_4717,N_4494,N_4236);
nor U4718 (N_4718,N_4295,N_4281);
nor U4719 (N_4719,N_4327,N_4427);
xnor U4720 (N_4720,N_4493,N_4278);
and U4721 (N_4721,N_4402,N_4436);
xnor U4722 (N_4722,N_4208,N_4350);
and U4723 (N_4723,N_4466,N_4417);
xnor U4724 (N_4724,N_4264,N_4378);
or U4725 (N_4725,N_4335,N_4372);
nor U4726 (N_4726,N_4234,N_4231);
and U4727 (N_4727,N_4279,N_4244);
nor U4728 (N_4728,N_4344,N_4207);
nand U4729 (N_4729,N_4243,N_4482);
and U4730 (N_4730,N_4291,N_4434);
nand U4731 (N_4731,N_4289,N_4219);
and U4732 (N_4732,N_4317,N_4323);
xnor U4733 (N_4733,N_4257,N_4455);
or U4734 (N_4734,N_4226,N_4330);
or U4735 (N_4735,N_4385,N_4276);
xor U4736 (N_4736,N_4456,N_4213);
nand U4737 (N_4737,N_4210,N_4309);
nand U4738 (N_4738,N_4384,N_4455);
or U4739 (N_4739,N_4263,N_4495);
and U4740 (N_4740,N_4383,N_4387);
nor U4741 (N_4741,N_4424,N_4254);
xnor U4742 (N_4742,N_4379,N_4411);
nand U4743 (N_4743,N_4357,N_4260);
nor U4744 (N_4744,N_4417,N_4412);
nor U4745 (N_4745,N_4271,N_4353);
or U4746 (N_4746,N_4411,N_4213);
xor U4747 (N_4747,N_4316,N_4280);
and U4748 (N_4748,N_4433,N_4432);
nor U4749 (N_4749,N_4236,N_4400);
xor U4750 (N_4750,N_4239,N_4275);
xnor U4751 (N_4751,N_4450,N_4268);
xnor U4752 (N_4752,N_4350,N_4247);
xnor U4753 (N_4753,N_4493,N_4332);
or U4754 (N_4754,N_4418,N_4402);
and U4755 (N_4755,N_4266,N_4378);
and U4756 (N_4756,N_4295,N_4334);
xor U4757 (N_4757,N_4441,N_4256);
and U4758 (N_4758,N_4256,N_4248);
xor U4759 (N_4759,N_4289,N_4317);
nor U4760 (N_4760,N_4415,N_4475);
nand U4761 (N_4761,N_4486,N_4317);
and U4762 (N_4762,N_4445,N_4236);
xnor U4763 (N_4763,N_4434,N_4234);
nor U4764 (N_4764,N_4228,N_4471);
xor U4765 (N_4765,N_4386,N_4203);
nand U4766 (N_4766,N_4348,N_4231);
or U4767 (N_4767,N_4214,N_4231);
or U4768 (N_4768,N_4430,N_4470);
and U4769 (N_4769,N_4244,N_4479);
nand U4770 (N_4770,N_4470,N_4328);
or U4771 (N_4771,N_4249,N_4405);
xor U4772 (N_4772,N_4284,N_4410);
or U4773 (N_4773,N_4417,N_4444);
and U4774 (N_4774,N_4227,N_4261);
xor U4775 (N_4775,N_4296,N_4309);
nand U4776 (N_4776,N_4249,N_4410);
nor U4777 (N_4777,N_4387,N_4414);
or U4778 (N_4778,N_4458,N_4362);
and U4779 (N_4779,N_4482,N_4356);
and U4780 (N_4780,N_4412,N_4238);
or U4781 (N_4781,N_4294,N_4357);
nor U4782 (N_4782,N_4386,N_4262);
nand U4783 (N_4783,N_4386,N_4321);
or U4784 (N_4784,N_4427,N_4433);
xnor U4785 (N_4785,N_4461,N_4310);
and U4786 (N_4786,N_4495,N_4287);
or U4787 (N_4787,N_4348,N_4325);
xnor U4788 (N_4788,N_4289,N_4367);
nand U4789 (N_4789,N_4438,N_4498);
nand U4790 (N_4790,N_4344,N_4282);
or U4791 (N_4791,N_4480,N_4418);
or U4792 (N_4792,N_4271,N_4448);
nand U4793 (N_4793,N_4355,N_4425);
xor U4794 (N_4794,N_4252,N_4436);
nand U4795 (N_4795,N_4411,N_4212);
nor U4796 (N_4796,N_4325,N_4203);
xor U4797 (N_4797,N_4225,N_4462);
nand U4798 (N_4798,N_4202,N_4359);
and U4799 (N_4799,N_4228,N_4282);
xor U4800 (N_4800,N_4625,N_4701);
or U4801 (N_4801,N_4736,N_4654);
and U4802 (N_4802,N_4716,N_4587);
nand U4803 (N_4803,N_4551,N_4526);
nor U4804 (N_4804,N_4776,N_4600);
and U4805 (N_4805,N_4574,N_4616);
nand U4806 (N_4806,N_4764,N_4674);
nor U4807 (N_4807,N_4770,N_4647);
nor U4808 (N_4808,N_4681,N_4698);
xnor U4809 (N_4809,N_4612,N_4718);
nand U4810 (N_4810,N_4753,N_4566);
nor U4811 (N_4811,N_4680,N_4672);
nand U4812 (N_4812,N_4585,N_4638);
nand U4813 (N_4813,N_4735,N_4781);
xor U4814 (N_4814,N_4741,N_4678);
nand U4815 (N_4815,N_4709,N_4529);
and U4816 (N_4816,N_4583,N_4596);
or U4817 (N_4817,N_4729,N_4758);
nor U4818 (N_4818,N_4670,N_4794);
or U4819 (N_4819,N_4584,N_4588);
or U4820 (N_4820,N_4653,N_4514);
nor U4821 (N_4821,N_4541,N_4522);
xor U4822 (N_4822,N_4582,N_4747);
nor U4823 (N_4823,N_4699,N_4534);
or U4824 (N_4824,N_4724,N_4766);
or U4825 (N_4825,N_4501,N_4705);
or U4826 (N_4826,N_4737,N_4604);
xor U4827 (N_4827,N_4704,N_4533);
nor U4828 (N_4828,N_4785,N_4520);
xor U4829 (N_4829,N_4564,N_4605);
or U4830 (N_4830,N_4796,N_4739);
and U4831 (N_4831,N_4688,N_4570);
nand U4832 (N_4832,N_4744,N_4641);
nand U4833 (N_4833,N_4777,N_4527);
nor U4834 (N_4834,N_4710,N_4554);
and U4835 (N_4835,N_4515,N_4530);
or U4836 (N_4836,N_4627,N_4686);
nand U4837 (N_4837,N_4679,N_4504);
and U4838 (N_4838,N_4548,N_4611);
nor U4839 (N_4839,N_4664,N_4599);
nand U4840 (N_4840,N_4798,N_4591);
nor U4841 (N_4841,N_4676,N_4542);
nor U4842 (N_4842,N_4707,N_4610);
nor U4843 (N_4843,N_4789,N_4742);
nor U4844 (N_4844,N_4563,N_4618);
or U4845 (N_4845,N_4717,N_4594);
xnor U4846 (N_4846,N_4606,N_4784);
and U4847 (N_4847,N_4626,N_4669);
or U4848 (N_4848,N_4667,N_4524);
or U4849 (N_4849,N_4757,N_4525);
nor U4850 (N_4850,N_4666,N_4769);
nand U4851 (N_4851,N_4791,N_4763);
xor U4852 (N_4852,N_4761,N_4683);
xor U4853 (N_4853,N_4608,N_4652);
and U4854 (N_4854,N_4569,N_4531);
xor U4855 (N_4855,N_4727,N_4692);
nand U4856 (N_4856,N_4571,N_4767);
or U4857 (N_4857,N_4507,N_4519);
or U4858 (N_4858,N_4714,N_4685);
or U4859 (N_4859,N_4510,N_4556);
and U4860 (N_4860,N_4628,N_4511);
xor U4861 (N_4861,N_4722,N_4500);
and U4862 (N_4862,N_4620,N_4545);
xnor U4863 (N_4863,N_4706,N_4636);
and U4864 (N_4864,N_4642,N_4546);
and U4865 (N_4865,N_4773,N_4694);
and U4866 (N_4866,N_4740,N_4622);
nor U4867 (N_4867,N_4660,N_4517);
and U4868 (N_4868,N_4675,N_4601);
xor U4869 (N_4869,N_4644,N_4684);
xnor U4870 (N_4870,N_4691,N_4700);
xnor U4871 (N_4871,N_4573,N_4663);
and U4872 (N_4872,N_4568,N_4711);
xor U4873 (N_4873,N_4790,N_4795);
nor U4874 (N_4874,N_4759,N_4687);
or U4875 (N_4875,N_4577,N_4731);
nand U4876 (N_4876,N_4779,N_4762);
and U4877 (N_4877,N_4629,N_4640);
nand U4878 (N_4878,N_4590,N_4578);
nand U4879 (N_4879,N_4593,N_4508);
xor U4880 (N_4880,N_4543,N_4512);
xnor U4881 (N_4881,N_4615,N_4723);
and U4882 (N_4882,N_4536,N_4792);
nor U4883 (N_4883,N_4658,N_4575);
xor U4884 (N_4884,N_4713,N_4637);
nor U4885 (N_4885,N_4502,N_4657);
nand U4886 (N_4886,N_4634,N_4765);
nand U4887 (N_4887,N_4528,N_4567);
nand U4888 (N_4888,N_4673,N_4597);
and U4889 (N_4889,N_4728,N_4797);
or U4890 (N_4890,N_4774,N_4513);
nor U4891 (N_4891,N_4756,N_4668);
or U4892 (N_4892,N_4748,N_4539);
or U4893 (N_4893,N_4607,N_4521);
xor U4894 (N_4894,N_4621,N_4743);
nand U4895 (N_4895,N_4755,N_4689);
nor U4896 (N_4896,N_4592,N_4659);
xor U4897 (N_4897,N_4544,N_4661);
xor U4898 (N_4898,N_4738,N_4589);
xor U4899 (N_4899,N_4523,N_4586);
xnor U4900 (N_4900,N_4535,N_4550);
nand U4901 (N_4901,N_4633,N_4712);
nand U4902 (N_4902,N_4703,N_4775);
and U4903 (N_4903,N_4505,N_4751);
or U4904 (N_4904,N_4677,N_4750);
or U4905 (N_4905,N_4624,N_4553);
xnor U4906 (N_4906,N_4561,N_4643);
or U4907 (N_4907,N_4518,N_4726);
or U4908 (N_4908,N_4752,N_4708);
nand U4909 (N_4909,N_4749,N_4787);
nand U4910 (N_4910,N_4623,N_4580);
xor U4911 (N_4911,N_4503,N_4565);
nor U4912 (N_4912,N_4632,N_4772);
or U4913 (N_4913,N_4613,N_4609);
nand U4914 (N_4914,N_4646,N_4732);
or U4915 (N_4915,N_4595,N_4648);
nor U4916 (N_4916,N_4562,N_4733);
nor U4917 (N_4917,N_4576,N_4695);
or U4918 (N_4918,N_4579,N_4651);
nand U4919 (N_4919,N_4537,N_4690);
xor U4920 (N_4920,N_4506,N_4720);
xor U4921 (N_4921,N_4581,N_4549);
or U4922 (N_4922,N_4760,N_4682);
or U4923 (N_4923,N_4665,N_4509);
xnor U4924 (N_4924,N_4598,N_4619);
xnor U4925 (N_4925,N_4639,N_4721);
or U4926 (N_4926,N_4783,N_4719);
and U4927 (N_4927,N_4725,N_4754);
and U4928 (N_4928,N_4771,N_4547);
or U4929 (N_4929,N_4560,N_4558);
or U4930 (N_4930,N_4662,N_4788);
nor U4931 (N_4931,N_4603,N_4635);
xnor U4932 (N_4932,N_4734,N_4799);
nor U4933 (N_4933,N_4617,N_4572);
xnor U4934 (N_4934,N_4697,N_4631);
nor U4935 (N_4935,N_4559,N_4786);
or U4936 (N_4936,N_4693,N_4746);
and U4937 (N_4937,N_4778,N_4696);
xor U4938 (N_4938,N_4715,N_4768);
and U4939 (N_4939,N_4671,N_4540);
nand U4940 (N_4940,N_4645,N_4557);
xnor U4941 (N_4941,N_4650,N_4555);
xor U4942 (N_4942,N_4780,N_4614);
nand U4943 (N_4943,N_4538,N_4630);
or U4944 (N_4944,N_4730,N_4656);
or U4945 (N_4945,N_4745,N_4655);
nand U4946 (N_4946,N_4793,N_4532);
nand U4947 (N_4947,N_4552,N_4516);
nor U4948 (N_4948,N_4602,N_4702);
and U4949 (N_4949,N_4782,N_4649);
and U4950 (N_4950,N_4763,N_4792);
nor U4951 (N_4951,N_4799,N_4646);
and U4952 (N_4952,N_4780,N_4733);
xnor U4953 (N_4953,N_4524,N_4641);
nor U4954 (N_4954,N_4783,N_4757);
or U4955 (N_4955,N_4625,N_4789);
xnor U4956 (N_4956,N_4675,N_4797);
xor U4957 (N_4957,N_4600,N_4595);
xor U4958 (N_4958,N_4696,N_4782);
nand U4959 (N_4959,N_4672,N_4636);
nand U4960 (N_4960,N_4576,N_4509);
and U4961 (N_4961,N_4504,N_4528);
or U4962 (N_4962,N_4674,N_4759);
or U4963 (N_4963,N_4555,N_4541);
nor U4964 (N_4964,N_4748,N_4720);
and U4965 (N_4965,N_4526,N_4561);
nor U4966 (N_4966,N_4669,N_4585);
or U4967 (N_4967,N_4534,N_4679);
nand U4968 (N_4968,N_4536,N_4703);
or U4969 (N_4969,N_4568,N_4765);
or U4970 (N_4970,N_4552,N_4580);
nor U4971 (N_4971,N_4595,N_4517);
and U4972 (N_4972,N_4520,N_4715);
nand U4973 (N_4973,N_4790,N_4558);
nor U4974 (N_4974,N_4575,N_4536);
nor U4975 (N_4975,N_4511,N_4566);
xnor U4976 (N_4976,N_4526,N_4709);
and U4977 (N_4977,N_4736,N_4642);
or U4978 (N_4978,N_4688,N_4654);
or U4979 (N_4979,N_4760,N_4692);
or U4980 (N_4980,N_4699,N_4582);
and U4981 (N_4981,N_4783,N_4569);
nor U4982 (N_4982,N_4694,N_4593);
xor U4983 (N_4983,N_4780,N_4598);
and U4984 (N_4984,N_4744,N_4758);
nor U4985 (N_4985,N_4633,N_4683);
nand U4986 (N_4986,N_4646,N_4504);
and U4987 (N_4987,N_4506,N_4503);
xnor U4988 (N_4988,N_4502,N_4559);
or U4989 (N_4989,N_4579,N_4646);
and U4990 (N_4990,N_4649,N_4537);
xor U4991 (N_4991,N_4612,N_4691);
and U4992 (N_4992,N_4550,N_4770);
and U4993 (N_4993,N_4770,N_4757);
nand U4994 (N_4994,N_4553,N_4691);
xor U4995 (N_4995,N_4597,N_4546);
xor U4996 (N_4996,N_4650,N_4569);
xnor U4997 (N_4997,N_4794,N_4547);
and U4998 (N_4998,N_4692,N_4513);
nor U4999 (N_4999,N_4640,N_4627);
xnor U5000 (N_5000,N_4527,N_4531);
and U5001 (N_5001,N_4581,N_4659);
or U5002 (N_5002,N_4644,N_4591);
nand U5003 (N_5003,N_4602,N_4745);
nand U5004 (N_5004,N_4651,N_4739);
xor U5005 (N_5005,N_4770,N_4744);
nor U5006 (N_5006,N_4609,N_4724);
or U5007 (N_5007,N_4541,N_4535);
and U5008 (N_5008,N_4745,N_4730);
nand U5009 (N_5009,N_4662,N_4799);
xor U5010 (N_5010,N_4796,N_4733);
nand U5011 (N_5011,N_4527,N_4521);
xnor U5012 (N_5012,N_4614,N_4688);
xor U5013 (N_5013,N_4746,N_4657);
xnor U5014 (N_5014,N_4646,N_4699);
nor U5015 (N_5015,N_4567,N_4608);
and U5016 (N_5016,N_4591,N_4604);
or U5017 (N_5017,N_4586,N_4657);
and U5018 (N_5018,N_4764,N_4566);
and U5019 (N_5019,N_4639,N_4756);
xnor U5020 (N_5020,N_4606,N_4702);
or U5021 (N_5021,N_4665,N_4598);
and U5022 (N_5022,N_4783,N_4539);
nand U5023 (N_5023,N_4783,N_4721);
or U5024 (N_5024,N_4716,N_4692);
nor U5025 (N_5025,N_4648,N_4541);
or U5026 (N_5026,N_4759,N_4697);
nand U5027 (N_5027,N_4606,N_4756);
and U5028 (N_5028,N_4583,N_4710);
and U5029 (N_5029,N_4778,N_4722);
or U5030 (N_5030,N_4515,N_4729);
xor U5031 (N_5031,N_4641,N_4622);
xor U5032 (N_5032,N_4635,N_4639);
xor U5033 (N_5033,N_4688,N_4632);
and U5034 (N_5034,N_4674,N_4601);
nand U5035 (N_5035,N_4582,N_4619);
or U5036 (N_5036,N_4691,N_4501);
and U5037 (N_5037,N_4581,N_4568);
nand U5038 (N_5038,N_4686,N_4747);
xnor U5039 (N_5039,N_4609,N_4573);
xnor U5040 (N_5040,N_4713,N_4716);
xor U5041 (N_5041,N_4589,N_4575);
nor U5042 (N_5042,N_4690,N_4699);
xnor U5043 (N_5043,N_4717,N_4601);
xnor U5044 (N_5044,N_4652,N_4774);
or U5045 (N_5045,N_4591,N_4642);
and U5046 (N_5046,N_4755,N_4765);
nand U5047 (N_5047,N_4754,N_4721);
xor U5048 (N_5048,N_4719,N_4679);
nand U5049 (N_5049,N_4751,N_4546);
nor U5050 (N_5050,N_4606,N_4711);
nor U5051 (N_5051,N_4675,N_4791);
nand U5052 (N_5052,N_4754,N_4707);
nand U5053 (N_5053,N_4584,N_4716);
or U5054 (N_5054,N_4538,N_4729);
or U5055 (N_5055,N_4709,N_4767);
nor U5056 (N_5056,N_4744,N_4546);
nand U5057 (N_5057,N_4628,N_4673);
and U5058 (N_5058,N_4568,N_4750);
nand U5059 (N_5059,N_4770,N_4606);
nand U5060 (N_5060,N_4640,N_4718);
nand U5061 (N_5061,N_4503,N_4713);
and U5062 (N_5062,N_4578,N_4507);
and U5063 (N_5063,N_4616,N_4689);
xnor U5064 (N_5064,N_4770,N_4673);
and U5065 (N_5065,N_4772,N_4736);
xor U5066 (N_5066,N_4592,N_4773);
and U5067 (N_5067,N_4551,N_4599);
xor U5068 (N_5068,N_4595,N_4544);
and U5069 (N_5069,N_4536,N_4690);
nor U5070 (N_5070,N_4664,N_4638);
or U5071 (N_5071,N_4744,N_4717);
nand U5072 (N_5072,N_4686,N_4723);
nor U5073 (N_5073,N_4627,N_4737);
or U5074 (N_5074,N_4690,N_4663);
xor U5075 (N_5075,N_4761,N_4774);
and U5076 (N_5076,N_4525,N_4602);
or U5077 (N_5077,N_4625,N_4552);
xor U5078 (N_5078,N_4567,N_4578);
or U5079 (N_5079,N_4673,N_4737);
and U5080 (N_5080,N_4535,N_4698);
xor U5081 (N_5081,N_4649,N_4691);
nor U5082 (N_5082,N_4648,N_4515);
nand U5083 (N_5083,N_4730,N_4602);
xnor U5084 (N_5084,N_4733,N_4669);
and U5085 (N_5085,N_4593,N_4559);
nor U5086 (N_5086,N_4633,N_4605);
nor U5087 (N_5087,N_4540,N_4610);
nand U5088 (N_5088,N_4595,N_4584);
or U5089 (N_5089,N_4665,N_4771);
nand U5090 (N_5090,N_4505,N_4537);
xor U5091 (N_5091,N_4690,N_4521);
or U5092 (N_5092,N_4667,N_4745);
xor U5093 (N_5093,N_4557,N_4770);
xnor U5094 (N_5094,N_4699,N_4796);
xor U5095 (N_5095,N_4629,N_4665);
nor U5096 (N_5096,N_4676,N_4532);
or U5097 (N_5097,N_4689,N_4687);
xor U5098 (N_5098,N_4675,N_4689);
and U5099 (N_5099,N_4535,N_4778);
nor U5100 (N_5100,N_4925,N_4888);
xor U5101 (N_5101,N_5021,N_5091);
or U5102 (N_5102,N_4970,N_5073);
or U5103 (N_5103,N_4989,N_5087);
or U5104 (N_5104,N_4893,N_5004);
nor U5105 (N_5105,N_5020,N_5025);
nand U5106 (N_5106,N_5012,N_4811);
nand U5107 (N_5107,N_4987,N_5046);
nand U5108 (N_5108,N_5051,N_4871);
and U5109 (N_5109,N_4820,N_4861);
and U5110 (N_5110,N_4990,N_4876);
xnor U5111 (N_5111,N_5085,N_4931);
or U5112 (N_5112,N_4836,N_4992);
nor U5113 (N_5113,N_4806,N_5069);
nor U5114 (N_5114,N_4900,N_4884);
nor U5115 (N_5115,N_5003,N_4919);
nor U5116 (N_5116,N_5057,N_4897);
and U5117 (N_5117,N_4907,N_5006);
or U5118 (N_5118,N_4964,N_5045);
nor U5119 (N_5119,N_5029,N_4842);
xor U5120 (N_5120,N_4974,N_4874);
and U5121 (N_5121,N_4819,N_5080);
xor U5122 (N_5122,N_4872,N_5064);
nand U5123 (N_5123,N_4891,N_4980);
nand U5124 (N_5124,N_4911,N_4856);
or U5125 (N_5125,N_4933,N_5017);
and U5126 (N_5126,N_5093,N_4805);
nor U5127 (N_5127,N_4971,N_5037);
or U5128 (N_5128,N_5050,N_5082);
or U5129 (N_5129,N_4955,N_5042);
xor U5130 (N_5130,N_4831,N_4914);
or U5131 (N_5131,N_4939,N_4847);
nor U5132 (N_5132,N_5084,N_4943);
nand U5133 (N_5133,N_4951,N_4921);
or U5134 (N_5134,N_4881,N_4870);
nor U5135 (N_5135,N_5090,N_4928);
nor U5136 (N_5136,N_4882,N_4862);
and U5137 (N_5137,N_4969,N_4944);
xnor U5138 (N_5138,N_5086,N_4863);
xor U5139 (N_5139,N_4972,N_5065);
or U5140 (N_5140,N_5001,N_4804);
nor U5141 (N_5141,N_4910,N_4937);
or U5142 (N_5142,N_4952,N_5077);
xnor U5143 (N_5143,N_4993,N_5039);
nand U5144 (N_5144,N_4945,N_4983);
and U5145 (N_5145,N_5066,N_5008);
and U5146 (N_5146,N_5000,N_4817);
and U5147 (N_5147,N_4896,N_4843);
nor U5148 (N_5148,N_4926,N_5009);
xor U5149 (N_5149,N_4956,N_5019);
nand U5150 (N_5150,N_4946,N_4832);
nand U5151 (N_5151,N_4998,N_5055);
nor U5152 (N_5152,N_4865,N_4875);
nor U5153 (N_5153,N_4966,N_5088);
nor U5154 (N_5154,N_5010,N_4903);
nand U5155 (N_5155,N_5092,N_4853);
xnor U5156 (N_5156,N_5034,N_5096);
nor U5157 (N_5157,N_5030,N_5061);
and U5158 (N_5158,N_5005,N_4857);
nor U5159 (N_5159,N_5033,N_4938);
nand U5160 (N_5160,N_4880,N_4941);
and U5161 (N_5161,N_4878,N_4991);
xor U5162 (N_5162,N_4835,N_5072);
or U5163 (N_5163,N_4984,N_5074);
xor U5164 (N_5164,N_4909,N_4818);
nand U5165 (N_5165,N_4934,N_4995);
nand U5166 (N_5166,N_4829,N_4917);
nand U5167 (N_5167,N_4967,N_4958);
nand U5168 (N_5168,N_5081,N_4961);
or U5169 (N_5169,N_4962,N_4902);
and U5170 (N_5170,N_5068,N_4822);
xnor U5171 (N_5171,N_4994,N_4830);
or U5172 (N_5172,N_4976,N_4930);
and U5173 (N_5173,N_5049,N_4916);
and U5174 (N_5174,N_5059,N_4950);
nor U5175 (N_5175,N_4924,N_4846);
xor U5176 (N_5176,N_4942,N_4965);
nand U5177 (N_5177,N_4812,N_5013);
nor U5178 (N_5178,N_4895,N_4954);
xnor U5179 (N_5179,N_5014,N_5028);
or U5180 (N_5180,N_4833,N_4840);
and U5181 (N_5181,N_5007,N_4801);
nand U5182 (N_5182,N_5026,N_4890);
xnor U5183 (N_5183,N_4908,N_4883);
and U5184 (N_5184,N_4906,N_4999);
nor U5185 (N_5185,N_4923,N_4850);
or U5186 (N_5186,N_5038,N_5094);
and U5187 (N_5187,N_4827,N_4986);
or U5188 (N_5188,N_4885,N_4927);
nor U5189 (N_5189,N_4826,N_5060);
xor U5190 (N_5190,N_5054,N_4898);
xnor U5191 (N_5191,N_4816,N_5040);
xnor U5192 (N_5192,N_4851,N_4813);
or U5193 (N_5193,N_5032,N_4867);
xor U5194 (N_5194,N_4929,N_5044);
nor U5195 (N_5195,N_4912,N_4968);
and U5196 (N_5196,N_4815,N_5099);
and U5197 (N_5197,N_4957,N_5071);
nand U5198 (N_5198,N_5070,N_4838);
nor U5199 (N_5199,N_5018,N_4837);
nor U5200 (N_5200,N_5075,N_4981);
nand U5201 (N_5201,N_5089,N_5048);
nor U5202 (N_5202,N_4940,N_4859);
and U5203 (N_5203,N_4932,N_5024);
nand U5204 (N_5204,N_4948,N_5063);
xor U5205 (N_5205,N_4899,N_4821);
xnor U5206 (N_5206,N_4834,N_4982);
or U5207 (N_5207,N_4809,N_4860);
nand U5208 (N_5208,N_4879,N_4901);
and U5209 (N_5209,N_4841,N_4947);
and U5210 (N_5210,N_5036,N_5076);
or U5211 (N_5211,N_4960,N_4807);
xor U5212 (N_5212,N_4997,N_5067);
and U5213 (N_5213,N_5027,N_4953);
or U5214 (N_5214,N_4844,N_4922);
nand U5215 (N_5215,N_5041,N_4828);
and U5216 (N_5216,N_4873,N_5022);
or U5217 (N_5217,N_5097,N_5098);
xnor U5218 (N_5218,N_5023,N_4866);
and U5219 (N_5219,N_5015,N_4949);
nand U5220 (N_5220,N_4877,N_4825);
or U5221 (N_5221,N_5031,N_4886);
xor U5222 (N_5222,N_5079,N_4975);
nor U5223 (N_5223,N_4869,N_4904);
and U5224 (N_5224,N_4996,N_4824);
or U5225 (N_5225,N_5083,N_5095);
and U5226 (N_5226,N_4855,N_5052);
nor U5227 (N_5227,N_4887,N_4978);
nor U5228 (N_5228,N_5035,N_5056);
xor U5229 (N_5229,N_5062,N_4913);
nor U5230 (N_5230,N_4814,N_5043);
and U5231 (N_5231,N_4894,N_4803);
and U5232 (N_5232,N_4889,N_4920);
nand U5233 (N_5233,N_4800,N_4848);
nand U5234 (N_5234,N_4808,N_4988);
xnor U5235 (N_5235,N_4823,N_4849);
or U5236 (N_5236,N_4915,N_4868);
or U5237 (N_5237,N_4918,N_5053);
nor U5238 (N_5238,N_5047,N_4979);
xnor U5239 (N_5239,N_4977,N_5016);
or U5240 (N_5240,N_4854,N_5011);
and U5241 (N_5241,N_5058,N_4959);
nand U5242 (N_5242,N_4839,N_4905);
or U5243 (N_5243,N_5078,N_4985);
nor U5244 (N_5244,N_4810,N_4936);
nand U5245 (N_5245,N_4864,N_4852);
xor U5246 (N_5246,N_4935,N_5002);
and U5247 (N_5247,N_4973,N_4845);
and U5248 (N_5248,N_4858,N_4802);
nand U5249 (N_5249,N_4963,N_4892);
xor U5250 (N_5250,N_4842,N_4806);
or U5251 (N_5251,N_4944,N_4980);
or U5252 (N_5252,N_4910,N_4875);
or U5253 (N_5253,N_4985,N_4917);
or U5254 (N_5254,N_4990,N_4819);
or U5255 (N_5255,N_4917,N_4892);
or U5256 (N_5256,N_5006,N_4920);
nor U5257 (N_5257,N_4916,N_4842);
xor U5258 (N_5258,N_4864,N_5038);
nor U5259 (N_5259,N_5025,N_4922);
or U5260 (N_5260,N_5059,N_5000);
and U5261 (N_5261,N_4802,N_4895);
xnor U5262 (N_5262,N_4944,N_4883);
nor U5263 (N_5263,N_4933,N_4851);
nand U5264 (N_5264,N_4805,N_4807);
xor U5265 (N_5265,N_4947,N_5018);
xor U5266 (N_5266,N_4975,N_4944);
or U5267 (N_5267,N_4820,N_5094);
and U5268 (N_5268,N_5032,N_4837);
or U5269 (N_5269,N_4922,N_4928);
xor U5270 (N_5270,N_5016,N_4833);
xor U5271 (N_5271,N_5088,N_5064);
xor U5272 (N_5272,N_4992,N_4923);
and U5273 (N_5273,N_4908,N_5037);
and U5274 (N_5274,N_4813,N_5033);
and U5275 (N_5275,N_4998,N_4910);
or U5276 (N_5276,N_4899,N_4826);
xnor U5277 (N_5277,N_4976,N_5093);
nor U5278 (N_5278,N_4888,N_4801);
nand U5279 (N_5279,N_4811,N_4884);
or U5280 (N_5280,N_5055,N_4984);
xor U5281 (N_5281,N_4898,N_5090);
nand U5282 (N_5282,N_4841,N_4978);
xor U5283 (N_5283,N_4827,N_4950);
nand U5284 (N_5284,N_4908,N_5010);
xnor U5285 (N_5285,N_4811,N_5025);
nand U5286 (N_5286,N_5025,N_4954);
xor U5287 (N_5287,N_5088,N_5070);
nand U5288 (N_5288,N_5093,N_4992);
xnor U5289 (N_5289,N_4991,N_5037);
nand U5290 (N_5290,N_4981,N_4834);
nor U5291 (N_5291,N_5025,N_4982);
nand U5292 (N_5292,N_5052,N_4903);
and U5293 (N_5293,N_4893,N_4983);
or U5294 (N_5294,N_4820,N_5015);
or U5295 (N_5295,N_5033,N_4839);
nand U5296 (N_5296,N_5080,N_4816);
nor U5297 (N_5297,N_4847,N_4881);
xnor U5298 (N_5298,N_4930,N_5011);
nand U5299 (N_5299,N_4841,N_5024);
nor U5300 (N_5300,N_5052,N_4856);
nand U5301 (N_5301,N_4957,N_5058);
nor U5302 (N_5302,N_5087,N_5030);
and U5303 (N_5303,N_4993,N_4897);
or U5304 (N_5304,N_5035,N_4816);
or U5305 (N_5305,N_4863,N_5040);
or U5306 (N_5306,N_4932,N_5061);
nand U5307 (N_5307,N_4893,N_4803);
or U5308 (N_5308,N_4825,N_4923);
xnor U5309 (N_5309,N_4922,N_4996);
or U5310 (N_5310,N_5037,N_4939);
xnor U5311 (N_5311,N_4997,N_5023);
xor U5312 (N_5312,N_5098,N_4935);
nor U5313 (N_5313,N_4907,N_4922);
or U5314 (N_5314,N_4846,N_4933);
xnor U5315 (N_5315,N_4912,N_4963);
or U5316 (N_5316,N_4917,N_4814);
nor U5317 (N_5317,N_4961,N_4977);
nand U5318 (N_5318,N_4957,N_4873);
nand U5319 (N_5319,N_4804,N_5070);
or U5320 (N_5320,N_4801,N_4894);
and U5321 (N_5321,N_5032,N_5029);
nand U5322 (N_5322,N_4929,N_4957);
and U5323 (N_5323,N_4903,N_5027);
or U5324 (N_5324,N_4952,N_4857);
nand U5325 (N_5325,N_5002,N_4988);
or U5326 (N_5326,N_4996,N_4911);
nor U5327 (N_5327,N_4820,N_4817);
and U5328 (N_5328,N_4805,N_4987);
or U5329 (N_5329,N_4876,N_4826);
and U5330 (N_5330,N_5077,N_4944);
and U5331 (N_5331,N_4816,N_4851);
xnor U5332 (N_5332,N_4883,N_4806);
and U5333 (N_5333,N_4861,N_4935);
xor U5334 (N_5334,N_4926,N_5043);
and U5335 (N_5335,N_5096,N_4869);
nand U5336 (N_5336,N_5026,N_4953);
nand U5337 (N_5337,N_4982,N_4849);
xor U5338 (N_5338,N_4907,N_4876);
and U5339 (N_5339,N_4853,N_4841);
nand U5340 (N_5340,N_5066,N_4821);
xnor U5341 (N_5341,N_4940,N_4880);
nor U5342 (N_5342,N_4985,N_4973);
or U5343 (N_5343,N_4857,N_4859);
nand U5344 (N_5344,N_4816,N_4951);
xor U5345 (N_5345,N_4852,N_4811);
xor U5346 (N_5346,N_5018,N_5067);
xnor U5347 (N_5347,N_5003,N_4903);
nand U5348 (N_5348,N_4992,N_4898);
or U5349 (N_5349,N_4814,N_5066);
nor U5350 (N_5350,N_5058,N_5062);
nor U5351 (N_5351,N_4995,N_5017);
xor U5352 (N_5352,N_4991,N_5052);
and U5353 (N_5353,N_5063,N_4959);
or U5354 (N_5354,N_4938,N_5049);
xnor U5355 (N_5355,N_4876,N_4997);
and U5356 (N_5356,N_5055,N_4811);
or U5357 (N_5357,N_5084,N_4928);
xnor U5358 (N_5358,N_5069,N_4965);
or U5359 (N_5359,N_4899,N_4948);
nand U5360 (N_5360,N_5086,N_4936);
or U5361 (N_5361,N_5060,N_4926);
nor U5362 (N_5362,N_4985,N_4878);
nor U5363 (N_5363,N_5035,N_5052);
and U5364 (N_5364,N_5049,N_4836);
nand U5365 (N_5365,N_4992,N_5012);
nand U5366 (N_5366,N_4854,N_5034);
nand U5367 (N_5367,N_4970,N_4860);
and U5368 (N_5368,N_4954,N_4990);
xor U5369 (N_5369,N_4888,N_4805);
xnor U5370 (N_5370,N_4923,N_4852);
and U5371 (N_5371,N_4978,N_5026);
nand U5372 (N_5372,N_4978,N_4848);
or U5373 (N_5373,N_4809,N_4907);
xor U5374 (N_5374,N_5003,N_4955);
nand U5375 (N_5375,N_4855,N_4921);
and U5376 (N_5376,N_4886,N_4864);
nor U5377 (N_5377,N_5007,N_4858);
nand U5378 (N_5378,N_4885,N_4854);
and U5379 (N_5379,N_4874,N_4966);
nor U5380 (N_5380,N_5084,N_5083);
nand U5381 (N_5381,N_4819,N_4832);
or U5382 (N_5382,N_5038,N_5010);
or U5383 (N_5383,N_5017,N_4821);
xnor U5384 (N_5384,N_5000,N_5091);
nor U5385 (N_5385,N_4861,N_4830);
nand U5386 (N_5386,N_4888,N_4945);
or U5387 (N_5387,N_4900,N_4967);
nor U5388 (N_5388,N_4807,N_4921);
nand U5389 (N_5389,N_4946,N_5036);
xnor U5390 (N_5390,N_5078,N_5063);
and U5391 (N_5391,N_5013,N_5055);
nor U5392 (N_5392,N_4976,N_5031);
or U5393 (N_5393,N_4968,N_5046);
xor U5394 (N_5394,N_4894,N_4946);
nand U5395 (N_5395,N_5006,N_4923);
xor U5396 (N_5396,N_4926,N_4881);
nand U5397 (N_5397,N_4882,N_4813);
and U5398 (N_5398,N_4899,N_5071);
nand U5399 (N_5399,N_5081,N_4846);
nor U5400 (N_5400,N_5170,N_5320);
nor U5401 (N_5401,N_5119,N_5325);
nand U5402 (N_5402,N_5342,N_5285);
and U5403 (N_5403,N_5117,N_5245);
nand U5404 (N_5404,N_5139,N_5177);
and U5405 (N_5405,N_5392,N_5159);
or U5406 (N_5406,N_5153,N_5179);
nand U5407 (N_5407,N_5306,N_5209);
nand U5408 (N_5408,N_5293,N_5313);
or U5409 (N_5409,N_5379,N_5275);
and U5410 (N_5410,N_5335,N_5116);
nor U5411 (N_5411,N_5184,N_5394);
nand U5412 (N_5412,N_5270,N_5241);
nand U5413 (N_5413,N_5276,N_5175);
and U5414 (N_5414,N_5222,N_5229);
xnor U5415 (N_5415,N_5109,N_5143);
and U5416 (N_5416,N_5375,N_5346);
xnor U5417 (N_5417,N_5149,N_5213);
xor U5418 (N_5418,N_5107,N_5301);
nand U5419 (N_5419,N_5307,N_5311);
and U5420 (N_5420,N_5126,N_5395);
xnor U5421 (N_5421,N_5130,N_5137);
or U5422 (N_5422,N_5193,N_5176);
nand U5423 (N_5423,N_5356,N_5147);
nor U5424 (N_5424,N_5278,N_5210);
xor U5425 (N_5425,N_5273,N_5372);
nand U5426 (N_5426,N_5236,N_5361);
nor U5427 (N_5427,N_5380,N_5322);
xor U5428 (N_5428,N_5316,N_5219);
and U5429 (N_5429,N_5277,N_5103);
and U5430 (N_5430,N_5262,N_5183);
or U5431 (N_5431,N_5259,N_5102);
nand U5432 (N_5432,N_5283,N_5230);
nand U5433 (N_5433,N_5370,N_5118);
xnor U5434 (N_5434,N_5255,N_5336);
nand U5435 (N_5435,N_5133,N_5339);
or U5436 (N_5436,N_5299,N_5221);
nand U5437 (N_5437,N_5148,N_5291);
and U5438 (N_5438,N_5247,N_5224);
and U5439 (N_5439,N_5207,N_5376);
or U5440 (N_5440,N_5189,N_5263);
nand U5441 (N_5441,N_5101,N_5233);
nand U5442 (N_5442,N_5127,N_5238);
xnor U5443 (N_5443,N_5249,N_5141);
nand U5444 (N_5444,N_5371,N_5243);
nor U5445 (N_5445,N_5142,N_5114);
and U5446 (N_5446,N_5389,N_5374);
nand U5447 (N_5447,N_5220,N_5384);
or U5448 (N_5448,N_5146,N_5298);
nand U5449 (N_5449,N_5378,N_5156);
xor U5450 (N_5450,N_5287,N_5180);
and U5451 (N_5451,N_5171,N_5225);
nand U5452 (N_5452,N_5309,N_5359);
xnor U5453 (N_5453,N_5267,N_5111);
and U5454 (N_5454,N_5125,N_5385);
xnor U5455 (N_5455,N_5327,N_5155);
xor U5456 (N_5456,N_5203,N_5129);
nor U5457 (N_5457,N_5257,N_5305);
and U5458 (N_5458,N_5252,N_5152);
xor U5459 (N_5459,N_5333,N_5202);
nor U5460 (N_5460,N_5244,N_5188);
xor U5461 (N_5461,N_5261,N_5223);
or U5462 (N_5462,N_5338,N_5279);
and U5463 (N_5463,N_5154,N_5345);
nand U5464 (N_5464,N_5344,N_5218);
nor U5465 (N_5465,N_5382,N_5377);
nand U5466 (N_5466,N_5196,N_5271);
and U5467 (N_5467,N_5163,N_5348);
xor U5468 (N_5468,N_5303,N_5295);
xor U5469 (N_5469,N_5260,N_5134);
xor U5470 (N_5470,N_5312,N_5368);
nand U5471 (N_5471,N_5274,N_5248);
nor U5472 (N_5472,N_5166,N_5272);
or U5473 (N_5473,N_5214,N_5365);
nand U5474 (N_5474,N_5239,N_5264);
nand U5475 (N_5475,N_5317,N_5397);
xnor U5476 (N_5476,N_5104,N_5300);
and U5477 (N_5477,N_5200,N_5122);
nor U5478 (N_5478,N_5296,N_5396);
xnor U5479 (N_5479,N_5286,N_5237);
xor U5480 (N_5480,N_5319,N_5165);
xor U5481 (N_5481,N_5268,N_5204);
and U5482 (N_5482,N_5289,N_5235);
xor U5483 (N_5483,N_5355,N_5280);
xor U5484 (N_5484,N_5304,N_5297);
and U5485 (N_5485,N_5324,N_5367);
nand U5486 (N_5486,N_5173,N_5205);
and U5487 (N_5487,N_5121,N_5199);
nand U5488 (N_5488,N_5231,N_5323);
nand U5489 (N_5489,N_5105,N_5331);
nor U5490 (N_5490,N_5390,N_5211);
xnor U5491 (N_5491,N_5308,N_5251);
and U5492 (N_5492,N_5253,N_5284);
nand U5493 (N_5493,N_5250,N_5329);
nor U5494 (N_5494,N_5354,N_5341);
xnor U5495 (N_5495,N_5106,N_5131);
or U5496 (N_5496,N_5201,N_5144);
and U5497 (N_5497,N_5358,N_5321);
xnor U5498 (N_5498,N_5123,N_5388);
nand U5499 (N_5499,N_5349,N_5217);
or U5500 (N_5500,N_5351,N_5310);
or U5501 (N_5501,N_5330,N_5162);
nand U5502 (N_5502,N_5288,N_5269);
or U5503 (N_5503,N_5100,N_5246);
xnor U5504 (N_5504,N_5172,N_5332);
nand U5505 (N_5505,N_5178,N_5360);
xnor U5506 (N_5506,N_5386,N_5181);
or U5507 (N_5507,N_5208,N_5254);
and U5508 (N_5508,N_5357,N_5206);
and U5509 (N_5509,N_5383,N_5337);
or U5510 (N_5510,N_5212,N_5292);
nand U5511 (N_5511,N_5350,N_5167);
and U5512 (N_5512,N_5113,N_5326);
and U5513 (N_5513,N_5398,N_5168);
nand U5514 (N_5514,N_5314,N_5364);
and U5515 (N_5515,N_5216,N_5227);
and U5516 (N_5516,N_5315,N_5174);
nor U5517 (N_5517,N_5182,N_5138);
or U5518 (N_5518,N_5387,N_5110);
or U5519 (N_5519,N_5150,N_5343);
xor U5520 (N_5520,N_5158,N_5242);
or U5521 (N_5521,N_5145,N_5265);
or U5522 (N_5522,N_5192,N_5366);
or U5523 (N_5523,N_5169,N_5108);
nor U5524 (N_5524,N_5334,N_5187);
nor U5525 (N_5525,N_5234,N_5140);
nand U5526 (N_5526,N_5115,N_5399);
and U5527 (N_5527,N_5340,N_5124);
and U5528 (N_5528,N_5185,N_5160);
nand U5529 (N_5529,N_5256,N_5381);
nand U5530 (N_5530,N_5290,N_5195);
or U5531 (N_5531,N_5281,N_5228);
nor U5532 (N_5532,N_5161,N_5352);
nand U5533 (N_5533,N_5186,N_5240);
or U5534 (N_5534,N_5135,N_5151);
or U5535 (N_5535,N_5198,N_5369);
xor U5536 (N_5536,N_5258,N_5353);
or U5537 (N_5537,N_5373,N_5226);
nor U5538 (N_5538,N_5347,N_5136);
or U5539 (N_5539,N_5302,N_5318);
xor U5540 (N_5540,N_5120,N_5194);
nand U5541 (N_5541,N_5157,N_5266);
nand U5542 (N_5542,N_5164,N_5363);
xor U5543 (N_5543,N_5282,N_5362);
nor U5544 (N_5544,N_5393,N_5132);
nand U5545 (N_5545,N_5328,N_5215);
and U5546 (N_5546,N_5190,N_5128);
xor U5547 (N_5547,N_5232,N_5391);
nand U5548 (N_5548,N_5197,N_5294);
or U5549 (N_5549,N_5112,N_5191);
and U5550 (N_5550,N_5335,N_5361);
nor U5551 (N_5551,N_5337,N_5150);
xnor U5552 (N_5552,N_5309,N_5374);
xor U5553 (N_5553,N_5279,N_5264);
or U5554 (N_5554,N_5347,N_5276);
or U5555 (N_5555,N_5240,N_5336);
nand U5556 (N_5556,N_5389,N_5120);
xor U5557 (N_5557,N_5110,N_5312);
or U5558 (N_5558,N_5220,N_5164);
nor U5559 (N_5559,N_5373,N_5306);
and U5560 (N_5560,N_5155,N_5193);
xor U5561 (N_5561,N_5311,N_5182);
or U5562 (N_5562,N_5155,N_5317);
nor U5563 (N_5563,N_5137,N_5215);
nand U5564 (N_5564,N_5246,N_5183);
or U5565 (N_5565,N_5312,N_5372);
or U5566 (N_5566,N_5354,N_5277);
nor U5567 (N_5567,N_5146,N_5370);
nor U5568 (N_5568,N_5252,N_5134);
xnor U5569 (N_5569,N_5134,N_5121);
or U5570 (N_5570,N_5292,N_5119);
xnor U5571 (N_5571,N_5313,N_5175);
or U5572 (N_5572,N_5382,N_5191);
nor U5573 (N_5573,N_5393,N_5117);
nand U5574 (N_5574,N_5191,N_5127);
and U5575 (N_5575,N_5351,N_5256);
xnor U5576 (N_5576,N_5275,N_5160);
and U5577 (N_5577,N_5278,N_5231);
nand U5578 (N_5578,N_5364,N_5245);
xor U5579 (N_5579,N_5143,N_5389);
nand U5580 (N_5580,N_5371,N_5125);
or U5581 (N_5581,N_5356,N_5213);
and U5582 (N_5582,N_5116,N_5264);
nand U5583 (N_5583,N_5188,N_5382);
nor U5584 (N_5584,N_5355,N_5259);
and U5585 (N_5585,N_5179,N_5178);
or U5586 (N_5586,N_5160,N_5101);
nor U5587 (N_5587,N_5354,N_5263);
nand U5588 (N_5588,N_5209,N_5268);
nor U5589 (N_5589,N_5213,N_5340);
xor U5590 (N_5590,N_5107,N_5275);
xor U5591 (N_5591,N_5255,N_5145);
or U5592 (N_5592,N_5364,N_5248);
or U5593 (N_5593,N_5385,N_5174);
nor U5594 (N_5594,N_5241,N_5141);
xor U5595 (N_5595,N_5339,N_5283);
and U5596 (N_5596,N_5268,N_5301);
nor U5597 (N_5597,N_5126,N_5139);
or U5598 (N_5598,N_5244,N_5146);
or U5599 (N_5599,N_5240,N_5354);
and U5600 (N_5600,N_5317,N_5273);
nand U5601 (N_5601,N_5132,N_5134);
nand U5602 (N_5602,N_5374,N_5302);
nand U5603 (N_5603,N_5293,N_5182);
nor U5604 (N_5604,N_5198,N_5167);
nand U5605 (N_5605,N_5149,N_5320);
nand U5606 (N_5606,N_5392,N_5353);
xor U5607 (N_5607,N_5169,N_5172);
nor U5608 (N_5608,N_5350,N_5144);
xor U5609 (N_5609,N_5104,N_5136);
xor U5610 (N_5610,N_5328,N_5137);
or U5611 (N_5611,N_5135,N_5105);
nand U5612 (N_5612,N_5141,N_5110);
and U5613 (N_5613,N_5373,N_5168);
and U5614 (N_5614,N_5196,N_5384);
or U5615 (N_5615,N_5257,N_5341);
xnor U5616 (N_5616,N_5368,N_5128);
nand U5617 (N_5617,N_5177,N_5344);
nand U5618 (N_5618,N_5235,N_5241);
or U5619 (N_5619,N_5338,N_5349);
and U5620 (N_5620,N_5171,N_5367);
and U5621 (N_5621,N_5331,N_5221);
nor U5622 (N_5622,N_5336,N_5261);
or U5623 (N_5623,N_5102,N_5170);
nor U5624 (N_5624,N_5208,N_5174);
or U5625 (N_5625,N_5275,N_5343);
nand U5626 (N_5626,N_5242,N_5314);
and U5627 (N_5627,N_5207,N_5187);
or U5628 (N_5628,N_5357,N_5280);
or U5629 (N_5629,N_5215,N_5155);
nand U5630 (N_5630,N_5160,N_5289);
nand U5631 (N_5631,N_5335,N_5113);
nor U5632 (N_5632,N_5103,N_5355);
or U5633 (N_5633,N_5302,N_5213);
or U5634 (N_5634,N_5223,N_5121);
xor U5635 (N_5635,N_5248,N_5154);
or U5636 (N_5636,N_5392,N_5194);
xor U5637 (N_5637,N_5377,N_5165);
nand U5638 (N_5638,N_5285,N_5273);
nor U5639 (N_5639,N_5368,N_5294);
xnor U5640 (N_5640,N_5244,N_5301);
or U5641 (N_5641,N_5104,N_5176);
nor U5642 (N_5642,N_5344,N_5329);
xnor U5643 (N_5643,N_5164,N_5368);
xor U5644 (N_5644,N_5311,N_5180);
xnor U5645 (N_5645,N_5327,N_5200);
nor U5646 (N_5646,N_5213,N_5189);
nor U5647 (N_5647,N_5327,N_5262);
xnor U5648 (N_5648,N_5288,N_5370);
nand U5649 (N_5649,N_5226,N_5117);
or U5650 (N_5650,N_5117,N_5399);
xor U5651 (N_5651,N_5158,N_5368);
nand U5652 (N_5652,N_5275,N_5174);
and U5653 (N_5653,N_5189,N_5285);
and U5654 (N_5654,N_5375,N_5249);
xor U5655 (N_5655,N_5255,N_5228);
nand U5656 (N_5656,N_5362,N_5109);
nand U5657 (N_5657,N_5310,N_5335);
nand U5658 (N_5658,N_5254,N_5264);
nand U5659 (N_5659,N_5212,N_5329);
or U5660 (N_5660,N_5173,N_5272);
nor U5661 (N_5661,N_5281,N_5248);
xor U5662 (N_5662,N_5370,N_5267);
nand U5663 (N_5663,N_5186,N_5196);
and U5664 (N_5664,N_5104,N_5267);
or U5665 (N_5665,N_5309,N_5264);
or U5666 (N_5666,N_5376,N_5342);
and U5667 (N_5667,N_5303,N_5239);
and U5668 (N_5668,N_5115,N_5382);
and U5669 (N_5669,N_5316,N_5348);
or U5670 (N_5670,N_5272,N_5238);
xnor U5671 (N_5671,N_5154,N_5321);
nand U5672 (N_5672,N_5382,N_5334);
xnor U5673 (N_5673,N_5279,N_5360);
nor U5674 (N_5674,N_5345,N_5366);
nand U5675 (N_5675,N_5164,N_5179);
nor U5676 (N_5676,N_5306,N_5355);
and U5677 (N_5677,N_5285,N_5277);
nor U5678 (N_5678,N_5335,N_5333);
xor U5679 (N_5679,N_5329,N_5180);
nand U5680 (N_5680,N_5342,N_5310);
and U5681 (N_5681,N_5271,N_5109);
and U5682 (N_5682,N_5275,N_5391);
nand U5683 (N_5683,N_5143,N_5110);
nor U5684 (N_5684,N_5398,N_5275);
or U5685 (N_5685,N_5377,N_5257);
xor U5686 (N_5686,N_5137,N_5185);
nor U5687 (N_5687,N_5386,N_5339);
or U5688 (N_5688,N_5133,N_5349);
nor U5689 (N_5689,N_5219,N_5327);
and U5690 (N_5690,N_5170,N_5150);
nand U5691 (N_5691,N_5309,N_5112);
nand U5692 (N_5692,N_5135,N_5195);
and U5693 (N_5693,N_5119,N_5217);
xnor U5694 (N_5694,N_5210,N_5285);
nor U5695 (N_5695,N_5215,N_5191);
nand U5696 (N_5696,N_5128,N_5364);
xor U5697 (N_5697,N_5115,N_5204);
xnor U5698 (N_5698,N_5205,N_5162);
nand U5699 (N_5699,N_5184,N_5278);
nor U5700 (N_5700,N_5570,N_5495);
nand U5701 (N_5701,N_5473,N_5613);
and U5702 (N_5702,N_5439,N_5518);
nand U5703 (N_5703,N_5542,N_5586);
or U5704 (N_5704,N_5466,N_5440);
or U5705 (N_5705,N_5482,N_5535);
xor U5706 (N_5706,N_5643,N_5512);
xnor U5707 (N_5707,N_5515,N_5555);
and U5708 (N_5708,N_5417,N_5690);
or U5709 (N_5709,N_5657,N_5587);
and U5710 (N_5710,N_5626,N_5670);
nor U5711 (N_5711,N_5629,N_5623);
or U5712 (N_5712,N_5642,N_5599);
and U5713 (N_5713,N_5600,N_5451);
xor U5714 (N_5714,N_5589,N_5510);
xnor U5715 (N_5715,N_5562,N_5663);
nand U5716 (N_5716,N_5699,N_5454);
nor U5717 (N_5717,N_5694,N_5414);
and U5718 (N_5718,N_5572,N_5588);
xor U5719 (N_5719,N_5421,N_5524);
nor U5720 (N_5720,N_5689,N_5638);
and U5721 (N_5721,N_5499,N_5698);
xor U5722 (N_5722,N_5541,N_5616);
nand U5723 (N_5723,N_5617,N_5429);
or U5724 (N_5724,N_5428,N_5682);
or U5725 (N_5725,N_5457,N_5494);
xnor U5726 (N_5726,N_5654,N_5426);
and U5727 (N_5727,N_5450,N_5583);
and U5728 (N_5728,N_5575,N_5525);
nor U5729 (N_5729,N_5463,N_5416);
xor U5730 (N_5730,N_5564,N_5632);
nand U5731 (N_5731,N_5509,N_5635);
nor U5732 (N_5732,N_5423,N_5531);
nand U5733 (N_5733,N_5526,N_5513);
xnor U5734 (N_5734,N_5693,N_5485);
nor U5735 (N_5735,N_5559,N_5688);
nor U5736 (N_5736,N_5449,N_5409);
and U5737 (N_5737,N_5540,N_5605);
nor U5738 (N_5738,N_5578,N_5500);
xnor U5739 (N_5739,N_5476,N_5558);
xor U5740 (N_5740,N_5641,N_5432);
and U5741 (N_5741,N_5528,N_5601);
nor U5742 (N_5742,N_5661,N_5461);
and U5743 (N_5743,N_5594,N_5472);
xor U5744 (N_5744,N_5592,N_5610);
or U5745 (N_5745,N_5553,N_5506);
xor U5746 (N_5746,N_5406,N_5458);
nand U5747 (N_5747,N_5614,N_5656);
xnor U5748 (N_5748,N_5478,N_5595);
nor U5749 (N_5749,N_5539,N_5627);
or U5750 (N_5750,N_5590,N_5520);
or U5751 (N_5751,N_5567,N_5673);
xor U5752 (N_5752,N_5508,N_5696);
and U5753 (N_5753,N_5465,N_5644);
nor U5754 (N_5754,N_5637,N_5573);
or U5755 (N_5755,N_5549,N_5444);
or U5756 (N_5756,N_5552,N_5684);
or U5757 (N_5757,N_5554,N_5672);
and U5758 (N_5758,N_5674,N_5408);
xor U5759 (N_5759,N_5681,N_5563);
nand U5760 (N_5760,N_5668,N_5568);
or U5761 (N_5761,N_5566,N_5471);
nand U5762 (N_5762,N_5521,N_5665);
nor U5763 (N_5763,N_5504,N_5447);
nand U5764 (N_5764,N_5479,N_5557);
and U5765 (N_5765,N_5452,N_5658);
xor U5766 (N_5766,N_5606,N_5652);
nand U5767 (N_5767,N_5550,N_5456);
or U5768 (N_5768,N_5662,N_5622);
xnor U5769 (N_5769,N_5490,N_5676);
or U5770 (N_5770,N_5496,N_5608);
nor U5771 (N_5771,N_5460,N_5430);
and U5772 (N_5772,N_5481,N_5529);
nand U5773 (N_5773,N_5593,N_5486);
xnor U5774 (N_5774,N_5691,N_5647);
or U5775 (N_5775,N_5653,N_5505);
nor U5776 (N_5776,N_5425,N_5602);
or U5777 (N_5777,N_5646,N_5420);
and U5778 (N_5778,N_5462,N_5574);
xor U5779 (N_5779,N_5427,N_5407);
nand U5780 (N_5780,N_5640,N_5669);
xnor U5781 (N_5781,N_5402,N_5679);
nor U5782 (N_5782,N_5493,N_5561);
nor U5783 (N_5783,N_5400,N_5683);
or U5784 (N_5784,N_5624,N_5446);
nor U5785 (N_5785,N_5651,N_5604);
xor U5786 (N_5786,N_5501,N_5618);
nand U5787 (N_5787,N_5659,N_5422);
xor U5788 (N_5788,N_5438,N_5403);
nor U5789 (N_5789,N_5413,N_5453);
and U5790 (N_5790,N_5569,N_5579);
nand U5791 (N_5791,N_5467,N_5609);
and U5792 (N_5792,N_5523,N_5437);
nand U5793 (N_5793,N_5410,N_5418);
nand U5794 (N_5794,N_5433,N_5639);
nand U5795 (N_5795,N_5544,N_5419);
nand U5796 (N_5796,N_5582,N_5516);
nor U5797 (N_5797,N_5630,N_5695);
or U5798 (N_5798,N_5680,N_5650);
nand U5799 (N_5799,N_5633,N_5671);
or U5800 (N_5800,N_5546,N_5470);
or U5801 (N_5801,N_5580,N_5631);
xnor U5802 (N_5802,N_5664,N_5443);
and U5803 (N_5803,N_5543,N_5483);
xnor U5804 (N_5804,N_5442,N_5538);
xor U5805 (N_5805,N_5660,N_5498);
or U5806 (N_5806,N_5678,N_5436);
xor U5807 (N_5807,N_5435,N_5455);
and U5808 (N_5808,N_5533,N_5556);
and U5809 (N_5809,N_5612,N_5655);
and U5810 (N_5810,N_5507,N_5615);
nor U5811 (N_5811,N_5489,N_5607);
nor U5812 (N_5812,N_5697,N_5459);
nand U5813 (N_5813,N_5666,N_5534);
nand U5814 (N_5814,N_5527,N_5448);
nor U5815 (N_5815,N_5537,N_5611);
and U5816 (N_5816,N_5474,N_5469);
and U5817 (N_5817,N_5645,N_5571);
or U5818 (N_5818,N_5487,N_5625);
nor U5819 (N_5819,N_5598,N_5675);
or U5820 (N_5820,N_5503,N_5511);
nand U5821 (N_5821,N_5581,N_5628);
and U5822 (N_5822,N_5441,N_5597);
or U5823 (N_5823,N_5404,N_5621);
xnor U5824 (N_5824,N_5415,N_5431);
nand U5825 (N_5825,N_5522,N_5685);
or U5826 (N_5826,N_5565,N_5484);
nand U5827 (N_5827,N_5551,N_5545);
or U5828 (N_5828,N_5667,N_5497);
nor U5829 (N_5829,N_5401,N_5584);
xor U5830 (N_5830,N_5686,N_5577);
and U5831 (N_5831,N_5517,N_5585);
or U5832 (N_5832,N_5591,N_5620);
nand U5833 (N_5833,N_5634,N_5412);
or U5834 (N_5834,N_5424,N_5492);
xnor U5835 (N_5835,N_5603,N_5536);
nor U5836 (N_5836,N_5576,N_5619);
nand U5837 (N_5837,N_5491,N_5445);
nor U5838 (N_5838,N_5464,N_5405);
and U5839 (N_5839,N_5648,N_5468);
nor U5840 (N_5840,N_5692,N_5547);
or U5841 (N_5841,N_5596,N_5502);
xor U5842 (N_5842,N_5548,N_5636);
or U5843 (N_5843,N_5532,N_5411);
nor U5844 (N_5844,N_5480,N_5560);
and U5845 (N_5845,N_5488,N_5434);
or U5846 (N_5846,N_5519,N_5687);
nand U5847 (N_5847,N_5649,N_5477);
nor U5848 (N_5848,N_5475,N_5514);
and U5849 (N_5849,N_5677,N_5530);
or U5850 (N_5850,N_5476,N_5590);
xor U5851 (N_5851,N_5442,N_5458);
nor U5852 (N_5852,N_5683,N_5483);
or U5853 (N_5853,N_5508,N_5530);
xor U5854 (N_5854,N_5693,N_5514);
and U5855 (N_5855,N_5540,N_5476);
nor U5856 (N_5856,N_5633,N_5446);
and U5857 (N_5857,N_5568,N_5654);
nand U5858 (N_5858,N_5682,N_5479);
and U5859 (N_5859,N_5567,N_5443);
or U5860 (N_5860,N_5677,N_5639);
nor U5861 (N_5861,N_5634,N_5522);
xnor U5862 (N_5862,N_5405,N_5694);
and U5863 (N_5863,N_5474,N_5509);
nand U5864 (N_5864,N_5481,N_5605);
xnor U5865 (N_5865,N_5557,N_5401);
nor U5866 (N_5866,N_5587,N_5422);
nor U5867 (N_5867,N_5430,N_5409);
or U5868 (N_5868,N_5676,N_5563);
or U5869 (N_5869,N_5571,N_5638);
nor U5870 (N_5870,N_5471,N_5550);
or U5871 (N_5871,N_5502,N_5693);
xnor U5872 (N_5872,N_5602,N_5414);
and U5873 (N_5873,N_5453,N_5597);
nand U5874 (N_5874,N_5630,N_5408);
nor U5875 (N_5875,N_5548,N_5673);
nor U5876 (N_5876,N_5425,N_5634);
xor U5877 (N_5877,N_5683,N_5604);
or U5878 (N_5878,N_5564,N_5543);
and U5879 (N_5879,N_5543,N_5684);
or U5880 (N_5880,N_5416,N_5468);
or U5881 (N_5881,N_5481,N_5488);
nor U5882 (N_5882,N_5578,N_5595);
and U5883 (N_5883,N_5446,N_5447);
nand U5884 (N_5884,N_5550,N_5448);
or U5885 (N_5885,N_5699,N_5599);
nor U5886 (N_5886,N_5532,N_5630);
xor U5887 (N_5887,N_5445,N_5667);
xor U5888 (N_5888,N_5603,N_5471);
and U5889 (N_5889,N_5668,N_5651);
or U5890 (N_5890,N_5639,N_5598);
nand U5891 (N_5891,N_5635,N_5474);
or U5892 (N_5892,N_5414,N_5579);
and U5893 (N_5893,N_5483,N_5490);
or U5894 (N_5894,N_5639,N_5685);
xor U5895 (N_5895,N_5569,N_5507);
nand U5896 (N_5896,N_5576,N_5502);
or U5897 (N_5897,N_5406,N_5621);
and U5898 (N_5898,N_5598,N_5684);
nand U5899 (N_5899,N_5589,N_5695);
and U5900 (N_5900,N_5602,N_5586);
nand U5901 (N_5901,N_5632,N_5407);
nor U5902 (N_5902,N_5538,N_5409);
xnor U5903 (N_5903,N_5506,N_5632);
and U5904 (N_5904,N_5419,N_5690);
or U5905 (N_5905,N_5409,N_5506);
or U5906 (N_5906,N_5451,N_5590);
xnor U5907 (N_5907,N_5671,N_5523);
nor U5908 (N_5908,N_5582,N_5635);
or U5909 (N_5909,N_5567,N_5551);
nor U5910 (N_5910,N_5603,N_5604);
or U5911 (N_5911,N_5416,N_5699);
nor U5912 (N_5912,N_5637,N_5667);
and U5913 (N_5913,N_5571,N_5642);
or U5914 (N_5914,N_5508,N_5453);
xnor U5915 (N_5915,N_5512,N_5688);
and U5916 (N_5916,N_5501,N_5475);
nand U5917 (N_5917,N_5672,N_5564);
and U5918 (N_5918,N_5667,N_5633);
nand U5919 (N_5919,N_5431,N_5494);
nor U5920 (N_5920,N_5627,N_5451);
nor U5921 (N_5921,N_5572,N_5626);
xor U5922 (N_5922,N_5500,N_5440);
nor U5923 (N_5923,N_5446,N_5564);
nand U5924 (N_5924,N_5455,N_5443);
and U5925 (N_5925,N_5415,N_5557);
xor U5926 (N_5926,N_5650,N_5560);
or U5927 (N_5927,N_5650,N_5555);
xor U5928 (N_5928,N_5642,N_5625);
xor U5929 (N_5929,N_5469,N_5640);
xnor U5930 (N_5930,N_5649,N_5431);
nor U5931 (N_5931,N_5416,N_5679);
xnor U5932 (N_5932,N_5546,N_5438);
nand U5933 (N_5933,N_5620,N_5542);
nand U5934 (N_5934,N_5525,N_5670);
or U5935 (N_5935,N_5621,N_5477);
and U5936 (N_5936,N_5693,N_5447);
or U5937 (N_5937,N_5474,N_5592);
and U5938 (N_5938,N_5440,N_5667);
xnor U5939 (N_5939,N_5417,N_5534);
or U5940 (N_5940,N_5599,N_5664);
or U5941 (N_5941,N_5536,N_5638);
or U5942 (N_5942,N_5628,N_5471);
or U5943 (N_5943,N_5524,N_5616);
nor U5944 (N_5944,N_5514,N_5468);
nand U5945 (N_5945,N_5580,N_5570);
or U5946 (N_5946,N_5510,N_5512);
or U5947 (N_5947,N_5624,N_5657);
or U5948 (N_5948,N_5697,N_5584);
or U5949 (N_5949,N_5425,N_5473);
nor U5950 (N_5950,N_5523,N_5521);
nand U5951 (N_5951,N_5470,N_5612);
xnor U5952 (N_5952,N_5414,N_5652);
nand U5953 (N_5953,N_5436,N_5635);
or U5954 (N_5954,N_5588,N_5699);
and U5955 (N_5955,N_5557,N_5674);
nor U5956 (N_5956,N_5441,N_5486);
nand U5957 (N_5957,N_5411,N_5512);
and U5958 (N_5958,N_5639,N_5422);
xnor U5959 (N_5959,N_5445,N_5414);
nand U5960 (N_5960,N_5407,N_5475);
nand U5961 (N_5961,N_5496,N_5430);
nand U5962 (N_5962,N_5526,N_5586);
nor U5963 (N_5963,N_5557,N_5678);
or U5964 (N_5964,N_5584,N_5683);
nor U5965 (N_5965,N_5470,N_5692);
and U5966 (N_5966,N_5657,N_5553);
and U5967 (N_5967,N_5556,N_5479);
and U5968 (N_5968,N_5487,N_5427);
xor U5969 (N_5969,N_5560,N_5607);
nand U5970 (N_5970,N_5421,N_5519);
xor U5971 (N_5971,N_5649,N_5468);
nand U5972 (N_5972,N_5574,N_5549);
nand U5973 (N_5973,N_5481,N_5677);
nor U5974 (N_5974,N_5409,N_5672);
and U5975 (N_5975,N_5516,N_5465);
or U5976 (N_5976,N_5572,N_5633);
nor U5977 (N_5977,N_5671,N_5477);
and U5978 (N_5978,N_5449,N_5470);
xnor U5979 (N_5979,N_5555,N_5662);
xor U5980 (N_5980,N_5524,N_5534);
nand U5981 (N_5981,N_5452,N_5556);
xor U5982 (N_5982,N_5522,N_5624);
or U5983 (N_5983,N_5428,N_5559);
nand U5984 (N_5984,N_5693,N_5541);
nor U5985 (N_5985,N_5567,N_5453);
nor U5986 (N_5986,N_5622,N_5551);
nand U5987 (N_5987,N_5438,N_5556);
nor U5988 (N_5988,N_5678,N_5579);
nand U5989 (N_5989,N_5428,N_5582);
and U5990 (N_5990,N_5400,N_5500);
xnor U5991 (N_5991,N_5455,N_5487);
or U5992 (N_5992,N_5588,N_5673);
nor U5993 (N_5993,N_5450,N_5499);
or U5994 (N_5994,N_5587,N_5430);
xor U5995 (N_5995,N_5567,N_5535);
nor U5996 (N_5996,N_5621,N_5521);
nand U5997 (N_5997,N_5465,N_5579);
or U5998 (N_5998,N_5635,N_5646);
nand U5999 (N_5999,N_5479,N_5404);
and U6000 (N_6000,N_5707,N_5899);
and U6001 (N_6001,N_5997,N_5882);
nor U6002 (N_6002,N_5913,N_5918);
or U6003 (N_6003,N_5809,N_5821);
nor U6004 (N_6004,N_5836,N_5860);
nor U6005 (N_6005,N_5756,N_5924);
nor U6006 (N_6006,N_5921,N_5830);
xnor U6007 (N_6007,N_5896,N_5722);
or U6008 (N_6008,N_5846,N_5715);
nor U6009 (N_6009,N_5868,N_5930);
xor U6010 (N_6010,N_5964,N_5724);
xor U6011 (N_6011,N_5703,N_5827);
or U6012 (N_6012,N_5876,N_5853);
nand U6013 (N_6013,N_5966,N_5768);
nand U6014 (N_6014,N_5718,N_5959);
xnor U6015 (N_6015,N_5794,N_5817);
xor U6016 (N_6016,N_5828,N_5877);
nand U6017 (N_6017,N_5739,N_5976);
nor U6018 (N_6018,N_5986,N_5951);
nand U6019 (N_6019,N_5990,N_5791);
and U6020 (N_6020,N_5814,N_5970);
or U6021 (N_6021,N_5942,N_5806);
or U6022 (N_6022,N_5772,N_5844);
and U6023 (N_6023,N_5710,N_5985);
nor U6024 (N_6024,N_5738,N_5788);
nor U6025 (N_6025,N_5734,N_5841);
xnor U6026 (N_6026,N_5885,N_5781);
xor U6027 (N_6027,N_5701,N_5889);
nor U6028 (N_6028,N_5870,N_5880);
xnor U6029 (N_6029,N_5748,N_5826);
xor U6030 (N_6030,N_5850,N_5898);
xnor U6031 (N_6031,N_5866,N_5953);
nand U6032 (N_6032,N_5937,N_5927);
and U6033 (N_6033,N_5727,N_5716);
nor U6034 (N_6034,N_5883,N_5736);
xnor U6035 (N_6035,N_5775,N_5910);
xor U6036 (N_6036,N_5878,N_5996);
and U6037 (N_6037,N_5792,N_5746);
and U6038 (N_6038,N_5713,N_5934);
xnor U6039 (N_6039,N_5816,N_5785);
nor U6040 (N_6040,N_5919,N_5749);
nor U6041 (N_6041,N_5799,N_5787);
xor U6042 (N_6042,N_5995,N_5929);
xnor U6043 (N_6043,N_5780,N_5893);
xor U6044 (N_6044,N_5725,N_5755);
nand U6045 (N_6045,N_5873,N_5831);
xor U6046 (N_6046,N_5980,N_5906);
nor U6047 (N_6047,N_5797,N_5782);
nor U6048 (N_6048,N_5954,N_5917);
nor U6049 (N_6049,N_5867,N_5773);
nor U6050 (N_6050,N_5938,N_5948);
or U6051 (N_6051,N_5705,N_5881);
and U6052 (N_6052,N_5798,N_5887);
or U6053 (N_6053,N_5952,N_5769);
and U6054 (N_6054,N_5891,N_5793);
xor U6055 (N_6055,N_5994,N_5956);
and U6056 (N_6056,N_5884,N_5900);
xor U6057 (N_6057,N_5947,N_5897);
xor U6058 (N_6058,N_5911,N_5901);
nand U6059 (N_6059,N_5928,N_5865);
xor U6060 (N_6060,N_5983,N_5998);
nand U6061 (N_6061,N_5702,N_5704);
nand U6062 (N_6062,N_5759,N_5904);
xor U6063 (N_6063,N_5751,N_5712);
and U6064 (N_6064,N_5862,N_5820);
nor U6065 (N_6065,N_5895,N_5700);
nand U6066 (N_6066,N_5825,N_5766);
nor U6067 (N_6067,N_5914,N_5812);
nor U6068 (N_6068,N_5949,N_5774);
nor U6069 (N_6069,N_5750,N_5907);
nand U6070 (N_6070,N_5915,N_5778);
and U6071 (N_6071,N_5863,N_5745);
nor U6072 (N_6072,N_5786,N_5757);
or U6073 (N_6073,N_5717,N_5838);
and U6074 (N_6074,N_5943,N_5872);
or U6075 (N_6075,N_5946,N_5857);
nand U6076 (N_6076,N_5842,N_5925);
nor U6077 (N_6077,N_5987,N_5848);
nor U6078 (N_6078,N_5741,N_5975);
or U6079 (N_6079,N_5731,N_5832);
nand U6080 (N_6080,N_5758,N_5721);
nand U6081 (N_6081,N_5902,N_5847);
or U6082 (N_6082,N_5805,N_5926);
nor U6083 (N_6083,N_5789,N_5988);
nor U6084 (N_6084,N_5923,N_5808);
and U6085 (N_6085,N_5935,N_5804);
and U6086 (N_6086,N_5807,N_5909);
xor U6087 (N_6087,N_5856,N_5708);
and U6088 (N_6088,N_5855,N_5819);
xor U6089 (N_6089,N_5810,N_5761);
and U6090 (N_6090,N_5965,N_5754);
xor U6091 (N_6091,N_5871,N_5869);
or U6092 (N_6092,N_5803,N_5971);
nand U6093 (N_6093,N_5973,N_5961);
or U6094 (N_6094,N_5955,N_5962);
and U6095 (N_6095,N_5905,N_5932);
nor U6096 (N_6096,N_5779,N_5892);
nor U6097 (N_6097,N_5922,N_5709);
and U6098 (N_6098,N_5908,N_5967);
xor U6099 (N_6099,N_5960,N_5992);
or U6100 (N_6100,N_5824,N_5843);
xnor U6101 (N_6101,N_5760,N_5835);
and U6102 (N_6102,N_5875,N_5972);
nor U6103 (N_6103,N_5999,N_5800);
and U6104 (N_6104,N_5706,N_5818);
and U6105 (N_6105,N_5737,N_5764);
nor U6106 (N_6106,N_5762,N_5969);
and U6107 (N_6107,N_5729,N_5936);
nor U6108 (N_6108,N_5858,N_5851);
xor U6109 (N_6109,N_5916,N_5742);
nand U6110 (N_6110,N_5833,N_5974);
and U6111 (N_6111,N_5783,N_5735);
or U6112 (N_6112,N_5979,N_5864);
or U6113 (N_6113,N_5747,N_5859);
nor U6114 (N_6114,N_5845,N_5837);
xor U6115 (N_6115,N_5958,N_5740);
nor U6116 (N_6116,N_5982,N_5777);
nor U6117 (N_6117,N_5767,N_5776);
xor U6118 (N_6118,N_5763,N_5815);
xnor U6119 (N_6119,N_5726,N_5944);
or U6120 (N_6120,N_5861,N_5894);
xnor U6121 (N_6121,N_5903,N_5854);
nor U6122 (N_6122,N_5931,N_5977);
nor U6123 (N_6123,N_5732,N_5950);
and U6124 (N_6124,N_5743,N_5784);
or U6125 (N_6125,N_5890,N_5981);
and U6126 (N_6126,N_5795,N_5978);
or U6127 (N_6127,N_5991,N_5852);
and U6128 (N_6128,N_5886,N_5941);
xnor U6129 (N_6129,N_5912,N_5730);
or U6130 (N_6130,N_5752,N_5823);
nor U6131 (N_6131,N_5874,N_5723);
nand U6132 (N_6132,N_5957,N_5822);
and U6133 (N_6133,N_5802,N_5714);
and U6134 (N_6134,N_5765,N_5796);
nand U6135 (N_6135,N_5720,N_5753);
or U6136 (N_6136,N_5920,N_5719);
and U6137 (N_6137,N_5829,N_5790);
nand U6138 (N_6138,N_5888,N_5801);
nor U6139 (N_6139,N_5834,N_5728);
or U6140 (N_6140,N_5879,N_5963);
nor U6141 (N_6141,N_5933,N_5993);
or U6142 (N_6142,N_5849,N_5770);
xnor U6143 (N_6143,N_5811,N_5939);
or U6144 (N_6144,N_5839,N_5984);
xor U6145 (N_6145,N_5945,N_5989);
nor U6146 (N_6146,N_5711,N_5968);
xnor U6147 (N_6147,N_5733,N_5840);
and U6148 (N_6148,N_5771,N_5940);
xor U6149 (N_6149,N_5813,N_5744);
xor U6150 (N_6150,N_5895,N_5780);
nand U6151 (N_6151,N_5942,N_5788);
nor U6152 (N_6152,N_5812,N_5897);
nand U6153 (N_6153,N_5717,N_5702);
or U6154 (N_6154,N_5871,N_5975);
nor U6155 (N_6155,N_5861,N_5712);
or U6156 (N_6156,N_5874,N_5753);
nor U6157 (N_6157,N_5928,N_5852);
nor U6158 (N_6158,N_5958,N_5718);
nand U6159 (N_6159,N_5991,N_5794);
or U6160 (N_6160,N_5733,N_5954);
or U6161 (N_6161,N_5842,N_5852);
or U6162 (N_6162,N_5772,N_5870);
or U6163 (N_6163,N_5816,N_5718);
nand U6164 (N_6164,N_5867,N_5954);
nor U6165 (N_6165,N_5866,N_5975);
or U6166 (N_6166,N_5971,N_5767);
nor U6167 (N_6167,N_5711,N_5942);
and U6168 (N_6168,N_5942,N_5921);
or U6169 (N_6169,N_5841,N_5788);
or U6170 (N_6170,N_5989,N_5747);
nor U6171 (N_6171,N_5900,N_5871);
and U6172 (N_6172,N_5991,N_5933);
nor U6173 (N_6173,N_5816,N_5790);
nor U6174 (N_6174,N_5855,N_5976);
nand U6175 (N_6175,N_5968,N_5763);
and U6176 (N_6176,N_5772,N_5752);
xor U6177 (N_6177,N_5747,N_5840);
xor U6178 (N_6178,N_5912,N_5886);
and U6179 (N_6179,N_5991,N_5739);
nor U6180 (N_6180,N_5968,N_5976);
nor U6181 (N_6181,N_5785,N_5723);
nand U6182 (N_6182,N_5843,N_5865);
nand U6183 (N_6183,N_5856,N_5903);
or U6184 (N_6184,N_5847,N_5772);
nor U6185 (N_6185,N_5907,N_5944);
and U6186 (N_6186,N_5719,N_5768);
nor U6187 (N_6187,N_5885,N_5924);
xor U6188 (N_6188,N_5757,N_5842);
and U6189 (N_6189,N_5980,N_5702);
and U6190 (N_6190,N_5892,N_5869);
or U6191 (N_6191,N_5907,N_5880);
nor U6192 (N_6192,N_5823,N_5926);
and U6193 (N_6193,N_5848,N_5762);
or U6194 (N_6194,N_5949,N_5843);
nor U6195 (N_6195,N_5936,N_5819);
xnor U6196 (N_6196,N_5732,N_5921);
xor U6197 (N_6197,N_5983,N_5861);
nand U6198 (N_6198,N_5911,N_5939);
xor U6199 (N_6199,N_5847,N_5901);
or U6200 (N_6200,N_5916,N_5740);
and U6201 (N_6201,N_5784,N_5950);
or U6202 (N_6202,N_5956,N_5900);
xor U6203 (N_6203,N_5915,N_5958);
and U6204 (N_6204,N_5734,N_5816);
nor U6205 (N_6205,N_5711,N_5703);
or U6206 (N_6206,N_5738,N_5887);
nor U6207 (N_6207,N_5757,N_5730);
or U6208 (N_6208,N_5886,N_5873);
nor U6209 (N_6209,N_5970,N_5917);
nor U6210 (N_6210,N_5855,N_5806);
or U6211 (N_6211,N_5750,N_5981);
or U6212 (N_6212,N_5857,N_5937);
and U6213 (N_6213,N_5779,N_5789);
or U6214 (N_6214,N_5770,N_5899);
or U6215 (N_6215,N_5786,N_5888);
nor U6216 (N_6216,N_5896,N_5726);
nand U6217 (N_6217,N_5749,N_5944);
nor U6218 (N_6218,N_5940,N_5715);
or U6219 (N_6219,N_5886,N_5927);
nand U6220 (N_6220,N_5740,N_5894);
or U6221 (N_6221,N_5916,N_5871);
xor U6222 (N_6222,N_5897,N_5964);
or U6223 (N_6223,N_5867,N_5759);
xnor U6224 (N_6224,N_5810,N_5767);
xnor U6225 (N_6225,N_5869,N_5754);
or U6226 (N_6226,N_5982,N_5718);
and U6227 (N_6227,N_5770,N_5803);
nand U6228 (N_6228,N_5934,N_5791);
xnor U6229 (N_6229,N_5823,N_5865);
nand U6230 (N_6230,N_5985,N_5975);
nand U6231 (N_6231,N_5714,N_5975);
nor U6232 (N_6232,N_5703,N_5733);
and U6233 (N_6233,N_5710,N_5938);
nor U6234 (N_6234,N_5834,N_5802);
nand U6235 (N_6235,N_5903,N_5927);
nor U6236 (N_6236,N_5900,N_5845);
nand U6237 (N_6237,N_5726,N_5739);
nand U6238 (N_6238,N_5927,N_5992);
and U6239 (N_6239,N_5916,N_5858);
xnor U6240 (N_6240,N_5853,N_5852);
nand U6241 (N_6241,N_5785,N_5885);
nor U6242 (N_6242,N_5877,N_5774);
xor U6243 (N_6243,N_5889,N_5936);
and U6244 (N_6244,N_5880,N_5961);
nor U6245 (N_6245,N_5829,N_5817);
nand U6246 (N_6246,N_5911,N_5960);
xor U6247 (N_6247,N_5798,N_5937);
and U6248 (N_6248,N_5762,N_5967);
and U6249 (N_6249,N_5743,N_5701);
or U6250 (N_6250,N_5908,N_5907);
or U6251 (N_6251,N_5917,N_5889);
nand U6252 (N_6252,N_5949,N_5926);
or U6253 (N_6253,N_5958,N_5988);
nand U6254 (N_6254,N_5831,N_5762);
xor U6255 (N_6255,N_5941,N_5851);
nand U6256 (N_6256,N_5924,N_5966);
or U6257 (N_6257,N_5712,N_5859);
xor U6258 (N_6258,N_5961,N_5750);
nand U6259 (N_6259,N_5962,N_5812);
or U6260 (N_6260,N_5965,N_5761);
nor U6261 (N_6261,N_5906,N_5969);
xor U6262 (N_6262,N_5946,N_5861);
nor U6263 (N_6263,N_5948,N_5754);
xor U6264 (N_6264,N_5725,N_5896);
xor U6265 (N_6265,N_5761,N_5804);
and U6266 (N_6266,N_5996,N_5772);
nand U6267 (N_6267,N_5862,N_5732);
nor U6268 (N_6268,N_5721,N_5896);
and U6269 (N_6269,N_5891,N_5985);
xnor U6270 (N_6270,N_5939,N_5885);
and U6271 (N_6271,N_5822,N_5782);
nor U6272 (N_6272,N_5744,N_5705);
or U6273 (N_6273,N_5770,N_5841);
or U6274 (N_6274,N_5881,N_5760);
and U6275 (N_6275,N_5867,N_5780);
and U6276 (N_6276,N_5942,N_5864);
or U6277 (N_6277,N_5824,N_5746);
nor U6278 (N_6278,N_5890,N_5801);
nor U6279 (N_6279,N_5796,N_5972);
or U6280 (N_6280,N_5851,N_5763);
nand U6281 (N_6281,N_5768,N_5733);
nand U6282 (N_6282,N_5832,N_5739);
xor U6283 (N_6283,N_5824,N_5981);
or U6284 (N_6284,N_5866,N_5988);
nand U6285 (N_6285,N_5824,N_5769);
or U6286 (N_6286,N_5825,N_5999);
nand U6287 (N_6287,N_5794,N_5743);
nor U6288 (N_6288,N_5985,N_5798);
nand U6289 (N_6289,N_5803,N_5880);
xnor U6290 (N_6290,N_5957,N_5934);
nand U6291 (N_6291,N_5709,N_5968);
and U6292 (N_6292,N_5788,N_5846);
or U6293 (N_6293,N_5779,N_5955);
nor U6294 (N_6294,N_5766,N_5849);
nor U6295 (N_6295,N_5853,N_5906);
xnor U6296 (N_6296,N_5945,N_5958);
xor U6297 (N_6297,N_5754,N_5775);
or U6298 (N_6298,N_5902,N_5803);
nor U6299 (N_6299,N_5990,N_5775);
and U6300 (N_6300,N_6056,N_6182);
nor U6301 (N_6301,N_6090,N_6032);
xnor U6302 (N_6302,N_6287,N_6290);
and U6303 (N_6303,N_6134,N_6133);
nor U6304 (N_6304,N_6183,N_6249);
or U6305 (N_6305,N_6034,N_6064);
nand U6306 (N_6306,N_6123,N_6130);
or U6307 (N_6307,N_6279,N_6169);
nand U6308 (N_6308,N_6233,N_6283);
and U6309 (N_6309,N_6068,N_6266);
or U6310 (N_6310,N_6288,N_6272);
nand U6311 (N_6311,N_6122,N_6057);
nor U6312 (N_6312,N_6031,N_6170);
and U6313 (N_6313,N_6291,N_6231);
xnor U6314 (N_6314,N_6007,N_6275);
nor U6315 (N_6315,N_6158,N_6069);
and U6316 (N_6316,N_6222,N_6281);
nor U6317 (N_6317,N_6033,N_6001);
and U6318 (N_6318,N_6053,N_6005);
xor U6319 (N_6319,N_6148,N_6145);
nand U6320 (N_6320,N_6025,N_6129);
and U6321 (N_6321,N_6294,N_6297);
or U6322 (N_6322,N_6230,N_6255);
or U6323 (N_6323,N_6116,N_6024);
nor U6324 (N_6324,N_6191,N_6100);
xor U6325 (N_6325,N_6017,N_6235);
xnor U6326 (N_6326,N_6175,N_6135);
nor U6327 (N_6327,N_6040,N_6105);
nor U6328 (N_6328,N_6271,N_6195);
or U6329 (N_6329,N_6089,N_6298);
xor U6330 (N_6330,N_6002,N_6225);
and U6331 (N_6331,N_6164,N_6015);
nand U6332 (N_6332,N_6193,N_6120);
and U6333 (N_6333,N_6160,N_6054);
xor U6334 (N_6334,N_6150,N_6096);
xor U6335 (N_6335,N_6264,N_6192);
xor U6336 (N_6336,N_6085,N_6003);
or U6337 (N_6337,N_6016,N_6178);
nand U6338 (N_6338,N_6119,N_6239);
or U6339 (N_6339,N_6111,N_6062);
and U6340 (N_6340,N_6186,N_6240);
xnor U6341 (N_6341,N_6000,N_6167);
or U6342 (N_6342,N_6189,N_6163);
nor U6343 (N_6343,N_6241,N_6204);
and U6344 (N_6344,N_6126,N_6087);
xnor U6345 (N_6345,N_6285,N_6083);
nand U6346 (N_6346,N_6152,N_6194);
and U6347 (N_6347,N_6156,N_6095);
nor U6348 (N_6348,N_6277,N_6099);
or U6349 (N_6349,N_6199,N_6070);
or U6350 (N_6350,N_6219,N_6282);
xnor U6351 (N_6351,N_6209,N_6008);
nor U6352 (N_6352,N_6196,N_6212);
or U6353 (N_6353,N_6045,N_6162);
or U6354 (N_6354,N_6102,N_6121);
and U6355 (N_6355,N_6037,N_6161);
xnor U6356 (N_6356,N_6112,N_6205);
or U6357 (N_6357,N_6187,N_6103);
or U6358 (N_6358,N_6038,N_6139);
xnor U6359 (N_6359,N_6289,N_6220);
xnor U6360 (N_6360,N_6088,N_6251);
or U6361 (N_6361,N_6092,N_6246);
and U6362 (N_6362,N_6138,N_6014);
nor U6363 (N_6363,N_6159,N_6080);
and U6364 (N_6364,N_6206,N_6118);
and U6365 (N_6365,N_6259,N_6256);
or U6366 (N_6366,N_6276,N_6079);
or U6367 (N_6367,N_6197,N_6278);
or U6368 (N_6368,N_6261,N_6142);
nand U6369 (N_6369,N_6201,N_6188);
and U6370 (N_6370,N_6210,N_6208);
xor U6371 (N_6371,N_6023,N_6022);
nor U6372 (N_6372,N_6166,N_6232);
xnor U6373 (N_6373,N_6216,N_6243);
xor U6374 (N_6374,N_6157,N_6009);
xor U6375 (N_6375,N_6097,N_6078);
xnor U6376 (N_6376,N_6151,N_6213);
and U6377 (N_6377,N_6013,N_6149);
or U6378 (N_6378,N_6153,N_6248);
nor U6379 (N_6379,N_6128,N_6245);
nand U6380 (N_6380,N_6190,N_6106);
or U6381 (N_6381,N_6073,N_6052);
or U6382 (N_6382,N_6082,N_6146);
nor U6383 (N_6383,N_6177,N_6094);
nor U6384 (N_6384,N_6200,N_6262);
xor U6385 (N_6385,N_6039,N_6026);
xnor U6386 (N_6386,N_6173,N_6211);
and U6387 (N_6387,N_6066,N_6081);
or U6388 (N_6388,N_6260,N_6051);
or U6389 (N_6389,N_6048,N_6144);
xor U6390 (N_6390,N_6136,N_6113);
nand U6391 (N_6391,N_6067,N_6027);
nand U6392 (N_6392,N_6084,N_6036);
xor U6393 (N_6393,N_6254,N_6218);
or U6394 (N_6394,N_6242,N_6109);
and U6395 (N_6395,N_6041,N_6217);
or U6396 (N_6396,N_6234,N_6131);
nand U6397 (N_6397,N_6270,N_6117);
nand U6398 (N_6398,N_6093,N_6280);
nor U6399 (N_6399,N_6250,N_6165);
nor U6400 (N_6400,N_6274,N_6171);
and U6401 (N_6401,N_6006,N_6252);
nor U6402 (N_6402,N_6228,N_6143);
xor U6403 (N_6403,N_6107,N_6207);
nand U6404 (N_6404,N_6059,N_6044);
or U6405 (N_6405,N_6286,N_6202);
or U6406 (N_6406,N_6018,N_6077);
and U6407 (N_6407,N_6176,N_6227);
nand U6408 (N_6408,N_6299,N_6247);
nor U6409 (N_6409,N_6020,N_6168);
and U6410 (N_6410,N_6257,N_6074);
and U6411 (N_6411,N_6137,N_6236);
nor U6412 (N_6412,N_6238,N_6114);
nor U6413 (N_6413,N_6125,N_6035);
and U6414 (N_6414,N_6141,N_6058);
nor U6415 (N_6415,N_6091,N_6147);
nor U6416 (N_6416,N_6075,N_6229);
and U6417 (N_6417,N_6174,N_6098);
or U6418 (N_6418,N_6019,N_6071);
nor U6419 (N_6419,N_6004,N_6042);
nor U6420 (N_6420,N_6172,N_6110);
or U6421 (N_6421,N_6104,N_6203);
and U6422 (N_6422,N_6223,N_6132);
xnor U6423 (N_6423,N_6292,N_6224);
xor U6424 (N_6424,N_6076,N_6108);
nor U6425 (N_6425,N_6061,N_6127);
or U6426 (N_6426,N_6215,N_6010);
nand U6427 (N_6427,N_6124,N_6180);
nor U6428 (N_6428,N_6060,N_6226);
or U6429 (N_6429,N_6030,N_6185);
and U6430 (N_6430,N_6181,N_6214);
or U6431 (N_6431,N_6293,N_6029);
and U6432 (N_6432,N_6063,N_6237);
or U6433 (N_6433,N_6179,N_6268);
or U6434 (N_6434,N_6043,N_6140);
nor U6435 (N_6435,N_6273,N_6263);
or U6436 (N_6436,N_6046,N_6047);
xnor U6437 (N_6437,N_6284,N_6184);
and U6438 (N_6438,N_6198,N_6086);
nand U6439 (N_6439,N_6011,N_6295);
xor U6440 (N_6440,N_6265,N_6021);
nor U6441 (N_6441,N_6012,N_6267);
or U6442 (N_6442,N_6028,N_6049);
nand U6443 (N_6443,N_6296,N_6221);
nor U6444 (N_6444,N_6055,N_6269);
nand U6445 (N_6445,N_6244,N_6115);
nor U6446 (N_6446,N_6072,N_6101);
nand U6447 (N_6447,N_6253,N_6154);
nor U6448 (N_6448,N_6050,N_6065);
nand U6449 (N_6449,N_6155,N_6258);
nand U6450 (N_6450,N_6185,N_6127);
nor U6451 (N_6451,N_6139,N_6154);
or U6452 (N_6452,N_6223,N_6104);
nor U6453 (N_6453,N_6158,N_6137);
nand U6454 (N_6454,N_6046,N_6122);
nand U6455 (N_6455,N_6040,N_6071);
nand U6456 (N_6456,N_6020,N_6231);
or U6457 (N_6457,N_6149,N_6260);
or U6458 (N_6458,N_6221,N_6277);
and U6459 (N_6459,N_6264,N_6207);
nor U6460 (N_6460,N_6203,N_6246);
or U6461 (N_6461,N_6149,N_6111);
xnor U6462 (N_6462,N_6069,N_6066);
nor U6463 (N_6463,N_6182,N_6197);
nand U6464 (N_6464,N_6286,N_6199);
nor U6465 (N_6465,N_6249,N_6274);
and U6466 (N_6466,N_6033,N_6067);
xor U6467 (N_6467,N_6034,N_6199);
xor U6468 (N_6468,N_6128,N_6109);
or U6469 (N_6469,N_6255,N_6122);
xor U6470 (N_6470,N_6081,N_6097);
or U6471 (N_6471,N_6079,N_6148);
or U6472 (N_6472,N_6159,N_6236);
nand U6473 (N_6473,N_6026,N_6127);
xnor U6474 (N_6474,N_6204,N_6175);
and U6475 (N_6475,N_6104,N_6190);
nor U6476 (N_6476,N_6118,N_6097);
xor U6477 (N_6477,N_6287,N_6158);
nand U6478 (N_6478,N_6214,N_6100);
nand U6479 (N_6479,N_6202,N_6053);
or U6480 (N_6480,N_6115,N_6051);
and U6481 (N_6481,N_6107,N_6223);
or U6482 (N_6482,N_6122,N_6055);
nand U6483 (N_6483,N_6228,N_6071);
nor U6484 (N_6484,N_6002,N_6081);
nand U6485 (N_6485,N_6060,N_6194);
and U6486 (N_6486,N_6180,N_6199);
nor U6487 (N_6487,N_6289,N_6104);
and U6488 (N_6488,N_6098,N_6198);
nand U6489 (N_6489,N_6116,N_6046);
xor U6490 (N_6490,N_6056,N_6175);
nand U6491 (N_6491,N_6217,N_6074);
nor U6492 (N_6492,N_6123,N_6116);
and U6493 (N_6493,N_6027,N_6101);
xor U6494 (N_6494,N_6225,N_6061);
or U6495 (N_6495,N_6252,N_6213);
nor U6496 (N_6496,N_6236,N_6070);
and U6497 (N_6497,N_6179,N_6129);
nor U6498 (N_6498,N_6005,N_6071);
nand U6499 (N_6499,N_6216,N_6090);
nand U6500 (N_6500,N_6284,N_6285);
or U6501 (N_6501,N_6248,N_6044);
xor U6502 (N_6502,N_6146,N_6208);
nand U6503 (N_6503,N_6012,N_6026);
nand U6504 (N_6504,N_6223,N_6263);
nor U6505 (N_6505,N_6256,N_6274);
nor U6506 (N_6506,N_6251,N_6109);
nand U6507 (N_6507,N_6178,N_6002);
nor U6508 (N_6508,N_6288,N_6065);
nand U6509 (N_6509,N_6109,N_6173);
nand U6510 (N_6510,N_6198,N_6150);
nand U6511 (N_6511,N_6182,N_6031);
or U6512 (N_6512,N_6286,N_6192);
or U6513 (N_6513,N_6232,N_6188);
or U6514 (N_6514,N_6022,N_6139);
nand U6515 (N_6515,N_6228,N_6094);
xnor U6516 (N_6516,N_6253,N_6298);
or U6517 (N_6517,N_6208,N_6186);
nor U6518 (N_6518,N_6133,N_6187);
and U6519 (N_6519,N_6023,N_6052);
nand U6520 (N_6520,N_6259,N_6069);
nand U6521 (N_6521,N_6276,N_6072);
nand U6522 (N_6522,N_6039,N_6075);
nor U6523 (N_6523,N_6011,N_6117);
nor U6524 (N_6524,N_6087,N_6181);
and U6525 (N_6525,N_6272,N_6178);
nor U6526 (N_6526,N_6171,N_6039);
and U6527 (N_6527,N_6261,N_6279);
xor U6528 (N_6528,N_6210,N_6209);
nand U6529 (N_6529,N_6103,N_6260);
or U6530 (N_6530,N_6252,N_6240);
or U6531 (N_6531,N_6269,N_6035);
xnor U6532 (N_6532,N_6251,N_6047);
xor U6533 (N_6533,N_6186,N_6196);
nand U6534 (N_6534,N_6108,N_6014);
and U6535 (N_6535,N_6039,N_6260);
nor U6536 (N_6536,N_6091,N_6279);
xor U6537 (N_6537,N_6021,N_6256);
xor U6538 (N_6538,N_6240,N_6046);
and U6539 (N_6539,N_6002,N_6014);
nor U6540 (N_6540,N_6238,N_6207);
nand U6541 (N_6541,N_6103,N_6119);
and U6542 (N_6542,N_6173,N_6188);
xor U6543 (N_6543,N_6093,N_6158);
nand U6544 (N_6544,N_6052,N_6059);
and U6545 (N_6545,N_6289,N_6154);
xnor U6546 (N_6546,N_6135,N_6057);
and U6547 (N_6547,N_6298,N_6281);
nand U6548 (N_6548,N_6246,N_6021);
xnor U6549 (N_6549,N_6142,N_6117);
nand U6550 (N_6550,N_6185,N_6063);
and U6551 (N_6551,N_6180,N_6140);
and U6552 (N_6552,N_6051,N_6161);
nand U6553 (N_6553,N_6137,N_6081);
nor U6554 (N_6554,N_6068,N_6167);
nor U6555 (N_6555,N_6011,N_6249);
and U6556 (N_6556,N_6198,N_6189);
xnor U6557 (N_6557,N_6288,N_6165);
nor U6558 (N_6558,N_6264,N_6137);
nor U6559 (N_6559,N_6114,N_6251);
nor U6560 (N_6560,N_6019,N_6281);
and U6561 (N_6561,N_6240,N_6038);
or U6562 (N_6562,N_6022,N_6097);
or U6563 (N_6563,N_6176,N_6125);
nor U6564 (N_6564,N_6284,N_6259);
xnor U6565 (N_6565,N_6130,N_6202);
nand U6566 (N_6566,N_6111,N_6252);
nand U6567 (N_6567,N_6169,N_6290);
nand U6568 (N_6568,N_6291,N_6289);
or U6569 (N_6569,N_6133,N_6171);
nor U6570 (N_6570,N_6049,N_6103);
nor U6571 (N_6571,N_6029,N_6064);
or U6572 (N_6572,N_6094,N_6217);
nor U6573 (N_6573,N_6297,N_6232);
or U6574 (N_6574,N_6299,N_6217);
and U6575 (N_6575,N_6023,N_6042);
nor U6576 (N_6576,N_6025,N_6258);
xnor U6577 (N_6577,N_6122,N_6086);
nor U6578 (N_6578,N_6192,N_6076);
xor U6579 (N_6579,N_6292,N_6216);
xor U6580 (N_6580,N_6167,N_6252);
or U6581 (N_6581,N_6083,N_6154);
or U6582 (N_6582,N_6271,N_6289);
or U6583 (N_6583,N_6052,N_6228);
and U6584 (N_6584,N_6153,N_6143);
nand U6585 (N_6585,N_6226,N_6178);
and U6586 (N_6586,N_6272,N_6069);
nor U6587 (N_6587,N_6173,N_6243);
or U6588 (N_6588,N_6137,N_6079);
nand U6589 (N_6589,N_6221,N_6018);
or U6590 (N_6590,N_6259,N_6196);
nor U6591 (N_6591,N_6207,N_6149);
or U6592 (N_6592,N_6283,N_6004);
nand U6593 (N_6593,N_6063,N_6187);
or U6594 (N_6594,N_6152,N_6271);
nor U6595 (N_6595,N_6097,N_6089);
nand U6596 (N_6596,N_6152,N_6062);
nor U6597 (N_6597,N_6167,N_6044);
and U6598 (N_6598,N_6120,N_6251);
or U6599 (N_6599,N_6279,N_6054);
and U6600 (N_6600,N_6492,N_6578);
or U6601 (N_6601,N_6309,N_6437);
nand U6602 (N_6602,N_6331,N_6398);
xor U6603 (N_6603,N_6342,N_6462);
and U6604 (N_6604,N_6587,N_6314);
nand U6605 (N_6605,N_6470,N_6304);
or U6606 (N_6606,N_6411,N_6307);
xnor U6607 (N_6607,N_6420,N_6491);
nor U6608 (N_6608,N_6426,N_6343);
nor U6609 (N_6609,N_6341,N_6313);
or U6610 (N_6610,N_6523,N_6532);
and U6611 (N_6611,N_6524,N_6529);
or U6612 (N_6612,N_6402,N_6436);
nand U6613 (N_6613,N_6427,N_6435);
and U6614 (N_6614,N_6486,N_6338);
and U6615 (N_6615,N_6424,N_6458);
xor U6616 (N_6616,N_6315,N_6325);
nand U6617 (N_6617,N_6548,N_6444);
nor U6618 (N_6618,N_6316,N_6335);
nor U6619 (N_6619,N_6405,N_6319);
or U6620 (N_6620,N_6336,N_6599);
nand U6621 (N_6621,N_6536,N_6428);
nor U6622 (N_6622,N_6355,N_6417);
and U6623 (N_6623,N_6590,N_6572);
nor U6624 (N_6624,N_6303,N_6448);
nand U6625 (N_6625,N_6544,N_6456);
nand U6626 (N_6626,N_6347,N_6306);
and U6627 (N_6627,N_6585,N_6445);
or U6628 (N_6628,N_6570,N_6305);
or U6629 (N_6629,N_6418,N_6328);
nor U6630 (N_6630,N_6369,N_6332);
nor U6631 (N_6631,N_6494,N_6560);
xnor U6632 (N_6632,N_6518,N_6395);
nand U6633 (N_6633,N_6477,N_6324);
nor U6634 (N_6634,N_6597,N_6553);
or U6635 (N_6635,N_6408,N_6471);
or U6636 (N_6636,N_6479,N_6483);
nor U6637 (N_6637,N_6413,N_6583);
xor U6638 (N_6638,N_6528,N_6360);
nand U6639 (N_6639,N_6357,N_6453);
xnor U6640 (N_6640,N_6521,N_6459);
xnor U6641 (N_6641,N_6511,N_6588);
or U6642 (N_6642,N_6412,N_6488);
and U6643 (N_6643,N_6441,N_6401);
nand U6644 (N_6644,N_6558,N_6562);
and U6645 (N_6645,N_6559,N_6500);
and U6646 (N_6646,N_6551,N_6541);
and U6647 (N_6647,N_6552,N_6454);
nand U6648 (N_6648,N_6443,N_6502);
or U6649 (N_6649,N_6537,N_6423);
xnor U6650 (N_6650,N_6564,N_6384);
nor U6651 (N_6651,N_6480,N_6390);
xor U6652 (N_6652,N_6352,N_6584);
nand U6653 (N_6653,N_6365,N_6340);
and U6654 (N_6654,N_6493,N_6510);
xor U6655 (N_6655,N_6375,N_6556);
and U6656 (N_6656,N_6586,N_6526);
or U6657 (N_6657,N_6542,N_6362);
or U6658 (N_6658,N_6574,N_6466);
and U6659 (N_6659,N_6476,N_6378);
and U6660 (N_6660,N_6356,N_6465);
and U6661 (N_6661,N_6414,N_6487);
xnor U6662 (N_6662,N_6387,N_6563);
nand U6663 (N_6663,N_6374,N_6457);
xor U6664 (N_6664,N_6580,N_6391);
and U6665 (N_6665,N_6567,N_6593);
or U6666 (N_6666,N_6372,N_6345);
and U6667 (N_6667,N_6344,N_6368);
nand U6668 (N_6668,N_6379,N_6533);
and U6669 (N_6669,N_6359,N_6392);
xnor U6670 (N_6670,N_6404,N_6400);
nor U6671 (N_6671,N_6576,N_6527);
nand U6672 (N_6672,N_6485,N_6531);
xor U6673 (N_6673,N_6322,N_6376);
nand U6674 (N_6674,N_6538,N_6535);
nor U6675 (N_6675,N_6380,N_6449);
nand U6676 (N_6676,N_6482,N_6589);
nand U6677 (N_6677,N_6358,N_6591);
nor U6678 (N_6678,N_6351,N_6568);
or U6679 (N_6679,N_6549,N_6433);
or U6680 (N_6680,N_6547,N_6419);
nand U6681 (N_6681,N_6311,N_6489);
or U6682 (N_6682,N_6321,N_6337);
or U6683 (N_6683,N_6403,N_6429);
nor U6684 (N_6684,N_6468,N_6582);
and U6685 (N_6685,N_6312,N_6410);
nor U6686 (N_6686,N_6363,N_6354);
nor U6687 (N_6687,N_6506,N_6475);
nand U6688 (N_6688,N_6478,N_6383);
nand U6689 (N_6689,N_6349,N_6519);
nand U6690 (N_6690,N_6407,N_6498);
nor U6691 (N_6691,N_6543,N_6460);
nand U6692 (N_6692,N_6434,N_6496);
or U6693 (N_6693,N_6490,N_6565);
nor U6694 (N_6694,N_6495,N_6333);
or U6695 (N_6695,N_6366,N_6571);
and U6696 (N_6696,N_6432,N_6581);
nor U6697 (N_6697,N_6422,N_6421);
nor U6698 (N_6698,N_6416,N_6330);
or U6699 (N_6699,N_6353,N_6598);
or U6700 (N_6700,N_6439,N_6509);
or U6701 (N_6701,N_6323,N_6367);
nor U6702 (N_6702,N_6517,N_6442);
nand U6703 (N_6703,N_6450,N_6302);
xnor U6704 (N_6704,N_6399,N_6447);
nor U6705 (N_6705,N_6569,N_6546);
nand U6706 (N_6706,N_6361,N_6516);
nor U6707 (N_6707,N_6440,N_6386);
or U6708 (N_6708,N_6566,N_6555);
nand U6709 (N_6709,N_6388,N_6455);
nand U6710 (N_6710,N_6438,N_6310);
xnor U6711 (N_6711,N_6451,N_6515);
nand U6712 (N_6712,N_6406,N_6525);
and U6713 (N_6713,N_6463,N_6393);
nor U6714 (N_6714,N_6339,N_6539);
and U6715 (N_6715,N_6503,N_6575);
nor U6716 (N_6716,N_6484,N_6320);
nand U6717 (N_6717,N_6594,N_6508);
or U6718 (N_6718,N_6327,N_6308);
and U6719 (N_6719,N_6514,N_6377);
nand U6720 (N_6720,N_6512,N_6394);
xor U6721 (N_6721,N_6317,N_6497);
and U6722 (N_6722,N_6329,N_6334);
nand U6723 (N_6723,N_6431,N_6467);
nor U6724 (N_6724,N_6504,N_6561);
nand U6725 (N_6725,N_6592,N_6550);
nor U6726 (N_6726,N_6326,N_6596);
nand U6727 (N_6727,N_6513,N_6481);
xnor U6728 (N_6728,N_6425,N_6579);
and U6729 (N_6729,N_6385,N_6446);
and U6730 (N_6730,N_6505,N_6534);
nand U6731 (N_6731,N_6499,N_6573);
and U6732 (N_6732,N_6472,N_6373);
nand U6733 (N_6733,N_6522,N_6554);
and U6734 (N_6734,N_6545,N_6430);
xnor U6735 (N_6735,N_6577,N_6409);
nand U6736 (N_6736,N_6507,N_6530);
xnor U6737 (N_6737,N_6381,N_6389);
and U6738 (N_6738,N_6371,N_6540);
and U6739 (N_6739,N_6397,N_6469);
and U6740 (N_6740,N_6348,N_6520);
xnor U6741 (N_6741,N_6300,N_6464);
nand U6742 (N_6742,N_6595,N_6452);
nand U6743 (N_6743,N_6473,N_6318);
nand U6744 (N_6744,N_6474,N_6350);
xor U6745 (N_6745,N_6461,N_6557);
xor U6746 (N_6746,N_6396,N_6415);
nor U6747 (N_6747,N_6346,N_6301);
nand U6748 (N_6748,N_6501,N_6364);
nand U6749 (N_6749,N_6382,N_6370);
nand U6750 (N_6750,N_6359,N_6533);
and U6751 (N_6751,N_6544,N_6567);
nor U6752 (N_6752,N_6311,N_6403);
nand U6753 (N_6753,N_6469,N_6598);
nor U6754 (N_6754,N_6535,N_6558);
nor U6755 (N_6755,N_6424,N_6358);
nor U6756 (N_6756,N_6339,N_6395);
and U6757 (N_6757,N_6325,N_6410);
or U6758 (N_6758,N_6492,N_6477);
and U6759 (N_6759,N_6584,N_6365);
or U6760 (N_6760,N_6404,N_6535);
or U6761 (N_6761,N_6455,N_6312);
or U6762 (N_6762,N_6493,N_6431);
and U6763 (N_6763,N_6414,N_6309);
nand U6764 (N_6764,N_6513,N_6355);
nor U6765 (N_6765,N_6591,N_6477);
or U6766 (N_6766,N_6452,N_6434);
or U6767 (N_6767,N_6348,N_6314);
nand U6768 (N_6768,N_6513,N_6501);
and U6769 (N_6769,N_6512,N_6352);
and U6770 (N_6770,N_6503,N_6322);
and U6771 (N_6771,N_6373,N_6541);
or U6772 (N_6772,N_6348,N_6456);
xnor U6773 (N_6773,N_6485,N_6526);
nor U6774 (N_6774,N_6461,N_6564);
and U6775 (N_6775,N_6444,N_6406);
nand U6776 (N_6776,N_6474,N_6555);
nor U6777 (N_6777,N_6451,N_6327);
nand U6778 (N_6778,N_6388,N_6576);
nand U6779 (N_6779,N_6588,N_6453);
and U6780 (N_6780,N_6443,N_6590);
or U6781 (N_6781,N_6397,N_6399);
nand U6782 (N_6782,N_6473,N_6364);
nor U6783 (N_6783,N_6449,N_6422);
or U6784 (N_6784,N_6564,N_6326);
and U6785 (N_6785,N_6354,N_6404);
nand U6786 (N_6786,N_6499,N_6300);
xnor U6787 (N_6787,N_6553,N_6332);
nor U6788 (N_6788,N_6549,N_6476);
nand U6789 (N_6789,N_6599,N_6348);
nor U6790 (N_6790,N_6440,N_6432);
xor U6791 (N_6791,N_6340,N_6371);
or U6792 (N_6792,N_6522,N_6417);
or U6793 (N_6793,N_6473,N_6326);
or U6794 (N_6794,N_6529,N_6562);
nor U6795 (N_6795,N_6363,N_6401);
nand U6796 (N_6796,N_6503,N_6348);
nor U6797 (N_6797,N_6487,N_6466);
nand U6798 (N_6798,N_6572,N_6520);
xnor U6799 (N_6799,N_6421,N_6394);
xnor U6800 (N_6800,N_6395,N_6375);
xor U6801 (N_6801,N_6415,N_6538);
xnor U6802 (N_6802,N_6446,N_6499);
nand U6803 (N_6803,N_6428,N_6453);
nor U6804 (N_6804,N_6388,N_6533);
or U6805 (N_6805,N_6543,N_6438);
nor U6806 (N_6806,N_6465,N_6377);
nor U6807 (N_6807,N_6563,N_6311);
or U6808 (N_6808,N_6406,N_6440);
and U6809 (N_6809,N_6469,N_6382);
xnor U6810 (N_6810,N_6321,N_6585);
xnor U6811 (N_6811,N_6515,N_6346);
nor U6812 (N_6812,N_6545,N_6363);
and U6813 (N_6813,N_6584,N_6427);
and U6814 (N_6814,N_6463,N_6453);
xor U6815 (N_6815,N_6575,N_6446);
nand U6816 (N_6816,N_6349,N_6374);
and U6817 (N_6817,N_6595,N_6535);
or U6818 (N_6818,N_6410,N_6371);
and U6819 (N_6819,N_6492,N_6589);
or U6820 (N_6820,N_6359,N_6349);
xnor U6821 (N_6821,N_6311,N_6576);
nor U6822 (N_6822,N_6376,N_6399);
xnor U6823 (N_6823,N_6468,N_6361);
and U6824 (N_6824,N_6491,N_6439);
nand U6825 (N_6825,N_6430,N_6552);
or U6826 (N_6826,N_6487,N_6308);
and U6827 (N_6827,N_6320,N_6572);
and U6828 (N_6828,N_6596,N_6425);
xnor U6829 (N_6829,N_6513,N_6338);
or U6830 (N_6830,N_6578,N_6590);
and U6831 (N_6831,N_6351,N_6495);
nand U6832 (N_6832,N_6333,N_6508);
nand U6833 (N_6833,N_6515,N_6489);
xor U6834 (N_6834,N_6549,N_6323);
and U6835 (N_6835,N_6428,N_6559);
or U6836 (N_6836,N_6353,N_6373);
nand U6837 (N_6837,N_6327,N_6454);
nor U6838 (N_6838,N_6385,N_6369);
and U6839 (N_6839,N_6379,N_6471);
xnor U6840 (N_6840,N_6511,N_6418);
nor U6841 (N_6841,N_6478,N_6419);
xor U6842 (N_6842,N_6444,N_6514);
xnor U6843 (N_6843,N_6315,N_6408);
and U6844 (N_6844,N_6395,N_6393);
xor U6845 (N_6845,N_6546,N_6558);
nand U6846 (N_6846,N_6532,N_6570);
nor U6847 (N_6847,N_6367,N_6511);
or U6848 (N_6848,N_6319,N_6444);
and U6849 (N_6849,N_6461,N_6464);
or U6850 (N_6850,N_6330,N_6373);
and U6851 (N_6851,N_6497,N_6593);
and U6852 (N_6852,N_6503,N_6445);
xnor U6853 (N_6853,N_6331,N_6542);
and U6854 (N_6854,N_6419,N_6571);
or U6855 (N_6855,N_6554,N_6369);
nand U6856 (N_6856,N_6405,N_6355);
nand U6857 (N_6857,N_6436,N_6517);
and U6858 (N_6858,N_6342,N_6425);
nor U6859 (N_6859,N_6541,N_6542);
nand U6860 (N_6860,N_6387,N_6517);
xor U6861 (N_6861,N_6449,N_6468);
and U6862 (N_6862,N_6374,N_6472);
nor U6863 (N_6863,N_6373,N_6502);
nor U6864 (N_6864,N_6536,N_6326);
nand U6865 (N_6865,N_6522,N_6494);
xnor U6866 (N_6866,N_6487,N_6453);
xor U6867 (N_6867,N_6481,N_6358);
and U6868 (N_6868,N_6536,N_6425);
or U6869 (N_6869,N_6394,N_6508);
and U6870 (N_6870,N_6554,N_6327);
and U6871 (N_6871,N_6308,N_6407);
nand U6872 (N_6872,N_6545,N_6533);
or U6873 (N_6873,N_6534,N_6312);
nand U6874 (N_6874,N_6380,N_6375);
or U6875 (N_6875,N_6366,N_6568);
nand U6876 (N_6876,N_6582,N_6360);
or U6877 (N_6877,N_6566,N_6514);
nand U6878 (N_6878,N_6563,N_6394);
and U6879 (N_6879,N_6541,N_6355);
nor U6880 (N_6880,N_6504,N_6599);
nand U6881 (N_6881,N_6498,N_6527);
nand U6882 (N_6882,N_6579,N_6449);
nor U6883 (N_6883,N_6422,N_6361);
nor U6884 (N_6884,N_6312,N_6472);
and U6885 (N_6885,N_6535,N_6326);
nand U6886 (N_6886,N_6527,N_6404);
and U6887 (N_6887,N_6322,N_6442);
and U6888 (N_6888,N_6532,N_6574);
nor U6889 (N_6889,N_6504,N_6392);
or U6890 (N_6890,N_6356,N_6387);
xnor U6891 (N_6891,N_6356,N_6352);
or U6892 (N_6892,N_6453,N_6479);
nand U6893 (N_6893,N_6322,N_6539);
nand U6894 (N_6894,N_6444,N_6563);
nor U6895 (N_6895,N_6426,N_6553);
or U6896 (N_6896,N_6341,N_6478);
xor U6897 (N_6897,N_6304,N_6592);
or U6898 (N_6898,N_6442,N_6426);
nor U6899 (N_6899,N_6364,N_6349);
or U6900 (N_6900,N_6724,N_6716);
xor U6901 (N_6901,N_6699,N_6812);
and U6902 (N_6902,N_6683,N_6695);
nand U6903 (N_6903,N_6611,N_6770);
or U6904 (N_6904,N_6826,N_6800);
xnor U6905 (N_6905,N_6743,N_6814);
nor U6906 (N_6906,N_6613,N_6701);
nor U6907 (N_6907,N_6720,N_6831);
nor U6908 (N_6908,N_6628,N_6792);
xnor U6909 (N_6909,N_6672,N_6677);
nor U6910 (N_6910,N_6860,N_6855);
nand U6911 (N_6911,N_6868,N_6865);
nor U6912 (N_6912,N_6687,N_6633);
xor U6913 (N_6913,N_6734,N_6846);
nand U6914 (N_6914,N_6882,N_6785);
xor U6915 (N_6915,N_6619,N_6775);
and U6916 (N_6916,N_6781,N_6784);
and U6917 (N_6917,N_6804,N_6685);
or U6918 (N_6918,N_6643,N_6732);
or U6919 (N_6919,N_6815,N_6834);
xnor U6920 (N_6920,N_6614,N_6742);
xnor U6921 (N_6921,N_6862,N_6825);
or U6922 (N_6922,N_6659,N_6631);
nor U6923 (N_6923,N_6881,N_6893);
or U6924 (N_6924,N_6853,N_6736);
nand U6925 (N_6925,N_6609,N_6783);
nor U6926 (N_6926,N_6746,N_6637);
and U6927 (N_6927,N_6771,N_6837);
or U6928 (N_6928,N_6618,N_6680);
or U6929 (N_6929,N_6874,N_6646);
or U6930 (N_6930,N_6719,N_6739);
nor U6931 (N_6931,N_6884,N_6735);
or U6932 (N_6932,N_6610,N_6635);
nor U6933 (N_6933,N_6895,N_6844);
nand U6934 (N_6934,N_6790,N_6811);
nor U6935 (N_6935,N_6888,N_6828);
or U6936 (N_6936,N_6755,N_6647);
nor U6937 (N_6937,N_6808,N_6702);
nand U6938 (N_6938,N_6816,N_6833);
nand U6939 (N_6939,N_6607,N_6711);
nor U6940 (N_6940,N_6648,N_6839);
xor U6941 (N_6941,N_6891,N_6713);
xnor U6942 (N_6942,N_6678,N_6887);
and U6943 (N_6943,N_6866,N_6896);
xor U6944 (N_6944,N_6823,N_6747);
nor U6945 (N_6945,N_6665,N_6799);
nor U6946 (N_6946,N_6653,N_6669);
or U6947 (N_6947,N_6819,N_6776);
or U6948 (N_6948,N_6670,N_6726);
or U6949 (N_6949,N_6845,N_6754);
xor U6950 (N_6950,N_6621,N_6892);
and U6951 (N_6951,N_6897,N_6774);
xor U6952 (N_6952,N_6753,N_6675);
nor U6953 (N_6953,N_6706,N_6709);
nor U6954 (N_6954,N_6717,N_6782);
nor U6955 (N_6955,N_6615,N_6793);
and U6956 (N_6956,N_6870,N_6880);
and U6957 (N_6957,N_6883,N_6843);
or U6958 (N_6958,N_6886,N_6772);
or U6959 (N_6959,N_6662,N_6821);
and U6960 (N_6960,N_6767,N_6617);
nor U6961 (N_6961,N_6681,N_6813);
and U6962 (N_6962,N_6838,N_6822);
or U6963 (N_6963,N_6798,N_6651);
and U6964 (N_6964,N_6802,N_6778);
xor U6965 (N_6965,N_6714,N_6602);
or U6966 (N_6966,N_6649,N_6723);
xnor U6967 (N_6967,N_6829,N_6626);
nor U6968 (N_6968,N_6750,N_6780);
nor U6969 (N_6969,N_6697,N_6601);
nor U6970 (N_6970,N_6629,N_6807);
or U6971 (N_6971,N_6765,N_6638);
nand U6972 (N_6972,N_6885,N_6809);
nor U6973 (N_6973,N_6818,N_6787);
and U6974 (N_6974,N_6867,N_6803);
or U6975 (N_6975,N_6875,N_6738);
and U6976 (N_6976,N_6655,N_6759);
nor U6977 (N_6977,N_6622,N_6620);
and U6978 (N_6978,N_6877,N_6854);
and U6979 (N_6979,N_6795,N_6763);
or U6980 (N_6980,N_6715,N_6636);
nand U6981 (N_6981,N_6623,N_6700);
nor U6982 (N_6982,N_6864,N_6773);
and U6983 (N_6983,N_6805,N_6890);
nand U6984 (N_6984,N_6756,N_6645);
nor U6985 (N_6985,N_6757,N_6625);
nand U6986 (N_6986,N_6642,N_6797);
and U6987 (N_6987,N_6801,N_6725);
or U6988 (N_6988,N_6703,N_6894);
nor U6989 (N_6989,N_6796,N_6612);
and U6990 (N_6990,N_6667,N_6693);
or U6991 (N_6991,N_6654,N_6603);
nor U6992 (N_6992,N_6630,N_6737);
nand U6993 (N_6993,N_6820,N_6721);
nand U6994 (N_6994,N_6729,N_6730);
nor U6995 (N_6995,N_6824,N_6861);
xor U6996 (N_6996,N_6727,N_6663);
nand U6997 (N_6997,N_6690,N_6777);
xnor U6998 (N_6998,N_6722,N_6806);
nand U6999 (N_6999,N_6688,N_6710);
or U7000 (N_7000,N_6858,N_6879);
nor U7001 (N_7001,N_6758,N_6707);
nor U7002 (N_7002,N_6851,N_6664);
nor U7003 (N_7003,N_6691,N_6668);
or U7004 (N_7004,N_6657,N_6761);
xnor U7005 (N_7005,N_6842,N_6872);
or U7006 (N_7006,N_6682,N_6673);
nand U7007 (N_7007,N_6836,N_6731);
or U7008 (N_7008,N_6676,N_6639);
and U7009 (N_7009,N_6686,N_6658);
nand U7010 (N_7010,N_6789,N_6650);
and U7011 (N_7011,N_6627,N_6752);
nor U7012 (N_7012,N_6733,N_6661);
nand U7013 (N_7013,N_6744,N_6841);
xor U7014 (N_7014,N_6869,N_6656);
xnor U7015 (N_7015,N_6671,N_6779);
xnor U7016 (N_7016,N_6786,N_6704);
nor U7017 (N_7017,N_6689,N_6898);
xnor U7018 (N_7018,N_6679,N_6718);
nor U7019 (N_7019,N_6694,N_6764);
and U7020 (N_7020,N_6768,N_6769);
and U7021 (N_7021,N_6728,N_6641);
nor U7022 (N_7022,N_6794,N_6624);
xnor U7023 (N_7023,N_6632,N_6600);
nor U7024 (N_7024,N_6847,N_6871);
xor U7025 (N_7025,N_6741,N_6810);
nand U7026 (N_7026,N_6745,N_6840);
nor U7027 (N_7027,N_6835,N_6640);
xnor U7028 (N_7028,N_6712,N_6698);
nand U7029 (N_7029,N_6832,N_6899);
nor U7030 (N_7030,N_6705,N_6788);
xor U7031 (N_7031,N_6604,N_6766);
and U7032 (N_7032,N_6848,N_6740);
nand U7033 (N_7033,N_6876,N_6748);
nand U7034 (N_7034,N_6634,N_6863);
nand U7035 (N_7035,N_6827,N_6849);
and U7036 (N_7036,N_6644,N_6708);
and U7037 (N_7037,N_6616,N_6751);
and U7038 (N_7038,N_6674,N_6878);
or U7039 (N_7039,N_6873,N_6859);
nand U7040 (N_7040,N_6857,N_6608);
nand U7041 (N_7041,N_6852,N_6652);
xor U7042 (N_7042,N_6856,N_6660);
nor U7043 (N_7043,N_6889,N_6749);
and U7044 (N_7044,N_6762,N_6760);
xnor U7045 (N_7045,N_6605,N_6684);
or U7046 (N_7046,N_6830,N_6692);
or U7047 (N_7047,N_6850,N_6791);
or U7048 (N_7048,N_6666,N_6696);
or U7049 (N_7049,N_6817,N_6606);
nor U7050 (N_7050,N_6674,N_6830);
nand U7051 (N_7051,N_6751,N_6777);
xor U7052 (N_7052,N_6604,N_6675);
nor U7053 (N_7053,N_6716,N_6651);
nor U7054 (N_7054,N_6616,N_6633);
nand U7055 (N_7055,N_6802,N_6700);
nor U7056 (N_7056,N_6744,N_6669);
and U7057 (N_7057,N_6801,N_6866);
nor U7058 (N_7058,N_6750,N_6678);
or U7059 (N_7059,N_6717,N_6800);
and U7060 (N_7060,N_6692,N_6843);
or U7061 (N_7061,N_6657,N_6830);
and U7062 (N_7062,N_6606,N_6754);
nand U7063 (N_7063,N_6798,N_6830);
xor U7064 (N_7064,N_6659,N_6772);
and U7065 (N_7065,N_6811,N_6843);
and U7066 (N_7066,N_6807,N_6704);
nand U7067 (N_7067,N_6859,N_6883);
or U7068 (N_7068,N_6854,N_6646);
nor U7069 (N_7069,N_6703,N_6631);
nor U7070 (N_7070,N_6648,N_6818);
nand U7071 (N_7071,N_6875,N_6660);
and U7072 (N_7072,N_6657,N_6602);
or U7073 (N_7073,N_6745,N_6661);
and U7074 (N_7074,N_6664,N_6778);
or U7075 (N_7075,N_6844,N_6642);
or U7076 (N_7076,N_6801,N_6857);
and U7077 (N_7077,N_6884,N_6643);
nand U7078 (N_7078,N_6675,N_6743);
and U7079 (N_7079,N_6784,N_6809);
xnor U7080 (N_7080,N_6838,N_6633);
or U7081 (N_7081,N_6888,N_6642);
and U7082 (N_7082,N_6825,N_6691);
or U7083 (N_7083,N_6694,N_6888);
xor U7084 (N_7084,N_6677,N_6744);
nand U7085 (N_7085,N_6649,N_6872);
or U7086 (N_7086,N_6898,N_6886);
or U7087 (N_7087,N_6602,N_6638);
xor U7088 (N_7088,N_6878,N_6611);
and U7089 (N_7089,N_6688,N_6743);
nor U7090 (N_7090,N_6604,N_6635);
xnor U7091 (N_7091,N_6797,N_6709);
nand U7092 (N_7092,N_6797,N_6762);
nor U7093 (N_7093,N_6823,N_6629);
xor U7094 (N_7094,N_6643,N_6835);
and U7095 (N_7095,N_6716,N_6702);
and U7096 (N_7096,N_6794,N_6717);
nand U7097 (N_7097,N_6776,N_6842);
nand U7098 (N_7098,N_6826,N_6624);
nand U7099 (N_7099,N_6684,N_6804);
xnor U7100 (N_7100,N_6796,N_6785);
nand U7101 (N_7101,N_6869,N_6892);
nand U7102 (N_7102,N_6797,N_6606);
nor U7103 (N_7103,N_6802,N_6799);
xnor U7104 (N_7104,N_6867,N_6856);
xnor U7105 (N_7105,N_6813,N_6849);
nor U7106 (N_7106,N_6718,N_6628);
nor U7107 (N_7107,N_6879,N_6697);
nand U7108 (N_7108,N_6694,N_6812);
nor U7109 (N_7109,N_6623,N_6709);
and U7110 (N_7110,N_6646,N_6865);
or U7111 (N_7111,N_6710,N_6741);
or U7112 (N_7112,N_6826,N_6741);
nand U7113 (N_7113,N_6841,N_6610);
nor U7114 (N_7114,N_6859,N_6709);
nand U7115 (N_7115,N_6880,N_6749);
or U7116 (N_7116,N_6888,N_6871);
nand U7117 (N_7117,N_6626,N_6831);
nor U7118 (N_7118,N_6671,N_6684);
xnor U7119 (N_7119,N_6895,N_6656);
xnor U7120 (N_7120,N_6634,N_6722);
nand U7121 (N_7121,N_6875,N_6815);
xor U7122 (N_7122,N_6699,N_6624);
and U7123 (N_7123,N_6687,N_6847);
nor U7124 (N_7124,N_6675,N_6605);
or U7125 (N_7125,N_6736,N_6835);
nor U7126 (N_7126,N_6739,N_6628);
nand U7127 (N_7127,N_6877,N_6658);
nand U7128 (N_7128,N_6894,N_6815);
or U7129 (N_7129,N_6861,N_6627);
or U7130 (N_7130,N_6762,N_6866);
nor U7131 (N_7131,N_6671,N_6735);
or U7132 (N_7132,N_6665,N_6709);
or U7133 (N_7133,N_6649,N_6776);
or U7134 (N_7134,N_6605,N_6854);
or U7135 (N_7135,N_6768,N_6600);
and U7136 (N_7136,N_6833,N_6608);
and U7137 (N_7137,N_6745,N_6832);
xnor U7138 (N_7138,N_6861,N_6746);
or U7139 (N_7139,N_6748,N_6815);
nand U7140 (N_7140,N_6667,N_6676);
nand U7141 (N_7141,N_6652,N_6673);
and U7142 (N_7142,N_6852,N_6849);
and U7143 (N_7143,N_6873,N_6891);
nand U7144 (N_7144,N_6762,N_6880);
nand U7145 (N_7145,N_6785,N_6831);
and U7146 (N_7146,N_6788,N_6742);
or U7147 (N_7147,N_6626,N_6632);
or U7148 (N_7148,N_6879,N_6725);
nand U7149 (N_7149,N_6814,N_6832);
xnor U7150 (N_7150,N_6706,N_6679);
nor U7151 (N_7151,N_6704,N_6763);
nor U7152 (N_7152,N_6635,N_6618);
and U7153 (N_7153,N_6809,N_6808);
or U7154 (N_7154,N_6811,N_6758);
nand U7155 (N_7155,N_6863,N_6650);
xnor U7156 (N_7156,N_6745,N_6698);
or U7157 (N_7157,N_6895,N_6852);
xnor U7158 (N_7158,N_6686,N_6644);
or U7159 (N_7159,N_6820,N_6604);
xnor U7160 (N_7160,N_6853,N_6767);
xor U7161 (N_7161,N_6766,N_6632);
nand U7162 (N_7162,N_6736,N_6665);
nor U7163 (N_7163,N_6845,N_6721);
nand U7164 (N_7164,N_6779,N_6860);
nand U7165 (N_7165,N_6647,N_6764);
nand U7166 (N_7166,N_6632,N_6827);
or U7167 (N_7167,N_6858,N_6607);
nand U7168 (N_7168,N_6894,N_6758);
nor U7169 (N_7169,N_6677,N_6621);
xnor U7170 (N_7170,N_6698,N_6840);
and U7171 (N_7171,N_6639,N_6894);
xor U7172 (N_7172,N_6806,N_6848);
nor U7173 (N_7173,N_6870,N_6676);
nor U7174 (N_7174,N_6656,N_6735);
or U7175 (N_7175,N_6773,N_6853);
nor U7176 (N_7176,N_6750,N_6849);
and U7177 (N_7177,N_6691,N_6627);
and U7178 (N_7178,N_6778,N_6642);
and U7179 (N_7179,N_6735,N_6699);
nor U7180 (N_7180,N_6678,N_6827);
xor U7181 (N_7181,N_6675,N_6760);
or U7182 (N_7182,N_6610,N_6701);
or U7183 (N_7183,N_6677,N_6866);
and U7184 (N_7184,N_6633,N_6614);
nor U7185 (N_7185,N_6702,N_6656);
nand U7186 (N_7186,N_6626,N_6740);
and U7187 (N_7187,N_6748,N_6897);
or U7188 (N_7188,N_6886,N_6749);
or U7189 (N_7189,N_6678,N_6674);
nor U7190 (N_7190,N_6630,N_6651);
nand U7191 (N_7191,N_6661,N_6873);
or U7192 (N_7192,N_6658,N_6829);
or U7193 (N_7193,N_6881,N_6687);
xor U7194 (N_7194,N_6667,N_6804);
and U7195 (N_7195,N_6675,N_6782);
xor U7196 (N_7196,N_6740,N_6698);
and U7197 (N_7197,N_6619,N_6786);
nor U7198 (N_7198,N_6853,N_6677);
nor U7199 (N_7199,N_6780,N_6813);
nand U7200 (N_7200,N_7097,N_7194);
nand U7201 (N_7201,N_7124,N_7080);
nand U7202 (N_7202,N_7193,N_7185);
and U7203 (N_7203,N_7164,N_7074);
or U7204 (N_7204,N_7147,N_7101);
xor U7205 (N_7205,N_7054,N_7116);
and U7206 (N_7206,N_7166,N_7069);
nor U7207 (N_7207,N_7184,N_7034);
xnor U7208 (N_7208,N_6931,N_6904);
or U7209 (N_7209,N_7198,N_7102);
and U7210 (N_7210,N_7149,N_7012);
or U7211 (N_7211,N_6959,N_7130);
or U7212 (N_7212,N_6970,N_6977);
or U7213 (N_7213,N_7025,N_7073);
xor U7214 (N_7214,N_6972,N_7044);
nand U7215 (N_7215,N_7160,N_7107);
and U7216 (N_7216,N_7146,N_6907);
and U7217 (N_7217,N_7026,N_7190);
and U7218 (N_7218,N_7145,N_7156);
and U7219 (N_7219,N_6963,N_7125);
xnor U7220 (N_7220,N_7072,N_7133);
xnor U7221 (N_7221,N_7121,N_6980);
and U7222 (N_7222,N_7091,N_6994);
nand U7223 (N_7223,N_7174,N_7047);
or U7224 (N_7224,N_7070,N_7129);
and U7225 (N_7225,N_7159,N_7151);
and U7226 (N_7226,N_6953,N_7056);
and U7227 (N_7227,N_7103,N_7171);
and U7228 (N_7228,N_6917,N_7168);
and U7229 (N_7229,N_7096,N_7017);
xnor U7230 (N_7230,N_6915,N_7144);
or U7231 (N_7231,N_7010,N_7098);
nand U7232 (N_7232,N_7083,N_7188);
or U7233 (N_7233,N_6903,N_7018);
and U7234 (N_7234,N_7094,N_7182);
or U7235 (N_7235,N_6909,N_7016);
or U7236 (N_7236,N_7055,N_6945);
and U7237 (N_7237,N_6993,N_7046);
nor U7238 (N_7238,N_6998,N_7162);
or U7239 (N_7239,N_6971,N_7021);
or U7240 (N_7240,N_7057,N_7082);
nor U7241 (N_7241,N_7170,N_7084);
and U7242 (N_7242,N_6938,N_7136);
xnor U7243 (N_7243,N_7095,N_6973);
or U7244 (N_7244,N_7173,N_7137);
nor U7245 (N_7245,N_6932,N_7120);
nor U7246 (N_7246,N_7195,N_7112);
and U7247 (N_7247,N_7126,N_6961);
or U7248 (N_7248,N_7150,N_7002);
and U7249 (N_7249,N_6954,N_6996);
nor U7250 (N_7250,N_6950,N_6900);
and U7251 (N_7251,N_6920,N_7053);
xor U7252 (N_7252,N_6955,N_7175);
or U7253 (N_7253,N_7143,N_7020);
or U7254 (N_7254,N_6951,N_6958);
nand U7255 (N_7255,N_6986,N_6901);
and U7256 (N_7256,N_7135,N_7163);
nor U7257 (N_7257,N_6935,N_7059);
and U7258 (N_7258,N_7060,N_6934);
or U7259 (N_7259,N_7148,N_7109);
nand U7260 (N_7260,N_7113,N_7140);
nand U7261 (N_7261,N_7092,N_6960);
and U7262 (N_7262,N_7177,N_6947);
nand U7263 (N_7263,N_6989,N_7030);
nand U7264 (N_7264,N_6914,N_7036);
xnor U7265 (N_7265,N_6956,N_6990);
xor U7266 (N_7266,N_7153,N_6979);
nand U7267 (N_7267,N_7139,N_6910);
and U7268 (N_7268,N_7192,N_6924);
xnor U7269 (N_7269,N_6982,N_7076);
or U7270 (N_7270,N_6952,N_7077);
and U7271 (N_7271,N_7038,N_7086);
or U7272 (N_7272,N_7052,N_7009);
nand U7273 (N_7273,N_7037,N_6921);
or U7274 (N_7274,N_7042,N_7049);
and U7275 (N_7275,N_7186,N_6930);
and U7276 (N_7276,N_7157,N_7063);
nand U7277 (N_7277,N_7006,N_6912);
xor U7278 (N_7278,N_6948,N_7003);
xor U7279 (N_7279,N_7031,N_7141);
or U7280 (N_7280,N_6957,N_7062);
nor U7281 (N_7281,N_6939,N_6926);
and U7282 (N_7282,N_7014,N_6902);
and U7283 (N_7283,N_7099,N_7169);
or U7284 (N_7284,N_6988,N_7104);
nand U7285 (N_7285,N_6927,N_7068);
nand U7286 (N_7286,N_7040,N_7011);
or U7287 (N_7287,N_6997,N_7050);
nand U7288 (N_7288,N_7079,N_6922);
or U7289 (N_7289,N_7075,N_7004);
nor U7290 (N_7290,N_7093,N_6919);
nor U7291 (N_7291,N_7114,N_7127);
xor U7292 (N_7292,N_7165,N_6936);
xor U7293 (N_7293,N_7111,N_6908);
nand U7294 (N_7294,N_6981,N_7088);
nor U7295 (N_7295,N_6995,N_7119);
or U7296 (N_7296,N_6946,N_7045);
nor U7297 (N_7297,N_7051,N_7176);
xnor U7298 (N_7298,N_7039,N_7172);
nand U7299 (N_7299,N_6964,N_6929);
xnor U7300 (N_7300,N_6911,N_6943);
nor U7301 (N_7301,N_6928,N_7001);
xnor U7302 (N_7302,N_6965,N_6969);
xnor U7303 (N_7303,N_7123,N_6905);
and U7304 (N_7304,N_7067,N_7032);
nand U7305 (N_7305,N_6987,N_7035);
nand U7306 (N_7306,N_7019,N_7013);
and U7307 (N_7307,N_6975,N_6913);
or U7308 (N_7308,N_6992,N_6978);
nand U7309 (N_7309,N_6974,N_7100);
or U7310 (N_7310,N_7064,N_7142);
nor U7311 (N_7311,N_7132,N_7007);
nor U7312 (N_7312,N_7008,N_7041);
nor U7313 (N_7313,N_7161,N_7183);
and U7314 (N_7314,N_7043,N_6999);
xor U7315 (N_7315,N_7110,N_6916);
nor U7316 (N_7316,N_7106,N_7134);
nor U7317 (N_7317,N_7048,N_7000);
and U7318 (N_7318,N_7118,N_7105);
xnor U7319 (N_7319,N_7167,N_6976);
or U7320 (N_7320,N_7196,N_7027);
and U7321 (N_7321,N_7115,N_7131);
and U7322 (N_7322,N_6937,N_7155);
nand U7323 (N_7323,N_7005,N_7033);
or U7324 (N_7324,N_7029,N_7181);
xnor U7325 (N_7325,N_6962,N_7078);
xnor U7326 (N_7326,N_7065,N_7061);
and U7327 (N_7327,N_7024,N_7089);
and U7328 (N_7328,N_7015,N_7087);
nand U7329 (N_7329,N_7138,N_7189);
nor U7330 (N_7330,N_7128,N_7152);
nor U7331 (N_7331,N_7197,N_7122);
xnor U7332 (N_7332,N_7066,N_7081);
xor U7333 (N_7333,N_6933,N_7028);
nand U7334 (N_7334,N_7158,N_6941);
or U7335 (N_7335,N_6949,N_7108);
or U7336 (N_7336,N_7023,N_6906);
xnor U7337 (N_7337,N_7058,N_7022);
or U7338 (N_7338,N_6925,N_6984);
or U7339 (N_7339,N_6985,N_7180);
and U7340 (N_7340,N_7117,N_6942);
nand U7341 (N_7341,N_6923,N_7187);
xnor U7342 (N_7342,N_7085,N_6918);
nand U7343 (N_7343,N_7090,N_7071);
or U7344 (N_7344,N_6944,N_7199);
and U7345 (N_7345,N_7154,N_6966);
or U7346 (N_7346,N_6991,N_6983);
nand U7347 (N_7347,N_6968,N_7191);
nand U7348 (N_7348,N_6940,N_6967);
xnor U7349 (N_7349,N_7179,N_7178);
xor U7350 (N_7350,N_6955,N_6954);
xor U7351 (N_7351,N_6939,N_6900);
and U7352 (N_7352,N_7199,N_6992);
xnor U7353 (N_7353,N_7096,N_6973);
and U7354 (N_7354,N_6955,N_6945);
nor U7355 (N_7355,N_7082,N_6951);
nor U7356 (N_7356,N_7130,N_7180);
or U7357 (N_7357,N_6991,N_7113);
and U7358 (N_7358,N_7078,N_6928);
or U7359 (N_7359,N_7025,N_7056);
nand U7360 (N_7360,N_7004,N_6947);
nand U7361 (N_7361,N_6969,N_7063);
or U7362 (N_7362,N_7047,N_6914);
or U7363 (N_7363,N_7024,N_6941);
nand U7364 (N_7364,N_7060,N_6952);
nand U7365 (N_7365,N_7076,N_7137);
or U7366 (N_7366,N_7182,N_7015);
and U7367 (N_7367,N_7197,N_6970);
xnor U7368 (N_7368,N_7129,N_7103);
or U7369 (N_7369,N_7137,N_6999);
nor U7370 (N_7370,N_7070,N_6974);
nand U7371 (N_7371,N_7135,N_6935);
or U7372 (N_7372,N_6967,N_7152);
or U7373 (N_7373,N_7134,N_7167);
and U7374 (N_7374,N_6997,N_7075);
xnor U7375 (N_7375,N_6951,N_7042);
nor U7376 (N_7376,N_6902,N_6924);
xnor U7377 (N_7377,N_7175,N_6934);
and U7378 (N_7378,N_7131,N_7140);
nor U7379 (N_7379,N_6973,N_7108);
or U7380 (N_7380,N_7127,N_6993);
or U7381 (N_7381,N_6994,N_7121);
xor U7382 (N_7382,N_6923,N_7140);
nand U7383 (N_7383,N_6993,N_7065);
nand U7384 (N_7384,N_6964,N_7003);
nand U7385 (N_7385,N_7016,N_6900);
and U7386 (N_7386,N_6970,N_7063);
nand U7387 (N_7387,N_6936,N_6921);
or U7388 (N_7388,N_6940,N_6911);
nand U7389 (N_7389,N_7019,N_7146);
and U7390 (N_7390,N_6911,N_6919);
nand U7391 (N_7391,N_7016,N_6954);
and U7392 (N_7392,N_6990,N_7160);
nand U7393 (N_7393,N_6910,N_7081);
and U7394 (N_7394,N_6976,N_7135);
nor U7395 (N_7395,N_7063,N_7101);
nand U7396 (N_7396,N_7027,N_6948);
or U7397 (N_7397,N_7099,N_7111);
nor U7398 (N_7398,N_7095,N_7168);
nor U7399 (N_7399,N_7173,N_7134);
nor U7400 (N_7400,N_7027,N_6918);
nand U7401 (N_7401,N_7040,N_7082);
nand U7402 (N_7402,N_7144,N_6979);
nand U7403 (N_7403,N_7170,N_7071);
or U7404 (N_7404,N_6990,N_7030);
nand U7405 (N_7405,N_6921,N_7031);
nand U7406 (N_7406,N_7064,N_7042);
nand U7407 (N_7407,N_7076,N_7195);
nor U7408 (N_7408,N_7125,N_7051);
or U7409 (N_7409,N_7072,N_6969);
nand U7410 (N_7410,N_6920,N_7151);
nand U7411 (N_7411,N_7067,N_6907);
and U7412 (N_7412,N_7112,N_6995);
nand U7413 (N_7413,N_6931,N_7057);
and U7414 (N_7414,N_7125,N_7161);
xor U7415 (N_7415,N_7093,N_7105);
xnor U7416 (N_7416,N_6964,N_7077);
and U7417 (N_7417,N_6990,N_7053);
xor U7418 (N_7418,N_7008,N_7015);
xor U7419 (N_7419,N_7170,N_7182);
or U7420 (N_7420,N_7119,N_6982);
and U7421 (N_7421,N_7074,N_6987);
or U7422 (N_7422,N_7049,N_7018);
nand U7423 (N_7423,N_7003,N_6919);
xor U7424 (N_7424,N_7047,N_7052);
xor U7425 (N_7425,N_6970,N_6962);
xnor U7426 (N_7426,N_7181,N_7191);
nor U7427 (N_7427,N_7060,N_6908);
nand U7428 (N_7428,N_6999,N_7090);
and U7429 (N_7429,N_7059,N_7027);
or U7430 (N_7430,N_7053,N_7073);
nor U7431 (N_7431,N_7096,N_6907);
xnor U7432 (N_7432,N_7031,N_7034);
and U7433 (N_7433,N_6902,N_7082);
xor U7434 (N_7434,N_7031,N_7196);
nand U7435 (N_7435,N_6988,N_7136);
xor U7436 (N_7436,N_6937,N_6974);
and U7437 (N_7437,N_7113,N_7129);
nand U7438 (N_7438,N_6912,N_7137);
nand U7439 (N_7439,N_6961,N_7082);
xnor U7440 (N_7440,N_6926,N_7008);
and U7441 (N_7441,N_7176,N_7048);
and U7442 (N_7442,N_7130,N_7025);
or U7443 (N_7443,N_7001,N_6948);
and U7444 (N_7444,N_7080,N_6915);
and U7445 (N_7445,N_7075,N_6951);
xor U7446 (N_7446,N_7199,N_7112);
nand U7447 (N_7447,N_6956,N_6968);
nor U7448 (N_7448,N_7044,N_6919);
nand U7449 (N_7449,N_6998,N_7022);
or U7450 (N_7450,N_6922,N_6990);
or U7451 (N_7451,N_6972,N_6955);
nand U7452 (N_7452,N_6998,N_7118);
xor U7453 (N_7453,N_6924,N_6934);
or U7454 (N_7454,N_7144,N_7053);
or U7455 (N_7455,N_7050,N_6974);
or U7456 (N_7456,N_6944,N_6994);
and U7457 (N_7457,N_7183,N_6904);
nor U7458 (N_7458,N_7025,N_7167);
nand U7459 (N_7459,N_7065,N_7171);
xor U7460 (N_7460,N_7085,N_7006);
and U7461 (N_7461,N_6926,N_7142);
and U7462 (N_7462,N_6973,N_7137);
or U7463 (N_7463,N_7071,N_7130);
nor U7464 (N_7464,N_6994,N_6968);
and U7465 (N_7465,N_7005,N_7159);
nand U7466 (N_7466,N_7053,N_6994);
nand U7467 (N_7467,N_6983,N_7182);
xor U7468 (N_7468,N_7129,N_7172);
xor U7469 (N_7469,N_6938,N_6945);
or U7470 (N_7470,N_7056,N_7090);
or U7471 (N_7471,N_7144,N_6973);
or U7472 (N_7472,N_6996,N_6935);
nand U7473 (N_7473,N_6908,N_7191);
nand U7474 (N_7474,N_7098,N_7020);
xor U7475 (N_7475,N_7022,N_6903);
nand U7476 (N_7476,N_6930,N_6908);
nand U7477 (N_7477,N_6993,N_7081);
nor U7478 (N_7478,N_7128,N_7085);
and U7479 (N_7479,N_7169,N_6967);
nand U7480 (N_7480,N_7075,N_7073);
xor U7481 (N_7481,N_7188,N_6946);
nor U7482 (N_7482,N_7163,N_6994);
or U7483 (N_7483,N_6944,N_6943);
nand U7484 (N_7484,N_6962,N_7012);
nor U7485 (N_7485,N_7156,N_6998);
nand U7486 (N_7486,N_7091,N_7009);
xnor U7487 (N_7487,N_6910,N_7095);
nor U7488 (N_7488,N_6906,N_7126);
or U7489 (N_7489,N_7002,N_7160);
or U7490 (N_7490,N_6990,N_6906);
and U7491 (N_7491,N_7082,N_6929);
or U7492 (N_7492,N_7160,N_7154);
or U7493 (N_7493,N_7094,N_7172);
xnor U7494 (N_7494,N_7095,N_6907);
nor U7495 (N_7495,N_7016,N_7197);
xor U7496 (N_7496,N_7018,N_7028);
or U7497 (N_7497,N_7070,N_7142);
and U7498 (N_7498,N_7011,N_7018);
or U7499 (N_7499,N_7172,N_7030);
nor U7500 (N_7500,N_7220,N_7432);
and U7501 (N_7501,N_7393,N_7307);
and U7502 (N_7502,N_7239,N_7446);
nor U7503 (N_7503,N_7406,N_7224);
nor U7504 (N_7504,N_7315,N_7421);
xor U7505 (N_7505,N_7440,N_7473);
xnor U7506 (N_7506,N_7385,N_7203);
nand U7507 (N_7507,N_7262,N_7227);
xor U7508 (N_7508,N_7388,N_7304);
and U7509 (N_7509,N_7368,N_7338);
and U7510 (N_7510,N_7383,N_7288);
xor U7511 (N_7511,N_7434,N_7350);
nand U7512 (N_7512,N_7223,N_7379);
nand U7513 (N_7513,N_7285,N_7492);
and U7514 (N_7514,N_7390,N_7452);
nand U7515 (N_7515,N_7218,N_7387);
and U7516 (N_7516,N_7327,N_7256);
xnor U7517 (N_7517,N_7330,N_7472);
nor U7518 (N_7518,N_7280,N_7303);
and U7519 (N_7519,N_7289,N_7284);
and U7520 (N_7520,N_7347,N_7210);
and U7521 (N_7521,N_7247,N_7437);
and U7522 (N_7522,N_7279,N_7323);
xnor U7523 (N_7523,N_7275,N_7415);
nor U7524 (N_7524,N_7345,N_7322);
nor U7525 (N_7525,N_7229,N_7399);
nand U7526 (N_7526,N_7252,N_7242);
nand U7527 (N_7527,N_7202,N_7445);
xor U7528 (N_7528,N_7470,N_7295);
nor U7529 (N_7529,N_7319,N_7422);
and U7530 (N_7530,N_7276,N_7353);
and U7531 (N_7531,N_7246,N_7266);
nor U7532 (N_7532,N_7412,N_7310);
nand U7533 (N_7533,N_7233,N_7346);
nor U7534 (N_7534,N_7357,N_7259);
nor U7535 (N_7535,N_7367,N_7403);
nand U7536 (N_7536,N_7290,N_7249);
nor U7537 (N_7537,N_7364,N_7389);
nor U7538 (N_7538,N_7483,N_7213);
and U7539 (N_7539,N_7419,N_7248);
xor U7540 (N_7540,N_7464,N_7365);
or U7541 (N_7541,N_7306,N_7463);
xnor U7542 (N_7542,N_7320,N_7298);
or U7543 (N_7543,N_7370,N_7458);
and U7544 (N_7544,N_7362,N_7337);
or U7545 (N_7545,N_7456,N_7352);
or U7546 (N_7546,N_7312,N_7297);
xor U7547 (N_7547,N_7386,N_7372);
xor U7548 (N_7548,N_7216,N_7438);
and U7549 (N_7549,N_7411,N_7225);
and U7550 (N_7550,N_7380,N_7324);
nand U7551 (N_7551,N_7444,N_7294);
nand U7552 (N_7552,N_7344,N_7495);
xnor U7553 (N_7553,N_7299,N_7436);
nor U7554 (N_7554,N_7207,N_7425);
nor U7555 (N_7555,N_7251,N_7237);
nand U7556 (N_7556,N_7355,N_7471);
nor U7557 (N_7557,N_7433,N_7486);
nor U7558 (N_7558,N_7427,N_7361);
and U7559 (N_7559,N_7359,N_7475);
and U7560 (N_7560,N_7351,N_7395);
nor U7561 (N_7561,N_7377,N_7429);
nor U7562 (N_7562,N_7499,N_7292);
nand U7563 (N_7563,N_7360,N_7270);
xnor U7564 (N_7564,N_7479,N_7494);
and U7565 (N_7565,N_7235,N_7363);
nand U7566 (N_7566,N_7455,N_7241);
and U7567 (N_7567,N_7405,N_7269);
nor U7568 (N_7568,N_7261,N_7480);
nand U7569 (N_7569,N_7443,N_7417);
nand U7570 (N_7570,N_7325,N_7414);
or U7571 (N_7571,N_7481,N_7407);
nor U7572 (N_7572,N_7451,N_7382);
or U7573 (N_7573,N_7243,N_7293);
nand U7574 (N_7574,N_7468,N_7410);
nand U7575 (N_7575,N_7373,N_7491);
xnor U7576 (N_7576,N_7428,N_7408);
nor U7577 (N_7577,N_7420,N_7281);
nor U7578 (N_7578,N_7374,N_7442);
nand U7579 (N_7579,N_7416,N_7371);
nor U7580 (N_7580,N_7469,N_7335);
or U7581 (N_7581,N_7485,N_7318);
xor U7582 (N_7582,N_7236,N_7231);
nor U7583 (N_7583,N_7300,N_7384);
nand U7584 (N_7584,N_7254,N_7448);
nor U7585 (N_7585,N_7212,N_7354);
nand U7586 (N_7586,N_7234,N_7206);
nand U7587 (N_7587,N_7278,N_7497);
or U7588 (N_7588,N_7466,N_7214);
and U7589 (N_7589,N_7305,N_7404);
and U7590 (N_7590,N_7204,N_7277);
and U7591 (N_7591,N_7267,N_7439);
nor U7592 (N_7592,N_7426,N_7488);
xor U7593 (N_7593,N_7490,N_7447);
nor U7594 (N_7594,N_7316,N_7311);
or U7595 (N_7595,N_7487,N_7402);
and U7596 (N_7596,N_7313,N_7205);
xnor U7597 (N_7597,N_7423,N_7282);
and U7598 (N_7598,N_7339,N_7308);
or U7599 (N_7599,N_7232,N_7476);
nor U7600 (N_7600,N_7394,N_7333);
nand U7601 (N_7601,N_7268,N_7465);
xnor U7602 (N_7602,N_7484,N_7302);
and U7603 (N_7603,N_7331,N_7461);
nand U7604 (N_7604,N_7271,N_7453);
and U7605 (N_7605,N_7200,N_7400);
xor U7606 (N_7606,N_7392,N_7441);
nor U7607 (N_7607,N_7498,N_7431);
nand U7608 (N_7608,N_7343,N_7334);
or U7609 (N_7609,N_7454,N_7260);
nor U7610 (N_7610,N_7215,N_7369);
and U7611 (N_7611,N_7238,N_7228);
or U7612 (N_7612,N_7450,N_7250);
and U7613 (N_7613,N_7460,N_7349);
nor U7614 (N_7614,N_7240,N_7258);
xor U7615 (N_7615,N_7366,N_7273);
xor U7616 (N_7616,N_7301,N_7321);
or U7617 (N_7617,N_7348,N_7462);
xnor U7618 (N_7618,N_7221,N_7244);
or U7619 (N_7619,N_7457,N_7459);
nor U7620 (N_7620,N_7317,N_7332);
nand U7621 (N_7621,N_7219,N_7493);
nor U7622 (N_7622,N_7477,N_7376);
xnor U7623 (N_7623,N_7217,N_7341);
nor U7624 (N_7624,N_7245,N_7253);
and U7625 (N_7625,N_7329,N_7264);
and U7626 (N_7626,N_7378,N_7274);
or U7627 (N_7627,N_7375,N_7342);
or U7628 (N_7628,N_7263,N_7340);
nor U7629 (N_7629,N_7467,N_7449);
xor U7630 (N_7630,N_7209,N_7496);
xnor U7631 (N_7631,N_7309,N_7226);
or U7632 (N_7632,N_7474,N_7489);
and U7633 (N_7633,N_7409,N_7230);
and U7634 (N_7634,N_7358,N_7222);
nand U7635 (N_7635,N_7381,N_7283);
xnor U7636 (N_7636,N_7287,N_7255);
or U7637 (N_7637,N_7418,N_7272);
or U7638 (N_7638,N_7257,N_7356);
or U7639 (N_7639,N_7424,N_7435);
nand U7640 (N_7640,N_7396,N_7336);
nand U7641 (N_7641,N_7314,N_7413);
nor U7642 (N_7642,N_7430,N_7478);
or U7643 (N_7643,N_7286,N_7201);
and U7644 (N_7644,N_7398,N_7397);
or U7645 (N_7645,N_7326,N_7328);
nand U7646 (N_7646,N_7482,N_7391);
or U7647 (N_7647,N_7291,N_7401);
nor U7648 (N_7648,N_7211,N_7296);
and U7649 (N_7649,N_7208,N_7265);
nand U7650 (N_7650,N_7202,N_7446);
xnor U7651 (N_7651,N_7469,N_7331);
and U7652 (N_7652,N_7238,N_7498);
or U7653 (N_7653,N_7474,N_7438);
nand U7654 (N_7654,N_7382,N_7398);
xor U7655 (N_7655,N_7430,N_7358);
or U7656 (N_7656,N_7402,N_7236);
or U7657 (N_7657,N_7363,N_7439);
nand U7658 (N_7658,N_7365,N_7381);
nor U7659 (N_7659,N_7201,N_7345);
nor U7660 (N_7660,N_7378,N_7424);
xnor U7661 (N_7661,N_7363,N_7278);
nor U7662 (N_7662,N_7234,N_7372);
and U7663 (N_7663,N_7249,N_7401);
xnor U7664 (N_7664,N_7307,N_7313);
and U7665 (N_7665,N_7262,N_7292);
nand U7666 (N_7666,N_7224,N_7443);
and U7667 (N_7667,N_7453,N_7230);
xnor U7668 (N_7668,N_7474,N_7230);
and U7669 (N_7669,N_7475,N_7458);
nor U7670 (N_7670,N_7360,N_7328);
and U7671 (N_7671,N_7492,N_7478);
xor U7672 (N_7672,N_7218,N_7259);
nand U7673 (N_7673,N_7424,N_7391);
and U7674 (N_7674,N_7398,N_7414);
nand U7675 (N_7675,N_7264,N_7393);
nand U7676 (N_7676,N_7294,N_7200);
nand U7677 (N_7677,N_7377,N_7440);
nor U7678 (N_7678,N_7420,N_7304);
or U7679 (N_7679,N_7283,N_7465);
and U7680 (N_7680,N_7481,N_7200);
nand U7681 (N_7681,N_7303,N_7353);
and U7682 (N_7682,N_7208,N_7273);
and U7683 (N_7683,N_7333,N_7379);
xor U7684 (N_7684,N_7248,N_7202);
nor U7685 (N_7685,N_7470,N_7253);
nor U7686 (N_7686,N_7378,N_7213);
nor U7687 (N_7687,N_7255,N_7302);
nor U7688 (N_7688,N_7471,N_7240);
or U7689 (N_7689,N_7318,N_7334);
nand U7690 (N_7690,N_7320,N_7463);
and U7691 (N_7691,N_7381,N_7215);
xnor U7692 (N_7692,N_7320,N_7339);
nand U7693 (N_7693,N_7285,N_7243);
and U7694 (N_7694,N_7231,N_7298);
or U7695 (N_7695,N_7356,N_7291);
or U7696 (N_7696,N_7200,N_7446);
and U7697 (N_7697,N_7391,N_7272);
nand U7698 (N_7698,N_7271,N_7385);
nor U7699 (N_7699,N_7444,N_7343);
and U7700 (N_7700,N_7357,N_7394);
or U7701 (N_7701,N_7209,N_7315);
or U7702 (N_7702,N_7491,N_7498);
or U7703 (N_7703,N_7349,N_7264);
and U7704 (N_7704,N_7334,N_7352);
or U7705 (N_7705,N_7403,N_7373);
and U7706 (N_7706,N_7278,N_7251);
and U7707 (N_7707,N_7417,N_7260);
xnor U7708 (N_7708,N_7331,N_7496);
nor U7709 (N_7709,N_7329,N_7284);
and U7710 (N_7710,N_7383,N_7243);
and U7711 (N_7711,N_7459,N_7258);
or U7712 (N_7712,N_7395,N_7428);
nor U7713 (N_7713,N_7301,N_7233);
and U7714 (N_7714,N_7276,N_7313);
nand U7715 (N_7715,N_7209,N_7239);
nor U7716 (N_7716,N_7460,N_7254);
or U7717 (N_7717,N_7467,N_7463);
or U7718 (N_7718,N_7256,N_7447);
and U7719 (N_7719,N_7326,N_7449);
and U7720 (N_7720,N_7452,N_7438);
nand U7721 (N_7721,N_7461,N_7240);
nor U7722 (N_7722,N_7464,N_7347);
xnor U7723 (N_7723,N_7260,N_7368);
nor U7724 (N_7724,N_7492,N_7388);
xor U7725 (N_7725,N_7360,N_7493);
nor U7726 (N_7726,N_7479,N_7261);
xor U7727 (N_7727,N_7210,N_7373);
and U7728 (N_7728,N_7363,N_7373);
or U7729 (N_7729,N_7241,N_7364);
nor U7730 (N_7730,N_7362,N_7220);
and U7731 (N_7731,N_7278,N_7422);
xnor U7732 (N_7732,N_7369,N_7211);
xor U7733 (N_7733,N_7463,N_7277);
and U7734 (N_7734,N_7261,N_7469);
nor U7735 (N_7735,N_7201,N_7233);
nand U7736 (N_7736,N_7356,N_7417);
nand U7737 (N_7737,N_7434,N_7402);
and U7738 (N_7738,N_7367,N_7317);
xor U7739 (N_7739,N_7302,N_7259);
nor U7740 (N_7740,N_7365,N_7243);
xnor U7741 (N_7741,N_7434,N_7360);
xnor U7742 (N_7742,N_7410,N_7320);
xnor U7743 (N_7743,N_7223,N_7451);
nand U7744 (N_7744,N_7419,N_7477);
or U7745 (N_7745,N_7252,N_7221);
xnor U7746 (N_7746,N_7263,N_7429);
and U7747 (N_7747,N_7403,N_7394);
xnor U7748 (N_7748,N_7236,N_7396);
nor U7749 (N_7749,N_7365,N_7346);
nand U7750 (N_7750,N_7478,N_7374);
nand U7751 (N_7751,N_7318,N_7340);
and U7752 (N_7752,N_7296,N_7375);
xnor U7753 (N_7753,N_7334,N_7342);
xor U7754 (N_7754,N_7401,N_7455);
nand U7755 (N_7755,N_7386,N_7281);
or U7756 (N_7756,N_7318,N_7427);
or U7757 (N_7757,N_7207,N_7325);
nor U7758 (N_7758,N_7460,N_7278);
or U7759 (N_7759,N_7218,N_7293);
and U7760 (N_7760,N_7361,N_7385);
xnor U7761 (N_7761,N_7292,N_7436);
and U7762 (N_7762,N_7259,N_7398);
or U7763 (N_7763,N_7312,N_7368);
nor U7764 (N_7764,N_7218,N_7267);
and U7765 (N_7765,N_7280,N_7355);
xnor U7766 (N_7766,N_7211,N_7312);
nor U7767 (N_7767,N_7230,N_7227);
xnor U7768 (N_7768,N_7278,N_7381);
nand U7769 (N_7769,N_7338,N_7351);
and U7770 (N_7770,N_7289,N_7499);
nor U7771 (N_7771,N_7320,N_7394);
nand U7772 (N_7772,N_7438,N_7416);
xnor U7773 (N_7773,N_7216,N_7483);
nand U7774 (N_7774,N_7275,N_7333);
or U7775 (N_7775,N_7498,N_7322);
xnor U7776 (N_7776,N_7292,N_7377);
or U7777 (N_7777,N_7219,N_7385);
and U7778 (N_7778,N_7458,N_7448);
or U7779 (N_7779,N_7455,N_7378);
nand U7780 (N_7780,N_7480,N_7225);
and U7781 (N_7781,N_7204,N_7205);
and U7782 (N_7782,N_7283,N_7210);
and U7783 (N_7783,N_7463,N_7384);
or U7784 (N_7784,N_7473,N_7381);
nor U7785 (N_7785,N_7436,N_7461);
or U7786 (N_7786,N_7446,N_7374);
xnor U7787 (N_7787,N_7366,N_7276);
nor U7788 (N_7788,N_7453,N_7423);
or U7789 (N_7789,N_7201,N_7239);
nand U7790 (N_7790,N_7499,N_7341);
and U7791 (N_7791,N_7386,N_7371);
nand U7792 (N_7792,N_7453,N_7364);
or U7793 (N_7793,N_7444,N_7457);
xnor U7794 (N_7794,N_7246,N_7272);
nand U7795 (N_7795,N_7340,N_7406);
nor U7796 (N_7796,N_7429,N_7278);
and U7797 (N_7797,N_7459,N_7391);
xor U7798 (N_7798,N_7385,N_7278);
or U7799 (N_7799,N_7481,N_7439);
or U7800 (N_7800,N_7524,N_7572);
or U7801 (N_7801,N_7639,N_7570);
and U7802 (N_7802,N_7681,N_7569);
and U7803 (N_7803,N_7561,N_7558);
xnor U7804 (N_7804,N_7757,N_7529);
xor U7805 (N_7805,N_7533,N_7598);
and U7806 (N_7806,N_7535,N_7698);
xnor U7807 (N_7807,N_7732,N_7623);
and U7808 (N_7808,N_7611,N_7505);
xor U7809 (N_7809,N_7607,N_7734);
nor U7810 (N_7810,N_7509,N_7768);
nor U7811 (N_7811,N_7714,N_7543);
and U7812 (N_7812,N_7599,N_7584);
nor U7813 (N_7813,N_7673,N_7617);
or U7814 (N_7814,N_7510,N_7513);
and U7815 (N_7815,N_7526,N_7578);
nand U7816 (N_7816,N_7713,N_7666);
xnor U7817 (N_7817,N_7756,N_7538);
nor U7818 (N_7818,N_7554,N_7679);
xnor U7819 (N_7819,N_7655,N_7548);
nand U7820 (N_7820,N_7641,N_7691);
and U7821 (N_7821,N_7575,N_7706);
and U7822 (N_7822,N_7622,N_7615);
nand U7823 (N_7823,N_7557,N_7542);
nor U7824 (N_7824,N_7507,N_7752);
or U7825 (N_7825,N_7614,N_7724);
nor U7826 (N_7826,N_7736,N_7596);
nor U7827 (N_7827,N_7503,N_7587);
nand U7828 (N_7828,N_7571,N_7669);
nand U7829 (N_7829,N_7523,N_7667);
nand U7830 (N_7830,N_7780,N_7580);
xnor U7831 (N_7831,N_7647,N_7630);
nand U7832 (N_7832,N_7668,N_7773);
or U7833 (N_7833,N_7789,N_7586);
nand U7834 (N_7834,N_7795,N_7699);
and U7835 (N_7835,N_7775,N_7602);
or U7836 (N_7836,N_7762,N_7717);
nand U7837 (N_7837,N_7688,N_7730);
or U7838 (N_7838,N_7771,N_7733);
and U7839 (N_7839,N_7595,N_7729);
nor U7840 (N_7840,N_7566,N_7727);
nor U7841 (N_7841,N_7612,N_7700);
or U7842 (N_7842,N_7606,N_7740);
nor U7843 (N_7843,N_7627,N_7755);
nor U7844 (N_7844,N_7689,N_7520);
nand U7845 (N_7845,N_7545,N_7674);
nand U7846 (N_7846,N_7620,N_7675);
and U7847 (N_7847,N_7551,N_7697);
and U7848 (N_7848,N_7646,N_7785);
and U7849 (N_7849,N_7648,N_7796);
nor U7850 (N_7850,N_7565,N_7650);
xor U7851 (N_7851,N_7657,N_7659);
nor U7852 (N_7852,N_7685,N_7704);
and U7853 (N_7853,N_7741,N_7760);
nand U7854 (N_7854,N_7683,N_7726);
or U7855 (N_7855,N_7553,N_7577);
and U7856 (N_7856,N_7568,N_7703);
nor U7857 (N_7857,N_7608,N_7731);
or U7858 (N_7858,N_7636,N_7672);
nor U7859 (N_7859,N_7552,N_7573);
nor U7860 (N_7860,N_7787,N_7506);
and U7861 (N_7861,N_7754,N_7634);
or U7862 (N_7862,N_7522,N_7531);
xor U7863 (N_7863,N_7582,N_7585);
xor U7864 (N_7864,N_7626,N_7676);
nor U7865 (N_7865,N_7799,N_7514);
or U7866 (N_7866,N_7723,N_7656);
nor U7867 (N_7867,N_7564,N_7663);
xor U7868 (N_7868,N_7654,N_7652);
nor U7869 (N_7869,N_7784,N_7778);
and U7870 (N_7870,N_7750,N_7525);
xnor U7871 (N_7871,N_7791,N_7766);
or U7872 (N_7872,N_7537,N_7753);
xor U7873 (N_7873,N_7701,N_7748);
nand U7874 (N_7874,N_7738,N_7696);
nand U7875 (N_7875,N_7677,N_7519);
or U7876 (N_7876,N_7769,N_7643);
nor U7877 (N_7877,N_7761,N_7720);
nand U7878 (N_7878,N_7546,N_7781);
and U7879 (N_7879,N_7516,N_7550);
nor U7880 (N_7880,N_7604,N_7770);
xor U7881 (N_7881,N_7504,N_7702);
nor U7882 (N_7882,N_7593,N_7744);
nand U7883 (N_7883,N_7635,N_7745);
nor U7884 (N_7884,N_7767,N_7782);
nor U7885 (N_7885,N_7678,N_7665);
or U7886 (N_7886,N_7690,N_7613);
nor U7887 (N_7887,N_7621,N_7722);
or U7888 (N_7888,N_7544,N_7649);
nor U7889 (N_7889,N_7605,N_7783);
and U7890 (N_7890,N_7747,N_7528);
or U7891 (N_7891,N_7707,N_7776);
and U7892 (N_7892,N_7628,N_7786);
xnor U7893 (N_7893,N_7680,N_7549);
nor U7894 (N_7894,N_7695,N_7772);
nor U7895 (N_7895,N_7594,N_7798);
nand U7896 (N_7896,N_7728,N_7642);
and U7897 (N_7897,N_7590,N_7779);
nand U7898 (N_7898,N_7721,N_7682);
or U7899 (N_7899,N_7739,N_7500);
nor U7900 (N_7900,N_7579,N_7793);
or U7901 (N_7901,N_7746,N_7711);
or U7902 (N_7902,N_7742,N_7653);
nand U7903 (N_7903,N_7518,N_7644);
xor U7904 (N_7904,N_7664,N_7616);
nor U7905 (N_7905,N_7631,N_7794);
or U7906 (N_7906,N_7719,N_7600);
and U7907 (N_7907,N_7591,N_7661);
and U7908 (N_7908,N_7556,N_7512);
nand U7909 (N_7909,N_7624,N_7662);
and U7910 (N_7910,N_7709,N_7708);
xor U7911 (N_7911,N_7532,N_7694);
xnor U7912 (N_7912,N_7547,N_7692);
nand U7913 (N_7913,N_7511,N_7592);
or U7914 (N_7914,N_7777,N_7581);
xor U7915 (N_7915,N_7640,N_7797);
nor U7916 (N_7916,N_7637,N_7588);
nor U7917 (N_7917,N_7687,N_7671);
xor U7918 (N_7918,N_7765,N_7743);
nand U7919 (N_7919,N_7788,N_7758);
nor U7920 (N_7920,N_7763,N_7660);
and U7921 (N_7921,N_7560,N_7693);
nor U7922 (N_7922,N_7521,N_7710);
or U7923 (N_7923,N_7684,N_7563);
xnor U7924 (N_7924,N_7574,N_7629);
and U7925 (N_7925,N_7759,N_7737);
and U7926 (N_7926,N_7619,N_7589);
nor U7927 (N_7927,N_7517,N_7534);
nand U7928 (N_7928,N_7601,N_7638);
xnor U7929 (N_7929,N_7749,N_7718);
xnor U7930 (N_7930,N_7536,N_7576);
nand U7931 (N_7931,N_7632,N_7764);
or U7932 (N_7932,N_7715,N_7610);
and U7933 (N_7933,N_7645,N_7597);
or U7934 (N_7934,N_7792,N_7625);
and U7935 (N_7935,N_7559,N_7530);
and U7936 (N_7936,N_7515,N_7502);
or U7937 (N_7937,N_7751,N_7501);
nand U7938 (N_7938,N_7541,N_7735);
xor U7939 (N_7939,N_7539,N_7705);
xnor U7940 (N_7940,N_7725,N_7583);
or U7941 (N_7941,N_7567,N_7508);
and U7942 (N_7942,N_7618,N_7658);
or U7943 (N_7943,N_7670,N_7774);
xnor U7944 (N_7944,N_7527,N_7603);
nand U7945 (N_7945,N_7555,N_7790);
nor U7946 (N_7946,N_7651,N_7712);
nor U7947 (N_7947,N_7686,N_7540);
or U7948 (N_7948,N_7716,N_7633);
and U7949 (N_7949,N_7562,N_7609);
and U7950 (N_7950,N_7644,N_7531);
or U7951 (N_7951,N_7782,N_7554);
or U7952 (N_7952,N_7600,N_7573);
nor U7953 (N_7953,N_7504,N_7552);
nor U7954 (N_7954,N_7640,N_7695);
nor U7955 (N_7955,N_7793,N_7745);
nand U7956 (N_7956,N_7538,N_7534);
or U7957 (N_7957,N_7571,N_7506);
xor U7958 (N_7958,N_7671,N_7607);
or U7959 (N_7959,N_7686,N_7688);
or U7960 (N_7960,N_7622,N_7754);
and U7961 (N_7961,N_7761,N_7717);
nor U7962 (N_7962,N_7655,N_7773);
nand U7963 (N_7963,N_7719,N_7598);
nand U7964 (N_7964,N_7710,N_7795);
nand U7965 (N_7965,N_7722,N_7539);
and U7966 (N_7966,N_7701,N_7640);
nand U7967 (N_7967,N_7547,N_7798);
xor U7968 (N_7968,N_7686,N_7530);
nor U7969 (N_7969,N_7765,N_7702);
nand U7970 (N_7970,N_7573,N_7786);
and U7971 (N_7971,N_7758,N_7522);
or U7972 (N_7972,N_7588,N_7765);
nand U7973 (N_7973,N_7668,N_7682);
nand U7974 (N_7974,N_7535,N_7584);
xnor U7975 (N_7975,N_7749,N_7660);
nand U7976 (N_7976,N_7501,N_7585);
nand U7977 (N_7977,N_7786,N_7519);
or U7978 (N_7978,N_7726,N_7704);
xor U7979 (N_7979,N_7742,N_7798);
and U7980 (N_7980,N_7595,N_7525);
nand U7981 (N_7981,N_7725,N_7754);
nor U7982 (N_7982,N_7669,N_7677);
and U7983 (N_7983,N_7544,N_7748);
nor U7984 (N_7984,N_7519,N_7599);
nor U7985 (N_7985,N_7638,N_7656);
nor U7986 (N_7986,N_7745,N_7740);
nor U7987 (N_7987,N_7785,N_7555);
or U7988 (N_7988,N_7706,N_7781);
nor U7989 (N_7989,N_7759,N_7622);
nor U7990 (N_7990,N_7537,N_7599);
or U7991 (N_7991,N_7519,N_7587);
and U7992 (N_7992,N_7696,N_7737);
nand U7993 (N_7993,N_7793,N_7665);
nor U7994 (N_7994,N_7789,N_7737);
and U7995 (N_7995,N_7760,N_7544);
or U7996 (N_7996,N_7723,N_7746);
xnor U7997 (N_7997,N_7784,N_7775);
and U7998 (N_7998,N_7629,N_7550);
nand U7999 (N_7999,N_7689,N_7780);
xnor U8000 (N_8000,N_7776,N_7716);
xnor U8001 (N_8001,N_7508,N_7624);
nor U8002 (N_8002,N_7769,N_7736);
or U8003 (N_8003,N_7505,N_7664);
and U8004 (N_8004,N_7547,N_7527);
nor U8005 (N_8005,N_7574,N_7791);
xnor U8006 (N_8006,N_7738,N_7695);
nand U8007 (N_8007,N_7560,N_7644);
xnor U8008 (N_8008,N_7594,N_7505);
xnor U8009 (N_8009,N_7780,N_7721);
and U8010 (N_8010,N_7710,N_7721);
nand U8011 (N_8011,N_7707,N_7628);
xor U8012 (N_8012,N_7728,N_7547);
nand U8013 (N_8013,N_7715,N_7652);
and U8014 (N_8014,N_7519,N_7578);
nor U8015 (N_8015,N_7775,N_7794);
nor U8016 (N_8016,N_7628,N_7683);
and U8017 (N_8017,N_7662,N_7720);
nand U8018 (N_8018,N_7540,N_7797);
and U8019 (N_8019,N_7656,N_7501);
nand U8020 (N_8020,N_7559,N_7698);
nor U8021 (N_8021,N_7647,N_7669);
nand U8022 (N_8022,N_7557,N_7624);
or U8023 (N_8023,N_7536,N_7521);
or U8024 (N_8024,N_7684,N_7581);
xor U8025 (N_8025,N_7711,N_7772);
xor U8026 (N_8026,N_7691,N_7563);
or U8027 (N_8027,N_7647,N_7542);
xor U8028 (N_8028,N_7749,N_7799);
and U8029 (N_8029,N_7737,N_7534);
nand U8030 (N_8030,N_7799,N_7732);
or U8031 (N_8031,N_7587,N_7525);
xor U8032 (N_8032,N_7574,N_7692);
xnor U8033 (N_8033,N_7675,N_7600);
nand U8034 (N_8034,N_7767,N_7676);
xnor U8035 (N_8035,N_7594,N_7746);
nand U8036 (N_8036,N_7553,N_7568);
and U8037 (N_8037,N_7642,N_7708);
xnor U8038 (N_8038,N_7526,N_7625);
nor U8039 (N_8039,N_7624,N_7764);
or U8040 (N_8040,N_7632,N_7702);
nand U8041 (N_8041,N_7710,N_7702);
nand U8042 (N_8042,N_7639,N_7576);
and U8043 (N_8043,N_7731,N_7743);
or U8044 (N_8044,N_7555,N_7593);
or U8045 (N_8045,N_7798,N_7584);
nand U8046 (N_8046,N_7718,N_7584);
nand U8047 (N_8047,N_7526,N_7706);
xor U8048 (N_8048,N_7644,N_7596);
or U8049 (N_8049,N_7560,N_7572);
nor U8050 (N_8050,N_7535,N_7503);
xor U8051 (N_8051,N_7662,N_7705);
nand U8052 (N_8052,N_7720,N_7661);
and U8053 (N_8053,N_7671,N_7519);
or U8054 (N_8054,N_7772,N_7586);
xnor U8055 (N_8055,N_7563,N_7722);
or U8056 (N_8056,N_7536,N_7592);
nand U8057 (N_8057,N_7580,N_7630);
xnor U8058 (N_8058,N_7647,N_7777);
or U8059 (N_8059,N_7559,N_7611);
or U8060 (N_8060,N_7746,N_7724);
and U8061 (N_8061,N_7797,N_7735);
and U8062 (N_8062,N_7623,N_7671);
and U8063 (N_8063,N_7673,N_7720);
or U8064 (N_8064,N_7614,N_7601);
nor U8065 (N_8065,N_7630,N_7556);
and U8066 (N_8066,N_7692,N_7713);
xor U8067 (N_8067,N_7677,N_7601);
nor U8068 (N_8068,N_7582,N_7595);
and U8069 (N_8069,N_7542,N_7552);
or U8070 (N_8070,N_7678,N_7674);
nor U8071 (N_8071,N_7514,N_7711);
and U8072 (N_8072,N_7668,N_7554);
nand U8073 (N_8073,N_7591,N_7506);
and U8074 (N_8074,N_7747,N_7703);
nand U8075 (N_8075,N_7559,N_7799);
nor U8076 (N_8076,N_7545,N_7526);
nand U8077 (N_8077,N_7540,N_7550);
and U8078 (N_8078,N_7719,N_7575);
or U8079 (N_8079,N_7783,N_7616);
nand U8080 (N_8080,N_7534,N_7565);
xor U8081 (N_8081,N_7610,N_7789);
nor U8082 (N_8082,N_7553,N_7569);
or U8083 (N_8083,N_7595,N_7631);
nor U8084 (N_8084,N_7550,N_7567);
or U8085 (N_8085,N_7689,N_7762);
nand U8086 (N_8086,N_7590,N_7658);
nand U8087 (N_8087,N_7669,N_7599);
nand U8088 (N_8088,N_7782,N_7747);
xnor U8089 (N_8089,N_7516,N_7787);
and U8090 (N_8090,N_7723,N_7735);
or U8091 (N_8091,N_7554,N_7541);
nand U8092 (N_8092,N_7683,N_7600);
xnor U8093 (N_8093,N_7591,N_7713);
nand U8094 (N_8094,N_7744,N_7759);
nor U8095 (N_8095,N_7791,N_7673);
and U8096 (N_8096,N_7699,N_7580);
nor U8097 (N_8097,N_7537,N_7548);
and U8098 (N_8098,N_7673,N_7639);
nand U8099 (N_8099,N_7616,N_7673);
nand U8100 (N_8100,N_7997,N_8050);
nor U8101 (N_8101,N_7943,N_7800);
nor U8102 (N_8102,N_7861,N_8045);
nand U8103 (N_8103,N_8080,N_7944);
or U8104 (N_8104,N_7959,N_8078);
nor U8105 (N_8105,N_8085,N_8028);
and U8106 (N_8106,N_7852,N_7870);
and U8107 (N_8107,N_8011,N_7864);
nor U8108 (N_8108,N_7805,N_7847);
nand U8109 (N_8109,N_7890,N_7947);
or U8110 (N_8110,N_8067,N_7949);
nand U8111 (N_8111,N_7950,N_7830);
nand U8112 (N_8112,N_8072,N_7993);
nor U8113 (N_8113,N_7863,N_7908);
or U8114 (N_8114,N_7801,N_8084);
nand U8115 (N_8115,N_7874,N_7853);
and U8116 (N_8116,N_7882,N_7922);
nand U8117 (N_8117,N_8030,N_7906);
or U8118 (N_8118,N_7992,N_7854);
nor U8119 (N_8119,N_7967,N_8086);
nor U8120 (N_8120,N_7820,N_7904);
nand U8121 (N_8121,N_8026,N_8032);
xnor U8122 (N_8122,N_8059,N_7851);
nor U8123 (N_8123,N_7955,N_7807);
nor U8124 (N_8124,N_7828,N_8062);
xor U8125 (N_8125,N_8002,N_7822);
nand U8126 (N_8126,N_7860,N_7891);
nor U8127 (N_8127,N_8015,N_7975);
and U8128 (N_8128,N_7920,N_7946);
and U8129 (N_8129,N_8018,N_8000);
xor U8130 (N_8130,N_7948,N_7990);
nand U8131 (N_8131,N_8037,N_8031);
or U8132 (N_8132,N_7982,N_7827);
nor U8133 (N_8133,N_7895,N_8040);
and U8134 (N_8134,N_7921,N_7818);
nor U8135 (N_8135,N_8025,N_7829);
nor U8136 (N_8136,N_8035,N_7928);
nor U8137 (N_8137,N_7978,N_8066);
nand U8138 (N_8138,N_8090,N_7925);
or U8139 (N_8139,N_7994,N_7848);
or U8140 (N_8140,N_7979,N_7867);
nor U8141 (N_8141,N_7932,N_8082);
nor U8142 (N_8142,N_7842,N_8024);
xor U8143 (N_8143,N_7998,N_7927);
nor U8144 (N_8144,N_8083,N_7869);
or U8145 (N_8145,N_8075,N_7883);
and U8146 (N_8146,N_7880,N_7831);
and U8147 (N_8147,N_7862,N_7840);
xnor U8148 (N_8148,N_7878,N_8048);
nand U8149 (N_8149,N_8047,N_7802);
nand U8150 (N_8150,N_7907,N_7939);
xnor U8151 (N_8151,N_8088,N_7887);
xnor U8152 (N_8152,N_7892,N_8053);
xnor U8153 (N_8153,N_8034,N_7938);
and U8154 (N_8154,N_7855,N_7876);
xnor U8155 (N_8155,N_8017,N_8043);
or U8156 (N_8156,N_8003,N_7817);
nor U8157 (N_8157,N_7912,N_8089);
nand U8158 (N_8158,N_7889,N_7875);
nand U8159 (N_8159,N_8007,N_7850);
and U8160 (N_8160,N_7957,N_7872);
or U8161 (N_8161,N_7812,N_8019);
or U8162 (N_8162,N_8004,N_7885);
or U8163 (N_8163,N_7806,N_7923);
or U8164 (N_8164,N_8014,N_7886);
xor U8165 (N_8165,N_7859,N_7811);
xor U8166 (N_8166,N_8074,N_7819);
and U8167 (N_8167,N_7898,N_8052);
or U8168 (N_8168,N_7896,N_7962);
and U8169 (N_8169,N_8038,N_8060);
and U8170 (N_8170,N_7824,N_7914);
or U8171 (N_8171,N_7841,N_7846);
nor U8172 (N_8172,N_7910,N_7970);
xor U8173 (N_8173,N_7804,N_7952);
nor U8174 (N_8174,N_7972,N_7971);
or U8175 (N_8175,N_7984,N_8013);
and U8176 (N_8176,N_8012,N_7953);
nand U8177 (N_8177,N_7905,N_8022);
and U8178 (N_8178,N_7836,N_7936);
nor U8179 (N_8179,N_7868,N_7940);
xor U8180 (N_8180,N_7826,N_7999);
and U8181 (N_8181,N_7873,N_8095);
xnor U8182 (N_8182,N_7963,N_7816);
xor U8183 (N_8183,N_7931,N_7930);
or U8184 (N_8184,N_7969,N_7900);
or U8185 (N_8185,N_7991,N_7866);
nor U8186 (N_8186,N_8029,N_7894);
nand U8187 (N_8187,N_7808,N_7986);
and U8188 (N_8188,N_7919,N_7958);
xnor U8189 (N_8189,N_8077,N_7917);
nand U8190 (N_8190,N_7835,N_7985);
nor U8191 (N_8191,N_8016,N_7966);
and U8192 (N_8192,N_7834,N_7954);
and U8193 (N_8193,N_7995,N_7964);
xnor U8194 (N_8194,N_7934,N_8008);
or U8195 (N_8195,N_7942,N_7911);
or U8196 (N_8196,N_8044,N_7929);
nand U8197 (N_8197,N_8070,N_8051);
nand U8198 (N_8198,N_8079,N_7832);
nor U8199 (N_8199,N_7961,N_8021);
xor U8200 (N_8200,N_7987,N_7937);
nor U8201 (N_8201,N_8068,N_7844);
nand U8202 (N_8202,N_8027,N_8058);
nor U8203 (N_8203,N_8097,N_8005);
nor U8204 (N_8204,N_7918,N_7996);
xor U8205 (N_8205,N_7951,N_8009);
and U8206 (N_8206,N_8093,N_8055);
nor U8207 (N_8207,N_7803,N_7915);
nor U8208 (N_8208,N_7976,N_7973);
xor U8209 (N_8209,N_7843,N_8010);
or U8210 (N_8210,N_8023,N_8073);
nor U8211 (N_8211,N_7857,N_8054);
and U8212 (N_8212,N_7988,N_8063);
and U8213 (N_8213,N_8061,N_7881);
and U8214 (N_8214,N_8069,N_7945);
nand U8215 (N_8215,N_8094,N_8020);
nor U8216 (N_8216,N_8033,N_8098);
or U8217 (N_8217,N_8099,N_8092);
and U8218 (N_8218,N_7879,N_7933);
nor U8219 (N_8219,N_7809,N_7814);
or U8220 (N_8220,N_7849,N_7815);
and U8221 (N_8221,N_8064,N_7965);
and U8222 (N_8222,N_8087,N_8065);
xnor U8223 (N_8223,N_7899,N_8056);
or U8224 (N_8224,N_7821,N_7893);
xnor U8225 (N_8225,N_7902,N_7838);
or U8226 (N_8226,N_7926,N_7871);
nor U8227 (N_8227,N_7833,N_7825);
and U8228 (N_8228,N_7924,N_8049);
and U8229 (N_8229,N_7913,N_7903);
and U8230 (N_8230,N_8036,N_7845);
or U8231 (N_8231,N_7968,N_8071);
nor U8232 (N_8232,N_8081,N_7823);
and U8233 (N_8233,N_8091,N_7981);
nand U8234 (N_8234,N_7897,N_7956);
xnor U8235 (N_8235,N_7983,N_8041);
xnor U8236 (N_8236,N_7813,N_8039);
or U8237 (N_8237,N_7974,N_7865);
xnor U8238 (N_8238,N_7989,N_7909);
nand U8239 (N_8239,N_8057,N_7888);
nand U8240 (N_8240,N_7839,N_8006);
xor U8241 (N_8241,N_7901,N_8042);
nor U8242 (N_8242,N_7858,N_7856);
and U8243 (N_8243,N_7980,N_7884);
xor U8244 (N_8244,N_7810,N_7916);
nor U8245 (N_8245,N_8096,N_8001);
and U8246 (N_8246,N_7941,N_7877);
or U8247 (N_8247,N_7960,N_7977);
or U8248 (N_8248,N_8076,N_7935);
nor U8249 (N_8249,N_7837,N_8046);
xnor U8250 (N_8250,N_8022,N_7831);
nand U8251 (N_8251,N_7998,N_8024);
nand U8252 (N_8252,N_7911,N_8075);
or U8253 (N_8253,N_7828,N_7865);
nor U8254 (N_8254,N_7951,N_7967);
or U8255 (N_8255,N_7971,N_7821);
nor U8256 (N_8256,N_8003,N_7809);
nand U8257 (N_8257,N_7954,N_8090);
nor U8258 (N_8258,N_8020,N_8055);
nand U8259 (N_8259,N_7935,N_7909);
or U8260 (N_8260,N_7954,N_7965);
and U8261 (N_8261,N_8089,N_7978);
xnor U8262 (N_8262,N_7867,N_7852);
nor U8263 (N_8263,N_7867,N_7911);
xnor U8264 (N_8264,N_7925,N_8035);
or U8265 (N_8265,N_8061,N_8024);
nand U8266 (N_8266,N_8069,N_8074);
or U8267 (N_8267,N_7811,N_7834);
nor U8268 (N_8268,N_8037,N_8041);
xnor U8269 (N_8269,N_7957,N_8000);
nand U8270 (N_8270,N_8076,N_7838);
xnor U8271 (N_8271,N_8066,N_7827);
nor U8272 (N_8272,N_7878,N_8035);
xnor U8273 (N_8273,N_7894,N_7922);
xor U8274 (N_8274,N_7849,N_7964);
or U8275 (N_8275,N_7835,N_7990);
nand U8276 (N_8276,N_7817,N_8022);
nand U8277 (N_8277,N_8039,N_8040);
and U8278 (N_8278,N_7835,N_7828);
xnor U8279 (N_8279,N_7804,N_8093);
and U8280 (N_8280,N_7829,N_7860);
xnor U8281 (N_8281,N_7875,N_8086);
xnor U8282 (N_8282,N_7829,N_7883);
or U8283 (N_8283,N_7978,N_7854);
nand U8284 (N_8284,N_8056,N_7926);
xnor U8285 (N_8285,N_7850,N_7804);
and U8286 (N_8286,N_7945,N_7938);
xor U8287 (N_8287,N_7909,N_7899);
nor U8288 (N_8288,N_7821,N_8031);
nand U8289 (N_8289,N_7957,N_7951);
xnor U8290 (N_8290,N_7994,N_7999);
and U8291 (N_8291,N_7892,N_7899);
xnor U8292 (N_8292,N_7840,N_8022);
or U8293 (N_8293,N_7917,N_7935);
and U8294 (N_8294,N_8051,N_7823);
xnor U8295 (N_8295,N_7861,N_7819);
and U8296 (N_8296,N_7980,N_8095);
and U8297 (N_8297,N_8070,N_7998);
and U8298 (N_8298,N_7904,N_7843);
xnor U8299 (N_8299,N_7914,N_7823);
or U8300 (N_8300,N_7851,N_8067);
xnor U8301 (N_8301,N_8094,N_7851);
or U8302 (N_8302,N_7805,N_7947);
nand U8303 (N_8303,N_7871,N_7873);
nor U8304 (N_8304,N_7969,N_7920);
or U8305 (N_8305,N_7981,N_7822);
nor U8306 (N_8306,N_7969,N_7814);
nand U8307 (N_8307,N_7945,N_8017);
or U8308 (N_8308,N_7840,N_8050);
nor U8309 (N_8309,N_7841,N_7944);
and U8310 (N_8310,N_7879,N_7919);
nor U8311 (N_8311,N_7976,N_7883);
and U8312 (N_8312,N_7954,N_7827);
nor U8313 (N_8313,N_7848,N_7821);
nor U8314 (N_8314,N_8075,N_7810);
or U8315 (N_8315,N_8084,N_7908);
nand U8316 (N_8316,N_7966,N_7802);
or U8317 (N_8317,N_7889,N_7941);
nand U8318 (N_8318,N_8026,N_7980);
and U8319 (N_8319,N_8036,N_7972);
xnor U8320 (N_8320,N_7973,N_7978);
nor U8321 (N_8321,N_7800,N_7920);
nor U8322 (N_8322,N_7944,N_7901);
xor U8323 (N_8323,N_7804,N_8021);
nor U8324 (N_8324,N_7822,N_7848);
or U8325 (N_8325,N_7887,N_8031);
xor U8326 (N_8326,N_8018,N_8039);
nor U8327 (N_8327,N_8018,N_7836);
or U8328 (N_8328,N_7943,N_7985);
nor U8329 (N_8329,N_7965,N_7855);
or U8330 (N_8330,N_8077,N_8058);
nand U8331 (N_8331,N_8049,N_8028);
nor U8332 (N_8332,N_7836,N_7808);
nand U8333 (N_8333,N_8032,N_7867);
xnor U8334 (N_8334,N_7895,N_7842);
nor U8335 (N_8335,N_8005,N_7961);
nand U8336 (N_8336,N_7869,N_7910);
or U8337 (N_8337,N_7974,N_7827);
nor U8338 (N_8338,N_7960,N_7860);
xor U8339 (N_8339,N_7970,N_7984);
xnor U8340 (N_8340,N_7875,N_8000);
or U8341 (N_8341,N_7860,N_7989);
xnor U8342 (N_8342,N_7943,N_7817);
or U8343 (N_8343,N_8020,N_8059);
xor U8344 (N_8344,N_7818,N_7918);
xor U8345 (N_8345,N_7811,N_7990);
and U8346 (N_8346,N_7916,N_8034);
nor U8347 (N_8347,N_7963,N_7812);
nor U8348 (N_8348,N_8029,N_7909);
nand U8349 (N_8349,N_7843,N_7818);
and U8350 (N_8350,N_7837,N_7990);
or U8351 (N_8351,N_7989,N_8037);
xor U8352 (N_8352,N_8035,N_7931);
xnor U8353 (N_8353,N_8039,N_7838);
and U8354 (N_8354,N_8045,N_7929);
or U8355 (N_8355,N_7813,N_7854);
or U8356 (N_8356,N_7844,N_8033);
or U8357 (N_8357,N_7814,N_8078);
xor U8358 (N_8358,N_7858,N_8020);
or U8359 (N_8359,N_7891,N_7812);
nor U8360 (N_8360,N_8043,N_8003);
nor U8361 (N_8361,N_8070,N_7901);
and U8362 (N_8362,N_8043,N_7968);
or U8363 (N_8363,N_7918,N_8083);
nand U8364 (N_8364,N_7830,N_7981);
xnor U8365 (N_8365,N_8023,N_8040);
and U8366 (N_8366,N_8042,N_7921);
and U8367 (N_8367,N_7870,N_7885);
nor U8368 (N_8368,N_7982,N_8042);
or U8369 (N_8369,N_8042,N_7920);
nand U8370 (N_8370,N_7983,N_7901);
and U8371 (N_8371,N_8085,N_7938);
nand U8372 (N_8372,N_8006,N_7809);
or U8373 (N_8373,N_7943,N_8085);
nor U8374 (N_8374,N_7964,N_7911);
or U8375 (N_8375,N_7910,N_8078);
or U8376 (N_8376,N_8070,N_7909);
nand U8377 (N_8377,N_8083,N_8088);
nand U8378 (N_8378,N_7897,N_7860);
and U8379 (N_8379,N_8004,N_7896);
xnor U8380 (N_8380,N_8079,N_7856);
xor U8381 (N_8381,N_7832,N_8084);
xnor U8382 (N_8382,N_7962,N_7815);
or U8383 (N_8383,N_7811,N_7916);
nor U8384 (N_8384,N_7921,N_7939);
nor U8385 (N_8385,N_7923,N_7817);
xor U8386 (N_8386,N_7947,N_7976);
nor U8387 (N_8387,N_7812,N_7924);
nand U8388 (N_8388,N_7934,N_8091);
and U8389 (N_8389,N_7875,N_7876);
and U8390 (N_8390,N_8005,N_8004);
nand U8391 (N_8391,N_7964,N_7965);
nand U8392 (N_8392,N_7815,N_8073);
and U8393 (N_8393,N_7989,N_8086);
nand U8394 (N_8394,N_7943,N_7994);
and U8395 (N_8395,N_7930,N_7818);
xnor U8396 (N_8396,N_7841,N_7892);
xor U8397 (N_8397,N_7836,N_7883);
and U8398 (N_8398,N_7822,N_8001);
nand U8399 (N_8399,N_7970,N_7994);
nand U8400 (N_8400,N_8267,N_8326);
xnor U8401 (N_8401,N_8145,N_8140);
xor U8402 (N_8402,N_8307,N_8252);
nor U8403 (N_8403,N_8177,N_8121);
xnor U8404 (N_8404,N_8189,N_8208);
nand U8405 (N_8405,N_8325,N_8146);
nor U8406 (N_8406,N_8188,N_8175);
and U8407 (N_8407,N_8352,N_8336);
nand U8408 (N_8408,N_8180,N_8260);
nand U8409 (N_8409,N_8291,N_8297);
and U8410 (N_8410,N_8216,N_8360);
nor U8411 (N_8411,N_8295,N_8112);
xor U8412 (N_8412,N_8251,N_8293);
xor U8413 (N_8413,N_8356,N_8378);
nand U8414 (N_8414,N_8332,N_8113);
nand U8415 (N_8415,N_8205,N_8284);
or U8416 (N_8416,N_8320,N_8393);
xor U8417 (N_8417,N_8160,N_8290);
nand U8418 (N_8418,N_8289,N_8167);
xnor U8419 (N_8419,N_8234,N_8117);
nor U8420 (N_8420,N_8330,N_8166);
or U8421 (N_8421,N_8328,N_8294);
or U8422 (N_8422,N_8346,N_8310);
or U8423 (N_8423,N_8181,N_8190);
nand U8424 (N_8424,N_8338,N_8244);
and U8425 (N_8425,N_8229,N_8220);
and U8426 (N_8426,N_8334,N_8395);
nand U8427 (N_8427,N_8182,N_8271);
xnor U8428 (N_8428,N_8381,N_8256);
nor U8429 (N_8429,N_8217,N_8374);
xnor U8430 (N_8430,N_8351,N_8298);
and U8431 (N_8431,N_8344,N_8274);
or U8432 (N_8432,N_8169,N_8357);
nand U8433 (N_8433,N_8387,N_8191);
xor U8434 (N_8434,N_8253,N_8266);
nand U8435 (N_8435,N_8211,N_8394);
and U8436 (N_8436,N_8315,N_8200);
and U8437 (N_8437,N_8236,N_8218);
xor U8438 (N_8438,N_8142,N_8309);
and U8439 (N_8439,N_8154,N_8390);
nand U8440 (N_8440,N_8138,N_8255);
nand U8441 (N_8441,N_8209,N_8385);
nand U8442 (N_8442,N_8304,N_8179);
nand U8443 (N_8443,N_8238,N_8322);
and U8444 (N_8444,N_8354,N_8375);
nor U8445 (N_8445,N_8345,N_8116);
nor U8446 (N_8446,N_8366,N_8141);
nand U8447 (N_8447,N_8300,N_8231);
nand U8448 (N_8448,N_8161,N_8162);
nand U8449 (N_8449,N_8153,N_8157);
xnor U8450 (N_8450,N_8143,N_8319);
xor U8451 (N_8451,N_8163,N_8224);
nand U8452 (N_8452,N_8386,N_8353);
and U8453 (N_8453,N_8324,N_8119);
xor U8454 (N_8454,N_8221,N_8235);
xnor U8455 (N_8455,N_8249,N_8342);
xor U8456 (N_8456,N_8135,N_8268);
xnor U8457 (N_8457,N_8228,N_8118);
xnor U8458 (N_8458,N_8213,N_8199);
xor U8459 (N_8459,N_8323,N_8137);
nand U8460 (N_8460,N_8287,N_8275);
or U8461 (N_8461,N_8281,N_8292);
nor U8462 (N_8462,N_8184,N_8120);
or U8463 (N_8463,N_8302,N_8288);
or U8464 (N_8464,N_8369,N_8358);
and U8465 (N_8465,N_8373,N_8149);
xor U8466 (N_8466,N_8331,N_8214);
and U8467 (N_8467,N_8222,N_8176);
or U8468 (N_8468,N_8318,N_8258);
and U8469 (N_8469,N_8193,N_8259);
xor U8470 (N_8470,N_8202,N_8399);
nor U8471 (N_8471,N_8283,N_8359);
and U8472 (N_8472,N_8278,N_8276);
nor U8473 (N_8473,N_8367,N_8349);
xnor U8474 (N_8474,N_8102,N_8333);
or U8475 (N_8475,N_8183,N_8243);
xnor U8476 (N_8476,N_8206,N_8311);
nand U8477 (N_8477,N_8391,N_8261);
nand U8478 (N_8478,N_8159,N_8272);
nor U8479 (N_8479,N_8262,N_8109);
nand U8480 (N_8480,N_8370,N_8170);
nand U8481 (N_8481,N_8158,N_8398);
nor U8482 (N_8482,N_8144,N_8316);
and U8483 (N_8483,N_8148,N_8123);
or U8484 (N_8484,N_8111,N_8246);
nor U8485 (N_8485,N_8263,N_8348);
or U8486 (N_8486,N_8172,N_8329);
and U8487 (N_8487,N_8174,N_8233);
and U8488 (N_8488,N_8377,N_8350);
or U8489 (N_8489,N_8270,N_8128);
or U8490 (N_8490,N_8203,N_8339);
nor U8491 (N_8491,N_8337,N_8282);
or U8492 (N_8492,N_8132,N_8107);
nand U8493 (N_8493,N_8226,N_8365);
or U8494 (N_8494,N_8204,N_8372);
or U8495 (N_8495,N_8382,N_8237);
and U8496 (N_8496,N_8397,N_8273);
nor U8497 (N_8497,N_8156,N_8227);
or U8498 (N_8498,N_8240,N_8198);
nand U8499 (N_8499,N_8389,N_8219);
nand U8500 (N_8500,N_8306,N_8379);
xor U8501 (N_8501,N_8305,N_8388);
or U8502 (N_8502,N_8101,N_8313);
nor U8503 (N_8503,N_8127,N_8106);
or U8504 (N_8504,N_8103,N_8384);
or U8505 (N_8505,N_8317,N_8364);
nor U8506 (N_8506,N_8242,N_8257);
and U8507 (N_8507,N_8327,N_8165);
xor U8508 (N_8508,N_8363,N_8343);
or U8509 (N_8509,N_8114,N_8321);
xnor U8510 (N_8510,N_8303,N_8314);
xnor U8511 (N_8511,N_8368,N_8269);
nand U8512 (N_8512,N_8392,N_8215);
xor U8513 (N_8513,N_8280,N_8164);
and U8514 (N_8514,N_8230,N_8340);
nand U8515 (N_8515,N_8301,N_8104);
and U8516 (N_8516,N_8134,N_8241);
xor U8517 (N_8517,N_8299,N_8129);
or U8518 (N_8518,N_8210,N_8115);
and U8519 (N_8519,N_8131,N_8185);
nand U8520 (N_8520,N_8396,N_8187);
or U8521 (N_8521,N_8245,N_8296);
nor U8522 (N_8522,N_8380,N_8248);
xnor U8523 (N_8523,N_8122,N_8133);
xor U8524 (N_8524,N_8347,N_8376);
and U8525 (N_8525,N_8383,N_8105);
xor U8526 (N_8526,N_8225,N_8151);
xor U8527 (N_8527,N_8194,N_8335);
nand U8528 (N_8528,N_8341,N_8250);
xor U8529 (N_8529,N_8136,N_8239);
nor U8530 (N_8530,N_8308,N_8150);
and U8531 (N_8531,N_8355,N_8223);
nor U8532 (N_8532,N_8286,N_8247);
nand U8533 (N_8533,N_8212,N_8173);
and U8534 (N_8534,N_8197,N_8124);
or U8535 (N_8535,N_8201,N_8147);
and U8536 (N_8536,N_8168,N_8195);
nand U8537 (N_8537,N_8362,N_8361);
and U8538 (N_8538,N_8186,N_8108);
and U8539 (N_8539,N_8265,N_8207);
nand U8540 (N_8540,N_8110,N_8254);
or U8541 (N_8541,N_8155,N_8371);
or U8542 (N_8542,N_8126,N_8130);
nand U8543 (N_8543,N_8277,N_8100);
and U8544 (N_8544,N_8312,N_8285);
or U8545 (N_8545,N_8178,N_8196);
xnor U8546 (N_8546,N_8264,N_8192);
and U8547 (N_8547,N_8139,N_8171);
nand U8548 (N_8548,N_8125,N_8152);
nand U8549 (N_8549,N_8279,N_8232);
or U8550 (N_8550,N_8379,N_8369);
nor U8551 (N_8551,N_8266,N_8396);
nand U8552 (N_8552,N_8161,N_8116);
and U8553 (N_8553,N_8298,N_8273);
nor U8554 (N_8554,N_8288,N_8360);
and U8555 (N_8555,N_8273,N_8108);
nor U8556 (N_8556,N_8117,N_8317);
nor U8557 (N_8557,N_8282,N_8252);
or U8558 (N_8558,N_8279,N_8247);
or U8559 (N_8559,N_8158,N_8165);
or U8560 (N_8560,N_8387,N_8274);
xnor U8561 (N_8561,N_8134,N_8150);
xor U8562 (N_8562,N_8357,N_8170);
or U8563 (N_8563,N_8355,N_8202);
and U8564 (N_8564,N_8396,N_8278);
nand U8565 (N_8565,N_8361,N_8284);
nor U8566 (N_8566,N_8269,N_8225);
and U8567 (N_8567,N_8298,N_8342);
xor U8568 (N_8568,N_8244,N_8253);
nor U8569 (N_8569,N_8369,N_8378);
nor U8570 (N_8570,N_8363,N_8329);
xor U8571 (N_8571,N_8265,N_8164);
or U8572 (N_8572,N_8110,N_8245);
nor U8573 (N_8573,N_8294,N_8136);
nor U8574 (N_8574,N_8130,N_8152);
nor U8575 (N_8575,N_8160,N_8317);
or U8576 (N_8576,N_8357,N_8210);
and U8577 (N_8577,N_8162,N_8318);
nor U8578 (N_8578,N_8138,N_8157);
or U8579 (N_8579,N_8131,N_8201);
and U8580 (N_8580,N_8373,N_8313);
or U8581 (N_8581,N_8311,N_8338);
or U8582 (N_8582,N_8100,N_8117);
or U8583 (N_8583,N_8114,N_8335);
nand U8584 (N_8584,N_8159,N_8113);
nand U8585 (N_8585,N_8359,N_8272);
or U8586 (N_8586,N_8255,N_8125);
nor U8587 (N_8587,N_8283,N_8275);
nand U8588 (N_8588,N_8378,N_8349);
xor U8589 (N_8589,N_8341,N_8275);
nand U8590 (N_8590,N_8360,N_8148);
xnor U8591 (N_8591,N_8223,N_8206);
nor U8592 (N_8592,N_8147,N_8177);
or U8593 (N_8593,N_8304,N_8217);
and U8594 (N_8594,N_8126,N_8362);
nor U8595 (N_8595,N_8195,N_8218);
nor U8596 (N_8596,N_8179,N_8218);
nand U8597 (N_8597,N_8168,N_8358);
xor U8598 (N_8598,N_8267,N_8292);
and U8599 (N_8599,N_8320,N_8396);
and U8600 (N_8600,N_8149,N_8250);
or U8601 (N_8601,N_8161,N_8321);
xnor U8602 (N_8602,N_8116,N_8341);
nor U8603 (N_8603,N_8188,N_8157);
nand U8604 (N_8604,N_8195,N_8358);
xnor U8605 (N_8605,N_8306,N_8149);
nand U8606 (N_8606,N_8144,N_8341);
nand U8607 (N_8607,N_8151,N_8251);
or U8608 (N_8608,N_8399,N_8355);
xor U8609 (N_8609,N_8262,N_8357);
or U8610 (N_8610,N_8253,N_8170);
or U8611 (N_8611,N_8191,N_8383);
nand U8612 (N_8612,N_8130,N_8238);
and U8613 (N_8613,N_8354,N_8146);
or U8614 (N_8614,N_8387,N_8208);
and U8615 (N_8615,N_8242,N_8156);
nand U8616 (N_8616,N_8100,N_8184);
or U8617 (N_8617,N_8331,N_8175);
nand U8618 (N_8618,N_8171,N_8314);
nor U8619 (N_8619,N_8111,N_8363);
nor U8620 (N_8620,N_8124,N_8287);
and U8621 (N_8621,N_8385,N_8197);
and U8622 (N_8622,N_8315,N_8280);
nor U8623 (N_8623,N_8112,N_8225);
and U8624 (N_8624,N_8301,N_8166);
or U8625 (N_8625,N_8180,N_8124);
xor U8626 (N_8626,N_8395,N_8233);
xor U8627 (N_8627,N_8246,N_8174);
or U8628 (N_8628,N_8153,N_8285);
or U8629 (N_8629,N_8186,N_8373);
nor U8630 (N_8630,N_8185,N_8165);
nor U8631 (N_8631,N_8354,N_8309);
and U8632 (N_8632,N_8118,N_8358);
or U8633 (N_8633,N_8155,N_8305);
nand U8634 (N_8634,N_8397,N_8379);
xnor U8635 (N_8635,N_8274,N_8351);
xor U8636 (N_8636,N_8314,N_8218);
and U8637 (N_8637,N_8178,N_8131);
xnor U8638 (N_8638,N_8127,N_8253);
and U8639 (N_8639,N_8274,N_8125);
and U8640 (N_8640,N_8351,N_8197);
xor U8641 (N_8641,N_8129,N_8174);
and U8642 (N_8642,N_8169,N_8266);
and U8643 (N_8643,N_8115,N_8391);
nand U8644 (N_8644,N_8340,N_8311);
nor U8645 (N_8645,N_8344,N_8338);
and U8646 (N_8646,N_8352,N_8295);
nand U8647 (N_8647,N_8154,N_8269);
or U8648 (N_8648,N_8214,N_8370);
nand U8649 (N_8649,N_8128,N_8310);
and U8650 (N_8650,N_8346,N_8174);
or U8651 (N_8651,N_8214,N_8383);
and U8652 (N_8652,N_8189,N_8236);
xor U8653 (N_8653,N_8243,N_8362);
nand U8654 (N_8654,N_8294,N_8119);
or U8655 (N_8655,N_8167,N_8151);
and U8656 (N_8656,N_8139,N_8297);
nand U8657 (N_8657,N_8203,N_8263);
and U8658 (N_8658,N_8257,N_8189);
or U8659 (N_8659,N_8124,N_8245);
and U8660 (N_8660,N_8372,N_8369);
nor U8661 (N_8661,N_8177,N_8318);
xnor U8662 (N_8662,N_8304,N_8139);
nor U8663 (N_8663,N_8165,N_8355);
and U8664 (N_8664,N_8280,N_8367);
xor U8665 (N_8665,N_8167,N_8229);
or U8666 (N_8666,N_8147,N_8274);
nand U8667 (N_8667,N_8388,N_8374);
nor U8668 (N_8668,N_8375,N_8170);
nor U8669 (N_8669,N_8219,N_8225);
or U8670 (N_8670,N_8355,N_8185);
nor U8671 (N_8671,N_8205,N_8324);
nand U8672 (N_8672,N_8120,N_8223);
xor U8673 (N_8673,N_8359,N_8390);
nand U8674 (N_8674,N_8119,N_8187);
and U8675 (N_8675,N_8386,N_8276);
nor U8676 (N_8676,N_8397,N_8212);
and U8677 (N_8677,N_8364,N_8299);
or U8678 (N_8678,N_8292,N_8198);
and U8679 (N_8679,N_8235,N_8289);
xnor U8680 (N_8680,N_8364,N_8235);
nor U8681 (N_8681,N_8129,N_8339);
xnor U8682 (N_8682,N_8145,N_8167);
or U8683 (N_8683,N_8341,N_8211);
xor U8684 (N_8684,N_8142,N_8195);
xnor U8685 (N_8685,N_8199,N_8190);
xnor U8686 (N_8686,N_8258,N_8280);
xnor U8687 (N_8687,N_8149,N_8122);
xnor U8688 (N_8688,N_8263,N_8236);
nor U8689 (N_8689,N_8137,N_8138);
xor U8690 (N_8690,N_8182,N_8384);
nand U8691 (N_8691,N_8298,N_8195);
nand U8692 (N_8692,N_8328,N_8353);
and U8693 (N_8693,N_8313,N_8260);
nor U8694 (N_8694,N_8373,N_8325);
and U8695 (N_8695,N_8330,N_8217);
or U8696 (N_8696,N_8392,N_8289);
or U8697 (N_8697,N_8104,N_8153);
or U8698 (N_8698,N_8136,N_8338);
and U8699 (N_8699,N_8265,N_8341);
nand U8700 (N_8700,N_8681,N_8684);
nand U8701 (N_8701,N_8643,N_8579);
nand U8702 (N_8702,N_8473,N_8452);
or U8703 (N_8703,N_8433,N_8449);
nand U8704 (N_8704,N_8488,N_8647);
nor U8705 (N_8705,N_8622,N_8442);
xor U8706 (N_8706,N_8561,N_8650);
and U8707 (N_8707,N_8629,N_8554);
or U8708 (N_8708,N_8674,N_8479);
or U8709 (N_8709,N_8631,N_8691);
nor U8710 (N_8710,N_8645,N_8608);
xnor U8711 (N_8711,N_8653,N_8489);
nor U8712 (N_8712,N_8617,N_8616);
and U8713 (N_8713,N_8601,N_8538);
and U8714 (N_8714,N_8472,N_8576);
or U8715 (N_8715,N_8414,N_8676);
xor U8716 (N_8716,N_8470,N_8527);
and U8717 (N_8717,N_8604,N_8408);
or U8718 (N_8718,N_8533,N_8420);
nor U8719 (N_8719,N_8458,N_8666);
or U8720 (N_8720,N_8531,N_8422);
xnor U8721 (N_8721,N_8583,N_8438);
or U8722 (N_8722,N_8459,N_8501);
nand U8723 (N_8723,N_8564,N_8520);
nand U8724 (N_8724,N_8588,N_8614);
xnor U8725 (N_8725,N_8627,N_8405);
and U8726 (N_8726,N_8566,N_8518);
nor U8727 (N_8727,N_8569,N_8672);
or U8728 (N_8728,N_8580,N_8648);
or U8729 (N_8729,N_8620,N_8652);
xnor U8730 (N_8730,N_8659,N_8439);
or U8731 (N_8731,N_8547,N_8665);
or U8732 (N_8732,N_8613,N_8661);
nand U8733 (N_8733,N_8656,N_8611);
xor U8734 (N_8734,N_8628,N_8453);
nor U8735 (N_8735,N_8693,N_8594);
or U8736 (N_8736,N_8475,N_8544);
xnor U8737 (N_8737,N_8492,N_8609);
xnor U8738 (N_8738,N_8536,N_8448);
nor U8739 (N_8739,N_8556,N_8486);
or U8740 (N_8740,N_8465,N_8549);
or U8741 (N_8741,N_8424,N_8502);
or U8742 (N_8742,N_8657,N_8655);
xnor U8743 (N_8743,N_8532,N_8410);
xor U8744 (N_8744,N_8673,N_8572);
and U8745 (N_8745,N_8568,N_8619);
and U8746 (N_8746,N_8560,N_8679);
or U8747 (N_8747,N_8494,N_8495);
or U8748 (N_8748,N_8567,N_8491);
nor U8749 (N_8749,N_8625,N_8641);
and U8750 (N_8750,N_8697,N_8678);
and U8751 (N_8751,N_8537,N_8668);
xor U8752 (N_8752,N_8654,N_8523);
xnor U8753 (N_8753,N_8670,N_8419);
and U8754 (N_8754,N_8680,N_8637);
nand U8755 (N_8755,N_8407,N_8496);
nor U8756 (N_8756,N_8635,N_8460);
xnor U8757 (N_8757,N_8677,N_8513);
or U8758 (N_8758,N_8529,N_8558);
or U8759 (N_8759,N_8667,N_8546);
nor U8760 (N_8760,N_8401,N_8437);
xor U8761 (N_8761,N_8582,N_8514);
or U8762 (N_8762,N_8418,N_8624);
xor U8763 (N_8763,N_8688,N_8550);
and U8764 (N_8764,N_8699,N_8632);
and U8765 (N_8765,N_8522,N_8417);
and U8766 (N_8766,N_8525,N_8462);
nor U8767 (N_8767,N_8552,N_8591);
nor U8768 (N_8768,N_8698,N_8535);
nor U8769 (N_8769,N_8528,N_8503);
or U8770 (N_8770,N_8456,N_8490);
nand U8771 (N_8771,N_8406,N_8526);
nor U8772 (N_8772,N_8545,N_8573);
xor U8773 (N_8773,N_8493,N_8639);
xnor U8774 (N_8774,N_8530,N_8484);
nand U8775 (N_8775,N_8485,N_8469);
or U8776 (N_8776,N_8497,N_8630);
or U8777 (N_8777,N_8570,N_8463);
nand U8778 (N_8778,N_8660,N_8563);
and U8779 (N_8779,N_8606,N_8642);
nand U8780 (N_8780,N_8507,N_8555);
nor U8781 (N_8781,N_8516,N_8455);
or U8782 (N_8782,N_8441,N_8587);
nand U8783 (N_8783,N_8464,N_8429);
xor U8784 (N_8784,N_8603,N_8450);
xor U8785 (N_8785,N_8483,N_8415);
xor U8786 (N_8786,N_8474,N_8578);
and U8787 (N_8787,N_8689,N_8574);
nor U8788 (N_8788,N_8445,N_8506);
xor U8789 (N_8789,N_8499,N_8542);
xor U8790 (N_8790,N_8477,N_8471);
xor U8791 (N_8791,N_8586,N_8548);
or U8792 (N_8792,N_8435,N_8412);
nor U8793 (N_8793,N_8431,N_8658);
or U8794 (N_8794,N_8605,N_8589);
nor U8795 (N_8795,N_8457,N_8482);
and U8796 (N_8796,N_8595,N_8686);
xnor U8797 (N_8797,N_8468,N_8426);
nand U8798 (N_8798,N_8610,N_8682);
nor U8799 (N_8799,N_8519,N_8626);
nor U8800 (N_8800,N_8559,N_8649);
and U8801 (N_8801,N_8683,N_8663);
and U8802 (N_8802,N_8510,N_8597);
and U8803 (N_8803,N_8553,N_8466);
nor U8804 (N_8804,N_8581,N_8557);
nand U8805 (N_8805,N_8618,N_8512);
xor U8806 (N_8806,N_8593,N_8521);
or U8807 (N_8807,N_8675,N_8540);
xnor U8808 (N_8808,N_8565,N_8461);
xnor U8809 (N_8809,N_8577,N_8664);
or U8810 (N_8810,N_8427,N_8644);
and U8811 (N_8811,N_8590,N_8571);
and U8812 (N_8812,N_8487,N_8432);
xor U8813 (N_8813,N_8596,N_8694);
nor U8814 (N_8814,N_8669,N_8543);
and U8815 (N_8815,N_8444,N_8500);
nand U8816 (N_8816,N_8434,N_8481);
or U8817 (N_8817,N_8498,N_8508);
or U8818 (N_8818,N_8423,N_8695);
xnor U8819 (N_8819,N_8612,N_8505);
or U8820 (N_8820,N_8436,N_8662);
nor U8821 (N_8821,N_8685,N_8640);
nor U8822 (N_8822,N_8425,N_8584);
xnor U8823 (N_8823,N_8411,N_8607);
xor U8824 (N_8824,N_8671,N_8598);
xor U8825 (N_8825,N_8541,N_8621);
or U8826 (N_8826,N_8696,N_8467);
nor U8827 (N_8827,N_8416,N_8404);
nor U8828 (N_8828,N_8447,N_8638);
nand U8829 (N_8829,N_8646,N_8428);
nor U8830 (N_8830,N_8509,N_8592);
nor U8831 (N_8831,N_8480,N_8600);
xor U8832 (N_8832,N_8633,N_8409);
or U8833 (N_8833,N_8615,N_8515);
or U8834 (N_8834,N_8421,N_8692);
and U8835 (N_8835,N_8539,N_8534);
and U8836 (N_8836,N_8585,N_8403);
nand U8837 (N_8837,N_8623,N_8478);
nand U8838 (N_8838,N_8524,N_8602);
or U8839 (N_8839,N_8440,N_8634);
or U8840 (N_8840,N_8402,N_8454);
xnor U8841 (N_8841,N_8443,N_8511);
and U8842 (N_8842,N_8400,N_8599);
and U8843 (N_8843,N_8690,N_8451);
nor U8844 (N_8844,N_8651,N_8636);
nor U8845 (N_8845,N_8446,N_8504);
or U8846 (N_8846,N_8575,N_8430);
xnor U8847 (N_8847,N_8551,N_8687);
and U8848 (N_8848,N_8517,N_8413);
nor U8849 (N_8849,N_8476,N_8562);
or U8850 (N_8850,N_8406,N_8634);
xnor U8851 (N_8851,N_8430,N_8567);
or U8852 (N_8852,N_8466,N_8462);
nor U8853 (N_8853,N_8621,N_8557);
and U8854 (N_8854,N_8687,N_8445);
or U8855 (N_8855,N_8578,N_8636);
nor U8856 (N_8856,N_8428,N_8557);
xor U8857 (N_8857,N_8577,N_8656);
nor U8858 (N_8858,N_8547,N_8460);
nand U8859 (N_8859,N_8621,N_8429);
and U8860 (N_8860,N_8684,N_8459);
xnor U8861 (N_8861,N_8467,N_8426);
and U8862 (N_8862,N_8497,N_8553);
xor U8863 (N_8863,N_8591,N_8601);
nor U8864 (N_8864,N_8663,N_8430);
or U8865 (N_8865,N_8491,N_8507);
nor U8866 (N_8866,N_8682,N_8458);
or U8867 (N_8867,N_8692,N_8401);
xor U8868 (N_8868,N_8639,N_8533);
xnor U8869 (N_8869,N_8611,N_8403);
or U8870 (N_8870,N_8480,N_8512);
or U8871 (N_8871,N_8603,N_8680);
xor U8872 (N_8872,N_8668,N_8670);
xor U8873 (N_8873,N_8680,N_8597);
or U8874 (N_8874,N_8424,N_8493);
xnor U8875 (N_8875,N_8425,N_8640);
xnor U8876 (N_8876,N_8495,N_8681);
nor U8877 (N_8877,N_8520,N_8570);
nand U8878 (N_8878,N_8437,N_8626);
xnor U8879 (N_8879,N_8576,N_8687);
nor U8880 (N_8880,N_8685,N_8482);
nor U8881 (N_8881,N_8514,N_8595);
nor U8882 (N_8882,N_8520,N_8458);
nand U8883 (N_8883,N_8565,N_8412);
or U8884 (N_8884,N_8479,N_8575);
nand U8885 (N_8885,N_8457,N_8621);
nand U8886 (N_8886,N_8498,N_8679);
and U8887 (N_8887,N_8649,N_8642);
nand U8888 (N_8888,N_8419,N_8524);
and U8889 (N_8889,N_8490,N_8564);
nor U8890 (N_8890,N_8623,N_8690);
or U8891 (N_8891,N_8587,N_8595);
nand U8892 (N_8892,N_8530,N_8513);
and U8893 (N_8893,N_8448,N_8683);
and U8894 (N_8894,N_8571,N_8609);
nand U8895 (N_8895,N_8654,N_8651);
or U8896 (N_8896,N_8448,N_8645);
and U8897 (N_8897,N_8604,N_8609);
nor U8898 (N_8898,N_8414,N_8484);
nor U8899 (N_8899,N_8674,N_8499);
nor U8900 (N_8900,N_8568,N_8449);
or U8901 (N_8901,N_8439,N_8523);
nor U8902 (N_8902,N_8529,N_8683);
nor U8903 (N_8903,N_8586,N_8526);
nor U8904 (N_8904,N_8625,N_8536);
nor U8905 (N_8905,N_8680,N_8415);
xnor U8906 (N_8906,N_8427,N_8694);
or U8907 (N_8907,N_8448,N_8621);
and U8908 (N_8908,N_8585,N_8590);
or U8909 (N_8909,N_8445,N_8650);
and U8910 (N_8910,N_8432,N_8502);
xor U8911 (N_8911,N_8661,N_8668);
and U8912 (N_8912,N_8488,N_8649);
xnor U8913 (N_8913,N_8568,N_8587);
or U8914 (N_8914,N_8569,N_8432);
nor U8915 (N_8915,N_8559,N_8424);
xnor U8916 (N_8916,N_8441,N_8642);
or U8917 (N_8917,N_8652,N_8499);
or U8918 (N_8918,N_8500,N_8667);
nand U8919 (N_8919,N_8686,N_8658);
and U8920 (N_8920,N_8419,N_8586);
nand U8921 (N_8921,N_8451,N_8647);
xor U8922 (N_8922,N_8458,N_8415);
or U8923 (N_8923,N_8593,N_8636);
nor U8924 (N_8924,N_8434,N_8432);
or U8925 (N_8925,N_8507,N_8468);
nand U8926 (N_8926,N_8525,N_8488);
and U8927 (N_8927,N_8499,N_8434);
xor U8928 (N_8928,N_8503,N_8519);
or U8929 (N_8929,N_8516,N_8505);
nor U8930 (N_8930,N_8470,N_8407);
xor U8931 (N_8931,N_8562,N_8664);
and U8932 (N_8932,N_8543,N_8633);
nor U8933 (N_8933,N_8478,N_8558);
nor U8934 (N_8934,N_8441,N_8551);
nor U8935 (N_8935,N_8412,N_8467);
or U8936 (N_8936,N_8686,N_8512);
or U8937 (N_8937,N_8677,N_8426);
or U8938 (N_8938,N_8608,N_8401);
nor U8939 (N_8939,N_8693,N_8577);
nor U8940 (N_8940,N_8418,N_8617);
nor U8941 (N_8941,N_8529,N_8467);
and U8942 (N_8942,N_8404,N_8564);
nand U8943 (N_8943,N_8656,N_8452);
nor U8944 (N_8944,N_8604,N_8480);
and U8945 (N_8945,N_8572,N_8652);
and U8946 (N_8946,N_8444,N_8545);
or U8947 (N_8947,N_8589,N_8428);
or U8948 (N_8948,N_8480,N_8425);
nor U8949 (N_8949,N_8456,N_8636);
and U8950 (N_8950,N_8492,N_8503);
nor U8951 (N_8951,N_8522,N_8534);
or U8952 (N_8952,N_8413,N_8678);
and U8953 (N_8953,N_8684,N_8623);
nor U8954 (N_8954,N_8695,N_8592);
nand U8955 (N_8955,N_8547,N_8458);
xor U8956 (N_8956,N_8659,N_8403);
or U8957 (N_8957,N_8606,N_8548);
nor U8958 (N_8958,N_8671,N_8617);
nor U8959 (N_8959,N_8657,N_8432);
and U8960 (N_8960,N_8559,N_8590);
nor U8961 (N_8961,N_8416,N_8423);
xnor U8962 (N_8962,N_8425,N_8523);
or U8963 (N_8963,N_8629,N_8633);
xor U8964 (N_8964,N_8692,N_8643);
nor U8965 (N_8965,N_8664,N_8472);
xnor U8966 (N_8966,N_8484,N_8411);
nand U8967 (N_8967,N_8454,N_8414);
nand U8968 (N_8968,N_8580,N_8404);
xnor U8969 (N_8969,N_8550,N_8505);
nor U8970 (N_8970,N_8670,N_8693);
nand U8971 (N_8971,N_8607,N_8435);
nand U8972 (N_8972,N_8562,N_8561);
xor U8973 (N_8973,N_8524,N_8680);
xor U8974 (N_8974,N_8691,N_8605);
nor U8975 (N_8975,N_8604,N_8646);
or U8976 (N_8976,N_8656,N_8564);
and U8977 (N_8977,N_8628,N_8511);
and U8978 (N_8978,N_8672,N_8401);
nand U8979 (N_8979,N_8653,N_8482);
nand U8980 (N_8980,N_8620,N_8506);
and U8981 (N_8981,N_8579,N_8658);
and U8982 (N_8982,N_8488,N_8558);
nor U8983 (N_8983,N_8614,N_8691);
nand U8984 (N_8984,N_8665,N_8644);
or U8985 (N_8985,N_8524,N_8426);
or U8986 (N_8986,N_8424,N_8626);
and U8987 (N_8987,N_8566,N_8584);
or U8988 (N_8988,N_8555,N_8671);
nand U8989 (N_8989,N_8515,N_8406);
or U8990 (N_8990,N_8625,N_8497);
or U8991 (N_8991,N_8430,N_8592);
and U8992 (N_8992,N_8660,N_8637);
xor U8993 (N_8993,N_8651,N_8460);
xor U8994 (N_8994,N_8561,N_8510);
and U8995 (N_8995,N_8656,N_8434);
nand U8996 (N_8996,N_8520,N_8413);
xor U8997 (N_8997,N_8660,N_8455);
and U8998 (N_8998,N_8543,N_8553);
and U8999 (N_8999,N_8546,N_8623);
or U9000 (N_9000,N_8751,N_8957);
nor U9001 (N_9001,N_8834,N_8809);
nand U9002 (N_9002,N_8730,N_8922);
and U9003 (N_9003,N_8852,N_8725);
xor U9004 (N_9004,N_8705,N_8918);
or U9005 (N_9005,N_8975,N_8797);
or U9006 (N_9006,N_8754,N_8897);
nor U9007 (N_9007,N_8927,N_8825);
nand U9008 (N_9008,N_8937,N_8771);
xor U9009 (N_9009,N_8729,N_8710);
nand U9010 (N_9010,N_8945,N_8946);
xnor U9011 (N_9011,N_8909,N_8917);
or U9012 (N_9012,N_8719,N_8798);
nand U9013 (N_9013,N_8989,N_8902);
nand U9014 (N_9014,N_8805,N_8838);
nor U9015 (N_9015,N_8837,N_8704);
nor U9016 (N_9016,N_8905,N_8858);
or U9017 (N_9017,N_8815,N_8867);
nor U9018 (N_9018,N_8864,N_8877);
or U9019 (N_9019,N_8987,N_8854);
xor U9020 (N_9020,N_8804,N_8847);
nand U9021 (N_9021,N_8747,N_8986);
nor U9022 (N_9022,N_8718,N_8776);
and U9023 (N_9023,N_8748,N_8742);
nand U9024 (N_9024,N_8703,N_8930);
or U9025 (N_9025,N_8994,N_8795);
or U9026 (N_9026,N_8788,N_8843);
or U9027 (N_9027,N_8898,N_8876);
nor U9028 (N_9028,N_8723,N_8781);
nor U9029 (N_9029,N_8882,N_8701);
nor U9030 (N_9030,N_8850,N_8941);
and U9031 (N_9031,N_8961,N_8849);
xnor U9032 (N_9032,N_8855,N_8801);
nand U9033 (N_9033,N_8911,N_8728);
xor U9034 (N_9034,N_8949,N_8839);
nor U9035 (N_9035,N_8840,N_8991);
nor U9036 (N_9036,N_8845,N_8870);
nand U9037 (N_9037,N_8908,N_8965);
nand U9038 (N_9038,N_8915,N_8831);
nor U9039 (N_9039,N_8868,N_8836);
xnor U9040 (N_9040,N_8958,N_8889);
nor U9041 (N_9041,N_8990,N_8980);
or U9042 (N_9042,N_8977,N_8765);
and U9043 (N_9043,N_8966,N_8921);
nor U9044 (N_9044,N_8952,N_8794);
nand U9045 (N_9045,N_8919,N_8786);
nand U9046 (N_9046,N_8924,N_8873);
nand U9047 (N_9047,N_8779,N_8862);
xor U9048 (N_9048,N_8819,N_8931);
xnor U9049 (N_9049,N_8861,N_8820);
xor U9050 (N_9050,N_8948,N_8724);
or U9051 (N_9051,N_8829,N_8901);
or U9052 (N_9052,N_8981,N_8762);
xor U9053 (N_9053,N_8740,N_8885);
and U9054 (N_9054,N_8846,N_8892);
xor U9055 (N_9055,N_8928,N_8722);
or U9056 (N_9056,N_8835,N_8973);
nand U9057 (N_9057,N_8733,N_8950);
nor U9058 (N_9058,N_8817,N_8960);
nand U9059 (N_9059,N_8784,N_8851);
or U9060 (N_9060,N_8974,N_8772);
and U9061 (N_9061,N_8875,N_8992);
xor U9062 (N_9062,N_8793,N_8976);
nor U9063 (N_9063,N_8899,N_8757);
nand U9064 (N_9064,N_8709,N_8964);
nor U9065 (N_9065,N_8844,N_8866);
and U9066 (N_9066,N_8770,N_8821);
nor U9067 (N_9067,N_8741,N_8893);
nand U9068 (N_9068,N_8979,N_8951);
xor U9069 (N_9069,N_8983,N_8760);
or U9070 (N_9070,N_8953,N_8783);
xor U9071 (N_9071,N_8803,N_8763);
xnor U9072 (N_9072,N_8887,N_8932);
nor U9073 (N_9073,N_8860,N_8780);
nor U9074 (N_9074,N_8954,N_8929);
nor U9075 (N_9075,N_8947,N_8886);
or U9076 (N_9076,N_8792,N_8942);
or U9077 (N_9077,N_8714,N_8769);
nand U9078 (N_9078,N_8894,N_8767);
and U9079 (N_9079,N_8939,N_8743);
or U9080 (N_9080,N_8832,N_8717);
xnor U9081 (N_9081,N_8735,N_8796);
nand U9082 (N_9082,N_8972,N_8824);
xor U9083 (N_9083,N_8857,N_8826);
nor U9084 (N_9084,N_8955,N_8700);
xor U9085 (N_9085,N_8906,N_8812);
and U9086 (N_9086,N_8785,N_8750);
or U9087 (N_9087,N_8993,N_8853);
nand U9088 (N_9088,N_8920,N_8995);
and U9089 (N_9089,N_8807,N_8752);
nand U9090 (N_9090,N_8956,N_8841);
or U9091 (N_9091,N_8738,N_8896);
and U9092 (N_9092,N_8878,N_8884);
nor U9093 (N_9093,N_8782,N_8967);
or U9094 (N_9094,N_8895,N_8944);
nand U9095 (N_9095,N_8963,N_8764);
nor U9096 (N_9096,N_8802,N_8913);
and U9097 (N_9097,N_8823,N_8758);
nand U9098 (N_9098,N_8756,N_8914);
or U9099 (N_9099,N_8736,N_8806);
nor U9100 (N_9100,N_8856,N_8891);
and U9101 (N_9101,N_8833,N_8810);
xor U9102 (N_9102,N_8934,N_8745);
or U9103 (N_9103,N_8962,N_8936);
or U9104 (N_9104,N_8923,N_8814);
nor U9105 (N_9105,N_8808,N_8778);
nor U9106 (N_9106,N_8985,N_8737);
xor U9107 (N_9107,N_8706,N_8938);
nor U9108 (N_9108,N_8871,N_8800);
or U9109 (N_9109,N_8744,N_8789);
nand U9110 (N_9110,N_8720,N_8926);
and U9111 (N_9111,N_8818,N_8900);
or U9112 (N_9112,N_8982,N_8816);
nand U9113 (N_9113,N_8726,N_8734);
nor U9114 (N_9114,N_8827,N_8880);
or U9115 (N_9115,N_8865,N_8761);
or U9116 (N_9116,N_8910,N_8707);
nor U9117 (N_9117,N_8766,N_8969);
and U9118 (N_9118,N_8996,N_8881);
nand U9119 (N_9119,N_8890,N_8925);
nor U9120 (N_9120,N_8916,N_8848);
or U9121 (N_9121,N_8904,N_8903);
and U9122 (N_9122,N_8759,N_8768);
nand U9123 (N_9123,N_8716,N_8732);
nor U9124 (N_9124,N_8999,N_8988);
nand U9125 (N_9125,N_8940,N_8912);
xnor U9126 (N_9126,N_8883,N_8830);
xor U9127 (N_9127,N_8859,N_8813);
nor U9128 (N_9128,N_8787,N_8774);
or U9129 (N_9129,N_8721,N_8874);
nor U9130 (N_9130,N_8775,N_8777);
xor U9131 (N_9131,N_8799,N_8888);
or U9132 (N_9132,N_8746,N_8978);
or U9133 (N_9133,N_8739,N_8822);
nor U9134 (N_9134,N_8943,N_8755);
and U9135 (N_9135,N_8879,N_8997);
nand U9136 (N_9136,N_8907,N_8811);
nand U9137 (N_9137,N_8872,N_8828);
and U9138 (N_9138,N_8790,N_8968);
and U9139 (N_9139,N_8984,N_8708);
nand U9140 (N_9140,N_8711,N_8842);
and U9141 (N_9141,N_8773,N_8749);
and U9142 (N_9142,N_8970,N_8791);
nand U9143 (N_9143,N_8935,N_8933);
xor U9144 (N_9144,N_8971,N_8712);
xnor U9145 (N_9145,N_8998,N_8715);
xnor U9146 (N_9146,N_8863,N_8731);
nand U9147 (N_9147,N_8869,N_8727);
nand U9148 (N_9148,N_8959,N_8753);
or U9149 (N_9149,N_8713,N_8702);
nor U9150 (N_9150,N_8995,N_8782);
and U9151 (N_9151,N_8795,N_8933);
nor U9152 (N_9152,N_8885,N_8879);
or U9153 (N_9153,N_8863,N_8940);
and U9154 (N_9154,N_8839,N_8779);
or U9155 (N_9155,N_8839,N_8785);
xor U9156 (N_9156,N_8958,N_8794);
and U9157 (N_9157,N_8985,N_8855);
nand U9158 (N_9158,N_8772,N_8713);
xnor U9159 (N_9159,N_8774,N_8943);
or U9160 (N_9160,N_8868,N_8747);
or U9161 (N_9161,N_8823,N_8861);
and U9162 (N_9162,N_8976,N_8886);
nand U9163 (N_9163,N_8819,N_8860);
and U9164 (N_9164,N_8750,N_8905);
nor U9165 (N_9165,N_8934,N_8941);
or U9166 (N_9166,N_8915,N_8851);
nor U9167 (N_9167,N_8834,N_8728);
and U9168 (N_9168,N_8862,N_8750);
or U9169 (N_9169,N_8767,N_8808);
nor U9170 (N_9170,N_8948,N_8810);
nor U9171 (N_9171,N_8841,N_8833);
nand U9172 (N_9172,N_8724,N_8860);
and U9173 (N_9173,N_8731,N_8988);
and U9174 (N_9174,N_8972,N_8706);
or U9175 (N_9175,N_8780,N_8841);
and U9176 (N_9176,N_8700,N_8932);
nor U9177 (N_9177,N_8784,N_8902);
and U9178 (N_9178,N_8996,N_8849);
xnor U9179 (N_9179,N_8895,N_8869);
or U9180 (N_9180,N_8925,N_8870);
or U9181 (N_9181,N_8822,N_8722);
nand U9182 (N_9182,N_8933,N_8943);
nor U9183 (N_9183,N_8790,N_8944);
nor U9184 (N_9184,N_8889,N_8919);
xnor U9185 (N_9185,N_8872,N_8732);
nor U9186 (N_9186,N_8847,N_8839);
nor U9187 (N_9187,N_8815,N_8912);
xor U9188 (N_9188,N_8992,N_8840);
or U9189 (N_9189,N_8908,N_8847);
xor U9190 (N_9190,N_8963,N_8819);
nor U9191 (N_9191,N_8727,N_8822);
and U9192 (N_9192,N_8926,N_8782);
xnor U9193 (N_9193,N_8795,N_8791);
nor U9194 (N_9194,N_8781,N_8727);
xnor U9195 (N_9195,N_8890,N_8850);
xnor U9196 (N_9196,N_8749,N_8734);
nor U9197 (N_9197,N_8707,N_8778);
and U9198 (N_9198,N_8879,N_8860);
or U9199 (N_9199,N_8936,N_8715);
or U9200 (N_9200,N_8714,N_8771);
nor U9201 (N_9201,N_8743,N_8973);
xnor U9202 (N_9202,N_8855,N_8792);
xor U9203 (N_9203,N_8976,N_8978);
xor U9204 (N_9204,N_8782,N_8994);
nand U9205 (N_9205,N_8722,N_8920);
nand U9206 (N_9206,N_8870,N_8985);
nand U9207 (N_9207,N_8778,N_8844);
xnor U9208 (N_9208,N_8969,N_8789);
xnor U9209 (N_9209,N_8730,N_8775);
xor U9210 (N_9210,N_8837,N_8917);
nor U9211 (N_9211,N_8871,N_8787);
xnor U9212 (N_9212,N_8786,N_8868);
and U9213 (N_9213,N_8913,N_8797);
nand U9214 (N_9214,N_8887,N_8742);
and U9215 (N_9215,N_8925,N_8989);
nand U9216 (N_9216,N_8800,N_8945);
and U9217 (N_9217,N_8958,N_8744);
nand U9218 (N_9218,N_8855,N_8881);
nor U9219 (N_9219,N_8925,N_8929);
and U9220 (N_9220,N_8790,N_8959);
nand U9221 (N_9221,N_8716,N_8833);
or U9222 (N_9222,N_8724,N_8919);
or U9223 (N_9223,N_8830,N_8784);
nor U9224 (N_9224,N_8938,N_8968);
xnor U9225 (N_9225,N_8926,N_8738);
nor U9226 (N_9226,N_8953,N_8889);
nor U9227 (N_9227,N_8723,N_8720);
and U9228 (N_9228,N_8730,N_8851);
and U9229 (N_9229,N_8882,N_8781);
xor U9230 (N_9230,N_8924,N_8729);
xor U9231 (N_9231,N_8940,N_8991);
xnor U9232 (N_9232,N_8890,N_8837);
nor U9233 (N_9233,N_8821,N_8710);
and U9234 (N_9234,N_8904,N_8890);
or U9235 (N_9235,N_8756,N_8860);
nand U9236 (N_9236,N_8927,N_8784);
or U9237 (N_9237,N_8726,N_8731);
or U9238 (N_9238,N_8971,N_8931);
and U9239 (N_9239,N_8931,N_8759);
nand U9240 (N_9240,N_8822,N_8756);
xor U9241 (N_9241,N_8908,N_8860);
nand U9242 (N_9242,N_8796,N_8875);
xor U9243 (N_9243,N_8867,N_8899);
nor U9244 (N_9244,N_8932,N_8795);
nor U9245 (N_9245,N_8940,N_8794);
nand U9246 (N_9246,N_8900,N_8765);
xor U9247 (N_9247,N_8735,N_8826);
nor U9248 (N_9248,N_8910,N_8830);
or U9249 (N_9249,N_8976,N_8945);
or U9250 (N_9250,N_8942,N_8811);
and U9251 (N_9251,N_8989,N_8829);
and U9252 (N_9252,N_8952,N_8763);
nand U9253 (N_9253,N_8720,N_8849);
nand U9254 (N_9254,N_8997,N_8751);
xnor U9255 (N_9255,N_8927,N_8742);
or U9256 (N_9256,N_8898,N_8723);
and U9257 (N_9257,N_8771,N_8873);
nand U9258 (N_9258,N_8968,N_8882);
nand U9259 (N_9259,N_8795,N_8902);
or U9260 (N_9260,N_8976,N_8825);
or U9261 (N_9261,N_8701,N_8727);
nand U9262 (N_9262,N_8738,N_8727);
xor U9263 (N_9263,N_8894,N_8836);
nand U9264 (N_9264,N_8938,N_8957);
nor U9265 (N_9265,N_8716,N_8850);
nor U9266 (N_9266,N_8895,N_8717);
and U9267 (N_9267,N_8780,N_8919);
and U9268 (N_9268,N_8970,N_8715);
xor U9269 (N_9269,N_8877,N_8851);
xnor U9270 (N_9270,N_8745,N_8947);
nor U9271 (N_9271,N_8837,N_8767);
xor U9272 (N_9272,N_8775,N_8872);
or U9273 (N_9273,N_8732,N_8819);
or U9274 (N_9274,N_8756,N_8839);
nor U9275 (N_9275,N_8726,N_8702);
nor U9276 (N_9276,N_8907,N_8980);
and U9277 (N_9277,N_8810,N_8991);
nand U9278 (N_9278,N_8841,N_8876);
nor U9279 (N_9279,N_8758,N_8828);
and U9280 (N_9280,N_8962,N_8922);
or U9281 (N_9281,N_8946,N_8800);
nor U9282 (N_9282,N_8886,N_8863);
and U9283 (N_9283,N_8796,N_8968);
nor U9284 (N_9284,N_8720,N_8967);
xnor U9285 (N_9285,N_8848,N_8862);
and U9286 (N_9286,N_8958,N_8975);
and U9287 (N_9287,N_8806,N_8793);
xor U9288 (N_9288,N_8814,N_8855);
or U9289 (N_9289,N_8783,N_8967);
nor U9290 (N_9290,N_8885,N_8867);
nand U9291 (N_9291,N_8793,N_8974);
xnor U9292 (N_9292,N_8908,N_8702);
nand U9293 (N_9293,N_8983,N_8778);
nand U9294 (N_9294,N_8932,N_8905);
or U9295 (N_9295,N_8729,N_8904);
and U9296 (N_9296,N_8944,N_8896);
nor U9297 (N_9297,N_8758,N_8858);
and U9298 (N_9298,N_8700,N_8764);
xnor U9299 (N_9299,N_8801,N_8907);
nand U9300 (N_9300,N_9071,N_9141);
and U9301 (N_9301,N_9139,N_9003);
nor U9302 (N_9302,N_9197,N_9276);
nor U9303 (N_9303,N_9115,N_9161);
and U9304 (N_9304,N_9093,N_9210);
xor U9305 (N_9305,N_9116,N_9050);
xor U9306 (N_9306,N_9207,N_9005);
nand U9307 (N_9307,N_9124,N_9002);
nor U9308 (N_9308,N_9034,N_9281);
and U9309 (N_9309,N_9042,N_9246);
xor U9310 (N_9310,N_9275,N_9140);
xor U9311 (N_9311,N_9172,N_9152);
nor U9312 (N_9312,N_9015,N_9279);
and U9313 (N_9313,N_9258,N_9126);
and U9314 (N_9314,N_9128,N_9021);
xnor U9315 (N_9315,N_9202,N_9066);
and U9316 (N_9316,N_9223,N_9182);
or U9317 (N_9317,N_9144,N_9186);
nor U9318 (N_9318,N_9272,N_9104);
or U9319 (N_9319,N_9195,N_9047);
nor U9320 (N_9320,N_9263,N_9082);
nand U9321 (N_9321,N_9067,N_9100);
nor U9322 (N_9322,N_9029,N_9169);
nand U9323 (N_9323,N_9170,N_9127);
nand U9324 (N_9324,N_9296,N_9295);
or U9325 (N_9325,N_9048,N_9287);
nor U9326 (N_9326,N_9038,N_9228);
xnor U9327 (N_9327,N_9226,N_9289);
nor U9328 (N_9328,N_9249,N_9240);
and U9329 (N_9329,N_9111,N_9282);
or U9330 (N_9330,N_9168,N_9227);
and U9331 (N_9331,N_9030,N_9268);
and U9332 (N_9332,N_9065,N_9235);
and U9333 (N_9333,N_9175,N_9114);
or U9334 (N_9334,N_9262,N_9232);
nand U9335 (N_9335,N_9159,N_9057);
nor U9336 (N_9336,N_9173,N_9132);
nand U9337 (N_9337,N_9131,N_9203);
xnor U9338 (N_9338,N_9072,N_9251);
or U9339 (N_9339,N_9119,N_9062);
xor U9340 (N_9340,N_9183,N_9255);
nand U9341 (N_9341,N_9288,N_9294);
nor U9342 (N_9342,N_9107,N_9120);
xor U9343 (N_9343,N_9108,N_9266);
and U9344 (N_9344,N_9110,N_9181);
or U9345 (N_9345,N_9176,N_9166);
xor U9346 (N_9346,N_9164,N_9280);
xor U9347 (N_9347,N_9222,N_9095);
nand U9348 (N_9348,N_9200,N_9103);
or U9349 (N_9349,N_9134,N_9231);
or U9350 (N_9350,N_9081,N_9083);
or U9351 (N_9351,N_9112,N_9022);
or U9352 (N_9352,N_9009,N_9193);
xnor U9353 (N_9353,N_9273,N_9269);
nand U9354 (N_9354,N_9135,N_9089);
or U9355 (N_9355,N_9234,N_9055);
or U9356 (N_9356,N_9018,N_9201);
nand U9357 (N_9357,N_9059,N_9061);
nor U9358 (N_9358,N_9239,N_9291);
nand U9359 (N_9359,N_9122,N_9014);
nor U9360 (N_9360,N_9206,N_9220);
nand U9361 (N_9361,N_9041,N_9293);
nor U9362 (N_9362,N_9233,N_9040);
and U9363 (N_9363,N_9218,N_9253);
or U9364 (N_9364,N_9184,N_9180);
and U9365 (N_9365,N_9052,N_9292);
or U9366 (N_9366,N_9084,N_9221);
nand U9367 (N_9367,N_9213,N_9076);
and U9368 (N_9368,N_9162,N_9241);
and U9369 (N_9369,N_9204,N_9118);
nor U9370 (N_9370,N_9027,N_9211);
nor U9371 (N_9371,N_9219,N_9187);
nand U9372 (N_9372,N_9056,N_9199);
nand U9373 (N_9373,N_9045,N_9245);
and U9374 (N_9374,N_9121,N_9020);
nand U9375 (N_9375,N_9259,N_9019);
xor U9376 (N_9376,N_9033,N_9063);
nor U9377 (N_9377,N_9123,N_9088);
or U9378 (N_9378,N_9286,N_9190);
nor U9379 (N_9379,N_9277,N_9043);
and U9380 (N_9380,N_9230,N_9053);
and U9381 (N_9381,N_9174,N_9085);
and U9382 (N_9382,N_9150,N_9224);
or U9383 (N_9383,N_9004,N_9125);
nor U9384 (N_9384,N_9192,N_9148);
nor U9385 (N_9385,N_9205,N_9060);
nor U9386 (N_9386,N_9297,N_9189);
or U9387 (N_9387,N_9285,N_9080);
nand U9388 (N_9388,N_9267,N_9260);
and U9389 (N_9389,N_9145,N_9007);
nand U9390 (N_9390,N_9079,N_9271);
and U9391 (N_9391,N_9151,N_9244);
xor U9392 (N_9392,N_9087,N_9215);
nor U9393 (N_9393,N_9248,N_9264);
nor U9394 (N_9394,N_9133,N_9237);
xor U9395 (N_9395,N_9212,N_9137);
nor U9396 (N_9396,N_9142,N_9031);
and U9397 (N_9397,N_9178,N_9208);
nor U9398 (N_9398,N_9153,N_9252);
nor U9399 (N_9399,N_9035,N_9278);
and U9400 (N_9400,N_9086,N_9191);
xnor U9401 (N_9401,N_9026,N_9024);
nor U9402 (N_9402,N_9070,N_9250);
nand U9403 (N_9403,N_9194,N_9000);
nand U9404 (N_9404,N_9049,N_9146);
and U9405 (N_9405,N_9274,N_9214);
nor U9406 (N_9406,N_9163,N_9097);
nor U9407 (N_9407,N_9036,N_9265);
and U9408 (N_9408,N_9037,N_9078);
and U9409 (N_9409,N_9069,N_9068);
nand U9410 (N_9410,N_9028,N_9058);
nor U9411 (N_9411,N_9270,N_9136);
xnor U9412 (N_9412,N_9147,N_9098);
nor U9413 (N_9413,N_9074,N_9298);
xnor U9414 (N_9414,N_9243,N_9023);
or U9415 (N_9415,N_9032,N_9094);
and U9416 (N_9416,N_9051,N_9257);
nand U9417 (N_9417,N_9238,N_9109);
nand U9418 (N_9418,N_9171,N_9016);
or U9419 (N_9419,N_9091,N_9188);
or U9420 (N_9420,N_9077,N_9283);
nor U9421 (N_9421,N_9113,N_9001);
xor U9422 (N_9422,N_9101,N_9256);
or U9423 (N_9423,N_9198,N_9158);
nor U9424 (N_9424,N_9129,N_9130);
nand U9425 (N_9425,N_9154,N_9160);
and U9426 (N_9426,N_9254,N_9225);
and U9427 (N_9427,N_9143,N_9236);
and U9428 (N_9428,N_9284,N_9149);
and U9429 (N_9429,N_9054,N_9177);
nand U9430 (N_9430,N_9044,N_9229);
and U9431 (N_9431,N_9099,N_9011);
nand U9432 (N_9432,N_9106,N_9092);
and U9433 (N_9433,N_9261,N_9299);
or U9434 (N_9434,N_9138,N_9247);
and U9435 (N_9435,N_9008,N_9217);
nand U9436 (N_9436,N_9010,N_9290);
and U9437 (N_9437,N_9196,N_9185);
nand U9438 (N_9438,N_9179,N_9102);
xnor U9439 (N_9439,N_9096,N_9209);
or U9440 (N_9440,N_9039,N_9155);
nor U9441 (N_9441,N_9117,N_9216);
and U9442 (N_9442,N_9167,N_9105);
nand U9443 (N_9443,N_9156,N_9073);
nor U9444 (N_9444,N_9017,N_9012);
or U9445 (N_9445,N_9090,N_9157);
nor U9446 (N_9446,N_9025,N_9013);
and U9447 (N_9447,N_9006,N_9064);
and U9448 (N_9448,N_9242,N_9165);
nand U9449 (N_9449,N_9046,N_9075);
or U9450 (N_9450,N_9294,N_9299);
and U9451 (N_9451,N_9137,N_9082);
or U9452 (N_9452,N_9223,N_9126);
nand U9453 (N_9453,N_9123,N_9049);
nand U9454 (N_9454,N_9090,N_9136);
and U9455 (N_9455,N_9204,N_9068);
xnor U9456 (N_9456,N_9085,N_9257);
or U9457 (N_9457,N_9237,N_9147);
nand U9458 (N_9458,N_9001,N_9165);
nand U9459 (N_9459,N_9031,N_9188);
nor U9460 (N_9460,N_9105,N_9288);
and U9461 (N_9461,N_9181,N_9221);
nor U9462 (N_9462,N_9288,N_9179);
or U9463 (N_9463,N_9188,N_9027);
nor U9464 (N_9464,N_9238,N_9290);
xor U9465 (N_9465,N_9275,N_9219);
xnor U9466 (N_9466,N_9103,N_9297);
xnor U9467 (N_9467,N_9088,N_9265);
xnor U9468 (N_9468,N_9071,N_9271);
or U9469 (N_9469,N_9218,N_9110);
and U9470 (N_9470,N_9167,N_9051);
nor U9471 (N_9471,N_9004,N_9285);
nor U9472 (N_9472,N_9298,N_9009);
nor U9473 (N_9473,N_9286,N_9241);
xor U9474 (N_9474,N_9252,N_9299);
or U9475 (N_9475,N_9236,N_9090);
or U9476 (N_9476,N_9228,N_9294);
or U9477 (N_9477,N_9093,N_9286);
xor U9478 (N_9478,N_9140,N_9137);
xnor U9479 (N_9479,N_9083,N_9037);
xnor U9480 (N_9480,N_9255,N_9018);
nor U9481 (N_9481,N_9195,N_9247);
nand U9482 (N_9482,N_9286,N_9024);
xor U9483 (N_9483,N_9231,N_9235);
or U9484 (N_9484,N_9233,N_9242);
or U9485 (N_9485,N_9087,N_9238);
xor U9486 (N_9486,N_9174,N_9058);
nand U9487 (N_9487,N_9049,N_9024);
xor U9488 (N_9488,N_9161,N_9255);
nor U9489 (N_9489,N_9122,N_9240);
or U9490 (N_9490,N_9079,N_9130);
and U9491 (N_9491,N_9263,N_9204);
or U9492 (N_9492,N_9271,N_9058);
or U9493 (N_9493,N_9042,N_9061);
or U9494 (N_9494,N_9021,N_9130);
nor U9495 (N_9495,N_9149,N_9275);
nand U9496 (N_9496,N_9219,N_9149);
nand U9497 (N_9497,N_9177,N_9086);
nand U9498 (N_9498,N_9151,N_9080);
and U9499 (N_9499,N_9212,N_9036);
and U9500 (N_9500,N_9058,N_9260);
and U9501 (N_9501,N_9191,N_9118);
xor U9502 (N_9502,N_9020,N_9001);
xnor U9503 (N_9503,N_9148,N_9235);
nor U9504 (N_9504,N_9030,N_9123);
and U9505 (N_9505,N_9170,N_9033);
xor U9506 (N_9506,N_9013,N_9157);
xor U9507 (N_9507,N_9299,N_9150);
and U9508 (N_9508,N_9235,N_9007);
or U9509 (N_9509,N_9057,N_9202);
nand U9510 (N_9510,N_9286,N_9140);
nor U9511 (N_9511,N_9240,N_9183);
or U9512 (N_9512,N_9074,N_9296);
xor U9513 (N_9513,N_9238,N_9299);
nor U9514 (N_9514,N_9222,N_9154);
nor U9515 (N_9515,N_9286,N_9273);
nor U9516 (N_9516,N_9006,N_9054);
or U9517 (N_9517,N_9159,N_9137);
nor U9518 (N_9518,N_9288,N_9184);
nand U9519 (N_9519,N_9040,N_9212);
nor U9520 (N_9520,N_9021,N_9105);
and U9521 (N_9521,N_9214,N_9124);
nor U9522 (N_9522,N_9247,N_9113);
nor U9523 (N_9523,N_9267,N_9038);
nand U9524 (N_9524,N_9116,N_9073);
and U9525 (N_9525,N_9101,N_9033);
or U9526 (N_9526,N_9034,N_9175);
and U9527 (N_9527,N_9165,N_9079);
and U9528 (N_9528,N_9129,N_9188);
nor U9529 (N_9529,N_9176,N_9197);
and U9530 (N_9530,N_9144,N_9085);
or U9531 (N_9531,N_9209,N_9279);
and U9532 (N_9532,N_9084,N_9211);
and U9533 (N_9533,N_9021,N_9272);
or U9534 (N_9534,N_9034,N_9190);
and U9535 (N_9535,N_9070,N_9166);
nand U9536 (N_9536,N_9198,N_9239);
or U9537 (N_9537,N_9031,N_9010);
and U9538 (N_9538,N_9106,N_9056);
or U9539 (N_9539,N_9198,N_9135);
nor U9540 (N_9540,N_9186,N_9157);
or U9541 (N_9541,N_9163,N_9090);
xnor U9542 (N_9542,N_9147,N_9203);
nand U9543 (N_9543,N_9202,N_9028);
xor U9544 (N_9544,N_9035,N_9270);
nor U9545 (N_9545,N_9039,N_9152);
nor U9546 (N_9546,N_9060,N_9219);
nand U9547 (N_9547,N_9246,N_9175);
nor U9548 (N_9548,N_9191,N_9242);
nor U9549 (N_9549,N_9251,N_9041);
nand U9550 (N_9550,N_9109,N_9031);
or U9551 (N_9551,N_9278,N_9225);
or U9552 (N_9552,N_9296,N_9190);
or U9553 (N_9553,N_9151,N_9279);
xnor U9554 (N_9554,N_9019,N_9163);
nand U9555 (N_9555,N_9104,N_9120);
and U9556 (N_9556,N_9050,N_9051);
or U9557 (N_9557,N_9203,N_9241);
xor U9558 (N_9558,N_9160,N_9032);
nand U9559 (N_9559,N_9053,N_9257);
nand U9560 (N_9560,N_9103,N_9275);
nor U9561 (N_9561,N_9181,N_9235);
nor U9562 (N_9562,N_9115,N_9010);
or U9563 (N_9563,N_9149,N_9260);
nand U9564 (N_9564,N_9253,N_9250);
nand U9565 (N_9565,N_9239,N_9179);
and U9566 (N_9566,N_9263,N_9075);
nand U9567 (N_9567,N_9131,N_9296);
and U9568 (N_9568,N_9257,N_9166);
xnor U9569 (N_9569,N_9178,N_9214);
and U9570 (N_9570,N_9162,N_9152);
nand U9571 (N_9571,N_9134,N_9140);
and U9572 (N_9572,N_9046,N_9032);
and U9573 (N_9573,N_9248,N_9104);
xor U9574 (N_9574,N_9142,N_9282);
and U9575 (N_9575,N_9001,N_9172);
and U9576 (N_9576,N_9235,N_9272);
nor U9577 (N_9577,N_9263,N_9288);
or U9578 (N_9578,N_9266,N_9100);
xor U9579 (N_9579,N_9207,N_9121);
nand U9580 (N_9580,N_9279,N_9145);
xnor U9581 (N_9581,N_9109,N_9000);
and U9582 (N_9582,N_9163,N_9149);
nor U9583 (N_9583,N_9299,N_9272);
or U9584 (N_9584,N_9210,N_9281);
and U9585 (N_9585,N_9085,N_9265);
xor U9586 (N_9586,N_9132,N_9213);
or U9587 (N_9587,N_9292,N_9100);
and U9588 (N_9588,N_9001,N_9109);
nor U9589 (N_9589,N_9106,N_9164);
nor U9590 (N_9590,N_9158,N_9214);
xnor U9591 (N_9591,N_9292,N_9272);
nor U9592 (N_9592,N_9291,N_9094);
nand U9593 (N_9593,N_9082,N_9186);
xnor U9594 (N_9594,N_9297,N_9168);
nand U9595 (N_9595,N_9197,N_9286);
nand U9596 (N_9596,N_9069,N_9217);
xor U9597 (N_9597,N_9042,N_9211);
and U9598 (N_9598,N_9162,N_9248);
nand U9599 (N_9599,N_9142,N_9158);
xnor U9600 (N_9600,N_9380,N_9493);
or U9601 (N_9601,N_9442,N_9490);
xor U9602 (N_9602,N_9571,N_9338);
or U9603 (N_9603,N_9535,N_9530);
nor U9604 (N_9604,N_9556,N_9585);
or U9605 (N_9605,N_9504,N_9435);
and U9606 (N_9606,N_9433,N_9588);
nand U9607 (N_9607,N_9545,N_9508);
xnor U9608 (N_9608,N_9596,N_9353);
nand U9609 (N_9609,N_9402,N_9472);
xor U9610 (N_9610,N_9500,N_9441);
xor U9611 (N_9611,N_9482,N_9356);
and U9612 (N_9612,N_9572,N_9448);
xor U9613 (N_9613,N_9319,N_9497);
and U9614 (N_9614,N_9534,N_9593);
or U9615 (N_9615,N_9552,N_9546);
xnor U9616 (N_9616,N_9479,N_9328);
or U9617 (N_9617,N_9345,N_9503);
xnor U9618 (N_9618,N_9458,N_9595);
and U9619 (N_9619,N_9540,N_9502);
xnor U9620 (N_9620,N_9410,N_9586);
and U9621 (N_9621,N_9457,N_9374);
or U9622 (N_9622,N_9450,N_9468);
or U9623 (N_9623,N_9412,N_9592);
nand U9624 (N_9624,N_9553,N_9409);
or U9625 (N_9625,N_9339,N_9337);
or U9626 (N_9626,N_9569,N_9373);
or U9627 (N_9627,N_9360,N_9528);
and U9628 (N_9628,N_9300,N_9317);
nand U9629 (N_9629,N_9559,N_9510);
nor U9630 (N_9630,N_9427,N_9459);
nor U9631 (N_9631,N_9513,N_9393);
nor U9632 (N_9632,N_9349,N_9444);
xor U9633 (N_9633,N_9564,N_9599);
nand U9634 (N_9634,N_9413,N_9543);
or U9635 (N_9635,N_9415,N_9426);
and U9636 (N_9636,N_9547,N_9536);
or U9637 (N_9637,N_9396,N_9488);
nor U9638 (N_9638,N_9359,N_9453);
xnor U9639 (N_9639,N_9423,N_9587);
or U9640 (N_9640,N_9509,N_9548);
or U9641 (N_9641,N_9514,N_9470);
nor U9642 (N_9642,N_9542,N_9362);
nand U9643 (N_9643,N_9463,N_9521);
xor U9644 (N_9644,N_9471,N_9538);
nand U9645 (N_9645,N_9473,N_9496);
xnor U9646 (N_9646,N_9340,N_9336);
nor U9647 (N_9647,N_9562,N_9467);
nor U9648 (N_9648,N_9314,N_9558);
or U9649 (N_9649,N_9430,N_9570);
or U9650 (N_9650,N_9367,N_9375);
or U9651 (N_9651,N_9446,N_9478);
nor U9652 (N_9652,N_9310,N_9304);
xnor U9653 (N_9653,N_9485,N_9580);
nor U9654 (N_9654,N_9511,N_9404);
nor U9655 (N_9655,N_9407,N_9437);
xor U9656 (N_9656,N_9321,N_9418);
nor U9657 (N_9657,N_9389,N_9575);
and U9658 (N_9658,N_9567,N_9487);
or U9659 (N_9659,N_9388,N_9400);
or U9660 (N_9660,N_9512,N_9320);
nand U9661 (N_9661,N_9422,N_9454);
and U9662 (N_9662,N_9366,N_9520);
xor U9663 (N_9663,N_9591,N_9577);
xor U9664 (N_9664,N_9489,N_9439);
xnor U9665 (N_9665,N_9476,N_9597);
nor U9666 (N_9666,N_9498,N_9392);
xnor U9667 (N_9667,N_9384,N_9358);
xnor U9668 (N_9668,N_9405,N_9507);
xnor U9669 (N_9669,N_9350,N_9408);
and U9670 (N_9670,N_9395,N_9371);
nor U9671 (N_9671,N_9451,N_9421);
or U9672 (N_9672,N_9369,N_9334);
nand U9673 (N_9673,N_9329,N_9447);
and U9674 (N_9674,N_9305,N_9312);
or U9675 (N_9675,N_9486,N_9589);
nor U9676 (N_9676,N_9398,N_9576);
nor U9677 (N_9677,N_9414,N_9363);
xor U9678 (N_9678,N_9594,N_9331);
or U9679 (N_9679,N_9440,N_9311);
xor U9680 (N_9680,N_9424,N_9560);
and U9681 (N_9681,N_9462,N_9505);
or U9682 (N_9682,N_9325,N_9361);
xor U9683 (N_9683,N_9568,N_9399);
xor U9684 (N_9684,N_9522,N_9573);
xnor U9685 (N_9685,N_9581,N_9555);
xor U9686 (N_9686,N_9434,N_9324);
and U9687 (N_9687,N_9544,N_9531);
xnor U9688 (N_9688,N_9313,N_9347);
or U9689 (N_9689,N_9537,N_9460);
xor U9690 (N_9690,N_9394,N_9355);
xor U9691 (N_9691,N_9365,N_9343);
and U9692 (N_9692,N_9480,N_9376);
or U9693 (N_9693,N_9483,N_9309);
xor U9694 (N_9694,N_9370,N_9332);
and U9695 (N_9695,N_9382,N_9477);
or U9696 (N_9696,N_9308,N_9406);
or U9697 (N_9697,N_9494,N_9518);
nor U9698 (N_9698,N_9529,N_9532);
and U9699 (N_9699,N_9372,N_9333);
and U9700 (N_9700,N_9401,N_9419);
xor U9701 (N_9701,N_9425,N_9351);
nor U9702 (N_9702,N_9533,N_9525);
nor U9703 (N_9703,N_9301,N_9383);
and U9704 (N_9704,N_9306,N_9390);
xor U9705 (N_9705,N_9456,N_9524);
or U9706 (N_9706,N_9403,N_9598);
nor U9707 (N_9707,N_9364,N_9475);
nor U9708 (N_9708,N_9566,N_9432);
nand U9709 (N_9709,N_9443,N_9436);
and U9710 (N_9710,N_9517,N_9315);
nor U9711 (N_9711,N_9550,N_9465);
xnor U9712 (N_9712,N_9484,N_9561);
nand U9713 (N_9713,N_9539,N_9354);
nor U9714 (N_9714,N_9326,N_9344);
nor U9715 (N_9715,N_9495,N_9348);
xor U9716 (N_9716,N_9506,N_9515);
xnor U9717 (N_9717,N_9416,N_9466);
nand U9718 (N_9718,N_9526,N_9357);
or U9719 (N_9719,N_9499,N_9381);
nor U9720 (N_9720,N_9417,N_9452);
xor U9721 (N_9721,N_9346,N_9377);
or U9722 (N_9722,N_9341,N_9368);
nor U9723 (N_9723,N_9378,N_9335);
or U9724 (N_9724,N_9420,N_9481);
nand U9725 (N_9725,N_9554,N_9385);
nand U9726 (N_9726,N_9469,N_9578);
or U9727 (N_9727,N_9318,N_9583);
xor U9728 (N_9728,N_9551,N_9327);
nor U9729 (N_9729,N_9302,N_9428);
or U9730 (N_9730,N_9492,N_9386);
nor U9731 (N_9731,N_9429,N_9519);
nor U9732 (N_9732,N_9574,N_9307);
nand U9733 (N_9733,N_9455,N_9316);
xnor U9734 (N_9734,N_9342,N_9445);
nand U9735 (N_9735,N_9397,N_9523);
and U9736 (N_9736,N_9582,N_9449);
and U9737 (N_9737,N_9323,N_9431);
nand U9738 (N_9738,N_9411,N_9352);
and U9739 (N_9739,N_9557,N_9330);
and U9740 (N_9740,N_9565,N_9379);
xnor U9741 (N_9741,N_9474,N_9438);
xnor U9742 (N_9742,N_9387,N_9590);
nand U9743 (N_9743,N_9391,N_9584);
or U9744 (N_9744,N_9491,N_9322);
nand U9745 (N_9745,N_9516,N_9527);
nand U9746 (N_9746,N_9464,N_9563);
and U9747 (N_9747,N_9501,N_9541);
nor U9748 (N_9748,N_9579,N_9549);
xor U9749 (N_9749,N_9461,N_9303);
nor U9750 (N_9750,N_9328,N_9538);
xor U9751 (N_9751,N_9397,N_9584);
nor U9752 (N_9752,N_9508,N_9369);
and U9753 (N_9753,N_9546,N_9401);
nor U9754 (N_9754,N_9454,N_9582);
and U9755 (N_9755,N_9304,N_9541);
nand U9756 (N_9756,N_9463,N_9406);
xor U9757 (N_9757,N_9380,N_9405);
or U9758 (N_9758,N_9532,N_9443);
nand U9759 (N_9759,N_9443,N_9565);
or U9760 (N_9760,N_9524,N_9354);
or U9761 (N_9761,N_9442,N_9597);
nand U9762 (N_9762,N_9359,N_9539);
nand U9763 (N_9763,N_9558,N_9509);
xor U9764 (N_9764,N_9381,N_9473);
and U9765 (N_9765,N_9409,N_9312);
or U9766 (N_9766,N_9493,N_9554);
or U9767 (N_9767,N_9476,N_9345);
or U9768 (N_9768,N_9413,N_9423);
or U9769 (N_9769,N_9440,N_9580);
or U9770 (N_9770,N_9399,N_9584);
nor U9771 (N_9771,N_9535,N_9446);
nor U9772 (N_9772,N_9329,N_9327);
nor U9773 (N_9773,N_9561,N_9598);
or U9774 (N_9774,N_9343,N_9448);
nor U9775 (N_9775,N_9370,N_9438);
and U9776 (N_9776,N_9375,N_9579);
xor U9777 (N_9777,N_9586,N_9574);
or U9778 (N_9778,N_9384,N_9501);
and U9779 (N_9779,N_9571,N_9452);
nand U9780 (N_9780,N_9331,N_9587);
or U9781 (N_9781,N_9534,N_9500);
and U9782 (N_9782,N_9438,N_9552);
nor U9783 (N_9783,N_9341,N_9581);
nor U9784 (N_9784,N_9492,N_9399);
or U9785 (N_9785,N_9563,N_9381);
xnor U9786 (N_9786,N_9491,N_9358);
or U9787 (N_9787,N_9450,N_9455);
xnor U9788 (N_9788,N_9463,N_9532);
nor U9789 (N_9789,N_9489,N_9305);
nand U9790 (N_9790,N_9563,N_9449);
and U9791 (N_9791,N_9345,N_9587);
nor U9792 (N_9792,N_9366,N_9458);
or U9793 (N_9793,N_9558,N_9446);
xnor U9794 (N_9794,N_9301,N_9579);
xor U9795 (N_9795,N_9382,N_9378);
or U9796 (N_9796,N_9592,N_9347);
and U9797 (N_9797,N_9343,N_9468);
and U9798 (N_9798,N_9405,N_9451);
or U9799 (N_9799,N_9429,N_9574);
and U9800 (N_9800,N_9385,N_9397);
and U9801 (N_9801,N_9384,N_9567);
and U9802 (N_9802,N_9536,N_9433);
nor U9803 (N_9803,N_9386,N_9380);
xnor U9804 (N_9804,N_9570,N_9580);
nand U9805 (N_9805,N_9479,N_9599);
or U9806 (N_9806,N_9509,N_9502);
and U9807 (N_9807,N_9431,N_9430);
xor U9808 (N_9808,N_9487,N_9441);
xnor U9809 (N_9809,N_9333,N_9538);
and U9810 (N_9810,N_9593,N_9566);
nor U9811 (N_9811,N_9401,N_9465);
or U9812 (N_9812,N_9569,N_9566);
and U9813 (N_9813,N_9439,N_9566);
and U9814 (N_9814,N_9417,N_9523);
or U9815 (N_9815,N_9359,N_9549);
or U9816 (N_9816,N_9325,N_9501);
nor U9817 (N_9817,N_9334,N_9498);
and U9818 (N_9818,N_9514,N_9567);
nand U9819 (N_9819,N_9339,N_9465);
and U9820 (N_9820,N_9501,N_9348);
xor U9821 (N_9821,N_9519,N_9441);
nor U9822 (N_9822,N_9581,N_9597);
or U9823 (N_9823,N_9359,N_9567);
nand U9824 (N_9824,N_9411,N_9343);
and U9825 (N_9825,N_9596,N_9394);
xnor U9826 (N_9826,N_9575,N_9362);
or U9827 (N_9827,N_9455,N_9564);
nand U9828 (N_9828,N_9465,N_9543);
or U9829 (N_9829,N_9582,N_9520);
and U9830 (N_9830,N_9553,N_9477);
and U9831 (N_9831,N_9481,N_9453);
xor U9832 (N_9832,N_9507,N_9546);
and U9833 (N_9833,N_9339,N_9426);
or U9834 (N_9834,N_9567,N_9430);
xnor U9835 (N_9835,N_9438,N_9349);
and U9836 (N_9836,N_9378,N_9372);
and U9837 (N_9837,N_9443,N_9467);
xnor U9838 (N_9838,N_9584,N_9362);
nand U9839 (N_9839,N_9338,N_9483);
nor U9840 (N_9840,N_9501,N_9344);
xnor U9841 (N_9841,N_9356,N_9465);
and U9842 (N_9842,N_9577,N_9499);
nand U9843 (N_9843,N_9352,N_9343);
nand U9844 (N_9844,N_9497,N_9406);
nor U9845 (N_9845,N_9434,N_9323);
nand U9846 (N_9846,N_9443,N_9360);
nand U9847 (N_9847,N_9587,N_9336);
nand U9848 (N_9848,N_9522,N_9536);
and U9849 (N_9849,N_9336,N_9427);
nand U9850 (N_9850,N_9403,N_9323);
nand U9851 (N_9851,N_9599,N_9485);
and U9852 (N_9852,N_9378,N_9448);
xnor U9853 (N_9853,N_9474,N_9564);
and U9854 (N_9854,N_9596,N_9308);
nand U9855 (N_9855,N_9465,N_9482);
nand U9856 (N_9856,N_9434,N_9355);
xnor U9857 (N_9857,N_9451,N_9351);
and U9858 (N_9858,N_9489,N_9313);
and U9859 (N_9859,N_9503,N_9452);
xnor U9860 (N_9860,N_9320,N_9591);
nor U9861 (N_9861,N_9377,N_9528);
or U9862 (N_9862,N_9429,N_9315);
nor U9863 (N_9863,N_9333,N_9465);
and U9864 (N_9864,N_9386,N_9496);
nand U9865 (N_9865,N_9516,N_9433);
xnor U9866 (N_9866,N_9320,N_9492);
nand U9867 (N_9867,N_9424,N_9322);
xnor U9868 (N_9868,N_9463,N_9530);
or U9869 (N_9869,N_9504,N_9350);
or U9870 (N_9870,N_9435,N_9497);
nand U9871 (N_9871,N_9544,N_9301);
nand U9872 (N_9872,N_9391,N_9301);
nor U9873 (N_9873,N_9503,N_9515);
xor U9874 (N_9874,N_9540,N_9508);
or U9875 (N_9875,N_9462,N_9314);
nand U9876 (N_9876,N_9469,N_9580);
nand U9877 (N_9877,N_9331,N_9591);
and U9878 (N_9878,N_9441,N_9488);
nor U9879 (N_9879,N_9362,N_9598);
xor U9880 (N_9880,N_9307,N_9398);
and U9881 (N_9881,N_9410,N_9569);
xor U9882 (N_9882,N_9461,N_9457);
nand U9883 (N_9883,N_9370,N_9506);
xor U9884 (N_9884,N_9483,N_9514);
or U9885 (N_9885,N_9562,N_9389);
xnor U9886 (N_9886,N_9593,N_9444);
or U9887 (N_9887,N_9349,N_9319);
nor U9888 (N_9888,N_9302,N_9344);
xnor U9889 (N_9889,N_9404,N_9583);
or U9890 (N_9890,N_9358,N_9578);
or U9891 (N_9891,N_9541,N_9487);
nand U9892 (N_9892,N_9518,N_9346);
nand U9893 (N_9893,N_9424,N_9440);
or U9894 (N_9894,N_9510,N_9367);
nand U9895 (N_9895,N_9393,N_9361);
nor U9896 (N_9896,N_9417,N_9441);
xnor U9897 (N_9897,N_9550,N_9510);
xnor U9898 (N_9898,N_9480,N_9577);
xor U9899 (N_9899,N_9486,N_9563);
or U9900 (N_9900,N_9830,N_9744);
and U9901 (N_9901,N_9653,N_9606);
nor U9902 (N_9902,N_9674,N_9834);
nand U9903 (N_9903,N_9784,N_9721);
and U9904 (N_9904,N_9607,N_9665);
nand U9905 (N_9905,N_9732,N_9820);
xor U9906 (N_9906,N_9873,N_9673);
and U9907 (N_9907,N_9899,N_9775);
or U9908 (N_9908,N_9745,N_9838);
and U9909 (N_9909,N_9779,N_9773);
and U9910 (N_9910,N_9859,N_9614);
and U9911 (N_9911,N_9660,N_9648);
nor U9912 (N_9912,N_9768,N_9608);
and U9913 (N_9913,N_9646,N_9624);
nor U9914 (N_9914,N_9778,N_9839);
and U9915 (N_9915,N_9726,N_9875);
xnor U9916 (N_9916,N_9605,N_9704);
xor U9917 (N_9917,N_9831,N_9833);
nand U9918 (N_9918,N_9742,N_9749);
xor U9919 (N_9919,N_9853,N_9652);
and U9920 (N_9920,N_9626,N_9857);
nor U9921 (N_9921,N_9639,N_9752);
nor U9922 (N_9922,N_9891,N_9601);
nor U9923 (N_9923,N_9856,N_9709);
nor U9924 (N_9924,N_9881,N_9609);
and U9925 (N_9925,N_9718,N_9808);
and U9926 (N_9926,N_9724,N_9731);
nand U9927 (N_9927,N_9789,N_9885);
nor U9928 (N_9928,N_9656,N_9889);
nor U9929 (N_9929,N_9781,N_9760);
and U9930 (N_9930,N_9753,N_9854);
nor U9931 (N_9931,N_9705,N_9818);
nand U9932 (N_9932,N_9659,N_9793);
nand U9933 (N_9933,N_9620,N_9851);
nor U9934 (N_9934,N_9879,N_9611);
nor U9935 (N_9935,N_9772,N_9880);
nor U9936 (N_9936,N_9681,N_9668);
nand U9937 (N_9937,N_9628,N_9827);
nor U9938 (N_9938,N_9806,N_9671);
or U9939 (N_9939,N_9612,N_9619);
xor U9940 (N_9940,N_9877,N_9603);
or U9941 (N_9941,N_9722,N_9600);
nor U9942 (N_9942,N_9865,N_9675);
and U9943 (N_9943,N_9822,N_9643);
xor U9944 (N_9944,N_9819,N_9888);
and U9945 (N_9945,N_9890,N_9637);
nand U9946 (N_9946,N_9746,N_9871);
nand U9947 (N_9947,N_9698,N_9622);
nor U9948 (N_9948,N_9625,N_9751);
nand U9949 (N_9949,N_9706,N_9848);
nor U9950 (N_9950,N_9733,N_9790);
xor U9951 (N_9951,N_9780,N_9798);
nand U9952 (N_9952,N_9862,N_9821);
and U9953 (N_9953,N_9767,N_9774);
and U9954 (N_9954,N_9739,N_9644);
xnor U9955 (N_9955,N_9777,N_9747);
nand U9956 (N_9956,N_9736,N_9633);
nor U9957 (N_9957,N_9869,N_9863);
xor U9958 (N_9958,N_9641,N_9812);
or U9959 (N_9959,N_9743,N_9876);
or U9960 (N_9960,N_9766,N_9765);
and U9961 (N_9961,N_9723,N_9898);
nor U9962 (N_9962,N_9850,N_9682);
and U9963 (N_9963,N_9623,N_9713);
and U9964 (N_9964,N_9826,N_9651);
nor U9965 (N_9965,N_9823,N_9796);
nor U9966 (N_9966,N_9693,N_9680);
nand U9967 (N_9967,N_9791,N_9759);
and U9968 (N_9968,N_9836,N_9740);
nor U9969 (N_9969,N_9769,N_9717);
and U9970 (N_9970,N_9844,N_9701);
or U9971 (N_9971,N_9874,N_9832);
and U9972 (N_9972,N_9642,N_9800);
xor U9973 (N_9973,N_9632,N_9810);
xnor U9974 (N_9974,N_9697,N_9692);
nor U9975 (N_9975,N_9776,N_9720);
or U9976 (N_9976,N_9686,N_9663);
and U9977 (N_9977,N_9610,N_9689);
and U9978 (N_9978,N_9734,N_9771);
nor U9979 (N_9979,N_9829,N_9728);
nor U9980 (N_9980,N_9634,N_9758);
xnor U9981 (N_9981,N_9896,N_9841);
nand U9982 (N_9982,N_9866,N_9893);
and U9983 (N_9983,N_9664,N_9615);
nand U9984 (N_9984,N_9761,N_9755);
nand U9985 (N_9985,N_9762,N_9636);
nand U9986 (N_9986,N_9868,N_9645);
xor U9987 (N_9987,N_9696,N_9757);
or U9988 (N_9988,N_9878,N_9799);
and U9989 (N_9989,N_9805,N_9657);
nand U9990 (N_9990,N_9811,N_9691);
or U9991 (N_9991,N_9617,N_9792);
xnor U9992 (N_9992,N_9785,N_9687);
nand U9993 (N_9993,N_9788,N_9662);
and U9994 (N_9994,N_9654,N_9802);
xnor U9995 (N_9995,N_9883,N_9700);
nand U9996 (N_9996,N_9695,N_9770);
or U9997 (N_9997,N_9685,N_9794);
nand U9998 (N_9998,N_9658,N_9630);
or U9999 (N_9999,N_9725,N_9864);
or U10000 (N_10000,N_9678,N_9787);
nor U10001 (N_10001,N_9892,N_9649);
nor U10002 (N_10002,N_9647,N_9825);
nor U10003 (N_10003,N_9707,N_9714);
and U10004 (N_10004,N_9631,N_9764);
xnor U10005 (N_10005,N_9809,N_9886);
nand U10006 (N_10006,N_9884,N_9702);
nand U10007 (N_10007,N_9688,N_9824);
or U10008 (N_10008,N_9872,N_9640);
nand U10009 (N_10009,N_9783,N_9710);
or U10010 (N_10010,N_9801,N_9754);
and U10011 (N_10011,N_9894,N_9737);
nor U10012 (N_10012,N_9795,N_9711);
nand U10013 (N_10013,N_9679,N_9699);
and U10014 (N_10014,N_9694,N_9703);
nand U10015 (N_10015,N_9661,N_9672);
and U10016 (N_10016,N_9855,N_9719);
and U10017 (N_10017,N_9627,N_9815);
and U10018 (N_10018,N_9803,N_9715);
xor U10019 (N_10019,N_9604,N_9667);
and U10020 (N_10020,N_9716,N_9750);
nor U10021 (N_10021,N_9816,N_9756);
nor U10022 (N_10022,N_9729,N_9676);
xnor U10023 (N_10023,N_9813,N_9828);
or U10024 (N_10024,N_9748,N_9895);
or U10025 (N_10025,N_9861,N_9735);
or U10026 (N_10026,N_9613,N_9741);
nand U10027 (N_10027,N_9860,N_9655);
and U10028 (N_10028,N_9817,N_9616);
nand U10029 (N_10029,N_9786,N_9708);
nand U10030 (N_10030,N_9814,N_9621);
or U10031 (N_10031,N_9763,N_9840);
and U10032 (N_10032,N_9669,N_9837);
or U10033 (N_10033,N_9835,N_9797);
or U10034 (N_10034,N_9677,N_9635);
nand U10035 (N_10035,N_9852,N_9629);
xor U10036 (N_10036,N_9738,N_9849);
nand U10037 (N_10037,N_9602,N_9804);
nor U10038 (N_10038,N_9670,N_9727);
nand U10039 (N_10039,N_9867,N_9684);
nand U10040 (N_10040,N_9842,N_9712);
or U10041 (N_10041,N_9882,N_9650);
or U10042 (N_10042,N_9845,N_9638);
or U10043 (N_10043,N_9730,N_9858);
xnor U10044 (N_10044,N_9887,N_9666);
nor U10045 (N_10045,N_9847,N_9870);
nor U10046 (N_10046,N_9897,N_9690);
nand U10047 (N_10047,N_9843,N_9807);
nor U10048 (N_10048,N_9618,N_9782);
and U10049 (N_10049,N_9846,N_9683);
xnor U10050 (N_10050,N_9728,N_9671);
nor U10051 (N_10051,N_9603,N_9756);
nor U10052 (N_10052,N_9738,N_9892);
and U10053 (N_10053,N_9870,N_9635);
nor U10054 (N_10054,N_9685,N_9762);
nor U10055 (N_10055,N_9807,N_9671);
xnor U10056 (N_10056,N_9662,N_9647);
or U10057 (N_10057,N_9763,N_9829);
nor U10058 (N_10058,N_9730,N_9744);
nand U10059 (N_10059,N_9836,N_9882);
nand U10060 (N_10060,N_9807,N_9610);
xnor U10061 (N_10061,N_9871,N_9769);
nor U10062 (N_10062,N_9832,N_9643);
nor U10063 (N_10063,N_9692,N_9833);
and U10064 (N_10064,N_9613,N_9894);
nor U10065 (N_10065,N_9707,N_9698);
and U10066 (N_10066,N_9707,N_9618);
xor U10067 (N_10067,N_9718,N_9892);
xnor U10068 (N_10068,N_9668,N_9608);
xnor U10069 (N_10069,N_9746,N_9798);
nor U10070 (N_10070,N_9608,N_9869);
or U10071 (N_10071,N_9801,N_9600);
nor U10072 (N_10072,N_9639,N_9831);
nand U10073 (N_10073,N_9733,N_9847);
and U10074 (N_10074,N_9801,N_9647);
or U10075 (N_10075,N_9654,N_9602);
nor U10076 (N_10076,N_9681,N_9601);
nand U10077 (N_10077,N_9875,N_9723);
xor U10078 (N_10078,N_9643,N_9636);
nand U10079 (N_10079,N_9617,N_9623);
nor U10080 (N_10080,N_9717,N_9709);
nand U10081 (N_10081,N_9714,N_9896);
or U10082 (N_10082,N_9848,N_9755);
or U10083 (N_10083,N_9655,N_9785);
or U10084 (N_10084,N_9645,N_9723);
or U10085 (N_10085,N_9604,N_9727);
nand U10086 (N_10086,N_9678,N_9893);
or U10087 (N_10087,N_9877,N_9711);
and U10088 (N_10088,N_9791,N_9824);
nand U10089 (N_10089,N_9845,N_9841);
nand U10090 (N_10090,N_9673,N_9774);
or U10091 (N_10091,N_9892,N_9836);
nor U10092 (N_10092,N_9677,N_9762);
or U10093 (N_10093,N_9740,N_9787);
and U10094 (N_10094,N_9605,N_9655);
or U10095 (N_10095,N_9777,N_9629);
xnor U10096 (N_10096,N_9708,N_9703);
nor U10097 (N_10097,N_9602,N_9857);
nor U10098 (N_10098,N_9786,N_9650);
or U10099 (N_10099,N_9667,N_9813);
nand U10100 (N_10100,N_9856,N_9722);
nand U10101 (N_10101,N_9762,N_9852);
or U10102 (N_10102,N_9855,N_9780);
nor U10103 (N_10103,N_9755,N_9849);
nor U10104 (N_10104,N_9639,N_9769);
or U10105 (N_10105,N_9854,N_9799);
xnor U10106 (N_10106,N_9773,N_9656);
xor U10107 (N_10107,N_9611,N_9704);
nand U10108 (N_10108,N_9704,N_9869);
or U10109 (N_10109,N_9786,N_9717);
or U10110 (N_10110,N_9804,N_9610);
nand U10111 (N_10111,N_9847,N_9609);
xor U10112 (N_10112,N_9883,N_9888);
nor U10113 (N_10113,N_9817,N_9768);
nor U10114 (N_10114,N_9801,N_9744);
xor U10115 (N_10115,N_9628,N_9826);
or U10116 (N_10116,N_9715,N_9613);
nor U10117 (N_10117,N_9843,N_9623);
and U10118 (N_10118,N_9895,N_9609);
xnor U10119 (N_10119,N_9656,N_9645);
and U10120 (N_10120,N_9790,N_9873);
nand U10121 (N_10121,N_9623,N_9639);
and U10122 (N_10122,N_9745,N_9613);
nor U10123 (N_10123,N_9814,N_9742);
or U10124 (N_10124,N_9856,N_9837);
and U10125 (N_10125,N_9625,N_9699);
xnor U10126 (N_10126,N_9613,N_9820);
nand U10127 (N_10127,N_9726,N_9818);
nor U10128 (N_10128,N_9767,N_9724);
nand U10129 (N_10129,N_9649,N_9612);
or U10130 (N_10130,N_9606,N_9752);
nor U10131 (N_10131,N_9827,N_9812);
or U10132 (N_10132,N_9678,N_9638);
nor U10133 (N_10133,N_9611,N_9603);
or U10134 (N_10134,N_9863,N_9894);
or U10135 (N_10135,N_9662,N_9862);
or U10136 (N_10136,N_9890,N_9835);
or U10137 (N_10137,N_9835,N_9810);
xor U10138 (N_10138,N_9897,N_9644);
xor U10139 (N_10139,N_9699,N_9787);
and U10140 (N_10140,N_9728,N_9709);
and U10141 (N_10141,N_9854,N_9694);
or U10142 (N_10142,N_9769,N_9622);
or U10143 (N_10143,N_9741,N_9670);
and U10144 (N_10144,N_9734,N_9819);
or U10145 (N_10145,N_9726,N_9774);
or U10146 (N_10146,N_9803,N_9851);
nor U10147 (N_10147,N_9675,N_9711);
xnor U10148 (N_10148,N_9650,N_9654);
nor U10149 (N_10149,N_9632,N_9739);
and U10150 (N_10150,N_9810,N_9720);
xor U10151 (N_10151,N_9722,N_9737);
or U10152 (N_10152,N_9679,N_9844);
and U10153 (N_10153,N_9859,N_9690);
or U10154 (N_10154,N_9805,N_9754);
xnor U10155 (N_10155,N_9743,N_9872);
or U10156 (N_10156,N_9795,N_9857);
and U10157 (N_10157,N_9737,N_9800);
or U10158 (N_10158,N_9702,N_9640);
and U10159 (N_10159,N_9607,N_9658);
xnor U10160 (N_10160,N_9776,N_9820);
and U10161 (N_10161,N_9681,N_9622);
nand U10162 (N_10162,N_9824,N_9836);
and U10163 (N_10163,N_9668,N_9855);
xor U10164 (N_10164,N_9831,N_9699);
nor U10165 (N_10165,N_9814,N_9701);
and U10166 (N_10166,N_9840,N_9893);
and U10167 (N_10167,N_9757,N_9838);
or U10168 (N_10168,N_9898,N_9678);
nor U10169 (N_10169,N_9766,N_9882);
or U10170 (N_10170,N_9657,N_9643);
and U10171 (N_10171,N_9795,N_9785);
nor U10172 (N_10172,N_9646,N_9774);
nand U10173 (N_10173,N_9888,N_9689);
nor U10174 (N_10174,N_9805,N_9618);
nand U10175 (N_10175,N_9672,N_9740);
nor U10176 (N_10176,N_9688,N_9764);
nor U10177 (N_10177,N_9662,N_9779);
nor U10178 (N_10178,N_9801,N_9852);
or U10179 (N_10179,N_9772,N_9864);
xor U10180 (N_10180,N_9614,N_9632);
or U10181 (N_10181,N_9633,N_9637);
and U10182 (N_10182,N_9629,N_9871);
or U10183 (N_10183,N_9780,N_9838);
or U10184 (N_10184,N_9776,N_9861);
and U10185 (N_10185,N_9719,N_9889);
and U10186 (N_10186,N_9692,N_9776);
nand U10187 (N_10187,N_9833,N_9863);
nor U10188 (N_10188,N_9638,N_9760);
or U10189 (N_10189,N_9882,N_9792);
nand U10190 (N_10190,N_9604,N_9617);
nand U10191 (N_10191,N_9794,N_9688);
nand U10192 (N_10192,N_9892,N_9818);
nand U10193 (N_10193,N_9771,N_9650);
and U10194 (N_10194,N_9806,N_9664);
and U10195 (N_10195,N_9748,N_9654);
or U10196 (N_10196,N_9698,N_9652);
nand U10197 (N_10197,N_9632,N_9751);
and U10198 (N_10198,N_9697,N_9734);
xnor U10199 (N_10199,N_9710,N_9834);
and U10200 (N_10200,N_9913,N_10094);
nand U10201 (N_10201,N_10174,N_9954);
nor U10202 (N_10202,N_9985,N_9973);
nor U10203 (N_10203,N_9927,N_9959);
nor U10204 (N_10204,N_9990,N_10019);
nor U10205 (N_10205,N_10012,N_10099);
or U10206 (N_10206,N_10148,N_9991);
and U10207 (N_10207,N_10028,N_10044);
or U10208 (N_10208,N_10147,N_10186);
and U10209 (N_10209,N_10056,N_9997);
or U10210 (N_10210,N_10071,N_10022);
and U10211 (N_10211,N_10198,N_10140);
or U10212 (N_10212,N_9999,N_10087);
nor U10213 (N_10213,N_9917,N_10045);
xor U10214 (N_10214,N_10093,N_10073);
nor U10215 (N_10215,N_9958,N_10164);
xnor U10216 (N_10216,N_10014,N_9907);
xnor U10217 (N_10217,N_10064,N_10116);
and U10218 (N_10218,N_10163,N_10033);
or U10219 (N_10219,N_10095,N_9919);
nand U10220 (N_10220,N_10016,N_9933);
or U10221 (N_10221,N_10050,N_10107);
nand U10222 (N_10222,N_10021,N_10180);
and U10223 (N_10223,N_9974,N_9949);
nor U10224 (N_10224,N_9928,N_10039);
and U10225 (N_10225,N_9980,N_10066);
xnor U10226 (N_10226,N_9969,N_10126);
or U10227 (N_10227,N_9916,N_10146);
nor U10228 (N_10228,N_9937,N_9902);
xnor U10229 (N_10229,N_10196,N_10058);
or U10230 (N_10230,N_9951,N_10030);
or U10231 (N_10231,N_9940,N_10134);
nand U10232 (N_10232,N_10122,N_9998);
nand U10233 (N_10233,N_9978,N_10139);
xnor U10234 (N_10234,N_9956,N_9979);
or U10235 (N_10235,N_10067,N_10111);
nor U10236 (N_10236,N_10136,N_9924);
xor U10237 (N_10237,N_9987,N_10157);
xor U10238 (N_10238,N_10104,N_10096);
or U10239 (N_10239,N_10143,N_10042);
and U10240 (N_10240,N_10190,N_9950);
or U10241 (N_10241,N_10158,N_10061);
nand U10242 (N_10242,N_10070,N_10031);
nand U10243 (N_10243,N_9915,N_9934);
and U10244 (N_10244,N_10057,N_10117);
and U10245 (N_10245,N_10091,N_9909);
or U10246 (N_10246,N_10118,N_10151);
and U10247 (N_10247,N_10000,N_9925);
or U10248 (N_10248,N_9962,N_10176);
or U10249 (N_10249,N_10131,N_10006);
nand U10250 (N_10250,N_10130,N_10048);
or U10251 (N_10251,N_10038,N_10152);
and U10252 (N_10252,N_10034,N_10159);
and U10253 (N_10253,N_10185,N_10055);
or U10254 (N_10254,N_10177,N_10098);
nor U10255 (N_10255,N_10053,N_10032);
xor U10256 (N_10256,N_10110,N_9994);
nand U10257 (N_10257,N_10179,N_10109);
nand U10258 (N_10258,N_10154,N_10144);
or U10259 (N_10259,N_10193,N_10009);
or U10260 (N_10260,N_9921,N_10029);
nand U10261 (N_10261,N_10170,N_10085);
nand U10262 (N_10262,N_9929,N_10052);
or U10263 (N_10263,N_9918,N_10079);
xor U10264 (N_10264,N_9992,N_9977);
or U10265 (N_10265,N_10003,N_10168);
nand U10266 (N_10266,N_9944,N_9955);
or U10267 (N_10267,N_9935,N_10089);
nand U10268 (N_10268,N_10020,N_9904);
xnor U10269 (N_10269,N_10069,N_10119);
xnor U10270 (N_10270,N_9906,N_10043);
and U10271 (N_10271,N_9983,N_9926);
xor U10272 (N_10272,N_10138,N_9961);
nand U10273 (N_10273,N_10171,N_10083);
nand U10274 (N_10274,N_9981,N_9900);
nor U10275 (N_10275,N_10023,N_10128);
nand U10276 (N_10276,N_10187,N_9922);
or U10277 (N_10277,N_10125,N_10063);
nand U10278 (N_10278,N_9914,N_10194);
or U10279 (N_10279,N_9975,N_10124);
nor U10280 (N_10280,N_9931,N_10133);
xnor U10281 (N_10281,N_10082,N_9930);
nor U10282 (N_10282,N_10051,N_9988);
nand U10283 (N_10283,N_10097,N_10184);
xnor U10284 (N_10284,N_10035,N_10054);
nor U10285 (N_10285,N_10165,N_10153);
xnor U10286 (N_10286,N_10068,N_10047);
or U10287 (N_10287,N_10175,N_10004);
or U10288 (N_10288,N_10199,N_10017);
nor U10289 (N_10289,N_9972,N_9982);
or U10290 (N_10290,N_9963,N_10080);
xor U10291 (N_10291,N_9957,N_10182);
nor U10292 (N_10292,N_10167,N_10007);
and U10293 (N_10293,N_9905,N_9976);
and U10294 (N_10294,N_9901,N_10013);
and U10295 (N_10295,N_10018,N_10002);
xnor U10296 (N_10296,N_9911,N_10191);
nor U10297 (N_10297,N_10145,N_10195);
xor U10298 (N_10298,N_10076,N_10041);
and U10299 (N_10299,N_10011,N_10060);
or U10300 (N_10300,N_10075,N_10059);
nand U10301 (N_10301,N_9966,N_10114);
nor U10302 (N_10302,N_9923,N_10001);
xor U10303 (N_10303,N_10188,N_10142);
nor U10304 (N_10304,N_10166,N_10072);
nand U10305 (N_10305,N_10172,N_10027);
nand U10306 (N_10306,N_10156,N_10077);
xnor U10307 (N_10307,N_10189,N_10160);
and U10308 (N_10308,N_9953,N_9971);
nand U10309 (N_10309,N_10049,N_10015);
nor U10310 (N_10310,N_9989,N_10155);
nor U10311 (N_10311,N_10008,N_9947);
or U10312 (N_10312,N_10025,N_10137);
xnor U10313 (N_10313,N_10103,N_9938);
nand U10314 (N_10314,N_9995,N_10120);
or U10315 (N_10315,N_9932,N_10112);
xor U10316 (N_10316,N_10105,N_9920);
and U10317 (N_10317,N_9996,N_10086);
xnor U10318 (N_10318,N_10183,N_10169);
xor U10319 (N_10319,N_10115,N_9939);
nand U10320 (N_10320,N_9912,N_9968);
nand U10321 (N_10321,N_9946,N_10081);
nor U10322 (N_10322,N_10100,N_9970);
and U10323 (N_10323,N_10101,N_9908);
or U10324 (N_10324,N_9910,N_10102);
xor U10325 (N_10325,N_9960,N_9964);
or U10326 (N_10326,N_10040,N_10161);
or U10327 (N_10327,N_9967,N_9936);
xnor U10328 (N_10328,N_10123,N_10065);
xor U10329 (N_10329,N_10127,N_9942);
or U10330 (N_10330,N_10197,N_10005);
xor U10331 (N_10331,N_10192,N_9984);
nand U10332 (N_10332,N_10178,N_10010);
or U10333 (N_10333,N_10132,N_9943);
xor U10334 (N_10334,N_9986,N_9965);
nand U10335 (N_10335,N_10162,N_10037);
nand U10336 (N_10336,N_10036,N_9948);
or U10337 (N_10337,N_10046,N_10121);
and U10338 (N_10338,N_9945,N_10150);
or U10339 (N_10339,N_10149,N_9903);
and U10340 (N_10340,N_10181,N_10084);
nor U10341 (N_10341,N_10088,N_10090);
nand U10342 (N_10342,N_10092,N_10078);
xor U10343 (N_10343,N_10173,N_10074);
and U10344 (N_10344,N_10135,N_10062);
nor U10345 (N_10345,N_9993,N_10113);
nand U10346 (N_10346,N_10129,N_10108);
xnor U10347 (N_10347,N_10106,N_10024);
or U10348 (N_10348,N_9952,N_10026);
and U10349 (N_10349,N_10141,N_9941);
nor U10350 (N_10350,N_9923,N_10098);
nand U10351 (N_10351,N_9986,N_9915);
or U10352 (N_10352,N_9996,N_9986);
xor U10353 (N_10353,N_10158,N_10132);
nor U10354 (N_10354,N_10012,N_10063);
nor U10355 (N_10355,N_10002,N_10023);
nor U10356 (N_10356,N_10147,N_9928);
or U10357 (N_10357,N_10199,N_10028);
nand U10358 (N_10358,N_10013,N_10158);
or U10359 (N_10359,N_10091,N_9930);
nor U10360 (N_10360,N_10126,N_10133);
nor U10361 (N_10361,N_9976,N_10118);
or U10362 (N_10362,N_9983,N_10107);
or U10363 (N_10363,N_10013,N_9939);
nor U10364 (N_10364,N_10024,N_9970);
nand U10365 (N_10365,N_10167,N_10111);
nor U10366 (N_10366,N_9935,N_9970);
xnor U10367 (N_10367,N_10030,N_9914);
and U10368 (N_10368,N_10017,N_10085);
or U10369 (N_10369,N_10050,N_10102);
nor U10370 (N_10370,N_10197,N_10161);
nor U10371 (N_10371,N_10072,N_10164);
xor U10372 (N_10372,N_10089,N_10050);
xor U10373 (N_10373,N_9916,N_9901);
xor U10374 (N_10374,N_10164,N_10033);
nor U10375 (N_10375,N_10102,N_10092);
nor U10376 (N_10376,N_9911,N_10171);
nor U10377 (N_10377,N_9932,N_10115);
nand U10378 (N_10378,N_10085,N_10052);
xor U10379 (N_10379,N_9926,N_10145);
and U10380 (N_10380,N_9967,N_10158);
or U10381 (N_10381,N_10129,N_10089);
nor U10382 (N_10382,N_10092,N_9945);
and U10383 (N_10383,N_10002,N_9966);
nor U10384 (N_10384,N_10037,N_10171);
nand U10385 (N_10385,N_10042,N_10080);
xor U10386 (N_10386,N_9969,N_10054);
xor U10387 (N_10387,N_10163,N_10115);
or U10388 (N_10388,N_10016,N_10061);
xor U10389 (N_10389,N_10092,N_9991);
or U10390 (N_10390,N_10162,N_9934);
and U10391 (N_10391,N_9941,N_9992);
nand U10392 (N_10392,N_10142,N_9952);
xor U10393 (N_10393,N_9903,N_10159);
nor U10394 (N_10394,N_9971,N_10045);
nand U10395 (N_10395,N_10033,N_10115);
or U10396 (N_10396,N_10129,N_10094);
nor U10397 (N_10397,N_9925,N_10078);
and U10398 (N_10398,N_10096,N_10144);
or U10399 (N_10399,N_10165,N_9956);
or U10400 (N_10400,N_9927,N_10168);
nor U10401 (N_10401,N_9949,N_9934);
nand U10402 (N_10402,N_10128,N_9917);
nor U10403 (N_10403,N_9974,N_9950);
or U10404 (N_10404,N_10122,N_10059);
nand U10405 (N_10405,N_9916,N_9997);
nand U10406 (N_10406,N_9998,N_9912);
and U10407 (N_10407,N_10193,N_10166);
nor U10408 (N_10408,N_10104,N_9919);
and U10409 (N_10409,N_10076,N_10176);
or U10410 (N_10410,N_10054,N_9963);
nor U10411 (N_10411,N_10045,N_10019);
nand U10412 (N_10412,N_10009,N_10097);
xor U10413 (N_10413,N_9976,N_10035);
nand U10414 (N_10414,N_9945,N_10001);
nand U10415 (N_10415,N_9977,N_9928);
nor U10416 (N_10416,N_10152,N_10181);
nor U10417 (N_10417,N_10159,N_10058);
or U10418 (N_10418,N_10027,N_10042);
nor U10419 (N_10419,N_9930,N_10094);
or U10420 (N_10420,N_9939,N_9936);
xor U10421 (N_10421,N_10052,N_10093);
nand U10422 (N_10422,N_10066,N_10082);
nand U10423 (N_10423,N_10193,N_9945);
xor U10424 (N_10424,N_10141,N_9940);
xor U10425 (N_10425,N_10029,N_10097);
xor U10426 (N_10426,N_9904,N_10008);
and U10427 (N_10427,N_10106,N_10179);
and U10428 (N_10428,N_10147,N_9917);
nand U10429 (N_10429,N_9957,N_10014);
nor U10430 (N_10430,N_10127,N_10059);
or U10431 (N_10431,N_10075,N_10159);
and U10432 (N_10432,N_10161,N_10162);
or U10433 (N_10433,N_10046,N_10116);
xnor U10434 (N_10434,N_9943,N_9957);
xnor U10435 (N_10435,N_10192,N_10150);
nand U10436 (N_10436,N_10049,N_10178);
xor U10437 (N_10437,N_10165,N_9913);
nand U10438 (N_10438,N_9933,N_10073);
xor U10439 (N_10439,N_10043,N_9909);
or U10440 (N_10440,N_10126,N_10106);
xor U10441 (N_10441,N_10019,N_10117);
nand U10442 (N_10442,N_9943,N_10139);
or U10443 (N_10443,N_10098,N_10112);
nor U10444 (N_10444,N_10179,N_10167);
nor U10445 (N_10445,N_10086,N_10040);
or U10446 (N_10446,N_9917,N_10056);
or U10447 (N_10447,N_9957,N_10097);
and U10448 (N_10448,N_10139,N_10135);
or U10449 (N_10449,N_9941,N_9970);
nor U10450 (N_10450,N_10108,N_10193);
nor U10451 (N_10451,N_10115,N_10109);
and U10452 (N_10452,N_10060,N_9976);
nor U10453 (N_10453,N_9926,N_10075);
and U10454 (N_10454,N_10134,N_10073);
xor U10455 (N_10455,N_10154,N_10109);
and U10456 (N_10456,N_9988,N_10002);
nand U10457 (N_10457,N_10163,N_10018);
and U10458 (N_10458,N_9964,N_9914);
or U10459 (N_10459,N_10008,N_9967);
nand U10460 (N_10460,N_10022,N_10111);
nand U10461 (N_10461,N_10182,N_9968);
xor U10462 (N_10462,N_10073,N_9905);
nor U10463 (N_10463,N_10172,N_10093);
nor U10464 (N_10464,N_9953,N_9974);
xor U10465 (N_10465,N_9933,N_10069);
nand U10466 (N_10466,N_9924,N_10031);
nand U10467 (N_10467,N_10196,N_10022);
xnor U10468 (N_10468,N_9922,N_9933);
nor U10469 (N_10469,N_9948,N_9915);
and U10470 (N_10470,N_10162,N_10065);
or U10471 (N_10471,N_10156,N_10192);
and U10472 (N_10472,N_10129,N_10023);
and U10473 (N_10473,N_10076,N_10100);
and U10474 (N_10474,N_9974,N_9978);
nand U10475 (N_10475,N_10170,N_9960);
xnor U10476 (N_10476,N_10008,N_9938);
xor U10477 (N_10477,N_10043,N_10085);
nand U10478 (N_10478,N_10103,N_10060);
nand U10479 (N_10479,N_9995,N_10137);
xor U10480 (N_10480,N_10037,N_10091);
and U10481 (N_10481,N_10004,N_10053);
or U10482 (N_10482,N_10061,N_10002);
or U10483 (N_10483,N_10151,N_9907);
and U10484 (N_10484,N_9983,N_10160);
xor U10485 (N_10485,N_9987,N_10093);
nor U10486 (N_10486,N_9998,N_9993);
or U10487 (N_10487,N_10167,N_9902);
or U10488 (N_10488,N_9908,N_10176);
and U10489 (N_10489,N_10066,N_10056);
xnor U10490 (N_10490,N_10196,N_10160);
xor U10491 (N_10491,N_10045,N_9955);
or U10492 (N_10492,N_10090,N_10035);
nand U10493 (N_10493,N_10190,N_10125);
xor U10494 (N_10494,N_10147,N_10156);
xor U10495 (N_10495,N_9917,N_10008);
nand U10496 (N_10496,N_10023,N_10082);
xor U10497 (N_10497,N_10085,N_10126);
nor U10498 (N_10498,N_10051,N_10042);
nand U10499 (N_10499,N_9933,N_10049);
or U10500 (N_10500,N_10212,N_10272);
xor U10501 (N_10501,N_10357,N_10391);
xor U10502 (N_10502,N_10288,N_10316);
xnor U10503 (N_10503,N_10482,N_10282);
nor U10504 (N_10504,N_10224,N_10378);
or U10505 (N_10505,N_10325,N_10499);
nand U10506 (N_10506,N_10445,N_10351);
xor U10507 (N_10507,N_10238,N_10225);
nand U10508 (N_10508,N_10363,N_10240);
xor U10509 (N_10509,N_10346,N_10490);
or U10510 (N_10510,N_10323,N_10301);
or U10511 (N_10511,N_10223,N_10242);
nand U10512 (N_10512,N_10468,N_10459);
xor U10513 (N_10513,N_10353,N_10333);
and U10514 (N_10514,N_10229,N_10483);
nor U10515 (N_10515,N_10373,N_10406);
nor U10516 (N_10516,N_10486,N_10447);
nor U10517 (N_10517,N_10294,N_10492);
nand U10518 (N_10518,N_10420,N_10324);
xnor U10519 (N_10519,N_10422,N_10414);
or U10520 (N_10520,N_10397,N_10304);
nor U10521 (N_10521,N_10404,N_10408);
nand U10522 (N_10522,N_10307,N_10350);
xnor U10523 (N_10523,N_10376,N_10298);
nand U10524 (N_10524,N_10417,N_10285);
nand U10525 (N_10525,N_10395,N_10443);
xor U10526 (N_10526,N_10308,N_10368);
and U10527 (N_10527,N_10211,N_10437);
and U10528 (N_10528,N_10379,N_10204);
nand U10529 (N_10529,N_10394,N_10329);
nand U10530 (N_10530,N_10331,N_10388);
and U10531 (N_10531,N_10244,N_10476);
and U10532 (N_10532,N_10365,N_10338);
xor U10533 (N_10533,N_10231,N_10465);
nor U10534 (N_10534,N_10366,N_10415);
nand U10535 (N_10535,N_10206,N_10336);
and U10536 (N_10536,N_10385,N_10384);
and U10537 (N_10537,N_10435,N_10264);
and U10538 (N_10538,N_10403,N_10339);
and U10539 (N_10539,N_10359,N_10421);
or U10540 (N_10540,N_10386,N_10208);
nor U10541 (N_10541,N_10202,N_10234);
and U10542 (N_10542,N_10252,N_10372);
and U10543 (N_10543,N_10265,N_10480);
or U10544 (N_10544,N_10269,N_10203);
nor U10545 (N_10545,N_10491,N_10249);
xnor U10546 (N_10546,N_10296,N_10402);
or U10547 (N_10547,N_10389,N_10342);
nor U10548 (N_10548,N_10464,N_10398);
nor U10549 (N_10549,N_10456,N_10283);
and U10550 (N_10550,N_10474,N_10449);
nor U10551 (N_10551,N_10340,N_10248);
nand U10552 (N_10552,N_10488,N_10303);
or U10553 (N_10553,N_10473,N_10452);
nand U10554 (N_10554,N_10251,N_10300);
or U10555 (N_10555,N_10232,N_10462);
or U10556 (N_10556,N_10345,N_10419);
or U10557 (N_10557,N_10467,N_10327);
nor U10558 (N_10558,N_10418,N_10457);
xor U10559 (N_10559,N_10455,N_10305);
nor U10560 (N_10560,N_10320,N_10302);
and U10561 (N_10561,N_10216,N_10262);
xor U10562 (N_10562,N_10217,N_10278);
nor U10563 (N_10563,N_10469,N_10470);
xnor U10564 (N_10564,N_10201,N_10215);
nand U10565 (N_10565,N_10487,N_10281);
nand U10566 (N_10566,N_10337,N_10409);
or U10567 (N_10567,N_10429,N_10237);
nor U10568 (N_10568,N_10259,N_10263);
nor U10569 (N_10569,N_10375,N_10255);
and U10570 (N_10570,N_10258,N_10433);
nor U10571 (N_10571,N_10377,N_10214);
xnor U10572 (N_10572,N_10362,N_10434);
xnor U10573 (N_10573,N_10222,N_10383);
nor U10574 (N_10574,N_10430,N_10330);
or U10575 (N_10575,N_10411,N_10479);
or U10576 (N_10576,N_10254,N_10367);
or U10577 (N_10577,N_10380,N_10267);
nor U10578 (N_10578,N_10322,N_10235);
nand U10579 (N_10579,N_10387,N_10364);
nand U10580 (N_10580,N_10312,N_10451);
or U10581 (N_10581,N_10458,N_10289);
and U10582 (N_10582,N_10390,N_10432);
nor U10583 (N_10583,N_10275,N_10354);
and U10584 (N_10584,N_10493,N_10343);
nor U10585 (N_10585,N_10311,N_10356);
xor U10586 (N_10586,N_10328,N_10205);
or U10587 (N_10587,N_10219,N_10497);
xor U10588 (N_10588,N_10370,N_10349);
nand U10589 (N_10589,N_10371,N_10247);
nor U10590 (N_10590,N_10230,N_10374);
or U10591 (N_10591,N_10318,N_10268);
and U10592 (N_10592,N_10442,N_10266);
or U10593 (N_10593,N_10423,N_10369);
and U10594 (N_10594,N_10334,N_10292);
and U10595 (N_10595,N_10256,N_10489);
or U10596 (N_10596,N_10413,N_10287);
or U10597 (N_10597,N_10286,N_10315);
nand U10598 (N_10598,N_10436,N_10471);
nor U10599 (N_10599,N_10317,N_10213);
xor U10600 (N_10600,N_10405,N_10253);
nor U10601 (N_10601,N_10257,N_10475);
nand U10602 (N_10602,N_10313,N_10407);
and U10603 (N_10603,N_10477,N_10396);
nand U10604 (N_10604,N_10293,N_10400);
nand U10605 (N_10605,N_10261,N_10291);
nand U10606 (N_10606,N_10271,N_10412);
or U10607 (N_10607,N_10310,N_10494);
nand U10608 (N_10608,N_10299,N_10341);
xnor U10609 (N_10609,N_10484,N_10431);
nand U10610 (N_10610,N_10236,N_10450);
xnor U10611 (N_10611,N_10314,N_10348);
and U10612 (N_10612,N_10274,N_10270);
xor U10613 (N_10613,N_10495,N_10226);
xnor U10614 (N_10614,N_10227,N_10361);
and U10615 (N_10615,N_10446,N_10358);
nor U10616 (N_10616,N_10220,N_10439);
nor U10617 (N_10617,N_10280,N_10453);
nand U10618 (N_10618,N_10355,N_10321);
or U10619 (N_10619,N_10207,N_10454);
or U10620 (N_10620,N_10461,N_10221);
nand U10621 (N_10621,N_10410,N_10200);
xor U10622 (N_10622,N_10319,N_10309);
nand U10623 (N_10623,N_10401,N_10246);
nor U10624 (N_10624,N_10239,N_10218);
nand U10625 (N_10625,N_10245,N_10279);
or U10626 (N_10626,N_10392,N_10347);
xnor U10627 (N_10627,N_10472,N_10427);
and U10628 (N_10628,N_10444,N_10295);
or U10629 (N_10629,N_10260,N_10233);
nand U10630 (N_10630,N_10277,N_10250);
xor U10631 (N_10631,N_10399,N_10332);
xnor U10632 (N_10632,N_10297,N_10424);
xor U10633 (N_10633,N_10441,N_10485);
and U10634 (N_10634,N_10498,N_10352);
nand U10635 (N_10635,N_10466,N_10360);
and U10636 (N_10636,N_10284,N_10426);
nand U10637 (N_10637,N_10290,N_10243);
or U10638 (N_10638,N_10428,N_10276);
nand U10639 (N_10639,N_10344,N_10448);
or U10640 (N_10640,N_10381,N_10440);
or U10641 (N_10641,N_10326,N_10393);
or U10642 (N_10642,N_10228,N_10460);
and U10643 (N_10643,N_10273,N_10425);
or U10644 (N_10644,N_10416,N_10438);
or U10645 (N_10645,N_10463,N_10210);
xor U10646 (N_10646,N_10481,N_10478);
xnor U10647 (N_10647,N_10382,N_10209);
or U10648 (N_10648,N_10496,N_10306);
and U10649 (N_10649,N_10335,N_10241);
or U10650 (N_10650,N_10333,N_10447);
or U10651 (N_10651,N_10490,N_10220);
and U10652 (N_10652,N_10367,N_10260);
or U10653 (N_10653,N_10415,N_10482);
and U10654 (N_10654,N_10253,N_10401);
or U10655 (N_10655,N_10390,N_10347);
and U10656 (N_10656,N_10247,N_10258);
xor U10657 (N_10657,N_10354,N_10335);
and U10658 (N_10658,N_10406,N_10296);
nand U10659 (N_10659,N_10299,N_10278);
or U10660 (N_10660,N_10348,N_10250);
or U10661 (N_10661,N_10280,N_10342);
or U10662 (N_10662,N_10428,N_10331);
nor U10663 (N_10663,N_10434,N_10415);
and U10664 (N_10664,N_10467,N_10252);
nor U10665 (N_10665,N_10238,N_10424);
xor U10666 (N_10666,N_10461,N_10243);
or U10667 (N_10667,N_10361,N_10241);
xor U10668 (N_10668,N_10399,N_10372);
xor U10669 (N_10669,N_10272,N_10271);
nand U10670 (N_10670,N_10455,N_10405);
or U10671 (N_10671,N_10249,N_10406);
nand U10672 (N_10672,N_10385,N_10337);
nor U10673 (N_10673,N_10284,N_10471);
nand U10674 (N_10674,N_10412,N_10461);
and U10675 (N_10675,N_10480,N_10378);
or U10676 (N_10676,N_10240,N_10219);
or U10677 (N_10677,N_10370,N_10223);
xor U10678 (N_10678,N_10470,N_10319);
and U10679 (N_10679,N_10210,N_10279);
or U10680 (N_10680,N_10231,N_10257);
or U10681 (N_10681,N_10383,N_10387);
nor U10682 (N_10682,N_10373,N_10242);
or U10683 (N_10683,N_10468,N_10425);
or U10684 (N_10684,N_10265,N_10282);
xnor U10685 (N_10685,N_10352,N_10286);
and U10686 (N_10686,N_10496,N_10240);
and U10687 (N_10687,N_10328,N_10453);
nor U10688 (N_10688,N_10225,N_10421);
and U10689 (N_10689,N_10262,N_10343);
or U10690 (N_10690,N_10380,N_10363);
xnor U10691 (N_10691,N_10224,N_10302);
and U10692 (N_10692,N_10285,N_10378);
nand U10693 (N_10693,N_10256,N_10380);
xor U10694 (N_10694,N_10410,N_10499);
and U10695 (N_10695,N_10268,N_10405);
xnor U10696 (N_10696,N_10247,N_10260);
nor U10697 (N_10697,N_10346,N_10464);
or U10698 (N_10698,N_10323,N_10224);
and U10699 (N_10699,N_10448,N_10224);
or U10700 (N_10700,N_10339,N_10415);
xnor U10701 (N_10701,N_10359,N_10440);
nor U10702 (N_10702,N_10292,N_10251);
nand U10703 (N_10703,N_10411,N_10351);
xnor U10704 (N_10704,N_10236,N_10345);
and U10705 (N_10705,N_10230,N_10426);
xnor U10706 (N_10706,N_10392,N_10357);
xor U10707 (N_10707,N_10361,N_10364);
or U10708 (N_10708,N_10370,N_10200);
and U10709 (N_10709,N_10372,N_10423);
nand U10710 (N_10710,N_10457,N_10209);
xor U10711 (N_10711,N_10343,N_10490);
xnor U10712 (N_10712,N_10214,N_10497);
nor U10713 (N_10713,N_10393,N_10274);
xnor U10714 (N_10714,N_10219,N_10245);
and U10715 (N_10715,N_10472,N_10380);
or U10716 (N_10716,N_10353,N_10281);
xnor U10717 (N_10717,N_10419,N_10448);
and U10718 (N_10718,N_10346,N_10281);
or U10719 (N_10719,N_10363,N_10416);
or U10720 (N_10720,N_10438,N_10263);
and U10721 (N_10721,N_10451,N_10322);
nand U10722 (N_10722,N_10265,N_10378);
and U10723 (N_10723,N_10473,N_10387);
and U10724 (N_10724,N_10252,N_10336);
and U10725 (N_10725,N_10245,N_10363);
nor U10726 (N_10726,N_10326,N_10359);
nor U10727 (N_10727,N_10367,N_10425);
xor U10728 (N_10728,N_10330,N_10306);
and U10729 (N_10729,N_10341,N_10268);
xnor U10730 (N_10730,N_10338,N_10442);
and U10731 (N_10731,N_10297,N_10213);
xnor U10732 (N_10732,N_10252,N_10202);
nor U10733 (N_10733,N_10378,N_10366);
and U10734 (N_10734,N_10429,N_10291);
xor U10735 (N_10735,N_10229,N_10253);
and U10736 (N_10736,N_10373,N_10232);
nor U10737 (N_10737,N_10304,N_10485);
xor U10738 (N_10738,N_10287,N_10428);
and U10739 (N_10739,N_10439,N_10463);
nor U10740 (N_10740,N_10329,N_10200);
or U10741 (N_10741,N_10450,N_10410);
nor U10742 (N_10742,N_10229,N_10336);
and U10743 (N_10743,N_10352,N_10457);
and U10744 (N_10744,N_10279,N_10207);
xor U10745 (N_10745,N_10365,N_10385);
or U10746 (N_10746,N_10247,N_10318);
xor U10747 (N_10747,N_10402,N_10336);
or U10748 (N_10748,N_10257,N_10469);
nor U10749 (N_10749,N_10346,N_10396);
xnor U10750 (N_10750,N_10231,N_10202);
nor U10751 (N_10751,N_10340,N_10289);
nand U10752 (N_10752,N_10364,N_10446);
nor U10753 (N_10753,N_10224,N_10309);
nor U10754 (N_10754,N_10402,N_10210);
xor U10755 (N_10755,N_10212,N_10300);
xnor U10756 (N_10756,N_10351,N_10240);
xnor U10757 (N_10757,N_10439,N_10449);
and U10758 (N_10758,N_10333,N_10303);
nand U10759 (N_10759,N_10335,N_10250);
or U10760 (N_10760,N_10367,N_10258);
nand U10761 (N_10761,N_10303,N_10471);
nand U10762 (N_10762,N_10271,N_10496);
nand U10763 (N_10763,N_10286,N_10430);
and U10764 (N_10764,N_10382,N_10365);
xor U10765 (N_10765,N_10210,N_10481);
nor U10766 (N_10766,N_10364,N_10244);
nor U10767 (N_10767,N_10200,N_10355);
or U10768 (N_10768,N_10239,N_10202);
and U10769 (N_10769,N_10355,N_10287);
and U10770 (N_10770,N_10312,N_10244);
or U10771 (N_10771,N_10386,N_10364);
xnor U10772 (N_10772,N_10311,N_10421);
nor U10773 (N_10773,N_10203,N_10248);
nor U10774 (N_10774,N_10422,N_10358);
nand U10775 (N_10775,N_10263,N_10233);
xnor U10776 (N_10776,N_10210,N_10261);
or U10777 (N_10777,N_10250,N_10360);
nand U10778 (N_10778,N_10305,N_10343);
and U10779 (N_10779,N_10323,N_10266);
and U10780 (N_10780,N_10217,N_10465);
nand U10781 (N_10781,N_10214,N_10281);
xor U10782 (N_10782,N_10241,N_10292);
and U10783 (N_10783,N_10314,N_10264);
and U10784 (N_10784,N_10265,N_10477);
nand U10785 (N_10785,N_10377,N_10421);
and U10786 (N_10786,N_10422,N_10389);
nand U10787 (N_10787,N_10291,N_10371);
and U10788 (N_10788,N_10211,N_10233);
and U10789 (N_10789,N_10333,N_10361);
nand U10790 (N_10790,N_10235,N_10413);
or U10791 (N_10791,N_10372,N_10453);
nand U10792 (N_10792,N_10267,N_10288);
and U10793 (N_10793,N_10499,N_10486);
nand U10794 (N_10794,N_10283,N_10451);
or U10795 (N_10795,N_10445,N_10341);
or U10796 (N_10796,N_10400,N_10203);
or U10797 (N_10797,N_10410,N_10454);
nand U10798 (N_10798,N_10260,N_10280);
or U10799 (N_10799,N_10299,N_10435);
and U10800 (N_10800,N_10558,N_10652);
or U10801 (N_10801,N_10671,N_10581);
or U10802 (N_10802,N_10718,N_10756);
and U10803 (N_10803,N_10527,N_10621);
xnor U10804 (N_10804,N_10759,N_10644);
nor U10805 (N_10805,N_10665,N_10568);
nor U10806 (N_10806,N_10552,N_10594);
nor U10807 (N_10807,N_10775,N_10702);
nand U10808 (N_10808,N_10647,N_10721);
and U10809 (N_10809,N_10653,N_10667);
xor U10810 (N_10810,N_10708,N_10618);
and U10811 (N_10811,N_10760,N_10731);
nor U10812 (N_10812,N_10692,N_10535);
nor U10813 (N_10813,N_10545,N_10749);
and U10814 (N_10814,N_10709,N_10559);
xnor U10815 (N_10815,N_10534,N_10758);
xnor U10816 (N_10816,N_10579,N_10543);
nand U10817 (N_10817,N_10640,N_10599);
or U10818 (N_10818,N_10502,N_10727);
nor U10819 (N_10819,N_10521,N_10525);
or U10820 (N_10820,N_10530,N_10738);
or U10821 (N_10821,N_10726,N_10714);
xor U10822 (N_10822,N_10791,N_10508);
or U10823 (N_10823,N_10607,N_10588);
nand U10824 (N_10824,N_10522,N_10503);
or U10825 (N_10825,N_10734,N_10752);
nand U10826 (N_10826,N_10757,N_10693);
nand U10827 (N_10827,N_10748,N_10732);
and U10828 (N_10828,N_10565,N_10542);
and U10829 (N_10829,N_10638,N_10600);
xnor U10830 (N_10830,N_10747,N_10639);
and U10831 (N_10831,N_10571,N_10694);
nand U10832 (N_10832,N_10628,N_10511);
or U10833 (N_10833,N_10541,N_10561);
and U10834 (N_10834,N_10645,N_10664);
or U10835 (N_10835,N_10532,N_10793);
xnor U10836 (N_10836,N_10792,N_10669);
nand U10837 (N_10837,N_10509,N_10625);
nand U10838 (N_10838,N_10507,N_10728);
or U10839 (N_10839,N_10700,N_10668);
nand U10840 (N_10840,N_10583,N_10706);
or U10841 (N_10841,N_10554,N_10710);
or U10842 (N_10842,N_10787,N_10678);
nand U10843 (N_10843,N_10570,N_10557);
or U10844 (N_10844,N_10587,N_10670);
xnor U10845 (N_10845,N_10797,N_10707);
nand U10846 (N_10846,N_10604,N_10737);
nand U10847 (N_10847,N_10646,N_10553);
xnor U10848 (N_10848,N_10696,N_10540);
nand U10849 (N_10849,N_10631,N_10586);
and U10850 (N_10850,N_10705,N_10697);
nor U10851 (N_10851,N_10769,N_10677);
nand U10852 (N_10852,N_10575,N_10770);
nand U10853 (N_10853,N_10567,N_10780);
nor U10854 (N_10854,N_10582,N_10562);
nor U10855 (N_10855,N_10741,N_10506);
nor U10856 (N_10856,N_10563,N_10674);
xor U10857 (N_10857,N_10516,N_10673);
xnor U10858 (N_10858,N_10578,N_10635);
or U10859 (N_10859,N_10572,N_10795);
nor U10860 (N_10860,N_10514,N_10690);
xor U10861 (N_10861,N_10596,N_10622);
xnor U10862 (N_10862,N_10623,N_10611);
and U10863 (N_10863,N_10650,N_10739);
nor U10864 (N_10864,N_10755,N_10574);
and U10865 (N_10865,N_10781,N_10753);
nor U10866 (N_10866,N_10501,N_10699);
nand U10867 (N_10867,N_10589,N_10722);
and U10868 (N_10868,N_10679,N_10617);
nand U10869 (N_10869,N_10736,N_10536);
or U10870 (N_10870,N_10765,N_10729);
or U10871 (N_10871,N_10666,N_10768);
and U10872 (N_10872,N_10661,N_10680);
and U10873 (N_10873,N_10681,N_10515);
nand U10874 (N_10874,N_10790,N_10691);
or U10875 (N_10875,N_10688,N_10569);
nor U10876 (N_10876,N_10637,N_10751);
nand U10877 (N_10877,N_10658,N_10539);
and U10878 (N_10878,N_10512,N_10523);
and U10879 (N_10879,N_10740,N_10610);
xnor U10880 (N_10880,N_10641,N_10774);
and U10881 (N_10881,N_10533,N_10730);
xnor U10882 (N_10882,N_10733,N_10655);
xnor U10883 (N_10883,N_10613,N_10779);
or U10884 (N_10884,N_10636,N_10783);
and U10885 (N_10885,N_10609,N_10689);
xor U10886 (N_10886,N_10684,N_10616);
and U10887 (N_10887,N_10773,N_10672);
and U10888 (N_10888,N_10750,N_10551);
nand U10889 (N_10889,N_10510,N_10789);
nand U10890 (N_10890,N_10742,N_10663);
or U10891 (N_10891,N_10606,N_10698);
and U10892 (N_10892,N_10767,N_10717);
xor U10893 (N_10893,N_10573,N_10794);
nand U10894 (N_10894,N_10782,N_10585);
nand U10895 (N_10895,N_10785,N_10746);
nor U10896 (N_10896,N_10643,N_10743);
nand U10897 (N_10897,N_10719,N_10626);
nand U10898 (N_10898,N_10505,N_10654);
or U10899 (N_10899,N_10786,N_10788);
nor U10900 (N_10900,N_10686,N_10685);
and U10901 (N_10901,N_10528,N_10524);
nor U10902 (N_10902,N_10598,N_10675);
nor U10903 (N_10903,N_10584,N_10619);
nor U10904 (N_10904,N_10517,N_10630);
xor U10905 (N_10905,N_10519,N_10546);
nand U10906 (N_10906,N_10591,N_10762);
and U10907 (N_10907,N_10615,N_10576);
or U10908 (N_10908,N_10590,N_10687);
nor U10909 (N_10909,N_10798,N_10634);
nor U10910 (N_10910,N_10597,N_10724);
nand U10911 (N_10911,N_10547,N_10766);
nor U10912 (N_10912,N_10796,N_10712);
or U10913 (N_10913,N_10725,N_10526);
nor U10914 (N_10914,N_10662,N_10772);
nor U10915 (N_10915,N_10744,N_10715);
xnor U10916 (N_10916,N_10548,N_10603);
nor U10917 (N_10917,N_10704,N_10538);
nand U10918 (N_10918,N_10593,N_10651);
nor U10919 (N_10919,N_10633,N_10555);
and U10920 (N_10920,N_10577,N_10520);
or U10921 (N_10921,N_10556,N_10754);
nand U10922 (N_10922,N_10657,N_10632);
and U10923 (N_10923,N_10602,N_10682);
or U10924 (N_10924,N_10761,N_10550);
or U10925 (N_10925,N_10544,N_10778);
xor U10926 (N_10926,N_10564,N_10642);
nor U10927 (N_10927,N_10595,N_10713);
and U10928 (N_10928,N_10656,N_10580);
nand U10929 (N_10929,N_10701,N_10500);
xor U10930 (N_10930,N_10745,N_10799);
nor U10931 (N_10931,N_10649,N_10735);
and U10932 (N_10932,N_10560,N_10659);
xor U10933 (N_10933,N_10608,N_10605);
nor U10934 (N_10934,N_10676,N_10683);
or U10935 (N_10935,N_10648,N_10614);
nand U10936 (N_10936,N_10612,N_10723);
and U10937 (N_10937,N_10620,N_10720);
and U10938 (N_10938,N_10711,N_10771);
or U10939 (N_10939,N_10566,N_10537);
xor U10940 (N_10940,N_10592,N_10764);
nand U10941 (N_10941,N_10529,N_10777);
nand U10942 (N_10942,N_10627,N_10601);
and U10943 (N_10943,N_10549,N_10518);
or U10944 (N_10944,N_10695,N_10629);
xor U10945 (N_10945,N_10763,N_10531);
nand U10946 (N_10946,N_10716,N_10703);
and U10947 (N_10947,N_10784,N_10776);
and U10948 (N_10948,N_10513,N_10624);
nand U10949 (N_10949,N_10504,N_10660);
nor U10950 (N_10950,N_10616,N_10675);
xor U10951 (N_10951,N_10538,N_10725);
or U10952 (N_10952,N_10668,N_10625);
nor U10953 (N_10953,N_10517,N_10515);
nor U10954 (N_10954,N_10607,N_10782);
nor U10955 (N_10955,N_10596,N_10594);
and U10956 (N_10956,N_10608,N_10601);
nand U10957 (N_10957,N_10630,N_10560);
nand U10958 (N_10958,N_10503,N_10684);
nor U10959 (N_10959,N_10748,N_10523);
nand U10960 (N_10960,N_10585,N_10677);
nor U10961 (N_10961,N_10570,N_10708);
and U10962 (N_10962,N_10561,N_10511);
xor U10963 (N_10963,N_10775,N_10517);
nand U10964 (N_10964,N_10719,N_10551);
and U10965 (N_10965,N_10699,N_10764);
nand U10966 (N_10966,N_10530,N_10677);
nor U10967 (N_10967,N_10615,N_10651);
xor U10968 (N_10968,N_10598,N_10630);
and U10969 (N_10969,N_10784,N_10651);
or U10970 (N_10970,N_10736,N_10789);
nand U10971 (N_10971,N_10739,N_10678);
and U10972 (N_10972,N_10772,N_10766);
and U10973 (N_10973,N_10568,N_10696);
or U10974 (N_10974,N_10652,N_10596);
xor U10975 (N_10975,N_10509,N_10540);
and U10976 (N_10976,N_10654,N_10728);
nor U10977 (N_10977,N_10612,N_10619);
xor U10978 (N_10978,N_10564,N_10690);
nor U10979 (N_10979,N_10695,N_10771);
nand U10980 (N_10980,N_10738,N_10574);
nand U10981 (N_10981,N_10780,N_10562);
xnor U10982 (N_10982,N_10559,N_10761);
nor U10983 (N_10983,N_10793,N_10608);
and U10984 (N_10984,N_10648,N_10739);
xor U10985 (N_10985,N_10619,N_10537);
nand U10986 (N_10986,N_10525,N_10623);
nor U10987 (N_10987,N_10623,N_10584);
xnor U10988 (N_10988,N_10643,N_10688);
nor U10989 (N_10989,N_10605,N_10654);
nand U10990 (N_10990,N_10691,N_10525);
nor U10991 (N_10991,N_10588,N_10563);
nor U10992 (N_10992,N_10555,N_10615);
nor U10993 (N_10993,N_10684,N_10529);
xnor U10994 (N_10994,N_10506,N_10561);
nor U10995 (N_10995,N_10505,N_10714);
or U10996 (N_10996,N_10609,N_10621);
nor U10997 (N_10997,N_10522,N_10581);
xnor U10998 (N_10998,N_10500,N_10525);
xnor U10999 (N_10999,N_10561,N_10500);
and U11000 (N_11000,N_10656,N_10551);
xor U11001 (N_11001,N_10567,N_10666);
nand U11002 (N_11002,N_10652,N_10772);
xor U11003 (N_11003,N_10586,N_10595);
and U11004 (N_11004,N_10501,N_10750);
nor U11005 (N_11005,N_10713,N_10736);
and U11006 (N_11006,N_10633,N_10758);
nand U11007 (N_11007,N_10555,N_10715);
or U11008 (N_11008,N_10749,N_10584);
nor U11009 (N_11009,N_10552,N_10757);
and U11010 (N_11010,N_10707,N_10575);
xnor U11011 (N_11011,N_10584,N_10598);
nor U11012 (N_11012,N_10610,N_10694);
and U11013 (N_11013,N_10583,N_10508);
or U11014 (N_11014,N_10511,N_10571);
xor U11015 (N_11015,N_10624,N_10642);
or U11016 (N_11016,N_10617,N_10514);
and U11017 (N_11017,N_10527,N_10791);
nor U11018 (N_11018,N_10743,N_10719);
or U11019 (N_11019,N_10511,N_10752);
nor U11020 (N_11020,N_10673,N_10707);
or U11021 (N_11021,N_10762,N_10703);
nand U11022 (N_11022,N_10591,N_10781);
and U11023 (N_11023,N_10745,N_10776);
nor U11024 (N_11024,N_10521,N_10708);
nand U11025 (N_11025,N_10638,N_10688);
or U11026 (N_11026,N_10587,N_10689);
xnor U11027 (N_11027,N_10748,N_10782);
or U11028 (N_11028,N_10745,N_10655);
xor U11029 (N_11029,N_10782,N_10662);
or U11030 (N_11030,N_10714,N_10560);
or U11031 (N_11031,N_10790,N_10554);
xnor U11032 (N_11032,N_10616,N_10548);
nor U11033 (N_11033,N_10599,N_10613);
and U11034 (N_11034,N_10583,N_10546);
nand U11035 (N_11035,N_10588,N_10686);
or U11036 (N_11036,N_10687,N_10508);
xnor U11037 (N_11037,N_10567,N_10717);
nor U11038 (N_11038,N_10507,N_10583);
and U11039 (N_11039,N_10660,N_10621);
nor U11040 (N_11040,N_10511,N_10576);
nand U11041 (N_11041,N_10541,N_10656);
xnor U11042 (N_11042,N_10786,N_10618);
nand U11043 (N_11043,N_10557,N_10757);
nand U11044 (N_11044,N_10744,N_10629);
or U11045 (N_11045,N_10619,N_10796);
or U11046 (N_11046,N_10676,N_10784);
nor U11047 (N_11047,N_10693,N_10504);
xor U11048 (N_11048,N_10525,N_10722);
xnor U11049 (N_11049,N_10567,N_10742);
xor U11050 (N_11050,N_10791,N_10665);
nor U11051 (N_11051,N_10638,N_10625);
xor U11052 (N_11052,N_10775,N_10602);
xor U11053 (N_11053,N_10688,N_10737);
or U11054 (N_11054,N_10630,N_10561);
and U11055 (N_11055,N_10779,N_10632);
or U11056 (N_11056,N_10724,N_10568);
xor U11057 (N_11057,N_10753,N_10681);
nand U11058 (N_11058,N_10646,N_10767);
nand U11059 (N_11059,N_10683,N_10629);
and U11060 (N_11060,N_10581,N_10609);
xor U11061 (N_11061,N_10683,N_10705);
nand U11062 (N_11062,N_10750,N_10528);
nor U11063 (N_11063,N_10577,N_10774);
xnor U11064 (N_11064,N_10523,N_10730);
xor U11065 (N_11065,N_10681,N_10684);
nor U11066 (N_11066,N_10799,N_10788);
nor U11067 (N_11067,N_10778,N_10677);
xor U11068 (N_11068,N_10796,N_10719);
xnor U11069 (N_11069,N_10635,N_10727);
and U11070 (N_11070,N_10728,N_10790);
nor U11071 (N_11071,N_10761,N_10688);
or U11072 (N_11072,N_10500,N_10579);
nor U11073 (N_11073,N_10672,N_10737);
and U11074 (N_11074,N_10691,N_10528);
or U11075 (N_11075,N_10755,N_10611);
xnor U11076 (N_11076,N_10651,N_10513);
nor U11077 (N_11077,N_10792,N_10729);
nor U11078 (N_11078,N_10526,N_10612);
nor U11079 (N_11079,N_10681,N_10797);
xor U11080 (N_11080,N_10671,N_10603);
nand U11081 (N_11081,N_10646,N_10584);
or U11082 (N_11082,N_10673,N_10570);
nand U11083 (N_11083,N_10609,N_10745);
xor U11084 (N_11084,N_10521,N_10670);
and U11085 (N_11085,N_10540,N_10781);
xnor U11086 (N_11086,N_10581,N_10533);
nor U11087 (N_11087,N_10525,N_10656);
xor U11088 (N_11088,N_10534,N_10723);
and U11089 (N_11089,N_10749,N_10554);
xor U11090 (N_11090,N_10704,N_10756);
or U11091 (N_11091,N_10548,N_10589);
or U11092 (N_11092,N_10776,N_10721);
nand U11093 (N_11093,N_10560,N_10763);
or U11094 (N_11094,N_10730,N_10548);
nand U11095 (N_11095,N_10745,N_10523);
xnor U11096 (N_11096,N_10729,N_10544);
nand U11097 (N_11097,N_10529,N_10658);
nor U11098 (N_11098,N_10703,N_10708);
or U11099 (N_11099,N_10781,N_10691);
xnor U11100 (N_11100,N_10882,N_11014);
and U11101 (N_11101,N_11091,N_10925);
and U11102 (N_11102,N_10855,N_10864);
nand U11103 (N_11103,N_10867,N_10815);
nand U11104 (N_11104,N_10871,N_11005);
nor U11105 (N_11105,N_10939,N_11042);
and U11106 (N_11106,N_10987,N_11067);
and U11107 (N_11107,N_10954,N_11012);
xor U11108 (N_11108,N_10991,N_11078);
nor U11109 (N_11109,N_10953,N_10847);
xnor U11110 (N_11110,N_10914,N_10965);
nand U11111 (N_11111,N_10898,N_11089);
nor U11112 (N_11112,N_11028,N_10988);
xor U11113 (N_11113,N_10934,N_10892);
nand U11114 (N_11114,N_11055,N_11024);
xnor U11115 (N_11115,N_10935,N_11038);
nor U11116 (N_11116,N_10904,N_10959);
xor U11117 (N_11117,N_10802,N_11016);
nor U11118 (N_11118,N_10908,N_11083);
xnor U11119 (N_11119,N_10944,N_10857);
xnor U11120 (N_11120,N_11035,N_10861);
and U11121 (N_11121,N_10902,N_10933);
nand U11122 (N_11122,N_10969,N_11013);
nor U11123 (N_11123,N_10929,N_10818);
nor U11124 (N_11124,N_10996,N_10907);
xor U11125 (N_11125,N_10984,N_11070);
and U11126 (N_11126,N_10844,N_10838);
nor U11127 (N_11127,N_10806,N_10900);
and U11128 (N_11128,N_10896,N_10903);
nand U11129 (N_11129,N_11074,N_11066);
or U11130 (N_11130,N_10848,N_10852);
or U11131 (N_11131,N_10877,N_10997);
and U11132 (N_11132,N_10856,N_11011);
nand U11133 (N_11133,N_11047,N_10941);
nand U11134 (N_11134,N_11052,N_10891);
nand U11135 (N_11135,N_11079,N_10917);
xor U11136 (N_11136,N_11040,N_11021);
nand U11137 (N_11137,N_10943,N_11077);
nor U11138 (N_11138,N_10961,N_10950);
nand U11139 (N_11139,N_10971,N_11023);
and U11140 (N_11140,N_11098,N_10957);
and U11141 (N_11141,N_11076,N_10865);
nor U11142 (N_11142,N_10849,N_10975);
xor U11143 (N_11143,N_10827,N_10909);
nor U11144 (N_11144,N_10817,N_11072);
or U11145 (N_11145,N_10809,N_10912);
nor U11146 (N_11146,N_11015,N_10811);
nand U11147 (N_11147,N_11039,N_10833);
and U11148 (N_11148,N_10862,N_11082);
and U11149 (N_11149,N_11032,N_11007);
or U11150 (N_11150,N_11092,N_11059);
and U11151 (N_11151,N_10949,N_10938);
and U11152 (N_11152,N_10993,N_10834);
nand U11153 (N_11153,N_10889,N_10966);
nand U11154 (N_11154,N_10859,N_11003);
nand U11155 (N_11155,N_10986,N_11001);
nor U11156 (N_11156,N_11054,N_10905);
nor U11157 (N_11157,N_10926,N_10853);
xnor U11158 (N_11158,N_10860,N_10958);
xor U11159 (N_11159,N_10928,N_10921);
or U11160 (N_11160,N_10951,N_10843);
xor U11161 (N_11161,N_10835,N_11053);
nor U11162 (N_11162,N_11010,N_10879);
and U11163 (N_11163,N_10816,N_10890);
xnor U11164 (N_11164,N_11090,N_11056);
and U11165 (N_11165,N_10812,N_10845);
nor U11166 (N_11166,N_10911,N_11033);
xor U11167 (N_11167,N_10805,N_10895);
xnor U11168 (N_11168,N_11050,N_10869);
xnor U11169 (N_11169,N_11064,N_10999);
nand U11170 (N_11170,N_10878,N_11019);
nand U11171 (N_11171,N_10854,N_11022);
and U11172 (N_11172,N_10936,N_10937);
nor U11173 (N_11173,N_10880,N_10897);
and U11174 (N_11174,N_10918,N_11017);
and U11175 (N_11175,N_10899,N_11073);
or U11176 (N_11176,N_10825,N_10875);
nor U11177 (N_11177,N_10823,N_10820);
or U11178 (N_11178,N_10989,N_10821);
nand U11179 (N_11179,N_10876,N_10832);
xnor U11180 (N_11180,N_10866,N_10828);
nand U11181 (N_11181,N_11044,N_10894);
or U11182 (N_11182,N_11000,N_11086);
nand U11183 (N_11183,N_10826,N_11049);
nor U11184 (N_11184,N_10945,N_10927);
and U11185 (N_11185,N_10808,N_11030);
xor U11186 (N_11186,N_11087,N_11099);
or U11187 (N_11187,N_10955,N_10964);
and U11188 (N_11188,N_10956,N_10901);
nand U11189 (N_11189,N_10923,N_10801);
and U11190 (N_11190,N_10840,N_11029);
nand U11191 (N_11191,N_10906,N_10974);
nor U11192 (N_11192,N_10973,N_10983);
nand U11193 (N_11193,N_11020,N_10804);
nand U11194 (N_11194,N_10831,N_10888);
or U11195 (N_11195,N_11068,N_10998);
nor U11196 (N_11196,N_11061,N_10851);
and U11197 (N_11197,N_11063,N_10994);
or U11198 (N_11198,N_11025,N_11080);
xor U11199 (N_11199,N_10976,N_11081);
nand U11200 (N_11200,N_11051,N_11060);
or U11201 (N_11201,N_11048,N_10979);
or U11202 (N_11202,N_10887,N_10824);
xor U11203 (N_11203,N_10800,N_10872);
and U11204 (N_11204,N_11034,N_11026);
nor U11205 (N_11205,N_10873,N_10916);
xnor U11206 (N_11206,N_11088,N_11093);
nand U11207 (N_11207,N_10822,N_11046);
nor U11208 (N_11208,N_10995,N_10980);
or U11209 (N_11209,N_11036,N_10846);
nand U11210 (N_11210,N_10807,N_11009);
and U11211 (N_11211,N_10977,N_11069);
xor U11212 (N_11212,N_11095,N_11037);
nor U11213 (N_11213,N_10910,N_10893);
nor U11214 (N_11214,N_10972,N_10982);
xor U11215 (N_11215,N_10813,N_10924);
xor U11216 (N_11216,N_10985,N_10870);
and U11217 (N_11217,N_10968,N_10837);
or U11218 (N_11218,N_10829,N_10814);
xor U11219 (N_11219,N_10884,N_10960);
xnor U11220 (N_11220,N_10819,N_10922);
and U11221 (N_11221,N_11004,N_10913);
xnor U11222 (N_11222,N_10842,N_11041);
nor U11223 (N_11223,N_11085,N_10962);
nand U11224 (N_11224,N_11065,N_11018);
or U11225 (N_11225,N_10830,N_10992);
xor U11226 (N_11226,N_10940,N_10883);
or U11227 (N_11227,N_11043,N_10886);
or U11228 (N_11228,N_11006,N_10981);
nor U11229 (N_11229,N_10850,N_10948);
nand U11230 (N_11230,N_10803,N_10963);
or U11231 (N_11231,N_10952,N_11094);
nor U11232 (N_11232,N_10920,N_10881);
or U11233 (N_11233,N_10931,N_11027);
nor U11234 (N_11234,N_11084,N_10946);
nor U11235 (N_11235,N_10947,N_10858);
or U11236 (N_11236,N_10942,N_11031);
and U11237 (N_11237,N_10932,N_10868);
and U11238 (N_11238,N_10839,N_10841);
nand U11239 (N_11239,N_11057,N_11096);
nand U11240 (N_11240,N_10970,N_10990);
nand U11241 (N_11241,N_10919,N_11008);
nor U11242 (N_11242,N_10885,N_11058);
nor U11243 (N_11243,N_11075,N_10967);
nor U11244 (N_11244,N_10930,N_11071);
xnor U11245 (N_11245,N_11045,N_10836);
and U11246 (N_11246,N_10978,N_10863);
xnor U11247 (N_11247,N_11097,N_11062);
or U11248 (N_11248,N_10874,N_11002);
nor U11249 (N_11249,N_10915,N_10810);
xnor U11250 (N_11250,N_10921,N_10885);
nor U11251 (N_11251,N_10944,N_10941);
nor U11252 (N_11252,N_11001,N_11094);
or U11253 (N_11253,N_11025,N_11010);
nor U11254 (N_11254,N_10912,N_11029);
and U11255 (N_11255,N_11007,N_11071);
and U11256 (N_11256,N_11025,N_11070);
or U11257 (N_11257,N_11001,N_10979);
and U11258 (N_11258,N_11037,N_10994);
nand U11259 (N_11259,N_11050,N_10872);
or U11260 (N_11260,N_11014,N_10982);
nand U11261 (N_11261,N_10893,N_11036);
xor U11262 (N_11262,N_11009,N_10870);
nor U11263 (N_11263,N_10844,N_11019);
nand U11264 (N_11264,N_10846,N_10989);
or U11265 (N_11265,N_10972,N_11054);
nand U11266 (N_11266,N_10905,N_10813);
and U11267 (N_11267,N_10932,N_10869);
xor U11268 (N_11268,N_10898,N_11099);
nand U11269 (N_11269,N_10875,N_10908);
or U11270 (N_11270,N_11006,N_10826);
nand U11271 (N_11271,N_11083,N_11026);
nor U11272 (N_11272,N_11091,N_11011);
or U11273 (N_11273,N_10871,N_11025);
and U11274 (N_11274,N_10967,N_11047);
nand U11275 (N_11275,N_11061,N_10947);
nand U11276 (N_11276,N_11020,N_11029);
nand U11277 (N_11277,N_11074,N_10857);
nand U11278 (N_11278,N_11068,N_10909);
xnor U11279 (N_11279,N_10828,N_10994);
nor U11280 (N_11280,N_11088,N_10868);
and U11281 (N_11281,N_10810,N_10842);
nor U11282 (N_11282,N_10933,N_10944);
nor U11283 (N_11283,N_11072,N_10814);
nand U11284 (N_11284,N_10800,N_11062);
xor U11285 (N_11285,N_11075,N_10959);
nand U11286 (N_11286,N_11081,N_11001);
xor U11287 (N_11287,N_10869,N_10830);
or U11288 (N_11288,N_10992,N_11032);
nor U11289 (N_11289,N_10883,N_11045);
nor U11290 (N_11290,N_11066,N_11095);
and U11291 (N_11291,N_10875,N_10921);
and U11292 (N_11292,N_11072,N_10980);
nor U11293 (N_11293,N_10973,N_10916);
and U11294 (N_11294,N_11012,N_10837);
or U11295 (N_11295,N_10980,N_11033);
and U11296 (N_11296,N_11075,N_10823);
nand U11297 (N_11297,N_11010,N_10859);
nor U11298 (N_11298,N_10807,N_10928);
nor U11299 (N_11299,N_10892,N_10844);
and U11300 (N_11300,N_11097,N_10825);
and U11301 (N_11301,N_11098,N_10878);
or U11302 (N_11302,N_10983,N_10816);
and U11303 (N_11303,N_10873,N_10941);
xnor U11304 (N_11304,N_10856,N_10847);
or U11305 (N_11305,N_10802,N_10806);
nor U11306 (N_11306,N_11084,N_10832);
xnor U11307 (N_11307,N_11001,N_10917);
xnor U11308 (N_11308,N_10846,N_10823);
or U11309 (N_11309,N_11053,N_10983);
xnor U11310 (N_11310,N_10848,N_10901);
xor U11311 (N_11311,N_10985,N_10840);
and U11312 (N_11312,N_10900,N_10930);
and U11313 (N_11313,N_10986,N_11013);
xnor U11314 (N_11314,N_11047,N_11004);
nand U11315 (N_11315,N_10828,N_10918);
and U11316 (N_11316,N_10992,N_10873);
nand U11317 (N_11317,N_10852,N_11065);
or U11318 (N_11318,N_10827,N_10829);
nor U11319 (N_11319,N_10857,N_10838);
xnor U11320 (N_11320,N_10849,N_10920);
nand U11321 (N_11321,N_11098,N_10818);
xnor U11322 (N_11322,N_10902,N_11095);
and U11323 (N_11323,N_10906,N_10981);
and U11324 (N_11324,N_10959,N_10989);
and U11325 (N_11325,N_11029,N_10881);
nand U11326 (N_11326,N_11019,N_10821);
nor U11327 (N_11327,N_10926,N_11089);
nor U11328 (N_11328,N_10903,N_10975);
nand U11329 (N_11329,N_11078,N_10920);
or U11330 (N_11330,N_10955,N_10849);
xnor U11331 (N_11331,N_10829,N_10944);
or U11332 (N_11332,N_10904,N_10980);
nand U11333 (N_11333,N_10951,N_11042);
nand U11334 (N_11334,N_11097,N_10936);
or U11335 (N_11335,N_10868,N_10838);
nor U11336 (N_11336,N_10816,N_11008);
and U11337 (N_11337,N_11096,N_10877);
or U11338 (N_11338,N_11077,N_11092);
nor U11339 (N_11339,N_11050,N_10812);
xor U11340 (N_11340,N_11025,N_11064);
or U11341 (N_11341,N_11022,N_11090);
nand U11342 (N_11342,N_10819,N_10923);
xnor U11343 (N_11343,N_10834,N_11009);
or U11344 (N_11344,N_11027,N_10850);
and U11345 (N_11345,N_10905,N_11026);
and U11346 (N_11346,N_10859,N_11066);
nand U11347 (N_11347,N_10886,N_10887);
and U11348 (N_11348,N_10950,N_10850);
xor U11349 (N_11349,N_11095,N_10845);
and U11350 (N_11350,N_10940,N_11078);
nor U11351 (N_11351,N_10979,N_10927);
xnor U11352 (N_11352,N_10980,N_11058);
or U11353 (N_11353,N_10965,N_11019);
nand U11354 (N_11354,N_10914,N_11074);
or U11355 (N_11355,N_11064,N_10873);
nand U11356 (N_11356,N_11074,N_11045);
or U11357 (N_11357,N_10820,N_10809);
nor U11358 (N_11358,N_10994,N_11070);
xnor U11359 (N_11359,N_11009,N_10959);
nor U11360 (N_11360,N_10833,N_10835);
nand U11361 (N_11361,N_11049,N_10918);
nand U11362 (N_11362,N_10815,N_10902);
and U11363 (N_11363,N_10819,N_10925);
or U11364 (N_11364,N_11011,N_10869);
and U11365 (N_11365,N_10815,N_10905);
or U11366 (N_11366,N_11097,N_10983);
xnor U11367 (N_11367,N_11070,N_10833);
nor U11368 (N_11368,N_11088,N_10944);
or U11369 (N_11369,N_11020,N_11076);
nor U11370 (N_11370,N_10880,N_11035);
nor U11371 (N_11371,N_10820,N_10869);
nand U11372 (N_11372,N_11072,N_10876);
nand U11373 (N_11373,N_10861,N_11043);
xor U11374 (N_11374,N_11001,N_11084);
and U11375 (N_11375,N_11099,N_10930);
nor U11376 (N_11376,N_10992,N_11054);
and U11377 (N_11377,N_11084,N_10889);
or U11378 (N_11378,N_10945,N_10850);
nor U11379 (N_11379,N_11096,N_11045);
nor U11380 (N_11380,N_11060,N_10823);
nand U11381 (N_11381,N_10891,N_11087);
nor U11382 (N_11382,N_11003,N_10906);
and U11383 (N_11383,N_11048,N_11003);
nand U11384 (N_11384,N_10804,N_10806);
nor U11385 (N_11385,N_10967,N_11028);
nor U11386 (N_11386,N_10803,N_11050);
nand U11387 (N_11387,N_10898,N_10816);
and U11388 (N_11388,N_10996,N_10965);
nor U11389 (N_11389,N_10950,N_11021);
nor U11390 (N_11390,N_10884,N_10828);
and U11391 (N_11391,N_10853,N_10847);
nor U11392 (N_11392,N_11075,N_10854);
and U11393 (N_11393,N_11061,N_11072);
nand U11394 (N_11394,N_11049,N_10933);
and U11395 (N_11395,N_11065,N_11063);
nor U11396 (N_11396,N_10927,N_11012);
or U11397 (N_11397,N_11011,N_10833);
and U11398 (N_11398,N_10821,N_11075);
and U11399 (N_11399,N_11089,N_10889);
and U11400 (N_11400,N_11109,N_11325);
nor U11401 (N_11401,N_11294,N_11137);
and U11402 (N_11402,N_11237,N_11371);
or U11403 (N_11403,N_11159,N_11378);
or U11404 (N_11404,N_11197,N_11281);
xnor U11405 (N_11405,N_11280,N_11307);
nand U11406 (N_11406,N_11279,N_11171);
nand U11407 (N_11407,N_11315,N_11338);
nand U11408 (N_11408,N_11234,N_11322);
xor U11409 (N_11409,N_11351,N_11270);
and U11410 (N_11410,N_11125,N_11146);
and U11411 (N_11411,N_11272,N_11214);
nand U11412 (N_11412,N_11106,N_11180);
nand U11413 (N_11413,N_11126,N_11347);
and U11414 (N_11414,N_11103,N_11285);
and U11415 (N_11415,N_11190,N_11114);
xor U11416 (N_11416,N_11264,N_11364);
nor U11417 (N_11417,N_11273,N_11184);
nand U11418 (N_11418,N_11334,N_11191);
nor U11419 (N_11419,N_11222,N_11302);
nor U11420 (N_11420,N_11374,N_11120);
or U11421 (N_11421,N_11110,N_11149);
nand U11422 (N_11422,N_11253,N_11203);
nor U11423 (N_11423,N_11221,N_11301);
or U11424 (N_11424,N_11292,N_11132);
and U11425 (N_11425,N_11376,N_11358);
xor U11426 (N_11426,N_11323,N_11179);
nand U11427 (N_11427,N_11233,N_11356);
xor U11428 (N_11428,N_11123,N_11399);
and U11429 (N_11429,N_11368,N_11207);
and U11430 (N_11430,N_11181,N_11161);
or U11431 (N_11431,N_11274,N_11202);
xor U11432 (N_11432,N_11306,N_11308);
xor U11433 (N_11433,N_11176,N_11187);
xnor U11434 (N_11434,N_11258,N_11138);
nor U11435 (N_11435,N_11134,N_11116);
nor U11436 (N_11436,N_11113,N_11393);
nand U11437 (N_11437,N_11101,N_11236);
or U11438 (N_11438,N_11199,N_11166);
nand U11439 (N_11439,N_11131,N_11341);
nand U11440 (N_11440,N_11316,N_11185);
and U11441 (N_11441,N_11350,N_11250);
nor U11442 (N_11442,N_11304,N_11319);
and U11443 (N_11443,N_11267,N_11271);
or U11444 (N_11444,N_11365,N_11303);
and U11445 (N_11445,N_11102,N_11108);
nand U11446 (N_11446,N_11130,N_11175);
xnor U11447 (N_11447,N_11295,N_11357);
nor U11448 (N_11448,N_11249,N_11195);
and U11449 (N_11449,N_11335,N_11167);
or U11450 (N_11450,N_11311,N_11331);
nor U11451 (N_11451,N_11259,N_11395);
nand U11452 (N_11452,N_11154,N_11160);
and U11453 (N_11453,N_11139,N_11381);
and U11454 (N_11454,N_11100,N_11328);
xnor U11455 (N_11455,N_11383,N_11387);
nor U11456 (N_11456,N_11300,N_11366);
and U11457 (N_11457,N_11115,N_11119);
and U11458 (N_11458,N_11291,N_11193);
and U11459 (N_11459,N_11299,N_11248);
and U11460 (N_11460,N_11204,N_11118);
nor U11461 (N_11461,N_11330,N_11255);
and U11462 (N_11462,N_11235,N_11163);
nor U11463 (N_11463,N_11104,N_11168);
or U11464 (N_11464,N_11290,N_11242);
xor U11465 (N_11465,N_11396,N_11162);
and U11466 (N_11466,N_11140,N_11337);
and U11467 (N_11467,N_11165,N_11286);
nor U11468 (N_11468,N_11243,N_11225);
nand U11469 (N_11469,N_11397,N_11170);
and U11470 (N_11470,N_11282,N_11135);
or U11471 (N_11471,N_11200,N_11345);
and U11472 (N_11472,N_11239,N_11196);
nor U11473 (N_11473,N_11318,N_11359);
and U11474 (N_11474,N_11133,N_11192);
or U11475 (N_11475,N_11212,N_11394);
and U11476 (N_11476,N_11367,N_11127);
nor U11477 (N_11477,N_11151,N_11217);
xnor U11478 (N_11478,N_11340,N_11178);
nor U11479 (N_11479,N_11326,N_11155);
nor U11480 (N_11480,N_11241,N_11260);
and U11481 (N_11481,N_11232,N_11287);
nor U11482 (N_11482,N_11173,N_11391);
xnor U11483 (N_11483,N_11372,N_11229);
and U11484 (N_11484,N_11208,N_11388);
or U11485 (N_11485,N_11215,N_11211);
xor U11486 (N_11486,N_11320,N_11240);
xor U11487 (N_11487,N_11321,N_11389);
or U11488 (N_11488,N_11220,N_11205);
or U11489 (N_11489,N_11148,N_11293);
nand U11490 (N_11490,N_11327,N_11355);
or U11491 (N_11491,N_11362,N_11231);
nand U11492 (N_11492,N_11268,N_11201);
nor U11493 (N_11493,N_11153,N_11361);
or U11494 (N_11494,N_11370,N_11329);
or U11495 (N_11495,N_11157,N_11144);
or U11496 (N_11496,N_11386,N_11247);
nor U11497 (N_11497,N_11112,N_11332);
nor U11498 (N_11498,N_11254,N_11111);
xnor U11499 (N_11499,N_11219,N_11141);
and U11500 (N_11500,N_11346,N_11256);
and U11501 (N_11501,N_11218,N_11238);
and U11502 (N_11502,N_11354,N_11379);
xor U11503 (N_11503,N_11230,N_11186);
nor U11504 (N_11504,N_11392,N_11373);
xor U11505 (N_11505,N_11183,N_11188);
xnor U11506 (N_11506,N_11164,N_11129);
nor U11507 (N_11507,N_11275,N_11384);
nand U11508 (N_11508,N_11172,N_11289);
or U11509 (N_11509,N_11360,N_11174);
nor U11510 (N_11510,N_11348,N_11224);
or U11511 (N_11511,N_11158,N_11339);
and U11512 (N_11512,N_11128,N_11312);
or U11513 (N_11513,N_11210,N_11297);
nor U11514 (N_11514,N_11377,N_11363);
xnor U11515 (N_11515,N_11105,N_11369);
nor U11516 (N_11516,N_11269,N_11390);
xor U11517 (N_11517,N_11310,N_11182);
xnor U11518 (N_11518,N_11313,N_11317);
and U11519 (N_11519,N_11226,N_11398);
and U11520 (N_11520,N_11194,N_11213);
xor U11521 (N_11521,N_11216,N_11276);
nor U11522 (N_11522,N_11252,N_11296);
nand U11523 (N_11523,N_11246,N_11227);
nor U11524 (N_11524,N_11136,N_11209);
nor U11525 (N_11525,N_11324,N_11263);
or U11526 (N_11526,N_11342,N_11333);
nand U11527 (N_11527,N_11343,N_11385);
nor U11528 (N_11528,N_11198,N_11309);
and U11529 (N_11529,N_11380,N_11122);
nor U11530 (N_11530,N_11352,N_11266);
and U11531 (N_11531,N_11156,N_11257);
nand U11532 (N_11532,N_11283,N_11314);
nor U11533 (N_11533,N_11206,N_11298);
and U11534 (N_11534,N_11284,N_11107);
nor U11535 (N_11535,N_11121,N_11124);
or U11536 (N_11536,N_11142,N_11152);
or U11537 (N_11537,N_11305,N_11336);
nor U11538 (N_11538,N_11189,N_11223);
nand U11539 (N_11539,N_11251,N_11349);
and U11540 (N_11540,N_11261,N_11117);
and U11541 (N_11541,N_11244,N_11353);
nor U11542 (N_11542,N_11288,N_11265);
xor U11543 (N_11543,N_11277,N_11278);
and U11544 (N_11544,N_11177,N_11228);
and U11545 (N_11545,N_11262,N_11375);
xor U11546 (N_11546,N_11145,N_11169);
nand U11547 (N_11547,N_11147,N_11245);
and U11548 (N_11548,N_11382,N_11150);
nor U11549 (N_11549,N_11143,N_11344);
nor U11550 (N_11550,N_11271,N_11140);
nand U11551 (N_11551,N_11138,N_11309);
xor U11552 (N_11552,N_11116,N_11342);
xor U11553 (N_11553,N_11240,N_11209);
nor U11554 (N_11554,N_11279,N_11119);
or U11555 (N_11555,N_11305,N_11316);
or U11556 (N_11556,N_11336,N_11232);
and U11557 (N_11557,N_11397,N_11386);
xor U11558 (N_11558,N_11111,N_11143);
nand U11559 (N_11559,N_11178,N_11130);
and U11560 (N_11560,N_11148,N_11106);
nor U11561 (N_11561,N_11177,N_11346);
xor U11562 (N_11562,N_11257,N_11212);
or U11563 (N_11563,N_11303,N_11184);
nor U11564 (N_11564,N_11171,N_11168);
and U11565 (N_11565,N_11327,N_11131);
nor U11566 (N_11566,N_11138,N_11159);
nand U11567 (N_11567,N_11177,N_11200);
or U11568 (N_11568,N_11240,N_11346);
xor U11569 (N_11569,N_11333,N_11372);
or U11570 (N_11570,N_11255,N_11377);
nor U11571 (N_11571,N_11166,N_11146);
or U11572 (N_11572,N_11154,N_11274);
nand U11573 (N_11573,N_11208,N_11115);
or U11574 (N_11574,N_11224,N_11375);
xor U11575 (N_11575,N_11195,N_11246);
or U11576 (N_11576,N_11171,N_11151);
nor U11577 (N_11577,N_11367,N_11217);
xor U11578 (N_11578,N_11259,N_11354);
and U11579 (N_11579,N_11204,N_11283);
nand U11580 (N_11580,N_11313,N_11192);
nor U11581 (N_11581,N_11258,N_11268);
or U11582 (N_11582,N_11360,N_11221);
or U11583 (N_11583,N_11364,N_11239);
or U11584 (N_11584,N_11359,N_11354);
nand U11585 (N_11585,N_11138,N_11121);
nor U11586 (N_11586,N_11245,N_11345);
or U11587 (N_11587,N_11335,N_11298);
or U11588 (N_11588,N_11234,N_11253);
or U11589 (N_11589,N_11143,N_11237);
nand U11590 (N_11590,N_11149,N_11233);
and U11591 (N_11591,N_11257,N_11316);
or U11592 (N_11592,N_11309,N_11178);
nand U11593 (N_11593,N_11176,N_11189);
xor U11594 (N_11594,N_11208,N_11193);
nand U11595 (N_11595,N_11241,N_11290);
xnor U11596 (N_11596,N_11221,N_11198);
xor U11597 (N_11597,N_11210,N_11139);
nor U11598 (N_11598,N_11289,N_11309);
and U11599 (N_11599,N_11107,N_11267);
and U11600 (N_11600,N_11317,N_11236);
nand U11601 (N_11601,N_11378,N_11365);
nand U11602 (N_11602,N_11149,N_11336);
xor U11603 (N_11603,N_11328,N_11369);
or U11604 (N_11604,N_11309,N_11274);
nor U11605 (N_11605,N_11303,N_11366);
nor U11606 (N_11606,N_11356,N_11240);
and U11607 (N_11607,N_11215,N_11262);
nand U11608 (N_11608,N_11195,N_11216);
nand U11609 (N_11609,N_11333,N_11353);
xor U11610 (N_11610,N_11154,N_11246);
xnor U11611 (N_11611,N_11381,N_11247);
nand U11612 (N_11612,N_11223,N_11216);
or U11613 (N_11613,N_11174,N_11380);
nand U11614 (N_11614,N_11398,N_11364);
nand U11615 (N_11615,N_11337,N_11177);
nor U11616 (N_11616,N_11211,N_11172);
nor U11617 (N_11617,N_11382,N_11214);
xnor U11618 (N_11618,N_11291,N_11175);
and U11619 (N_11619,N_11153,N_11327);
nand U11620 (N_11620,N_11298,N_11284);
or U11621 (N_11621,N_11254,N_11351);
nand U11622 (N_11622,N_11181,N_11268);
nor U11623 (N_11623,N_11234,N_11134);
nor U11624 (N_11624,N_11168,N_11158);
or U11625 (N_11625,N_11201,N_11264);
and U11626 (N_11626,N_11202,N_11166);
and U11627 (N_11627,N_11189,N_11102);
or U11628 (N_11628,N_11228,N_11392);
and U11629 (N_11629,N_11129,N_11391);
and U11630 (N_11630,N_11140,N_11135);
nor U11631 (N_11631,N_11326,N_11318);
and U11632 (N_11632,N_11378,N_11148);
nor U11633 (N_11633,N_11206,N_11340);
xor U11634 (N_11634,N_11385,N_11218);
xor U11635 (N_11635,N_11256,N_11393);
xor U11636 (N_11636,N_11354,N_11391);
and U11637 (N_11637,N_11199,N_11266);
or U11638 (N_11638,N_11391,N_11337);
nor U11639 (N_11639,N_11340,N_11339);
xnor U11640 (N_11640,N_11241,N_11314);
and U11641 (N_11641,N_11134,N_11369);
or U11642 (N_11642,N_11115,N_11364);
and U11643 (N_11643,N_11249,N_11301);
nor U11644 (N_11644,N_11373,N_11259);
and U11645 (N_11645,N_11371,N_11329);
nor U11646 (N_11646,N_11193,N_11366);
xnor U11647 (N_11647,N_11358,N_11216);
or U11648 (N_11648,N_11218,N_11300);
xor U11649 (N_11649,N_11216,N_11275);
xnor U11650 (N_11650,N_11316,N_11277);
and U11651 (N_11651,N_11393,N_11336);
and U11652 (N_11652,N_11345,N_11112);
and U11653 (N_11653,N_11130,N_11120);
or U11654 (N_11654,N_11398,N_11373);
nor U11655 (N_11655,N_11161,N_11107);
and U11656 (N_11656,N_11250,N_11236);
xor U11657 (N_11657,N_11144,N_11230);
nor U11658 (N_11658,N_11271,N_11261);
nor U11659 (N_11659,N_11307,N_11393);
nand U11660 (N_11660,N_11140,N_11217);
xor U11661 (N_11661,N_11264,N_11103);
nand U11662 (N_11662,N_11205,N_11170);
and U11663 (N_11663,N_11269,N_11344);
xnor U11664 (N_11664,N_11340,N_11328);
and U11665 (N_11665,N_11256,N_11230);
xor U11666 (N_11666,N_11131,N_11367);
nor U11667 (N_11667,N_11144,N_11155);
nor U11668 (N_11668,N_11134,N_11127);
xor U11669 (N_11669,N_11210,N_11104);
xor U11670 (N_11670,N_11300,N_11290);
nor U11671 (N_11671,N_11194,N_11160);
or U11672 (N_11672,N_11335,N_11371);
xnor U11673 (N_11673,N_11316,N_11204);
nor U11674 (N_11674,N_11142,N_11374);
or U11675 (N_11675,N_11262,N_11341);
nor U11676 (N_11676,N_11248,N_11321);
xnor U11677 (N_11677,N_11313,N_11180);
and U11678 (N_11678,N_11173,N_11313);
nor U11679 (N_11679,N_11167,N_11149);
nor U11680 (N_11680,N_11225,N_11375);
xnor U11681 (N_11681,N_11206,N_11338);
nand U11682 (N_11682,N_11241,N_11291);
xor U11683 (N_11683,N_11325,N_11182);
nand U11684 (N_11684,N_11375,N_11141);
xnor U11685 (N_11685,N_11384,N_11128);
xnor U11686 (N_11686,N_11243,N_11114);
nor U11687 (N_11687,N_11280,N_11218);
or U11688 (N_11688,N_11143,N_11139);
and U11689 (N_11689,N_11300,N_11205);
xnor U11690 (N_11690,N_11241,N_11386);
or U11691 (N_11691,N_11201,N_11305);
or U11692 (N_11692,N_11345,N_11362);
nor U11693 (N_11693,N_11337,N_11396);
and U11694 (N_11694,N_11352,N_11110);
xor U11695 (N_11695,N_11156,N_11228);
and U11696 (N_11696,N_11199,N_11189);
nor U11697 (N_11697,N_11303,N_11244);
nand U11698 (N_11698,N_11100,N_11262);
xor U11699 (N_11699,N_11241,N_11189);
or U11700 (N_11700,N_11466,N_11414);
or U11701 (N_11701,N_11649,N_11676);
xnor U11702 (N_11702,N_11537,N_11621);
or U11703 (N_11703,N_11441,N_11685);
nand U11704 (N_11704,N_11447,N_11540);
or U11705 (N_11705,N_11661,N_11642);
xnor U11706 (N_11706,N_11611,N_11574);
nor U11707 (N_11707,N_11511,N_11677);
nor U11708 (N_11708,N_11613,N_11525);
or U11709 (N_11709,N_11693,N_11630);
xnor U11710 (N_11710,N_11597,N_11549);
and U11711 (N_11711,N_11560,N_11485);
nand U11712 (N_11712,N_11631,N_11476);
nand U11713 (N_11713,N_11519,N_11694);
and U11714 (N_11714,N_11527,N_11581);
xnor U11715 (N_11715,N_11532,N_11451);
xnor U11716 (N_11716,N_11595,N_11641);
nand U11717 (N_11717,N_11552,N_11638);
and U11718 (N_11718,N_11425,N_11563);
nor U11719 (N_11719,N_11433,N_11696);
nor U11720 (N_11720,N_11573,N_11653);
xor U11721 (N_11721,N_11428,N_11583);
xor U11722 (N_11722,N_11697,N_11556);
and U11723 (N_11723,N_11550,N_11582);
and U11724 (N_11724,N_11543,N_11643);
nor U11725 (N_11725,N_11603,N_11413);
and U11726 (N_11726,N_11684,N_11673);
xnor U11727 (N_11727,N_11558,N_11486);
xor U11728 (N_11728,N_11571,N_11454);
or U11729 (N_11729,N_11546,N_11438);
nand U11730 (N_11730,N_11617,N_11623);
xnor U11731 (N_11731,N_11467,N_11610);
and U11732 (N_11732,N_11609,N_11406);
and U11733 (N_11733,N_11465,N_11488);
nor U11734 (N_11734,N_11509,N_11420);
nand U11735 (N_11735,N_11529,N_11660);
nor U11736 (N_11736,N_11615,N_11471);
nor U11737 (N_11737,N_11536,N_11645);
nand U11738 (N_11738,N_11477,N_11654);
nand U11739 (N_11739,N_11487,N_11589);
or U11740 (N_11740,N_11469,N_11481);
or U11741 (N_11741,N_11551,N_11491);
nand U11742 (N_11742,N_11568,N_11593);
xnor U11743 (N_11743,N_11699,N_11542);
nor U11744 (N_11744,N_11579,N_11590);
and U11745 (N_11745,N_11484,N_11691);
and U11746 (N_11746,N_11565,N_11600);
xor U11747 (N_11747,N_11668,N_11423);
or U11748 (N_11748,N_11671,N_11405);
nand U11749 (N_11749,N_11416,N_11427);
xor U11750 (N_11750,N_11401,N_11678);
nor U11751 (N_11751,N_11524,N_11458);
nand U11752 (N_11752,N_11497,N_11639);
and U11753 (N_11753,N_11470,N_11500);
or U11754 (N_11754,N_11652,N_11670);
xnor U11755 (N_11755,N_11584,N_11667);
and U11756 (N_11756,N_11429,N_11442);
nand U11757 (N_11757,N_11569,N_11503);
and U11758 (N_11758,N_11572,N_11690);
or U11759 (N_11759,N_11629,N_11612);
xnor U11760 (N_11760,N_11686,N_11426);
and U11761 (N_11761,N_11682,N_11403);
xnor U11762 (N_11762,N_11514,N_11459);
or U11763 (N_11763,N_11518,N_11580);
or U11764 (N_11764,N_11436,N_11555);
nand U11765 (N_11765,N_11695,N_11417);
xnor U11766 (N_11766,N_11530,N_11535);
nand U11767 (N_11767,N_11587,N_11679);
xnor U11768 (N_11768,N_11510,N_11544);
xor U11769 (N_11769,N_11460,N_11517);
nor U11770 (N_11770,N_11548,N_11462);
and U11771 (N_11771,N_11435,N_11541);
nor U11772 (N_11772,N_11404,N_11614);
nand U11773 (N_11773,N_11657,N_11501);
nand U11774 (N_11774,N_11650,N_11636);
nor U11775 (N_11775,N_11626,N_11431);
xnor U11776 (N_11776,N_11683,N_11473);
and U11777 (N_11777,N_11596,N_11412);
or U11778 (N_11778,N_11545,N_11424);
nor U11779 (N_11779,N_11616,N_11410);
nor U11780 (N_11780,N_11439,N_11482);
xnor U11781 (N_11781,N_11464,N_11437);
nor U11782 (N_11782,N_11434,N_11480);
and U11783 (N_11783,N_11674,N_11662);
or U11784 (N_11784,N_11498,N_11570);
xor U11785 (N_11785,N_11606,N_11578);
or U11786 (N_11786,N_11655,N_11504);
nor U11787 (N_11787,N_11452,N_11534);
xnor U11788 (N_11788,N_11496,N_11415);
nor U11789 (N_11789,N_11627,N_11506);
nand U11790 (N_11790,N_11647,N_11591);
nand U11791 (N_11791,N_11619,N_11522);
and U11792 (N_11792,N_11664,N_11687);
or U11793 (N_11793,N_11605,N_11648);
xor U11794 (N_11794,N_11494,N_11675);
or U11795 (N_11795,N_11402,N_11628);
nor U11796 (N_11796,N_11608,N_11656);
nand U11797 (N_11797,N_11586,N_11513);
nand U11798 (N_11798,N_11567,N_11561);
or U11799 (N_11799,N_11457,N_11502);
and U11800 (N_11800,N_11489,N_11456);
xor U11801 (N_11801,N_11472,N_11625);
xnor U11802 (N_11802,N_11411,N_11445);
xnor U11803 (N_11803,N_11577,N_11521);
nand U11804 (N_11804,N_11554,N_11499);
nor U11805 (N_11805,N_11520,N_11493);
and U11806 (N_11806,N_11508,N_11526);
nor U11807 (N_11807,N_11455,N_11419);
and U11808 (N_11808,N_11680,N_11468);
and U11809 (N_11809,N_11539,N_11632);
nor U11810 (N_11810,N_11599,N_11562);
nor U11811 (N_11811,N_11622,N_11634);
xor U11812 (N_11812,N_11478,N_11533);
nor U11813 (N_11813,N_11432,N_11620);
and U11814 (N_11814,N_11492,N_11444);
nand U11815 (N_11815,N_11483,N_11698);
nor U11816 (N_11816,N_11564,N_11618);
nor U11817 (N_11817,N_11495,N_11666);
nor U11818 (N_11818,N_11688,N_11449);
or U11819 (N_11819,N_11507,N_11576);
xnor U11820 (N_11820,N_11594,N_11559);
xor U11821 (N_11821,N_11400,N_11531);
and U11822 (N_11822,N_11646,N_11461);
and U11823 (N_11823,N_11692,N_11443);
and U11824 (N_11824,N_11505,N_11448);
and U11825 (N_11825,N_11624,N_11681);
or U11826 (N_11826,N_11588,N_11665);
nor U11827 (N_11827,N_11575,N_11602);
or U11828 (N_11828,N_11672,N_11658);
nand U11829 (N_11829,N_11598,N_11515);
nand U11830 (N_11830,N_11553,N_11409);
nand U11831 (N_11831,N_11516,N_11418);
xnor U11832 (N_11832,N_11689,N_11663);
and U11833 (N_11833,N_11479,N_11659);
xor U11834 (N_11834,N_11490,N_11446);
nand U11835 (N_11835,N_11407,N_11463);
or U11836 (N_11836,N_11538,N_11592);
nand U11837 (N_11837,N_11601,N_11633);
nand U11838 (N_11838,N_11453,N_11422);
or U11839 (N_11839,N_11585,N_11408);
and U11840 (N_11840,N_11644,N_11475);
or U11841 (N_11841,N_11607,N_11474);
or U11842 (N_11842,N_11523,N_11512);
xnor U11843 (N_11843,N_11547,N_11669);
or U11844 (N_11844,N_11430,N_11651);
and U11845 (N_11845,N_11440,N_11450);
nand U11846 (N_11846,N_11637,N_11421);
xor U11847 (N_11847,N_11604,N_11635);
or U11848 (N_11848,N_11557,N_11640);
and U11849 (N_11849,N_11566,N_11528);
nand U11850 (N_11850,N_11672,N_11507);
xor U11851 (N_11851,N_11642,N_11455);
and U11852 (N_11852,N_11413,N_11498);
xnor U11853 (N_11853,N_11434,N_11437);
xor U11854 (N_11854,N_11663,N_11685);
or U11855 (N_11855,N_11536,N_11559);
nand U11856 (N_11856,N_11583,N_11516);
or U11857 (N_11857,N_11471,N_11616);
or U11858 (N_11858,N_11625,N_11584);
or U11859 (N_11859,N_11404,N_11480);
or U11860 (N_11860,N_11681,N_11580);
or U11861 (N_11861,N_11568,N_11581);
or U11862 (N_11862,N_11406,N_11659);
and U11863 (N_11863,N_11445,N_11449);
nand U11864 (N_11864,N_11465,N_11697);
nand U11865 (N_11865,N_11452,N_11599);
nand U11866 (N_11866,N_11477,N_11627);
nand U11867 (N_11867,N_11609,N_11669);
xor U11868 (N_11868,N_11691,N_11689);
nand U11869 (N_11869,N_11410,N_11658);
nand U11870 (N_11870,N_11537,N_11595);
xor U11871 (N_11871,N_11512,N_11688);
nand U11872 (N_11872,N_11442,N_11488);
and U11873 (N_11873,N_11673,N_11442);
nor U11874 (N_11874,N_11626,N_11616);
and U11875 (N_11875,N_11491,N_11526);
xor U11876 (N_11876,N_11664,N_11565);
nand U11877 (N_11877,N_11470,N_11623);
or U11878 (N_11878,N_11522,N_11403);
nor U11879 (N_11879,N_11657,N_11650);
nand U11880 (N_11880,N_11453,N_11619);
nand U11881 (N_11881,N_11519,N_11412);
nor U11882 (N_11882,N_11656,N_11524);
and U11883 (N_11883,N_11432,N_11622);
xnor U11884 (N_11884,N_11545,N_11427);
or U11885 (N_11885,N_11675,N_11595);
or U11886 (N_11886,N_11610,N_11662);
or U11887 (N_11887,N_11655,N_11495);
xnor U11888 (N_11888,N_11660,N_11672);
or U11889 (N_11889,N_11633,N_11669);
nand U11890 (N_11890,N_11638,N_11525);
nor U11891 (N_11891,N_11584,N_11551);
or U11892 (N_11892,N_11582,N_11455);
nor U11893 (N_11893,N_11472,N_11597);
and U11894 (N_11894,N_11546,N_11521);
xor U11895 (N_11895,N_11525,N_11447);
nor U11896 (N_11896,N_11645,N_11624);
xor U11897 (N_11897,N_11692,N_11410);
nand U11898 (N_11898,N_11679,N_11493);
and U11899 (N_11899,N_11643,N_11685);
xnor U11900 (N_11900,N_11420,N_11479);
nand U11901 (N_11901,N_11563,N_11461);
and U11902 (N_11902,N_11650,N_11487);
nand U11903 (N_11903,N_11470,N_11481);
xor U11904 (N_11904,N_11550,N_11405);
and U11905 (N_11905,N_11427,N_11419);
nor U11906 (N_11906,N_11609,N_11551);
nand U11907 (N_11907,N_11460,N_11558);
xnor U11908 (N_11908,N_11433,N_11606);
nor U11909 (N_11909,N_11569,N_11402);
and U11910 (N_11910,N_11504,N_11472);
nand U11911 (N_11911,N_11443,N_11585);
or U11912 (N_11912,N_11650,N_11663);
nor U11913 (N_11913,N_11436,N_11535);
and U11914 (N_11914,N_11669,N_11517);
nand U11915 (N_11915,N_11693,N_11464);
xnor U11916 (N_11916,N_11411,N_11589);
nor U11917 (N_11917,N_11466,N_11510);
nor U11918 (N_11918,N_11653,N_11637);
xor U11919 (N_11919,N_11619,N_11649);
nand U11920 (N_11920,N_11637,N_11474);
or U11921 (N_11921,N_11534,N_11473);
xnor U11922 (N_11922,N_11534,N_11620);
and U11923 (N_11923,N_11693,N_11609);
and U11924 (N_11924,N_11482,N_11421);
or U11925 (N_11925,N_11645,N_11677);
or U11926 (N_11926,N_11661,N_11696);
xor U11927 (N_11927,N_11426,N_11555);
or U11928 (N_11928,N_11696,N_11428);
and U11929 (N_11929,N_11464,N_11565);
or U11930 (N_11930,N_11517,N_11409);
and U11931 (N_11931,N_11455,N_11452);
or U11932 (N_11932,N_11557,N_11625);
nand U11933 (N_11933,N_11456,N_11577);
xor U11934 (N_11934,N_11476,N_11518);
xnor U11935 (N_11935,N_11627,N_11432);
xnor U11936 (N_11936,N_11683,N_11427);
nor U11937 (N_11937,N_11611,N_11406);
xnor U11938 (N_11938,N_11593,N_11455);
and U11939 (N_11939,N_11655,N_11550);
and U11940 (N_11940,N_11570,N_11535);
nor U11941 (N_11941,N_11587,N_11561);
and U11942 (N_11942,N_11680,N_11402);
or U11943 (N_11943,N_11606,N_11531);
nand U11944 (N_11944,N_11565,N_11643);
xor U11945 (N_11945,N_11496,N_11416);
nand U11946 (N_11946,N_11620,N_11538);
nor U11947 (N_11947,N_11659,N_11592);
or U11948 (N_11948,N_11566,N_11654);
nand U11949 (N_11949,N_11592,N_11572);
and U11950 (N_11950,N_11497,N_11445);
or U11951 (N_11951,N_11678,N_11524);
xor U11952 (N_11952,N_11472,N_11603);
or U11953 (N_11953,N_11697,N_11566);
nand U11954 (N_11954,N_11589,N_11492);
and U11955 (N_11955,N_11673,N_11512);
or U11956 (N_11956,N_11636,N_11535);
nand U11957 (N_11957,N_11441,N_11496);
nand U11958 (N_11958,N_11607,N_11445);
nand U11959 (N_11959,N_11639,N_11606);
nor U11960 (N_11960,N_11452,N_11692);
xor U11961 (N_11961,N_11607,N_11487);
nor U11962 (N_11962,N_11461,N_11507);
and U11963 (N_11963,N_11499,N_11597);
xor U11964 (N_11964,N_11565,N_11435);
or U11965 (N_11965,N_11411,N_11414);
xor U11966 (N_11966,N_11477,N_11613);
nor U11967 (N_11967,N_11615,N_11683);
or U11968 (N_11968,N_11487,N_11494);
and U11969 (N_11969,N_11484,N_11672);
nand U11970 (N_11970,N_11625,N_11498);
nor U11971 (N_11971,N_11606,N_11505);
xnor U11972 (N_11972,N_11485,N_11520);
nor U11973 (N_11973,N_11511,N_11616);
or U11974 (N_11974,N_11567,N_11412);
nand U11975 (N_11975,N_11696,N_11497);
nand U11976 (N_11976,N_11561,N_11443);
or U11977 (N_11977,N_11649,N_11657);
nor U11978 (N_11978,N_11456,N_11418);
and U11979 (N_11979,N_11416,N_11584);
or U11980 (N_11980,N_11436,N_11651);
xnor U11981 (N_11981,N_11581,N_11446);
and U11982 (N_11982,N_11532,N_11540);
xor U11983 (N_11983,N_11625,N_11553);
xnor U11984 (N_11984,N_11608,N_11555);
xor U11985 (N_11985,N_11520,N_11602);
nand U11986 (N_11986,N_11586,N_11617);
xnor U11987 (N_11987,N_11483,N_11627);
or U11988 (N_11988,N_11547,N_11627);
or U11989 (N_11989,N_11674,N_11454);
nor U11990 (N_11990,N_11536,N_11466);
xor U11991 (N_11991,N_11579,N_11426);
and U11992 (N_11992,N_11629,N_11514);
nand U11993 (N_11993,N_11633,N_11483);
and U11994 (N_11994,N_11414,N_11663);
nand U11995 (N_11995,N_11486,N_11514);
and U11996 (N_11996,N_11437,N_11440);
or U11997 (N_11997,N_11566,N_11576);
and U11998 (N_11998,N_11411,N_11430);
nand U11999 (N_11999,N_11556,N_11437);
and U12000 (N_12000,N_11873,N_11800);
or U12001 (N_12001,N_11890,N_11821);
nor U12002 (N_12002,N_11768,N_11799);
or U12003 (N_12003,N_11989,N_11831);
and U12004 (N_12004,N_11816,N_11779);
or U12005 (N_12005,N_11752,N_11726);
and U12006 (N_12006,N_11881,N_11709);
and U12007 (N_12007,N_11967,N_11741);
or U12008 (N_12008,N_11785,N_11828);
or U12009 (N_12009,N_11913,N_11906);
or U12010 (N_12010,N_11946,N_11887);
xor U12011 (N_12011,N_11889,N_11791);
or U12012 (N_12012,N_11888,N_11736);
or U12013 (N_12013,N_11937,N_11815);
and U12014 (N_12014,N_11760,N_11842);
xor U12015 (N_12015,N_11823,N_11919);
nor U12016 (N_12016,N_11729,N_11928);
or U12017 (N_12017,N_11972,N_11879);
xor U12018 (N_12018,N_11774,N_11701);
nor U12019 (N_12019,N_11813,N_11744);
and U12020 (N_12020,N_11761,N_11820);
xnor U12021 (N_12021,N_11865,N_11924);
nand U12022 (N_12022,N_11720,N_11796);
nand U12023 (N_12023,N_11914,N_11978);
and U12024 (N_12024,N_11730,N_11893);
xor U12025 (N_12025,N_11804,N_11860);
xor U12026 (N_12026,N_11921,N_11737);
nand U12027 (N_12027,N_11925,N_11982);
and U12028 (N_12028,N_11704,N_11746);
nor U12029 (N_12029,N_11991,N_11735);
xor U12030 (N_12030,N_11973,N_11974);
and U12031 (N_12031,N_11712,N_11780);
or U12032 (N_12032,N_11975,N_11859);
or U12033 (N_12033,N_11909,N_11999);
xor U12034 (N_12034,N_11797,N_11874);
and U12035 (N_12035,N_11740,N_11944);
nand U12036 (N_12036,N_11771,N_11711);
xor U12037 (N_12037,N_11957,N_11886);
or U12038 (N_12038,N_11835,N_11903);
nand U12039 (N_12039,N_11722,N_11868);
and U12040 (N_12040,N_11824,N_11786);
or U12041 (N_12041,N_11856,N_11731);
nor U12042 (N_12042,N_11772,N_11794);
nor U12043 (N_12043,N_11995,N_11847);
and U12044 (N_12044,N_11819,N_11810);
or U12045 (N_12045,N_11969,N_11857);
or U12046 (N_12046,N_11979,N_11915);
nor U12047 (N_12047,N_11878,N_11802);
nand U12048 (N_12048,N_11728,N_11977);
nand U12049 (N_12049,N_11861,N_11808);
or U12050 (N_12050,N_11918,N_11814);
nand U12051 (N_12051,N_11725,N_11962);
nand U12052 (N_12052,N_11985,N_11745);
or U12053 (N_12053,N_11723,N_11826);
nor U12054 (N_12054,N_11756,N_11943);
xor U12055 (N_12055,N_11758,N_11992);
xnor U12056 (N_12056,N_11936,N_11922);
xnor U12057 (N_12057,N_11714,N_11951);
nand U12058 (N_12058,N_11777,N_11895);
and U12059 (N_12059,N_11930,N_11721);
or U12060 (N_12060,N_11883,N_11703);
and U12061 (N_12061,N_11852,N_11892);
or U12062 (N_12062,N_11894,N_11952);
or U12063 (N_12063,N_11884,N_11832);
xnor U12064 (N_12064,N_11834,N_11953);
and U12065 (N_12065,N_11920,N_11927);
xnor U12066 (N_12066,N_11983,N_11750);
nand U12067 (N_12067,N_11926,N_11940);
or U12068 (N_12068,N_11898,N_11837);
xor U12069 (N_12069,N_11980,N_11836);
or U12070 (N_12070,N_11717,N_11942);
and U12071 (N_12071,N_11792,N_11770);
nand U12072 (N_12072,N_11862,N_11965);
or U12073 (N_12073,N_11864,N_11742);
nor U12074 (N_12074,N_11912,N_11941);
and U12075 (N_12075,N_11964,N_11702);
nor U12076 (N_12076,N_11707,N_11773);
nand U12077 (N_12077,N_11904,N_11990);
and U12078 (N_12078,N_11870,N_11933);
or U12079 (N_12079,N_11748,N_11949);
xor U12080 (N_12080,N_11900,N_11775);
nand U12081 (N_12081,N_11759,N_11954);
and U12082 (N_12082,N_11955,N_11733);
nor U12083 (N_12083,N_11938,N_11948);
xnor U12084 (N_12084,N_11840,N_11896);
nor U12085 (N_12085,N_11769,N_11902);
xor U12086 (N_12086,N_11743,N_11963);
or U12087 (N_12087,N_11715,N_11970);
and U12088 (N_12088,N_11935,N_11917);
and U12089 (N_12089,N_11793,N_11986);
xnor U12090 (N_12090,N_11956,N_11907);
and U12091 (N_12091,N_11845,N_11945);
nand U12092 (N_12092,N_11809,N_11981);
nor U12093 (N_12093,N_11968,N_11825);
nor U12094 (N_12094,N_11848,N_11778);
nand U12095 (N_12095,N_11734,N_11781);
nand U12096 (N_12096,N_11776,N_11858);
and U12097 (N_12097,N_11899,N_11971);
and U12098 (N_12098,N_11706,N_11806);
and U12099 (N_12099,N_11783,N_11872);
nor U12100 (N_12100,N_11749,N_11976);
nor U12101 (N_12101,N_11908,N_11998);
xnor U12102 (N_12102,N_11716,N_11766);
and U12103 (N_12103,N_11798,N_11988);
xnor U12104 (N_12104,N_11724,N_11960);
xor U12105 (N_12105,N_11851,N_11854);
xor U12106 (N_12106,N_11747,N_11763);
or U12107 (N_12107,N_11853,N_11993);
xor U12108 (N_12108,N_11866,N_11867);
and U12109 (N_12109,N_11788,N_11996);
nand U12110 (N_12110,N_11830,N_11863);
or U12111 (N_12111,N_11710,N_11850);
or U12112 (N_12112,N_11891,N_11757);
or U12113 (N_12113,N_11910,N_11934);
xnor U12114 (N_12114,N_11923,N_11811);
xor U12115 (N_12115,N_11739,N_11876);
xor U12116 (N_12116,N_11829,N_11869);
nor U12117 (N_12117,N_11855,N_11875);
and U12118 (N_12118,N_11817,N_11961);
xor U12119 (N_12119,N_11751,N_11838);
xnor U12120 (N_12120,N_11987,N_11764);
nor U12121 (N_12121,N_11753,N_11932);
or U12122 (N_12122,N_11738,N_11966);
xor U12123 (N_12123,N_11877,N_11700);
and U12124 (N_12124,N_11885,N_11997);
or U12125 (N_12125,N_11790,N_11765);
nor U12126 (N_12126,N_11959,N_11841);
nor U12127 (N_12127,N_11822,N_11767);
xor U12128 (N_12128,N_11958,N_11801);
nand U12129 (N_12129,N_11827,N_11950);
nor U12130 (N_12130,N_11916,N_11929);
xor U12131 (N_12131,N_11846,N_11880);
or U12132 (N_12132,N_11719,N_11713);
xnor U12133 (N_12133,N_11984,N_11784);
or U12134 (N_12134,N_11833,N_11705);
or U12135 (N_12135,N_11805,N_11994);
nor U12136 (N_12136,N_11849,N_11755);
nor U12137 (N_12137,N_11843,N_11911);
or U12138 (N_12138,N_11882,N_11812);
xnor U12139 (N_12139,N_11708,N_11787);
nand U12140 (N_12140,N_11795,N_11727);
nor U12141 (N_12141,N_11818,N_11901);
and U12142 (N_12142,N_11947,N_11754);
or U12143 (N_12143,N_11718,N_11782);
or U12144 (N_12144,N_11789,N_11803);
nand U12145 (N_12145,N_11807,N_11931);
and U12146 (N_12146,N_11762,N_11897);
xnor U12147 (N_12147,N_11871,N_11939);
nor U12148 (N_12148,N_11905,N_11732);
or U12149 (N_12149,N_11844,N_11839);
xnor U12150 (N_12150,N_11864,N_11817);
xnor U12151 (N_12151,N_11916,N_11807);
xnor U12152 (N_12152,N_11997,N_11748);
nand U12153 (N_12153,N_11974,N_11943);
or U12154 (N_12154,N_11766,N_11802);
nand U12155 (N_12155,N_11838,N_11892);
nor U12156 (N_12156,N_11869,N_11778);
and U12157 (N_12157,N_11820,N_11900);
xor U12158 (N_12158,N_11822,N_11800);
nand U12159 (N_12159,N_11891,N_11852);
nor U12160 (N_12160,N_11968,N_11798);
and U12161 (N_12161,N_11958,N_11783);
or U12162 (N_12162,N_11787,N_11955);
xnor U12163 (N_12163,N_11788,N_11863);
nand U12164 (N_12164,N_11998,N_11792);
xor U12165 (N_12165,N_11775,N_11884);
nand U12166 (N_12166,N_11795,N_11902);
nor U12167 (N_12167,N_11859,N_11837);
and U12168 (N_12168,N_11744,N_11927);
or U12169 (N_12169,N_11831,N_11822);
or U12170 (N_12170,N_11860,N_11890);
or U12171 (N_12171,N_11728,N_11743);
nand U12172 (N_12172,N_11831,N_11817);
xor U12173 (N_12173,N_11814,N_11859);
or U12174 (N_12174,N_11943,N_11935);
nor U12175 (N_12175,N_11790,N_11961);
xnor U12176 (N_12176,N_11904,N_11835);
nand U12177 (N_12177,N_11767,N_11852);
nor U12178 (N_12178,N_11881,N_11878);
or U12179 (N_12179,N_11721,N_11706);
or U12180 (N_12180,N_11912,N_11773);
nor U12181 (N_12181,N_11902,N_11756);
nor U12182 (N_12182,N_11818,N_11783);
nand U12183 (N_12183,N_11918,N_11957);
and U12184 (N_12184,N_11775,N_11999);
xnor U12185 (N_12185,N_11867,N_11825);
nor U12186 (N_12186,N_11741,N_11826);
nand U12187 (N_12187,N_11947,N_11708);
nor U12188 (N_12188,N_11880,N_11931);
nor U12189 (N_12189,N_11910,N_11945);
nand U12190 (N_12190,N_11791,N_11933);
nor U12191 (N_12191,N_11821,N_11724);
nor U12192 (N_12192,N_11870,N_11729);
and U12193 (N_12193,N_11890,N_11764);
and U12194 (N_12194,N_11894,N_11962);
nand U12195 (N_12195,N_11908,N_11821);
xor U12196 (N_12196,N_11727,N_11959);
nor U12197 (N_12197,N_11975,N_11720);
and U12198 (N_12198,N_11915,N_11976);
xnor U12199 (N_12199,N_11765,N_11913);
or U12200 (N_12200,N_11778,N_11790);
and U12201 (N_12201,N_11949,N_11788);
and U12202 (N_12202,N_11794,N_11907);
or U12203 (N_12203,N_11854,N_11769);
or U12204 (N_12204,N_11789,N_11818);
or U12205 (N_12205,N_11812,N_11821);
and U12206 (N_12206,N_11803,N_11816);
or U12207 (N_12207,N_11797,N_11865);
xnor U12208 (N_12208,N_11998,N_11706);
or U12209 (N_12209,N_11803,N_11770);
xnor U12210 (N_12210,N_11700,N_11984);
nand U12211 (N_12211,N_11918,N_11770);
or U12212 (N_12212,N_11781,N_11854);
nor U12213 (N_12213,N_11985,N_11904);
nor U12214 (N_12214,N_11836,N_11744);
xnor U12215 (N_12215,N_11755,N_11889);
nor U12216 (N_12216,N_11752,N_11744);
nor U12217 (N_12217,N_11716,N_11743);
or U12218 (N_12218,N_11893,N_11882);
nand U12219 (N_12219,N_11858,N_11937);
or U12220 (N_12220,N_11895,N_11734);
and U12221 (N_12221,N_11813,N_11741);
nand U12222 (N_12222,N_11740,N_11753);
nor U12223 (N_12223,N_11787,N_11999);
nand U12224 (N_12224,N_11917,N_11948);
xor U12225 (N_12225,N_11972,N_11938);
nand U12226 (N_12226,N_11741,N_11955);
and U12227 (N_12227,N_11951,N_11881);
or U12228 (N_12228,N_11946,N_11755);
or U12229 (N_12229,N_11997,N_11750);
or U12230 (N_12230,N_11813,N_11851);
and U12231 (N_12231,N_11859,N_11990);
nand U12232 (N_12232,N_11811,N_11935);
and U12233 (N_12233,N_11732,N_11771);
nand U12234 (N_12234,N_11999,N_11819);
and U12235 (N_12235,N_11943,N_11867);
nand U12236 (N_12236,N_11877,N_11749);
xnor U12237 (N_12237,N_11730,N_11977);
and U12238 (N_12238,N_11935,N_11778);
or U12239 (N_12239,N_11914,N_11876);
nand U12240 (N_12240,N_11777,N_11782);
xor U12241 (N_12241,N_11818,N_11975);
nand U12242 (N_12242,N_11849,N_11747);
and U12243 (N_12243,N_11799,N_11999);
nand U12244 (N_12244,N_11744,N_11950);
or U12245 (N_12245,N_11888,N_11704);
nand U12246 (N_12246,N_11790,N_11933);
nand U12247 (N_12247,N_11816,N_11893);
or U12248 (N_12248,N_11731,N_11988);
nor U12249 (N_12249,N_11871,N_11787);
and U12250 (N_12250,N_11891,N_11915);
and U12251 (N_12251,N_11870,N_11847);
or U12252 (N_12252,N_11949,N_11730);
nand U12253 (N_12253,N_11743,N_11757);
or U12254 (N_12254,N_11919,N_11849);
or U12255 (N_12255,N_11791,N_11978);
nand U12256 (N_12256,N_11982,N_11821);
and U12257 (N_12257,N_11974,N_11959);
and U12258 (N_12258,N_11939,N_11824);
nor U12259 (N_12259,N_11887,N_11803);
or U12260 (N_12260,N_11935,N_11720);
nor U12261 (N_12261,N_11886,N_11792);
and U12262 (N_12262,N_11703,N_11755);
or U12263 (N_12263,N_11836,N_11833);
or U12264 (N_12264,N_11741,N_11995);
xor U12265 (N_12265,N_11718,N_11776);
or U12266 (N_12266,N_11749,N_11943);
xor U12267 (N_12267,N_11905,N_11726);
nor U12268 (N_12268,N_11790,N_11716);
nor U12269 (N_12269,N_11940,N_11959);
xnor U12270 (N_12270,N_11762,N_11939);
nand U12271 (N_12271,N_11929,N_11750);
nor U12272 (N_12272,N_11706,N_11886);
nand U12273 (N_12273,N_11759,N_11976);
nor U12274 (N_12274,N_11737,N_11980);
xnor U12275 (N_12275,N_11927,N_11928);
or U12276 (N_12276,N_11802,N_11900);
or U12277 (N_12277,N_11912,N_11712);
nand U12278 (N_12278,N_11757,N_11798);
xnor U12279 (N_12279,N_11751,N_11724);
nor U12280 (N_12280,N_11934,N_11957);
or U12281 (N_12281,N_11765,N_11923);
nand U12282 (N_12282,N_11719,N_11999);
or U12283 (N_12283,N_11879,N_11701);
xnor U12284 (N_12284,N_11971,N_11749);
xnor U12285 (N_12285,N_11868,N_11875);
and U12286 (N_12286,N_11970,N_11940);
nand U12287 (N_12287,N_11873,N_11778);
nand U12288 (N_12288,N_11736,N_11779);
xnor U12289 (N_12289,N_11963,N_11721);
or U12290 (N_12290,N_11803,N_11981);
or U12291 (N_12291,N_11929,N_11738);
and U12292 (N_12292,N_11965,N_11800);
nand U12293 (N_12293,N_11804,N_11858);
nor U12294 (N_12294,N_11810,N_11915);
nor U12295 (N_12295,N_11800,N_11723);
xnor U12296 (N_12296,N_11869,N_11985);
nand U12297 (N_12297,N_11912,N_11943);
and U12298 (N_12298,N_11758,N_11942);
and U12299 (N_12299,N_11722,N_11915);
or U12300 (N_12300,N_12026,N_12181);
nand U12301 (N_12301,N_12095,N_12076);
xor U12302 (N_12302,N_12242,N_12289);
nor U12303 (N_12303,N_12091,N_12213);
nor U12304 (N_12304,N_12121,N_12165);
nor U12305 (N_12305,N_12141,N_12147);
xnor U12306 (N_12306,N_12187,N_12068);
and U12307 (N_12307,N_12285,N_12084);
nand U12308 (N_12308,N_12249,N_12240);
nor U12309 (N_12309,N_12158,N_12299);
or U12310 (N_12310,N_12049,N_12042);
nand U12311 (N_12311,N_12111,N_12295);
nor U12312 (N_12312,N_12248,N_12170);
and U12313 (N_12313,N_12169,N_12216);
nor U12314 (N_12314,N_12260,N_12077);
nor U12315 (N_12315,N_12006,N_12236);
xnor U12316 (N_12316,N_12131,N_12264);
nor U12317 (N_12317,N_12228,N_12103);
xor U12318 (N_12318,N_12041,N_12258);
nand U12319 (N_12319,N_12254,N_12197);
or U12320 (N_12320,N_12100,N_12144);
xor U12321 (N_12321,N_12119,N_12220);
or U12322 (N_12322,N_12233,N_12276);
xor U12323 (N_12323,N_12027,N_12268);
and U12324 (N_12324,N_12073,N_12033);
nor U12325 (N_12325,N_12237,N_12206);
nor U12326 (N_12326,N_12174,N_12163);
and U12327 (N_12327,N_12140,N_12288);
nor U12328 (N_12328,N_12253,N_12192);
and U12329 (N_12329,N_12110,N_12136);
or U12330 (N_12330,N_12247,N_12129);
nand U12331 (N_12331,N_12018,N_12161);
nor U12332 (N_12332,N_12124,N_12164);
nor U12333 (N_12333,N_12062,N_12172);
or U12334 (N_12334,N_12244,N_12278);
xnor U12335 (N_12335,N_12135,N_12005);
and U12336 (N_12336,N_12117,N_12284);
and U12337 (N_12337,N_12120,N_12063);
nor U12338 (N_12338,N_12200,N_12231);
and U12339 (N_12339,N_12032,N_12191);
and U12340 (N_12340,N_12015,N_12051);
or U12341 (N_12341,N_12043,N_12024);
nor U12342 (N_12342,N_12105,N_12039);
nor U12343 (N_12343,N_12047,N_12019);
nor U12344 (N_12344,N_12167,N_12003);
or U12345 (N_12345,N_12186,N_12107);
and U12346 (N_12346,N_12149,N_12070);
or U12347 (N_12347,N_12229,N_12146);
nand U12348 (N_12348,N_12177,N_12035);
nor U12349 (N_12349,N_12023,N_12296);
and U12350 (N_12350,N_12160,N_12090);
nand U12351 (N_12351,N_12071,N_12016);
or U12352 (N_12352,N_12112,N_12209);
nor U12353 (N_12353,N_12065,N_12214);
xnor U12354 (N_12354,N_12223,N_12128);
and U12355 (N_12355,N_12145,N_12116);
and U12356 (N_12356,N_12044,N_12168);
nor U12357 (N_12357,N_12273,N_12226);
nand U12358 (N_12358,N_12277,N_12179);
xnor U12359 (N_12359,N_12234,N_12265);
xnor U12360 (N_12360,N_12297,N_12125);
nand U12361 (N_12361,N_12011,N_12182);
xnor U12362 (N_12362,N_12137,N_12086);
and U12363 (N_12363,N_12029,N_12053);
xor U12364 (N_12364,N_12020,N_12132);
or U12365 (N_12365,N_12245,N_12098);
xnor U12366 (N_12366,N_12250,N_12152);
nor U12367 (N_12367,N_12075,N_12217);
xor U12368 (N_12368,N_12055,N_12087);
xnor U12369 (N_12369,N_12287,N_12109);
or U12370 (N_12370,N_12008,N_12263);
and U12371 (N_12371,N_12238,N_12202);
nand U12372 (N_12372,N_12294,N_12183);
xnor U12373 (N_12373,N_12155,N_12166);
and U12374 (N_12374,N_12034,N_12219);
nand U12375 (N_12375,N_12002,N_12298);
xor U12376 (N_12376,N_12104,N_12004);
xnor U12377 (N_12377,N_12232,N_12143);
xnor U12378 (N_12378,N_12211,N_12162);
and U12379 (N_12379,N_12012,N_12227);
and U12380 (N_12380,N_12079,N_12082);
xnor U12381 (N_12381,N_12115,N_12282);
nor U12382 (N_12382,N_12218,N_12259);
or U12383 (N_12383,N_12126,N_12266);
xor U12384 (N_12384,N_12072,N_12052);
nor U12385 (N_12385,N_12099,N_12203);
xnor U12386 (N_12386,N_12185,N_12290);
nor U12387 (N_12387,N_12060,N_12272);
nand U12388 (N_12388,N_12198,N_12291);
nor U12389 (N_12389,N_12275,N_12134);
xor U12390 (N_12390,N_12207,N_12212);
xnor U12391 (N_12391,N_12093,N_12235);
or U12392 (N_12392,N_12114,N_12176);
nor U12393 (N_12393,N_12028,N_12215);
nand U12394 (N_12394,N_12036,N_12173);
nor U12395 (N_12395,N_12088,N_12222);
nor U12396 (N_12396,N_12180,N_12094);
and U12397 (N_12397,N_12097,N_12286);
nand U12398 (N_12398,N_12038,N_12083);
or U12399 (N_12399,N_12013,N_12118);
nand U12400 (N_12400,N_12138,N_12092);
xnor U12401 (N_12401,N_12050,N_12221);
and U12402 (N_12402,N_12127,N_12017);
nor U12403 (N_12403,N_12271,N_12096);
nand U12404 (N_12404,N_12054,N_12101);
or U12405 (N_12405,N_12113,N_12133);
and U12406 (N_12406,N_12059,N_12045);
nand U12407 (N_12407,N_12195,N_12014);
or U12408 (N_12408,N_12175,N_12267);
nand U12409 (N_12409,N_12066,N_12037);
nor U12410 (N_12410,N_12064,N_12102);
nand U12411 (N_12411,N_12021,N_12078);
xor U12412 (N_12412,N_12257,N_12061);
nor U12413 (N_12413,N_12190,N_12230);
and U12414 (N_12414,N_12293,N_12274);
nor U12415 (N_12415,N_12283,N_12178);
or U12416 (N_12416,N_12251,N_12153);
nor U12417 (N_12417,N_12031,N_12069);
and U12418 (N_12418,N_12193,N_12194);
nand U12419 (N_12419,N_12252,N_12046);
or U12420 (N_12420,N_12205,N_12081);
or U12421 (N_12421,N_12239,N_12139);
and U12422 (N_12422,N_12280,N_12156);
nand U12423 (N_12423,N_12001,N_12089);
nand U12424 (N_12424,N_12171,N_12000);
nor U12425 (N_12425,N_12058,N_12056);
nand U12426 (N_12426,N_12151,N_12269);
xnor U12427 (N_12427,N_12108,N_12189);
and U12428 (N_12428,N_12246,N_12281);
nand U12429 (N_12429,N_12085,N_12188);
nand U12430 (N_12430,N_12106,N_12201);
nor U12431 (N_12431,N_12007,N_12150);
or U12432 (N_12432,N_12148,N_12270);
and U12433 (N_12433,N_12224,N_12074);
and U12434 (N_12434,N_12080,N_12159);
nand U12435 (N_12435,N_12208,N_12010);
nor U12436 (N_12436,N_12057,N_12009);
nor U12437 (N_12437,N_12122,N_12184);
and U12438 (N_12438,N_12067,N_12256);
nor U12439 (N_12439,N_12279,N_12025);
nand U12440 (N_12440,N_12030,N_12225);
and U12441 (N_12441,N_12142,N_12243);
and U12442 (N_12442,N_12123,N_12040);
nand U12443 (N_12443,N_12241,N_12048);
nor U12444 (N_12444,N_12204,N_12261);
or U12445 (N_12445,N_12210,N_12262);
and U12446 (N_12446,N_12130,N_12199);
and U12447 (N_12447,N_12196,N_12157);
and U12448 (N_12448,N_12255,N_12292);
or U12449 (N_12449,N_12022,N_12154);
nor U12450 (N_12450,N_12221,N_12041);
xor U12451 (N_12451,N_12292,N_12074);
nor U12452 (N_12452,N_12027,N_12098);
xnor U12453 (N_12453,N_12060,N_12074);
nand U12454 (N_12454,N_12216,N_12152);
or U12455 (N_12455,N_12095,N_12064);
nor U12456 (N_12456,N_12084,N_12151);
nand U12457 (N_12457,N_12271,N_12210);
or U12458 (N_12458,N_12097,N_12185);
nor U12459 (N_12459,N_12122,N_12151);
and U12460 (N_12460,N_12126,N_12011);
nand U12461 (N_12461,N_12136,N_12211);
xnor U12462 (N_12462,N_12132,N_12176);
nand U12463 (N_12463,N_12067,N_12181);
or U12464 (N_12464,N_12070,N_12141);
nand U12465 (N_12465,N_12013,N_12009);
nand U12466 (N_12466,N_12260,N_12236);
and U12467 (N_12467,N_12028,N_12022);
or U12468 (N_12468,N_12071,N_12112);
nor U12469 (N_12469,N_12278,N_12023);
nor U12470 (N_12470,N_12203,N_12148);
nor U12471 (N_12471,N_12036,N_12125);
nand U12472 (N_12472,N_12090,N_12073);
nand U12473 (N_12473,N_12275,N_12282);
and U12474 (N_12474,N_12211,N_12222);
and U12475 (N_12475,N_12190,N_12185);
and U12476 (N_12476,N_12057,N_12276);
xnor U12477 (N_12477,N_12203,N_12265);
xnor U12478 (N_12478,N_12190,N_12099);
and U12479 (N_12479,N_12123,N_12252);
nor U12480 (N_12480,N_12085,N_12116);
or U12481 (N_12481,N_12074,N_12022);
nor U12482 (N_12482,N_12002,N_12063);
nor U12483 (N_12483,N_12017,N_12186);
nand U12484 (N_12484,N_12047,N_12038);
or U12485 (N_12485,N_12150,N_12151);
xnor U12486 (N_12486,N_12285,N_12021);
nor U12487 (N_12487,N_12054,N_12091);
nand U12488 (N_12488,N_12097,N_12099);
nand U12489 (N_12489,N_12262,N_12176);
nor U12490 (N_12490,N_12035,N_12182);
and U12491 (N_12491,N_12018,N_12060);
or U12492 (N_12492,N_12053,N_12222);
nand U12493 (N_12493,N_12103,N_12191);
or U12494 (N_12494,N_12279,N_12119);
or U12495 (N_12495,N_12239,N_12176);
nor U12496 (N_12496,N_12162,N_12186);
or U12497 (N_12497,N_12255,N_12166);
and U12498 (N_12498,N_12249,N_12293);
nand U12499 (N_12499,N_12060,N_12223);
xnor U12500 (N_12500,N_12237,N_12257);
nor U12501 (N_12501,N_12025,N_12054);
nor U12502 (N_12502,N_12280,N_12289);
nand U12503 (N_12503,N_12106,N_12094);
or U12504 (N_12504,N_12136,N_12084);
xnor U12505 (N_12505,N_12162,N_12025);
nor U12506 (N_12506,N_12140,N_12003);
or U12507 (N_12507,N_12204,N_12035);
nor U12508 (N_12508,N_12117,N_12137);
nand U12509 (N_12509,N_12213,N_12162);
nor U12510 (N_12510,N_12094,N_12086);
or U12511 (N_12511,N_12254,N_12099);
or U12512 (N_12512,N_12060,N_12090);
nor U12513 (N_12513,N_12083,N_12110);
and U12514 (N_12514,N_12088,N_12092);
and U12515 (N_12515,N_12272,N_12274);
nor U12516 (N_12516,N_12127,N_12282);
or U12517 (N_12517,N_12056,N_12245);
nand U12518 (N_12518,N_12075,N_12137);
and U12519 (N_12519,N_12255,N_12057);
or U12520 (N_12520,N_12269,N_12078);
or U12521 (N_12521,N_12025,N_12137);
nor U12522 (N_12522,N_12006,N_12091);
and U12523 (N_12523,N_12280,N_12178);
nor U12524 (N_12524,N_12219,N_12115);
nor U12525 (N_12525,N_12186,N_12098);
nor U12526 (N_12526,N_12208,N_12066);
and U12527 (N_12527,N_12086,N_12063);
or U12528 (N_12528,N_12075,N_12141);
nand U12529 (N_12529,N_12021,N_12182);
xnor U12530 (N_12530,N_12258,N_12220);
nor U12531 (N_12531,N_12274,N_12070);
xor U12532 (N_12532,N_12073,N_12177);
nor U12533 (N_12533,N_12120,N_12091);
xnor U12534 (N_12534,N_12182,N_12181);
or U12535 (N_12535,N_12140,N_12213);
nand U12536 (N_12536,N_12164,N_12219);
nor U12537 (N_12537,N_12254,N_12108);
nand U12538 (N_12538,N_12127,N_12018);
nand U12539 (N_12539,N_12183,N_12027);
xnor U12540 (N_12540,N_12173,N_12295);
nand U12541 (N_12541,N_12106,N_12235);
or U12542 (N_12542,N_12012,N_12135);
nand U12543 (N_12543,N_12034,N_12212);
and U12544 (N_12544,N_12063,N_12023);
xnor U12545 (N_12545,N_12115,N_12095);
and U12546 (N_12546,N_12046,N_12178);
nand U12547 (N_12547,N_12124,N_12271);
and U12548 (N_12548,N_12127,N_12191);
nand U12549 (N_12549,N_12118,N_12279);
or U12550 (N_12550,N_12241,N_12227);
nor U12551 (N_12551,N_12059,N_12086);
or U12552 (N_12552,N_12053,N_12233);
and U12553 (N_12553,N_12182,N_12149);
and U12554 (N_12554,N_12041,N_12031);
xnor U12555 (N_12555,N_12030,N_12241);
nand U12556 (N_12556,N_12141,N_12047);
xor U12557 (N_12557,N_12257,N_12140);
nor U12558 (N_12558,N_12279,N_12198);
nand U12559 (N_12559,N_12115,N_12108);
nor U12560 (N_12560,N_12098,N_12022);
nor U12561 (N_12561,N_12067,N_12008);
or U12562 (N_12562,N_12133,N_12085);
or U12563 (N_12563,N_12266,N_12008);
or U12564 (N_12564,N_12076,N_12124);
xnor U12565 (N_12565,N_12277,N_12178);
nand U12566 (N_12566,N_12225,N_12150);
nor U12567 (N_12567,N_12165,N_12285);
nor U12568 (N_12568,N_12257,N_12128);
nor U12569 (N_12569,N_12237,N_12179);
or U12570 (N_12570,N_12180,N_12226);
nand U12571 (N_12571,N_12087,N_12095);
nor U12572 (N_12572,N_12135,N_12297);
and U12573 (N_12573,N_12143,N_12156);
xor U12574 (N_12574,N_12165,N_12122);
and U12575 (N_12575,N_12137,N_12073);
xnor U12576 (N_12576,N_12271,N_12298);
and U12577 (N_12577,N_12235,N_12145);
and U12578 (N_12578,N_12192,N_12086);
or U12579 (N_12579,N_12183,N_12018);
and U12580 (N_12580,N_12132,N_12018);
xnor U12581 (N_12581,N_12230,N_12144);
nand U12582 (N_12582,N_12236,N_12218);
nand U12583 (N_12583,N_12008,N_12016);
xor U12584 (N_12584,N_12123,N_12251);
xor U12585 (N_12585,N_12047,N_12153);
and U12586 (N_12586,N_12190,N_12155);
and U12587 (N_12587,N_12217,N_12139);
xnor U12588 (N_12588,N_12063,N_12092);
and U12589 (N_12589,N_12074,N_12078);
and U12590 (N_12590,N_12110,N_12113);
nand U12591 (N_12591,N_12174,N_12290);
nand U12592 (N_12592,N_12018,N_12023);
nor U12593 (N_12593,N_12256,N_12252);
nor U12594 (N_12594,N_12288,N_12030);
nor U12595 (N_12595,N_12113,N_12146);
nand U12596 (N_12596,N_12137,N_12156);
or U12597 (N_12597,N_12239,N_12119);
or U12598 (N_12598,N_12155,N_12233);
or U12599 (N_12599,N_12247,N_12016);
xor U12600 (N_12600,N_12463,N_12413);
nor U12601 (N_12601,N_12348,N_12583);
nor U12602 (N_12602,N_12562,N_12330);
nor U12603 (N_12603,N_12527,N_12598);
xnor U12604 (N_12604,N_12590,N_12320);
nor U12605 (N_12605,N_12465,N_12381);
or U12606 (N_12606,N_12338,N_12452);
xor U12607 (N_12607,N_12444,N_12480);
xor U12608 (N_12608,N_12534,N_12363);
nor U12609 (N_12609,N_12579,N_12459);
and U12610 (N_12610,N_12325,N_12387);
or U12611 (N_12611,N_12508,N_12371);
xor U12612 (N_12612,N_12448,N_12585);
and U12613 (N_12613,N_12319,N_12567);
or U12614 (N_12614,N_12362,N_12396);
nor U12615 (N_12615,N_12344,N_12443);
xor U12616 (N_12616,N_12312,N_12592);
xor U12617 (N_12617,N_12536,N_12461);
or U12618 (N_12618,N_12565,N_12507);
or U12619 (N_12619,N_12324,N_12431);
nand U12620 (N_12620,N_12561,N_12424);
xnor U12621 (N_12621,N_12485,N_12403);
or U12622 (N_12622,N_12380,N_12449);
or U12623 (N_12623,N_12525,N_12394);
nand U12624 (N_12624,N_12315,N_12580);
and U12625 (N_12625,N_12535,N_12505);
nand U12626 (N_12626,N_12367,N_12372);
nor U12627 (N_12627,N_12593,N_12314);
or U12628 (N_12628,N_12430,N_12307);
nor U12629 (N_12629,N_12441,N_12386);
nor U12630 (N_12630,N_12342,N_12417);
or U12631 (N_12631,N_12486,N_12494);
nand U12632 (N_12632,N_12464,N_12478);
and U12633 (N_12633,N_12317,N_12309);
nor U12634 (N_12634,N_12341,N_12428);
and U12635 (N_12635,N_12421,N_12397);
or U12636 (N_12636,N_12333,N_12420);
and U12637 (N_12637,N_12569,N_12487);
or U12638 (N_12638,N_12356,N_12364);
or U12639 (N_12639,N_12543,N_12490);
and U12640 (N_12640,N_12301,N_12555);
and U12641 (N_12641,N_12369,N_12450);
nor U12642 (N_12642,N_12393,N_12438);
or U12643 (N_12643,N_12568,N_12492);
or U12644 (N_12644,N_12577,N_12326);
or U12645 (N_12645,N_12361,N_12586);
or U12646 (N_12646,N_12323,N_12336);
nor U12647 (N_12647,N_12349,N_12340);
or U12648 (N_12648,N_12538,N_12425);
xor U12649 (N_12649,N_12556,N_12500);
or U12650 (N_12650,N_12522,N_12451);
nand U12651 (N_12651,N_12318,N_12509);
nand U12652 (N_12652,N_12392,N_12405);
or U12653 (N_12653,N_12375,N_12533);
nor U12654 (N_12654,N_12594,N_12495);
nor U12655 (N_12655,N_12496,N_12512);
or U12656 (N_12656,N_12337,N_12359);
or U12657 (N_12657,N_12584,N_12322);
and U12658 (N_12658,N_12347,N_12378);
nor U12659 (N_12659,N_12304,N_12475);
xnor U12660 (N_12660,N_12571,N_12458);
or U12661 (N_12661,N_12373,N_12520);
xor U12662 (N_12662,N_12357,N_12557);
and U12663 (N_12663,N_12422,N_12541);
or U12664 (N_12664,N_12550,N_12412);
and U12665 (N_12665,N_12313,N_12334);
and U12666 (N_12666,N_12582,N_12532);
nor U12667 (N_12667,N_12454,N_12504);
and U12668 (N_12668,N_12546,N_12382);
nand U12669 (N_12669,N_12308,N_12379);
or U12670 (N_12670,N_12488,N_12368);
nor U12671 (N_12671,N_12406,N_12414);
nor U12672 (N_12672,N_12306,N_12433);
xnor U12673 (N_12673,N_12474,N_12399);
and U12674 (N_12674,N_12457,N_12531);
nand U12675 (N_12675,N_12491,N_12560);
xor U12676 (N_12676,N_12390,N_12552);
nor U12677 (N_12677,N_12513,N_12423);
and U12678 (N_12678,N_12553,N_12479);
or U12679 (N_12679,N_12370,N_12416);
nand U12680 (N_12680,N_12383,N_12332);
nand U12681 (N_12681,N_12503,N_12434);
or U12682 (N_12682,N_12551,N_12385);
or U12683 (N_12683,N_12411,N_12517);
nand U12684 (N_12684,N_12437,N_12483);
or U12685 (N_12685,N_12511,N_12400);
nor U12686 (N_12686,N_12366,N_12510);
xnor U12687 (N_12687,N_12542,N_12410);
nor U12688 (N_12688,N_12345,N_12502);
nand U12689 (N_12689,N_12576,N_12595);
xnor U12690 (N_12690,N_12559,N_12402);
and U12691 (N_12691,N_12499,N_12409);
or U12692 (N_12692,N_12581,N_12548);
and U12693 (N_12693,N_12388,N_12391);
and U12694 (N_12694,N_12300,N_12401);
nor U12695 (N_12695,N_12426,N_12456);
nor U12696 (N_12696,N_12482,N_12339);
nor U12697 (N_12697,N_12572,N_12305);
xor U12698 (N_12698,N_12429,N_12472);
and U12699 (N_12699,N_12516,N_12440);
xnor U12700 (N_12700,N_12526,N_12469);
nor U12701 (N_12701,N_12481,N_12321);
and U12702 (N_12702,N_12574,N_12597);
nor U12703 (N_12703,N_12419,N_12528);
xnor U12704 (N_12704,N_12343,N_12468);
nor U12705 (N_12705,N_12549,N_12493);
nand U12706 (N_12706,N_12303,N_12302);
xor U12707 (N_12707,N_12316,N_12596);
nor U12708 (N_12708,N_12365,N_12404);
xnor U12709 (N_12709,N_12374,N_12462);
nand U12710 (N_12710,N_12563,N_12453);
xor U12711 (N_12711,N_12427,N_12588);
and U12712 (N_12712,N_12418,N_12436);
and U12713 (N_12713,N_12435,N_12355);
or U12714 (N_12714,N_12376,N_12589);
nand U12715 (N_12715,N_12415,N_12477);
xnor U12716 (N_12716,N_12537,N_12529);
or U12717 (N_12717,N_12467,N_12329);
nor U12718 (N_12718,N_12439,N_12515);
xor U12719 (N_12719,N_12573,N_12311);
xnor U12720 (N_12720,N_12498,N_12335);
nor U12721 (N_12721,N_12484,N_12466);
nor U12722 (N_12722,N_12350,N_12497);
nand U12723 (N_12723,N_12389,N_12506);
or U12724 (N_12724,N_12599,N_12540);
and U12725 (N_12725,N_12518,N_12310);
nand U12726 (N_12726,N_12442,N_12460);
or U12727 (N_12727,N_12328,N_12360);
or U12728 (N_12728,N_12471,N_12558);
nor U12729 (N_12729,N_12570,N_12470);
nor U12730 (N_12730,N_12530,N_12407);
nand U12731 (N_12731,N_12544,N_12377);
and U12732 (N_12732,N_12346,N_12591);
and U12733 (N_12733,N_12587,N_12395);
and U12734 (N_12734,N_12566,N_12476);
nand U12735 (N_12735,N_12524,N_12519);
or U12736 (N_12736,N_12358,N_12352);
nand U12737 (N_12737,N_12523,N_12578);
and U12738 (N_12738,N_12514,N_12521);
xor U12739 (N_12739,N_12354,N_12501);
nor U12740 (N_12740,N_12547,N_12447);
nand U12741 (N_12741,N_12351,N_12489);
nor U12742 (N_12742,N_12384,N_12353);
xor U12743 (N_12743,N_12473,N_12331);
or U12744 (N_12744,N_12455,N_12539);
xnor U12745 (N_12745,N_12554,N_12432);
nor U12746 (N_12746,N_12408,N_12445);
and U12747 (N_12747,N_12545,N_12327);
or U12748 (N_12748,N_12564,N_12398);
xnor U12749 (N_12749,N_12446,N_12575);
and U12750 (N_12750,N_12483,N_12587);
nor U12751 (N_12751,N_12394,N_12581);
nor U12752 (N_12752,N_12411,N_12579);
or U12753 (N_12753,N_12492,N_12374);
and U12754 (N_12754,N_12426,N_12522);
and U12755 (N_12755,N_12321,N_12424);
or U12756 (N_12756,N_12336,N_12529);
nand U12757 (N_12757,N_12325,N_12573);
and U12758 (N_12758,N_12426,N_12457);
or U12759 (N_12759,N_12492,N_12513);
nand U12760 (N_12760,N_12411,N_12372);
nand U12761 (N_12761,N_12483,N_12595);
nor U12762 (N_12762,N_12521,N_12465);
nor U12763 (N_12763,N_12446,N_12503);
and U12764 (N_12764,N_12538,N_12351);
xor U12765 (N_12765,N_12406,N_12505);
xnor U12766 (N_12766,N_12563,N_12581);
nand U12767 (N_12767,N_12415,N_12551);
xnor U12768 (N_12768,N_12404,N_12495);
nand U12769 (N_12769,N_12456,N_12580);
nor U12770 (N_12770,N_12497,N_12507);
xor U12771 (N_12771,N_12543,N_12351);
or U12772 (N_12772,N_12391,N_12585);
xnor U12773 (N_12773,N_12466,N_12473);
nor U12774 (N_12774,N_12558,N_12394);
xor U12775 (N_12775,N_12510,N_12462);
and U12776 (N_12776,N_12506,N_12404);
or U12777 (N_12777,N_12439,N_12348);
nor U12778 (N_12778,N_12436,N_12440);
nor U12779 (N_12779,N_12341,N_12439);
nor U12780 (N_12780,N_12499,N_12598);
nor U12781 (N_12781,N_12513,N_12347);
or U12782 (N_12782,N_12499,N_12527);
nand U12783 (N_12783,N_12430,N_12524);
and U12784 (N_12784,N_12389,N_12561);
nor U12785 (N_12785,N_12565,N_12452);
and U12786 (N_12786,N_12573,N_12576);
nor U12787 (N_12787,N_12527,N_12466);
xor U12788 (N_12788,N_12324,N_12552);
nor U12789 (N_12789,N_12548,N_12380);
or U12790 (N_12790,N_12456,N_12490);
and U12791 (N_12791,N_12484,N_12305);
nor U12792 (N_12792,N_12340,N_12390);
xnor U12793 (N_12793,N_12307,N_12551);
nand U12794 (N_12794,N_12498,N_12323);
nand U12795 (N_12795,N_12493,N_12598);
xnor U12796 (N_12796,N_12473,N_12416);
nor U12797 (N_12797,N_12317,N_12336);
nor U12798 (N_12798,N_12538,N_12457);
and U12799 (N_12799,N_12432,N_12517);
xor U12800 (N_12800,N_12508,N_12496);
or U12801 (N_12801,N_12493,N_12599);
xnor U12802 (N_12802,N_12454,N_12551);
and U12803 (N_12803,N_12429,N_12452);
and U12804 (N_12804,N_12561,N_12452);
xor U12805 (N_12805,N_12599,N_12306);
and U12806 (N_12806,N_12452,N_12402);
nor U12807 (N_12807,N_12508,N_12595);
and U12808 (N_12808,N_12334,N_12441);
or U12809 (N_12809,N_12373,N_12442);
xor U12810 (N_12810,N_12399,N_12315);
and U12811 (N_12811,N_12530,N_12352);
and U12812 (N_12812,N_12354,N_12420);
or U12813 (N_12813,N_12501,N_12507);
nor U12814 (N_12814,N_12357,N_12568);
or U12815 (N_12815,N_12429,N_12500);
nor U12816 (N_12816,N_12532,N_12422);
and U12817 (N_12817,N_12527,N_12468);
xor U12818 (N_12818,N_12452,N_12417);
or U12819 (N_12819,N_12544,N_12376);
xnor U12820 (N_12820,N_12578,N_12383);
and U12821 (N_12821,N_12335,N_12528);
nor U12822 (N_12822,N_12510,N_12393);
xor U12823 (N_12823,N_12481,N_12519);
or U12824 (N_12824,N_12431,N_12570);
nor U12825 (N_12825,N_12347,N_12317);
or U12826 (N_12826,N_12436,N_12562);
xor U12827 (N_12827,N_12351,N_12488);
xor U12828 (N_12828,N_12547,N_12583);
nor U12829 (N_12829,N_12573,N_12447);
nor U12830 (N_12830,N_12545,N_12301);
nor U12831 (N_12831,N_12583,N_12538);
nand U12832 (N_12832,N_12454,N_12346);
xnor U12833 (N_12833,N_12345,N_12416);
and U12834 (N_12834,N_12482,N_12542);
or U12835 (N_12835,N_12422,N_12323);
nor U12836 (N_12836,N_12538,N_12529);
xnor U12837 (N_12837,N_12522,N_12582);
xor U12838 (N_12838,N_12357,N_12573);
nor U12839 (N_12839,N_12446,N_12304);
nor U12840 (N_12840,N_12372,N_12518);
nand U12841 (N_12841,N_12317,N_12405);
xor U12842 (N_12842,N_12378,N_12374);
xnor U12843 (N_12843,N_12523,N_12472);
and U12844 (N_12844,N_12528,N_12537);
or U12845 (N_12845,N_12458,N_12450);
nor U12846 (N_12846,N_12443,N_12386);
nor U12847 (N_12847,N_12473,N_12556);
nor U12848 (N_12848,N_12453,N_12342);
and U12849 (N_12849,N_12546,N_12576);
nor U12850 (N_12850,N_12580,N_12474);
nand U12851 (N_12851,N_12451,N_12454);
and U12852 (N_12852,N_12385,N_12453);
xnor U12853 (N_12853,N_12313,N_12336);
and U12854 (N_12854,N_12341,N_12416);
or U12855 (N_12855,N_12378,N_12581);
nand U12856 (N_12856,N_12413,N_12348);
xor U12857 (N_12857,N_12555,N_12339);
or U12858 (N_12858,N_12538,N_12423);
xnor U12859 (N_12859,N_12503,N_12511);
or U12860 (N_12860,N_12566,N_12300);
nand U12861 (N_12861,N_12395,N_12380);
or U12862 (N_12862,N_12549,N_12367);
xor U12863 (N_12863,N_12442,N_12311);
xor U12864 (N_12864,N_12543,N_12368);
or U12865 (N_12865,N_12352,N_12480);
or U12866 (N_12866,N_12598,N_12378);
and U12867 (N_12867,N_12311,N_12547);
nand U12868 (N_12868,N_12335,N_12598);
nor U12869 (N_12869,N_12557,N_12353);
and U12870 (N_12870,N_12327,N_12330);
nand U12871 (N_12871,N_12416,N_12365);
nor U12872 (N_12872,N_12516,N_12348);
and U12873 (N_12873,N_12458,N_12477);
or U12874 (N_12874,N_12485,N_12307);
or U12875 (N_12875,N_12585,N_12326);
nor U12876 (N_12876,N_12547,N_12588);
nor U12877 (N_12877,N_12557,N_12498);
xor U12878 (N_12878,N_12378,N_12550);
nor U12879 (N_12879,N_12594,N_12352);
and U12880 (N_12880,N_12404,N_12352);
or U12881 (N_12881,N_12412,N_12599);
or U12882 (N_12882,N_12526,N_12505);
nor U12883 (N_12883,N_12499,N_12498);
nor U12884 (N_12884,N_12536,N_12386);
xnor U12885 (N_12885,N_12312,N_12402);
or U12886 (N_12886,N_12325,N_12578);
xnor U12887 (N_12887,N_12584,N_12466);
nand U12888 (N_12888,N_12423,N_12320);
and U12889 (N_12889,N_12556,N_12499);
xnor U12890 (N_12890,N_12360,N_12509);
nand U12891 (N_12891,N_12321,N_12476);
xnor U12892 (N_12892,N_12597,N_12496);
nand U12893 (N_12893,N_12375,N_12418);
and U12894 (N_12894,N_12581,N_12528);
nor U12895 (N_12895,N_12582,N_12442);
nor U12896 (N_12896,N_12434,N_12381);
nor U12897 (N_12897,N_12452,N_12323);
nor U12898 (N_12898,N_12548,N_12309);
nand U12899 (N_12899,N_12514,N_12346);
nor U12900 (N_12900,N_12810,N_12884);
xnor U12901 (N_12901,N_12898,N_12638);
and U12902 (N_12902,N_12658,N_12762);
nor U12903 (N_12903,N_12686,N_12604);
or U12904 (N_12904,N_12792,N_12794);
or U12905 (N_12905,N_12709,N_12789);
nor U12906 (N_12906,N_12832,N_12679);
and U12907 (N_12907,N_12728,N_12715);
nand U12908 (N_12908,N_12678,N_12666);
nand U12909 (N_12909,N_12739,N_12886);
nand U12910 (N_12910,N_12890,N_12719);
or U12911 (N_12911,N_12615,N_12864);
nand U12912 (N_12912,N_12616,N_12773);
nand U12913 (N_12913,N_12816,N_12871);
xnor U12914 (N_12914,N_12880,N_12836);
nor U12915 (N_12915,N_12701,N_12878);
xor U12916 (N_12916,N_12869,N_12748);
xor U12917 (N_12917,N_12820,N_12895);
xor U12918 (N_12918,N_12600,N_12607);
and U12919 (N_12919,N_12841,N_12775);
xor U12920 (N_12920,N_12851,N_12778);
and U12921 (N_12921,N_12606,N_12687);
and U12922 (N_12922,N_12807,N_12843);
nand U12923 (N_12923,N_12741,N_12763);
nand U12924 (N_12924,N_12743,N_12642);
nor U12925 (N_12925,N_12611,N_12722);
or U12926 (N_12926,N_12625,N_12784);
or U12927 (N_12927,N_12894,N_12873);
nand U12928 (N_12928,N_12724,N_12704);
xnor U12929 (N_12929,N_12755,N_12867);
xor U12930 (N_12930,N_12854,N_12729);
and U12931 (N_12931,N_12791,N_12747);
and U12932 (N_12932,N_12824,N_12602);
or U12933 (N_12933,N_12635,N_12840);
xor U12934 (N_12934,N_12689,N_12786);
nand U12935 (N_12935,N_12746,N_12696);
nor U12936 (N_12936,N_12835,N_12753);
nand U12937 (N_12937,N_12812,N_12779);
xnor U12938 (N_12938,N_12769,N_12668);
and U12939 (N_12939,N_12756,N_12818);
xnor U12940 (N_12940,N_12656,N_12688);
nor U12941 (N_12941,N_12819,N_12623);
and U12942 (N_12942,N_12630,N_12661);
or U12943 (N_12943,N_12727,N_12676);
or U12944 (N_12944,N_12817,N_12723);
or U12945 (N_12945,N_12643,N_12694);
nand U12946 (N_12946,N_12777,N_12655);
xor U12947 (N_12947,N_12830,N_12874);
and U12948 (N_12948,N_12647,N_12706);
nand U12949 (N_12949,N_12750,N_12761);
or U12950 (N_12950,N_12669,N_12781);
or U12951 (N_12951,N_12870,N_12813);
xnor U12952 (N_12952,N_12881,N_12716);
xnor U12953 (N_12953,N_12680,N_12752);
nor U12954 (N_12954,N_12685,N_12758);
or U12955 (N_12955,N_12603,N_12788);
and U12956 (N_12956,N_12660,N_12738);
nand U12957 (N_12957,N_12757,N_12751);
and U12958 (N_12958,N_12613,N_12866);
nor U12959 (N_12959,N_12713,N_12766);
nand U12960 (N_12960,N_12828,N_12842);
nor U12961 (N_12961,N_12804,N_12834);
and U12962 (N_12962,N_12649,N_12740);
nand U12963 (N_12963,N_12802,N_12673);
and U12964 (N_12964,N_12768,N_12754);
and U12965 (N_12965,N_12601,N_12893);
and U12966 (N_12966,N_12826,N_12891);
xnor U12967 (N_12967,N_12849,N_12693);
or U12968 (N_12968,N_12672,N_12897);
or U12969 (N_12969,N_12675,N_12862);
xor U12970 (N_12970,N_12695,N_12733);
or U12971 (N_12971,N_12806,N_12651);
and U12972 (N_12972,N_12707,N_12609);
xor U12973 (N_12973,N_12646,N_12805);
xnor U12974 (N_12974,N_12861,N_12872);
and U12975 (N_12975,N_12684,N_12650);
xor U12976 (N_12976,N_12865,N_12850);
xnor U12977 (N_12977,N_12896,N_12749);
or U12978 (N_12978,N_12774,N_12618);
and U12979 (N_12979,N_12662,N_12797);
or U12980 (N_12980,N_12714,N_12608);
and U12981 (N_12981,N_12814,N_12720);
or U12982 (N_12982,N_12620,N_12783);
nor U12983 (N_12983,N_12730,N_12859);
or U12984 (N_12984,N_12780,N_12795);
or U12985 (N_12985,N_12882,N_12736);
nand U12986 (N_12986,N_12631,N_12782);
nand U12987 (N_12987,N_12644,N_12735);
nor U12988 (N_12988,N_12856,N_12888);
or U12989 (N_12989,N_12622,N_12863);
nand U12990 (N_12990,N_12628,N_12674);
and U12991 (N_12991,N_12760,N_12653);
and U12992 (N_12992,N_12648,N_12692);
and U12993 (N_12993,N_12876,N_12892);
or U12994 (N_12994,N_12833,N_12665);
and U12995 (N_12995,N_12737,N_12699);
and U12996 (N_12996,N_12839,N_12772);
and U12997 (N_12997,N_12800,N_12857);
nand U12998 (N_12998,N_12776,N_12825);
and U12999 (N_12999,N_12711,N_12732);
nand U13000 (N_13000,N_12659,N_12845);
nand U13001 (N_13001,N_12744,N_12629);
and U13002 (N_13002,N_12612,N_12617);
and U13003 (N_13003,N_12670,N_12633);
and U13004 (N_13004,N_12858,N_12848);
and U13005 (N_13005,N_12889,N_12877);
nor U13006 (N_13006,N_12703,N_12799);
nor U13007 (N_13007,N_12624,N_12634);
xor U13008 (N_13008,N_12831,N_12705);
xnor U13009 (N_13009,N_12690,N_12726);
nand U13010 (N_13010,N_12664,N_12700);
or U13011 (N_13011,N_12852,N_12847);
xor U13012 (N_13012,N_12627,N_12637);
nand U13013 (N_13013,N_12667,N_12767);
and U13014 (N_13014,N_12641,N_12811);
nor U13015 (N_13015,N_12803,N_12745);
and U13016 (N_13016,N_12793,N_12682);
xnor U13017 (N_13017,N_12887,N_12734);
and U13018 (N_13018,N_12626,N_12885);
xor U13019 (N_13019,N_12614,N_12710);
nand U13020 (N_13020,N_12663,N_12771);
and U13021 (N_13021,N_12636,N_12712);
nor U13022 (N_13022,N_12731,N_12821);
nor U13023 (N_13023,N_12822,N_12785);
or U13024 (N_13024,N_12798,N_12742);
xor U13025 (N_13025,N_12605,N_12765);
nand U13026 (N_13026,N_12632,N_12671);
or U13027 (N_13027,N_12837,N_12621);
nand U13028 (N_13028,N_12639,N_12759);
xor U13029 (N_13029,N_12815,N_12691);
or U13030 (N_13030,N_12610,N_12827);
or U13031 (N_13031,N_12899,N_12883);
nor U13032 (N_13032,N_12721,N_12860);
or U13033 (N_13033,N_12640,N_12853);
xor U13034 (N_13034,N_12868,N_12619);
and U13035 (N_13035,N_12764,N_12787);
or U13036 (N_13036,N_12879,N_12846);
and U13037 (N_13037,N_12698,N_12770);
and U13038 (N_13038,N_12808,N_12829);
or U13039 (N_13039,N_12838,N_12654);
nor U13040 (N_13040,N_12875,N_12708);
or U13041 (N_13041,N_12809,N_12717);
nand U13042 (N_13042,N_12718,N_12823);
or U13043 (N_13043,N_12844,N_12801);
nor U13044 (N_13044,N_12677,N_12683);
nor U13045 (N_13045,N_12725,N_12645);
xnor U13046 (N_13046,N_12790,N_12652);
nand U13047 (N_13047,N_12681,N_12697);
xor U13048 (N_13048,N_12796,N_12657);
nor U13049 (N_13049,N_12855,N_12702);
xor U13050 (N_13050,N_12888,N_12799);
nor U13051 (N_13051,N_12612,N_12668);
and U13052 (N_13052,N_12688,N_12705);
xor U13053 (N_13053,N_12702,N_12818);
nor U13054 (N_13054,N_12771,N_12719);
nand U13055 (N_13055,N_12759,N_12751);
and U13056 (N_13056,N_12814,N_12733);
nor U13057 (N_13057,N_12612,N_12834);
nor U13058 (N_13058,N_12852,N_12833);
nand U13059 (N_13059,N_12824,N_12640);
and U13060 (N_13060,N_12707,N_12616);
xor U13061 (N_13061,N_12761,N_12642);
nor U13062 (N_13062,N_12609,N_12888);
xnor U13063 (N_13063,N_12766,N_12602);
nand U13064 (N_13064,N_12721,N_12727);
and U13065 (N_13065,N_12674,N_12660);
nand U13066 (N_13066,N_12856,N_12717);
nor U13067 (N_13067,N_12744,N_12749);
xnor U13068 (N_13068,N_12771,N_12866);
xor U13069 (N_13069,N_12732,N_12794);
nand U13070 (N_13070,N_12660,N_12841);
nor U13071 (N_13071,N_12843,N_12638);
or U13072 (N_13072,N_12885,N_12803);
and U13073 (N_13073,N_12791,N_12695);
nand U13074 (N_13074,N_12607,N_12738);
or U13075 (N_13075,N_12637,N_12765);
and U13076 (N_13076,N_12728,N_12719);
and U13077 (N_13077,N_12749,N_12761);
xor U13078 (N_13078,N_12600,N_12739);
and U13079 (N_13079,N_12848,N_12673);
or U13080 (N_13080,N_12760,N_12744);
xnor U13081 (N_13081,N_12818,N_12815);
and U13082 (N_13082,N_12738,N_12875);
and U13083 (N_13083,N_12818,N_12634);
xor U13084 (N_13084,N_12854,N_12708);
nor U13085 (N_13085,N_12737,N_12886);
nand U13086 (N_13086,N_12811,N_12602);
and U13087 (N_13087,N_12688,N_12651);
and U13088 (N_13088,N_12790,N_12895);
nor U13089 (N_13089,N_12675,N_12824);
nor U13090 (N_13090,N_12686,N_12651);
xnor U13091 (N_13091,N_12845,N_12640);
or U13092 (N_13092,N_12850,N_12711);
nand U13093 (N_13093,N_12744,N_12877);
xor U13094 (N_13094,N_12747,N_12765);
and U13095 (N_13095,N_12894,N_12854);
xnor U13096 (N_13096,N_12797,N_12884);
and U13097 (N_13097,N_12805,N_12624);
xnor U13098 (N_13098,N_12790,N_12830);
nand U13099 (N_13099,N_12707,N_12738);
nor U13100 (N_13100,N_12615,N_12707);
and U13101 (N_13101,N_12762,N_12740);
nand U13102 (N_13102,N_12662,N_12684);
nor U13103 (N_13103,N_12825,N_12645);
or U13104 (N_13104,N_12821,N_12887);
nor U13105 (N_13105,N_12695,N_12661);
xnor U13106 (N_13106,N_12764,N_12833);
and U13107 (N_13107,N_12802,N_12779);
xnor U13108 (N_13108,N_12677,N_12847);
and U13109 (N_13109,N_12722,N_12717);
and U13110 (N_13110,N_12831,N_12833);
xnor U13111 (N_13111,N_12799,N_12722);
and U13112 (N_13112,N_12867,N_12696);
and U13113 (N_13113,N_12682,N_12614);
xor U13114 (N_13114,N_12619,N_12846);
nor U13115 (N_13115,N_12604,N_12767);
nor U13116 (N_13116,N_12641,N_12773);
nor U13117 (N_13117,N_12834,N_12750);
and U13118 (N_13118,N_12634,N_12747);
and U13119 (N_13119,N_12654,N_12873);
xor U13120 (N_13120,N_12716,N_12778);
nor U13121 (N_13121,N_12849,N_12603);
or U13122 (N_13122,N_12807,N_12633);
or U13123 (N_13123,N_12600,N_12854);
or U13124 (N_13124,N_12624,N_12864);
xor U13125 (N_13125,N_12752,N_12861);
nor U13126 (N_13126,N_12686,N_12717);
nor U13127 (N_13127,N_12728,N_12638);
and U13128 (N_13128,N_12853,N_12706);
nor U13129 (N_13129,N_12732,N_12601);
nor U13130 (N_13130,N_12697,N_12648);
nand U13131 (N_13131,N_12649,N_12721);
and U13132 (N_13132,N_12778,N_12727);
and U13133 (N_13133,N_12729,N_12807);
nor U13134 (N_13134,N_12634,N_12712);
and U13135 (N_13135,N_12652,N_12887);
nand U13136 (N_13136,N_12811,N_12726);
xnor U13137 (N_13137,N_12746,N_12758);
nor U13138 (N_13138,N_12893,N_12758);
and U13139 (N_13139,N_12635,N_12697);
nor U13140 (N_13140,N_12600,N_12788);
xor U13141 (N_13141,N_12861,N_12804);
xnor U13142 (N_13142,N_12663,N_12719);
xnor U13143 (N_13143,N_12656,N_12609);
xor U13144 (N_13144,N_12686,N_12657);
and U13145 (N_13145,N_12736,N_12892);
or U13146 (N_13146,N_12641,N_12752);
or U13147 (N_13147,N_12700,N_12832);
nor U13148 (N_13148,N_12612,N_12775);
and U13149 (N_13149,N_12770,N_12783);
xor U13150 (N_13150,N_12728,N_12852);
and U13151 (N_13151,N_12689,N_12863);
nor U13152 (N_13152,N_12605,N_12667);
or U13153 (N_13153,N_12651,N_12748);
xnor U13154 (N_13154,N_12788,N_12891);
xnor U13155 (N_13155,N_12809,N_12605);
or U13156 (N_13156,N_12894,N_12783);
and U13157 (N_13157,N_12608,N_12610);
xnor U13158 (N_13158,N_12608,N_12888);
nand U13159 (N_13159,N_12691,N_12616);
xnor U13160 (N_13160,N_12746,N_12682);
xor U13161 (N_13161,N_12713,N_12723);
nand U13162 (N_13162,N_12607,N_12852);
or U13163 (N_13163,N_12825,N_12871);
or U13164 (N_13164,N_12878,N_12712);
nor U13165 (N_13165,N_12688,N_12621);
and U13166 (N_13166,N_12634,N_12737);
or U13167 (N_13167,N_12810,N_12724);
and U13168 (N_13168,N_12713,N_12604);
nor U13169 (N_13169,N_12678,N_12760);
nand U13170 (N_13170,N_12856,N_12854);
xor U13171 (N_13171,N_12689,N_12765);
or U13172 (N_13172,N_12635,N_12703);
and U13173 (N_13173,N_12744,N_12600);
nor U13174 (N_13174,N_12708,N_12690);
nand U13175 (N_13175,N_12744,N_12818);
xnor U13176 (N_13176,N_12783,N_12766);
or U13177 (N_13177,N_12738,N_12860);
nand U13178 (N_13178,N_12853,N_12798);
xor U13179 (N_13179,N_12662,N_12762);
xor U13180 (N_13180,N_12610,N_12677);
nor U13181 (N_13181,N_12805,N_12788);
nand U13182 (N_13182,N_12863,N_12866);
and U13183 (N_13183,N_12895,N_12893);
and U13184 (N_13184,N_12762,N_12705);
or U13185 (N_13185,N_12859,N_12649);
nor U13186 (N_13186,N_12798,N_12675);
or U13187 (N_13187,N_12753,N_12814);
nand U13188 (N_13188,N_12892,N_12696);
xor U13189 (N_13189,N_12728,N_12888);
or U13190 (N_13190,N_12722,N_12616);
nand U13191 (N_13191,N_12843,N_12792);
or U13192 (N_13192,N_12892,N_12738);
nand U13193 (N_13193,N_12733,N_12887);
or U13194 (N_13194,N_12772,N_12761);
nand U13195 (N_13195,N_12790,N_12892);
xnor U13196 (N_13196,N_12765,N_12664);
xnor U13197 (N_13197,N_12775,N_12708);
or U13198 (N_13198,N_12865,N_12827);
and U13199 (N_13199,N_12774,N_12643);
nor U13200 (N_13200,N_13174,N_13106);
or U13201 (N_13201,N_13116,N_13166);
and U13202 (N_13202,N_13057,N_13175);
and U13203 (N_13203,N_13115,N_13038);
or U13204 (N_13204,N_13156,N_13194);
or U13205 (N_13205,N_13046,N_13125);
and U13206 (N_13206,N_13127,N_13162);
nor U13207 (N_13207,N_13058,N_12967);
xor U13208 (N_13208,N_12974,N_12933);
nand U13209 (N_13209,N_13160,N_13149);
or U13210 (N_13210,N_13132,N_13075);
xor U13211 (N_13211,N_12906,N_12916);
nand U13212 (N_13212,N_13150,N_13024);
nand U13213 (N_13213,N_13042,N_12951);
xor U13214 (N_13214,N_13029,N_13197);
nor U13215 (N_13215,N_12950,N_13159);
xnor U13216 (N_13216,N_13154,N_12909);
xor U13217 (N_13217,N_13118,N_13059);
or U13218 (N_13218,N_13001,N_12966);
nor U13219 (N_13219,N_13141,N_13086);
xnor U13220 (N_13220,N_13016,N_13140);
nand U13221 (N_13221,N_13173,N_13121);
and U13222 (N_13222,N_13037,N_12983);
and U13223 (N_13223,N_13062,N_13027);
and U13224 (N_13224,N_12994,N_12944);
xor U13225 (N_13225,N_12962,N_12975);
or U13226 (N_13226,N_12997,N_13080);
or U13227 (N_13227,N_12964,N_12921);
nand U13228 (N_13228,N_13126,N_13138);
nor U13229 (N_13229,N_12948,N_13097);
nand U13230 (N_13230,N_13066,N_13047);
xnor U13231 (N_13231,N_13088,N_13168);
xnor U13232 (N_13232,N_12984,N_13177);
nand U13233 (N_13233,N_12965,N_13050);
or U13234 (N_13234,N_13114,N_12923);
nor U13235 (N_13235,N_12902,N_13092);
and U13236 (N_13236,N_13072,N_13033);
and U13237 (N_13237,N_13148,N_12949);
nor U13238 (N_13238,N_12989,N_13190);
or U13239 (N_13239,N_13083,N_12912);
or U13240 (N_13240,N_12985,N_13153);
xor U13241 (N_13241,N_13052,N_13158);
or U13242 (N_13242,N_13195,N_12954);
nor U13243 (N_13243,N_12932,N_12968);
nor U13244 (N_13244,N_12917,N_13196);
xnor U13245 (N_13245,N_13049,N_13093);
and U13246 (N_13246,N_12907,N_13164);
xor U13247 (N_13247,N_13100,N_12979);
or U13248 (N_13248,N_13078,N_13020);
nand U13249 (N_13249,N_13103,N_12918);
and U13250 (N_13250,N_12910,N_13014);
nand U13251 (N_13251,N_13030,N_12999);
and U13252 (N_13252,N_13143,N_13105);
xor U13253 (N_13253,N_13176,N_13095);
nor U13254 (N_13254,N_12936,N_12972);
xnor U13255 (N_13255,N_12969,N_13139);
and U13256 (N_13256,N_13026,N_12940);
xnor U13257 (N_13257,N_13003,N_13112);
nor U13258 (N_13258,N_13188,N_13119);
nand U13259 (N_13259,N_13104,N_12952);
and U13260 (N_13260,N_13189,N_13018);
xor U13261 (N_13261,N_13110,N_13161);
xor U13262 (N_13262,N_12914,N_13094);
and U13263 (N_13263,N_12956,N_13034);
and U13264 (N_13264,N_13021,N_12938);
or U13265 (N_13265,N_12926,N_13186);
nand U13266 (N_13266,N_12947,N_13101);
nor U13267 (N_13267,N_13022,N_13151);
and U13268 (N_13268,N_12925,N_13193);
or U13269 (N_13269,N_13165,N_12941);
nor U13270 (N_13270,N_12990,N_12911);
or U13271 (N_13271,N_12992,N_13184);
nor U13272 (N_13272,N_13124,N_13053);
or U13273 (N_13273,N_13129,N_13007);
and U13274 (N_13274,N_12945,N_12996);
or U13275 (N_13275,N_13170,N_13045);
and U13276 (N_13276,N_13089,N_13043);
xor U13277 (N_13277,N_13180,N_13039);
nor U13278 (N_13278,N_13133,N_12981);
and U13279 (N_13279,N_13136,N_13123);
nand U13280 (N_13280,N_13064,N_13025);
and U13281 (N_13281,N_13000,N_13051);
xnor U13282 (N_13282,N_12937,N_13090);
nor U13283 (N_13283,N_12908,N_12905);
nand U13284 (N_13284,N_12943,N_13061);
nand U13285 (N_13285,N_12963,N_13067);
xnor U13286 (N_13286,N_13036,N_13005);
nor U13287 (N_13287,N_13108,N_12959);
or U13288 (N_13288,N_13107,N_13035);
nand U13289 (N_13289,N_12971,N_13031);
xnor U13290 (N_13290,N_13073,N_13135);
or U13291 (N_13291,N_13147,N_12935);
nor U13292 (N_13292,N_13019,N_13152);
or U13293 (N_13293,N_12900,N_12903);
or U13294 (N_13294,N_13167,N_13023);
or U13295 (N_13295,N_13081,N_13185);
nor U13296 (N_13296,N_12993,N_12939);
and U13297 (N_13297,N_13040,N_13187);
or U13298 (N_13298,N_12957,N_13032);
or U13299 (N_13299,N_13117,N_13011);
and U13300 (N_13300,N_13198,N_13017);
and U13301 (N_13301,N_12901,N_12928);
and U13302 (N_13302,N_12913,N_13113);
and U13303 (N_13303,N_12961,N_13010);
xnor U13304 (N_13304,N_13065,N_13063);
and U13305 (N_13305,N_12970,N_13178);
nor U13306 (N_13306,N_13102,N_13074);
xnor U13307 (N_13307,N_13163,N_13015);
nor U13308 (N_13308,N_13076,N_13004);
xor U13309 (N_13309,N_13087,N_13069);
or U13310 (N_13310,N_12934,N_13120);
nor U13311 (N_13311,N_13142,N_12977);
or U13312 (N_13312,N_13084,N_13182);
nand U13313 (N_13313,N_12922,N_12946);
and U13314 (N_13314,N_13134,N_13191);
nand U13315 (N_13315,N_13070,N_13048);
or U13316 (N_13316,N_13172,N_13183);
nor U13317 (N_13317,N_12953,N_13131);
nor U13318 (N_13318,N_13055,N_12976);
nand U13319 (N_13319,N_13098,N_12958);
or U13320 (N_13320,N_13028,N_13071);
or U13321 (N_13321,N_13054,N_13192);
nor U13322 (N_13322,N_13128,N_12978);
and U13323 (N_13323,N_12927,N_12995);
and U13324 (N_13324,N_12991,N_13085);
nor U13325 (N_13325,N_13041,N_13155);
or U13326 (N_13326,N_13179,N_12988);
and U13327 (N_13327,N_12998,N_12973);
or U13328 (N_13328,N_13130,N_12904);
xnor U13329 (N_13329,N_13079,N_12986);
xor U13330 (N_13330,N_13056,N_13091);
and U13331 (N_13331,N_13171,N_12982);
xor U13332 (N_13332,N_13111,N_13099);
xor U13333 (N_13333,N_12930,N_13002);
nand U13334 (N_13334,N_13082,N_13181);
nor U13335 (N_13335,N_13146,N_12915);
xor U13336 (N_13336,N_13077,N_13009);
xnor U13337 (N_13337,N_12980,N_12942);
nor U13338 (N_13338,N_13169,N_13060);
xor U13339 (N_13339,N_13157,N_13012);
nand U13340 (N_13340,N_12919,N_12920);
xor U13341 (N_13341,N_12987,N_13137);
nor U13342 (N_13342,N_12929,N_13008);
or U13343 (N_13343,N_13144,N_13044);
nor U13344 (N_13344,N_13096,N_12931);
or U13345 (N_13345,N_12955,N_13109);
nand U13346 (N_13346,N_13006,N_12924);
nand U13347 (N_13347,N_13013,N_13122);
nand U13348 (N_13348,N_13145,N_12960);
nand U13349 (N_13349,N_13068,N_13199);
or U13350 (N_13350,N_13186,N_12973);
or U13351 (N_13351,N_12988,N_13012);
nor U13352 (N_13352,N_12947,N_13151);
xor U13353 (N_13353,N_13002,N_13173);
xnor U13354 (N_13354,N_12986,N_12950);
and U13355 (N_13355,N_13029,N_12964);
or U13356 (N_13356,N_12914,N_13080);
and U13357 (N_13357,N_13022,N_13081);
xor U13358 (N_13358,N_12922,N_13199);
nand U13359 (N_13359,N_13176,N_13124);
or U13360 (N_13360,N_13065,N_13094);
nor U13361 (N_13361,N_13023,N_13034);
or U13362 (N_13362,N_12953,N_13129);
nand U13363 (N_13363,N_12973,N_12978);
or U13364 (N_13364,N_12981,N_13165);
nor U13365 (N_13365,N_12973,N_13018);
xnor U13366 (N_13366,N_12976,N_13132);
and U13367 (N_13367,N_13085,N_13164);
and U13368 (N_13368,N_13140,N_13042);
or U13369 (N_13369,N_13157,N_13149);
nor U13370 (N_13370,N_13177,N_13033);
xor U13371 (N_13371,N_13197,N_13033);
nor U13372 (N_13372,N_13026,N_12944);
nand U13373 (N_13373,N_12969,N_13016);
or U13374 (N_13374,N_12955,N_13013);
nor U13375 (N_13375,N_12947,N_13188);
nand U13376 (N_13376,N_13131,N_13007);
nor U13377 (N_13377,N_13047,N_12910);
or U13378 (N_13378,N_12949,N_13078);
nand U13379 (N_13379,N_13032,N_13145);
or U13380 (N_13380,N_13153,N_12937);
nand U13381 (N_13381,N_12922,N_13118);
nand U13382 (N_13382,N_13035,N_12953);
xnor U13383 (N_13383,N_12926,N_13073);
xor U13384 (N_13384,N_13096,N_13136);
nand U13385 (N_13385,N_13122,N_13033);
nand U13386 (N_13386,N_13110,N_13113);
nand U13387 (N_13387,N_13047,N_13137);
nor U13388 (N_13388,N_13070,N_12989);
xnor U13389 (N_13389,N_13170,N_12968);
or U13390 (N_13390,N_12912,N_13188);
or U13391 (N_13391,N_12927,N_13158);
or U13392 (N_13392,N_13109,N_13042);
nor U13393 (N_13393,N_12923,N_13090);
and U13394 (N_13394,N_13177,N_12904);
xor U13395 (N_13395,N_13019,N_13080);
and U13396 (N_13396,N_12952,N_12990);
and U13397 (N_13397,N_13030,N_13122);
and U13398 (N_13398,N_12960,N_13061);
or U13399 (N_13399,N_12941,N_13036);
nand U13400 (N_13400,N_13098,N_12960);
nand U13401 (N_13401,N_13147,N_13083);
or U13402 (N_13402,N_13051,N_12938);
nand U13403 (N_13403,N_12959,N_13175);
or U13404 (N_13404,N_13064,N_13083);
or U13405 (N_13405,N_12946,N_13028);
nor U13406 (N_13406,N_13121,N_12990);
xor U13407 (N_13407,N_13146,N_12912);
xnor U13408 (N_13408,N_13010,N_13137);
nor U13409 (N_13409,N_13139,N_13018);
and U13410 (N_13410,N_13160,N_13096);
nand U13411 (N_13411,N_13069,N_13126);
nor U13412 (N_13412,N_12915,N_13091);
and U13413 (N_13413,N_13196,N_13071);
and U13414 (N_13414,N_13154,N_13161);
or U13415 (N_13415,N_12997,N_12958);
and U13416 (N_13416,N_13021,N_13058);
or U13417 (N_13417,N_12973,N_13036);
xnor U13418 (N_13418,N_12974,N_13139);
and U13419 (N_13419,N_13007,N_13066);
xnor U13420 (N_13420,N_13171,N_12951);
or U13421 (N_13421,N_13068,N_13153);
nand U13422 (N_13422,N_13048,N_12928);
xnor U13423 (N_13423,N_13081,N_12909);
or U13424 (N_13424,N_13061,N_13175);
xnor U13425 (N_13425,N_13000,N_13025);
nand U13426 (N_13426,N_12948,N_13067);
xnor U13427 (N_13427,N_13059,N_13173);
xnor U13428 (N_13428,N_13019,N_13168);
nand U13429 (N_13429,N_13003,N_13180);
or U13430 (N_13430,N_13030,N_12916);
or U13431 (N_13431,N_13085,N_13100);
or U13432 (N_13432,N_13062,N_12987);
nor U13433 (N_13433,N_13024,N_13161);
nand U13434 (N_13434,N_13039,N_13041);
and U13435 (N_13435,N_13010,N_13176);
xor U13436 (N_13436,N_13021,N_12977);
and U13437 (N_13437,N_13021,N_12972);
or U13438 (N_13438,N_13074,N_13075);
nand U13439 (N_13439,N_13054,N_13188);
nand U13440 (N_13440,N_13085,N_13035);
xor U13441 (N_13441,N_13110,N_13134);
nand U13442 (N_13442,N_13147,N_13048);
or U13443 (N_13443,N_13004,N_12944);
nand U13444 (N_13444,N_13001,N_12995);
xor U13445 (N_13445,N_13037,N_12942);
xor U13446 (N_13446,N_12934,N_13195);
nor U13447 (N_13447,N_13108,N_13129);
nor U13448 (N_13448,N_13015,N_13065);
nor U13449 (N_13449,N_12995,N_12948);
nor U13450 (N_13450,N_13146,N_13119);
and U13451 (N_13451,N_13124,N_13033);
xor U13452 (N_13452,N_13121,N_13034);
nand U13453 (N_13453,N_12979,N_13006);
xor U13454 (N_13454,N_12914,N_13058);
and U13455 (N_13455,N_13161,N_12936);
and U13456 (N_13456,N_13051,N_13080);
and U13457 (N_13457,N_12952,N_13093);
nand U13458 (N_13458,N_13169,N_12950);
or U13459 (N_13459,N_13040,N_12917);
xnor U13460 (N_13460,N_13199,N_12978);
xnor U13461 (N_13461,N_13139,N_12967);
or U13462 (N_13462,N_12986,N_12955);
or U13463 (N_13463,N_13193,N_12985);
nor U13464 (N_13464,N_12930,N_13140);
nand U13465 (N_13465,N_12975,N_13136);
nand U13466 (N_13466,N_13043,N_12991);
nand U13467 (N_13467,N_13108,N_13000);
and U13468 (N_13468,N_13082,N_13157);
xnor U13469 (N_13469,N_13172,N_13169);
nand U13470 (N_13470,N_12937,N_12982);
nand U13471 (N_13471,N_13038,N_12945);
nand U13472 (N_13472,N_13171,N_13110);
xnor U13473 (N_13473,N_12987,N_13049);
or U13474 (N_13474,N_12996,N_12960);
xnor U13475 (N_13475,N_12933,N_12939);
nor U13476 (N_13476,N_13181,N_13144);
or U13477 (N_13477,N_13012,N_13003);
and U13478 (N_13478,N_12998,N_12983);
nand U13479 (N_13479,N_12965,N_13103);
nor U13480 (N_13480,N_12944,N_13162);
and U13481 (N_13481,N_12949,N_13177);
xnor U13482 (N_13482,N_12923,N_12970);
nand U13483 (N_13483,N_12917,N_13111);
and U13484 (N_13484,N_13132,N_13072);
or U13485 (N_13485,N_13175,N_13180);
nand U13486 (N_13486,N_12983,N_13009);
nand U13487 (N_13487,N_13126,N_13028);
xnor U13488 (N_13488,N_13091,N_12950);
nor U13489 (N_13489,N_12960,N_13189);
nor U13490 (N_13490,N_13079,N_13078);
or U13491 (N_13491,N_12992,N_12994);
xnor U13492 (N_13492,N_13132,N_12910);
nor U13493 (N_13493,N_12985,N_13199);
nor U13494 (N_13494,N_13032,N_13042);
or U13495 (N_13495,N_13188,N_13163);
and U13496 (N_13496,N_13173,N_13176);
nand U13497 (N_13497,N_12986,N_13102);
and U13498 (N_13498,N_12930,N_13019);
and U13499 (N_13499,N_13045,N_13192);
nor U13500 (N_13500,N_13380,N_13322);
nor U13501 (N_13501,N_13242,N_13454);
nor U13502 (N_13502,N_13406,N_13271);
and U13503 (N_13503,N_13277,N_13264);
nor U13504 (N_13504,N_13486,N_13300);
nand U13505 (N_13505,N_13378,N_13289);
xnor U13506 (N_13506,N_13328,N_13464);
nor U13507 (N_13507,N_13362,N_13267);
nor U13508 (N_13508,N_13266,N_13246);
nor U13509 (N_13509,N_13471,N_13317);
nor U13510 (N_13510,N_13210,N_13403);
or U13511 (N_13511,N_13333,N_13435);
and U13512 (N_13512,N_13469,N_13290);
xor U13513 (N_13513,N_13462,N_13459);
and U13514 (N_13514,N_13433,N_13438);
nand U13515 (N_13515,N_13262,N_13395);
nand U13516 (N_13516,N_13237,N_13306);
or U13517 (N_13517,N_13226,N_13444);
and U13518 (N_13518,N_13234,N_13215);
or U13519 (N_13519,N_13304,N_13346);
and U13520 (N_13520,N_13302,N_13407);
nand U13521 (N_13521,N_13429,N_13483);
xnor U13522 (N_13522,N_13252,N_13309);
nand U13523 (N_13523,N_13364,N_13453);
xnor U13524 (N_13524,N_13335,N_13439);
nor U13525 (N_13525,N_13451,N_13205);
nand U13526 (N_13526,N_13381,N_13200);
and U13527 (N_13527,N_13458,N_13342);
xor U13528 (N_13528,N_13278,N_13313);
and U13529 (N_13529,N_13389,N_13321);
or U13530 (N_13530,N_13343,N_13474);
or U13531 (N_13531,N_13225,N_13355);
or U13532 (N_13532,N_13390,N_13298);
nor U13533 (N_13533,N_13365,N_13287);
nand U13534 (N_13534,N_13258,N_13347);
nor U13535 (N_13535,N_13385,N_13201);
xor U13536 (N_13536,N_13376,N_13467);
nor U13537 (N_13537,N_13479,N_13330);
xnor U13538 (N_13538,N_13257,N_13497);
xnor U13539 (N_13539,N_13478,N_13404);
nor U13540 (N_13540,N_13254,N_13485);
and U13541 (N_13541,N_13269,N_13452);
xnor U13542 (N_13542,N_13299,N_13415);
xnor U13543 (N_13543,N_13447,N_13220);
nand U13544 (N_13544,N_13379,N_13473);
nand U13545 (N_13545,N_13297,N_13394);
or U13546 (N_13546,N_13293,N_13224);
nor U13547 (N_13547,N_13386,N_13239);
xnor U13548 (N_13548,N_13426,N_13425);
xor U13549 (N_13549,N_13440,N_13268);
nor U13550 (N_13550,N_13291,N_13377);
nor U13551 (N_13551,N_13323,N_13339);
nor U13552 (N_13552,N_13375,N_13270);
xnor U13553 (N_13553,N_13236,N_13247);
and U13554 (N_13554,N_13431,N_13296);
nor U13555 (N_13555,N_13372,N_13332);
or U13556 (N_13556,N_13392,N_13230);
nand U13557 (N_13557,N_13314,N_13401);
nand U13558 (N_13558,N_13273,N_13318);
xnor U13559 (N_13559,N_13228,N_13427);
and U13560 (N_13560,N_13441,N_13256);
xor U13561 (N_13561,N_13382,N_13432);
nor U13562 (N_13562,N_13341,N_13495);
or U13563 (N_13563,N_13371,N_13437);
or U13564 (N_13564,N_13261,N_13461);
nand U13565 (N_13565,N_13494,N_13295);
nor U13566 (N_13566,N_13259,N_13449);
xnor U13567 (N_13567,N_13421,N_13217);
nor U13568 (N_13568,N_13481,N_13319);
nand U13569 (N_13569,N_13216,N_13249);
or U13570 (N_13570,N_13282,N_13465);
nand U13571 (N_13571,N_13410,N_13397);
xor U13572 (N_13572,N_13211,N_13482);
nor U13573 (N_13573,N_13233,N_13285);
nor U13574 (N_13574,N_13312,N_13276);
and U13575 (N_13575,N_13344,N_13260);
nor U13576 (N_13576,N_13475,N_13284);
nand U13577 (N_13577,N_13345,N_13214);
or U13578 (N_13578,N_13489,N_13402);
and U13579 (N_13579,N_13491,N_13253);
or U13580 (N_13580,N_13241,N_13434);
nand U13581 (N_13581,N_13206,N_13393);
xnor U13582 (N_13582,N_13367,N_13411);
and U13583 (N_13583,N_13487,N_13340);
xor U13584 (N_13584,N_13316,N_13466);
nor U13585 (N_13585,N_13408,N_13400);
nor U13586 (N_13586,N_13263,N_13373);
nor U13587 (N_13587,N_13456,N_13251);
xor U13588 (N_13588,N_13281,N_13272);
and U13589 (N_13589,N_13472,N_13476);
nand U13590 (N_13590,N_13255,N_13357);
nor U13591 (N_13591,N_13436,N_13325);
and U13592 (N_13592,N_13280,N_13238);
nand U13593 (N_13593,N_13274,N_13351);
nor U13594 (N_13594,N_13303,N_13480);
nand U13595 (N_13595,N_13396,N_13336);
nor U13596 (N_13596,N_13409,N_13391);
xor U13597 (N_13597,N_13331,N_13457);
and U13598 (N_13598,N_13398,N_13349);
or U13599 (N_13599,N_13450,N_13209);
and U13600 (N_13600,N_13477,N_13283);
xor U13601 (N_13601,N_13227,N_13202);
xor U13602 (N_13602,N_13366,N_13231);
and U13603 (N_13603,N_13310,N_13498);
or U13604 (N_13604,N_13219,N_13419);
or U13605 (N_13605,N_13488,N_13213);
and U13606 (N_13606,N_13455,N_13221);
or U13607 (N_13607,N_13265,N_13353);
or U13608 (N_13608,N_13207,N_13212);
nand U13609 (N_13609,N_13245,N_13423);
or U13610 (N_13610,N_13356,N_13240);
xor U13611 (N_13611,N_13416,N_13279);
nor U13612 (N_13612,N_13414,N_13223);
nor U13613 (N_13613,N_13496,N_13368);
nor U13614 (N_13614,N_13460,N_13484);
nor U13615 (N_13615,N_13204,N_13326);
nand U13616 (N_13616,N_13417,N_13354);
and U13617 (N_13617,N_13442,N_13232);
xor U13618 (N_13618,N_13413,N_13288);
and U13619 (N_13619,N_13374,N_13405);
xor U13620 (N_13620,N_13387,N_13352);
and U13621 (N_13621,N_13350,N_13470);
xor U13622 (N_13622,N_13203,N_13235);
and U13623 (N_13623,N_13301,N_13338);
or U13624 (N_13624,N_13218,N_13412);
and U13625 (N_13625,N_13250,N_13430);
or U13626 (N_13626,N_13320,N_13334);
and U13627 (N_13627,N_13337,N_13358);
or U13628 (N_13628,N_13286,N_13244);
xnor U13629 (N_13629,N_13248,N_13308);
nand U13630 (N_13630,N_13305,N_13383);
and U13631 (N_13631,N_13388,N_13490);
xor U13632 (N_13632,N_13492,N_13363);
or U13633 (N_13633,N_13307,N_13292);
and U13634 (N_13634,N_13222,N_13443);
or U13635 (N_13635,N_13208,N_13445);
and U13636 (N_13636,N_13315,N_13243);
and U13637 (N_13637,N_13348,N_13384);
xor U13638 (N_13638,N_13360,N_13329);
nand U13639 (N_13639,N_13294,N_13446);
nor U13640 (N_13640,N_13369,N_13428);
or U13641 (N_13641,N_13370,N_13399);
and U13642 (N_13642,N_13311,N_13327);
nor U13643 (N_13643,N_13463,N_13424);
xnor U13644 (N_13644,N_13422,N_13324);
nand U13645 (N_13645,N_13420,N_13448);
and U13646 (N_13646,N_13493,N_13361);
xnor U13647 (N_13647,N_13468,N_13359);
nor U13648 (N_13648,N_13499,N_13229);
xor U13649 (N_13649,N_13275,N_13418);
nor U13650 (N_13650,N_13425,N_13448);
nand U13651 (N_13651,N_13237,N_13342);
and U13652 (N_13652,N_13238,N_13460);
xnor U13653 (N_13653,N_13261,N_13454);
xnor U13654 (N_13654,N_13460,N_13470);
nand U13655 (N_13655,N_13298,N_13362);
xnor U13656 (N_13656,N_13390,N_13380);
or U13657 (N_13657,N_13421,N_13359);
nand U13658 (N_13658,N_13253,N_13417);
nand U13659 (N_13659,N_13251,N_13227);
nand U13660 (N_13660,N_13299,N_13345);
or U13661 (N_13661,N_13268,N_13472);
nor U13662 (N_13662,N_13433,N_13418);
nand U13663 (N_13663,N_13202,N_13464);
nand U13664 (N_13664,N_13443,N_13269);
xnor U13665 (N_13665,N_13456,N_13281);
or U13666 (N_13666,N_13438,N_13452);
nor U13667 (N_13667,N_13242,N_13248);
nand U13668 (N_13668,N_13456,N_13288);
nand U13669 (N_13669,N_13466,N_13457);
nor U13670 (N_13670,N_13406,N_13353);
nor U13671 (N_13671,N_13316,N_13465);
nor U13672 (N_13672,N_13216,N_13461);
or U13673 (N_13673,N_13398,N_13480);
nand U13674 (N_13674,N_13278,N_13488);
xnor U13675 (N_13675,N_13308,N_13271);
nand U13676 (N_13676,N_13254,N_13471);
or U13677 (N_13677,N_13379,N_13362);
nor U13678 (N_13678,N_13412,N_13305);
or U13679 (N_13679,N_13352,N_13349);
nand U13680 (N_13680,N_13200,N_13219);
xor U13681 (N_13681,N_13381,N_13303);
nand U13682 (N_13682,N_13274,N_13347);
xor U13683 (N_13683,N_13281,N_13469);
xor U13684 (N_13684,N_13484,N_13278);
or U13685 (N_13685,N_13321,N_13417);
nand U13686 (N_13686,N_13448,N_13309);
or U13687 (N_13687,N_13336,N_13232);
xnor U13688 (N_13688,N_13222,N_13314);
nand U13689 (N_13689,N_13386,N_13265);
and U13690 (N_13690,N_13440,N_13231);
nor U13691 (N_13691,N_13405,N_13496);
xnor U13692 (N_13692,N_13393,N_13447);
nand U13693 (N_13693,N_13438,N_13216);
nor U13694 (N_13694,N_13453,N_13404);
nor U13695 (N_13695,N_13302,N_13256);
nand U13696 (N_13696,N_13208,N_13361);
or U13697 (N_13697,N_13289,N_13228);
xnor U13698 (N_13698,N_13355,N_13409);
nand U13699 (N_13699,N_13363,N_13340);
nor U13700 (N_13700,N_13300,N_13451);
or U13701 (N_13701,N_13327,N_13369);
and U13702 (N_13702,N_13435,N_13363);
nand U13703 (N_13703,N_13488,N_13322);
nor U13704 (N_13704,N_13324,N_13300);
and U13705 (N_13705,N_13430,N_13324);
and U13706 (N_13706,N_13351,N_13421);
or U13707 (N_13707,N_13418,N_13216);
or U13708 (N_13708,N_13464,N_13432);
or U13709 (N_13709,N_13368,N_13318);
nor U13710 (N_13710,N_13402,N_13271);
xor U13711 (N_13711,N_13494,N_13379);
nor U13712 (N_13712,N_13399,N_13368);
nand U13713 (N_13713,N_13467,N_13469);
xnor U13714 (N_13714,N_13229,N_13330);
nand U13715 (N_13715,N_13268,N_13477);
nand U13716 (N_13716,N_13474,N_13331);
and U13717 (N_13717,N_13296,N_13390);
or U13718 (N_13718,N_13437,N_13460);
nand U13719 (N_13719,N_13247,N_13414);
nor U13720 (N_13720,N_13265,N_13465);
or U13721 (N_13721,N_13223,N_13432);
xor U13722 (N_13722,N_13290,N_13216);
nor U13723 (N_13723,N_13398,N_13408);
and U13724 (N_13724,N_13452,N_13398);
or U13725 (N_13725,N_13260,N_13372);
and U13726 (N_13726,N_13272,N_13321);
or U13727 (N_13727,N_13372,N_13343);
and U13728 (N_13728,N_13316,N_13234);
nor U13729 (N_13729,N_13471,N_13470);
nor U13730 (N_13730,N_13287,N_13385);
nand U13731 (N_13731,N_13202,N_13255);
xor U13732 (N_13732,N_13259,N_13485);
nor U13733 (N_13733,N_13238,N_13413);
nor U13734 (N_13734,N_13339,N_13249);
and U13735 (N_13735,N_13470,N_13238);
xnor U13736 (N_13736,N_13430,N_13228);
or U13737 (N_13737,N_13465,N_13329);
xor U13738 (N_13738,N_13412,N_13235);
nor U13739 (N_13739,N_13484,N_13330);
nor U13740 (N_13740,N_13220,N_13352);
xor U13741 (N_13741,N_13460,N_13397);
or U13742 (N_13742,N_13421,N_13284);
nor U13743 (N_13743,N_13294,N_13292);
nor U13744 (N_13744,N_13478,N_13451);
nor U13745 (N_13745,N_13326,N_13478);
or U13746 (N_13746,N_13275,N_13491);
xor U13747 (N_13747,N_13287,N_13463);
nor U13748 (N_13748,N_13262,N_13276);
nor U13749 (N_13749,N_13333,N_13330);
and U13750 (N_13750,N_13243,N_13332);
xnor U13751 (N_13751,N_13402,N_13387);
nand U13752 (N_13752,N_13202,N_13285);
and U13753 (N_13753,N_13243,N_13394);
xor U13754 (N_13754,N_13343,N_13266);
xor U13755 (N_13755,N_13435,N_13403);
nor U13756 (N_13756,N_13279,N_13373);
or U13757 (N_13757,N_13343,N_13254);
xor U13758 (N_13758,N_13484,N_13458);
xnor U13759 (N_13759,N_13486,N_13258);
nor U13760 (N_13760,N_13476,N_13396);
xnor U13761 (N_13761,N_13430,N_13258);
nand U13762 (N_13762,N_13384,N_13437);
xor U13763 (N_13763,N_13477,N_13417);
nand U13764 (N_13764,N_13414,N_13319);
nand U13765 (N_13765,N_13347,N_13282);
and U13766 (N_13766,N_13345,N_13473);
xor U13767 (N_13767,N_13467,N_13371);
xnor U13768 (N_13768,N_13410,N_13236);
and U13769 (N_13769,N_13325,N_13474);
nor U13770 (N_13770,N_13399,N_13392);
xnor U13771 (N_13771,N_13426,N_13324);
or U13772 (N_13772,N_13296,N_13486);
nand U13773 (N_13773,N_13313,N_13324);
or U13774 (N_13774,N_13498,N_13241);
and U13775 (N_13775,N_13274,N_13492);
nand U13776 (N_13776,N_13475,N_13430);
nor U13777 (N_13777,N_13341,N_13417);
and U13778 (N_13778,N_13271,N_13472);
nor U13779 (N_13779,N_13280,N_13363);
xnor U13780 (N_13780,N_13423,N_13457);
nor U13781 (N_13781,N_13461,N_13353);
or U13782 (N_13782,N_13400,N_13417);
nand U13783 (N_13783,N_13487,N_13455);
or U13784 (N_13784,N_13392,N_13450);
nand U13785 (N_13785,N_13425,N_13258);
or U13786 (N_13786,N_13316,N_13264);
nor U13787 (N_13787,N_13244,N_13377);
nor U13788 (N_13788,N_13372,N_13218);
nand U13789 (N_13789,N_13388,N_13207);
or U13790 (N_13790,N_13201,N_13299);
and U13791 (N_13791,N_13259,N_13462);
and U13792 (N_13792,N_13330,N_13417);
nor U13793 (N_13793,N_13387,N_13312);
and U13794 (N_13794,N_13398,N_13224);
xnor U13795 (N_13795,N_13307,N_13265);
or U13796 (N_13796,N_13412,N_13433);
nor U13797 (N_13797,N_13436,N_13301);
nor U13798 (N_13798,N_13423,N_13393);
nand U13799 (N_13799,N_13252,N_13373);
nor U13800 (N_13800,N_13693,N_13573);
nor U13801 (N_13801,N_13722,N_13561);
nand U13802 (N_13802,N_13636,N_13565);
nand U13803 (N_13803,N_13773,N_13676);
or U13804 (N_13804,N_13723,N_13580);
xnor U13805 (N_13805,N_13519,N_13584);
nand U13806 (N_13806,N_13560,N_13550);
xnor U13807 (N_13807,N_13675,N_13583);
or U13808 (N_13808,N_13623,N_13517);
xor U13809 (N_13809,N_13787,N_13671);
nor U13810 (N_13810,N_13670,N_13632);
and U13811 (N_13811,N_13566,N_13709);
nor U13812 (N_13812,N_13653,N_13741);
nor U13813 (N_13813,N_13521,N_13512);
nor U13814 (N_13814,N_13790,N_13549);
and U13815 (N_13815,N_13527,N_13554);
or U13816 (N_13816,N_13640,N_13626);
nor U13817 (N_13817,N_13620,N_13768);
xnor U13818 (N_13818,N_13513,N_13673);
and U13819 (N_13819,N_13766,N_13639);
or U13820 (N_13820,N_13799,N_13765);
xor U13821 (N_13821,N_13572,N_13694);
nor U13822 (N_13822,N_13501,N_13736);
nand U13823 (N_13823,N_13665,N_13792);
nor U13824 (N_13824,N_13578,N_13570);
or U13825 (N_13825,N_13717,N_13514);
and U13826 (N_13826,N_13551,N_13544);
nor U13827 (N_13827,N_13699,N_13760);
nor U13828 (N_13828,N_13726,N_13508);
nand U13829 (N_13829,N_13780,N_13732);
and U13830 (N_13830,N_13615,N_13633);
or U13831 (N_13831,N_13656,N_13602);
nand U13832 (N_13832,N_13581,N_13710);
or U13833 (N_13833,N_13651,N_13716);
or U13834 (N_13834,N_13770,N_13646);
and U13835 (N_13835,N_13610,N_13534);
xor U13836 (N_13836,N_13753,N_13711);
nor U13837 (N_13837,N_13727,N_13531);
and U13838 (N_13838,N_13569,N_13721);
or U13839 (N_13839,N_13645,N_13685);
xor U13840 (N_13840,N_13637,N_13571);
nor U13841 (N_13841,N_13702,N_13795);
nand U13842 (N_13842,N_13526,N_13631);
or U13843 (N_13843,N_13611,N_13720);
xor U13844 (N_13844,N_13729,N_13731);
nand U13845 (N_13845,N_13597,N_13648);
nand U13846 (N_13846,N_13662,N_13627);
nor U13847 (N_13847,N_13754,N_13593);
nor U13848 (N_13848,N_13713,N_13666);
xor U13849 (N_13849,N_13771,N_13558);
and U13850 (N_13850,N_13506,N_13746);
and U13851 (N_13851,N_13567,N_13748);
nor U13852 (N_13852,N_13655,N_13781);
nor U13853 (N_13853,N_13797,N_13784);
or U13854 (N_13854,N_13756,N_13618);
nand U13855 (N_13855,N_13705,N_13577);
nor U13856 (N_13856,N_13616,N_13661);
xor U13857 (N_13857,N_13734,N_13778);
and U13858 (N_13858,N_13791,N_13511);
and U13859 (N_13859,N_13603,N_13677);
xor U13860 (N_13860,N_13530,N_13532);
and U13861 (N_13861,N_13755,N_13798);
nand U13862 (N_13862,N_13613,N_13762);
or U13863 (N_13863,N_13547,N_13520);
nand U13864 (N_13864,N_13657,N_13706);
and U13865 (N_13865,N_13647,N_13692);
nor U13866 (N_13866,N_13700,N_13642);
nand U13867 (N_13867,N_13579,N_13604);
and U13868 (N_13868,N_13704,N_13782);
nor U13869 (N_13869,N_13539,N_13529);
nand U13870 (N_13870,N_13769,N_13739);
or U13871 (N_13871,N_13678,N_13759);
nand U13872 (N_13872,N_13767,N_13664);
nor U13873 (N_13873,N_13764,N_13614);
or U13874 (N_13874,N_13674,N_13747);
or U13875 (N_13875,N_13537,N_13546);
or U13876 (N_13876,N_13590,N_13629);
or U13877 (N_13877,N_13591,N_13689);
xor U13878 (N_13878,N_13559,N_13745);
and U13879 (N_13879,N_13742,N_13545);
or U13880 (N_13880,N_13718,N_13644);
nor U13881 (N_13881,N_13543,N_13660);
nand U13882 (N_13882,N_13641,N_13536);
and U13883 (N_13883,N_13687,N_13761);
and U13884 (N_13884,N_13505,N_13680);
and U13885 (N_13885,N_13786,N_13601);
or U13886 (N_13886,N_13749,N_13625);
and U13887 (N_13887,N_13598,N_13617);
or U13888 (N_13888,N_13743,N_13599);
nor U13889 (N_13889,N_13524,N_13703);
or U13890 (N_13890,N_13735,N_13777);
nor U13891 (N_13891,N_13533,N_13542);
xnor U13892 (N_13892,N_13679,N_13562);
or U13893 (N_13893,N_13667,N_13776);
or U13894 (N_13894,N_13563,N_13690);
nand U13895 (N_13895,N_13619,N_13585);
or U13896 (N_13896,N_13523,N_13630);
or U13897 (N_13897,N_13587,N_13503);
and U13898 (N_13898,N_13714,N_13758);
nand U13899 (N_13899,N_13596,N_13793);
nor U13900 (N_13900,N_13775,N_13698);
and U13901 (N_13901,N_13715,N_13740);
xor U13902 (N_13902,N_13606,N_13600);
or U13903 (N_13903,N_13502,N_13672);
nand U13904 (N_13904,N_13555,N_13535);
nand U13905 (N_13905,N_13658,N_13682);
nand U13906 (N_13906,N_13540,N_13719);
nor U13907 (N_13907,N_13634,N_13785);
nand U13908 (N_13908,N_13688,N_13507);
nor U13909 (N_13909,N_13522,N_13643);
xnor U13910 (N_13910,N_13725,N_13744);
nor U13911 (N_13911,N_13635,N_13538);
nand U13912 (N_13912,N_13712,N_13528);
nor U13913 (N_13913,N_13668,N_13652);
and U13914 (N_13914,N_13621,N_13707);
xor U13915 (N_13915,N_13774,N_13504);
xnor U13916 (N_13916,N_13605,N_13763);
nand U13917 (N_13917,N_13592,N_13576);
nor U13918 (N_13918,N_13552,N_13669);
nor U13919 (N_13919,N_13574,N_13575);
nand U13920 (N_13920,N_13696,N_13541);
or U13921 (N_13921,N_13772,N_13654);
xnor U13922 (N_13922,N_13750,N_13564);
and U13923 (N_13923,N_13789,N_13622);
xnor U13924 (N_13924,N_13697,N_13624);
and U13925 (N_13925,N_13701,N_13730);
nor U13926 (N_13926,N_13695,N_13516);
nor U13927 (N_13927,N_13683,N_13738);
nor U13928 (N_13928,N_13628,N_13649);
nand U13929 (N_13929,N_13609,N_13684);
nor U13930 (N_13930,N_13708,N_13548);
nor U13931 (N_13931,N_13796,N_13608);
and U13932 (N_13932,N_13686,N_13659);
xnor U13933 (N_13933,N_13509,N_13500);
xor U13934 (N_13934,N_13751,N_13607);
nor U13935 (N_13935,N_13663,N_13582);
and U13936 (N_13936,N_13525,N_13728);
nor U13937 (N_13937,N_13783,N_13733);
xnor U13938 (N_13938,N_13752,N_13556);
nor U13939 (N_13939,N_13681,N_13757);
and U13940 (N_13940,N_13594,N_13553);
nand U13941 (N_13941,N_13691,N_13612);
nand U13942 (N_13942,N_13737,N_13568);
nor U13943 (N_13943,N_13595,N_13724);
and U13944 (N_13944,N_13638,N_13510);
or U13945 (N_13945,N_13788,N_13588);
and U13946 (N_13946,N_13557,N_13515);
and U13947 (N_13947,N_13650,N_13779);
xnor U13948 (N_13948,N_13589,N_13586);
or U13949 (N_13949,N_13794,N_13518);
xnor U13950 (N_13950,N_13584,N_13743);
xor U13951 (N_13951,N_13639,N_13744);
and U13952 (N_13952,N_13645,N_13562);
or U13953 (N_13953,N_13711,N_13723);
xnor U13954 (N_13954,N_13783,N_13718);
or U13955 (N_13955,N_13755,N_13757);
nand U13956 (N_13956,N_13628,N_13721);
or U13957 (N_13957,N_13535,N_13698);
nor U13958 (N_13958,N_13627,N_13621);
nand U13959 (N_13959,N_13746,N_13533);
or U13960 (N_13960,N_13782,N_13728);
and U13961 (N_13961,N_13594,N_13790);
nand U13962 (N_13962,N_13514,N_13594);
nor U13963 (N_13963,N_13554,N_13783);
or U13964 (N_13964,N_13782,N_13605);
and U13965 (N_13965,N_13708,N_13632);
xor U13966 (N_13966,N_13686,N_13549);
nor U13967 (N_13967,N_13794,N_13521);
nor U13968 (N_13968,N_13578,N_13627);
xnor U13969 (N_13969,N_13510,N_13660);
nor U13970 (N_13970,N_13674,N_13719);
or U13971 (N_13971,N_13688,N_13692);
nor U13972 (N_13972,N_13705,N_13662);
nand U13973 (N_13973,N_13767,N_13717);
and U13974 (N_13974,N_13638,N_13777);
nor U13975 (N_13975,N_13768,N_13541);
or U13976 (N_13976,N_13718,N_13622);
nand U13977 (N_13977,N_13713,N_13557);
and U13978 (N_13978,N_13560,N_13590);
and U13979 (N_13979,N_13568,N_13570);
xor U13980 (N_13980,N_13751,N_13672);
nor U13981 (N_13981,N_13545,N_13537);
and U13982 (N_13982,N_13655,N_13704);
and U13983 (N_13983,N_13501,N_13625);
and U13984 (N_13984,N_13506,N_13518);
xnor U13985 (N_13985,N_13564,N_13539);
or U13986 (N_13986,N_13508,N_13622);
nand U13987 (N_13987,N_13550,N_13754);
nor U13988 (N_13988,N_13778,N_13703);
xnor U13989 (N_13989,N_13673,N_13719);
or U13990 (N_13990,N_13562,N_13686);
nand U13991 (N_13991,N_13708,N_13783);
or U13992 (N_13992,N_13594,N_13724);
nand U13993 (N_13993,N_13618,N_13511);
nor U13994 (N_13994,N_13631,N_13768);
and U13995 (N_13995,N_13751,N_13697);
or U13996 (N_13996,N_13686,N_13772);
and U13997 (N_13997,N_13686,N_13602);
or U13998 (N_13998,N_13666,N_13572);
or U13999 (N_13999,N_13603,N_13763);
nor U14000 (N_14000,N_13500,N_13764);
nor U14001 (N_14001,N_13537,N_13737);
nor U14002 (N_14002,N_13684,N_13642);
xor U14003 (N_14003,N_13723,N_13623);
and U14004 (N_14004,N_13648,N_13608);
or U14005 (N_14005,N_13639,N_13607);
or U14006 (N_14006,N_13574,N_13536);
and U14007 (N_14007,N_13536,N_13664);
or U14008 (N_14008,N_13785,N_13521);
and U14009 (N_14009,N_13673,N_13704);
and U14010 (N_14010,N_13642,N_13588);
xnor U14011 (N_14011,N_13731,N_13678);
nor U14012 (N_14012,N_13610,N_13511);
nor U14013 (N_14013,N_13762,N_13583);
or U14014 (N_14014,N_13539,N_13582);
xor U14015 (N_14015,N_13676,N_13623);
nor U14016 (N_14016,N_13587,N_13527);
nor U14017 (N_14017,N_13623,N_13573);
nor U14018 (N_14018,N_13525,N_13683);
or U14019 (N_14019,N_13618,N_13545);
or U14020 (N_14020,N_13521,N_13571);
nor U14021 (N_14021,N_13579,N_13766);
and U14022 (N_14022,N_13778,N_13787);
or U14023 (N_14023,N_13764,N_13513);
nand U14024 (N_14024,N_13788,N_13718);
nand U14025 (N_14025,N_13723,N_13585);
nor U14026 (N_14026,N_13571,N_13596);
or U14027 (N_14027,N_13636,N_13611);
or U14028 (N_14028,N_13699,N_13661);
nor U14029 (N_14029,N_13618,N_13716);
and U14030 (N_14030,N_13633,N_13515);
nand U14031 (N_14031,N_13682,N_13785);
nand U14032 (N_14032,N_13684,N_13783);
xnor U14033 (N_14033,N_13760,N_13622);
or U14034 (N_14034,N_13790,N_13754);
nand U14035 (N_14035,N_13624,N_13641);
or U14036 (N_14036,N_13654,N_13705);
nor U14037 (N_14037,N_13572,N_13656);
and U14038 (N_14038,N_13544,N_13673);
or U14039 (N_14039,N_13760,N_13675);
nand U14040 (N_14040,N_13673,N_13730);
xnor U14041 (N_14041,N_13689,N_13763);
and U14042 (N_14042,N_13701,N_13583);
nand U14043 (N_14043,N_13514,N_13504);
or U14044 (N_14044,N_13732,N_13665);
and U14045 (N_14045,N_13766,N_13564);
and U14046 (N_14046,N_13786,N_13670);
xor U14047 (N_14047,N_13755,N_13678);
nand U14048 (N_14048,N_13528,N_13722);
nand U14049 (N_14049,N_13531,N_13689);
and U14050 (N_14050,N_13512,N_13736);
and U14051 (N_14051,N_13612,N_13551);
and U14052 (N_14052,N_13774,N_13719);
and U14053 (N_14053,N_13645,N_13657);
or U14054 (N_14054,N_13610,N_13748);
nor U14055 (N_14055,N_13513,N_13794);
nand U14056 (N_14056,N_13707,N_13582);
or U14057 (N_14057,N_13695,N_13712);
nor U14058 (N_14058,N_13716,N_13784);
and U14059 (N_14059,N_13587,N_13706);
or U14060 (N_14060,N_13642,N_13799);
or U14061 (N_14061,N_13584,N_13597);
nand U14062 (N_14062,N_13798,N_13732);
nor U14063 (N_14063,N_13695,N_13551);
nor U14064 (N_14064,N_13759,N_13709);
nand U14065 (N_14065,N_13732,N_13655);
or U14066 (N_14066,N_13707,N_13519);
or U14067 (N_14067,N_13736,N_13789);
xor U14068 (N_14068,N_13540,N_13559);
xnor U14069 (N_14069,N_13620,N_13762);
or U14070 (N_14070,N_13501,N_13758);
and U14071 (N_14071,N_13711,N_13573);
and U14072 (N_14072,N_13596,N_13656);
and U14073 (N_14073,N_13610,N_13744);
nor U14074 (N_14074,N_13610,N_13530);
xnor U14075 (N_14075,N_13738,N_13547);
and U14076 (N_14076,N_13672,N_13713);
nor U14077 (N_14077,N_13754,N_13564);
or U14078 (N_14078,N_13616,N_13698);
and U14079 (N_14079,N_13640,N_13597);
nand U14080 (N_14080,N_13694,N_13727);
nand U14081 (N_14081,N_13715,N_13656);
xor U14082 (N_14082,N_13522,N_13741);
xnor U14083 (N_14083,N_13694,N_13710);
nand U14084 (N_14084,N_13601,N_13596);
nand U14085 (N_14085,N_13674,N_13515);
or U14086 (N_14086,N_13735,N_13771);
and U14087 (N_14087,N_13547,N_13719);
nand U14088 (N_14088,N_13689,N_13789);
nor U14089 (N_14089,N_13698,N_13662);
xnor U14090 (N_14090,N_13555,N_13608);
nor U14091 (N_14091,N_13750,N_13722);
xnor U14092 (N_14092,N_13764,N_13539);
xor U14093 (N_14093,N_13517,N_13622);
xor U14094 (N_14094,N_13673,N_13688);
or U14095 (N_14095,N_13538,N_13602);
or U14096 (N_14096,N_13734,N_13676);
nand U14097 (N_14097,N_13646,N_13699);
nor U14098 (N_14098,N_13574,N_13754);
xnor U14099 (N_14099,N_13776,N_13740);
xnor U14100 (N_14100,N_13978,N_13818);
xnor U14101 (N_14101,N_13969,N_13868);
or U14102 (N_14102,N_14023,N_13949);
nor U14103 (N_14103,N_13959,N_13816);
or U14104 (N_14104,N_14092,N_13827);
and U14105 (N_14105,N_13916,N_13835);
and U14106 (N_14106,N_13992,N_13815);
or U14107 (N_14107,N_14043,N_14055);
nor U14108 (N_14108,N_13880,N_13857);
xnor U14109 (N_14109,N_14014,N_14056);
nand U14110 (N_14110,N_13933,N_13824);
nor U14111 (N_14111,N_13891,N_13802);
nor U14112 (N_14112,N_13850,N_13892);
xnor U14113 (N_14113,N_14018,N_13828);
nand U14114 (N_14114,N_14086,N_13830);
nand U14115 (N_14115,N_13953,N_13973);
xor U14116 (N_14116,N_13847,N_14067);
nor U14117 (N_14117,N_13820,N_13865);
and U14118 (N_14118,N_13908,N_13956);
nor U14119 (N_14119,N_13900,N_13927);
and U14120 (N_14120,N_14080,N_13941);
xnor U14121 (N_14121,N_14006,N_13987);
or U14122 (N_14122,N_14029,N_13814);
nand U14123 (N_14123,N_13998,N_14064);
or U14124 (N_14124,N_14083,N_13926);
xnor U14125 (N_14125,N_14028,N_14052);
nand U14126 (N_14126,N_13906,N_13833);
or U14127 (N_14127,N_13968,N_13960);
or U14128 (N_14128,N_14072,N_13986);
and U14129 (N_14129,N_14033,N_13917);
or U14130 (N_14130,N_14008,N_14085);
or U14131 (N_14131,N_13938,N_14002);
xnor U14132 (N_14132,N_13909,N_13976);
nand U14133 (N_14133,N_13910,N_14045);
or U14134 (N_14134,N_13902,N_13903);
nand U14135 (N_14135,N_13876,N_13871);
nand U14136 (N_14136,N_14032,N_13947);
nor U14137 (N_14137,N_14093,N_14041);
nand U14138 (N_14138,N_14034,N_13836);
nor U14139 (N_14139,N_14057,N_13955);
nor U14140 (N_14140,N_13838,N_13928);
xnor U14141 (N_14141,N_13901,N_13943);
or U14142 (N_14142,N_13980,N_13832);
nand U14143 (N_14143,N_13885,N_14099);
and U14144 (N_14144,N_13993,N_14098);
xor U14145 (N_14145,N_14016,N_14074);
nor U14146 (N_14146,N_14066,N_13844);
or U14147 (N_14147,N_13883,N_13979);
or U14148 (N_14148,N_13849,N_13930);
nor U14149 (N_14149,N_13935,N_13813);
nand U14150 (N_14150,N_13840,N_13826);
or U14151 (N_14151,N_13867,N_13878);
xnor U14152 (N_14152,N_13874,N_13940);
or U14153 (N_14153,N_13817,N_13972);
and U14154 (N_14154,N_13803,N_14001);
or U14155 (N_14155,N_13869,N_14031);
and U14156 (N_14156,N_13983,N_13807);
or U14157 (N_14157,N_14077,N_13897);
xor U14158 (N_14158,N_14065,N_13848);
nor U14159 (N_14159,N_13948,N_13967);
or U14160 (N_14160,N_13913,N_13859);
xor U14161 (N_14161,N_13811,N_13918);
nor U14162 (N_14162,N_13936,N_13825);
nand U14163 (N_14163,N_14069,N_13988);
nand U14164 (N_14164,N_13889,N_13999);
and U14165 (N_14165,N_13864,N_14075);
xor U14166 (N_14166,N_13942,N_13886);
nand U14167 (N_14167,N_14047,N_14042);
and U14168 (N_14168,N_13887,N_14070);
nand U14169 (N_14169,N_13924,N_13881);
xnor U14170 (N_14170,N_13970,N_14020);
nor U14171 (N_14171,N_14089,N_14054);
or U14172 (N_14172,N_14050,N_13995);
nor U14173 (N_14173,N_14012,N_13934);
or U14174 (N_14174,N_13985,N_13895);
nor U14175 (N_14175,N_14021,N_14000);
nand U14176 (N_14176,N_14097,N_13842);
nand U14177 (N_14177,N_13806,N_13861);
and U14178 (N_14178,N_14003,N_14087);
xnor U14179 (N_14179,N_13898,N_13965);
or U14180 (N_14180,N_13921,N_13879);
and U14181 (N_14181,N_14038,N_14022);
and U14182 (N_14182,N_13872,N_13971);
nor U14183 (N_14183,N_13911,N_14060);
nor U14184 (N_14184,N_13801,N_14079);
nand U14185 (N_14185,N_13896,N_13888);
and U14186 (N_14186,N_13915,N_13862);
nor U14187 (N_14187,N_13804,N_13856);
or U14188 (N_14188,N_14046,N_13812);
and U14189 (N_14189,N_13805,N_13984);
xnor U14190 (N_14190,N_13991,N_14090);
and U14191 (N_14191,N_13954,N_13890);
or U14192 (N_14192,N_14013,N_13893);
and U14193 (N_14193,N_14076,N_14082);
or U14194 (N_14194,N_14005,N_13894);
or U14195 (N_14195,N_13843,N_13929);
and U14196 (N_14196,N_13958,N_14051);
or U14197 (N_14197,N_14024,N_13957);
and U14198 (N_14198,N_13860,N_13834);
nand U14199 (N_14199,N_13904,N_14063);
or U14200 (N_14200,N_13907,N_13875);
and U14201 (N_14201,N_14095,N_13990);
and U14202 (N_14202,N_13839,N_13937);
nor U14203 (N_14203,N_14049,N_14053);
nand U14204 (N_14204,N_14068,N_13997);
xor U14205 (N_14205,N_13851,N_13837);
or U14206 (N_14206,N_13873,N_13962);
and U14207 (N_14207,N_13846,N_13899);
nor U14208 (N_14208,N_14011,N_13852);
or U14209 (N_14209,N_14071,N_13950);
xnor U14210 (N_14210,N_13945,N_13981);
or U14211 (N_14211,N_13982,N_13975);
and U14212 (N_14212,N_14081,N_13877);
or U14213 (N_14213,N_13977,N_14009);
nand U14214 (N_14214,N_13994,N_14017);
nand U14215 (N_14215,N_13961,N_14010);
nor U14216 (N_14216,N_13989,N_14004);
nand U14217 (N_14217,N_13810,N_13931);
xor U14218 (N_14218,N_13951,N_13905);
nand U14219 (N_14219,N_14096,N_14094);
nor U14220 (N_14220,N_14039,N_14019);
xnor U14221 (N_14221,N_13963,N_14036);
or U14222 (N_14222,N_13863,N_13841);
xnor U14223 (N_14223,N_14040,N_14015);
xnor U14224 (N_14224,N_13845,N_13870);
nor U14225 (N_14225,N_13966,N_14048);
nor U14226 (N_14226,N_14091,N_13822);
or U14227 (N_14227,N_14037,N_13866);
nor U14228 (N_14228,N_13996,N_13819);
or U14229 (N_14229,N_13912,N_13823);
xor U14230 (N_14230,N_14078,N_13855);
nor U14231 (N_14231,N_13914,N_13854);
nor U14232 (N_14232,N_13952,N_14088);
or U14233 (N_14233,N_13920,N_14027);
or U14234 (N_14234,N_13821,N_14058);
and U14235 (N_14235,N_14026,N_13919);
nand U14236 (N_14236,N_13974,N_14030);
or U14237 (N_14237,N_13831,N_13829);
nor U14238 (N_14238,N_13939,N_14059);
and U14239 (N_14239,N_14061,N_14062);
and U14240 (N_14240,N_14025,N_13925);
nor U14241 (N_14241,N_13964,N_13858);
nor U14242 (N_14242,N_13946,N_13882);
or U14243 (N_14243,N_13932,N_14007);
and U14244 (N_14244,N_13944,N_13809);
and U14245 (N_14245,N_13922,N_14044);
nand U14246 (N_14246,N_14073,N_13800);
or U14247 (N_14247,N_13808,N_14084);
or U14248 (N_14248,N_13853,N_13923);
or U14249 (N_14249,N_13884,N_14035);
xor U14250 (N_14250,N_13843,N_13881);
and U14251 (N_14251,N_13927,N_13840);
and U14252 (N_14252,N_13905,N_13890);
nand U14253 (N_14253,N_13829,N_13808);
nor U14254 (N_14254,N_13859,N_14029);
and U14255 (N_14255,N_14017,N_13991);
nor U14256 (N_14256,N_13946,N_14026);
xor U14257 (N_14257,N_13812,N_14052);
nand U14258 (N_14258,N_14018,N_13809);
and U14259 (N_14259,N_13883,N_13990);
or U14260 (N_14260,N_13994,N_14055);
nor U14261 (N_14261,N_14044,N_13867);
xor U14262 (N_14262,N_13875,N_13883);
or U14263 (N_14263,N_13890,N_14025);
xnor U14264 (N_14264,N_13835,N_13925);
xnor U14265 (N_14265,N_14092,N_13835);
nand U14266 (N_14266,N_13838,N_13872);
nor U14267 (N_14267,N_14067,N_13893);
nor U14268 (N_14268,N_14035,N_13975);
nor U14269 (N_14269,N_13994,N_14083);
xor U14270 (N_14270,N_13829,N_14068);
or U14271 (N_14271,N_14009,N_13813);
and U14272 (N_14272,N_14066,N_14098);
xnor U14273 (N_14273,N_13963,N_13895);
xor U14274 (N_14274,N_13900,N_14083);
nand U14275 (N_14275,N_13850,N_13900);
nand U14276 (N_14276,N_14037,N_13944);
and U14277 (N_14277,N_14096,N_13875);
nor U14278 (N_14278,N_14050,N_13900);
or U14279 (N_14279,N_13919,N_14070);
xor U14280 (N_14280,N_13984,N_14082);
and U14281 (N_14281,N_13851,N_13876);
nor U14282 (N_14282,N_13910,N_13926);
or U14283 (N_14283,N_14096,N_13872);
or U14284 (N_14284,N_14061,N_13898);
xor U14285 (N_14285,N_13927,N_13866);
nor U14286 (N_14286,N_13831,N_14070);
and U14287 (N_14287,N_13811,N_13837);
nand U14288 (N_14288,N_13829,N_13912);
nor U14289 (N_14289,N_14087,N_14047);
and U14290 (N_14290,N_13978,N_13976);
and U14291 (N_14291,N_13992,N_14068);
nand U14292 (N_14292,N_13911,N_14009);
xnor U14293 (N_14293,N_14075,N_13809);
and U14294 (N_14294,N_13887,N_13833);
xor U14295 (N_14295,N_14088,N_13816);
or U14296 (N_14296,N_13987,N_14050);
and U14297 (N_14297,N_13885,N_13800);
nand U14298 (N_14298,N_13927,N_13836);
and U14299 (N_14299,N_14024,N_14069);
or U14300 (N_14300,N_13956,N_13901);
nand U14301 (N_14301,N_14020,N_14023);
nand U14302 (N_14302,N_13889,N_13930);
nand U14303 (N_14303,N_14099,N_14044);
nand U14304 (N_14304,N_13910,N_13907);
nand U14305 (N_14305,N_13963,N_13800);
xnor U14306 (N_14306,N_14032,N_13874);
nand U14307 (N_14307,N_13959,N_13970);
nor U14308 (N_14308,N_13801,N_13923);
and U14309 (N_14309,N_14098,N_13880);
and U14310 (N_14310,N_13876,N_13863);
nand U14311 (N_14311,N_13875,N_13828);
nand U14312 (N_14312,N_13936,N_13805);
and U14313 (N_14313,N_14010,N_14083);
or U14314 (N_14314,N_14091,N_13999);
and U14315 (N_14315,N_13850,N_13851);
and U14316 (N_14316,N_13806,N_13949);
nor U14317 (N_14317,N_14085,N_13893);
nor U14318 (N_14318,N_14027,N_14067);
nand U14319 (N_14319,N_13986,N_14051);
or U14320 (N_14320,N_13915,N_13816);
and U14321 (N_14321,N_14051,N_13831);
nand U14322 (N_14322,N_13922,N_13903);
nand U14323 (N_14323,N_14059,N_13827);
xnor U14324 (N_14324,N_13888,N_13956);
and U14325 (N_14325,N_13847,N_14078);
or U14326 (N_14326,N_14089,N_13844);
xor U14327 (N_14327,N_14044,N_13877);
and U14328 (N_14328,N_13972,N_13801);
xnor U14329 (N_14329,N_13945,N_13906);
and U14330 (N_14330,N_13876,N_14088);
or U14331 (N_14331,N_13929,N_14037);
or U14332 (N_14332,N_13889,N_13951);
xnor U14333 (N_14333,N_14021,N_13993);
nand U14334 (N_14334,N_14093,N_13847);
or U14335 (N_14335,N_13805,N_14013);
xor U14336 (N_14336,N_14024,N_14058);
and U14337 (N_14337,N_13990,N_13958);
and U14338 (N_14338,N_14071,N_14072);
nand U14339 (N_14339,N_13975,N_13856);
nand U14340 (N_14340,N_14039,N_13928);
nand U14341 (N_14341,N_14016,N_13828);
nor U14342 (N_14342,N_13898,N_13882);
or U14343 (N_14343,N_14034,N_13851);
nor U14344 (N_14344,N_14099,N_13858);
nor U14345 (N_14345,N_14094,N_13840);
and U14346 (N_14346,N_13835,N_13806);
xor U14347 (N_14347,N_13856,N_14020);
xor U14348 (N_14348,N_13901,N_14017);
and U14349 (N_14349,N_14043,N_13968);
nand U14350 (N_14350,N_13856,N_13941);
nand U14351 (N_14351,N_13802,N_13803);
or U14352 (N_14352,N_13933,N_13848);
or U14353 (N_14353,N_13958,N_13898);
or U14354 (N_14354,N_14044,N_14010);
nand U14355 (N_14355,N_13954,N_13941);
nor U14356 (N_14356,N_13985,N_14096);
nand U14357 (N_14357,N_13831,N_13982);
nand U14358 (N_14358,N_13882,N_14020);
or U14359 (N_14359,N_13821,N_14004);
or U14360 (N_14360,N_14058,N_13867);
nor U14361 (N_14361,N_13903,N_13944);
nor U14362 (N_14362,N_13907,N_13995);
xor U14363 (N_14363,N_13821,N_14006);
or U14364 (N_14364,N_13822,N_13951);
nor U14365 (N_14365,N_13965,N_13802);
or U14366 (N_14366,N_13936,N_13963);
nand U14367 (N_14367,N_13999,N_13865);
nand U14368 (N_14368,N_14025,N_13954);
nor U14369 (N_14369,N_14067,N_14066);
xnor U14370 (N_14370,N_13890,N_13806);
nand U14371 (N_14371,N_13919,N_13969);
nand U14372 (N_14372,N_13889,N_14000);
nand U14373 (N_14373,N_14077,N_13963);
and U14374 (N_14374,N_13892,N_13963);
nand U14375 (N_14375,N_13955,N_13813);
nand U14376 (N_14376,N_14068,N_13879);
or U14377 (N_14377,N_13901,N_13989);
nor U14378 (N_14378,N_14041,N_14085);
or U14379 (N_14379,N_14089,N_13851);
or U14380 (N_14380,N_13877,N_13816);
nor U14381 (N_14381,N_14078,N_13950);
or U14382 (N_14382,N_13838,N_13837);
nand U14383 (N_14383,N_13878,N_13910);
and U14384 (N_14384,N_13831,N_14079);
and U14385 (N_14385,N_14015,N_14049);
xnor U14386 (N_14386,N_13847,N_13849);
and U14387 (N_14387,N_14089,N_13823);
nand U14388 (N_14388,N_13976,N_13948);
and U14389 (N_14389,N_14008,N_14020);
nor U14390 (N_14390,N_13977,N_14084);
nor U14391 (N_14391,N_13907,N_13964);
nor U14392 (N_14392,N_13932,N_13891);
and U14393 (N_14393,N_13829,N_13813);
nand U14394 (N_14394,N_14078,N_14012);
and U14395 (N_14395,N_13836,N_13979);
nand U14396 (N_14396,N_13940,N_13819);
and U14397 (N_14397,N_14033,N_14080);
nor U14398 (N_14398,N_13845,N_14025);
and U14399 (N_14399,N_13918,N_13962);
nand U14400 (N_14400,N_14377,N_14167);
nor U14401 (N_14401,N_14114,N_14144);
or U14402 (N_14402,N_14360,N_14319);
or U14403 (N_14403,N_14315,N_14300);
nor U14404 (N_14404,N_14332,N_14340);
nand U14405 (N_14405,N_14223,N_14248);
or U14406 (N_14406,N_14250,N_14101);
nor U14407 (N_14407,N_14181,N_14294);
or U14408 (N_14408,N_14358,N_14229);
xor U14409 (N_14409,N_14322,N_14105);
nor U14410 (N_14410,N_14232,N_14234);
nand U14411 (N_14411,N_14190,N_14176);
nand U14412 (N_14412,N_14328,N_14110);
nand U14413 (N_14413,N_14126,N_14109);
nand U14414 (N_14414,N_14203,N_14194);
and U14415 (N_14415,N_14306,N_14266);
and U14416 (N_14416,N_14214,N_14254);
nand U14417 (N_14417,N_14382,N_14218);
nor U14418 (N_14418,N_14173,N_14333);
nand U14419 (N_14419,N_14125,N_14225);
and U14420 (N_14420,N_14261,N_14122);
xor U14421 (N_14421,N_14169,N_14163);
or U14422 (N_14422,N_14281,N_14345);
and U14423 (N_14423,N_14133,N_14280);
or U14424 (N_14424,N_14213,N_14212);
and U14425 (N_14425,N_14104,N_14171);
or U14426 (N_14426,N_14397,N_14244);
nor U14427 (N_14427,N_14170,N_14310);
and U14428 (N_14428,N_14269,N_14188);
or U14429 (N_14429,N_14222,N_14390);
or U14430 (N_14430,N_14320,N_14326);
xor U14431 (N_14431,N_14161,N_14355);
nand U14432 (N_14432,N_14151,N_14195);
and U14433 (N_14433,N_14327,N_14305);
and U14434 (N_14434,N_14227,N_14165);
or U14435 (N_14435,N_14153,N_14219);
nor U14436 (N_14436,N_14235,N_14143);
or U14437 (N_14437,N_14150,N_14283);
xor U14438 (N_14438,N_14210,N_14350);
and U14439 (N_14439,N_14359,N_14155);
nor U14440 (N_14440,N_14295,N_14289);
nor U14441 (N_14441,N_14292,N_14121);
xor U14442 (N_14442,N_14273,N_14318);
and U14443 (N_14443,N_14392,N_14338);
and U14444 (N_14444,N_14399,N_14282);
xnor U14445 (N_14445,N_14145,N_14346);
xor U14446 (N_14446,N_14367,N_14113);
or U14447 (N_14447,N_14226,N_14348);
xor U14448 (N_14448,N_14245,N_14287);
xnor U14449 (N_14449,N_14172,N_14231);
xor U14450 (N_14450,N_14362,N_14311);
nor U14451 (N_14451,N_14196,N_14380);
nand U14452 (N_14452,N_14263,N_14182);
nor U14453 (N_14453,N_14132,N_14260);
xnor U14454 (N_14454,N_14236,N_14271);
xor U14455 (N_14455,N_14383,N_14233);
xnor U14456 (N_14456,N_14308,N_14291);
and U14457 (N_14457,N_14100,N_14309);
nand U14458 (N_14458,N_14240,N_14381);
or U14459 (N_14459,N_14356,N_14174);
nor U14460 (N_14460,N_14258,N_14389);
nor U14461 (N_14461,N_14387,N_14352);
xnor U14462 (N_14462,N_14123,N_14374);
and U14463 (N_14463,N_14206,N_14279);
xor U14464 (N_14464,N_14243,N_14102);
nand U14465 (N_14465,N_14290,N_14317);
or U14466 (N_14466,N_14135,N_14168);
nor U14467 (N_14467,N_14252,N_14142);
and U14468 (N_14468,N_14321,N_14349);
nor U14469 (N_14469,N_14154,N_14303);
nand U14470 (N_14470,N_14127,N_14136);
nor U14471 (N_14471,N_14147,N_14187);
xor U14472 (N_14472,N_14118,N_14293);
nor U14473 (N_14473,N_14111,N_14204);
xor U14474 (N_14474,N_14164,N_14302);
and U14475 (N_14475,N_14334,N_14199);
nor U14476 (N_14476,N_14372,N_14158);
nor U14477 (N_14477,N_14301,N_14241);
nor U14478 (N_14478,N_14270,N_14185);
nand U14479 (N_14479,N_14140,N_14313);
xnor U14480 (N_14480,N_14298,N_14197);
and U14481 (N_14481,N_14146,N_14296);
xor U14482 (N_14482,N_14186,N_14156);
nor U14483 (N_14483,N_14242,N_14388);
xor U14484 (N_14484,N_14265,N_14139);
or U14485 (N_14485,N_14353,N_14286);
and U14486 (N_14486,N_14276,N_14278);
xnor U14487 (N_14487,N_14128,N_14157);
and U14488 (N_14488,N_14207,N_14189);
nor U14489 (N_14489,N_14220,N_14339);
or U14490 (N_14490,N_14344,N_14354);
or U14491 (N_14491,N_14217,N_14343);
nor U14492 (N_14492,N_14379,N_14394);
nand U14493 (N_14493,N_14268,N_14239);
xnor U14494 (N_14494,N_14277,N_14264);
and U14495 (N_14495,N_14272,N_14115);
or U14496 (N_14496,N_14341,N_14391);
and U14497 (N_14497,N_14216,N_14202);
nor U14498 (N_14498,N_14357,N_14209);
xor U14499 (N_14499,N_14112,N_14162);
nor U14500 (N_14500,N_14160,N_14325);
or U14501 (N_14501,N_14256,N_14373);
nand U14502 (N_14502,N_14347,N_14175);
or U14503 (N_14503,N_14205,N_14274);
or U14504 (N_14504,N_14342,N_14361);
xor U14505 (N_14505,N_14184,N_14363);
or U14506 (N_14506,N_14201,N_14335);
and U14507 (N_14507,N_14238,N_14108);
or U14508 (N_14508,N_14369,N_14124);
nor U14509 (N_14509,N_14183,N_14331);
xnor U14510 (N_14510,N_14370,N_14323);
nand U14511 (N_14511,N_14237,N_14259);
and U14512 (N_14512,N_14284,N_14221);
and U14513 (N_14513,N_14103,N_14191);
nor U14514 (N_14514,N_14178,N_14152);
and U14515 (N_14515,N_14368,N_14365);
and U14516 (N_14516,N_14288,N_14330);
xnor U14517 (N_14517,N_14230,N_14384);
nor U14518 (N_14518,N_14247,N_14398);
xnor U14519 (N_14519,N_14375,N_14116);
nand U14520 (N_14520,N_14299,N_14211);
nor U14521 (N_14521,N_14193,N_14149);
or U14522 (N_14522,N_14179,N_14378);
and U14523 (N_14523,N_14386,N_14200);
and U14524 (N_14524,N_14192,N_14215);
or U14525 (N_14525,N_14198,N_14285);
xnor U14526 (N_14526,N_14275,N_14249);
and U14527 (N_14527,N_14138,N_14366);
nor U14528 (N_14528,N_14267,N_14351);
nand U14529 (N_14529,N_14117,N_14107);
nand U14530 (N_14530,N_14134,N_14137);
nand U14531 (N_14531,N_14120,N_14129);
nor U14532 (N_14532,N_14329,N_14255);
and U14533 (N_14533,N_14324,N_14314);
nand U14534 (N_14534,N_14364,N_14312);
and U14535 (N_14535,N_14159,N_14251);
or U14536 (N_14536,N_14208,N_14180);
xor U14537 (N_14537,N_14376,N_14307);
nand U14538 (N_14538,N_14119,N_14395);
nand U14539 (N_14539,N_14166,N_14246);
or U14540 (N_14540,N_14130,N_14337);
nand U14541 (N_14541,N_14262,N_14396);
nand U14542 (N_14542,N_14371,N_14141);
xnor U14543 (N_14543,N_14228,N_14304);
or U14544 (N_14544,N_14385,N_14253);
xor U14545 (N_14545,N_14297,N_14316);
or U14546 (N_14546,N_14177,N_14336);
nor U14547 (N_14547,N_14106,N_14224);
nand U14548 (N_14548,N_14393,N_14257);
nor U14549 (N_14549,N_14131,N_14148);
nand U14550 (N_14550,N_14235,N_14188);
and U14551 (N_14551,N_14346,N_14283);
nor U14552 (N_14552,N_14328,N_14353);
nor U14553 (N_14553,N_14361,N_14161);
nor U14554 (N_14554,N_14281,N_14327);
nor U14555 (N_14555,N_14330,N_14146);
and U14556 (N_14556,N_14146,N_14363);
and U14557 (N_14557,N_14291,N_14123);
nand U14558 (N_14558,N_14111,N_14272);
or U14559 (N_14559,N_14110,N_14271);
or U14560 (N_14560,N_14295,N_14369);
nor U14561 (N_14561,N_14232,N_14156);
or U14562 (N_14562,N_14359,N_14269);
xor U14563 (N_14563,N_14133,N_14309);
xnor U14564 (N_14564,N_14115,N_14111);
or U14565 (N_14565,N_14382,N_14270);
xnor U14566 (N_14566,N_14178,N_14355);
nor U14567 (N_14567,N_14261,N_14162);
xor U14568 (N_14568,N_14278,N_14207);
xor U14569 (N_14569,N_14336,N_14185);
and U14570 (N_14570,N_14136,N_14388);
or U14571 (N_14571,N_14223,N_14391);
or U14572 (N_14572,N_14103,N_14334);
nand U14573 (N_14573,N_14299,N_14146);
or U14574 (N_14574,N_14199,N_14295);
xnor U14575 (N_14575,N_14141,N_14355);
or U14576 (N_14576,N_14182,N_14115);
nor U14577 (N_14577,N_14143,N_14240);
nand U14578 (N_14578,N_14268,N_14152);
and U14579 (N_14579,N_14272,N_14184);
nor U14580 (N_14580,N_14390,N_14238);
xnor U14581 (N_14581,N_14145,N_14152);
or U14582 (N_14582,N_14323,N_14207);
or U14583 (N_14583,N_14233,N_14102);
xor U14584 (N_14584,N_14112,N_14294);
and U14585 (N_14585,N_14388,N_14319);
nand U14586 (N_14586,N_14156,N_14365);
xor U14587 (N_14587,N_14264,N_14160);
nor U14588 (N_14588,N_14336,N_14205);
nand U14589 (N_14589,N_14107,N_14268);
xnor U14590 (N_14590,N_14147,N_14163);
nor U14591 (N_14591,N_14189,N_14193);
xnor U14592 (N_14592,N_14332,N_14274);
nor U14593 (N_14593,N_14311,N_14282);
xnor U14594 (N_14594,N_14109,N_14271);
nor U14595 (N_14595,N_14279,N_14356);
or U14596 (N_14596,N_14275,N_14161);
nand U14597 (N_14597,N_14342,N_14137);
and U14598 (N_14598,N_14141,N_14205);
or U14599 (N_14599,N_14327,N_14229);
xnor U14600 (N_14600,N_14247,N_14382);
nand U14601 (N_14601,N_14270,N_14307);
nor U14602 (N_14602,N_14205,N_14276);
and U14603 (N_14603,N_14190,N_14293);
xor U14604 (N_14604,N_14330,N_14162);
nand U14605 (N_14605,N_14250,N_14236);
nand U14606 (N_14606,N_14100,N_14135);
xnor U14607 (N_14607,N_14327,N_14117);
xor U14608 (N_14608,N_14281,N_14234);
nor U14609 (N_14609,N_14271,N_14144);
and U14610 (N_14610,N_14320,N_14268);
nor U14611 (N_14611,N_14369,N_14255);
or U14612 (N_14612,N_14325,N_14200);
nand U14613 (N_14613,N_14126,N_14337);
nand U14614 (N_14614,N_14394,N_14142);
xnor U14615 (N_14615,N_14201,N_14360);
nand U14616 (N_14616,N_14186,N_14109);
nand U14617 (N_14617,N_14126,N_14245);
nand U14618 (N_14618,N_14294,N_14139);
nand U14619 (N_14619,N_14251,N_14241);
nor U14620 (N_14620,N_14290,N_14269);
and U14621 (N_14621,N_14389,N_14104);
xnor U14622 (N_14622,N_14174,N_14263);
or U14623 (N_14623,N_14258,N_14163);
and U14624 (N_14624,N_14155,N_14166);
or U14625 (N_14625,N_14150,N_14370);
or U14626 (N_14626,N_14203,N_14328);
nor U14627 (N_14627,N_14312,N_14161);
nand U14628 (N_14628,N_14226,N_14392);
and U14629 (N_14629,N_14312,N_14131);
xor U14630 (N_14630,N_14325,N_14377);
or U14631 (N_14631,N_14295,N_14216);
nor U14632 (N_14632,N_14134,N_14232);
nor U14633 (N_14633,N_14351,N_14311);
nand U14634 (N_14634,N_14152,N_14171);
xor U14635 (N_14635,N_14390,N_14352);
or U14636 (N_14636,N_14172,N_14216);
and U14637 (N_14637,N_14314,N_14181);
or U14638 (N_14638,N_14163,N_14249);
nand U14639 (N_14639,N_14365,N_14281);
and U14640 (N_14640,N_14132,N_14315);
or U14641 (N_14641,N_14208,N_14118);
or U14642 (N_14642,N_14305,N_14336);
nand U14643 (N_14643,N_14301,N_14120);
nor U14644 (N_14644,N_14218,N_14358);
and U14645 (N_14645,N_14157,N_14354);
or U14646 (N_14646,N_14382,N_14110);
xor U14647 (N_14647,N_14386,N_14192);
nor U14648 (N_14648,N_14334,N_14170);
xnor U14649 (N_14649,N_14159,N_14195);
or U14650 (N_14650,N_14241,N_14355);
or U14651 (N_14651,N_14314,N_14306);
and U14652 (N_14652,N_14369,N_14387);
nor U14653 (N_14653,N_14296,N_14374);
or U14654 (N_14654,N_14215,N_14319);
nor U14655 (N_14655,N_14251,N_14111);
xor U14656 (N_14656,N_14163,N_14113);
xnor U14657 (N_14657,N_14398,N_14177);
and U14658 (N_14658,N_14327,N_14105);
nor U14659 (N_14659,N_14151,N_14207);
or U14660 (N_14660,N_14147,N_14341);
or U14661 (N_14661,N_14108,N_14389);
or U14662 (N_14662,N_14244,N_14366);
nor U14663 (N_14663,N_14148,N_14184);
or U14664 (N_14664,N_14196,N_14234);
or U14665 (N_14665,N_14378,N_14207);
or U14666 (N_14666,N_14211,N_14191);
or U14667 (N_14667,N_14324,N_14124);
or U14668 (N_14668,N_14114,N_14366);
xor U14669 (N_14669,N_14127,N_14189);
or U14670 (N_14670,N_14295,N_14316);
nand U14671 (N_14671,N_14204,N_14366);
or U14672 (N_14672,N_14157,N_14314);
and U14673 (N_14673,N_14274,N_14366);
nor U14674 (N_14674,N_14356,N_14315);
nand U14675 (N_14675,N_14291,N_14320);
xor U14676 (N_14676,N_14100,N_14396);
nand U14677 (N_14677,N_14322,N_14392);
xor U14678 (N_14678,N_14167,N_14199);
and U14679 (N_14679,N_14129,N_14168);
and U14680 (N_14680,N_14243,N_14103);
and U14681 (N_14681,N_14131,N_14153);
xnor U14682 (N_14682,N_14364,N_14238);
nand U14683 (N_14683,N_14209,N_14300);
and U14684 (N_14684,N_14304,N_14130);
or U14685 (N_14685,N_14335,N_14186);
xnor U14686 (N_14686,N_14279,N_14357);
and U14687 (N_14687,N_14370,N_14158);
nand U14688 (N_14688,N_14393,N_14361);
or U14689 (N_14689,N_14180,N_14289);
nand U14690 (N_14690,N_14209,N_14319);
nor U14691 (N_14691,N_14236,N_14247);
or U14692 (N_14692,N_14228,N_14191);
or U14693 (N_14693,N_14197,N_14354);
nand U14694 (N_14694,N_14211,N_14276);
xnor U14695 (N_14695,N_14388,N_14345);
xor U14696 (N_14696,N_14152,N_14204);
xor U14697 (N_14697,N_14137,N_14121);
xnor U14698 (N_14698,N_14321,N_14366);
xor U14699 (N_14699,N_14188,N_14340);
or U14700 (N_14700,N_14593,N_14613);
and U14701 (N_14701,N_14590,N_14610);
nor U14702 (N_14702,N_14543,N_14499);
nor U14703 (N_14703,N_14554,N_14415);
nand U14704 (N_14704,N_14609,N_14502);
xor U14705 (N_14705,N_14454,N_14421);
xor U14706 (N_14706,N_14433,N_14653);
nand U14707 (N_14707,N_14620,N_14444);
nor U14708 (N_14708,N_14650,N_14580);
xnor U14709 (N_14709,N_14474,N_14511);
xnor U14710 (N_14710,N_14440,N_14513);
nand U14711 (N_14711,N_14697,N_14498);
nor U14712 (N_14712,N_14638,N_14460);
and U14713 (N_14713,N_14503,N_14633);
or U14714 (N_14714,N_14642,N_14425);
nor U14715 (N_14715,N_14501,N_14473);
xor U14716 (N_14716,N_14693,N_14599);
nor U14717 (N_14717,N_14528,N_14657);
xor U14718 (N_14718,N_14504,N_14521);
xor U14719 (N_14719,N_14436,N_14644);
nand U14720 (N_14720,N_14438,N_14542);
xnor U14721 (N_14721,N_14641,N_14466);
nor U14722 (N_14722,N_14488,N_14594);
nor U14723 (N_14723,N_14408,N_14661);
and U14724 (N_14724,N_14598,N_14667);
or U14725 (N_14725,N_14495,N_14690);
and U14726 (N_14726,N_14637,N_14559);
nand U14727 (N_14727,N_14486,N_14648);
and U14728 (N_14728,N_14680,N_14519);
nand U14729 (N_14729,N_14500,N_14682);
xor U14730 (N_14730,N_14489,N_14573);
nand U14731 (N_14731,N_14403,N_14464);
nand U14732 (N_14732,N_14518,N_14691);
xor U14733 (N_14733,N_14683,N_14475);
xnor U14734 (N_14734,N_14537,N_14617);
nor U14735 (N_14735,N_14666,N_14558);
nor U14736 (N_14736,N_14484,N_14557);
nand U14737 (N_14737,N_14628,N_14417);
nand U14738 (N_14738,N_14562,N_14468);
xor U14739 (N_14739,N_14532,N_14688);
or U14740 (N_14740,N_14659,N_14626);
and U14741 (N_14741,N_14449,N_14566);
nand U14742 (N_14742,N_14527,N_14625);
and U14743 (N_14743,N_14509,N_14674);
nand U14744 (N_14744,N_14512,N_14589);
or U14745 (N_14745,N_14685,N_14616);
or U14746 (N_14746,N_14561,N_14526);
nor U14747 (N_14747,N_14608,N_14606);
or U14748 (N_14748,N_14665,N_14551);
nand U14749 (N_14749,N_14514,N_14675);
xnor U14750 (N_14750,N_14645,N_14535);
xnor U14751 (N_14751,N_14510,N_14420);
and U14752 (N_14752,N_14695,N_14586);
xnor U14753 (N_14753,N_14602,N_14406);
nor U14754 (N_14754,N_14435,N_14604);
or U14755 (N_14755,N_14465,N_14422);
or U14756 (N_14756,N_14699,N_14446);
nand U14757 (N_14757,N_14624,N_14471);
nand U14758 (N_14758,N_14605,N_14582);
nand U14759 (N_14759,N_14560,N_14478);
or U14760 (N_14760,N_14579,N_14467);
xor U14761 (N_14761,N_14640,N_14588);
nand U14762 (N_14762,N_14541,N_14545);
and U14763 (N_14763,N_14572,N_14552);
nor U14764 (N_14764,N_14441,N_14491);
nand U14765 (N_14765,N_14490,N_14540);
xor U14766 (N_14766,N_14568,N_14684);
xnor U14767 (N_14767,N_14564,N_14563);
and U14768 (N_14768,N_14450,N_14622);
nor U14769 (N_14769,N_14643,N_14458);
nor U14770 (N_14770,N_14480,N_14538);
nand U14771 (N_14771,N_14544,N_14612);
and U14772 (N_14772,N_14672,N_14636);
nand U14773 (N_14773,N_14445,N_14635);
nor U14774 (N_14774,N_14456,N_14439);
or U14775 (N_14775,N_14546,N_14671);
nor U14776 (N_14776,N_14429,N_14451);
xor U14777 (N_14777,N_14600,N_14427);
or U14778 (N_14778,N_14479,N_14487);
or U14779 (N_14779,N_14656,N_14505);
nand U14780 (N_14780,N_14404,N_14669);
and U14781 (N_14781,N_14461,N_14536);
nor U14782 (N_14782,N_14520,N_14426);
nand U14783 (N_14783,N_14418,N_14647);
and U14784 (N_14784,N_14492,N_14522);
or U14785 (N_14785,N_14658,N_14601);
xnor U14786 (N_14786,N_14575,N_14481);
or U14787 (N_14787,N_14569,N_14432);
nor U14788 (N_14788,N_14652,N_14632);
nand U14789 (N_14789,N_14419,N_14681);
or U14790 (N_14790,N_14677,N_14455);
or U14791 (N_14791,N_14494,N_14621);
and U14792 (N_14792,N_14649,N_14660);
nand U14793 (N_14793,N_14607,N_14452);
nor U14794 (N_14794,N_14443,N_14413);
and U14795 (N_14795,N_14430,N_14409);
nand U14796 (N_14796,N_14523,N_14623);
xor U14797 (N_14797,N_14547,N_14462);
and U14798 (N_14798,N_14634,N_14453);
nor U14799 (N_14799,N_14670,N_14470);
or U14800 (N_14800,N_14410,N_14407);
or U14801 (N_14801,N_14567,N_14463);
xnor U14802 (N_14802,N_14581,N_14549);
and U14803 (N_14803,N_14428,N_14459);
xor U14804 (N_14804,N_14577,N_14534);
nand U14805 (N_14805,N_14469,N_14485);
nand U14806 (N_14806,N_14571,N_14507);
xnor U14807 (N_14807,N_14556,N_14423);
nand U14808 (N_14808,N_14574,N_14506);
nor U14809 (N_14809,N_14664,N_14493);
and U14810 (N_14810,N_14411,N_14483);
nand U14811 (N_14811,N_14457,N_14629);
and U14812 (N_14812,N_14584,N_14663);
or U14813 (N_14813,N_14497,N_14482);
xnor U14814 (N_14814,N_14595,N_14583);
nor U14815 (N_14815,N_14401,N_14508);
xnor U14816 (N_14816,N_14694,N_14614);
xnor U14817 (N_14817,N_14565,N_14591);
nor U14818 (N_14818,N_14477,N_14578);
nand U14819 (N_14819,N_14550,N_14603);
nand U14820 (N_14820,N_14539,N_14442);
xnor U14821 (N_14821,N_14585,N_14596);
nand U14822 (N_14822,N_14627,N_14416);
and U14823 (N_14823,N_14531,N_14619);
and U14824 (N_14824,N_14679,N_14496);
nand U14825 (N_14825,N_14687,N_14525);
nand U14826 (N_14826,N_14548,N_14692);
nand U14827 (N_14827,N_14448,N_14696);
and U14828 (N_14828,N_14570,N_14587);
or U14829 (N_14829,N_14630,N_14424);
nand U14830 (N_14830,N_14592,N_14597);
and U14831 (N_14831,N_14524,N_14651);
nor U14832 (N_14832,N_14676,N_14405);
xor U14833 (N_14833,N_14515,N_14516);
and U14834 (N_14834,N_14402,N_14529);
nor U14835 (N_14835,N_14553,N_14412);
xnor U14836 (N_14836,N_14434,N_14678);
and U14837 (N_14837,N_14673,N_14639);
or U14838 (N_14838,N_14686,N_14631);
xor U14839 (N_14839,N_14437,N_14447);
nor U14840 (N_14840,N_14472,N_14476);
nor U14841 (N_14841,N_14400,N_14668);
xor U14842 (N_14842,N_14533,N_14654);
or U14843 (N_14843,N_14618,N_14655);
and U14844 (N_14844,N_14646,N_14615);
and U14845 (N_14845,N_14431,N_14662);
or U14846 (N_14846,N_14517,N_14530);
nand U14847 (N_14847,N_14414,N_14576);
and U14848 (N_14848,N_14689,N_14555);
xor U14849 (N_14849,N_14698,N_14611);
nor U14850 (N_14850,N_14456,N_14480);
xor U14851 (N_14851,N_14658,N_14635);
nand U14852 (N_14852,N_14527,N_14612);
or U14853 (N_14853,N_14526,N_14592);
nor U14854 (N_14854,N_14644,N_14606);
and U14855 (N_14855,N_14422,N_14669);
and U14856 (N_14856,N_14479,N_14434);
or U14857 (N_14857,N_14457,N_14573);
nor U14858 (N_14858,N_14456,N_14504);
xnor U14859 (N_14859,N_14412,N_14453);
or U14860 (N_14860,N_14434,N_14683);
nor U14861 (N_14861,N_14563,N_14573);
and U14862 (N_14862,N_14606,N_14671);
nor U14863 (N_14863,N_14605,N_14422);
xnor U14864 (N_14864,N_14518,N_14478);
nor U14865 (N_14865,N_14423,N_14409);
or U14866 (N_14866,N_14477,N_14471);
and U14867 (N_14867,N_14444,N_14439);
and U14868 (N_14868,N_14564,N_14633);
and U14869 (N_14869,N_14407,N_14450);
nor U14870 (N_14870,N_14487,N_14624);
nand U14871 (N_14871,N_14633,N_14563);
xor U14872 (N_14872,N_14410,N_14691);
nand U14873 (N_14873,N_14616,N_14648);
nand U14874 (N_14874,N_14656,N_14601);
xnor U14875 (N_14875,N_14622,N_14419);
nor U14876 (N_14876,N_14426,N_14627);
and U14877 (N_14877,N_14646,N_14674);
or U14878 (N_14878,N_14547,N_14482);
nand U14879 (N_14879,N_14427,N_14691);
nor U14880 (N_14880,N_14605,N_14678);
nor U14881 (N_14881,N_14404,N_14472);
and U14882 (N_14882,N_14591,N_14544);
nand U14883 (N_14883,N_14554,N_14453);
xnor U14884 (N_14884,N_14618,N_14641);
nand U14885 (N_14885,N_14430,N_14487);
and U14886 (N_14886,N_14425,N_14544);
xor U14887 (N_14887,N_14569,N_14682);
nand U14888 (N_14888,N_14638,N_14666);
xnor U14889 (N_14889,N_14607,N_14477);
xnor U14890 (N_14890,N_14499,N_14512);
nand U14891 (N_14891,N_14625,N_14484);
and U14892 (N_14892,N_14660,N_14602);
nor U14893 (N_14893,N_14581,N_14697);
and U14894 (N_14894,N_14489,N_14612);
and U14895 (N_14895,N_14560,N_14592);
or U14896 (N_14896,N_14524,N_14482);
xor U14897 (N_14897,N_14518,N_14557);
or U14898 (N_14898,N_14515,N_14408);
nor U14899 (N_14899,N_14529,N_14626);
xnor U14900 (N_14900,N_14543,N_14616);
nor U14901 (N_14901,N_14541,N_14432);
or U14902 (N_14902,N_14623,N_14456);
or U14903 (N_14903,N_14457,N_14486);
xor U14904 (N_14904,N_14475,N_14649);
xnor U14905 (N_14905,N_14543,N_14620);
or U14906 (N_14906,N_14607,N_14479);
or U14907 (N_14907,N_14503,N_14558);
nor U14908 (N_14908,N_14683,N_14467);
nand U14909 (N_14909,N_14416,N_14668);
xnor U14910 (N_14910,N_14612,N_14457);
nand U14911 (N_14911,N_14527,N_14448);
nor U14912 (N_14912,N_14647,N_14661);
xor U14913 (N_14913,N_14493,N_14453);
or U14914 (N_14914,N_14500,N_14475);
xnor U14915 (N_14915,N_14400,N_14462);
nor U14916 (N_14916,N_14623,N_14421);
xnor U14917 (N_14917,N_14586,N_14566);
nand U14918 (N_14918,N_14418,N_14571);
xor U14919 (N_14919,N_14440,N_14416);
and U14920 (N_14920,N_14567,N_14526);
nand U14921 (N_14921,N_14672,N_14666);
nor U14922 (N_14922,N_14579,N_14646);
nor U14923 (N_14923,N_14415,N_14510);
and U14924 (N_14924,N_14604,N_14453);
nand U14925 (N_14925,N_14671,N_14502);
and U14926 (N_14926,N_14657,N_14494);
xnor U14927 (N_14927,N_14403,N_14693);
xor U14928 (N_14928,N_14564,N_14454);
nor U14929 (N_14929,N_14619,N_14472);
and U14930 (N_14930,N_14432,N_14584);
and U14931 (N_14931,N_14488,N_14644);
and U14932 (N_14932,N_14584,N_14582);
or U14933 (N_14933,N_14535,N_14518);
nand U14934 (N_14934,N_14609,N_14593);
or U14935 (N_14935,N_14671,N_14442);
or U14936 (N_14936,N_14605,N_14631);
and U14937 (N_14937,N_14634,N_14699);
or U14938 (N_14938,N_14522,N_14443);
or U14939 (N_14939,N_14480,N_14552);
nand U14940 (N_14940,N_14520,N_14557);
xnor U14941 (N_14941,N_14542,N_14434);
xor U14942 (N_14942,N_14625,N_14566);
nor U14943 (N_14943,N_14694,N_14602);
nand U14944 (N_14944,N_14596,N_14513);
nor U14945 (N_14945,N_14670,N_14680);
nor U14946 (N_14946,N_14578,N_14425);
nor U14947 (N_14947,N_14569,N_14507);
and U14948 (N_14948,N_14407,N_14554);
or U14949 (N_14949,N_14533,N_14623);
nor U14950 (N_14950,N_14445,N_14478);
nor U14951 (N_14951,N_14581,N_14437);
or U14952 (N_14952,N_14659,N_14499);
nand U14953 (N_14953,N_14672,N_14557);
nor U14954 (N_14954,N_14688,N_14655);
xor U14955 (N_14955,N_14620,N_14428);
and U14956 (N_14956,N_14476,N_14641);
nor U14957 (N_14957,N_14516,N_14443);
and U14958 (N_14958,N_14413,N_14640);
and U14959 (N_14959,N_14445,N_14630);
xnor U14960 (N_14960,N_14473,N_14546);
xnor U14961 (N_14961,N_14643,N_14505);
xnor U14962 (N_14962,N_14609,N_14411);
xnor U14963 (N_14963,N_14610,N_14507);
xor U14964 (N_14964,N_14424,N_14518);
nor U14965 (N_14965,N_14449,N_14657);
xnor U14966 (N_14966,N_14624,N_14698);
nand U14967 (N_14967,N_14438,N_14464);
nand U14968 (N_14968,N_14480,N_14554);
and U14969 (N_14969,N_14602,N_14438);
nand U14970 (N_14970,N_14647,N_14569);
or U14971 (N_14971,N_14487,N_14472);
xor U14972 (N_14972,N_14689,N_14599);
and U14973 (N_14973,N_14699,N_14554);
nor U14974 (N_14974,N_14400,N_14697);
or U14975 (N_14975,N_14442,N_14483);
nand U14976 (N_14976,N_14586,N_14531);
and U14977 (N_14977,N_14595,N_14682);
nand U14978 (N_14978,N_14688,N_14485);
nand U14979 (N_14979,N_14573,N_14411);
xor U14980 (N_14980,N_14604,N_14569);
and U14981 (N_14981,N_14477,N_14594);
nor U14982 (N_14982,N_14477,N_14621);
nand U14983 (N_14983,N_14468,N_14510);
and U14984 (N_14984,N_14448,N_14498);
nor U14985 (N_14985,N_14644,N_14610);
or U14986 (N_14986,N_14435,N_14554);
nand U14987 (N_14987,N_14567,N_14401);
or U14988 (N_14988,N_14575,N_14568);
nor U14989 (N_14989,N_14488,N_14691);
or U14990 (N_14990,N_14473,N_14577);
nand U14991 (N_14991,N_14512,N_14682);
xor U14992 (N_14992,N_14409,N_14622);
and U14993 (N_14993,N_14511,N_14681);
nor U14994 (N_14994,N_14509,N_14443);
or U14995 (N_14995,N_14512,N_14671);
xor U14996 (N_14996,N_14520,N_14659);
nor U14997 (N_14997,N_14538,N_14477);
xor U14998 (N_14998,N_14588,N_14401);
or U14999 (N_14999,N_14520,N_14490);
nand UO_0 (O_0,N_14957,N_14922);
nor UO_1 (O_1,N_14927,N_14931);
nand UO_2 (O_2,N_14924,N_14987);
xnor UO_3 (O_3,N_14941,N_14755);
nor UO_4 (O_4,N_14965,N_14949);
nand UO_5 (O_5,N_14963,N_14792);
or UO_6 (O_6,N_14991,N_14892);
nor UO_7 (O_7,N_14801,N_14928);
xnor UO_8 (O_8,N_14764,N_14875);
nand UO_9 (O_9,N_14853,N_14909);
xor UO_10 (O_10,N_14935,N_14877);
xor UO_11 (O_11,N_14911,N_14727);
and UO_12 (O_12,N_14845,N_14769);
or UO_13 (O_13,N_14919,N_14710);
xnor UO_14 (O_14,N_14937,N_14902);
or UO_15 (O_15,N_14873,N_14956);
or UO_16 (O_16,N_14894,N_14700);
xor UO_17 (O_17,N_14901,N_14844);
nand UO_18 (O_18,N_14788,N_14772);
nand UO_19 (O_19,N_14910,N_14785);
xor UO_20 (O_20,N_14882,N_14849);
and UO_21 (O_21,N_14944,N_14802);
or UO_22 (O_22,N_14988,N_14899);
or UO_23 (O_23,N_14833,N_14945);
xor UO_24 (O_24,N_14846,N_14808);
nand UO_25 (O_25,N_14854,N_14748);
nor UO_26 (O_26,N_14930,N_14790);
nor UO_27 (O_27,N_14819,N_14992);
nand UO_28 (O_28,N_14774,N_14848);
and UO_29 (O_29,N_14806,N_14811);
xor UO_30 (O_30,N_14852,N_14722);
and UO_31 (O_31,N_14893,N_14820);
nor UO_32 (O_32,N_14870,N_14720);
nand UO_33 (O_33,N_14876,N_14714);
xor UO_34 (O_34,N_14797,N_14803);
nor UO_35 (O_35,N_14961,N_14867);
xor UO_36 (O_36,N_14721,N_14718);
xnor UO_37 (O_37,N_14864,N_14975);
nor UO_38 (O_38,N_14994,N_14998);
or UO_39 (O_39,N_14881,N_14871);
or UO_40 (O_40,N_14768,N_14952);
or UO_41 (O_41,N_14827,N_14923);
and UO_42 (O_42,N_14842,N_14766);
and UO_43 (O_43,N_14744,N_14787);
nor UO_44 (O_44,N_14725,N_14807);
nand UO_45 (O_45,N_14978,N_14891);
or UO_46 (O_46,N_14968,N_14799);
nor UO_47 (O_47,N_14783,N_14775);
or UO_48 (O_48,N_14826,N_14759);
xor UO_49 (O_49,N_14760,N_14989);
and UO_50 (O_50,N_14778,N_14859);
and UO_51 (O_51,N_14995,N_14861);
and UO_52 (O_52,N_14835,N_14789);
nor UO_53 (O_53,N_14750,N_14960);
nand UO_54 (O_54,N_14791,N_14883);
nand UO_55 (O_55,N_14834,N_14777);
nand UO_56 (O_56,N_14985,N_14981);
and UO_57 (O_57,N_14816,N_14967);
and UO_58 (O_58,N_14889,N_14798);
and UO_59 (O_59,N_14959,N_14817);
nand UO_60 (O_60,N_14925,N_14947);
and UO_61 (O_61,N_14724,N_14838);
nor UO_62 (O_62,N_14805,N_14885);
nor UO_63 (O_63,N_14869,N_14966);
nand UO_64 (O_64,N_14979,N_14784);
nand UO_65 (O_65,N_14762,N_14824);
and UO_66 (O_66,N_14971,N_14977);
nand UO_67 (O_67,N_14735,N_14962);
nand UO_68 (O_68,N_14916,N_14840);
nor UO_69 (O_69,N_14712,N_14708);
and UO_70 (O_70,N_14749,N_14950);
nand UO_71 (O_71,N_14898,N_14914);
or UO_72 (O_72,N_14936,N_14990);
or UO_73 (O_73,N_14993,N_14939);
and UO_74 (O_74,N_14831,N_14758);
and UO_75 (O_75,N_14955,N_14716);
nand UO_76 (O_76,N_14997,N_14886);
and UO_77 (O_77,N_14887,N_14739);
or UO_78 (O_78,N_14874,N_14756);
nor UO_79 (O_79,N_14776,N_14970);
and UO_80 (O_80,N_14974,N_14781);
xor UO_81 (O_81,N_14736,N_14723);
xnor UO_82 (O_82,N_14732,N_14743);
or UO_83 (O_83,N_14832,N_14953);
and UO_84 (O_84,N_14863,N_14813);
and UO_85 (O_85,N_14866,N_14706);
and UO_86 (O_86,N_14851,N_14946);
or UO_87 (O_87,N_14932,N_14913);
nor UO_88 (O_88,N_14809,N_14810);
and UO_89 (O_89,N_14983,N_14742);
xor UO_90 (O_90,N_14969,N_14976);
nand UO_91 (O_91,N_14929,N_14754);
nand UO_92 (O_92,N_14812,N_14704);
nor UO_93 (O_93,N_14707,N_14821);
nand UO_94 (O_94,N_14918,N_14940);
xor UO_95 (O_95,N_14713,N_14737);
nor UO_96 (O_96,N_14829,N_14763);
or UO_97 (O_97,N_14822,N_14715);
or UO_98 (O_98,N_14717,N_14841);
nor UO_99 (O_99,N_14839,N_14794);
and UO_100 (O_100,N_14795,N_14757);
nand UO_101 (O_101,N_14729,N_14830);
xor UO_102 (O_102,N_14917,N_14906);
xor UO_103 (O_103,N_14980,N_14709);
and UO_104 (O_104,N_14771,N_14765);
xor UO_105 (O_105,N_14986,N_14862);
nor UO_106 (O_106,N_14745,N_14879);
and UO_107 (O_107,N_14843,N_14746);
or UO_108 (O_108,N_14855,N_14825);
or UO_109 (O_109,N_14733,N_14999);
and UO_110 (O_110,N_14857,N_14740);
nor UO_111 (O_111,N_14815,N_14823);
nand UO_112 (O_112,N_14954,N_14761);
nor UO_113 (O_113,N_14878,N_14890);
and UO_114 (O_114,N_14782,N_14958);
or UO_115 (O_115,N_14731,N_14938);
and UO_116 (O_116,N_14793,N_14738);
xnor UO_117 (O_117,N_14752,N_14828);
and UO_118 (O_118,N_14888,N_14818);
nand UO_119 (O_119,N_14767,N_14734);
nor UO_120 (O_120,N_14933,N_14984);
xor UO_121 (O_121,N_14921,N_14858);
nor UO_122 (O_122,N_14711,N_14900);
or UO_123 (O_123,N_14880,N_14973);
nand UO_124 (O_124,N_14920,N_14896);
nor UO_125 (O_125,N_14747,N_14796);
xnor UO_126 (O_126,N_14856,N_14905);
and UO_127 (O_127,N_14860,N_14719);
nor UO_128 (O_128,N_14779,N_14753);
xnor UO_129 (O_129,N_14728,N_14703);
xnor UO_130 (O_130,N_14751,N_14912);
and UO_131 (O_131,N_14705,N_14926);
xor UO_132 (O_132,N_14996,N_14972);
and UO_133 (O_133,N_14726,N_14730);
nand UO_134 (O_134,N_14903,N_14908);
nor UO_135 (O_135,N_14837,N_14865);
nand UO_136 (O_136,N_14701,N_14895);
xnor UO_137 (O_137,N_14800,N_14942);
and UO_138 (O_138,N_14814,N_14897);
nor UO_139 (O_139,N_14915,N_14904);
and UO_140 (O_140,N_14804,N_14982);
or UO_141 (O_141,N_14773,N_14836);
xnor UO_142 (O_142,N_14702,N_14786);
nand UO_143 (O_143,N_14964,N_14847);
nand UO_144 (O_144,N_14884,N_14907);
xnor UO_145 (O_145,N_14770,N_14780);
nand UO_146 (O_146,N_14868,N_14934);
xnor UO_147 (O_147,N_14872,N_14741);
and UO_148 (O_148,N_14943,N_14951);
or UO_149 (O_149,N_14850,N_14948);
nor UO_150 (O_150,N_14968,N_14920);
or UO_151 (O_151,N_14743,N_14708);
or UO_152 (O_152,N_14863,N_14870);
nand UO_153 (O_153,N_14817,N_14763);
or UO_154 (O_154,N_14839,N_14873);
nand UO_155 (O_155,N_14990,N_14709);
and UO_156 (O_156,N_14811,N_14865);
or UO_157 (O_157,N_14800,N_14771);
nand UO_158 (O_158,N_14816,N_14715);
or UO_159 (O_159,N_14749,N_14944);
xor UO_160 (O_160,N_14853,N_14769);
and UO_161 (O_161,N_14841,N_14771);
and UO_162 (O_162,N_14890,N_14923);
or UO_163 (O_163,N_14701,N_14931);
and UO_164 (O_164,N_14795,N_14818);
nand UO_165 (O_165,N_14748,N_14723);
nor UO_166 (O_166,N_14789,N_14846);
and UO_167 (O_167,N_14833,N_14812);
and UO_168 (O_168,N_14987,N_14761);
nor UO_169 (O_169,N_14811,N_14928);
and UO_170 (O_170,N_14854,N_14714);
nand UO_171 (O_171,N_14921,N_14987);
xnor UO_172 (O_172,N_14984,N_14735);
or UO_173 (O_173,N_14785,N_14765);
nor UO_174 (O_174,N_14961,N_14722);
nor UO_175 (O_175,N_14832,N_14985);
or UO_176 (O_176,N_14773,N_14797);
nor UO_177 (O_177,N_14954,N_14708);
nand UO_178 (O_178,N_14833,N_14779);
and UO_179 (O_179,N_14878,N_14749);
and UO_180 (O_180,N_14948,N_14890);
xor UO_181 (O_181,N_14857,N_14802);
nor UO_182 (O_182,N_14705,N_14720);
and UO_183 (O_183,N_14967,N_14728);
xor UO_184 (O_184,N_14858,N_14819);
xnor UO_185 (O_185,N_14969,N_14840);
and UO_186 (O_186,N_14926,N_14858);
nor UO_187 (O_187,N_14955,N_14998);
or UO_188 (O_188,N_14730,N_14810);
or UO_189 (O_189,N_14858,N_14842);
or UO_190 (O_190,N_14828,N_14804);
nand UO_191 (O_191,N_14953,N_14943);
nor UO_192 (O_192,N_14950,N_14789);
or UO_193 (O_193,N_14755,N_14920);
xnor UO_194 (O_194,N_14785,N_14992);
nand UO_195 (O_195,N_14894,N_14853);
or UO_196 (O_196,N_14706,N_14928);
xor UO_197 (O_197,N_14805,N_14903);
xnor UO_198 (O_198,N_14710,N_14838);
or UO_199 (O_199,N_14934,N_14850);
and UO_200 (O_200,N_14862,N_14961);
xor UO_201 (O_201,N_14917,N_14771);
nand UO_202 (O_202,N_14911,N_14840);
nor UO_203 (O_203,N_14827,N_14774);
nor UO_204 (O_204,N_14843,N_14877);
and UO_205 (O_205,N_14707,N_14867);
xor UO_206 (O_206,N_14926,N_14872);
or UO_207 (O_207,N_14797,N_14826);
nand UO_208 (O_208,N_14969,N_14759);
and UO_209 (O_209,N_14709,N_14860);
and UO_210 (O_210,N_14731,N_14965);
or UO_211 (O_211,N_14981,N_14869);
or UO_212 (O_212,N_14942,N_14908);
and UO_213 (O_213,N_14787,N_14755);
nand UO_214 (O_214,N_14784,N_14933);
xor UO_215 (O_215,N_14945,N_14702);
nor UO_216 (O_216,N_14911,N_14905);
xnor UO_217 (O_217,N_14747,N_14718);
nand UO_218 (O_218,N_14730,N_14961);
xor UO_219 (O_219,N_14782,N_14883);
nor UO_220 (O_220,N_14756,N_14778);
and UO_221 (O_221,N_14963,N_14904);
nor UO_222 (O_222,N_14701,N_14733);
nor UO_223 (O_223,N_14984,N_14703);
or UO_224 (O_224,N_14843,N_14973);
xor UO_225 (O_225,N_14849,N_14771);
nand UO_226 (O_226,N_14772,N_14978);
nor UO_227 (O_227,N_14770,N_14981);
and UO_228 (O_228,N_14994,N_14926);
and UO_229 (O_229,N_14987,N_14714);
nor UO_230 (O_230,N_14936,N_14734);
nand UO_231 (O_231,N_14814,N_14781);
nand UO_232 (O_232,N_14776,N_14932);
nor UO_233 (O_233,N_14781,N_14778);
and UO_234 (O_234,N_14709,N_14833);
or UO_235 (O_235,N_14999,N_14856);
nand UO_236 (O_236,N_14893,N_14766);
or UO_237 (O_237,N_14718,N_14782);
nor UO_238 (O_238,N_14735,N_14723);
xnor UO_239 (O_239,N_14808,N_14989);
nor UO_240 (O_240,N_14744,N_14824);
or UO_241 (O_241,N_14715,N_14930);
xor UO_242 (O_242,N_14736,N_14967);
or UO_243 (O_243,N_14969,N_14926);
and UO_244 (O_244,N_14921,N_14710);
or UO_245 (O_245,N_14904,N_14961);
or UO_246 (O_246,N_14721,N_14769);
nand UO_247 (O_247,N_14713,N_14728);
or UO_248 (O_248,N_14849,N_14886);
and UO_249 (O_249,N_14857,N_14843);
or UO_250 (O_250,N_14769,N_14844);
nand UO_251 (O_251,N_14756,N_14939);
nand UO_252 (O_252,N_14897,N_14710);
nand UO_253 (O_253,N_14710,N_14773);
or UO_254 (O_254,N_14896,N_14703);
xnor UO_255 (O_255,N_14930,N_14712);
xor UO_256 (O_256,N_14994,N_14732);
or UO_257 (O_257,N_14721,N_14930);
xor UO_258 (O_258,N_14967,N_14959);
or UO_259 (O_259,N_14763,N_14881);
and UO_260 (O_260,N_14745,N_14805);
or UO_261 (O_261,N_14959,N_14878);
nor UO_262 (O_262,N_14919,N_14934);
xnor UO_263 (O_263,N_14705,N_14879);
nor UO_264 (O_264,N_14861,N_14978);
nand UO_265 (O_265,N_14887,N_14759);
nor UO_266 (O_266,N_14791,N_14794);
nor UO_267 (O_267,N_14769,N_14792);
and UO_268 (O_268,N_14938,N_14965);
xor UO_269 (O_269,N_14931,N_14829);
xnor UO_270 (O_270,N_14902,N_14868);
nand UO_271 (O_271,N_14956,N_14895);
and UO_272 (O_272,N_14873,N_14738);
and UO_273 (O_273,N_14992,N_14813);
xor UO_274 (O_274,N_14976,N_14796);
or UO_275 (O_275,N_14854,N_14815);
and UO_276 (O_276,N_14944,N_14792);
nor UO_277 (O_277,N_14760,N_14786);
nor UO_278 (O_278,N_14930,N_14835);
nor UO_279 (O_279,N_14798,N_14753);
and UO_280 (O_280,N_14888,N_14809);
and UO_281 (O_281,N_14724,N_14754);
nor UO_282 (O_282,N_14817,N_14771);
and UO_283 (O_283,N_14748,N_14724);
xor UO_284 (O_284,N_14711,N_14963);
xnor UO_285 (O_285,N_14709,N_14759);
or UO_286 (O_286,N_14764,N_14797);
and UO_287 (O_287,N_14833,N_14988);
nand UO_288 (O_288,N_14843,N_14710);
nand UO_289 (O_289,N_14828,N_14920);
xnor UO_290 (O_290,N_14770,N_14857);
xor UO_291 (O_291,N_14883,N_14860);
or UO_292 (O_292,N_14855,N_14805);
or UO_293 (O_293,N_14772,N_14813);
nor UO_294 (O_294,N_14714,N_14924);
and UO_295 (O_295,N_14824,N_14866);
nand UO_296 (O_296,N_14999,N_14724);
nor UO_297 (O_297,N_14955,N_14983);
xor UO_298 (O_298,N_14979,N_14702);
xor UO_299 (O_299,N_14786,N_14824);
or UO_300 (O_300,N_14800,N_14916);
or UO_301 (O_301,N_14941,N_14964);
or UO_302 (O_302,N_14728,N_14934);
nor UO_303 (O_303,N_14767,N_14927);
nand UO_304 (O_304,N_14738,N_14792);
nor UO_305 (O_305,N_14833,N_14733);
xor UO_306 (O_306,N_14830,N_14806);
or UO_307 (O_307,N_14762,N_14945);
or UO_308 (O_308,N_14879,N_14959);
nor UO_309 (O_309,N_14907,N_14969);
or UO_310 (O_310,N_14958,N_14998);
xnor UO_311 (O_311,N_14742,N_14980);
nor UO_312 (O_312,N_14745,N_14784);
xor UO_313 (O_313,N_14706,N_14849);
nor UO_314 (O_314,N_14812,N_14764);
xor UO_315 (O_315,N_14878,N_14874);
xnor UO_316 (O_316,N_14798,N_14872);
nor UO_317 (O_317,N_14895,N_14990);
nor UO_318 (O_318,N_14746,N_14917);
xor UO_319 (O_319,N_14712,N_14904);
nand UO_320 (O_320,N_14764,N_14776);
and UO_321 (O_321,N_14798,N_14882);
nor UO_322 (O_322,N_14815,N_14876);
and UO_323 (O_323,N_14902,N_14890);
nand UO_324 (O_324,N_14738,N_14894);
xnor UO_325 (O_325,N_14987,N_14764);
or UO_326 (O_326,N_14961,N_14829);
and UO_327 (O_327,N_14980,N_14724);
nand UO_328 (O_328,N_14855,N_14949);
xnor UO_329 (O_329,N_14953,N_14864);
nand UO_330 (O_330,N_14775,N_14983);
nor UO_331 (O_331,N_14928,N_14833);
nand UO_332 (O_332,N_14916,N_14747);
xor UO_333 (O_333,N_14880,N_14875);
nor UO_334 (O_334,N_14709,N_14952);
or UO_335 (O_335,N_14705,N_14851);
nand UO_336 (O_336,N_14960,N_14726);
xnor UO_337 (O_337,N_14865,N_14828);
xor UO_338 (O_338,N_14812,N_14935);
and UO_339 (O_339,N_14879,N_14829);
nand UO_340 (O_340,N_14782,N_14821);
xor UO_341 (O_341,N_14763,N_14752);
nand UO_342 (O_342,N_14838,N_14712);
or UO_343 (O_343,N_14999,N_14760);
or UO_344 (O_344,N_14801,N_14898);
or UO_345 (O_345,N_14901,N_14763);
nand UO_346 (O_346,N_14986,N_14991);
and UO_347 (O_347,N_14884,N_14721);
or UO_348 (O_348,N_14718,N_14708);
and UO_349 (O_349,N_14704,N_14996);
nor UO_350 (O_350,N_14780,N_14963);
and UO_351 (O_351,N_14758,N_14916);
and UO_352 (O_352,N_14785,N_14944);
xor UO_353 (O_353,N_14974,N_14841);
xnor UO_354 (O_354,N_14784,N_14823);
or UO_355 (O_355,N_14720,N_14981);
and UO_356 (O_356,N_14963,N_14761);
and UO_357 (O_357,N_14901,N_14932);
xnor UO_358 (O_358,N_14939,N_14927);
xnor UO_359 (O_359,N_14730,N_14909);
nand UO_360 (O_360,N_14736,N_14929);
nand UO_361 (O_361,N_14746,N_14928);
nor UO_362 (O_362,N_14888,N_14812);
nor UO_363 (O_363,N_14868,N_14916);
or UO_364 (O_364,N_14953,N_14705);
nor UO_365 (O_365,N_14784,N_14706);
nor UO_366 (O_366,N_14736,N_14883);
nand UO_367 (O_367,N_14963,N_14703);
nand UO_368 (O_368,N_14896,N_14805);
xnor UO_369 (O_369,N_14808,N_14985);
and UO_370 (O_370,N_14914,N_14722);
nand UO_371 (O_371,N_14710,N_14866);
nand UO_372 (O_372,N_14876,N_14810);
nand UO_373 (O_373,N_14927,N_14740);
nor UO_374 (O_374,N_14759,N_14882);
and UO_375 (O_375,N_14871,N_14855);
and UO_376 (O_376,N_14742,N_14788);
nand UO_377 (O_377,N_14748,N_14810);
xor UO_378 (O_378,N_14893,N_14843);
and UO_379 (O_379,N_14717,N_14736);
nor UO_380 (O_380,N_14948,N_14932);
nand UO_381 (O_381,N_14709,N_14873);
nand UO_382 (O_382,N_14807,N_14802);
xnor UO_383 (O_383,N_14827,N_14864);
and UO_384 (O_384,N_14984,N_14962);
nor UO_385 (O_385,N_14914,N_14899);
nor UO_386 (O_386,N_14785,N_14771);
or UO_387 (O_387,N_14908,N_14954);
xor UO_388 (O_388,N_14802,N_14822);
nor UO_389 (O_389,N_14866,N_14962);
nand UO_390 (O_390,N_14899,N_14748);
or UO_391 (O_391,N_14909,N_14775);
and UO_392 (O_392,N_14734,N_14796);
or UO_393 (O_393,N_14887,N_14718);
and UO_394 (O_394,N_14954,N_14789);
or UO_395 (O_395,N_14844,N_14796);
and UO_396 (O_396,N_14844,N_14708);
xor UO_397 (O_397,N_14774,N_14912);
or UO_398 (O_398,N_14755,N_14949);
and UO_399 (O_399,N_14961,N_14771);
xor UO_400 (O_400,N_14801,N_14807);
and UO_401 (O_401,N_14950,N_14761);
nand UO_402 (O_402,N_14987,N_14865);
nor UO_403 (O_403,N_14717,N_14799);
nand UO_404 (O_404,N_14896,N_14949);
or UO_405 (O_405,N_14929,N_14981);
and UO_406 (O_406,N_14821,N_14767);
nor UO_407 (O_407,N_14852,N_14702);
xnor UO_408 (O_408,N_14836,N_14700);
and UO_409 (O_409,N_14748,N_14884);
nor UO_410 (O_410,N_14990,N_14796);
nand UO_411 (O_411,N_14772,N_14886);
nor UO_412 (O_412,N_14984,N_14795);
and UO_413 (O_413,N_14729,N_14831);
xor UO_414 (O_414,N_14751,N_14829);
and UO_415 (O_415,N_14852,N_14949);
or UO_416 (O_416,N_14882,N_14876);
nand UO_417 (O_417,N_14745,N_14902);
nor UO_418 (O_418,N_14993,N_14761);
and UO_419 (O_419,N_14915,N_14983);
or UO_420 (O_420,N_14884,N_14954);
nand UO_421 (O_421,N_14781,N_14963);
or UO_422 (O_422,N_14869,N_14789);
xor UO_423 (O_423,N_14801,N_14909);
or UO_424 (O_424,N_14876,N_14931);
nor UO_425 (O_425,N_14820,N_14947);
nor UO_426 (O_426,N_14703,N_14899);
and UO_427 (O_427,N_14791,N_14984);
nor UO_428 (O_428,N_14827,N_14801);
or UO_429 (O_429,N_14998,N_14863);
nor UO_430 (O_430,N_14935,N_14706);
and UO_431 (O_431,N_14700,N_14883);
or UO_432 (O_432,N_14779,N_14937);
or UO_433 (O_433,N_14798,N_14915);
and UO_434 (O_434,N_14984,N_14817);
nor UO_435 (O_435,N_14769,N_14959);
and UO_436 (O_436,N_14719,N_14862);
and UO_437 (O_437,N_14795,N_14895);
nor UO_438 (O_438,N_14831,N_14896);
xnor UO_439 (O_439,N_14726,N_14715);
and UO_440 (O_440,N_14717,N_14719);
and UO_441 (O_441,N_14860,N_14713);
and UO_442 (O_442,N_14817,N_14861);
xor UO_443 (O_443,N_14811,N_14808);
nand UO_444 (O_444,N_14868,N_14774);
and UO_445 (O_445,N_14744,N_14906);
nand UO_446 (O_446,N_14952,N_14755);
and UO_447 (O_447,N_14725,N_14832);
nor UO_448 (O_448,N_14983,N_14859);
nand UO_449 (O_449,N_14945,N_14896);
nor UO_450 (O_450,N_14899,N_14872);
nand UO_451 (O_451,N_14967,N_14702);
or UO_452 (O_452,N_14965,N_14758);
xnor UO_453 (O_453,N_14811,N_14967);
or UO_454 (O_454,N_14839,N_14935);
and UO_455 (O_455,N_14868,N_14949);
nor UO_456 (O_456,N_14788,N_14759);
nand UO_457 (O_457,N_14813,N_14880);
and UO_458 (O_458,N_14826,N_14722);
xor UO_459 (O_459,N_14878,N_14711);
nor UO_460 (O_460,N_14742,N_14941);
xnor UO_461 (O_461,N_14815,N_14933);
and UO_462 (O_462,N_14876,N_14716);
xnor UO_463 (O_463,N_14994,N_14985);
xnor UO_464 (O_464,N_14911,N_14841);
nor UO_465 (O_465,N_14897,N_14753);
xnor UO_466 (O_466,N_14848,N_14892);
xnor UO_467 (O_467,N_14758,N_14933);
or UO_468 (O_468,N_14736,N_14845);
or UO_469 (O_469,N_14734,N_14744);
nand UO_470 (O_470,N_14727,N_14895);
or UO_471 (O_471,N_14717,N_14961);
or UO_472 (O_472,N_14855,N_14884);
nor UO_473 (O_473,N_14835,N_14796);
xor UO_474 (O_474,N_14924,N_14759);
and UO_475 (O_475,N_14852,N_14975);
nor UO_476 (O_476,N_14701,N_14902);
nor UO_477 (O_477,N_14802,N_14759);
and UO_478 (O_478,N_14936,N_14999);
or UO_479 (O_479,N_14860,N_14972);
xnor UO_480 (O_480,N_14830,N_14812);
or UO_481 (O_481,N_14780,N_14810);
nor UO_482 (O_482,N_14834,N_14706);
nand UO_483 (O_483,N_14858,N_14922);
nand UO_484 (O_484,N_14865,N_14798);
nand UO_485 (O_485,N_14735,N_14818);
nor UO_486 (O_486,N_14751,N_14714);
xnor UO_487 (O_487,N_14837,N_14790);
nor UO_488 (O_488,N_14925,N_14704);
xor UO_489 (O_489,N_14812,N_14846);
nor UO_490 (O_490,N_14958,N_14726);
and UO_491 (O_491,N_14744,N_14844);
or UO_492 (O_492,N_14879,N_14869);
and UO_493 (O_493,N_14919,N_14898);
or UO_494 (O_494,N_14999,N_14891);
or UO_495 (O_495,N_14858,N_14868);
xor UO_496 (O_496,N_14731,N_14972);
nand UO_497 (O_497,N_14891,N_14982);
nand UO_498 (O_498,N_14917,N_14729);
or UO_499 (O_499,N_14740,N_14911);
xnor UO_500 (O_500,N_14824,N_14834);
and UO_501 (O_501,N_14981,N_14951);
xnor UO_502 (O_502,N_14729,N_14748);
and UO_503 (O_503,N_14943,N_14758);
xor UO_504 (O_504,N_14797,N_14991);
nand UO_505 (O_505,N_14788,N_14767);
nor UO_506 (O_506,N_14959,N_14873);
xnor UO_507 (O_507,N_14899,N_14909);
nand UO_508 (O_508,N_14835,N_14942);
and UO_509 (O_509,N_14753,N_14863);
or UO_510 (O_510,N_14862,N_14922);
nand UO_511 (O_511,N_14766,N_14737);
and UO_512 (O_512,N_14857,N_14772);
nand UO_513 (O_513,N_14756,N_14873);
nand UO_514 (O_514,N_14781,N_14753);
xor UO_515 (O_515,N_14797,N_14958);
nor UO_516 (O_516,N_14755,N_14802);
and UO_517 (O_517,N_14780,N_14724);
nor UO_518 (O_518,N_14982,N_14857);
nor UO_519 (O_519,N_14851,N_14771);
nand UO_520 (O_520,N_14905,N_14904);
xor UO_521 (O_521,N_14725,N_14779);
or UO_522 (O_522,N_14917,N_14879);
and UO_523 (O_523,N_14750,N_14756);
nand UO_524 (O_524,N_14798,N_14749);
or UO_525 (O_525,N_14934,N_14770);
xor UO_526 (O_526,N_14733,N_14872);
xor UO_527 (O_527,N_14962,N_14821);
or UO_528 (O_528,N_14948,N_14865);
nand UO_529 (O_529,N_14987,N_14800);
xor UO_530 (O_530,N_14778,N_14947);
xor UO_531 (O_531,N_14757,N_14911);
xnor UO_532 (O_532,N_14862,N_14792);
and UO_533 (O_533,N_14838,N_14749);
and UO_534 (O_534,N_14739,N_14770);
nand UO_535 (O_535,N_14896,N_14855);
nand UO_536 (O_536,N_14843,N_14859);
nand UO_537 (O_537,N_14848,N_14824);
nand UO_538 (O_538,N_14901,N_14974);
nand UO_539 (O_539,N_14882,N_14778);
xnor UO_540 (O_540,N_14931,N_14906);
and UO_541 (O_541,N_14849,N_14709);
nand UO_542 (O_542,N_14784,N_14996);
and UO_543 (O_543,N_14814,N_14788);
nand UO_544 (O_544,N_14953,N_14959);
or UO_545 (O_545,N_14924,N_14889);
or UO_546 (O_546,N_14834,N_14843);
nor UO_547 (O_547,N_14949,N_14874);
xor UO_548 (O_548,N_14962,N_14773);
nor UO_549 (O_549,N_14814,N_14911);
or UO_550 (O_550,N_14829,N_14902);
or UO_551 (O_551,N_14893,N_14894);
nand UO_552 (O_552,N_14836,N_14893);
nand UO_553 (O_553,N_14770,N_14898);
nand UO_554 (O_554,N_14750,N_14871);
nor UO_555 (O_555,N_14861,N_14725);
and UO_556 (O_556,N_14869,N_14947);
xor UO_557 (O_557,N_14750,N_14880);
or UO_558 (O_558,N_14841,N_14814);
nor UO_559 (O_559,N_14878,N_14969);
xnor UO_560 (O_560,N_14758,N_14947);
and UO_561 (O_561,N_14779,N_14974);
and UO_562 (O_562,N_14903,N_14839);
xor UO_563 (O_563,N_14991,N_14883);
nor UO_564 (O_564,N_14908,N_14723);
or UO_565 (O_565,N_14957,N_14723);
nor UO_566 (O_566,N_14742,N_14924);
nor UO_567 (O_567,N_14992,N_14712);
xor UO_568 (O_568,N_14802,N_14907);
or UO_569 (O_569,N_14933,N_14740);
nand UO_570 (O_570,N_14996,N_14975);
or UO_571 (O_571,N_14929,N_14899);
and UO_572 (O_572,N_14952,N_14941);
or UO_573 (O_573,N_14978,N_14953);
and UO_574 (O_574,N_14892,N_14822);
nor UO_575 (O_575,N_14813,N_14819);
nor UO_576 (O_576,N_14790,N_14723);
xnor UO_577 (O_577,N_14738,N_14872);
and UO_578 (O_578,N_14908,N_14787);
nand UO_579 (O_579,N_14912,N_14883);
xnor UO_580 (O_580,N_14726,N_14984);
or UO_581 (O_581,N_14787,N_14914);
xor UO_582 (O_582,N_14900,N_14863);
or UO_583 (O_583,N_14990,N_14799);
or UO_584 (O_584,N_14760,N_14931);
nor UO_585 (O_585,N_14956,N_14739);
or UO_586 (O_586,N_14740,N_14822);
nand UO_587 (O_587,N_14727,N_14742);
and UO_588 (O_588,N_14714,N_14834);
nand UO_589 (O_589,N_14797,N_14741);
nand UO_590 (O_590,N_14802,N_14858);
nor UO_591 (O_591,N_14928,N_14834);
nand UO_592 (O_592,N_14797,N_14928);
nor UO_593 (O_593,N_14820,N_14991);
nand UO_594 (O_594,N_14778,N_14981);
xor UO_595 (O_595,N_14929,N_14795);
nand UO_596 (O_596,N_14835,N_14875);
or UO_597 (O_597,N_14744,N_14984);
or UO_598 (O_598,N_14889,N_14939);
xnor UO_599 (O_599,N_14722,N_14739);
and UO_600 (O_600,N_14723,N_14911);
nand UO_601 (O_601,N_14750,N_14810);
xor UO_602 (O_602,N_14929,N_14749);
or UO_603 (O_603,N_14780,N_14935);
xnor UO_604 (O_604,N_14784,N_14849);
nor UO_605 (O_605,N_14892,N_14722);
and UO_606 (O_606,N_14782,N_14866);
xnor UO_607 (O_607,N_14718,N_14970);
and UO_608 (O_608,N_14766,N_14885);
nand UO_609 (O_609,N_14961,N_14820);
nand UO_610 (O_610,N_14808,N_14930);
xnor UO_611 (O_611,N_14846,N_14717);
nand UO_612 (O_612,N_14924,N_14743);
and UO_613 (O_613,N_14995,N_14973);
and UO_614 (O_614,N_14795,N_14911);
xor UO_615 (O_615,N_14744,N_14784);
and UO_616 (O_616,N_14797,N_14892);
or UO_617 (O_617,N_14832,N_14933);
xor UO_618 (O_618,N_14888,N_14808);
or UO_619 (O_619,N_14762,N_14839);
nor UO_620 (O_620,N_14869,N_14759);
xor UO_621 (O_621,N_14969,N_14894);
or UO_622 (O_622,N_14949,N_14780);
xor UO_623 (O_623,N_14753,N_14735);
or UO_624 (O_624,N_14844,N_14775);
and UO_625 (O_625,N_14722,N_14969);
and UO_626 (O_626,N_14832,N_14891);
xor UO_627 (O_627,N_14956,N_14939);
and UO_628 (O_628,N_14964,N_14895);
or UO_629 (O_629,N_14975,N_14838);
nor UO_630 (O_630,N_14736,N_14935);
and UO_631 (O_631,N_14761,N_14720);
xor UO_632 (O_632,N_14717,N_14952);
nand UO_633 (O_633,N_14785,N_14972);
and UO_634 (O_634,N_14956,N_14945);
xor UO_635 (O_635,N_14770,N_14711);
and UO_636 (O_636,N_14886,N_14754);
and UO_637 (O_637,N_14962,N_14899);
nor UO_638 (O_638,N_14908,N_14920);
nor UO_639 (O_639,N_14859,N_14917);
nand UO_640 (O_640,N_14798,N_14919);
nand UO_641 (O_641,N_14885,N_14950);
and UO_642 (O_642,N_14974,N_14845);
and UO_643 (O_643,N_14825,N_14985);
and UO_644 (O_644,N_14734,N_14851);
xor UO_645 (O_645,N_14884,N_14706);
nand UO_646 (O_646,N_14922,N_14888);
nor UO_647 (O_647,N_14762,N_14972);
nand UO_648 (O_648,N_14761,N_14744);
xor UO_649 (O_649,N_14947,N_14999);
xnor UO_650 (O_650,N_14769,N_14981);
nand UO_651 (O_651,N_14934,N_14715);
nor UO_652 (O_652,N_14837,N_14985);
or UO_653 (O_653,N_14880,N_14978);
nand UO_654 (O_654,N_14764,N_14843);
nand UO_655 (O_655,N_14936,N_14910);
xnor UO_656 (O_656,N_14769,N_14823);
xor UO_657 (O_657,N_14904,N_14812);
xnor UO_658 (O_658,N_14735,N_14702);
nand UO_659 (O_659,N_14918,N_14830);
and UO_660 (O_660,N_14710,N_14790);
nor UO_661 (O_661,N_14744,N_14896);
or UO_662 (O_662,N_14961,N_14980);
and UO_663 (O_663,N_14899,N_14815);
nor UO_664 (O_664,N_14944,N_14772);
nor UO_665 (O_665,N_14777,N_14844);
nor UO_666 (O_666,N_14733,N_14785);
and UO_667 (O_667,N_14821,N_14931);
and UO_668 (O_668,N_14938,N_14788);
or UO_669 (O_669,N_14908,N_14876);
nand UO_670 (O_670,N_14967,N_14884);
or UO_671 (O_671,N_14727,N_14718);
xor UO_672 (O_672,N_14708,N_14782);
nand UO_673 (O_673,N_14765,N_14842);
nor UO_674 (O_674,N_14741,N_14772);
or UO_675 (O_675,N_14803,N_14963);
nor UO_676 (O_676,N_14815,N_14705);
or UO_677 (O_677,N_14992,N_14983);
nor UO_678 (O_678,N_14751,N_14892);
and UO_679 (O_679,N_14928,N_14735);
nand UO_680 (O_680,N_14877,N_14904);
or UO_681 (O_681,N_14981,N_14785);
xor UO_682 (O_682,N_14931,N_14714);
and UO_683 (O_683,N_14862,N_14728);
nor UO_684 (O_684,N_14868,N_14888);
nor UO_685 (O_685,N_14921,N_14707);
nor UO_686 (O_686,N_14949,N_14823);
xor UO_687 (O_687,N_14916,N_14755);
nor UO_688 (O_688,N_14804,N_14917);
nand UO_689 (O_689,N_14795,N_14726);
xnor UO_690 (O_690,N_14861,N_14915);
or UO_691 (O_691,N_14946,N_14955);
and UO_692 (O_692,N_14747,N_14711);
or UO_693 (O_693,N_14796,N_14887);
nor UO_694 (O_694,N_14782,N_14767);
nand UO_695 (O_695,N_14908,N_14770);
nor UO_696 (O_696,N_14998,N_14876);
or UO_697 (O_697,N_14849,N_14931);
xnor UO_698 (O_698,N_14847,N_14996);
nand UO_699 (O_699,N_14708,N_14880);
and UO_700 (O_700,N_14790,N_14796);
xor UO_701 (O_701,N_14825,N_14741);
xor UO_702 (O_702,N_14721,N_14791);
and UO_703 (O_703,N_14900,N_14823);
nor UO_704 (O_704,N_14881,N_14997);
nand UO_705 (O_705,N_14876,N_14827);
or UO_706 (O_706,N_14758,N_14966);
and UO_707 (O_707,N_14855,N_14833);
nor UO_708 (O_708,N_14888,N_14776);
and UO_709 (O_709,N_14874,N_14830);
xor UO_710 (O_710,N_14802,N_14971);
and UO_711 (O_711,N_14776,N_14737);
and UO_712 (O_712,N_14741,N_14838);
nand UO_713 (O_713,N_14921,N_14998);
xor UO_714 (O_714,N_14766,N_14714);
and UO_715 (O_715,N_14841,N_14946);
xor UO_716 (O_716,N_14888,N_14910);
nand UO_717 (O_717,N_14862,N_14775);
nor UO_718 (O_718,N_14976,N_14962);
nand UO_719 (O_719,N_14985,N_14919);
nor UO_720 (O_720,N_14886,N_14716);
xnor UO_721 (O_721,N_14760,N_14960);
nand UO_722 (O_722,N_14926,N_14943);
or UO_723 (O_723,N_14701,N_14825);
nand UO_724 (O_724,N_14921,N_14904);
and UO_725 (O_725,N_14928,N_14814);
nand UO_726 (O_726,N_14838,N_14871);
or UO_727 (O_727,N_14926,N_14923);
or UO_728 (O_728,N_14995,N_14855);
nor UO_729 (O_729,N_14912,N_14963);
or UO_730 (O_730,N_14820,N_14976);
and UO_731 (O_731,N_14831,N_14862);
and UO_732 (O_732,N_14886,N_14863);
nand UO_733 (O_733,N_14744,N_14926);
nor UO_734 (O_734,N_14767,N_14963);
or UO_735 (O_735,N_14987,N_14744);
nor UO_736 (O_736,N_14915,N_14739);
xnor UO_737 (O_737,N_14936,N_14809);
xor UO_738 (O_738,N_14920,N_14710);
xor UO_739 (O_739,N_14782,N_14812);
nand UO_740 (O_740,N_14788,N_14879);
or UO_741 (O_741,N_14834,N_14862);
nor UO_742 (O_742,N_14897,N_14960);
nand UO_743 (O_743,N_14793,N_14947);
and UO_744 (O_744,N_14809,N_14704);
nand UO_745 (O_745,N_14977,N_14825);
nand UO_746 (O_746,N_14951,N_14716);
or UO_747 (O_747,N_14733,N_14887);
or UO_748 (O_748,N_14753,N_14921);
or UO_749 (O_749,N_14777,N_14996);
nor UO_750 (O_750,N_14880,N_14736);
xor UO_751 (O_751,N_14730,N_14979);
nor UO_752 (O_752,N_14729,N_14939);
nor UO_753 (O_753,N_14970,N_14806);
or UO_754 (O_754,N_14946,N_14732);
and UO_755 (O_755,N_14939,N_14792);
nor UO_756 (O_756,N_14818,N_14723);
or UO_757 (O_757,N_14989,N_14857);
and UO_758 (O_758,N_14936,N_14976);
nor UO_759 (O_759,N_14884,N_14784);
nand UO_760 (O_760,N_14980,N_14719);
nand UO_761 (O_761,N_14812,N_14820);
or UO_762 (O_762,N_14726,N_14810);
and UO_763 (O_763,N_14767,N_14893);
and UO_764 (O_764,N_14981,N_14975);
xnor UO_765 (O_765,N_14916,N_14974);
nor UO_766 (O_766,N_14987,N_14782);
xnor UO_767 (O_767,N_14821,N_14784);
xor UO_768 (O_768,N_14801,N_14858);
or UO_769 (O_769,N_14769,N_14915);
nand UO_770 (O_770,N_14801,N_14784);
nand UO_771 (O_771,N_14749,N_14894);
or UO_772 (O_772,N_14997,N_14956);
xor UO_773 (O_773,N_14972,N_14936);
nand UO_774 (O_774,N_14760,N_14891);
nand UO_775 (O_775,N_14768,N_14929);
nor UO_776 (O_776,N_14935,N_14815);
nor UO_777 (O_777,N_14946,N_14718);
and UO_778 (O_778,N_14708,N_14854);
nand UO_779 (O_779,N_14728,N_14860);
and UO_780 (O_780,N_14955,N_14785);
and UO_781 (O_781,N_14982,N_14822);
and UO_782 (O_782,N_14712,N_14906);
nor UO_783 (O_783,N_14982,N_14867);
nor UO_784 (O_784,N_14880,N_14999);
and UO_785 (O_785,N_14936,N_14909);
and UO_786 (O_786,N_14977,N_14863);
or UO_787 (O_787,N_14957,N_14856);
or UO_788 (O_788,N_14902,N_14806);
xor UO_789 (O_789,N_14754,N_14835);
xor UO_790 (O_790,N_14901,N_14803);
and UO_791 (O_791,N_14770,N_14920);
xnor UO_792 (O_792,N_14727,N_14918);
or UO_793 (O_793,N_14757,N_14792);
nand UO_794 (O_794,N_14951,N_14800);
and UO_795 (O_795,N_14834,N_14880);
xor UO_796 (O_796,N_14839,N_14742);
nand UO_797 (O_797,N_14835,N_14713);
xnor UO_798 (O_798,N_14763,N_14948);
and UO_799 (O_799,N_14923,N_14891);
xor UO_800 (O_800,N_14921,N_14825);
nor UO_801 (O_801,N_14757,N_14717);
or UO_802 (O_802,N_14780,N_14758);
or UO_803 (O_803,N_14894,N_14936);
and UO_804 (O_804,N_14781,N_14986);
nor UO_805 (O_805,N_14810,N_14861);
and UO_806 (O_806,N_14912,N_14951);
nor UO_807 (O_807,N_14742,N_14976);
xor UO_808 (O_808,N_14994,N_14983);
nand UO_809 (O_809,N_14930,N_14726);
or UO_810 (O_810,N_14715,N_14836);
nor UO_811 (O_811,N_14733,N_14894);
nor UO_812 (O_812,N_14909,N_14997);
and UO_813 (O_813,N_14770,N_14950);
and UO_814 (O_814,N_14845,N_14821);
xnor UO_815 (O_815,N_14851,N_14935);
or UO_816 (O_816,N_14964,N_14816);
or UO_817 (O_817,N_14764,N_14980);
or UO_818 (O_818,N_14948,N_14735);
xor UO_819 (O_819,N_14721,N_14758);
nor UO_820 (O_820,N_14727,N_14856);
nand UO_821 (O_821,N_14711,N_14826);
or UO_822 (O_822,N_14706,N_14970);
and UO_823 (O_823,N_14770,N_14811);
xor UO_824 (O_824,N_14841,N_14742);
and UO_825 (O_825,N_14877,N_14977);
xnor UO_826 (O_826,N_14716,N_14789);
nand UO_827 (O_827,N_14994,N_14750);
xor UO_828 (O_828,N_14829,N_14720);
or UO_829 (O_829,N_14808,N_14921);
xnor UO_830 (O_830,N_14793,N_14851);
xor UO_831 (O_831,N_14736,N_14755);
nand UO_832 (O_832,N_14779,N_14875);
and UO_833 (O_833,N_14709,N_14749);
or UO_834 (O_834,N_14863,N_14896);
xnor UO_835 (O_835,N_14987,N_14980);
nand UO_836 (O_836,N_14989,N_14862);
or UO_837 (O_837,N_14804,N_14745);
xor UO_838 (O_838,N_14873,N_14871);
nand UO_839 (O_839,N_14965,N_14954);
nand UO_840 (O_840,N_14871,N_14734);
nand UO_841 (O_841,N_14849,N_14923);
xnor UO_842 (O_842,N_14949,N_14828);
and UO_843 (O_843,N_14713,N_14775);
and UO_844 (O_844,N_14987,N_14991);
and UO_845 (O_845,N_14979,N_14981);
nor UO_846 (O_846,N_14821,N_14961);
and UO_847 (O_847,N_14999,N_14754);
nor UO_848 (O_848,N_14883,N_14951);
nor UO_849 (O_849,N_14740,N_14759);
xnor UO_850 (O_850,N_14889,N_14967);
or UO_851 (O_851,N_14715,N_14811);
xor UO_852 (O_852,N_14808,N_14724);
or UO_853 (O_853,N_14716,N_14819);
nand UO_854 (O_854,N_14795,N_14782);
and UO_855 (O_855,N_14778,N_14878);
or UO_856 (O_856,N_14908,N_14766);
nor UO_857 (O_857,N_14755,N_14862);
nand UO_858 (O_858,N_14708,N_14853);
and UO_859 (O_859,N_14786,N_14722);
or UO_860 (O_860,N_14707,N_14767);
xnor UO_861 (O_861,N_14781,N_14819);
nand UO_862 (O_862,N_14861,N_14980);
nor UO_863 (O_863,N_14739,N_14714);
xnor UO_864 (O_864,N_14827,N_14906);
and UO_865 (O_865,N_14819,N_14880);
xnor UO_866 (O_866,N_14720,N_14944);
or UO_867 (O_867,N_14870,N_14791);
xnor UO_868 (O_868,N_14859,N_14787);
nor UO_869 (O_869,N_14762,N_14907);
or UO_870 (O_870,N_14928,N_14740);
and UO_871 (O_871,N_14776,N_14894);
or UO_872 (O_872,N_14752,N_14725);
nand UO_873 (O_873,N_14760,N_14899);
and UO_874 (O_874,N_14985,N_14971);
nand UO_875 (O_875,N_14848,N_14913);
and UO_876 (O_876,N_14887,N_14839);
nor UO_877 (O_877,N_14919,N_14991);
and UO_878 (O_878,N_14840,N_14897);
or UO_879 (O_879,N_14709,N_14965);
nor UO_880 (O_880,N_14915,N_14927);
nand UO_881 (O_881,N_14967,N_14943);
and UO_882 (O_882,N_14715,N_14970);
nor UO_883 (O_883,N_14846,N_14963);
or UO_884 (O_884,N_14704,N_14860);
or UO_885 (O_885,N_14705,N_14703);
xnor UO_886 (O_886,N_14940,N_14994);
xor UO_887 (O_887,N_14832,N_14823);
xor UO_888 (O_888,N_14715,N_14929);
or UO_889 (O_889,N_14975,N_14773);
nand UO_890 (O_890,N_14875,N_14987);
and UO_891 (O_891,N_14769,N_14899);
xnor UO_892 (O_892,N_14739,N_14911);
and UO_893 (O_893,N_14808,N_14816);
and UO_894 (O_894,N_14750,N_14729);
nand UO_895 (O_895,N_14925,N_14838);
nand UO_896 (O_896,N_14814,N_14966);
xnor UO_897 (O_897,N_14717,N_14776);
and UO_898 (O_898,N_14837,N_14918);
and UO_899 (O_899,N_14765,N_14786);
or UO_900 (O_900,N_14802,N_14713);
and UO_901 (O_901,N_14918,N_14805);
nand UO_902 (O_902,N_14884,N_14819);
nand UO_903 (O_903,N_14713,N_14942);
and UO_904 (O_904,N_14846,N_14713);
or UO_905 (O_905,N_14936,N_14806);
xnor UO_906 (O_906,N_14874,N_14864);
nand UO_907 (O_907,N_14805,N_14857);
nand UO_908 (O_908,N_14878,N_14721);
and UO_909 (O_909,N_14928,N_14855);
or UO_910 (O_910,N_14994,N_14919);
or UO_911 (O_911,N_14737,N_14942);
nor UO_912 (O_912,N_14893,N_14782);
nand UO_913 (O_913,N_14983,N_14707);
nor UO_914 (O_914,N_14922,N_14992);
xnor UO_915 (O_915,N_14950,N_14793);
nor UO_916 (O_916,N_14832,N_14934);
nand UO_917 (O_917,N_14798,N_14789);
xor UO_918 (O_918,N_14908,N_14732);
or UO_919 (O_919,N_14941,N_14928);
xor UO_920 (O_920,N_14765,N_14837);
and UO_921 (O_921,N_14810,N_14874);
and UO_922 (O_922,N_14965,N_14820);
or UO_923 (O_923,N_14935,N_14782);
xor UO_924 (O_924,N_14860,N_14823);
xnor UO_925 (O_925,N_14917,N_14733);
xor UO_926 (O_926,N_14970,N_14724);
or UO_927 (O_927,N_14805,N_14910);
or UO_928 (O_928,N_14940,N_14972);
nand UO_929 (O_929,N_14760,N_14894);
or UO_930 (O_930,N_14918,N_14750);
or UO_931 (O_931,N_14940,N_14999);
nand UO_932 (O_932,N_14852,N_14750);
nand UO_933 (O_933,N_14937,N_14885);
and UO_934 (O_934,N_14792,N_14962);
and UO_935 (O_935,N_14865,N_14796);
or UO_936 (O_936,N_14895,N_14735);
xnor UO_937 (O_937,N_14919,N_14997);
xnor UO_938 (O_938,N_14943,N_14980);
or UO_939 (O_939,N_14901,N_14893);
xnor UO_940 (O_940,N_14881,N_14835);
xnor UO_941 (O_941,N_14987,N_14855);
nor UO_942 (O_942,N_14741,N_14929);
or UO_943 (O_943,N_14885,N_14859);
nor UO_944 (O_944,N_14912,N_14906);
nand UO_945 (O_945,N_14988,N_14706);
xnor UO_946 (O_946,N_14950,N_14816);
and UO_947 (O_947,N_14806,N_14916);
and UO_948 (O_948,N_14958,N_14828);
or UO_949 (O_949,N_14729,N_14926);
or UO_950 (O_950,N_14816,N_14747);
xnor UO_951 (O_951,N_14728,N_14954);
and UO_952 (O_952,N_14917,N_14961);
nor UO_953 (O_953,N_14892,N_14861);
and UO_954 (O_954,N_14838,N_14886);
and UO_955 (O_955,N_14776,N_14872);
xor UO_956 (O_956,N_14722,N_14749);
nor UO_957 (O_957,N_14808,N_14861);
xor UO_958 (O_958,N_14848,N_14875);
and UO_959 (O_959,N_14705,N_14982);
nand UO_960 (O_960,N_14706,N_14747);
nand UO_961 (O_961,N_14855,N_14941);
or UO_962 (O_962,N_14757,N_14737);
nor UO_963 (O_963,N_14808,N_14729);
nand UO_964 (O_964,N_14981,N_14994);
and UO_965 (O_965,N_14919,N_14776);
and UO_966 (O_966,N_14778,N_14847);
or UO_967 (O_967,N_14896,N_14764);
xor UO_968 (O_968,N_14826,N_14941);
and UO_969 (O_969,N_14970,N_14786);
xnor UO_970 (O_970,N_14807,N_14793);
nor UO_971 (O_971,N_14910,N_14794);
or UO_972 (O_972,N_14866,N_14917);
nand UO_973 (O_973,N_14746,N_14806);
xor UO_974 (O_974,N_14840,N_14744);
nor UO_975 (O_975,N_14962,N_14875);
or UO_976 (O_976,N_14982,N_14710);
xnor UO_977 (O_977,N_14716,N_14752);
nor UO_978 (O_978,N_14845,N_14873);
and UO_979 (O_979,N_14983,N_14735);
nor UO_980 (O_980,N_14965,N_14945);
xnor UO_981 (O_981,N_14852,N_14751);
and UO_982 (O_982,N_14811,N_14898);
and UO_983 (O_983,N_14702,N_14750);
or UO_984 (O_984,N_14874,N_14977);
nand UO_985 (O_985,N_14946,N_14858);
and UO_986 (O_986,N_14866,N_14859);
nand UO_987 (O_987,N_14863,N_14980);
or UO_988 (O_988,N_14781,N_14755);
nor UO_989 (O_989,N_14816,N_14723);
or UO_990 (O_990,N_14950,N_14732);
and UO_991 (O_991,N_14812,N_14864);
nand UO_992 (O_992,N_14711,N_14841);
xnor UO_993 (O_993,N_14874,N_14839);
nand UO_994 (O_994,N_14821,N_14996);
and UO_995 (O_995,N_14768,N_14823);
xor UO_996 (O_996,N_14857,N_14754);
nor UO_997 (O_997,N_14720,N_14940);
nor UO_998 (O_998,N_14793,N_14783);
xor UO_999 (O_999,N_14709,N_14913);
and UO_1000 (O_1000,N_14899,N_14961);
or UO_1001 (O_1001,N_14798,N_14855);
nand UO_1002 (O_1002,N_14949,N_14991);
nand UO_1003 (O_1003,N_14806,N_14880);
nand UO_1004 (O_1004,N_14957,N_14888);
or UO_1005 (O_1005,N_14827,N_14945);
and UO_1006 (O_1006,N_14966,N_14782);
or UO_1007 (O_1007,N_14737,N_14828);
xor UO_1008 (O_1008,N_14914,N_14973);
and UO_1009 (O_1009,N_14778,N_14849);
or UO_1010 (O_1010,N_14784,N_14854);
and UO_1011 (O_1011,N_14973,N_14867);
nand UO_1012 (O_1012,N_14902,N_14848);
nand UO_1013 (O_1013,N_14891,N_14933);
xnor UO_1014 (O_1014,N_14947,N_14774);
xor UO_1015 (O_1015,N_14991,N_14984);
and UO_1016 (O_1016,N_14888,N_14775);
or UO_1017 (O_1017,N_14975,N_14775);
xor UO_1018 (O_1018,N_14811,N_14845);
or UO_1019 (O_1019,N_14954,N_14876);
xor UO_1020 (O_1020,N_14854,N_14787);
and UO_1021 (O_1021,N_14747,N_14918);
nand UO_1022 (O_1022,N_14714,N_14907);
xor UO_1023 (O_1023,N_14938,N_14888);
nand UO_1024 (O_1024,N_14741,N_14906);
and UO_1025 (O_1025,N_14810,N_14901);
nand UO_1026 (O_1026,N_14701,N_14811);
or UO_1027 (O_1027,N_14784,N_14751);
nor UO_1028 (O_1028,N_14837,N_14925);
or UO_1029 (O_1029,N_14860,N_14986);
xnor UO_1030 (O_1030,N_14794,N_14799);
nand UO_1031 (O_1031,N_14832,N_14923);
and UO_1032 (O_1032,N_14744,N_14952);
or UO_1033 (O_1033,N_14969,N_14762);
nand UO_1034 (O_1034,N_14867,N_14836);
or UO_1035 (O_1035,N_14948,N_14999);
nor UO_1036 (O_1036,N_14808,N_14855);
or UO_1037 (O_1037,N_14960,N_14948);
nand UO_1038 (O_1038,N_14765,N_14822);
and UO_1039 (O_1039,N_14883,N_14834);
nor UO_1040 (O_1040,N_14712,N_14746);
and UO_1041 (O_1041,N_14700,N_14869);
or UO_1042 (O_1042,N_14749,N_14700);
or UO_1043 (O_1043,N_14751,N_14831);
or UO_1044 (O_1044,N_14963,N_14918);
nor UO_1045 (O_1045,N_14707,N_14752);
and UO_1046 (O_1046,N_14978,N_14812);
nand UO_1047 (O_1047,N_14750,N_14767);
and UO_1048 (O_1048,N_14985,N_14841);
and UO_1049 (O_1049,N_14950,N_14862);
nor UO_1050 (O_1050,N_14911,N_14990);
nand UO_1051 (O_1051,N_14994,N_14815);
and UO_1052 (O_1052,N_14809,N_14834);
nand UO_1053 (O_1053,N_14854,N_14957);
nor UO_1054 (O_1054,N_14980,N_14766);
and UO_1055 (O_1055,N_14760,N_14920);
and UO_1056 (O_1056,N_14973,N_14947);
and UO_1057 (O_1057,N_14770,N_14769);
nand UO_1058 (O_1058,N_14710,N_14845);
xnor UO_1059 (O_1059,N_14870,N_14776);
or UO_1060 (O_1060,N_14883,N_14952);
nand UO_1061 (O_1061,N_14899,N_14708);
and UO_1062 (O_1062,N_14734,N_14923);
nor UO_1063 (O_1063,N_14789,N_14930);
and UO_1064 (O_1064,N_14770,N_14710);
nand UO_1065 (O_1065,N_14803,N_14935);
xor UO_1066 (O_1066,N_14848,N_14861);
nand UO_1067 (O_1067,N_14721,N_14907);
and UO_1068 (O_1068,N_14836,N_14975);
xor UO_1069 (O_1069,N_14952,N_14847);
xnor UO_1070 (O_1070,N_14932,N_14812);
nor UO_1071 (O_1071,N_14899,N_14968);
nor UO_1072 (O_1072,N_14736,N_14838);
nand UO_1073 (O_1073,N_14751,N_14994);
and UO_1074 (O_1074,N_14736,N_14746);
nand UO_1075 (O_1075,N_14710,N_14798);
nand UO_1076 (O_1076,N_14835,N_14771);
nand UO_1077 (O_1077,N_14848,N_14719);
or UO_1078 (O_1078,N_14963,N_14993);
and UO_1079 (O_1079,N_14864,N_14807);
nor UO_1080 (O_1080,N_14806,N_14757);
or UO_1081 (O_1081,N_14820,N_14952);
and UO_1082 (O_1082,N_14994,N_14972);
nor UO_1083 (O_1083,N_14806,N_14855);
nor UO_1084 (O_1084,N_14808,N_14708);
nor UO_1085 (O_1085,N_14706,N_14728);
nor UO_1086 (O_1086,N_14732,N_14966);
nand UO_1087 (O_1087,N_14791,N_14846);
nand UO_1088 (O_1088,N_14852,N_14900);
nand UO_1089 (O_1089,N_14891,N_14825);
nor UO_1090 (O_1090,N_14978,N_14877);
xor UO_1091 (O_1091,N_14711,N_14996);
or UO_1092 (O_1092,N_14775,N_14943);
and UO_1093 (O_1093,N_14764,N_14732);
xnor UO_1094 (O_1094,N_14905,N_14768);
and UO_1095 (O_1095,N_14708,N_14736);
xnor UO_1096 (O_1096,N_14940,N_14723);
nand UO_1097 (O_1097,N_14746,N_14958);
nand UO_1098 (O_1098,N_14716,N_14705);
nand UO_1099 (O_1099,N_14825,N_14738);
and UO_1100 (O_1100,N_14930,N_14751);
xor UO_1101 (O_1101,N_14770,N_14801);
or UO_1102 (O_1102,N_14887,N_14855);
xnor UO_1103 (O_1103,N_14929,N_14923);
nor UO_1104 (O_1104,N_14739,N_14955);
and UO_1105 (O_1105,N_14700,N_14831);
nand UO_1106 (O_1106,N_14743,N_14925);
nor UO_1107 (O_1107,N_14781,N_14776);
and UO_1108 (O_1108,N_14936,N_14937);
nor UO_1109 (O_1109,N_14899,N_14797);
and UO_1110 (O_1110,N_14807,N_14711);
nand UO_1111 (O_1111,N_14848,N_14934);
nor UO_1112 (O_1112,N_14879,N_14720);
and UO_1113 (O_1113,N_14865,N_14756);
and UO_1114 (O_1114,N_14960,N_14865);
and UO_1115 (O_1115,N_14702,N_14730);
nand UO_1116 (O_1116,N_14743,N_14999);
nand UO_1117 (O_1117,N_14761,N_14836);
or UO_1118 (O_1118,N_14750,N_14967);
and UO_1119 (O_1119,N_14992,N_14716);
and UO_1120 (O_1120,N_14725,N_14926);
and UO_1121 (O_1121,N_14984,N_14873);
nand UO_1122 (O_1122,N_14892,N_14953);
xnor UO_1123 (O_1123,N_14950,N_14714);
and UO_1124 (O_1124,N_14910,N_14938);
or UO_1125 (O_1125,N_14902,N_14907);
nor UO_1126 (O_1126,N_14860,N_14960);
nor UO_1127 (O_1127,N_14884,N_14920);
nand UO_1128 (O_1128,N_14740,N_14887);
and UO_1129 (O_1129,N_14795,N_14746);
and UO_1130 (O_1130,N_14919,N_14995);
or UO_1131 (O_1131,N_14938,N_14790);
nor UO_1132 (O_1132,N_14890,N_14825);
nor UO_1133 (O_1133,N_14715,N_14815);
nor UO_1134 (O_1134,N_14803,N_14833);
and UO_1135 (O_1135,N_14800,N_14768);
and UO_1136 (O_1136,N_14713,N_14827);
and UO_1137 (O_1137,N_14924,N_14973);
or UO_1138 (O_1138,N_14923,N_14930);
nand UO_1139 (O_1139,N_14830,N_14815);
nor UO_1140 (O_1140,N_14915,N_14895);
nor UO_1141 (O_1141,N_14933,N_14767);
xor UO_1142 (O_1142,N_14743,N_14702);
nor UO_1143 (O_1143,N_14736,N_14989);
xnor UO_1144 (O_1144,N_14806,N_14747);
nand UO_1145 (O_1145,N_14862,N_14853);
or UO_1146 (O_1146,N_14726,N_14800);
nand UO_1147 (O_1147,N_14886,N_14986);
nand UO_1148 (O_1148,N_14885,N_14927);
or UO_1149 (O_1149,N_14993,N_14856);
xnor UO_1150 (O_1150,N_14805,N_14820);
xnor UO_1151 (O_1151,N_14993,N_14750);
or UO_1152 (O_1152,N_14857,N_14871);
nand UO_1153 (O_1153,N_14735,N_14921);
and UO_1154 (O_1154,N_14857,N_14994);
nor UO_1155 (O_1155,N_14752,N_14712);
or UO_1156 (O_1156,N_14876,N_14850);
and UO_1157 (O_1157,N_14804,N_14771);
and UO_1158 (O_1158,N_14710,N_14721);
or UO_1159 (O_1159,N_14814,N_14981);
nand UO_1160 (O_1160,N_14913,N_14984);
nand UO_1161 (O_1161,N_14809,N_14815);
nor UO_1162 (O_1162,N_14769,N_14709);
xor UO_1163 (O_1163,N_14900,N_14766);
xor UO_1164 (O_1164,N_14752,N_14985);
and UO_1165 (O_1165,N_14833,N_14871);
or UO_1166 (O_1166,N_14733,N_14929);
and UO_1167 (O_1167,N_14997,N_14759);
or UO_1168 (O_1168,N_14998,N_14952);
nand UO_1169 (O_1169,N_14713,N_14748);
xor UO_1170 (O_1170,N_14816,N_14746);
xor UO_1171 (O_1171,N_14896,N_14875);
xor UO_1172 (O_1172,N_14913,N_14722);
and UO_1173 (O_1173,N_14855,N_14885);
or UO_1174 (O_1174,N_14888,N_14968);
and UO_1175 (O_1175,N_14888,N_14761);
nand UO_1176 (O_1176,N_14883,N_14997);
xor UO_1177 (O_1177,N_14751,N_14722);
and UO_1178 (O_1178,N_14937,N_14755);
nand UO_1179 (O_1179,N_14735,N_14861);
nor UO_1180 (O_1180,N_14987,N_14922);
nor UO_1181 (O_1181,N_14806,N_14705);
nand UO_1182 (O_1182,N_14937,N_14714);
nand UO_1183 (O_1183,N_14906,N_14787);
or UO_1184 (O_1184,N_14736,N_14919);
nor UO_1185 (O_1185,N_14907,N_14847);
and UO_1186 (O_1186,N_14864,N_14726);
and UO_1187 (O_1187,N_14785,N_14901);
nor UO_1188 (O_1188,N_14845,N_14930);
xor UO_1189 (O_1189,N_14732,N_14809);
nor UO_1190 (O_1190,N_14928,N_14781);
or UO_1191 (O_1191,N_14932,N_14778);
nor UO_1192 (O_1192,N_14911,N_14791);
xor UO_1193 (O_1193,N_14759,N_14772);
nand UO_1194 (O_1194,N_14837,N_14927);
nand UO_1195 (O_1195,N_14982,N_14786);
nor UO_1196 (O_1196,N_14797,N_14778);
or UO_1197 (O_1197,N_14844,N_14993);
nand UO_1198 (O_1198,N_14912,N_14814);
and UO_1199 (O_1199,N_14897,N_14902);
nand UO_1200 (O_1200,N_14703,N_14823);
nor UO_1201 (O_1201,N_14815,N_14998);
or UO_1202 (O_1202,N_14880,N_14874);
and UO_1203 (O_1203,N_14976,N_14867);
and UO_1204 (O_1204,N_14871,N_14804);
nor UO_1205 (O_1205,N_14839,N_14909);
and UO_1206 (O_1206,N_14771,N_14930);
or UO_1207 (O_1207,N_14876,N_14700);
nor UO_1208 (O_1208,N_14869,N_14977);
or UO_1209 (O_1209,N_14749,N_14744);
nand UO_1210 (O_1210,N_14767,N_14816);
nor UO_1211 (O_1211,N_14770,N_14906);
nand UO_1212 (O_1212,N_14911,N_14992);
xor UO_1213 (O_1213,N_14953,N_14854);
xor UO_1214 (O_1214,N_14856,N_14942);
or UO_1215 (O_1215,N_14975,N_14986);
and UO_1216 (O_1216,N_14996,N_14744);
and UO_1217 (O_1217,N_14737,N_14891);
xor UO_1218 (O_1218,N_14979,N_14767);
xor UO_1219 (O_1219,N_14956,N_14862);
nor UO_1220 (O_1220,N_14991,N_14763);
xnor UO_1221 (O_1221,N_14809,N_14795);
or UO_1222 (O_1222,N_14898,N_14907);
or UO_1223 (O_1223,N_14898,N_14705);
nor UO_1224 (O_1224,N_14995,N_14949);
nand UO_1225 (O_1225,N_14780,N_14933);
xnor UO_1226 (O_1226,N_14782,N_14807);
nor UO_1227 (O_1227,N_14770,N_14976);
xor UO_1228 (O_1228,N_14918,N_14975);
nor UO_1229 (O_1229,N_14951,N_14753);
xnor UO_1230 (O_1230,N_14805,N_14966);
nand UO_1231 (O_1231,N_14764,N_14738);
or UO_1232 (O_1232,N_14964,N_14885);
xor UO_1233 (O_1233,N_14903,N_14831);
nand UO_1234 (O_1234,N_14715,N_14705);
or UO_1235 (O_1235,N_14772,N_14924);
xor UO_1236 (O_1236,N_14750,N_14901);
xor UO_1237 (O_1237,N_14830,N_14711);
nand UO_1238 (O_1238,N_14834,N_14819);
xnor UO_1239 (O_1239,N_14849,N_14987);
nor UO_1240 (O_1240,N_14746,N_14775);
nand UO_1241 (O_1241,N_14765,N_14752);
nor UO_1242 (O_1242,N_14843,N_14964);
and UO_1243 (O_1243,N_14934,N_14887);
and UO_1244 (O_1244,N_14742,N_14972);
and UO_1245 (O_1245,N_14795,N_14708);
and UO_1246 (O_1246,N_14903,N_14870);
and UO_1247 (O_1247,N_14849,N_14949);
nor UO_1248 (O_1248,N_14923,N_14815);
nand UO_1249 (O_1249,N_14710,N_14875);
and UO_1250 (O_1250,N_14836,N_14916);
xnor UO_1251 (O_1251,N_14759,N_14907);
nand UO_1252 (O_1252,N_14831,N_14773);
xor UO_1253 (O_1253,N_14876,N_14762);
nor UO_1254 (O_1254,N_14724,N_14912);
and UO_1255 (O_1255,N_14784,N_14851);
and UO_1256 (O_1256,N_14975,N_14873);
nor UO_1257 (O_1257,N_14875,N_14861);
and UO_1258 (O_1258,N_14903,N_14801);
nor UO_1259 (O_1259,N_14775,N_14992);
or UO_1260 (O_1260,N_14828,N_14756);
and UO_1261 (O_1261,N_14866,N_14920);
nand UO_1262 (O_1262,N_14981,N_14803);
nand UO_1263 (O_1263,N_14754,N_14753);
xnor UO_1264 (O_1264,N_14947,N_14804);
xor UO_1265 (O_1265,N_14789,N_14844);
xnor UO_1266 (O_1266,N_14808,N_14793);
and UO_1267 (O_1267,N_14810,N_14727);
and UO_1268 (O_1268,N_14917,N_14888);
nand UO_1269 (O_1269,N_14817,N_14880);
nand UO_1270 (O_1270,N_14931,N_14956);
xnor UO_1271 (O_1271,N_14854,N_14989);
nor UO_1272 (O_1272,N_14862,N_14870);
and UO_1273 (O_1273,N_14793,N_14913);
xnor UO_1274 (O_1274,N_14858,N_14938);
and UO_1275 (O_1275,N_14959,N_14897);
nand UO_1276 (O_1276,N_14753,N_14912);
nor UO_1277 (O_1277,N_14734,N_14843);
and UO_1278 (O_1278,N_14800,N_14709);
and UO_1279 (O_1279,N_14759,N_14816);
nand UO_1280 (O_1280,N_14709,N_14805);
nor UO_1281 (O_1281,N_14857,N_14939);
and UO_1282 (O_1282,N_14917,N_14893);
xnor UO_1283 (O_1283,N_14841,N_14833);
nor UO_1284 (O_1284,N_14931,N_14965);
nand UO_1285 (O_1285,N_14738,N_14923);
nand UO_1286 (O_1286,N_14900,N_14832);
or UO_1287 (O_1287,N_14810,N_14975);
nor UO_1288 (O_1288,N_14901,N_14813);
nand UO_1289 (O_1289,N_14908,N_14804);
xor UO_1290 (O_1290,N_14719,N_14845);
and UO_1291 (O_1291,N_14785,N_14945);
nand UO_1292 (O_1292,N_14825,N_14990);
or UO_1293 (O_1293,N_14838,N_14883);
nand UO_1294 (O_1294,N_14812,N_14989);
xor UO_1295 (O_1295,N_14879,N_14875);
nand UO_1296 (O_1296,N_14832,N_14906);
and UO_1297 (O_1297,N_14825,N_14811);
and UO_1298 (O_1298,N_14717,N_14850);
xor UO_1299 (O_1299,N_14762,N_14883);
nor UO_1300 (O_1300,N_14985,N_14749);
xor UO_1301 (O_1301,N_14923,N_14866);
and UO_1302 (O_1302,N_14923,N_14846);
and UO_1303 (O_1303,N_14745,N_14889);
or UO_1304 (O_1304,N_14983,N_14827);
and UO_1305 (O_1305,N_14922,N_14782);
and UO_1306 (O_1306,N_14981,N_14700);
nand UO_1307 (O_1307,N_14994,N_14727);
xnor UO_1308 (O_1308,N_14724,N_14906);
nor UO_1309 (O_1309,N_14848,N_14873);
nor UO_1310 (O_1310,N_14929,N_14936);
or UO_1311 (O_1311,N_14804,N_14709);
xnor UO_1312 (O_1312,N_14804,N_14813);
nor UO_1313 (O_1313,N_14708,N_14787);
and UO_1314 (O_1314,N_14902,N_14972);
or UO_1315 (O_1315,N_14836,N_14805);
nand UO_1316 (O_1316,N_14909,N_14883);
or UO_1317 (O_1317,N_14825,N_14951);
and UO_1318 (O_1318,N_14907,N_14777);
nand UO_1319 (O_1319,N_14921,N_14820);
nand UO_1320 (O_1320,N_14817,N_14783);
nor UO_1321 (O_1321,N_14893,N_14949);
and UO_1322 (O_1322,N_14847,N_14794);
or UO_1323 (O_1323,N_14704,N_14719);
and UO_1324 (O_1324,N_14722,N_14933);
xor UO_1325 (O_1325,N_14824,N_14728);
nand UO_1326 (O_1326,N_14788,N_14935);
or UO_1327 (O_1327,N_14760,N_14983);
and UO_1328 (O_1328,N_14750,N_14909);
and UO_1329 (O_1329,N_14726,N_14827);
xnor UO_1330 (O_1330,N_14792,N_14980);
or UO_1331 (O_1331,N_14865,N_14915);
nor UO_1332 (O_1332,N_14968,N_14738);
xnor UO_1333 (O_1333,N_14731,N_14782);
nand UO_1334 (O_1334,N_14918,N_14775);
xnor UO_1335 (O_1335,N_14969,N_14822);
nor UO_1336 (O_1336,N_14841,N_14842);
nand UO_1337 (O_1337,N_14854,N_14875);
and UO_1338 (O_1338,N_14862,N_14911);
or UO_1339 (O_1339,N_14872,N_14886);
and UO_1340 (O_1340,N_14812,N_14781);
and UO_1341 (O_1341,N_14788,N_14763);
nor UO_1342 (O_1342,N_14731,N_14746);
or UO_1343 (O_1343,N_14905,N_14848);
nand UO_1344 (O_1344,N_14776,N_14707);
or UO_1345 (O_1345,N_14852,N_14902);
and UO_1346 (O_1346,N_14749,N_14904);
nand UO_1347 (O_1347,N_14892,N_14746);
xor UO_1348 (O_1348,N_14736,N_14750);
nand UO_1349 (O_1349,N_14991,N_14940);
xor UO_1350 (O_1350,N_14811,N_14843);
and UO_1351 (O_1351,N_14781,N_14841);
nand UO_1352 (O_1352,N_14835,N_14810);
nand UO_1353 (O_1353,N_14927,N_14751);
nand UO_1354 (O_1354,N_14938,N_14704);
nor UO_1355 (O_1355,N_14974,N_14846);
nand UO_1356 (O_1356,N_14734,N_14885);
and UO_1357 (O_1357,N_14811,N_14924);
or UO_1358 (O_1358,N_14812,N_14743);
xor UO_1359 (O_1359,N_14997,N_14984);
or UO_1360 (O_1360,N_14818,N_14971);
and UO_1361 (O_1361,N_14851,N_14964);
nor UO_1362 (O_1362,N_14945,N_14799);
or UO_1363 (O_1363,N_14937,N_14883);
or UO_1364 (O_1364,N_14701,N_14871);
xnor UO_1365 (O_1365,N_14764,N_14836);
nand UO_1366 (O_1366,N_14890,N_14710);
nand UO_1367 (O_1367,N_14783,N_14943);
nand UO_1368 (O_1368,N_14887,N_14705);
and UO_1369 (O_1369,N_14927,N_14839);
nor UO_1370 (O_1370,N_14825,N_14824);
or UO_1371 (O_1371,N_14849,N_14935);
nand UO_1372 (O_1372,N_14816,N_14882);
xnor UO_1373 (O_1373,N_14968,N_14910);
or UO_1374 (O_1374,N_14876,N_14851);
nand UO_1375 (O_1375,N_14766,N_14807);
or UO_1376 (O_1376,N_14729,N_14790);
or UO_1377 (O_1377,N_14800,N_14952);
nor UO_1378 (O_1378,N_14722,N_14922);
xor UO_1379 (O_1379,N_14815,N_14940);
xnor UO_1380 (O_1380,N_14979,N_14904);
nand UO_1381 (O_1381,N_14728,N_14895);
nand UO_1382 (O_1382,N_14777,N_14913);
nor UO_1383 (O_1383,N_14750,N_14784);
nor UO_1384 (O_1384,N_14977,N_14832);
xnor UO_1385 (O_1385,N_14935,N_14739);
or UO_1386 (O_1386,N_14790,N_14737);
and UO_1387 (O_1387,N_14849,N_14745);
or UO_1388 (O_1388,N_14736,N_14738);
or UO_1389 (O_1389,N_14846,N_14804);
nor UO_1390 (O_1390,N_14986,N_14924);
or UO_1391 (O_1391,N_14764,N_14936);
and UO_1392 (O_1392,N_14778,N_14857);
and UO_1393 (O_1393,N_14731,N_14926);
nor UO_1394 (O_1394,N_14979,N_14893);
nand UO_1395 (O_1395,N_14793,N_14930);
and UO_1396 (O_1396,N_14856,N_14836);
and UO_1397 (O_1397,N_14725,N_14947);
nor UO_1398 (O_1398,N_14955,N_14746);
or UO_1399 (O_1399,N_14718,N_14872);
or UO_1400 (O_1400,N_14780,N_14730);
xor UO_1401 (O_1401,N_14830,N_14998);
nor UO_1402 (O_1402,N_14972,N_14806);
or UO_1403 (O_1403,N_14780,N_14860);
nand UO_1404 (O_1404,N_14846,N_14980);
nand UO_1405 (O_1405,N_14836,N_14878);
nor UO_1406 (O_1406,N_14867,N_14948);
nor UO_1407 (O_1407,N_14965,N_14906);
and UO_1408 (O_1408,N_14737,N_14976);
and UO_1409 (O_1409,N_14858,N_14852);
or UO_1410 (O_1410,N_14862,N_14735);
nor UO_1411 (O_1411,N_14862,N_14766);
nand UO_1412 (O_1412,N_14827,N_14710);
and UO_1413 (O_1413,N_14966,N_14726);
and UO_1414 (O_1414,N_14742,N_14854);
nand UO_1415 (O_1415,N_14788,N_14976);
or UO_1416 (O_1416,N_14917,N_14786);
nor UO_1417 (O_1417,N_14758,N_14977);
and UO_1418 (O_1418,N_14756,N_14912);
nand UO_1419 (O_1419,N_14721,N_14770);
nand UO_1420 (O_1420,N_14768,N_14922);
and UO_1421 (O_1421,N_14788,N_14977);
nand UO_1422 (O_1422,N_14752,N_14948);
nand UO_1423 (O_1423,N_14704,N_14781);
and UO_1424 (O_1424,N_14770,N_14862);
or UO_1425 (O_1425,N_14804,N_14897);
or UO_1426 (O_1426,N_14721,N_14775);
nor UO_1427 (O_1427,N_14812,N_14943);
or UO_1428 (O_1428,N_14986,N_14968);
nand UO_1429 (O_1429,N_14784,N_14714);
xor UO_1430 (O_1430,N_14727,N_14804);
nor UO_1431 (O_1431,N_14797,N_14877);
or UO_1432 (O_1432,N_14970,N_14737);
or UO_1433 (O_1433,N_14877,N_14914);
and UO_1434 (O_1434,N_14712,N_14926);
and UO_1435 (O_1435,N_14879,N_14915);
xnor UO_1436 (O_1436,N_14891,N_14769);
and UO_1437 (O_1437,N_14842,N_14931);
nand UO_1438 (O_1438,N_14845,N_14862);
nor UO_1439 (O_1439,N_14894,N_14774);
nand UO_1440 (O_1440,N_14827,N_14812);
xor UO_1441 (O_1441,N_14957,N_14990);
or UO_1442 (O_1442,N_14751,N_14771);
nand UO_1443 (O_1443,N_14717,N_14747);
xnor UO_1444 (O_1444,N_14840,N_14849);
xnor UO_1445 (O_1445,N_14929,N_14721);
nand UO_1446 (O_1446,N_14756,N_14914);
xor UO_1447 (O_1447,N_14952,N_14925);
nand UO_1448 (O_1448,N_14941,N_14966);
or UO_1449 (O_1449,N_14888,N_14836);
nand UO_1450 (O_1450,N_14763,N_14794);
or UO_1451 (O_1451,N_14979,N_14855);
nand UO_1452 (O_1452,N_14786,N_14874);
nor UO_1453 (O_1453,N_14721,N_14821);
xnor UO_1454 (O_1454,N_14878,N_14958);
nor UO_1455 (O_1455,N_14700,N_14839);
nand UO_1456 (O_1456,N_14875,N_14765);
and UO_1457 (O_1457,N_14737,N_14962);
nand UO_1458 (O_1458,N_14749,N_14714);
nand UO_1459 (O_1459,N_14949,N_14840);
or UO_1460 (O_1460,N_14765,N_14744);
and UO_1461 (O_1461,N_14760,N_14878);
and UO_1462 (O_1462,N_14832,N_14880);
nor UO_1463 (O_1463,N_14799,N_14703);
xnor UO_1464 (O_1464,N_14755,N_14919);
xnor UO_1465 (O_1465,N_14860,N_14729);
nor UO_1466 (O_1466,N_14809,N_14714);
and UO_1467 (O_1467,N_14893,N_14811);
or UO_1468 (O_1468,N_14714,N_14938);
xnor UO_1469 (O_1469,N_14751,N_14938);
nor UO_1470 (O_1470,N_14793,N_14706);
nand UO_1471 (O_1471,N_14877,N_14792);
xor UO_1472 (O_1472,N_14880,N_14959);
and UO_1473 (O_1473,N_14953,N_14715);
nor UO_1474 (O_1474,N_14735,N_14991);
nand UO_1475 (O_1475,N_14981,N_14933);
and UO_1476 (O_1476,N_14909,N_14746);
nor UO_1477 (O_1477,N_14861,N_14717);
xor UO_1478 (O_1478,N_14823,N_14750);
xor UO_1479 (O_1479,N_14901,N_14801);
and UO_1480 (O_1480,N_14737,N_14714);
or UO_1481 (O_1481,N_14765,N_14796);
xor UO_1482 (O_1482,N_14972,N_14993);
and UO_1483 (O_1483,N_14811,N_14800);
xnor UO_1484 (O_1484,N_14787,N_14874);
nor UO_1485 (O_1485,N_14964,N_14834);
and UO_1486 (O_1486,N_14869,N_14730);
or UO_1487 (O_1487,N_14742,N_14946);
or UO_1488 (O_1488,N_14819,N_14738);
nand UO_1489 (O_1489,N_14815,N_14806);
nand UO_1490 (O_1490,N_14897,N_14810);
and UO_1491 (O_1491,N_14857,N_14959);
nor UO_1492 (O_1492,N_14843,N_14929);
and UO_1493 (O_1493,N_14867,N_14776);
xor UO_1494 (O_1494,N_14944,N_14753);
nand UO_1495 (O_1495,N_14747,N_14881);
nor UO_1496 (O_1496,N_14776,N_14947);
nor UO_1497 (O_1497,N_14864,N_14775);
and UO_1498 (O_1498,N_14938,N_14823);
nand UO_1499 (O_1499,N_14967,N_14956);
or UO_1500 (O_1500,N_14916,N_14891);
nand UO_1501 (O_1501,N_14700,N_14911);
nor UO_1502 (O_1502,N_14899,N_14864);
xor UO_1503 (O_1503,N_14793,N_14812);
nor UO_1504 (O_1504,N_14934,N_14824);
or UO_1505 (O_1505,N_14722,N_14916);
or UO_1506 (O_1506,N_14826,N_14877);
nor UO_1507 (O_1507,N_14912,N_14817);
or UO_1508 (O_1508,N_14744,N_14829);
or UO_1509 (O_1509,N_14887,N_14991);
nor UO_1510 (O_1510,N_14994,N_14890);
and UO_1511 (O_1511,N_14882,N_14730);
and UO_1512 (O_1512,N_14880,N_14791);
xor UO_1513 (O_1513,N_14840,N_14866);
and UO_1514 (O_1514,N_14757,N_14848);
or UO_1515 (O_1515,N_14877,N_14835);
nand UO_1516 (O_1516,N_14949,N_14739);
and UO_1517 (O_1517,N_14873,N_14787);
nor UO_1518 (O_1518,N_14811,N_14892);
and UO_1519 (O_1519,N_14955,N_14891);
nand UO_1520 (O_1520,N_14961,N_14929);
or UO_1521 (O_1521,N_14951,N_14869);
or UO_1522 (O_1522,N_14949,N_14842);
nor UO_1523 (O_1523,N_14940,N_14820);
xnor UO_1524 (O_1524,N_14844,N_14819);
and UO_1525 (O_1525,N_14845,N_14835);
nand UO_1526 (O_1526,N_14780,N_14970);
xnor UO_1527 (O_1527,N_14815,N_14769);
and UO_1528 (O_1528,N_14747,N_14709);
nor UO_1529 (O_1529,N_14700,N_14890);
nand UO_1530 (O_1530,N_14967,N_14748);
xnor UO_1531 (O_1531,N_14752,N_14822);
nor UO_1532 (O_1532,N_14951,N_14848);
xnor UO_1533 (O_1533,N_14916,N_14832);
xor UO_1534 (O_1534,N_14930,N_14984);
and UO_1535 (O_1535,N_14924,N_14861);
or UO_1536 (O_1536,N_14992,N_14885);
nor UO_1537 (O_1537,N_14953,N_14726);
and UO_1538 (O_1538,N_14941,N_14808);
nand UO_1539 (O_1539,N_14725,N_14835);
nand UO_1540 (O_1540,N_14824,N_14730);
or UO_1541 (O_1541,N_14947,N_14744);
nor UO_1542 (O_1542,N_14906,N_14986);
and UO_1543 (O_1543,N_14786,N_14947);
xor UO_1544 (O_1544,N_14881,N_14772);
xnor UO_1545 (O_1545,N_14969,N_14869);
xor UO_1546 (O_1546,N_14798,N_14951);
nand UO_1547 (O_1547,N_14711,N_14874);
nor UO_1548 (O_1548,N_14815,N_14835);
nand UO_1549 (O_1549,N_14996,N_14915);
nand UO_1550 (O_1550,N_14837,N_14996);
nand UO_1551 (O_1551,N_14958,N_14750);
nor UO_1552 (O_1552,N_14704,N_14712);
nor UO_1553 (O_1553,N_14982,N_14859);
or UO_1554 (O_1554,N_14989,N_14965);
nand UO_1555 (O_1555,N_14966,N_14714);
or UO_1556 (O_1556,N_14800,N_14719);
nor UO_1557 (O_1557,N_14855,N_14828);
xnor UO_1558 (O_1558,N_14780,N_14876);
and UO_1559 (O_1559,N_14981,N_14791);
nand UO_1560 (O_1560,N_14853,N_14912);
or UO_1561 (O_1561,N_14846,N_14810);
nor UO_1562 (O_1562,N_14945,N_14948);
nand UO_1563 (O_1563,N_14986,N_14995);
or UO_1564 (O_1564,N_14826,N_14962);
and UO_1565 (O_1565,N_14706,N_14975);
or UO_1566 (O_1566,N_14703,N_14739);
or UO_1567 (O_1567,N_14941,N_14914);
nand UO_1568 (O_1568,N_14969,N_14867);
and UO_1569 (O_1569,N_14718,N_14739);
and UO_1570 (O_1570,N_14725,N_14946);
nor UO_1571 (O_1571,N_14982,N_14702);
nand UO_1572 (O_1572,N_14913,N_14711);
xnor UO_1573 (O_1573,N_14962,N_14742);
or UO_1574 (O_1574,N_14785,N_14719);
nor UO_1575 (O_1575,N_14751,N_14800);
or UO_1576 (O_1576,N_14746,N_14799);
and UO_1577 (O_1577,N_14766,N_14829);
nor UO_1578 (O_1578,N_14731,N_14915);
nor UO_1579 (O_1579,N_14911,N_14826);
nor UO_1580 (O_1580,N_14895,N_14838);
nor UO_1581 (O_1581,N_14890,N_14958);
or UO_1582 (O_1582,N_14841,N_14887);
or UO_1583 (O_1583,N_14888,N_14784);
nand UO_1584 (O_1584,N_14908,N_14866);
and UO_1585 (O_1585,N_14815,N_14853);
nor UO_1586 (O_1586,N_14949,N_14940);
nand UO_1587 (O_1587,N_14796,N_14968);
or UO_1588 (O_1588,N_14961,N_14840);
or UO_1589 (O_1589,N_14780,N_14756);
nand UO_1590 (O_1590,N_14896,N_14711);
xnor UO_1591 (O_1591,N_14807,N_14979);
and UO_1592 (O_1592,N_14811,N_14783);
nor UO_1593 (O_1593,N_14818,N_14913);
nor UO_1594 (O_1594,N_14958,N_14741);
xnor UO_1595 (O_1595,N_14914,N_14773);
xnor UO_1596 (O_1596,N_14999,N_14734);
nor UO_1597 (O_1597,N_14735,N_14944);
and UO_1598 (O_1598,N_14702,N_14724);
and UO_1599 (O_1599,N_14957,N_14835);
nor UO_1600 (O_1600,N_14890,N_14820);
xnor UO_1601 (O_1601,N_14950,N_14785);
or UO_1602 (O_1602,N_14845,N_14801);
nand UO_1603 (O_1603,N_14786,N_14983);
or UO_1604 (O_1604,N_14740,N_14891);
and UO_1605 (O_1605,N_14725,N_14908);
nor UO_1606 (O_1606,N_14750,N_14790);
and UO_1607 (O_1607,N_14718,N_14838);
xnor UO_1608 (O_1608,N_14980,N_14773);
or UO_1609 (O_1609,N_14703,N_14710);
and UO_1610 (O_1610,N_14957,N_14877);
and UO_1611 (O_1611,N_14799,N_14836);
nand UO_1612 (O_1612,N_14893,N_14850);
nand UO_1613 (O_1613,N_14828,N_14746);
nor UO_1614 (O_1614,N_14760,N_14876);
and UO_1615 (O_1615,N_14981,N_14921);
and UO_1616 (O_1616,N_14709,N_14966);
xnor UO_1617 (O_1617,N_14737,N_14919);
nor UO_1618 (O_1618,N_14837,N_14914);
or UO_1619 (O_1619,N_14717,N_14710);
xor UO_1620 (O_1620,N_14908,N_14823);
nand UO_1621 (O_1621,N_14848,N_14845);
nand UO_1622 (O_1622,N_14761,N_14740);
nor UO_1623 (O_1623,N_14870,N_14890);
and UO_1624 (O_1624,N_14718,N_14921);
nand UO_1625 (O_1625,N_14876,N_14985);
or UO_1626 (O_1626,N_14732,N_14783);
xor UO_1627 (O_1627,N_14895,N_14776);
or UO_1628 (O_1628,N_14820,N_14764);
and UO_1629 (O_1629,N_14986,N_14798);
xnor UO_1630 (O_1630,N_14793,N_14847);
nand UO_1631 (O_1631,N_14988,N_14775);
nand UO_1632 (O_1632,N_14961,N_14731);
xor UO_1633 (O_1633,N_14761,N_14763);
or UO_1634 (O_1634,N_14858,N_14965);
and UO_1635 (O_1635,N_14885,N_14996);
nor UO_1636 (O_1636,N_14728,N_14916);
xor UO_1637 (O_1637,N_14758,N_14759);
nor UO_1638 (O_1638,N_14867,N_14788);
and UO_1639 (O_1639,N_14765,N_14824);
and UO_1640 (O_1640,N_14990,N_14826);
and UO_1641 (O_1641,N_14903,N_14813);
and UO_1642 (O_1642,N_14845,N_14751);
and UO_1643 (O_1643,N_14792,N_14867);
xnor UO_1644 (O_1644,N_14794,N_14752);
nor UO_1645 (O_1645,N_14725,N_14822);
and UO_1646 (O_1646,N_14779,N_14723);
xnor UO_1647 (O_1647,N_14787,N_14957);
or UO_1648 (O_1648,N_14940,N_14969);
nand UO_1649 (O_1649,N_14715,N_14813);
or UO_1650 (O_1650,N_14763,N_14905);
nand UO_1651 (O_1651,N_14899,N_14959);
xnor UO_1652 (O_1652,N_14731,N_14992);
xor UO_1653 (O_1653,N_14819,N_14893);
nor UO_1654 (O_1654,N_14855,N_14971);
and UO_1655 (O_1655,N_14782,N_14707);
or UO_1656 (O_1656,N_14783,N_14975);
xnor UO_1657 (O_1657,N_14789,N_14767);
nand UO_1658 (O_1658,N_14847,N_14813);
nand UO_1659 (O_1659,N_14709,N_14921);
or UO_1660 (O_1660,N_14765,N_14852);
or UO_1661 (O_1661,N_14738,N_14786);
and UO_1662 (O_1662,N_14790,N_14755);
and UO_1663 (O_1663,N_14741,N_14780);
nor UO_1664 (O_1664,N_14911,N_14818);
or UO_1665 (O_1665,N_14918,N_14873);
xor UO_1666 (O_1666,N_14856,N_14772);
or UO_1667 (O_1667,N_14972,N_14732);
xor UO_1668 (O_1668,N_14934,N_14877);
nand UO_1669 (O_1669,N_14946,N_14720);
or UO_1670 (O_1670,N_14894,N_14912);
and UO_1671 (O_1671,N_14976,N_14839);
nand UO_1672 (O_1672,N_14820,N_14919);
nand UO_1673 (O_1673,N_14989,N_14739);
nand UO_1674 (O_1674,N_14997,N_14711);
nor UO_1675 (O_1675,N_14723,N_14941);
or UO_1676 (O_1676,N_14742,N_14871);
and UO_1677 (O_1677,N_14943,N_14955);
xnor UO_1678 (O_1678,N_14921,N_14780);
nand UO_1679 (O_1679,N_14891,N_14939);
xnor UO_1680 (O_1680,N_14787,N_14949);
nor UO_1681 (O_1681,N_14984,N_14832);
and UO_1682 (O_1682,N_14947,N_14784);
xor UO_1683 (O_1683,N_14996,N_14792);
nand UO_1684 (O_1684,N_14730,N_14826);
nand UO_1685 (O_1685,N_14721,N_14786);
nor UO_1686 (O_1686,N_14927,N_14892);
nand UO_1687 (O_1687,N_14765,N_14967);
nor UO_1688 (O_1688,N_14876,N_14930);
and UO_1689 (O_1689,N_14956,N_14926);
nor UO_1690 (O_1690,N_14701,N_14818);
xnor UO_1691 (O_1691,N_14748,N_14847);
nand UO_1692 (O_1692,N_14827,N_14702);
xor UO_1693 (O_1693,N_14711,N_14967);
or UO_1694 (O_1694,N_14821,N_14957);
nand UO_1695 (O_1695,N_14872,N_14949);
nor UO_1696 (O_1696,N_14883,N_14842);
or UO_1697 (O_1697,N_14755,N_14929);
xnor UO_1698 (O_1698,N_14959,N_14731);
or UO_1699 (O_1699,N_14855,N_14907);
xnor UO_1700 (O_1700,N_14922,N_14738);
and UO_1701 (O_1701,N_14706,N_14861);
nand UO_1702 (O_1702,N_14825,N_14815);
xor UO_1703 (O_1703,N_14820,N_14973);
and UO_1704 (O_1704,N_14918,N_14840);
nor UO_1705 (O_1705,N_14799,N_14711);
xnor UO_1706 (O_1706,N_14861,N_14824);
and UO_1707 (O_1707,N_14789,N_14707);
and UO_1708 (O_1708,N_14829,N_14843);
or UO_1709 (O_1709,N_14855,N_14821);
xnor UO_1710 (O_1710,N_14965,N_14818);
xor UO_1711 (O_1711,N_14911,N_14964);
nand UO_1712 (O_1712,N_14922,N_14855);
and UO_1713 (O_1713,N_14871,N_14944);
or UO_1714 (O_1714,N_14911,N_14918);
xnor UO_1715 (O_1715,N_14983,N_14739);
and UO_1716 (O_1716,N_14762,N_14991);
xor UO_1717 (O_1717,N_14849,N_14760);
nor UO_1718 (O_1718,N_14750,N_14932);
and UO_1719 (O_1719,N_14932,N_14796);
xnor UO_1720 (O_1720,N_14831,N_14906);
or UO_1721 (O_1721,N_14908,N_14953);
or UO_1722 (O_1722,N_14703,N_14853);
xnor UO_1723 (O_1723,N_14705,N_14788);
or UO_1724 (O_1724,N_14962,N_14763);
nor UO_1725 (O_1725,N_14735,N_14713);
or UO_1726 (O_1726,N_14960,N_14779);
and UO_1727 (O_1727,N_14736,N_14782);
xor UO_1728 (O_1728,N_14804,N_14751);
nand UO_1729 (O_1729,N_14701,N_14814);
and UO_1730 (O_1730,N_14856,N_14974);
nand UO_1731 (O_1731,N_14990,N_14993);
nor UO_1732 (O_1732,N_14956,N_14738);
and UO_1733 (O_1733,N_14774,N_14877);
xor UO_1734 (O_1734,N_14778,N_14826);
xor UO_1735 (O_1735,N_14848,N_14701);
or UO_1736 (O_1736,N_14704,N_14761);
and UO_1737 (O_1737,N_14853,N_14914);
and UO_1738 (O_1738,N_14796,N_14819);
xnor UO_1739 (O_1739,N_14841,N_14939);
and UO_1740 (O_1740,N_14772,N_14927);
or UO_1741 (O_1741,N_14999,N_14878);
nor UO_1742 (O_1742,N_14982,N_14917);
nor UO_1743 (O_1743,N_14797,N_14761);
nand UO_1744 (O_1744,N_14919,N_14735);
xnor UO_1745 (O_1745,N_14983,N_14717);
or UO_1746 (O_1746,N_14805,N_14938);
and UO_1747 (O_1747,N_14823,N_14990);
or UO_1748 (O_1748,N_14921,N_14946);
nor UO_1749 (O_1749,N_14792,N_14748);
and UO_1750 (O_1750,N_14962,N_14922);
nor UO_1751 (O_1751,N_14736,N_14773);
or UO_1752 (O_1752,N_14726,N_14942);
nand UO_1753 (O_1753,N_14853,N_14828);
nor UO_1754 (O_1754,N_14867,N_14972);
nand UO_1755 (O_1755,N_14791,N_14828);
nand UO_1756 (O_1756,N_14731,N_14814);
xor UO_1757 (O_1757,N_14800,N_14981);
nor UO_1758 (O_1758,N_14966,N_14784);
and UO_1759 (O_1759,N_14987,N_14742);
nand UO_1760 (O_1760,N_14933,N_14829);
nor UO_1761 (O_1761,N_14838,N_14863);
nand UO_1762 (O_1762,N_14772,N_14737);
nand UO_1763 (O_1763,N_14817,N_14976);
xor UO_1764 (O_1764,N_14963,N_14911);
nor UO_1765 (O_1765,N_14937,N_14736);
and UO_1766 (O_1766,N_14879,N_14995);
xnor UO_1767 (O_1767,N_14836,N_14979);
and UO_1768 (O_1768,N_14885,N_14736);
xor UO_1769 (O_1769,N_14776,N_14830);
xnor UO_1770 (O_1770,N_14998,N_14945);
and UO_1771 (O_1771,N_14848,N_14783);
nand UO_1772 (O_1772,N_14806,N_14911);
and UO_1773 (O_1773,N_14894,N_14767);
nor UO_1774 (O_1774,N_14849,N_14737);
or UO_1775 (O_1775,N_14701,N_14783);
nand UO_1776 (O_1776,N_14875,N_14819);
or UO_1777 (O_1777,N_14973,N_14989);
nand UO_1778 (O_1778,N_14923,N_14961);
nand UO_1779 (O_1779,N_14960,N_14768);
nand UO_1780 (O_1780,N_14805,N_14877);
xor UO_1781 (O_1781,N_14866,N_14941);
xor UO_1782 (O_1782,N_14735,N_14863);
nand UO_1783 (O_1783,N_14895,N_14766);
and UO_1784 (O_1784,N_14740,N_14820);
or UO_1785 (O_1785,N_14755,N_14845);
nor UO_1786 (O_1786,N_14720,N_14901);
xnor UO_1787 (O_1787,N_14869,N_14876);
and UO_1788 (O_1788,N_14761,N_14942);
nor UO_1789 (O_1789,N_14886,N_14953);
nand UO_1790 (O_1790,N_14815,N_14909);
nand UO_1791 (O_1791,N_14814,N_14745);
or UO_1792 (O_1792,N_14775,N_14989);
nor UO_1793 (O_1793,N_14942,N_14733);
and UO_1794 (O_1794,N_14954,N_14750);
and UO_1795 (O_1795,N_14771,N_14808);
nand UO_1796 (O_1796,N_14827,N_14742);
nor UO_1797 (O_1797,N_14879,N_14739);
nor UO_1798 (O_1798,N_14930,N_14813);
nand UO_1799 (O_1799,N_14948,N_14703);
or UO_1800 (O_1800,N_14751,N_14958);
nor UO_1801 (O_1801,N_14753,N_14801);
and UO_1802 (O_1802,N_14999,N_14756);
and UO_1803 (O_1803,N_14897,N_14854);
and UO_1804 (O_1804,N_14978,N_14965);
xnor UO_1805 (O_1805,N_14829,N_14924);
xor UO_1806 (O_1806,N_14922,N_14929);
nor UO_1807 (O_1807,N_14771,N_14830);
nand UO_1808 (O_1808,N_14959,N_14881);
xnor UO_1809 (O_1809,N_14809,N_14928);
nor UO_1810 (O_1810,N_14747,N_14978);
nor UO_1811 (O_1811,N_14751,N_14883);
xnor UO_1812 (O_1812,N_14992,N_14795);
xor UO_1813 (O_1813,N_14765,N_14835);
nor UO_1814 (O_1814,N_14724,N_14952);
or UO_1815 (O_1815,N_14898,N_14785);
or UO_1816 (O_1816,N_14954,N_14988);
or UO_1817 (O_1817,N_14974,N_14721);
and UO_1818 (O_1818,N_14925,N_14910);
or UO_1819 (O_1819,N_14908,N_14859);
and UO_1820 (O_1820,N_14822,N_14930);
or UO_1821 (O_1821,N_14812,N_14767);
and UO_1822 (O_1822,N_14908,N_14851);
and UO_1823 (O_1823,N_14970,N_14749);
xnor UO_1824 (O_1824,N_14893,N_14962);
or UO_1825 (O_1825,N_14894,N_14797);
or UO_1826 (O_1826,N_14825,N_14924);
and UO_1827 (O_1827,N_14829,N_14756);
nor UO_1828 (O_1828,N_14957,N_14760);
nand UO_1829 (O_1829,N_14729,N_14938);
nand UO_1830 (O_1830,N_14702,N_14924);
nand UO_1831 (O_1831,N_14795,N_14863);
and UO_1832 (O_1832,N_14976,N_14910);
nand UO_1833 (O_1833,N_14989,N_14745);
nand UO_1834 (O_1834,N_14803,N_14793);
nand UO_1835 (O_1835,N_14786,N_14742);
and UO_1836 (O_1836,N_14989,N_14960);
or UO_1837 (O_1837,N_14761,N_14741);
xor UO_1838 (O_1838,N_14972,N_14906);
nor UO_1839 (O_1839,N_14918,N_14718);
xnor UO_1840 (O_1840,N_14891,N_14901);
xnor UO_1841 (O_1841,N_14967,N_14858);
nand UO_1842 (O_1842,N_14766,N_14899);
xnor UO_1843 (O_1843,N_14899,N_14747);
xnor UO_1844 (O_1844,N_14800,N_14897);
nor UO_1845 (O_1845,N_14985,N_14928);
xnor UO_1846 (O_1846,N_14994,N_14970);
nand UO_1847 (O_1847,N_14735,N_14719);
or UO_1848 (O_1848,N_14792,N_14765);
xor UO_1849 (O_1849,N_14966,N_14985);
xnor UO_1850 (O_1850,N_14955,N_14715);
or UO_1851 (O_1851,N_14719,N_14946);
or UO_1852 (O_1852,N_14799,N_14919);
and UO_1853 (O_1853,N_14990,N_14886);
nor UO_1854 (O_1854,N_14905,N_14708);
nand UO_1855 (O_1855,N_14911,N_14967);
nor UO_1856 (O_1856,N_14888,N_14969);
or UO_1857 (O_1857,N_14792,N_14844);
and UO_1858 (O_1858,N_14855,N_14705);
nor UO_1859 (O_1859,N_14872,N_14993);
and UO_1860 (O_1860,N_14798,N_14778);
or UO_1861 (O_1861,N_14778,N_14931);
xor UO_1862 (O_1862,N_14770,N_14716);
or UO_1863 (O_1863,N_14812,N_14925);
nor UO_1864 (O_1864,N_14972,N_14878);
xor UO_1865 (O_1865,N_14964,N_14711);
and UO_1866 (O_1866,N_14932,N_14871);
nor UO_1867 (O_1867,N_14900,N_14806);
nor UO_1868 (O_1868,N_14988,N_14750);
nand UO_1869 (O_1869,N_14837,N_14959);
nor UO_1870 (O_1870,N_14734,N_14839);
xnor UO_1871 (O_1871,N_14741,N_14730);
xor UO_1872 (O_1872,N_14813,N_14866);
and UO_1873 (O_1873,N_14956,N_14974);
or UO_1874 (O_1874,N_14954,N_14984);
or UO_1875 (O_1875,N_14915,N_14743);
nand UO_1876 (O_1876,N_14901,N_14940);
or UO_1877 (O_1877,N_14998,N_14754);
or UO_1878 (O_1878,N_14979,N_14799);
or UO_1879 (O_1879,N_14821,N_14912);
and UO_1880 (O_1880,N_14888,N_14799);
nor UO_1881 (O_1881,N_14728,N_14921);
nand UO_1882 (O_1882,N_14813,N_14933);
xor UO_1883 (O_1883,N_14746,N_14804);
xnor UO_1884 (O_1884,N_14749,N_14772);
nand UO_1885 (O_1885,N_14711,N_14977);
nor UO_1886 (O_1886,N_14725,N_14796);
or UO_1887 (O_1887,N_14844,N_14860);
nor UO_1888 (O_1888,N_14971,N_14892);
xor UO_1889 (O_1889,N_14866,N_14823);
nand UO_1890 (O_1890,N_14796,N_14764);
nor UO_1891 (O_1891,N_14956,N_14986);
or UO_1892 (O_1892,N_14916,N_14887);
or UO_1893 (O_1893,N_14998,N_14862);
nor UO_1894 (O_1894,N_14875,N_14713);
nor UO_1895 (O_1895,N_14954,N_14744);
nand UO_1896 (O_1896,N_14984,N_14730);
or UO_1897 (O_1897,N_14935,N_14822);
xor UO_1898 (O_1898,N_14753,N_14727);
xnor UO_1899 (O_1899,N_14766,N_14825);
or UO_1900 (O_1900,N_14889,N_14947);
nor UO_1901 (O_1901,N_14846,N_14768);
nor UO_1902 (O_1902,N_14920,N_14916);
or UO_1903 (O_1903,N_14910,N_14811);
xor UO_1904 (O_1904,N_14938,N_14902);
xor UO_1905 (O_1905,N_14788,N_14849);
and UO_1906 (O_1906,N_14991,N_14710);
or UO_1907 (O_1907,N_14980,N_14966);
or UO_1908 (O_1908,N_14898,N_14890);
or UO_1909 (O_1909,N_14828,N_14882);
nor UO_1910 (O_1910,N_14805,N_14962);
nand UO_1911 (O_1911,N_14957,N_14970);
nor UO_1912 (O_1912,N_14716,N_14790);
or UO_1913 (O_1913,N_14931,N_14943);
xnor UO_1914 (O_1914,N_14960,N_14968);
nand UO_1915 (O_1915,N_14954,N_14981);
and UO_1916 (O_1916,N_14972,N_14774);
or UO_1917 (O_1917,N_14900,N_14894);
xor UO_1918 (O_1918,N_14824,N_14757);
and UO_1919 (O_1919,N_14835,N_14823);
xnor UO_1920 (O_1920,N_14726,N_14701);
or UO_1921 (O_1921,N_14916,N_14851);
and UO_1922 (O_1922,N_14711,N_14903);
nor UO_1923 (O_1923,N_14840,N_14848);
xor UO_1924 (O_1924,N_14721,N_14891);
nand UO_1925 (O_1925,N_14828,N_14808);
nand UO_1926 (O_1926,N_14765,N_14933);
nor UO_1927 (O_1927,N_14999,N_14887);
nand UO_1928 (O_1928,N_14929,N_14737);
or UO_1929 (O_1929,N_14997,N_14841);
xnor UO_1930 (O_1930,N_14775,N_14735);
nor UO_1931 (O_1931,N_14768,N_14856);
nand UO_1932 (O_1932,N_14877,N_14881);
and UO_1933 (O_1933,N_14887,N_14935);
nand UO_1934 (O_1934,N_14763,N_14773);
and UO_1935 (O_1935,N_14721,N_14932);
or UO_1936 (O_1936,N_14780,N_14982);
and UO_1937 (O_1937,N_14988,N_14705);
nor UO_1938 (O_1938,N_14950,N_14965);
xnor UO_1939 (O_1939,N_14881,N_14984);
nor UO_1940 (O_1940,N_14842,N_14871);
nor UO_1941 (O_1941,N_14902,N_14759);
and UO_1942 (O_1942,N_14752,N_14767);
nand UO_1943 (O_1943,N_14734,N_14942);
xnor UO_1944 (O_1944,N_14750,N_14734);
and UO_1945 (O_1945,N_14917,N_14894);
and UO_1946 (O_1946,N_14956,N_14891);
nand UO_1947 (O_1947,N_14955,N_14812);
nand UO_1948 (O_1948,N_14987,N_14780);
xnor UO_1949 (O_1949,N_14830,N_14853);
or UO_1950 (O_1950,N_14970,N_14704);
and UO_1951 (O_1951,N_14989,N_14707);
nand UO_1952 (O_1952,N_14988,N_14903);
xor UO_1953 (O_1953,N_14759,N_14793);
or UO_1954 (O_1954,N_14925,N_14786);
and UO_1955 (O_1955,N_14758,N_14894);
xor UO_1956 (O_1956,N_14956,N_14703);
or UO_1957 (O_1957,N_14854,N_14713);
nand UO_1958 (O_1958,N_14872,N_14887);
nand UO_1959 (O_1959,N_14976,N_14807);
nor UO_1960 (O_1960,N_14740,N_14897);
nor UO_1961 (O_1961,N_14759,N_14865);
and UO_1962 (O_1962,N_14790,N_14918);
and UO_1963 (O_1963,N_14772,N_14918);
xnor UO_1964 (O_1964,N_14727,N_14701);
xor UO_1965 (O_1965,N_14828,N_14862);
nand UO_1966 (O_1966,N_14890,N_14762);
xnor UO_1967 (O_1967,N_14796,N_14833);
nand UO_1968 (O_1968,N_14958,N_14713);
xor UO_1969 (O_1969,N_14737,N_14731);
nand UO_1970 (O_1970,N_14852,N_14842);
and UO_1971 (O_1971,N_14989,N_14875);
nand UO_1972 (O_1972,N_14771,N_14887);
nor UO_1973 (O_1973,N_14842,N_14928);
nor UO_1974 (O_1974,N_14881,N_14762);
nor UO_1975 (O_1975,N_14909,N_14715);
or UO_1976 (O_1976,N_14901,N_14977);
nand UO_1977 (O_1977,N_14757,N_14809);
xor UO_1978 (O_1978,N_14861,N_14898);
or UO_1979 (O_1979,N_14827,N_14954);
xnor UO_1980 (O_1980,N_14806,N_14941);
and UO_1981 (O_1981,N_14795,N_14758);
and UO_1982 (O_1982,N_14758,N_14899);
nor UO_1983 (O_1983,N_14937,N_14813);
and UO_1984 (O_1984,N_14786,N_14896);
nand UO_1985 (O_1985,N_14942,N_14701);
or UO_1986 (O_1986,N_14803,N_14745);
or UO_1987 (O_1987,N_14909,N_14862);
nand UO_1988 (O_1988,N_14928,N_14921);
or UO_1989 (O_1989,N_14876,N_14878);
or UO_1990 (O_1990,N_14936,N_14763);
and UO_1991 (O_1991,N_14842,N_14721);
nor UO_1992 (O_1992,N_14832,N_14839);
nand UO_1993 (O_1993,N_14821,N_14938);
and UO_1994 (O_1994,N_14962,N_14932);
and UO_1995 (O_1995,N_14918,N_14906);
and UO_1996 (O_1996,N_14996,N_14932);
nand UO_1997 (O_1997,N_14884,N_14887);
xor UO_1998 (O_1998,N_14785,N_14769);
and UO_1999 (O_1999,N_14713,N_14771);
endmodule