module basic_1000_10000_1500_2_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5002,N_5005,N_5007,N_5008,N_5010,N_5012,N_5013,N_5016,N_5017,N_5018,N_5019,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5029,N_5034,N_5035,N_5036,N_5037,N_5038,N_5040,N_5041,N_5042,N_5044,N_5045,N_5046,N_5047,N_5049,N_5050,N_5052,N_5055,N_5059,N_5060,N_5061,N_5062,N_5063,N_5066,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5078,N_5079,N_5080,N_5081,N_5083,N_5084,N_5086,N_5087,N_5089,N_5094,N_5095,N_5096,N_5097,N_5100,N_5102,N_5103,N_5104,N_5105,N_5107,N_5109,N_5110,N_5113,N_5115,N_5116,N_5117,N_5119,N_5122,N_5124,N_5125,N_5127,N_5128,N_5130,N_5131,N_5133,N_5138,N_5139,N_5144,N_5146,N_5147,N_5151,N_5152,N_5153,N_5154,N_5156,N_5157,N_5158,N_5160,N_5161,N_5162,N_5166,N_5169,N_5171,N_5172,N_5173,N_5174,N_5175,N_5178,N_5179,N_5180,N_5182,N_5183,N_5184,N_5186,N_5188,N_5189,N_5190,N_5195,N_5199,N_5200,N_5201,N_5203,N_5205,N_5207,N_5213,N_5216,N_5217,N_5221,N_5224,N_5225,N_5226,N_5228,N_5229,N_5230,N_5231,N_5233,N_5235,N_5239,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5251,N_5252,N_5255,N_5258,N_5259,N_5261,N_5263,N_5264,N_5266,N_5267,N_5269,N_5270,N_5271,N_5272,N_5274,N_5275,N_5276,N_5278,N_5279,N_5282,N_5283,N_5284,N_5286,N_5288,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5310,N_5311,N_5313,N_5314,N_5315,N_5316,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5327,N_5328,N_5329,N_5330,N_5332,N_5335,N_5336,N_5337,N_5340,N_5342,N_5343,N_5344,N_5345,N_5346,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5357,N_5359,N_5360,N_5361,N_5365,N_5366,N_5368,N_5373,N_5375,N_5376,N_5378,N_5379,N_5381,N_5382,N_5383,N_5384,N_5385,N_5387,N_5388,N_5389,N_5390,N_5391,N_5393,N_5397,N_5399,N_5402,N_5403,N_5404,N_5405,N_5408,N_5411,N_5412,N_5414,N_5415,N_5416,N_5417,N_5419,N_5422,N_5423,N_5430,N_5431,N_5433,N_5434,N_5436,N_5438,N_5440,N_5441,N_5446,N_5448,N_5449,N_5450,N_5452,N_5453,N_5454,N_5455,N_5456,N_5458,N_5461,N_5462,N_5464,N_5467,N_5468,N_5469,N_5471,N_5477,N_5479,N_5480,N_5481,N_5483,N_5485,N_5486,N_5487,N_5488,N_5491,N_5493,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5504,N_5505,N_5506,N_5507,N_5509,N_5510,N_5516,N_5517,N_5518,N_5519,N_5521,N_5523,N_5524,N_5525,N_5526,N_5527,N_5529,N_5530,N_5532,N_5533,N_5535,N_5537,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5547,N_5548,N_5549,N_5552,N_5553,N_5554,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5567,N_5569,N_5571,N_5572,N_5575,N_5576,N_5581,N_5582,N_5587,N_5589,N_5590,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5599,N_5600,N_5601,N_5604,N_5606,N_5609,N_5610,N_5611,N_5613,N_5614,N_5617,N_5618,N_5621,N_5622,N_5623,N_5624,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5634,N_5635,N_5636,N_5638,N_5640,N_5641,N_5642,N_5643,N_5644,N_5646,N_5647,N_5649,N_5650,N_5651,N_5652,N_5653,N_5655,N_5657,N_5658,N_5660,N_5662,N_5663,N_5664,N_5665,N_5666,N_5668,N_5669,N_5670,N_5672,N_5676,N_5678,N_5683,N_5684,N_5685,N_5686,N_5689,N_5690,N_5691,N_5693,N_5694,N_5696,N_5698,N_5699,N_5700,N_5701,N_5702,N_5704,N_5708,N_5712,N_5713,N_5715,N_5716,N_5717,N_5718,N_5720,N_5721,N_5722,N_5723,N_5724,N_5730,N_5731,N_5732,N_5735,N_5736,N_5737,N_5738,N_5739,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5750,N_5751,N_5752,N_5753,N_5755,N_5756,N_5757,N_5761,N_5762,N_5765,N_5767,N_5768,N_5771,N_5773,N_5774,N_5776,N_5777,N_5778,N_5780,N_5783,N_5784,N_5785,N_5787,N_5788,N_5789,N_5790,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5799,N_5801,N_5802,N_5803,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5819,N_5822,N_5823,N_5826,N_5827,N_5828,N_5830,N_5832,N_5833,N_5836,N_5837,N_5839,N_5840,N_5842,N_5845,N_5846,N_5847,N_5850,N_5851,N_5854,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5869,N_5871,N_5872,N_5874,N_5875,N_5876,N_5877,N_5878,N_5880,N_5882,N_5883,N_5885,N_5887,N_5892,N_5895,N_5897,N_5898,N_5902,N_5903,N_5905,N_5907,N_5911,N_5912,N_5913,N_5914,N_5916,N_5918,N_5919,N_5921,N_5922,N_5926,N_5928,N_5930,N_5931,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5941,N_5943,N_5944,N_5947,N_5949,N_5951,N_5953,N_5954,N_5957,N_5959,N_5966,N_5967,N_5968,N_5969,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5980,N_5981,N_5983,N_5984,N_5985,N_5987,N_5988,N_5990,N_5991,N_5992,N_5995,N_5996,N_5998,N_6001,N_6002,N_6006,N_6007,N_6009,N_6012,N_6013,N_6014,N_6016,N_6017,N_6019,N_6020,N_6021,N_6022,N_6024,N_6025,N_6026,N_6032,N_6033,N_6035,N_6036,N_6037,N_6040,N_6041,N_6042,N_6043,N_6046,N_6047,N_6048,N_6050,N_6052,N_6053,N_6054,N_6055,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6068,N_6071,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6086,N_6087,N_6088,N_6089,N_6090,N_6094,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6105,N_6107,N_6108,N_6110,N_6112,N_6113,N_6114,N_6115,N_6118,N_6119,N_6121,N_6123,N_6124,N_6125,N_6126,N_6128,N_6129,N_6130,N_6131,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6144,N_6146,N_6148,N_6150,N_6151,N_6152,N_6155,N_6156,N_6157,N_6158,N_6160,N_6161,N_6162,N_6164,N_6166,N_6167,N_6168,N_6169,N_6170,N_6175,N_6177,N_6178,N_6179,N_6181,N_6182,N_6183,N_6185,N_6187,N_6189,N_6190,N_6191,N_6192,N_6193,N_6195,N_6196,N_6197,N_6198,N_6205,N_6206,N_6207,N_6210,N_6211,N_6219,N_6221,N_6222,N_6223,N_6224,N_6229,N_6230,N_6231,N_6232,N_6234,N_6236,N_6239,N_6241,N_6242,N_6245,N_6248,N_6249,N_6252,N_6254,N_6256,N_6258,N_6259,N_6262,N_6264,N_6270,N_6271,N_6272,N_6275,N_6276,N_6278,N_6279,N_6280,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6289,N_6290,N_6291,N_6293,N_6295,N_6297,N_6298,N_6301,N_6303,N_6305,N_6306,N_6309,N_6310,N_6311,N_6313,N_6314,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6323,N_6325,N_6326,N_6327,N_6328,N_6334,N_6335,N_6337,N_6338,N_6339,N_6340,N_6341,N_6344,N_6347,N_6348,N_6350,N_6351,N_6352,N_6353,N_6354,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6395,N_6396,N_6397,N_6399,N_6402,N_6403,N_6405,N_6406,N_6407,N_6409,N_6411,N_6412,N_6413,N_6415,N_6417,N_6418,N_6419,N_6421,N_6422,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6432,N_6433,N_6434,N_6436,N_6439,N_6441,N_6442,N_6444,N_6445,N_6446,N_6447,N_6450,N_6452,N_6453,N_6454,N_6456,N_6457,N_6459,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6470,N_6472,N_6473,N_6475,N_6477,N_6478,N_6479,N_6483,N_6484,N_6487,N_6492,N_6494,N_6497,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6508,N_6511,N_6514,N_6515,N_6517,N_6519,N_6520,N_6521,N_6522,N_6524,N_6525,N_6526,N_6529,N_6530,N_6532,N_6533,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6545,N_6547,N_6548,N_6549,N_6550,N_6554,N_6555,N_6556,N_6557,N_6558,N_6560,N_6561,N_6562,N_6563,N_6566,N_6569,N_6570,N_6571,N_6575,N_6578,N_6579,N_6580,N_6582,N_6583,N_6586,N_6587,N_6589,N_6592,N_6594,N_6596,N_6597,N_6602,N_6603,N_6605,N_6607,N_6608,N_6610,N_6612,N_6615,N_6616,N_6618,N_6620,N_6621,N_6622,N_6623,N_6626,N_6629,N_6631,N_6632,N_6634,N_6636,N_6638,N_6639,N_6641,N_6643,N_6644,N_6645,N_6646,N_6648,N_6651,N_6654,N_6655,N_6656,N_6657,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6671,N_6673,N_6675,N_6677,N_6679,N_6684,N_6685,N_6686,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6696,N_6699,N_6701,N_6702,N_6704,N_6706,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6719,N_6721,N_6723,N_6726,N_6727,N_6728,N_6731,N_6732,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6744,N_6746,N_6748,N_6752,N_6753,N_6754,N_6758,N_6761,N_6762,N_6768,N_6769,N_6770,N_6771,N_6773,N_6774,N_6775,N_6777,N_6778,N_6779,N_6783,N_6784,N_6785,N_6787,N_6788,N_6790,N_6795,N_6796,N_6797,N_6800,N_6801,N_6804,N_6805,N_6807,N_6810,N_6813,N_6814,N_6815,N_6817,N_6819,N_6820,N_6821,N_6823,N_6824,N_6826,N_6828,N_6829,N_6830,N_6831,N_6833,N_6834,N_6836,N_6837,N_6838,N_6841,N_6842,N_6845,N_6846,N_6847,N_6848,N_6851,N_6852,N_6854,N_6855,N_6857,N_6858,N_6861,N_6864,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6875,N_6876,N_6880,N_6882,N_6883,N_6884,N_6885,N_6886,N_6888,N_6889,N_6890,N_6892,N_6895,N_6896,N_6897,N_6899,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6908,N_6909,N_6910,N_6911,N_6912,N_6914,N_6916,N_6917,N_6918,N_6919,N_6920,N_6922,N_6923,N_6924,N_6925,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6938,N_6939,N_6940,N_6941,N_6943,N_6944,N_6945,N_6947,N_6950,N_6951,N_6956,N_6957,N_6960,N_6962,N_6963,N_6964,N_6966,N_6967,N_6968,N_6971,N_6972,N_6973,N_6977,N_6978,N_6982,N_6983,N_6984,N_6985,N_6986,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6995,N_6997,N_6998,N_7000,N_7002,N_7003,N_7004,N_7005,N_7007,N_7009,N_7010,N_7016,N_7018,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7027,N_7028,N_7029,N_7030,N_7032,N_7033,N_7034,N_7035,N_7037,N_7038,N_7039,N_7042,N_7044,N_7045,N_7046,N_7047,N_7049,N_7051,N_7054,N_7055,N_7057,N_7061,N_7063,N_7067,N_7068,N_7069,N_7070,N_7071,N_7074,N_7075,N_7078,N_7079,N_7081,N_7082,N_7084,N_7085,N_7086,N_7088,N_7089,N_7091,N_7092,N_7094,N_7097,N_7098,N_7102,N_7104,N_7106,N_7112,N_7116,N_7118,N_7119,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7133,N_7134,N_7136,N_7137,N_7139,N_7140,N_7141,N_7142,N_7143,N_7145,N_7146,N_7147,N_7150,N_7152,N_7153,N_7156,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7165,N_7166,N_7167,N_7169,N_7171,N_7172,N_7174,N_7176,N_7178,N_7179,N_7181,N_7184,N_7185,N_7186,N_7187,N_7188,N_7190,N_7192,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7205,N_7207,N_7208,N_7209,N_7213,N_7218,N_7219,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7233,N_7234,N_7235,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7248,N_7249,N_7250,N_7252,N_7254,N_7257,N_7259,N_7261,N_7262,N_7263,N_7264,N_7266,N_7267,N_7269,N_7270,N_7272,N_7275,N_7277,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7292,N_7294,N_7295,N_7297,N_7298,N_7299,N_7302,N_7303,N_7304,N_7306,N_7307,N_7309,N_7310,N_7311,N_7312,N_7314,N_7316,N_7318,N_7319,N_7320,N_7323,N_7324,N_7327,N_7328,N_7330,N_7331,N_7332,N_7333,N_7335,N_7336,N_7339,N_7340,N_7341,N_7342,N_7343,N_7346,N_7347,N_7350,N_7351,N_7352,N_7353,N_7355,N_7356,N_7357,N_7360,N_7361,N_7362,N_7364,N_7366,N_7367,N_7369,N_7371,N_7372,N_7373,N_7376,N_7377,N_7378,N_7380,N_7381,N_7384,N_7386,N_7388,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7397,N_7398,N_7399,N_7401,N_7402,N_7403,N_7408,N_7410,N_7411,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7423,N_7427,N_7428,N_7429,N_7430,N_7432,N_7433,N_7434,N_7437,N_7439,N_7440,N_7441,N_7442,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7457,N_7460,N_7461,N_7462,N_7463,N_7465,N_7466,N_7468,N_7469,N_7470,N_7472,N_7480,N_7483,N_7485,N_7490,N_7497,N_7498,N_7504,N_7505,N_7508,N_7509,N_7511,N_7512,N_7515,N_7517,N_7518,N_7521,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7530,N_7532,N_7534,N_7535,N_7536,N_7539,N_7542,N_7546,N_7547,N_7555,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7565,N_7567,N_7570,N_7571,N_7573,N_7574,N_7577,N_7578,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7587,N_7591,N_7592,N_7593,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7605,N_7608,N_7611,N_7612,N_7613,N_7614,N_7615,N_7618,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7638,N_7639,N_7643,N_7644,N_7645,N_7646,N_7647,N_7649,N_7651,N_7652,N_7653,N_7657,N_7658,N_7663,N_7664,N_7666,N_7670,N_7671,N_7672,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7682,N_7683,N_7684,N_7686,N_7687,N_7689,N_7692,N_7694,N_7696,N_7697,N_7698,N_7701,N_7702,N_7703,N_7706,N_7707,N_7708,N_7709,N_7711,N_7713,N_7714,N_7715,N_7717,N_7719,N_7720,N_7721,N_7723,N_7725,N_7726,N_7727,N_7728,N_7729,N_7731,N_7732,N_7734,N_7735,N_7737,N_7738,N_7740,N_7741,N_7743,N_7744,N_7746,N_7747,N_7748,N_7750,N_7753,N_7754,N_7755,N_7756,N_7757,N_7759,N_7760,N_7761,N_7762,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7776,N_7778,N_7779,N_7781,N_7782,N_7783,N_7784,N_7787,N_7788,N_7790,N_7792,N_7793,N_7795,N_7796,N_7797,N_7798,N_7802,N_7803,N_7808,N_7809,N_7810,N_7811,N_7812,N_7814,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7825,N_7828,N_7829,N_7830,N_7835,N_7836,N_7837,N_7841,N_7843,N_7845,N_7846,N_7847,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7870,N_7872,N_7875,N_7876,N_7880,N_7882,N_7884,N_7887,N_7888,N_7890,N_7891,N_7893,N_7896,N_7897,N_7899,N_7900,N_7901,N_7902,N_7905,N_7906,N_7907,N_7908,N_7911,N_7913,N_7915,N_7916,N_7918,N_7920,N_7922,N_7923,N_7925,N_7927,N_7928,N_7930,N_7931,N_7933,N_7934,N_7935,N_7937,N_7938,N_7939,N_7940,N_7942,N_7946,N_7948,N_7950,N_7952,N_7953,N_7954,N_7955,N_7957,N_7958,N_7960,N_7961,N_7962,N_7964,N_7967,N_7968,N_7970,N_7971,N_7972,N_7975,N_7976,N_7979,N_7980,N_7983,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7992,N_7993,N_7995,N_7996,N_7997,N_7999,N_8000,N_8002,N_8003,N_8004,N_8005,N_8007,N_8008,N_8010,N_8012,N_8015,N_8016,N_8017,N_8018,N_8020,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8030,N_8031,N_8034,N_8037,N_8038,N_8042,N_8044,N_8046,N_8047,N_8048,N_8052,N_8056,N_8057,N_8058,N_8060,N_8061,N_8062,N_8063,N_8065,N_8067,N_8069,N_8070,N_8071,N_8073,N_8078,N_8079,N_8081,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8111,N_8113,N_8116,N_8118,N_8119,N_8121,N_8123,N_8124,N_8125,N_8128,N_8129,N_8130,N_8131,N_8133,N_8134,N_8135,N_8136,N_8138,N_8139,N_8142,N_8145,N_8147,N_8148,N_8149,N_8153,N_8155,N_8156,N_8157,N_8161,N_8162,N_8164,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8177,N_8181,N_8182,N_8183,N_8184,N_8187,N_8188,N_8189,N_8190,N_8191,N_8193,N_8194,N_8195,N_8197,N_8198,N_8200,N_8202,N_8203,N_8205,N_8206,N_8207,N_8209,N_8210,N_8212,N_8215,N_8218,N_8222,N_8225,N_8226,N_8227,N_8228,N_8229,N_8232,N_8234,N_8236,N_8238,N_8239,N_8243,N_8244,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8254,N_8255,N_8256,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8267,N_8268,N_8272,N_8273,N_8275,N_8276,N_8277,N_8281,N_8282,N_8283,N_8286,N_8287,N_8288,N_8290,N_8291,N_8294,N_8295,N_8296,N_8297,N_8301,N_8302,N_8303,N_8307,N_8308,N_8309,N_8311,N_8313,N_8314,N_8315,N_8316,N_8318,N_8320,N_8321,N_8324,N_8325,N_8326,N_8328,N_8329,N_8330,N_8332,N_8335,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8350,N_8351,N_8352,N_8353,N_8355,N_8356,N_8357,N_8358,N_8363,N_8364,N_8366,N_8368,N_8369,N_8371,N_8372,N_8376,N_8377,N_8378,N_8381,N_8382,N_8383,N_8387,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8397,N_8398,N_8400,N_8401,N_8403,N_8405,N_8407,N_8408,N_8411,N_8414,N_8415,N_8416,N_8417,N_8418,N_8423,N_8424,N_8427,N_8428,N_8429,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8448,N_8450,N_8451,N_8455,N_8459,N_8460,N_8461,N_8462,N_8464,N_8465,N_8466,N_8467,N_8469,N_8476,N_8479,N_8481,N_8486,N_8488,N_8490,N_8492,N_8493,N_8496,N_8497,N_8499,N_8500,N_8501,N_8502,N_8504,N_8508,N_8509,N_8511,N_8512,N_8514,N_8516,N_8517,N_8520,N_8521,N_8523,N_8524,N_8526,N_8528,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8537,N_8540,N_8542,N_8543,N_8544,N_8547,N_8548,N_8550,N_8551,N_8554,N_8555,N_8556,N_8559,N_8562,N_8563,N_8564,N_8567,N_8568,N_8570,N_8574,N_8575,N_8576,N_8578,N_8579,N_8580,N_8581,N_8583,N_8586,N_8587,N_8588,N_8589,N_8590,N_8592,N_8595,N_8596,N_8599,N_8600,N_8602,N_8604,N_8605,N_8606,N_8608,N_8610,N_8611,N_8614,N_8615,N_8616,N_8617,N_8618,N_8620,N_8622,N_8624,N_8625,N_8626,N_8629,N_8630,N_8634,N_8636,N_8637,N_8638,N_8641,N_8648,N_8649,N_8650,N_8652,N_8653,N_8654,N_8655,N_8657,N_8658,N_8659,N_8660,N_8663,N_8665,N_8666,N_8668,N_8669,N_8671,N_8674,N_8675,N_8676,N_8677,N_8679,N_8680,N_8681,N_8682,N_8685,N_8686,N_8687,N_8688,N_8691,N_8693,N_8694,N_8695,N_8696,N_8698,N_8699,N_8701,N_8704,N_8705,N_8706,N_8710,N_8711,N_8715,N_8716,N_8717,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8727,N_8732,N_8734,N_8735,N_8736,N_8737,N_8739,N_8740,N_8741,N_8742,N_8743,N_8745,N_8747,N_8748,N_8752,N_8754,N_8756,N_8758,N_8760,N_8762,N_8763,N_8765,N_8767,N_8768,N_8770,N_8771,N_8772,N_8774,N_8776,N_8778,N_8779,N_8783,N_8785,N_8786,N_8787,N_8788,N_8790,N_8793,N_8794,N_8795,N_8796,N_8798,N_8799,N_8801,N_8802,N_8804,N_8806,N_8808,N_8811,N_8812,N_8813,N_8815,N_8825,N_8826,N_8829,N_8830,N_8831,N_8832,N_8835,N_8836,N_8838,N_8839,N_8841,N_8842,N_8843,N_8844,N_8846,N_8847,N_8848,N_8850,N_8852,N_8854,N_8857,N_8859,N_8861,N_8862,N_8865,N_8869,N_8870,N_8871,N_8874,N_8876,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8885,N_8887,N_8890,N_8895,N_8896,N_8897,N_8898,N_8901,N_8902,N_8904,N_8905,N_8906,N_8908,N_8909,N_8910,N_8913,N_8917,N_8918,N_8920,N_8922,N_8925,N_8926,N_8927,N_8928,N_8930,N_8931,N_8932,N_8934,N_8935,N_8936,N_8938,N_8940,N_8942,N_8945,N_8947,N_8948,N_8950,N_8951,N_8954,N_8955,N_8957,N_8958,N_8961,N_8964,N_8965,N_8966,N_8967,N_8969,N_8970,N_8971,N_8973,N_8974,N_8976,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8998,N_8999,N_9000,N_9005,N_9006,N_9007,N_9010,N_9011,N_9015,N_9017,N_9020,N_9021,N_9023,N_9024,N_9025,N_9027,N_9028,N_9036,N_9038,N_9040,N_9042,N_9043,N_9044,N_9045,N_9047,N_9049,N_9052,N_9054,N_9055,N_9056,N_9057,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9075,N_9077,N_9080,N_9082,N_9084,N_9085,N_9090,N_9091,N_9093,N_9095,N_9098,N_9099,N_9101,N_9103,N_9104,N_9106,N_9108,N_9109,N_9110,N_9114,N_9116,N_9117,N_9118,N_9119,N_9121,N_9122,N_9123,N_9125,N_9126,N_9127,N_9128,N_9132,N_9134,N_9135,N_9136,N_9139,N_9140,N_9142,N_9143,N_9144,N_9145,N_9148,N_9149,N_9150,N_9155,N_9156,N_9158,N_9159,N_9160,N_9161,N_9162,N_9164,N_9165,N_9167,N_9170,N_9172,N_9174,N_9177,N_9178,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9187,N_9188,N_9189,N_9195,N_9196,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9208,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9219,N_9220,N_9222,N_9223,N_9227,N_9229,N_9230,N_9231,N_9232,N_9235,N_9236,N_9243,N_9244,N_9245,N_9247,N_9249,N_9251,N_9252,N_9253,N_9255,N_9260,N_9261,N_9266,N_9270,N_9273,N_9274,N_9276,N_9281,N_9283,N_9284,N_9285,N_9287,N_9289,N_9290,N_9292,N_9293,N_9294,N_9295,N_9296,N_9298,N_9299,N_9300,N_9301,N_9304,N_9305,N_9306,N_9307,N_9309,N_9311,N_9312,N_9316,N_9318,N_9319,N_9321,N_9324,N_9325,N_9326,N_9328,N_9329,N_9330,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9342,N_9343,N_9345,N_9347,N_9348,N_9349,N_9352,N_9355,N_9357,N_9358,N_9361,N_9364,N_9365,N_9367,N_9369,N_9370,N_9372,N_9374,N_9375,N_9376,N_9377,N_9378,N_9380,N_9381,N_9382,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9391,N_9395,N_9396,N_9397,N_9400,N_9404,N_9406,N_9407,N_9408,N_9409,N_9410,N_9413,N_9415,N_9416,N_9417,N_9418,N_9420,N_9425,N_9426,N_9427,N_9428,N_9429,N_9433,N_9435,N_9436,N_9438,N_9439,N_9440,N_9441,N_9443,N_9446,N_9447,N_9448,N_9452,N_9454,N_9458,N_9459,N_9460,N_9462,N_9467,N_9468,N_9469,N_9471,N_9473,N_9474,N_9476,N_9477,N_9478,N_9480,N_9481,N_9483,N_9484,N_9485,N_9487,N_9488,N_9492,N_9493,N_9494,N_9495,N_9499,N_9500,N_9503,N_9504,N_9505,N_9506,N_9507,N_9510,N_9513,N_9515,N_9516,N_9518,N_9521,N_9524,N_9525,N_9529,N_9531,N_9532,N_9533,N_9535,N_9536,N_9537,N_9538,N_9539,N_9542,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9556,N_9558,N_9560,N_9561,N_9562,N_9563,N_9565,N_9566,N_9567,N_9569,N_9571,N_9572,N_9574,N_9575,N_9578,N_9579,N_9582,N_9585,N_9587,N_9588,N_9590,N_9592,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9604,N_9606,N_9609,N_9612,N_9613,N_9614,N_9615,N_9616,N_9618,N_9620,N_9621,N_9622,N_9623,N_9625,N_9626,N_9627,N_9628,N_9631,N_9633,N_9634,N_9636,N_9642,N_9645,N_9646,N_9648,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9665,N_9666,N_9669,N_9670,N_9671,N_9682,N_9683,N_9684,N_9686,N_9687,N_9688,N_9689,N_9690,N_9692,N_9696,N_9699,N_9702,N_9703,N_9706,N_9707,N_9708,N_9709,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9721,N_9722,N_9724,N_9725,N_9729,N_9731,N_9733,N_9734,N_9735,N_9737,N_9738,N_9739,N_9742,N_9743,N_9744,N_9745,N_9748,N_9750,N_9751,N_9752,N_9753,N_9754,N_9758,N_9760,N_9761,N_9762,N_9763,N_9766,N_9768,N_9771,N_9772,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9782,N_9784,N_9786,N_9787,N_9790,N_9791,N_9792,N_9793,N_9795,N_9796,N_9797,N_9801,N_9803,N_9805,N_9806,N_9808,N_9809,N_9810,N_9811,N_9812,N_9814,N_9818,N_9821,N_9824,N_9825,N_9826,N_9829,N_9833,N_9834,N_9835,N_9836,N_9837,N_9839,N_9841,N_9842,N_9847,N_9848,N_9850,N_9852,N_9854,N_9855,N_9856,N_9858,N_9859,N_9861,N_9863,N_9864,N_9865,N_9867,N_9869,N_9870,N_9871,N_9872,N_9874,N_9875,N_9878,N_9879,N_9880,N_9886,N_9888,N_9889,N_9893,N_9894,N_9895,N_9896,N_9900,N_9903,N_9904,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9922,N_9923,N_9924,N_9929,N_9930,N_9931,N_9933,N_9934,N_9936,N_9938,N_9939,N_9940,N_9941,N_9942,N_9944,N_9945,N_9946,N_9947,N_9949,N_9950,N_9951,N_9953,N_9955,N_9959,N_9960,N_9961,N_9963,N_9964,N_9966,N_9968,N_9969,N_9971,N_9972,N_9974,N_9975,N_9976,N_9978,N_9979,N_9982,N_9983,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9993,N_9994,N_9998;
or U0 (N_0,In_68,In_866);
nand U1 (N_1,In_895,In_81);
xnor U2 (N_2,In_847,In_452);
nand U3 (N_3,In_231,In_518);
or U4 (N_4,In_929,In_900);
and U5 (N_5,In_152,In_430);
or U6 (N_6,In_826,In_100);
xnor U7 (N_7,In_611,In_647);
and U8 (N_8,In_379,In_437);
nand U9 (N_9,In_519,In_709);
or U10 (N_10,In_771,In_115);
nand U11 (N_11,In_477,In_793);
nand U12 (N_12,In_787,In_760);
and U13 (N_13,In_59,In_982);
and U14 (N_14,In_275,In_288);
or U15 (N_15,In_359,In_96);
nand U16 (N_16,In_914,In_448);
nand U17 (N_17,In_988,In_620);
and U18 (N_18,In_216,In_223);
nor U19 (N_19,In_892,In_204);
or U20 (N_20,In_72,In_487);
nand U21 (N_21,In_101,In_978);
or U22 (N_22,In_915,In_11);
nand U23 (N_23,In_292,In_874);
or U24 (N_24,In_489,In_88);
or U25 (N_25,In_175,In_530);
or U26 (N_26,In_859,In_956);
or U27 (N_27,In_698,In_786);
or U28 (N_28,In_187,In_837);
nand U29 (N_29,In_262,In_751);
nor U30 (N_30,In_381,In_280);
and U31 (N_31,In_741,In_964);
nand U32 (N_32,In_896,In_527);
or U33 (N_33,In_344,In_375);
or U34 (N_34,In_372,In_229);
and U35 (N_35,In_350,In_236);
nor U36 (N_36,In_774,In_0);
nor U37 (N_37,In_614,In_319);
nand U38 (N_38,In_93,In_693);
nand U39 (N_39,In_123,In_605);
nand U40 (N_40,In_161,In_177);
nor U41 (N_41,In_97,In_150);
nor U42 (N_42,In_443,In_290);
or U43 (N_43,In_742,In_120);
nand U44 (N_44,In_640,In_606);
nand U45 (N_45,In_248,In_271);
nor U46 (N_46,In_706,In_705);
nand U47 (N_47,In_545,In_746);
and U48 (N_48,In_572,In_190);
or U49 (N_49,In_540,In_788);
nand U50 (N_50,In_828,In_314);
xor U51 (N_51,In_308,In_525);
nor U52 (N_52,In_172,In_493);
nand U53 (N_53,In_71,In_549);
or U54 (N_54,In_266,In_778);
and U55 (N_55,In_708,In_352);
and U56 (N_56,In_596,In_599);
or U57 (N_57,In_414,In_383);
and U58 (N_58,In_580,In_591);
and U59 (N_59,In_146,In_64);
and U60 (N_60,In_12,In_848);
and U61 (N_61,In_125,In_282);
and U62 (N_62,In_846,In_878);
and U63 (N_63,In_163,In_176);
nor U64 (N_64,In_702,In_776);
nand U65 (N_65,In_536,In_75);
or U66 (N_66,In_70,In_348);
nor U67 (N_67,In_257,In_780);
nor U68 (N_68,In_717,In_634);
nor U69 (N_69,In_641,In_977);
or U70 (N_70,In_528,In_789);
nand U71 (N_71,In_650,In_14);
or U72 (N_72,In_601,In_940);
and U73 (N_73,In_22,In_950);
or U74 (N_74,In_646,In_357);
and U75 (N_75,In_110,In_853);
and U76 (N_76,In_965,In_585);
nor U77 (N_77,In_105,In_212);
and U78 (N_78,In_809,In_631);
nand U79 (N_79,In_36,In_905);
or U80 (N_80,In_712,In_30);
nand U81 (N_81,In_178,In_356);
nand U82 (N_82,In_845,In_241);
nor U83 (N_83,In_703,In_474);
nand U84 (N_84,In_73,In_365);
nand U85 (N_85,In_390,In_199);
nand U86 (N_86,In_391,In_668);
nand U87 (N_87,In_407,In_523);
nand U88 (N_88,In_332,In_636);
or U89 (N_89,In_941,In_34);
xor U90 (N_90,In_612,In_880);
nor U91 (N_91,In_336,In_65);
nor U92 (N_92,In_841,In_743);
nand U93 (N_93,In_728,In_856);
nor U94 (N_94,In_830,In_191);
nand U95 (N_95,In_87,In_274);
nor U96 (N_96,In_174,In_304);
or U97 (N_97,In_975,In_261);
nor U98 (N_98,In_948,In_165);
and U99 (N_99,In_425,In_171);
nor U100 (N_100,In_169,In_4);
and U101 (N_101,In_618,In_796);
or U102 (N_102,In_427,In_339);
nand U103 (N_103,In_898,In_461);
or U104 (N_104,In_683,In_39);
nor U105 (N_105,In_497,In_755);
or U106 (N_106,In_426,In_83);
or U107 (N_107,In_483,In_695);
nor U108 (N_108,In_974,In_863);
nand U109 (N_109,In_6,In_394);
nand U110 (N_110,In_299,In_450);
nand U111 (N_111,In_667,In_464);
nand U112 (N_112,In_347,In_817);
and U113 (N_113,In_727,In_358);
nand U114 (N_114,In_921,In_936);
nand U115 (N_115,In_648,In_400);
or U116 (N_116,In_13,In_607);
or U117 (N_117,In_769,In_27);
and U118 (N_118,In_168,In_864);
or U119 (N_119,In_360,In_302);
and U120 (N_120,In_860,In_423);
and U121 (N_121,In_315,In_925);
nand U122 (N_122,In_707,In_806);
nand U123 (N_123,In_902,In_484);
or U124 (N_124,In_587,In_522);
or U125 (N_125,In_663,In_716);
and U126 (N_126,In_259,In_584);
and U127 (N_127,In_680,In_367);
or U128 (N_128,In_321,In_958);
nand U129 (N_129,In_901,In_132);
or U130 (N_130,In_444,In_328);
and U131 (N_131,In_313,In_193);
nand U132 (N_132,In_777,In_721);
nor U133 (N_133,In_267,In_504);
xor U134 (N_134,In_691,In_408);
and U135 (N_135,In_598,In_481);
nor U136 (N_136,In_480,In_291);
nand U137 (N_137,In_277,In_84);
nor U138 (N_138,In_23,In_496);
nand U139 (N_139,In_111,In_127);
nand U140 (N_140,In_671,In_364);
xor U141 (N_141,In_201,In_836);
and U142 (N_142,In_340,In_939);
nor U143 (N_143,In_143,In_135);
nor U144 (N_144,In_129,In_827);
nand U145 (N_145,In_731,In_581);
nand U146 (N_146,In_722,In_569);
or U147 (N_147,In_38,In_972);
or U148 (N_148,In_305,In_815);
nor U149 (N_149,In_920,In_969);
nand U150 (N_150,In_109,In_342);
nor U151 (N_151,In_719,In_345);
xnor U152 (N_152,In_872,In_289);
nor U153 (N_153,In_215,In_593);
or U154 (N_154,In_749,In_933);
nand U155 (N_155,In_453,In_862);
xnor U156 (N_156,In_382,In_657);
or U157 (N_157,In_696,In_486);
nor U158 (N_158,In_724,In_419);
and U159 (N_159,In_151,In_625);
nand U160 (N_160,In_962,In_66);
or U161 (N_161,In_903,In_102);
and U162 (N_162,In_211,In_52);
and U163 (N_163,In_104,In_816);
nand U164 (N_164,In_779,In_882);
or U165 (N_165,In_674,In_48);
or U166 (N_166,In_369,In_77);
or U167 (N_167,In_44,In_960);
nand U168 (N_168,In_928,In_740);
nor U169 (N_169,In_516,In_871);
and U170 (N_170,In_296,In_517);
nand U171 (N_171,In_462,In_773);
nor U172 (N_172,In_227,In_553);
nand U173 (N_173,In_78,In_783);
nor U174 (N_174,In_819,In_476);
nor U175 (N_175,In_456,In_718);
and U176 (N_176,In_368,In_149);
and U177 (N_177,In_660,In_7);
or U178 (N_178,In_986,In_181);
and U179 (N_179,In_467,In_952);
nor U180 (N_180,In_715,In_922);
nand U181 (N_181,In_362,In_566);
or U182 (N_182,In_185,In_739);
and U183 (N_183,In_554,In_655);
nor U184 (N_184,In_239,In_337);
and U185 (N_185,In_258,In_684);
nand U186 (N_186,In_567,In_28);
or U187 (N_187,In_268,In_658);
or U188 (N_188,In_438,In_329);
nor U189 (N_189,In_147,In_548);
or U190 (N_190,In_403,In_694);
or U191 (N_191,In_335,In_432);
or U192 (N_192,In_55,In_158);
nand U193 (N_193,In_665,In_785);
nand U194 (N_194,In_85,In_162);
nor U195 (N_195,In_550,In_881);
or U196 (N_196,In_574,In_270);
and U197 (N_197,In_353,In_888);
nand U198 (N_198,In_173,In_953);
nand U199 (N_199,In_745,In_117);
and U200 (N_200,In_220,In_632);
nand U201 (N_201,In_10,In_961);
and U202 (N_202,In_124,In_492);
or U203 (N_203,In_752,In_679);
nand U204 (N_204,In_385,In_249);
and U205 (N_205,In_659,In_160);
nand U206 (N_206,In_15,In_202);
nor U207 (N_207,In_384,In_306);
nor U208 (N_208,In_8,In_226);
nor U209 (N_209,In_389,In_831);
nand U210 (N_210,In_5,In_170);
nand U211 (N_211,In_327,In_439);
nand U212 (N_212,In_479,In_116);
or U213 (N_213,In_812,In_472);
or U214 (N_214,In_370,In_959);
nor U215 (N_215,In_992,In_681);
and U216 (N_216,In_908,In_897);
and U217 (N_217,In_310,In_113);
nor U218 (N_218,In_945,In_583);
nand U219 (N_219,In_546,In_466);
nor U220 (N_220,In_565,In_990);
or U221 (N_221,In_894,In_429);
and U222 (N_222,In_912,In_676);
or U223 (N_223,In_51,In_562);
nand U224 (N_224,In_393,In_511);
nor U225 (N_225,In_577,In_373);
and U226 (N_226,In_985,In_738);
nand U227 (N_227,In_954,In_653);
or U228 (N_228,In_157,In_515);
nor U229 (N_229,In_74,In_850);
and U230 (N_230,In_732,In_852);
nor U231 (N_231,In_203,In_944);
nor U232 (N_232,In_320,In_782);
xnor U233 (N_233,In_592,In_509);
or U234 (N_234,In_207,In_142);
nor U235 (N_235,In_630,In_943);
and U236 (N_236,In_946,In_402);
or U237 (N_237,In_445,In_573);
and U238 (N_238,In_285,In_750);
nor U239 (N_239,In_700,In_436);
nor U240 (N_240,In_33,In_757);
nor U241 (N_241,In_713,In_338);
nor U242 (N_242,In_813,In_240);
nor U243 (N_243,In_699,In_798);
or U244 (N_244,In_851,In_194);
nand U245 (N_245,In_298,In_279);
or U246 (N_246,In_595,In_794);
nor U247 (N_247,In_558,In_198);
or U248 (N_248,In_995,In_451);
or U249 (N_249,In_494,In_322);
nor U250 (N_250,In_392,In_899);
nand U251 (N_251,In_60,In_19);
and U252 (N_252,In_455,In_119);
nand U253 (N_253,In_281,In_76);
nor U254 (N_254,In_735,In_366);
nor U255 (N_255,In_21,In_167);
or U256 (N_256,In_440,In_513);
and U257 (N_257,In_876,In_86);
or U258 (N_258,In_447,In_253);
and U259 (N_259,In_122,In_53);
and U260 (N_260,In_287,In_99);
and U261 (N_261,In_799,In_682);
nand U262 (N_262,In_238,In_206);
and U263 (N_263,In_797,In_537);
nor U264 (N_264,In_508,In_927);
nor U265 (N_265,In_300,In_998);
and U266 (N_266,In_415,In_690);
and U267 (N_267,In_269,In_459);
nor U268 (N_268,In_371,In_58);
and U269 (N_269,In_886,In_649);
and U270 (N_270,In_931,In_301);
and U271 (N_271,In_879,In_406);
and U272 (N_272,In_622,In_156);
and U273 (N_273,In_250,In_685);
nand U274 (N_274,In_865,In_870);
nor U275 (N_275,In_463,In_688);
and U276 (N_276,In_904,In_910);
and U277 (N_277,In_571,In_210);
and U278 (N_278,In_16,In_832);
nand U279 (N_279,In_552,In_615);
or U280 (N_280,In_811,In_95);
nor U281 (N_281,In_748,In_916);
nand U282 (N_282,In_645,In_80);
and U283 (N_283,In_997,In_222);
nand U284 (N_284,In_840,In_488);
or U285 (N_285,In_137,In_254);
nand U286 (N_286,In_526,In_531);
nor U287 (N_287,In_768,In_417);
nand U288 (N_288,In_376,In_795);
nor U289 (N_289,In_90,In_63);
nor U290 (N_290,In_485,In_465);
nor U291 (N_291,In_535,In_473);
and U292 (N_292,In_906,In_514);
nand U293 (N_293,In_764,In_503);
or U294 (N_294,In_891,In_600);
nor U295 (N_295,In_114,In_138);
xor U296 (N_296,In_854,In_624);
nand U297 (N_297,In_714,In_767);
or U298 (N_298,In_808,In_121);
or U299 (N_299,In_112,In_45);
or U300 (N_300,In_909,In_334);
and U301 (N_301,In_924,In_805);
or U302 (N_302,In_885,In_243);
nand U303 (N_303,In_661,In_29);
nor U304 (N_304,In_790,In_18);
nand U305 (N_305,In_237,In_541);
or U306 (N_306,In_633,In_524);
and U307 (N_307,In_482,In_993);
or U308 (N_308,In_999,In_295);
or U309 (N_309,In_802,In_454);
nand U310 (N_310,In_186,In_803);
nor U311 (N_311,In_723,In_92);
nand U312 (N_312,In_506,In_582);
nor U313 (N_313,In_857,In_31);
and U314 (N_314,In_967,In_505);
nand U315 (N_315,In_822,In_701);
nor U316 (N_316,In_981,In_228);
nor U317 (N_317,In_801,In_765);
and U318 (N_318,In_205,In_568);
or U319 (N_319,In_26,In_861);
and U320 (N_320,In_140,In_420);
nor U321 (N_321,In_907,In_677);
nor U322 (N_322,In_603,In_499);
nand U323 (N_323,In_635,In_844);
nand U324 (N_324,In_729,In_136);
nor U325 (N_325,In_433,In_208);
nand U326 (N_326,In_25,In_197);
or U327 (N_327,In_468,In_772);
and U328 (N_328,In_232,In_976);
nor U329 (N_329,In_182,In_838);
nor U330 (N_330,In_361,In_814);
and U331 (N_331,In_643,In_734);
nor U332 (N_332,In_937,In_996);
or U333 (N_333,In_260,In_244);
and U334 (N_334,In_297,In_20);
nor U335 (N_335,In_617,In_687);
nor U336 (N_336,In_286,In_781);
nor U337 (N_337,In_994,In_627);
and U338 (N_338,In_255,In_597);
or U339 (N_339,In_930,In_242);
nor U340 (N_340,In_639,In_756);
or U341 (N_341,In_890,In_1);
nand U342 (N_342,In_159,In_619);
nor U343 (N_343,In_884,In_230);
nor U344 (N_344,In_987,In_89);
or U345 (N_345,In_824,In_820);
or U346 (N_346,In_602,In_678);
nand U347 (N_347,In_98,In_221);
nand U348 (N_348,In_542,In_460);
or U349 (N_349,In_307,In_533);
nor U350 (N_350,In_67,In_457);
nand U351 (N_351,In_932,In_179);
nor U352 (N_352,In_926,In_642);
nor U353 (N_353,In_442,In_623);
and U354 (N_354,In_428,In_521);
and U355 (N_355,In_79,In_821);
and U356 (N_356,In_733,In_935);
or U357 (N_357,In_118,In_919);
and U358 (N_358,In_410,In_47);
and U359 (N_359,In_189,In_24);
nand U360 (N_360,In_766,In_252);
nand U361 (N_361,In_209,In_942);
nor U362 (N_362,In_225,In_911);
nand U363 (N_363,In_791,In_747);
or U364 (N_364,In_673,In_672);
nand U365 (N_365,In_61,In_247);
nor U366 (N_366,In_418,In_610);
and U367 (N_367,In_923,In_955);
nor U368 (N_368,In_164,In_388);
and U369 (N_369,In_57,In_246);
nand U370 (N_370,In_134,In_758);
nand U371 (N_371,In_431,In_534);
or U372 (N_372,In_458,In_744);
or U373 (N_373,In_991,In_106);
nand U374 (N_374,In_501,In_883);
or U375 (N_375,In_303,In_133);
nor U376 (N_376,In_435,In_251);
nand U377 (N_377,In_273,In_256);
or U378 (N_378,In_82,In_213);
nor U379 (N_379,In_726,In_3);
and U380 (N_380,In_405,In_730);
nor U381 (N_381,In_317,In_689);
and U382 (N_382,In_155,In_711);
nand U383 (N_383,In_842,In_323);
nand U384 (N_384,In_214,In_126);
nor U385 (N_385,In_355,In_833);
nand U386 (N_386,In_529,In_825);
or U387 (N_387,In_62,In_792);
nor U388 (N_388,In_478,In_154);
nor U389 (N_389,In_35,In_153);
nor U390 (N_390,In_983,In_800);
or U391 (N_391,In_559,In_654);
nor U392 (N_392,In_588,In_346);
nand U393 (N_393,In_543,In_720);
and U394 (N_394,In_500,In_692);
or U395 (N_395,In_867,In_770);
and U396 (N_396,In_575,In_103);
nor U397 (N_397,In_675,In_374);
nor U398 (N_398,In_564,In_416);
or U399 (N_399,In_264,In_495);
or U400 (N_400,In_265,In_188);
or U401 (N_401,In_128,In_763);
nand U402 (N_402,In_539,In_318);
nor U403 (N_403,In_412,In_823);
nand U404 (N_404,In_293,In_475);
nor U405 (N_405,In_9,In_396);
nor U406 (N_406,In_563,In_446);
nor U407 (N_407,In_148,In_325);
or U408 (N_408,In_520,In_354);
or U409 (N_409,In_507,In_245);
or U410 (N_410,In_272,In_377);
nand U411 (N_411,In_887,In_424);
nor U412 (N_412,In_670,In_704);
nand U413 (N_413,In_590,In_918);
and U414 (N_414,In_775,In_17);
and U415 (N_415,In_512,In_386);
nand U416 (N_416,In_666,In_387);
and U417 (N_417,In_980,In_604);
and U418 (N_418,In_873,In_609);
or U419 (N_419,In_637,In_651);
nor U420 (N_420,In_869,In_311);
nand U421 (N_421,In_312,In_107);
or U422 (N_422,In_725,In_608);
nor U423 (N_423,In_470,In_557);
nand U424 (N_424,In_855,In_192);
nor U425 (N_425,In_341,In_54);
xor U426 (N_426,In_141,In_973);
or U427 (N_427,In_434,In_947);
nor U428 (N_428,In_233,In_235);
or U429 (N_429,In_875,In_490);
and U430 (N_430,In_139,In_380);
or U431 (N_431,In_195,In_56);
nand U432 (N_432,In_638,In_839);
nand U433 (N_433,In_218,In_395);
nor U434 (N_434,In_398,In_889);
xnor U435 (N_435,In_399,In_551);
nand U436 (N_436,In_807,In_594);
nor U437 (N_437,In_37,In_877);
nand U438 (N_438,In_41,In_131);
or U439 (N_439,In_510,In_555);
or U440 (N_440,In_989,In_32);
nor U441 (N_441,In_586,In_351);
nor U442 (N_442,In_629,In_378);
and U443 (N_443,In_951,In_91);
nand U444 (N_444,In_411,In_621);
nand U445 (N_445,In_224,In_697);
or U446 (N_446,In_656,In_938);
nor U447 (N_447,In_363,In_686);
nand U448 (N_448,In_589,In_868);
nand U449 (N_449,In_810,In_849);
and U450 (N_450,In_560,In_50);
or U451 (N_451,In_234,In_471);
and U452 (N_452,In_759,In_710);
or U453 (N_453,In_979,In_284);
nand U454 (N_454,In_217,In_968);
nand U455 (N_455,In_893,In_2);
nor U456 (N_456,In_421,In_949);
nand U457 (N_457,In_491,In_184);
or U458 (N_458,In_200,In_196);
nand U459 (N_459,In_349,In_219);
or U460 (N_460,In_422,In_180);
nand U461 (N_461,In_616,In_469);
and U462 (N_462,In_934,In_449);
nand U463 (N_463,In_835,In_324);
and U464 (N_464,In_834,In_761);
xor U465 (N_465,In_544,In_43);
or U466 (N_466,In_736,In_613);
and U467 (N_467,In_46,In_644);
and U468 (N_468,In_578,In_49);
nor U469 (N_469,In_263,In_538);
nand U470 (N_470,In_628,In_397);
or U471 (N_471,In_753,In_957);
nand U472 (N_472,In_829,In_130);
and U473 (N_473,In_94,In_669);
nor U474 (N_474,In_970,In_754);
nor U475 (N_475,In_183,In_843);
nor U476 (N_476,In_664,In_42);
nor U477 (N_477,In_278,In_108);
or U478 (N_478,In_413,In_333);
or U479 (N_479,In_309,In_294);
nand U480 (N_480,In_917,In_662);
and U481 (N_481,In_626,In_326);
nand U482 (N_482,In_316,In_570);
and U483 (N_483,In_401,In_547);
or U484 (N_484,In_144,In_331);
or U485 (N_485,In_784,In_971);
or U486 (N_486,In_556,In_409);
and U487 (N_487,In_69,In_166);
or U488 (N_488,In_913,In_576);
nor U489 (N_489,In_283,In_579);
or U490 (N_490,In_966,In_40);
or U491 (N_491,In_498,In_804);
nor U492 (N_492,In_561,In_502);
and U493 (N_493,In_984,In_858);
nand U494 (N_494,In_145,In_532);
or U495 (N_495,In_343,In_818);
nor U496 (N_496,In_441,In_404);
nand U497 (N_497,In_737,In_652);
or U498 (N_498,In_762,In_330);
nor U499 (N_499,In_963,In_276);
nand U500 (N_500,In_46,In_313);
and U501 (N_501,In_417,In_948);
nor U502 (N_502,In_334,In_903);
xnor U503 (N_503,In_664,In_947);
and U504 (N_504,In_999,In_686);
nand U505 (N_505,In_500,In_290);
nor U506 (N_506,In_206,In_957);
or U507 (N_507,In_199,In_222);
or U508 (N_508,In_338,In_561);
nor U509 (N_509,In_152,In_493);
or U510 (N_510,In_484,In_782);
nor U511 (N_511,In_644,In_517);
nor U512 (N_512,In_529,In_937);
and U513 (N_513,In_471,In_790);
and U514 (N_514,In_355,In_470);
and U515 (N_515,In_344,In_930);
or U516 (N_516,In_447,In_48);
nand U517 (N_517,In_664,In_192);
nor U518 (N_518,In_977,In_104);
or U519 (N_519,In_953,In_554);
nor U520 (N_520,In_409,In_633);
nand U521 (N_521,In_789,In_47);
or U522 (N_522,In_802,In_218);
nor U523 (N_523,In_418,In_752);
and U524 (N_524,In_446,In_539);
xnor U525 (N_525,In_241,In_383);
or U526 (N_526,In_89,In_795);
and U527 (N_527,In_761,In_858);
nand U528 (N_528,In_154,In_893);
nand U529 (N_529,In_788,In_720);
xnor U530 (N_530,In_909,In_728);
and U531 (N_531,In_2,In_673);
nor U532 (N_532,In_853,In_233);
or U533 (N_533,In_524,In_637);
and U534 (N_534,In_614,In_103);
and U535 (N_535,In_438,In_503);
nand U536 (N_536,In_354,In_414);
nand U537 (N_537,In_815,In_871);
and U538 (N_538,In_367,In_912);
and U539 (N_539,In_618,In_762);
or U540 (N_540,In_680,In_432);
or U541 (N_541,In_554,In_543);
and U542 (N_542,In_619,In_817);
and U543 (N_543,In_98,In_359);
nor U544 (N_544,In_737,In_430);
nand U545 (N_545,In_385,In_21);
nand U546 (N_546,In_977,In_296);
nand U547 (N_547,In_514,In_316);
or U548 (N_548,In_698,In_425);
nor U549 (N_549,In_763,In_586);
nor U550 (N_550,In_640,In_497);
or U551 (N_551,In_326,In_938);
nand U552 (N_552,In_169,In_714);
or U553 (N_553,In_475,In_899);
and U554 (N_554,In_61,In_676);
and U555 (N_555,In_890,In_539);
or U556 (N_556,In_348,In_106);
and U557 (N_557,In_809,In_509);
and U558 (N_558,In_886,In_35);
nand U559 (N_559,In_452,In_53);
nor U560 (N_560,In_245,In_703);
or U561 (N_561,In_736,In_827);
nand U562 (N_562,In_350,In_176);
nor U563 (N_563,In_752,In_535);
or U564 (N_564,In_618,In_600);
nand U565 (N_565,In_319,In_119);
nor U566 (N_566,In_411,In_739);
nor U567 (N_567,In_341,In_69);
nor U568 (N_568,In_659,In_287);
or U569 (N_569,In_610,In_999);
or U570 (N_570,In_38,In_757);
nor U571 (N_571,In_607,In_545);
or U572 (N_572,In_81,In_723);
nand U573 (N_573,In_153,In_619);
or U574 (N_574,In_437,In_45);
nand U575 (N_575,In_840,In_562);
or U576 (N_576,In_434,In_32);
nor U577 (N_577,In_805,In_117);
or U578 (N_578,In_112,In_760);
or U579 (N_579,In_364,In_416);
nand U580 (N_580,In_455,In_421);
xor U581 (N_581,In_42,In_258);
nor U582 (N_582,In_946,In_400);
and U583 (N_583,In_907,In_494);
or U584 (N_584,In_42,In_13);
nand U585 (N_585,In_341,In_314);
nor U586 (N_586,In_88,In_962);
nor U587 (N_587,In_576,In_971);
nand U588 (N_588,In_831,In_563);
nor U589 (N_589,In_105,In_644);
nand U590 (N_590,In_751,In_159);
nand U591 (N_591,In_477,In_121);
nand U592 (N_592,In_280,In_158);
nor U593 (N_593,In_608,In_908);
nand U594 (N_594,In_576,In_392);
and U595 (N_595,In_456,In_133);
nand U596 (N_596,In_927,In_73);
nand U597 (N_597,In_787,In_582);
or U598 (N_598,In_391,In_102);
nand U599 (N_599,In_481,In_432);
or U600 (N_600,In_866,In_351);
nand U601 (N_601,In_157,In_507);
nor U602 (N_602,In_281,In_642);
or U603 (N_603,In_167,In_650);
or U604 (N_604,In_493,In_177);
and U605 (N_605,In_940,In_579);
or U606 (N_606,In_241,In_174);
nor U607 (N_607,In_433,In_653);
or U608 (N_608,In_783,In_715);
nand U609 (N_609,In_406,In_802);
or U610 (N_610,In_644,In_801);
nand U611 (N_611,In_753,In_178);
nand U612 (N_612,In_590,In_172);
nor U613 (N_613,In_390,In_352);
nand U614 (N_614,In_977,In_156);
nand U615 (N_615,In_121,In_23);
or U616 (N_616,In_821,In_705);
nand U617 (N_617,In_205,In_734);
or U618 (N_618,In_596,In_123);
nand U619 (N_619,In_250,In_371);
or U620 (N_620,In_68,In_23);
or U621 (N_621,In_544,In_33);
or U622 (N_622,In_188,In_844);
or U623 (N_623,In_417,In_692);
and U624 (N_624,In_402,In_39);
nor U625 (N_625,In_717,In_59);
and U626 (N_626,In_795,In_199);
and U627 (N_627,In_497,In_203);
or U628 (N_628,In_467,In_377);
or U629 (N_629,In_422,In_234);
or U630 (N_630,In_469,In_583);
nor U631 (N_631,In_199,In_422);
nand U632 (N_632,In_282,In_716);
or U633 (N_633,In_63,In_265);
nand U634 (N_634,In_784,In_581);
and U635 (N_635,In_319,In_547);
and U636 (N_636,In_399,In_921);
nor U637 (N_637,In_757,In_968);
and U638 (N_638,In_101,In_120);
nand U639 (N_639,In_924,In_432);
nor U640 (N_640,In_644,In_316);
and U641 (N_641,In_261,In_116);
nand U642 (N_642,In_443,In_306);
nand U643 (N_643,In_810,In_38);
nor U644 (N_644,In_840,In_251);
nor U645 (N_645,In_277,In_947);
nor U646 (N_646,In_177,In_39);
or U647 (N_647,In_224,In_790);
nand U648 (N_648,In_582,In_358);
nor U649 (N_649,In_670,In_492);
nor U650 (N_650,In_243,In_387);
and U651 (N_651,In_662,In_205);
nor U652 (N_652,In_889,In_874);
nand U653 (N_653,In_203,In_811);
or U654 (N_654,In_851,In_162);
or U655 (N_655,In_973,In_13);
or U656 (N_656,In_613,In_207);
or U657 (N_657,In_597,In_76);
nor U658 (N_658,In_760,In_266);
nor U659 (N_659,In_946,In_451);
nand U660 (N_660,In_845,In_475);
nor U661 (N_661,In_882,In_902);
nand U662 (N_662,In_313,In_924);
nand U663 (N_663,In_670,In_569);
nand U664 (N_664,In_604,In_492);
nor U665 (N_665,In_927,In_370);
and U666 (N_666,In_22,In_803);
or U667 (N_667,In_569,In_926);
xnor U668 (N_668,In_414,In_112);
nand U669 (N_669,In_47,In_865);
and U670 (N_670,In_473,In_716);
and U671 (N_671,In_258,In_30);
nand U672 (N_672,In_939,In_322);
or U673 (N_673,In_932,In_471);
and U674 (N_674,In_640,In_56);
nor U675 (N_675,In_990,In_44);
and U676 (N_676,In_998,In_573);
nor U677 (N_677,In_778,In_641);
and U678 (N_678,In_642,In_223);
nor U679 (N_679,In_150,In_52);
nor U680 (N_680,In_915,In_781);
nand U681 (N_681,In_212,In_312);
nand U682 (N_682,In_54,In_537);
nor U683 (N_683,In_868,In_45);
nand U684 (N_684,In_119,In_947);
nand U685 (N_685,In_88,In_660);
nor U686 (N_686,In_689,In_651);
nand U687 (N_687,In_421,In_238);
nor U688 (N_688,In_84,In_671);
and U689 (N_689,In_537,In_204);
and U690 (N_690,In_662,In_293);
nand U691 (N_691,In_89,In_48);
or U692 (N_692,In_290,In_888);
nor U693 (N_693,In_78,In_330);
xnor U694 (N_694,In_733,In_453);
nor U695 (N_695,In_710,In_135);
or U696 (N_696,In_946,In_749);
or U697 (N_697,In_566,In_499);
nor U698 (N_698,In_648,In_89);
nand U699 (N_699,In_416,In_576);
nor U700 (N_700,In_233,In_526);
or U701 (N_701,In_401,In_693);
nand U702 (N_702,In_631,In_348);
nor U703 (N_703,In_343,In_44);
nor U704 (N_704,In_72,In_512);
or U705 (N_705,In_422,In_740);
and U706 (N_706,In_383,In_168);
nor U707 (N_707,In_910,In_392);
or U708 (N_708,In_275,In_56);
nand U709 (N_709,In_35,In_96);
nand U710 (N_710,In_339,In_852);
nor U711 (N_711,In_208,In_903);
and U712 (N_712,In_331,In_786);
and U713 (N_713,In_622,In_116);
and U714 (N_714,In_81,In_463);
or U715 (N_715,In_596,In_661);
and U716 (N_716,In_747,In_814);
and U717 (N_717,In_502,In_856);
xnor U718 (N_718,In_209,In_259);
or U719 (N_719,In_811,In_358);
and U720 (N_720,In_204,In_167);
and U721 (N_721,In_633,In_228);
and U722 (N_722,In_713,In_987);
or U723 (N_723,In_844,In_541);
and U724 (N_724,In_807,In_133);
and U725 (N_725,In_2,In_454);
and U726 (N_726,In_854,In_782);
and U727 (N_727,In_43,In_181);
or U728 (N_728,In_788,In_970);
or U729 (N_729,In_417,In_5);
nor U730 (N_730,In_293,In_552);
nand U731 (N_731,In_635,In_339);
nor U732 (N_732,In_846,In_235);
and U733 (N_733,In_450,In_776);
and U734 (N_734,In_872,In_831);
nand U735 (N_735,In_940,In_202);
nor U736 (N_736,In_179,In_275);
or U737 (N_737,In_708,In_65);
or U738 (N_738,In_134,In_879);
nand U739 (N_739,In_657,In_546);
and U740 (N_740,In_660,In_786);
nor U741 (N_741,In_754,In_60);
and U742 (N_742,In_491,In_418);
nand U743 (N_743,In_177,In_632);
or U744 (N_744,In_529,In_856);
nand U745 (N_745,In_832,In_730);
nor U746 (N_746,In_645,In_79);
nor U747 (N_747,In_944,In_736);
and U748 (N_748,In_933,In_754);
nand U749 (N_749,In_835,In_831);
nand U750 (N_750,In_936,In_753);
nand U751 (N_751,In_482,In_269);
or U752 (N_752,In_821,In_508);
or U753 (N_753,In_231,In_597);
and U754 (N_754,In_833,In_531);
nand U755 (N_755,In_156,In_337);
nor U756 (N_756,In_771,In_418);
nand U757 (N_757,In_908,In_366);
nor U758 (N_758,In_522,In_59);
or U759 (N_759,In_439,In_849);
and U760 (N_760,In_16,In_969);
or U761 (N_761,In_942,In_717);
nand U762 (N_762,In_713,In_512);
and U763 (N_763,In_863,In_870);
nand U764 (N_764,In_396,In_487);
or U765 (N_765,In_791,In_868);
nor U766 (N_766,In_323,In_203);
nand U767 (N_767,In_785,In_279);
and U768 (N_768,In_249,In_581);
or U769 (N_769,In_956,In_403);
and U770 (N_770,In_906,In_35);
nor U771 (N_771,In_618,In_133);
nor U772 (N_772,In_564,In_959);
or U773 (N_773,In_33,In_860);
or U774 (N_774,In_452,In_222);
nand U775 (N_775,In_644,In_920);
nor U776 (N_776,In_834,In_469);
and U777 (N_777,In_471,In_636);
and U778 (N_778,In_312,In_296);
or U779 (N_779,In_815,In_661);
nor U780 (N_780,In_955,In_338);
and U781 (N_781,In_756,In_114);
or U782 (N_782,In_974,In_796);
and U783 (N_783,In_865,In_872);
nor U784 (N_784,In_13,In_338);
nor U785 (N_785,In_376,In_766);
nor U786 (N_786,In_861,In_189);
nor U787 (N_787,In_429,In_480);
nor U788 (N_788,In_147,In_15);
nor U789 (N_789,In_491,In_954);
and U790 (N_790,In_423,In_488);
nor U791 (N_791,In_58,In_805);
or U792 (N_792,In_357,In_331);
and U793 (N_793,In_801,In_917);
nand U794 (N_794,In_933,In_101);
xnor U795 (N_795,In_831,In_768);
and U796 (N_796,In_390,In_165);
and U797 (N_797,In_326,In_98);
and U798 (N_798,In_22,In_486);
nor U799 (N_799,In_176,In_410);
or U800 (N_800,In_817,In_1);
nand U801 (N_801,In_8,In_603);
and U802 (N_802,In_764,In_788);
nand U803 (N_803,In_211,In_157);
or U804 (N_804,In_464,In_274);
nand U805 (N_805,In_147,In_255);
and U806 (N_806,In_574,In_144);
and U807 (N_807,In_933,In_371);
nand U808 (N_808,In_862,In_858);
and U809 (N_809,In_194,In_766);
nor U810 (N_810,In_266,In_645);
or U811 (N_811,In_459,In_813);
and U812 (N_812,In_463,In_97);
or U813 (N_813,In_768,In_936);
xnor U814 (N_814,In_467,In_653);
nand U815 (N_815,In_234,In_646);
nand U816 (N_816,In_970,In_340);
nor U817 (N_817,In_993,In_63);
xnor U818 (N_818,In_790,In_906);
nand U819 (N_819,In_773,In_983);
and U820 (N_820,In_161,In_170);
nand U821 (N_821,In_679,In_534);
and U822 (N_822,In_989,In_691);
or U823 (N_823,In_596,In_519);
xnor U824 (N_824,In_633,In_441);
nand U825 (N_825,In_787,In_20);
nor U826 (N_826,In_610,In_595);
nor U827 (N_827,In_695,In_583);
or U828 (N_828,In_185,In_726);
nand U829 (N_829,In_270,In_438);
xor U830 (N_830,In_788,In_6);
or U831 (N_831,In_778,In_674);
nor U832 (N_832,In_202,In_279);
nand U833 (N_833,In_147,In_339);
nor U834 (N_834,In_397,In_760);
and U835 (N_835,In_595,In_17);
xnor U836 (N_836,In_781,In_649);
nor U837 (N_837,In_121,In_816);
or U838 (N_838,In_243,In_160);
nand U839 (N_839,In_272,In_896);
or U840 (N_840,In_310,In_644);
and U841 (N_841,In_313,In_756);
or U842 (N_842,In_883,In_67);
nand U843 (N_843,In_266,In_318);
and U844 (N_844,In_452,In_175);
nand U845 (N_845,In_615,In_324);
nor U846 (N_846,In_760,In_219);
or U847 (N_847,In_953,In_819);
nand U848 (N_848,In_23,In_970);
and U849 (N_849,In_945,In_960);
or U850 (N_850,In_864,In_611);
nor U851 (N_851,In_147,In_832);
nor U852 (N_852,In_334,In_240);
nor U853 (N_853,In_969,In_734);
nand U854 (N_854,In_716,In_386);
or U855 (N_855,In_313,In_293);
nand U856 (N_856,In_925,In_791);
and U857 (N_857,In_397,In_166);
and U858 (N_858,In_188,In_45);
and U859 (N_859,In_796,In_758);
nor U860 (N_860,In_967,In_880);
or U861 (N_861,In_39,In_398);
nand U862 (N_862,In_378,In_314);
nand U863 (N_863,In_468,In_217);
nor U864 (N_864,In_576,In_578);
nand U865 (N_865,In_501,In_829);
nor U866 (N_866,In_639,In_175);
nand U867 (N_867,In_357,In_386);
nand U868 (N_868,In_514,In_799);
nand U869 (N_869,In_630,In_160);
and U870 (N_870,In_810,In_327);
nand U871 (N_871,In_728,In_183);
nand U872 (N_872,In_445,In_886);
nand U873 (N_873,In_933,In_341);
nand U874 (N_874,In_541,In_283);
and U875 (N_875,In_181,In_930);
nor U876 (N_876,In_458,In_7);
nor U877 (N_877,In_309,In_678);
or U878 (N_878,In_832,In_606);
nor U879 (N_879,In_724,In_702);
and U880 (N_880,In_825,In_813);
nor U881 (N_881,In_416,In_434);
and U882 (N_882,In_772,In_482);
or U883 (N_883,In_795,In_161);
nor U884 (N_884,In_674,In_108);
nor U885 (N_885,In_781,In_773);
nand U886 (N_886,In_524,In_703);
nor U887 (N_887,In_528,In_755);
nor U888 (N_888,In_479,In_547);
or U889 (N_889,In_745,In_672);
and U890 (N_890,In_580,In_854);
nand U891 (N_891,In_409,In_928);
or U892 (N_892,In_95,In_5);
nand U893 (N_893,In_367,In_121);
nor U894 (N_894,In_393,In_201);
nor U895 (N_895,In_247,In_532);
and U896 (N_896,In_515,In_184);
nand U897 (N_897,In_346,In_101);
xnor U898 (N_898,In_390,In_327);
nor U899 (N_899,In_808,In_341);
and U900 (N_900,In_472,In_163);
xor U901 (N_901,In_711,In_691);
or U902 (N_902,In_161,In_23);
nand U903 (N_903,In_832,In_918);
xnor U904 (N_904,In_727,In_951);
or U905 (N_905,In_832,In_622);
or U906 (N_906,In_162,In_888);
xnor U907 (N_907,In_126,In_354);
nor U908 (N_908,In_435,In_936);
and U909 (N_909,In_921,In_948);
and U910 (N_910,In_52,In_709);
and U911 (N_911,In_594,In_26);
and U912 (N_912,In_933,In_840);
or U913 (N_913,In_677,In_781);
and U914 (N_914,In_19,In_612);
nand U915 (N_915,In_301,In_980);
nor U916 (N_916,In_468,In_124);
nor U917 (N_917,In_710,In_128);
nor U918 (N_918,In_678,In_443);
or U919 (N_919,In_270,In_366);
nand U920 (N_920,In_239,In_555);
nand U921 (N_921,In_807,In_739);
or U922 (N_922,In_853,In_102);
nor U923 (N_923,In_356,In_63);
nor U924 (N_924,In_365,In_500);
nand U925 (N_925,In_189,In_507);
or U926 (N_926,In_733,In_330);
nand U927 (N_927,In_293,In_192);
or U928 (N_928,In_344,In_209);
nand U929 (N_929,In_84,In_493);
and U930 (N_930,In_898,In_374);
nand U931 (N_931,In_213,In_650);
and U932 (N_932,In_980,In_228);
and U933 (N_933,In_975,In_852);
and U934 (N_934,In_817,In_951);
nand U935 (N_935,In_486,In_506);
nand U936 (N_936,In_965,In_350);
nand U937 (N_937,In_833,In_741);
nor U938 (N_938,In_47,In_589);
or U939 (N_939,In_662,In_199);
nor U940 (N_940,In_480,In_129);
nor U941 (N_941,In_719,In_656);
or U942 (N_942,In_497,In_801);
nand U943 (N_943,In_759,In_163);
nand U944 (N_944,In_751,In_598);
nand U945 (N_945,In_300,In_135);
or U946 (N_946,In_573,In_386);
and U947 (N_947,In_174,In_821);
or U948 (N_948,In_913,In_756);
and U949 (N_949,In_678,In_587);
nand U950 (N_950,In_509,In_520);
nand U951 (N_951,In_8,In_50);
xor U952 (N_952,In_627,In_282);
nand U953 (N_953,In_660,In_909);
nand U954 (N_954,In_884,In_55);
nor U955 (N_955,In_569,In_971);
nand U956 (N_956,In_786,In_257);
or U957 (N_957,In_98,In_764);
and U958 (N_958,In_801,In_909);
xor U959 (N_959,In_865,In_465);
nor U960 (N_960,In_164,In_199);
nor U961 (N_961,In_934,In_446);
and U962 (N_962,In_138,In_754);
nor U963 (N_963,In_102,In_958);
nand U964 (N_964,In_528,In_64);
nand U965 (N_965,In_81,In_414);
or U966 (N_966,In_355,In_261);
or U967 (N_967,In_138,In_151);
nor U968 (N_968,In_333,In_781);
or U969 (N_969,In_729,In_728);
nor U970 (N_970,In_781,In_366);
and U971 (N_971,In_240,In_839);
or U972 (N_972,In_556,In_370);
nand U973 (N_973,In_376,In_994);
nand U974 (N_974,In_769,In_390);
nor U975 (N_975,In_523,In_303);
nand U976 (N_976,In_973,In_476);
and U977 (N_977,In_978,In_351);
xor U978 (N_978,In_839,In_596);
nor U979 (N_979,In_897,In_500);
or U980 (N_980,In_267,In_53);
nor U981 (N_981,In_0,In_247);
nor U982 (N_982,In_780,In_146);
nand U983 (N_983,In_779,In_154);
nand U984 (N_984,In_865,In_558);
or U985 (N_985,In_503,In_653);
or U986 (N_986,In_357,In_255);
nor U987 (N_987,In_761,In_642);
nand U988 (N_988,In_456,In_970);
nor U989 (N_989,In_538,In_446);
or U990 (N_990,In_115,In_853);
and U991 (N_991,In_710,In_156);
xor U992 (N_992,In_923,In_971);
nor U993 (N_993,In_668,In_681);
nor U994 (N_994,In_538,In_628);
nand U995 (N_995,In_871,In_356);
nor U996 (N_996,In_243,In_907);
and U997 (N_997,In_68,In_375);
and U998 (N_998,In_961,In_898);
or U999 (N_999,In_252,In_615);
or U1000 (N_1000,In_282,In_780);
nor U1001 (N_1001,In_238,In_181);
or U1002 (N_1002,In_728,In_873);
nor U1003 (N_1003,In_489,In_69);
and U1004 (N_1004,In_387,In_631);
and U1005 (N_1005,In_487,In_878);
or U1006 (N_1006,In_353,In_34);
nor U1007 (N_1007,In_495,In_566);
or U1008 (N_1008,In_13,In_197);
nand U1009 (N_1009,In_520,In_801);
nor U1010 (N_1010,In_374,In_560);
and U1011 (N_1011,In_956,In_285);
nand U1012 (N_1012,In_444,In_969);
and U1013 (N_1013,In_581,In_160);
and U1014 (N_1014,In_972,In_879);
nor U1015 (N_1015,In_742,In_825);
xnor U1016 (N_1016,In_12,In_830);
and U1017 (N_1017,In_448,In_304);
nand U1018 (N_1018,In_476,In_125);
and U1019 (N_1019,In_704,In_560);
and U1020 (N_1020,In_115,In_901);
or U1021 (N_1021,In_703,In_469);
or U1022 (N_1022,In_595,In_147);
nor U1023 (N_1023,In_383,In_851);
and U1024 (N_1024,In_95,In_475);
nor U1025 (N_1025,In_416,In_515);
nand U1026 (N_1026,In_732,In_778);
or U1027 (N_1027,In_391,In_551);
xor U1028 (N_1028,In_679,In_2);
nand U1029 (N_1029,In_138,In_800);
or U1030 (N_1030,In_982,In_811);
nand U1031 (N_1031,In_116,In_212);
nand U1032 (N_1032,In_619,In_443);
nor U1033 (N_1033,In_453,In_915);
nand U1034 (N_1034,In_288,In_112);
nor U1035 (N_1035,In_951,In_527);
or U1036 (N_1036,In_333,In_959);
nand U1037 (N_1037,In_402,In_550);
or U1038 (N_1038,In_673,In_416);
nor U1039 (N_1039,In_61,In_293);
and U1040 (N_1040,In_558,In_318);
and U1041 (N_1041,In_173,In_200);
and U1042 (N_1042,In_896,In_161);
or U1043 (N_1043,In_427,In_607);
or U1044 (N_1044,In_338,In_876);
xor U1045 (N_1045,In_795,In_541);
and U1046 (N_1046,In_638,In_447);
nand U1047 (N_1047,In_466,In_965);
nor U1048 (N_1048,In_770,In_670);
nor U1049 (N_1049,In_249,In_297);
nor U1050 (N_1050,In_805,In_100);
and U1051 (N_1051,In_822,In_303);
nor U1052 (N_1052,In_42,In_434);
xor U1053 (N_1053,In_107,In_819);
nor U1054 (N_1054,In_767,In_137);
or U1055 (N_1055,In_580,In_306);
or U1056 (N_1056,In_262,In_465);
nand U1057 (N_1057,In_797,In_690);
nand U1058 (N_1058,In_638,In_45);
nor U1059 (N_1059,In_938,In_103);
or U1060 (N_1060,In_802,In_396);
xor U1061 (N_1061,In_248,In_344);
nor U1062 (N_1062,In_279,In_588);
nor U1063 (N_1063,In_351,In_993);
nor U1064 (N_1064,In_108,In_869);
nand U1065 (N_1065,In_863,In_802);
xor U1066 (N_1066,In_425,In_19);
nand U1067 (N_1067,In_983,In_135);
nand U1068 (N_1068,In_578,In_781);
and U1069 (N_1069,In_604,In_394);
nand U1070 (N_1070,In_479,In_319);
nor U1071 (N_1071,In_491,In_457);
and U1072 (N_1072,In_649,In_924);
or U1073 (N_1073,In_12,In_858);
and U1074 (N_1074,In_305,In_317);
and U1075 (N_1075,In_98,In_249);
or U1076 (N_1076,In_792,In_542);
nand U1077 (N_1077,In_478,In_184);
and U1078 (N_1078,In_390,In_9);
nand U1079 (N_1079,In_953,In_442);
and U1080 (N_1080,In_518,In_95);
and U1081 (N_1081,In_904,In_631);
nor U1082 (N_1082,In_917,In_420);
nor U1083 (N_1083,In_808,In_901);
or U1084 (N_1084,In_160,In_446);
nand U1085 (N_1085,In_555,In_534);
or U1086 (N_1086,In_348,In_720);
nand U1087 (N_1087,In_825,In_45);
xor U1088 (N_1088,In_662,In_587);
and U1089 (N_1089,In_760,In_339);
and U1090 (N_1090,In_108,In_494);
nand U1091 (N_1091,In_153,In_516);
or U1092 (N_1092,In_901,In_183);
nand U1093 (N_1093,In_358,In_513);
nand U1094 (N_1094,In_791,In_894);
or U1095 (N_1095,In_340,In_769);
nand U1096 (N_1096,In_104,In_627);
nor U1097 (N_1097,In_826,In_315);
nor U1098 (N_1098,In_864,In_518);
nor U1099 (N_1099,In_183,In_257);
nand U1100 (N_1100,In_462,In_975);
and U1101 (N_1101,In_285,In_853);
or U1102 (N_1102,In_694,In_567);
nand U1103 (N_1103,In_785,In_605);
nor U1104 (N_1104,In_643,In_695);
or U1105 (N_1105,In_869,In_600);
nor U1106 (N_1106,In_275,In_712);
or U1107 (N_1107,In_547,In_442);
nor U1108 (N_1108,In_773,In_979);
and U1109 (N_1109,In_285,In_913);
and U1110 (N_1110,In_180,In_609);
and U1111 (N_1111,In_976,In_776);
nand U1112 (N_1112,In_713,In_488);
and U1113 (N_1113,In_296,In_653);
or U1114 (N_1114,In_933,In_434);
nand U1115 (N_1115,In_904,In_646);
nor U1116 (N_1116,In_446,In_692);
and U1117 (N_1117,In_972,In_818);
nand U1118 (N_1118,In_455,In_619);
nor U1119 (N_1119,In_767,In_573);
nand U1120 (N_1120,In_824,In_876);
nor U1121 (N_1121,In_555,In_957);
nor U1122 (N_1122,In_44,In_306);
nor U1123 (N_1123,In_975,In_772);
nor U1124 (N_1124,In_193,In_493);
or U1125 (N_1125,In_442,In_12);
or U1126 (N_1126,In_248,In_129);
and U1127 (N_1127,In_670,In_965);
or U1128 (N_1128,In_470,In_718);
nor U1129 (N_1129,In_557,In_56);
and U1130 (N_1130,In_873,In_638);
or U1131 (N_1131,In_376,In_773);
nand U1132 (N_1132,In_962,In_668);
and U1133 (N_1133,In_597,In_145);
nor U1134 (N_1134,In_52,In_154);
or U1135 (N_1135,In_871,In_502);
nand U1136 (N_1136,In_0,In_563);
nand U1137 (N_1137,In_18,In_152);
nand U1138 (N_1138,In_743,In_92);
nor U1139 (N_1139,In_999,In_215);
and U1140 (N_1140,In_733,In_342);
and U1141 (N_1141,In_51,In_163);
or U1142 (N_1142,In_576,In_141);
and U1143 (N_1143,In_377,In_542);
nand U1144 (N_1144,In_73,In_382);
and U1145 (N_1145,In_838,In_614);
and U1146 (N_1146,In_342,In_517);
nor U1147 (N_1147,In_386,In_627);
nor U1148 (N_1148,In_416,In_756);
or U1149 (N_1149,In_774,In_264);
or U1150 (N_1150,In_336,In_454);
and U1151 (N_1151,In_40,In_423);
or U1152 (N_1152,In_377,In_687);
or U1153 (N_1153,In_818,In_980);
nand U1154 (N_1154,In_822,In_411);
or U1155 (N_1155,In_847,In_800);
nand U1156 (N_1156,In_682,In_605);
or U1157 (N_1157,In_289,In_81);
nor U1158 (N_1158,In_356,In_464);
or U1159 (N_1159,In_920,In_692);
and U1160 (N_1160,In_232,In_559);
or U1161 (N_1161,In_883,In_336);
nand U1162 (N_1162,In_973,In_948);
or U1163 (N_1163,In_748,In_565);
nor U1164 (N_1164,In_585,In_654);
nand U1165 (N_1165,In_257,In_239);
or U1166 (N_1166,In_376,In_234);
nor U1167 (N_1167,In_499,In_807);
or U1168 (N_1168,In_365,In_899);
nor U1169 (N_1169,In_227,In_98);
and U1170 (N_1170,In_956,In_463);
nor U1171 (N_1171,In_223,In_682);
nand U1172 (N_1172,In_487,In_738);
or U1173 (N_1173,In_48,In_477);
nand U1174 (N_1174,In_649,In_113);
xnor U1175 (N_1175,In_421,In_809);
and U1176 (N_1176,In_752,In_144);
and U1177 (N_1177,In_64,In_376);
and U1178 (N_1178,In_623,In_512);
nor U1179 (N_1179,In_452,In_603);
or U1180 (N_1180,In_490,In_551);
or U1181 (N_1181,In_179,In_815);
and U1182 (N_1182,In_69,In_563);
nand U1183 (N_1183,In_258,In_83);
nand U1184 (N_1184,In_325,In_142);
nand U1185 (N_1185,In_573,In_588);
and U1186 (N_1186,In_484,In_135);
or U1187 (N_1187,In_393,In_647);
and U1188 (N_1188,In_91,In_863);
and U1189 (N_1189,In_756,In_71);
nand U1190 (N_1190,In_988,In_906);
or U1191 (N_1191,In_322,In_231);
and U1192 (N_1192,In_715,In_25);
nor U1193 (N_1193,In_538,In_440);
nor U1194 (N_1194,In_502,In_591);
nor U1195 (N_1195,In_117,In_500);
nor U1196 (N_1196,In_881,In_892);
nor U1197 (N_1197,In_375,In_505);
xor U1198 (N_1198,In_572,In_58);
nand U1199 (N_1199,In_376,In_119);
and U1200 (N_1200,In_806,In_934);
nand U1201 (N_1201,In_829,In_383);
or U1202 (N_1202,In_995,In_354);
nand U1203 (N_1203,In_567,In_368);
nor U1204 (N_1204,In_494,In_55);
or U1205 (N_1205,In_485,In_294);
xor U1206 (N_1206,In_765,In_100);
or U1207 (N_1207,In_736,In_909);
and U1208 (N_1208,In_618,In_264);
nor U1209 (N_1209,In_563,In_190);
or U1210 (N_1210,In_910,In_976);
or U1211 (N_1211,In_102,In_155);
or U1212 (N_1212,In_214,In_644);
and U1213 (N_1213,In_440,In_844);
and U1214 (N_1214,In_794,In_940);
nand U1215 (N_1215,In_530,In_255);
and U1216 (N_1216,In_910,In_14);
or U1217 (N_1217,In_180,In_822);
and U1218 (N_1218,In_125,In_33);
or U1219 (N_1219,In_429,In_176);
nor U1220 (N_1220,In_20,In_146);
or U1221 (N_1221,In_997,In_128);
nand U1222 (N_1222,In_262,In_905);
or U1223 (N_1223,In_562,In_522);
nand U1224 (N_1224,In_349,In_831);
nor U1225 (N_1225,In_787,In_794);
nor U1226 (N_1226,In_593,In_688);
nor U1227 (N_1227,In_19,In_6);
nor U1228 (N_1228,In_841,In_830);
nor U1229 (N_1229,In_221,In_824);
or U1230 (N_1230,In_908,In_214);
nand U1231 (N_1231,In_796,In_771);
and U1232 (N_1232,In_734,In_244);
and U1233 (N_1233,In_578,In_178);
and U1234 (N_1234,In_655,In_302);
nor U1235 (N_1235,In_585,In_665);
or U1236 (N_1236,In_105,In_617);
and U1237 (N_1237,In_78,In_217);
and U1238 (N_1238,In_148,In_327);
or U1239 (N_1239,In_750,In_20);
or U1240 (N_1240,In_832,In_779);
or U1241 (N_1241,In_199,In_628);
nand U1242 (N_1242,In_648,In_515);
xnor U1243 (N_1243,In_437,In_293);
and U1244 (N_1244,In_687,In_850);
nor U1245 (N_1245,In_221,In_962);
and U1246 (N_1246,In_110,In_723);
nand U1247 (N_1247,In_866,In_984);
nor U1248 (N_1248,In_873,In_942);
nor U1249 (N_1249,In_66,In_417);
and U1250 (N_1250,In_343,In_776);
or U1251 (N_1251,In_53,In_699);
nand U1252 (N_1252,In_646,In_536);
or U1253 (N_1253,In_982,In_973);
nor U1254 (N_1254,In_447,In_13);
nand U1255 (N_1255,In_232,In_62);
and U1256 (N_1256,In_932,In_924);
nand U1257 (N_1257,In_506,In_992);
and U1258 (N_1258,In_526,In_978);
nor U1259 (N_1259,In_978,In_878);
xor U1260 (N_1260,In_898,In_376);
or U1261 (N_1261,In_460,In_110);
nor U1262 (N_1262,In_543,In_84);
nand U1263 (N_1263,In_403,In_480);
or U1264 (N_1264,In_82,In_752);
xor U1265 (N_1265,In_267,In_967);
nand U1266 (N_1266,In_707,In_102);
or U1267 (N_1267,In_729,In_374);
nand U1268 (N_1268,In_403,In_679);
or U1269 (N_1269,In_723,In_805);
nand U1270 (N_1270,In_443,In_631);
and U1271 (N_1271,In_625,In_239);
or U1272 (N_1272,In_148,In_41);
or U1273 (N_1273,In_642,In_840);
or U1274 (N_1274,In_403,In_761);
nor U1275 (N_1275,In_84,In_3);
nand U1276 (N_1276,In_854,In_538);
nand U1277 (N_1277,In_758,In_71);
nand U1278 (N_1278,In_605,In_554);
nand U1279 (N_1279,In_774,In_806);
nor U1280 (N_1280,In_430,In_722);
nand U1281 (N_1281,In_735,In_664);
and U1282 (N_1282,In_579,In_67);
nor U1283 (N_1283,In_743,In_705);
or U1284 (N_1284,In_495,In_45);
nand U1285 (N_1285,In_658,In_450);
nand U1286 (N_1286,In_686,In_790);
nand U1287 (N_1287,In_889,In_623);
or U1288 (N_1288,In_218,In_481);
nand U1289 (N_1289,In_408,In_651);
and U1290 (N_1290,In_499,In_297);
and U1291 (N_1291,In_790,In_722);
nand U1292 (N_1292,In_860,In_355);
and U1293 (N_1293,In_595,In_644);
and U1294 (N_1294,In_555,In_436);
nor U1295 (N_1295,In_990,In_152);
nand U1296 (N_1296,In_333,In_133);
nand U1297 (N_1297,In_153,In_442);
or U1298 (N_1298,In_672,In_519);
nand U1299 (N_1299,In_71,In_985);
nand U1300 (N_1300,In_627,In_338);
nand U1301 (N_1301,In_703,In_669);
and U1302 (N_1302,In_982,In_295);
nor U1303 (N_1303,In_647,In_695);
nand U1304 (N_1304,In_834,In_617);
and U1305 (N_1305,In_789,In_715);
or U1306 (N_1306,In_174,In_896);
nor U1307 (N_1307,In_537,In_519);
nor U1308 (N_1308,In_507,In_813);
nand U1309 (N_1309,In_424,In_600);
nor U1310 (N_1310,In_681,In_133);
nand U1311 (N_1311,In_49,In_813);
nor U1312 (N_1312,In_662,In_79);
nor U1313 (N_1313,In_985,In_750);
nand U1314 (N_1314,In_417,In_576);
nor U1315 (N_1315,In_319,In_150);
and U1316 (N_1316,In_293,In_719);
nor U1317 (N_1317,In_371,In_722);
and U1318 (N_1318,In_630,In_339);
nand U1319 (N_1319,In_259,In_236);
nor U1320 (N_1320,In_419,In_296);
or U1321 (N_1321,In_845,In_204);
and U1322 (N_1322,In_220,In_713);
nor U1323 (N_1323,In_161,In_54);
nand U1324 (N_1324,In_604,In_3);
nor U1325 (N_1325,In_482,In_152);
nor U1326 (N_1326,In_210,In_463);
nand U1327 (N_1327,In_35,In_282);
or U1328 (N_1328,In_925,In_116);
nor U1329 (N_1329,In_398,In_992);
and U1330 (N_1330,In_482,In_475);
nor U1331 (N_1331,In_589,In_358);
nor U1332 (N_1332,In_135,In_720);
nand U1333 (N_1333,In_536,In_307);
nand U1334 (N_1334,In_811,In_390);
nor U1335 (N_1335,In_433,In_343);
and U1336 (N_1336,In_395,In_427);
or U1337 (N_1337,In_775,In_198);
and U1338 (N_1338,In_76,In_838);
and U1339 (N_1339,In_807,In_124);
nor U1340 (N_1340,In_387,In_130);
nand U1341 (N_1341,In_597,In_616);
nor U1342 (N_1342,In_968,In_384);
nand U1343 (N_1343,In_709,In_374);
or U1344 (N_1344,In_462,In_981);
and U1345 (N_1345,In_394,In_954);
and U1346 (N_1346,In_261,In_590);
or U1347 (N_1347,In_560,In_861);
nor U1348 (N_1348,In_97,In_147);
nor U1349 (N_1349,In_519,In_456);
nor U1350 (N_1350,In_703,In_301);
nand U1351 (N_1351,In_322,In_602);
nand U1352 (N_1352,In_505,In_979);
or U1353 (N_1353,In_101,In_969);
and U1354 (N_1354,In_308,In_630);
nand U1355 (N_1355,In_670,In_874);
and U1356 (N_1356,In_293,In_375);
nand U1357 (N_1357,In_738,In_953);
nor U1358 (N_1358,In_955,In_548);
nand U1359 (N_1359,In_651,In_902);
nor U1360 (N_1360,In_367,In_603);
nand U1361 (N_1361,In_628,In_247);
or U1362 (N_1362,In_477,In_886);
or U1363 (N_1363,In_234,In_39);
nor U1364 (N_1364,In_439,In_61);
or U1365 (N_1365,In_678,In_632);
and U1366 (N_1366,In_858,In_51);
nand U1367 (N_1367,In_140,In_943);
nor U1368 (N_1368,In_454,In_362);
nand U1369 (N_1369,In_460,In_806);
nor U1370 (N_1370,In_395,In_615);
or U1371 (N_1371,In_697,In_7);
nor U1372 (N_1372,In_131,In_981);
nand U1373 (N_1373,In_112,In_610);
nor U1374 (N_1374,In_226,In_312);
or U1375 (N_1375,In_273,In_349);
nand U1376 (N_1376,In_551,In_847);
or U1377 (N_1377,In_896,In_442);
nand U1378 (N_1378,In_287,In_396);
or U1379 (N_1379,In_927,In_467);
nor U1380 (N_1380,In_110,In_366);
or U1381 (N_1381,In_180,In_475);
and U1382 (N_1382,In_570,In_388);
nor U1383 (N_1383,In_101,In_378);
xor U1384 (N_1384,In_768,In_843);
and U1385 (N_1385,In_698,In_363);
nor U1386 (N_1386,In_49,In_781);
nand U1387 (N_1387,In_228,In_55);
or U1388 (N_1388,In_8,In_932);
nand U1389 (N_1389,In_639,In_740);
nand U1390 (N_1390,In_520,In_979);
and U1391 (N_1391,In_752,In_521);
nand U1392 (N_1392,In_542,In_12);
or U1393 (N_1393,In_995,In_53);
nand U1394 (N_1394,In_4,In_571);
nand U1395 (N_1395,In_789,In_921);
nand U1396 (N_1396,In_599,In_246);
or U1397 (N_1397,In_672,In_357);
nand U1398 (N_1398,In_160,In_575);
and U1399 (N_1399,In_329,In_521);
and U1400 (N_1400,In_684,In_356);
or U1401 (N_1401,In_483,In_67);
and U1402 (N_1402,In_454,In_684);
nor U1403 (N_1403,In_361,In_794);
or U1404 (N_1404,In_750,In_856);
or U1405 (N_1405,In_362,In_690);
or U1406 (N_1406,In_11,In_217);
nor U1407 (N_1407,In_840,In_232);
nor U1408 (N_1408,In_500,In_471);
nor U1409 (N_1409,In_231,In_93);
nand U1410 (N_1410,In_357,In_944);
nand U1411 (N_1411,In_741,In_397);
nor U1412 (N_1412,In_377,In_201);
nand U1413 (N_1413,In_97,In_540);
nor U1414 (N_1414,In_280,In_638);
or U1415 (N_1415,In_649,In_7);
xnor U1416 (N_1416,In_59,In_983);
nand U1417 (N_1417,In_309,In_423);
nor U1418 (N_1418,In_461,In_703);
xor U1419 (N_1419,In_810,In_436);
nand U1420 (N_1420,In_816,In_651);
nor U1421 (N_1421,In_985,In_371);
nor U1422 (N_1422,In_0,In_886);
or U1423 (N_1423,In_876,In_433);
xor U1424 (N_1424,In_374,In_866);
nand U1425 (N_1425,In_80,In_128);
and U1426 (N_1426,In_117,In_434);
and U1427 (N_1427,In_743,In_486);
nand U1428 (N_1428,In_969,In_480);
and U1429 (N_1429,In_87,In_566);
and U1430 (N_1430,In_803,In_200);
nand U1431 (N_1431,In_364,In_73);
and U1432 (N_1432,In_35,In_140);
or U1433 (N_1433,In_713,In_634);
nor U1434 (N_1434,In_497,In_572);
nor U1435 (N_1435,In_118,In_915);
or U1436 (N_1436,In_105,In_739);
and U1437 (N_1437,In_939,In_560);
or U1438 (N_1438,In_133,In_696);
nor U1439 (N_1439,In_829,In_152);
or U1440 (N_1440,In_730,In_181);
nor U1441 (N_1441,In_339,In_625);
or U1442 (N_1442,In_404,In_406);
and U1443 (N_1443,In_880,In_204);
or U1444 (N_1444,In_830,In_541);
nor U1445 (N_1445,In_487,In_112);
or U1446 (N_1446,In_226,In_492);
nand U1447 (N_1447,In_694,In_266);
and U1448 (N_1448,In_63,In_765);
or U1449 (N_1449,In_31,In_964);
and U1450 (N_1450,In_646,In_237);
or U1451 (N_1451,In_436,In_853);
xor U1452 (N_1452,In_166,In_51);
xor U1453 (N_1453,In_832,In_490);
and U1454 (N_1454,In_510,In_76);
or U1455 (N_1455,In_491,In_581);
and U1456 (N_1456,In_709,In_71);
nor U1457 (N_1457,In_890,In_624);
nand U1458 (N_1458,In_444,In_948);
nand U1459 (N_1459,In_40,In_5);
or U1460 (N_1460,In_655,In_662);
and U1461 (N_1461,In_321,In_633);
nand U1462 (N_1462,In_41,In_543);
nand U1463 (N_1463,In_181,In_613);
nor U1464 (N_1464,In_169,In_115);
nor U1465 (N_1465,In_763,In_385);
nor U1466 (N_1466,In_605,In_862);
nor U1467 (N_1467,In_249,In_811);
nand U1468 (N_1468,In_534,In_160);
or U1469 (N_1469,In_487,In_745);
nand U1470 (N_1470,In_97,In_850);
nand U1471 (N_1471,In_460,In_474);
and U1472 (N_1472,In_41,In_633);
nand U1473 (N_1473,In_932,In_176);
and U1474 (N_1474,In_250,In_168);
nor U1475 (N_1475,In_366,In_104);
or U1476 (N_1476,In_840,In_821);
nor U1477 (N_1477,In_379,In_827);
nor U1478 (N_1478,In_668,In_557);
or U1479 (N_1479,In_988,In_72);
and U1480 (N_1480,In_509,In_427);
or U1481 (N_1481,In_65,In_588);
nor U1482 (N_1482,In_796,In_187);
or U1483 (N_1483,In_823,In_310);
nand U1484 (N_1484,In_278,In_680);
and U1485 (N_1485,In_112,In_930);
nand U1486 (N_1486,In_461,In_963);
nand U1487 (N_1487,In_535,In_30);
nand U1488 (N_1488,In_145,In_791);
nand U1489 (N_1489,In_719,In_613);
nor U1490 (N_1490,In_524,In_477);
or U1491 (N_1491,In_733,In_365);
nor U1492 (N_1492,In_751,In_932);
and U1493 (N_1493,In_699,In_992);
nor U1494 (N_1494,In_364,In_878);
or U1495 (N_1495,In_390,In_343);
or U1496 (N_1496,In_60,In_675);
nand U1497 (N_1497,In_755,In_825);
xnor U1498 (N_1498,In_587,In_85);
nor U1499 (N_1499,In_570,In_338);
xor U1500 (N_1500,In_744,In_520);
nand U1501 (N_1501,In_604,In_352);
nor U1502 (N_1502,In_11,In_474);
nand U1503 (N_1503,In_996,In_372);
or U1504 (N_1504,In_28,In_965);
and U1505 (N_1505,In_52,In_194);
nand U1506 (N_1506,In_143,In_19);
or U1507 (N_1507,In_459,In_166);
nor U1508 (N_1508,In_243,In_163);
nor U1509 (N_1509,In_784,In_676);
and U1510 (N_1510,In_832,In_344);
and U1511 (N_1511,In_569,In_287);
or U1512 (N_1512,In_54,In_879);
nor U1513 (N_1513,In_710,In_592);
nand U1514 (N_1514,In_800,In_85);
or U1515 (N_1515,In_535,In_62);
or U1516 (N_1516,In_747,In_927);
or U1517 (N_1517,In_540,In_111);
nand U1518 (N_1518,In_706,In_669);
and U1519 (N_1519,In_902,In_184);
nand U1520 (N_1520,In_270,In_90);
nor U1521 (N_1521,In_628,In_358);
nand U1522 (N_1522,In_804,In_651);
xor U1523 (N_1523,In_91,In_513);
nand U1524 (N_1524,In_127,In_511);
nand U1525 (N_1525,In_189,In_667);
and U1526 (N_1526,In_480,In_610);
or U1527 (N_1527,In_607,In_249);
or U1528 (N_1528,In_815,In_571);
nor U1529 (N_1529,In_437,In_3);
xnor U1530 (N_1530,In_616,In_524);
and U1531 (N_1531,In_379,In_947);
nand U1532 (N_1532,In_125,In_547);
or U1533 (N_1533,In_123,In_771);
nand U1534 (N_1534,In_302,In_44);
nand U1535 (N_1535,In_210,In_145);
nand U1536 (N_1536,In_573,In_154);
or U1537 (N_1537,In_354,In_180);
and U1538 (N_1538,In_739,In_769);
and U1539 (N_1539,In_619,In_685);
and U1540 (N_1540,In_475,In_957);
or U1541 (N_1541,In_439,In_282);
or U1542 (N_1542,In_365,In_77);
nand U1543 (N_1543,In_306,In_480);
and U1544 (N_1544,In_664,In_964);
nand U1545 (N_1545,In_965,In_123);
nor U1546 (N_1546,In_251,In_642);
and U1547 (N_1547,In_362,In_577);
and U1548 (N_1548,In_889,In_132);
nand U1549 (N_1549,In_910,In_570);
nor U1550 (N_1550,In_816,In_17);
and U1551 (N_1551,In_359,In_949);
nor U1552 (N_1552,In_68,In_970);
and U1553 (N_1553,In_210,In_148);
xor U1554 (N_1554,In_78,In_736);
nor U1555 (N_1555,In_298,In_585);
nand U1556 (N_1556,In_405,In_310);
nand U1557 (N_1557,In_924,In_144);
xor U1558 (N_1558,In_962,In_304);
nor U1559 (N_1559,In_87,In_701);
and U1560 (N_1560,In_912,In_887);
or U1561 (N_1561,In_24,In_665);
nor U1562 (N_1562,In_245,In_181);
nand U1563 (N_1563,In_579,In_685);
and U1564 (N_1564,In_937,In_95);
nand U1565 (N_1565,In_91,In_275);
nand U1566 (N_1566,In_89,In_622);
or U1567 (N_1567,In_544,In_866);
and U1568 (N_1568,In_19,In_703);
nand U1569 (N_1569,In_307,In_15);
nand U1570 (N_1570,In_971,In_694);
nor U1571 (N_1571,In_924,In_104);
or U1572 (N_1572,In_739,In_116);
nor U1573 (N_1573,In_430,In_288);
and U1574 (N_1574,In_634,In_781);
nor U1575 (N_1575,In_521,In_598);
or U1576 (N_1576,In_88,In_593);
or U1577 (N_1577,In_393,In_655);
and U1578 (N_1578,In_592,In_129);
nand U1579 (N_1579,In_694,In_873);
or U1580 (N_1580,In_781,In_253);
nor U1581 (N_1581,In_468,In_213);
nand U1582 (N_1582,In_769,In_622);
or U1583 (N_1583,In_697,In_250);
nand U1584 (N_1584,In_94,In_15);
nand U1585 (N_1585,In_517,In_2);
nor U1586 (N_1586,In_351,In_862);
or U1587 (N_1587,In_975,In_756);
nand U1588 (N_1588,In_178,In_414);
nand U1589 (N_1589,In_924,In_325);
and U1590 (N_1590,In_584,In_463);
nor U1591 (N_1591,In_591,In_994);
nand U1592 (N_1592,In_914,In_523);
nor U1593 (N_1593,In_684,In_767);
nand U1594 (N_1594,In_965,In_467);
nand U1595 (N_1595,In_172,In_936);
and U1596 (N_1596,In_162,In_338);
or U1597 (N_1597,In_841,In_291);
or U1598 (N_1598,In_699,In_479);
and U1599 (N_1599,In_720,In_876);
nand U1600 (N_1600,In_361,In_439);
nand U1601 (N_1601,In_666,In_215);
or U1602 (N_1602,In_458,In_471);
or U1603 (N_1603,In_311,In_22);
and U1604 (N_1604,In_684,In_307);
and U1605 (N_1605,In_973,In_442);
or U1606 (N_1606,In_480,In_472);
nand U1607 (N_1607,In_98,In_700);
nand U1608 (N_1608,In_714,In_895);
nand U1609 (N_1609,In_726,In_425);
or U1610 (N_1610,In_307,In_772);
nor U1611 (N_1611,In_131,In_588);
or U1612 (N_1612,In_258,In_478);
nand U1613 (N_1613,In_289,In_408);
nor U1614 (N_1614,In_280,In_543);
and U1615 (N_1615,In_903,In_867);
nand U1616 (N_1616,In_742,In_177);
nand U1617 (N_1617,In_372,In_412);
or U1618 (N_1618,In_736,In_866);
xnor U1619 (N_1619,In_833,In_848);
nand U1620 (N_1620,In_351,In_242);
and U1621 (N_1621,In_112,In_251);
and U1622 (N_1622,In_222,In_870);
or U1623 (N_1623,In_185,In_716);
and U1624 (N_1624,In_590,In_776);
nor U1625 (N_1625,In_57,In_242);
and U1626 (N_1626,In_833,In_951);
nor U1627 (N_1627,In_518,In_833);
xor U1628 (N_1628,In_619,In_859);
and U1629 (N_1629,In_156,In_795);
nand U1630 (N_1630,In_200,In_30);
nand U1631 (N_1631,In_270,In_925);
or U1632 (N_1632,In_857,In_533);
and U1633 (N_1633,In_273,In_632);
xor U1634 (N_1634,In_370,In_466);
nor U1635 (N_1635,In_571,In_791);
and U1636 (N_1636,In_315,In_346);
nor U1637 (N_1637,In_72,In_553);
nor U1638 (N_1638,In_545,In_432);
nor U1639 (N_1639,In_183,In_858);
nand U1640 (N_1640,In_421,In_531);
and U1641 (N_1641,In_172,In_900);
nand U1642 (N_1642,In_746,In_552);
or U1643 (N_1643,In_955,In_830);
nor U1644 (N_1644,In_441,In_943);
or U1645 (N_1645,In_503,In_145);
nand U1646 (N_1646,In_334,In_946);
nand U1647 (N_1647,In_262,In_353);
and U1648 (N_1648,In_651,In_688);
nor U1649 (N_1649,In_200,In_324);
xor U1650 (N_1650,In_236,In_213);
nor U1651 (N_1651,In_574,In_162);
and U1652 (N_1652,In_301,In_604);
nor U1653 (N_1653,In_324,In_527);
nor U1654 (N_1654,In_126,In_151);
and U1655 (N_1655,In_131,In_0);
nand U1656 (N_1656,In_543,In_193);
or U1657 (N_1657,In_923,In_888);
nand U1658 (N_1658,In_979,In_771);
nor U1659 (N_1659,In_701,In_691);
and U1660 (N_1660,In_859,In_3);
and U1661 (N_1661,In_477,In_353);
nor U1662 (N_1662,In_390,In_698);
or U1663 (N_1663,In_357,In_288);
nand U1664 (N_1664,In_882,In_475);
and U1665 (N_1665,In_820,In_887);
nand U1666 (N_1666,In_829,In_419);
or U1667 (N_1667,In_401,In_610);
nor U1668 (N_1668,In_590,In_964);
nor U1669 (N_1669,In_420,In_144);
nor U1670 (N_1670,In_652,In_798);
nand U1671 (N_1671,In_115,In_217);
nand U1672 (N_1672,In_705,In_439);
or U1673 (N_1673,In_894,In_187);
and U1674 (N_1674,In_576,In_138);
and U1675 (N_1675,In_58,In_689);
nor U1676 (N_1676,In_443,In_415);
xnor U1677 (N_1677,In_761,In_461);
xor U1678 (N_1678,In_266,In_749);
nand U1679 (N_1679,In_129,In_167);
nor U1680 (N_1680,In_538,In_595);
nand U1681 (N_1681,In_156,In_296);
or U1682 (N_1682,In_904,In_455);
nor U1683 (N_1683,In_806,In_661);
and U1684 (N_1684,In_450,In_550);
or U1685 (N_1685,In_708,In_353);
nand U1686 (N_1686,In_447,In_251);
and U1687 (N_1687,In_714,In_949);
nor U1688 (N_1688,In_271,In_102);
and U1689 (N_1689,In_983,In_684);
nand U1690 (N_1690,In_579,In_881);
or U1691 (N_1691,In_491,In_966);
nand U1692 (N_1692,In_132,In_661);
or U1693 (N_1693,In_243,In_433);
and U1694 (N_1694,In_978,In_407);
or U1695 (N_1695,In_565,In_501);
or U1696 (N_1696,In_626,In_700);
or U1697 (N_1697,In_633,In_482);
nor U1698 (N_1698,In_787,In_343);
nor U1699 (N_1699,In_139,In_146);
nand U1700 (N_1700,In_298,In_548);
nor U1701 (N_1701,In_0,In_522);
and U1702 (N_1702,In_418,In_285);
and U1703 (N_1703,In_68,In_891);
nor U1704 (N_1704,In_591,In_227);
and U1705 (N_1705,In_776,In_674);
nor U1706 (N_1706,In_174,In_13);
nor U1707 (N_1707,In_532,In_675);
or U1708 (N_1708,In_757,In_162);
and U1709 (N_1709,In_944,In_998);
nor U1710 (N_1710,In_38,In_968);
nor U1711 (N_1711,In_672,In_805);
and U1712 (N_1712,In_71,In_653);
nor U1713 (N_1713,In_546,In_901);
and U1714 (N_1714,In_175,In_804);
nand U1715 (N_1715,In_784,In_561);
or U1716 (N_1716,In_824,In_373);
xor U1717 (N_1717,In_748,In_727);
or U1718 (N_1718,In_65,In_426);
nand U1719 (N_1719,In_419,In_976);
and U1720 (N_1720,In_23,In_124);
nor U1721 (N_1721,In_231,In_327);
or U1722 (N_1722,In_948,In_5);
nor U1723 (N_1723,In_737,In_767);
nand U1724 (N_1724,In_43,In_791);
and U1725 (N_1725,In_169,In_325);
and U1726 (N_1726,In_193,In_253);
and U1727 (N_1727,In_348,In_687);
and U1728 (N_1728,In_564,In_88);
nand U1729 (N_1729,In_682,In_18);
nor U1730 (N_1730,In_20,In_745);
or U1731 (N_1731,In_484,In_944);
and U1732 (N_1732,In_839,In_426);
nor U1733 (N_1733,In_442,In_923);
and U1734 (N_1734,In_968,In_388);
or U1735 (N_1735,In_490,In_777);
or U1736 (N_1736,In_779,In_953);
nand U1737 (N_1737,In_388,In_471);
or U1738 (N_1738,In_623,In_598);
nand U1739 (N_1739,In_974,In_632);
and U1740 (N_1740,In_636,In_739);
nor U1741 (N_1741,In_319,In_381);
and U1742 (N_1742,In_835,In_981);
and U1743 (N_1743,In_530,In_375);
or U1744 (N_1744,In_257,In_422);
or U1745 (N_1745,In_242,In_94);
or U1746 (N_1746,In_448,In_586);
nor U1747 (N_1747,In_925,In_528);
or U1748 (N_1748,In_347,In_961);
nand U1749 (N_1749,In_81,In_374);
or U1750 (N_1750,In_87,In_992);
nor U1751 (N_1751,In_891,In_142);
and U1752 (N_1752,In_774,In_245);
or U1753 (N_1753,In_674,In_313);
or U1754 (N_1754,In_434,In_173);
nand U1755 (N_1755,In_329,In_913);
or U1756 (N_1756,In_537,In_624);
and U1757 (N_1757,In_101,In_613);
nand U1758 (N_1758,In_706,In_58);
nand U1759 (N_1759,In_325,In_105);
and U1760 (N_1760,In_258,In_483);
and U1761 (N_1761,In_239,In_786);
and U1762 (N_1762,In_186,In_520);
nor U1763 (N_1763,In_67,In_988);
or U1764 (N_1764,In_334,In_93);
and U1765 (N_1765,In_692,In_464);
nand U1766 (N_1766,In_95,In_339);
and U1767 (N_1767,In_516,In_254);
and U1768 (N_1768,In_615,In_488);
xor U1769 (N_1769,In_325,In_451);
nor U1770 (N_1770,In_108,In_63);
or U1771 (N_1771,In_346,In_71);
or U1772 (N_1772,In_144,In_227);
nor U1773 (N_1773,In_317,In_309);
nand U1774 (N_1774,In_932,In_623);
nor U1775 (N_1775,In_670,In_946);
or U1776 (N_1776,In_420,In_306);
or U1777 (N_1777,In_272,In_885);
nor U1778 (N_1778,In_104,In_718);
nand U1779 (N_1779,In_558,In_727);
or U1780 (N_1780,In_646,In_253);
nand U1781 (N_1781,In_141,In_815);
nor U1782 (N_1782,In_549,In_829);
nand U1783 (N_1783,In_192,In_187);
nor U1784 (N_1784,In_642,In_630);
nor U1785 (N_1785,In_213,In_231);
nand U1786 (N_1786,In_632,In_279);
nor U1787 (N_1787,In_352,In_462);
or U1788 (N_1788,In_348,In_307);
nor U1789 (N_1789,In_191,In_797);
and U1790 (N_1790,In_282,In_985);
nor U1791 (N_1791,In_756,In_58);
nor U1792 (N_1792,In_422,In_604);
nand U1793 (N_1793,In_593,In_216);
or U1794 (N_1794,In_33,In_344);
nor U1795 (N_1795,In_83,In_27);
nor U1796 (N_1796,In_204,In_153);
nor U1797 (N_1797,In_197,In_47);
nand U1798 (N_1798,In_195,In_842);
or U1799 (N_1799,In_4,In_632);
nand U1800 (N_1800,In_983,In_926);
nand U1801 (N_1801,In_923,In_652);
nor U1802 (N_1802,In_7,In_951);
or U1803 (N_1803,In_183,In_895);
nor U1804 (N_1804,In_133,In_610);
and U1805 (N_1805,In_35,In_451);
nor U1806 (N_1806,In_313,In_676);
or U1807 (N_1807,In_0,In_449);
and U1808 (N_1808,In_540,In_259);
nand U1809 (N_1809,In_400,In_227);
nand U1810 (N_1810,In_694,In_520);
nand U1811 (N_1811,In_907,In_52);
nand U1812 (N_1812,In_907,In_428);
and U1813 (N_1813,In_176,In_700);
nand U1814 (N_1814,In_986,In_827);
nor U1815 (N_1815,In_577,In_300);
or U1816 (N_1816,In_409,In_885);
or U1817 (N_1817,In_139,In_14);
nand U1818 (N_1818,In_578,In_98);
or U1819 (N_1819,In_705,In_827);
nand U1820 (N_1820,In_238,In_188);
or U1821 (N_1821,In_723,In_890);
or U1822 (N_1822,In_680,In_83);
and U1823 (N_1823,In_271,In_255);
and U1824 (N_1824,In_370,In_746);
and U1825 (N_1825,In_700,In_704);
and U1826 (N_1826,In_432,In_178);
nand U1827 (N_1827,In_411,In_911);
and U1828 (N_1828,In_909,In_647);
nor U1829 (N_1829,In_380,In_35);
or U1830 (N_1830,In_741,In_394);
and U1831 (N_1831,In_946,In_44);
nand U1832 (N_1832,In_196,In_723);
or U1833 (N_1833,In_177,In_710);
or U1834 (N_1834,In_822,In_176);
or U1835 (N_1835,In_330,In_679);
nand U1836 (N_1836,In_800,In_311);
and U1837 (N_1837,In_788,In_760);
nor U1838 (N_1838,In_988,In_929);
nand U1839 (N_1839,In_324,In_958);
or U1840 (N_1840,In_625,In_774);
nor U1841 (N_1841,In_64,In_958);
nand U1842 (N_1842,In_575,In_421);
nor U1843 (N_1843,In_527,In_619);
nor U1844 (N_1844,In_760,In_775);
nand U1845 (N_1845,In_687,In_61);
and U1846 (N_1846,In_495,In_232);
or U1847 (N_1847,In_592,In_345);
nand U1848 (N_1848,In_169,In_98);
or U1849 (N_1849,In_184,In_189);
nand U1850 (N_1850,In_339,In_198);
nand U1851 (N_1851,In_650,In_680);
or U1852 (N_1852,In_653,In_925);
or U1853 (N_1853,In_591,In_720);
or U1854 (N_1854,In_983,In_859);
and U1855 (N_1855,In_694,In_684);
and U1856 (N_1856,In_968,In_139);
nand U1857 (N_1857,In_597,In_338);
nor U1858 (N_1858,In_929,In_164);
or U1859 (N_1859,In_118,In_168);
nand U1860 (N_1860,In_416,In_312);
or U1861 (N_1861,In_835,In_327);
or U1862 (N_1862,In_616,In_864);
xor U1863 (N_1863,In_482,In_700);
or U1864 (N_1864,In_89,In_251);
and U1865 (N_1865,In_955,In_925);
and U1866 (N_1866,In_994,In_567);
and U1867 (N_1867,In_91,In_191);
nor U1868 (N_1868,In_358,In_938);
and U1869 (N_1869,In_423,In_65);
and U1870 (N_1870,In_755,In_104);
nor U1871 (N_1871,In_952,In_773);
and U1872 (N_1872,In_801,In_741);
xnor U1873 (N_1873,In_317,In_329);
nand U1874 (N_1874,In_949,In_224);
and U1875 (N_1875,In_432,In_45);
nand U1876 (N_1876,In_678,In_28);
or U1877 (N_1877,In_516,In_624);
nor U1878 (N_1878,In_916,In_951);
nand U1879 (N_1879,In_469,In_101);
nand U1880 (N_1880,In_927,In_126);
nor U1881 (N_1881,In_963,In_21);
nor U1882 (N_1882,In_542,In_345);
xnor U1883 (N_1883,In_835,In_918);
nor U1884 (N_1884,In_234,In_19);
or U1885 (N_1885,In_734,In_494);
or U1886 (N_1886,In_442,In_287);
nor U1887 (N_1887,In_449,In_440);
nand U1888 (N_1888,In_87,In_372);
nor U1889 (N_1889,In_739,In_856);
nor U1890 (N_1890,In_711,In_200);
nor U1891 (N_1891,In_570,In_225);
nor U1892 (N_1892,In_625,In_439);
nand U1893 (N_1893,In_734,In_574);
and U1894 (N_1894,In_468,In_325);
and U1895 (N_1895,In_399,In_13);
nor U1896 (N_1896,In_352,In_802);
nand U1897 (N_1897,In_816,In_681);
nor U1898 (N_1898,In_966,In_513);
xnor U1899 (N_1899,In_924,In_596);
nor U1900 (N_1900,In_440,In_608);
or U1901 (N_1901,In_96,In_524);
and U1902 (N_1902,In_781,In_570);
nand U1903 (N_1903,In_912,In_88);
or U1904 (N_1904,In_203,In_24);
nor U1905 (N_1905,In_848,In_799);
and U1906 (N_1906,In_498,In_307);
or U1907 (N_1907,In_840,In_85);
and U1908 (N_1908,In_347,In_881);
nor U1909 (N_1909,In_988,In_354);
nor U1910 (N_1910,In_958,In_808);
nand U1911 (N_1911,In_477,In_787);
or U1912 (N_1912,In_781,In_233);
nand U1913 (N_1913,In_16,In_343);
or U1914 (N_1914,In_572,In_675);
and U1915 (N_1915,In_500,In_369);
or U1916 (N_1916,In_721,In_675);
nand U1917 (N_1917,In_43,In_410);
nand U1918 (N_1918,In_88,In_270);
and U1919 (N_1919,In_813,In_930);
nand U1920 (N_1920,In_227,In_407);
and U1921 (N_1921,In_451,In_905);
and U1922 (N_1922,In_431,In_659);
or U1923 (N_1923,In_487,In_894);
or U1924 (N_1924,In_987,In_937);
nand U1925 (N_1925,In_776,In_245);
nor U1926 (N_1926,In_16,In_858);
or U1927 (N_1927,In_600,In_902);
xor U1928 (N_1928,In_197,In_121);
and U1929 (N_1929,In_92,In_967);
or U1930 (N_1930,In_41,In_306);
nor U1931 (N_1931,In_326,In_725);
nand U1932 (N_1932,In_943,In_781);
nor U1933 (N_1933,In_446,In_453);
nor U1934 (N_1934,In_864,In_479);
or U1935 (N_1935,In_283,In_154);
or U1936 (N_1936,In_399,In_743);
and U1937 (N_1937,In_189,In_213);
nor U1938 (N_1938,In_750,In_265);
nor U1939 (N_1939,In_405,In_452);
and U1940 (N_1940,In_861,In_468);
nand U1941 (N_1941,In_175,In_176);
nor U1942 (N_1942,In_350,In_564);
and U1943 (N_1943,In_857,In_825);
nor U1944 (N_1944,In_0,In_259);
and U1945 (N_1945,In_212,In_844);
nor U1946 (N_1946,In_901,In_311);
nor U1947 (N_1947,In_359,In_583);
nor U1948 (N_1948,In_185,In_987);
or U1949 (N_1949,In_95,In_247);
or U1950 (N_1950,In_838,In_486);
or U1951 (N_1951,In_390,In_751);
nor U1952 (N_1952,In_214,In_206);
and U1953 (N_1953,In_470,In_374);
nor U1954 (N_1954,In_488,In_654);
or U1955 (N_1955,In_555,In_59);
nand U1956 (N_1956,In_991,In_621);
nor U1957 (N_1957,In_439,In_216);
nor U1958 (N_1958,In_216,In_774);
nand U1959 (N_1959,In_869,In_593);
nand U1960 (N_1960,In_203,In_563);
nand U1961 (N_1961,In_878,In_746);
nor U1962 (N_1962,In_150,In_609);
nor U1963 (N_1963,In_331,In_8);
nand U1964 (N_1964,In_415,In_105);
nor U1965 (N_1965,In_584,In_795);
and U1966 (N_1966,In_413,In_278);
or U1967 (N_1967,In_204,In_115);
nand U1968 (N_1968,In_610,In_4);
or U1969 (N_1969,In_826,In_707);
and U1970 (N_1970,In_466,In_885);
nor U1971 (N_1971,In_947,In_929);
nand U1972 (N_1972,In_6,In_868);
or U1973 (N_1973,In_997,In_101);
nand U1974 (N_1974,In_550,In_969);
or U1975 (N_1975,In_917,In_828);
nor U1976 (N_1976,In_731,In_243);
nand U1977 (N_1977,In_642,In_109);
nand U1978 (N_1978,In_548,In_179);
nor U1979 (N_1979,In_583,In_940);
nand U1980 (N_1980,In_130,In_765);
or U1981 (N_1981,In_996,In_989);
and U1982 (N_1982,In_867,In_978);
or U1983 (N_1983,In_155,In_669);
and U1984 (N_1984,In_274,In_605);
nand U1985 (N_1985,In_422,In_205);
nor U1986 (N_1986,In_18,In_206);
and U1987 (N_1987,In_719,In_564);
and U1988 (N_1988,In_641,In_656);
and U1989 (N_1989,In_287,In_266);
nor U1990 (N_1990,In_576,In_168);
or U1991 (N_1991,In_959,In_301);
nor U1992 (N_1992,In_681,In_608);
nor U1993 (N_1993,In_837,In_73);
nor U1994 (N_1994,In_692,In_381);
nand U1995 (N_1995,In_336,In_281);
xor U1996 (N_1996,In_527,In_745);
and U1997 (N_1997,In_231,In_959);
or U1998 (N_1998,In_290,In_998);
nand U1999 (N_1999,In_839,In_307);
and U2000 (N_2000,In_405,In_443);
xnor U2001 (N_2001,In_844,In_163);
nand U2002 (N_2002,In_100,In_478);
nor U2003 (N_2003,In_15,In_162);
nor U2004 (N_2004,In_655,In_747);
nand U2005 (N_2005,In_882,In_562);
and U2006 (N_2006,In_479,In_807);
or U2007 (N_2007,In_984,In_717);
or U2008 (N_2008,In_188,In_159);
or U2009 (N_2009,In_480,In_261);
nor U2010 (N_2010,In_354,In_263);
and U2011 (N_2011,In_124,In_11);
and U2012 (N_2012,In_995,In_226);
nand U2013 (N_2013,In_318,In_926);
nand U2014 (N_2014,In_893,In_560);
and U2015 (N_2015,In_853,In_870);
and U2016 (N_2016,In_141,In_381);
and U2017 (N_2017,In_494,In_256);
or U2018 (N_2018,In_962,In_680);
nor U2019 (N_2019,In_349,In_769);
and U2020 (N_2020,In_654,In_796);
nor U2021 (N_2021,In_697,In_293);
xor U2022 (N_2022,In_981,In_73);
nor U2023 (N_2023,In_285,In_491);
nor U2024 (N_2024,In_785,In_687);
nand U2025 (N_2025,In_67,In_729);
xor U2026 (N_2026,In_86,In_420);
nand U2027 (N_2027,In_588,In_991);
or U2028 (N_2028,In_399,In_999);
and U2029 (N_2029,In_714,In_866);
or U2030 (N_2030,In_783,In_403);
nor U2031 (N_2031,In_696,In_367);
nand U2032 (N_2032,In_997,In_152);
nor U2033 (N_2033,In_318,In_381);
nand U2034 (N_2034,In_177,In_410);
nor U2035 (N_2035,In_332,In_446);
and U2036 (N_2036,In_526,In_122);
nand U2037 (N_2037,In_988,In_539);
nand U2038 (N_2038,In_733,In_89);
and U2039 (N_2039,In_69,In_646);
nand U2040 (N_2040,In_675,In_604);
and U2041 (N_2041,In_539,In_240);
nor U2042 (N_2042,In_436,In_842);
nor U2043 (N_2043,In_30,In_893);
nor U2044 (N_2044,In_209,In_173);
xnor U2045 (N_2045,In_941,In_11);
and U2046 (N_2046,In_963,In_936);
nor U2047 (N_2047,In_436,In_427);
or U2048 (N_2048,In_343,In_137);
nor U2049 (N_2049,In_152,In_156);
nor U2050 (N_2050,In_401,In_989);
or U2051 (N_2051,In_294,In_406);
nand U2052 (N_2052,In_743,In_977);
nor U2053 (N_2053,In_823,In_708);
nand U2054 (N_2054,In_733,In_636);
nand U2055 (N_2055,In_842,In_548);
and U2056 (N_2056,In_769,In_885);
nand U2057 (N_2057,In_199,In_618);
and U2058 (N_2058,In_826,In_249);
nor U2059 (N_2059,In_142,In_950);
xnor U2060 (N_2060,In_881,In_669);
or U2061 (N_2061,In_311,In_526);
nand U2062 (N_2062,In_904,In_940);
nand U2063 (N_2063,In_386,In_655);
or U2064 (N_2064,In_224,In_468);
nand U2065 (N_2065,In_383,In_205);
nand U2066 (N_2066,In_857,In_356);
and U2067 (N_2067,In_561,In_1);
nor U2068 (N_2068,In_915,In_345);
nand U2069 (N_2069,In_831,In_86);
or U2070 (N_2070,In_622,In_325);
nand U2071 (N_2071,In_630,In_64);
or U2072 (N_2072,In_67,In_184);
and U2073 (N_2073,In_49,In_964);
and U2074 (N_2074,In_620,In_424);
or U2075 (N_2075,In_439,In_546);
nand U2076 (N_2076,In_891,In_755);
and U2077 (N_2077,In_369,In_750);
nand U2078 (N_2078,In_604,In_393);
nor U2079 (N_2079,In_806,In_359);
nand U2080 (N_2080,In_511,In_204);
nand U2081 (N_2081,In_528,In_44);
and U2082 (N_2082,In_259,In_944);
and U2083 (N_2083,In_314,In_335);
nor U2084 (N_2084,In_48,In_896);
nor U2085 (N_2085,In_355,In_3);
and U2086 (N_2086,In_255,In_569);
or U2087 (N_2087,In_418,In_87);
and U2088 (N_2088,In_592,In_825);
nand U2089 (N_2089,In_29,In_6);
xnor U2090 (N_2090,In_605,In_858);
or U2091 (N_2091,In_996,In_466);
xnor U2092 (N_2092,In_919,In_52);
nor U2093 (N_2093,In_290,In_898);
nor U2094 (N_2094,In_891,In_116);
nand U2095 (N_2095,In_318,In_124);
or U2096 (N_2096,In_469,In_398);
xnor U2097 (N_2097,In_53,In_872);
xnor U2098 (N_2098,In_612,In_687);
nand U2099 (N_2099,In_146,In_712);
and U2100 (N_2100,In_975,In_315);
and U2101 (N_2101,In_630,In_440);
and U2102 (N_2102,In_617,In_457);
nand U2103 (N_2103,In_252,In_264);
nor U2104 (N_2104,In_429,In_780);
nor U2105 (N_2105,In_13,In_782);
or U2106 (N_2106,In_552,In_241);
nor U2107 (N_2107,In_193,In_239);
or U2108 (N_2108,In_346,In_4);
or U2109 (N_2109,In_496,In_772);
nor U2110 (N_2110,In_757,In_944);
or U2111 (N_2111,In_520,In_437);
nor U2112 (N_2112,In_627,In_169);
or U2113 (N_2113,In_329,In_111);
nor U2114 (N_2114,In_962,In_625);
and U2115 (N_2115,In_183,In_118);
xor U2116 (N_2116,In_735,In_516);
nand U2117 (N_2117,In_854,In_409);
nand U2118 (N_2118,In_336,In_662);
and U2119 (N_2119,In_950,In_201);
nor U2120 (N_2120,In_408,In_270);
or U2121 (N_2121,In_967,In_329);
nor U2122 (N_2122,In_85,In_496);
or U2123 (N_2123,In_86,In_417);
or U2124 (N_2124,In_945,In_877);
nand U2125 (N_2125,In_980,In_327);
and U2126 (N_2126,In_324,In_903);
and U2127 (N_2127,In_21,In_179);
nand U2128 (N_2128,In_750,In_203);
nor U2129 (N_2129,In_179,In_549);
nor U2130 (N_2130,In_407,In_77);
nand U2131 (N_2131,In_953,In_102);
or U2132 (N_2132,In_457,In_494);
or U2133 (N_2133,In_544,In_53);
nor U2134 (N_2134,In_517,In_275);
or U2135 (N_2135,In_363,In_831);
nor U2136 (N_2136,In_646,In_706);
nor U2137 (N_2137,In_48,In_18);
nand U2138 (N_2138,In_11,In_903);
or U2139 (N_2139,In_467,In_772);
nor U2140 (N_2140,In_353,In_7);
and U2141 (N_2141,In_907,In_296);
and U2142 (N_2142,In_33,In_277);
or U2143 (N_2143,In_943,In_639);
nor U2144 (N_2144,In_660,In_394);
nand U2145 (N_2145,In_535,In_751);
nand U2146 (N_2146,In_574,In_387);
or U2147 (N_2147,In_977,In_468);
nor U2148 (N_2148,In_491,In_352);
nand U2149 (N_2149,In_883,In_414);
and U2150 (N_2150,In_620,In_8);
and U2151 (N_2151,In_383,In_350);
nor U2152 (N_2152,In_155,In_949);
nand U2153 (N_2153,In_240,In_914);
and U2154 (N_2154,In_106,In_273);
or U2155 (N_2155,In_780,In_165);
and U2156 (N_2156,In_616,In_149);
nand U2157 (N_2157,In_524,In_580);
and U2158 (N_2158,In_69,In_397);
nor U2159 (N_2159,In_706,In_801);
or U2160 (N_2160,In_66,In_273);
or U2161 (N_2161,In_653,In_869);
or U2162 (N_2162,In_796,In_876);
or U2163 (N_2163,In_665,In_159);
nor U2164 (N_2164,In_634,In_111);
nand U2165 (N_2165,In_726,In_91);
and U2166 (N_2166,In_571,In_102);
nand U2167 (N_2167,In_300,In_281);
and U2168 (N_2168,In_216,In_320);
nor U2169 (N_2169,In_820,In_189);
or U2170 (N_2170,In_100,In_954);
and U2171 (N_2171,In_84,In_166);
nor U2172 (N_2172,In_24,In_680);
nor U2173 (N_2173,In_276,In_196);
nand U2174 (N_2174,In_554,In_728);
and U2175 (N_2175,In_815,In_40);
and U2176 (N_2176,In_918,In_911);
and U2177 (N_2177,In_317,In_595);
and U2178 (N_2178,In_285,In_338);
nor U2179 (N_2179,In_843,In_879);
nand U2180 (N_2180,In_815,In_28);
nand U2181 (N_2181,In_111,In_181);
or U2182 (N_2182,In_724,In_607);
nor U2183 (N_2183,In_185,In_297);
nor U2184 (N_2184,In_536,In_7);
or U2185 (N_2185,In_818,In_384);
nand U2186 (N_2186,In_679,In_478);
nand U2187 (N_2187,In_901,In_644);
nor U2188 (N_2188,In_499,In_911);
or U2189 (N_2189,In_219,In_235);
nand U2190 (N_2190,In_461,In_863);
or U2191 (N_2191,In_362,In_996);
nand U2192 (N_2192,In_193,In_213);
nand U2193 (N_2193,In_494,In_855);
nand U2194 (N_2194,In_153,In_316);
and U2195 (N_2195,In_15,In_736);
nor U2196 (N_2196,In_781,In_95);
and U2197 (N_2197,In_158,In_222);
nand U2198 (N_2198,In_872,In_98);
nor U2199 (N_2199,In_394,In_150);
or U2200 (N_2200,In_677,In_473);
and U2201 (N_2201,In_196,In_894);
and U2202 (N_2202,In_447,In_816);
nand U2203 (N_2203,In_499,In_310);
and U2204 (N_2204,In_488,In_127);
nand U2205 (N_2205,In_590,In_99);
nor U2206 (N_2206,In_933,In_817);
nor U2207 (N_2207,In_421,In_646);
nand U2208 (N_2208,In_32,In_435);
and U2209 (N_2209,In_982,In_124);
and U2210 (N_2210,In_480,In_938);
nand U2211 (N_2211,In_432,In_166);
nor U2212 (N_2212,In_827,In_347);
or U2213 (N_2213,In_88,In_386);
nor U2214 (N_2214,In_83,In_688);
nor U2215 (N_2215,In_407,In_492);
and U2216 (N_2216,In_328,In_664);
nand U2217 (N_2217,In_591,In_6);
or U2218 (N_2218,In_806,In_494);
nand U2219 (N_2219,In_331,In_955);
and U2220 (N_2220,In_127,In_990);
and U2221 (N_2221,In_862,In_613);
or U2222 (N_2222,In_678,In_189);
nand U2223 (N_2223,In_146,In_35);
and U2224 (N_2224,In_574,In_149);
or U2225 (N_2225,In_286,In_666);
nor U2226 (N_2226,In_354,In_852);
or U2227 (N_2227,In_497,In_326);
nor U2228 (N_2228,In_719,In_900);
or U2229 (N_2229,In_491,In_662);
and U2230 (N_2230,In_334,In_462);
nor U2231 (N_2231,In_641,In_962);
and U2232 (N_2232,In_908,In_96);
or U2233 (N_2233,In_305,In_415);
nor U2234 (N_2234,In_799,In_941);
nor U2235 (N_2235,In_880,In_960);
nand U2236 (N_2236,In_643,In_565);
nand U2237 (N_2237,In_94,In_678);
nand U2238 (N_2238,In_515,In_580);
and U2239 (N_2239,In_845,In_561);
and U2240 (N_2240,In_765,In_449);
nand U2241 (N_2241,In_982,In_744);
or U2242 (N_2242,In_711,In_316);
nor U2243 (N_2243,In_942,In_948);
or U2244 (N_2244,In_856,In_809);
nor U2245 (N_2245,In_390,In_63);
and U2246 (N_2246,In_366,In_422);
nor U2247 (N_2247,In_485,In_441);
nor U2248 (N_2248,In_357,In_866);
xnor U2249 (N_2249,In_890,In_908);
nor U2250 (N_2250,In_295,In_287);
or U2251 (N_2251,In_577,In_832);
and U2252 (N_2252,In_133,In_997);
and U2253 (N_2253,In_337,In_447);
nor U2254 (N_2254,In_177,In_59);
or U2255 (N_2255,In_512,In_297);
or U2256 (N_2256,In_642,In_333);
nand U2257 (N_2257,In_846,In_392);
or U2258 (N_2258,In_542,In_884);
nor U2259 (N_2259,In_882,In_966);
and U2260 (N_2260,In_198,In_930);
and U2261 (N_2261,In_717,In_387);
and U2262 (N_2262,In_52,In_103);
and U2263 (N_2263,In_377,In_790);
nand U2264 (N_2264,In_749,In_305);
nand U2265 (N_2265,In_344,In_395);
or U2266 (N_2266,In_602,In_688);
nand U2267 (N_2267,In_412,In_38);
or U2268 (N_2268,In_532,In_272);
nand U2269 (N_2269,In_402,In_766);
or U2270 (N_2270,In_925,In_125);
and U2271 (N_2271,In_54,In_845);
or U2272 (N_2272,In_393,In_938);
and U2273 (N_2273,In_549,In_160);
and U2274 (N_2274,In_45,In_260);
or U2275 (N_2275,In_929,In_547);
nor U2276 (N_2276,In_313,In_964);
nor U2277 (N_2277,In_76,In_52);
and U2278 (N_2278,In_64,In_845);
or U2279 (N_2279,In_811,In_722);
or U2280 (N_2280,In_153,In_159);
or U2281 (N_2281,In_927,In_56);
nand U2282 (N_2282,In_110,In_178);
nor U2283 (N_2283,In_288,In_710);
and U2284 (N_2284,In_834,In_285);
nand U2285 (N_2285,In_379,In_429);
nand U2286 (N_2286,In_93,In_658);
nand U2287 (N_2287,In_847,In_245);
or U2288 (N_2288,In_384,In_511);
and U2289 (N_2289,In_343,In_313);
or U2290 (N_2290,In_659,In_688);
and U2291 (N_2291,In_114,In_814);
and U2292 (N_2292,In_100,In_31);
nand U2293 (N_2293,In_440,In_432);
nand U2294 (N_2294,In_505,In_808);
nand U2295 (N_2295,In_677,In_4);
or U2296 (N_2296,In_795,In_923);
and U2297 (N_2297,In_959,In_72);
nand U2298 (N_2298,In_613,In_989);
and U2299 (N_2299,In_159,In_861);
nand U2300 (N_2300,In_293,In_557);
nand U2301 (N_2301,In_837,In_58);
or U2302 (N_2302,In_782,In_556);
and U2303 (N_2303,In_964,In_105);
and U2304 (N_2304,In_887,In_692);
and U2305 (N_2305,In_279,In_511);
nor U2306 (N_2306,In_644,In_752);
and U2307 (N_2307,In_792,In_662);
nand U2308 (N_2308,In_557,In_387);
and U2309 (N_2309,In_338,In_362);
nor U2310 (N_2310,In_815,In_672);
or U2311 (N_2311,In_206,In_54);
nor U2312 (N_2312,In_840,In_97);
or U2313 (N_2313,In_1,In_883);
nand U2314 (N_2314,In_916,In_668);
nand U2315 (N_2315,In_646,In_629);
or U2316 (N_2316,In_964,In_345);
and U2317 (N_2317,In_951,In_275);
or U2318 (N_2318,In_789,In_229);
nor U2319 (N_2319,In_814,In_725);
and U2320 (N_2320,In_376,In_785);
nor U2321 (N_2321,In_432,In_829);
nand U2322 (N_2322,In_760,In_334);
and U2323 (N_2323,In_464,In_735);
nand U2324 (N_2324,In_175,In_238);
and U2325 (N_2325,In_603,In_625);
nand U2326 (N_2326,In_81,In_147);
nand U2327 (N_2327,In_901,In_396);
nand U2328 (N_2328,In_88,In_485);
nand U2329 (N_2329,In_889,In_269);
or U2330 (N_2330,In_217,In_529);
nand U2331 (N_2331,In_598,In_85);
and U2332 (N_2332,In_369,In_42);
and U2333 (N_2333,In_521,In_350);
or U2334 (N_2334,In_358,In_116);
or U2335 (N_2335,In_741,In_174);
nand U2336 (N_2336,In_458,In_587);
or U2337 (N_2337,In_94,In_581);
or U2338 (N_2338,In_697,In_872);
nand U2339 (N_2339,In_197,In_280);
or U2340 (N_2340,In_593,In_32);
or U2341 (N_2341,In_957,In_391);
nor U2342 (N_2342,In_366,In_946);
or U2343 (N_2343,In_879,In_915);
nand U2344 (N_2344,In_292,In_340);
nor U2345 (N_2345,In_720,In_848);
and U2346 (N_2346,In_417,In_78);
or U2347 (N_2347,In_853,In_533);
nor U2348 (N_2348,In_106,In_321);
and U2349 (N_2349,In_773,In_479);
nand U2350 (N_2350,In_191,In_390);
or U2351 (N_2351,In_724,In_787);
xnor U2352 (N_2352,In_480,In_631);
nand U2353 (N_2353,In_984,In_462);
nor U2354 (N_2354,In_587,In_455);
nor U2355 (N_2355,In_233,In_810);
or U2356 (N_2356,In_333,In_231);
nand U2357 (N_2357,In_538,In_95);
nor U2358 (N_2358,In_659,In_939);
xor U2359 (N_2359,In_151,In_503);
xnor U2360 (N_2360,In_912,In_210);
nor U2361 (N_2361,In_742,In_777);
nand U2362 (N_2362,In_735,In_567);
xnor U2363 (N_2363,In_930,In_833);
and U2364 (N_2364,In_1,In_81);
nor U2365 (N_2365,In_687,In_684);
or U2366 (N_2366,In_494,In_293);
and U2367 (N_2367,In_532,In_35);
nand U2368 (N_2368,In_27,In_775);
and U2369 (N_2369,In_479,In_255);
nor U2370 (N_2370,In_565,In_442);
or U2371 (N_2371,In_95,In_828);
and U2372 (N_2372,In_44,In_128);
and U2373 (N_2373,In_892,In_263);
or U2374 (N_2374,In_638,In_477);
nor U2375 (N_2375,In_263,In_144);
xnor U2376 (N_2376,In_388,In_361);
nand U2377 (N_2377,In_498,In_295);
and U2378 (N_2378,In_270,In_227);
nor U2379 (N_2379,In_930,In_465);
nor U2380 (N_2380,In_34,In_638);
and U2381 (N_2381,In_336,In_692);
or U2382 (N_2382,In_512,In_572);
nor U2383 (N_2383,In_594,In_93);
or U2384 (N_2384,In_702,In_905);
nor U2385 (N_2385,In_825,In_868);
nor U2386 (N_2386,In_516,In_111);
or U2387 (N_2387,In_321,In_488);
or U2388 (N_2388,In_18,In_963);
nor U2389 (N_2389,In_904,In_199);
and U2390 (N_2390,In_669,In_581);
nand U2391 (N_2391,In_357,In_468);
nor U2392 (N_2392,In_823,In_990);
and U2393 (N_2393,In_19,In_201);
and U2394 (N_2394,In_735,In_228);
nand U2395 (N_2395,In_127,In_270);
or U2396 (N_2396,In_820,In_774);
and U2397 (N_2397,In_971,In_144);
and U2398 (N_2398,In_638,In_292);
nand U2399 (N_2399,In_849,In_6);
and U2400 (N_2400,In_866,In_302);
nor U2401 (N_2401,In_468,In_188);
and U2402 (N_2402,In_142,In_964);
nor U2403 (N_2403,In_529,In_787);
nand U2404 (N_2404,In_908,In_530);
and U2405 (N_2405,In_52,In_463);
nor U2406 (N_2406,In_595,In_677);
nand U2407 (N_2407,In_549,In_519);
or U2408 (N_2408,In_435,In_304);
nor U2409 (N_2409,In_756,In_308);
nand U2410 (N_2410,In_241,In_892);
and U2411 (N_2411,In_799,In_111);
nor U2412 (N_2412,In_935,In_267);
nor U2413 (N_2413,In_550,In_582);
and U2414 (N_2414,In_936,In_201);
nor U2415 (N_2415,In_644,In_80);
nor U2416 (N_2416,In_747,In_841);
nor U2417 (N_2417,In_251,In_292);
nand U2418 (N_2418,In_294,In_879);
or U2419 (N_2419,In_144,In_258);
and U2420 (N_2420,In_444,In_745);
nor U2421 (N_2421,In_166,In_747);
and U2422 (N_2422,In_314,In_783);
nand U2423 (N_2423,In_996,In_577);
or U2424 (N_2424,In_819,In_121);
nand U2425 (N_2425,In_79,In_917);
or U2426 (N_2426,In_892,In_817);
nand U2427 (N_2427,In_616,In_533);
nor U2428 (N_2428,In_11,In_506);
or U2429 (N_2429,In_544,In_688);
and U2430 (N_2430,In_100,In_536);
or U2431 (N_2431,In_773,In_213);
and U2432 (N_2432,In_750,In_400);
nand U2433 (N_2433,In_186,In_377);
nand U2434 (N_2434,In_750,In_792);
or U2435 (N_2435,In_238,In_367);
or U2436 (N_2436,In_274,In_322);
nand U2437 (N_2437,In_437,In_875);
nor U2438 (N_2438,In_739,In_967);
or U2439 (N_2439,In_556,In_172);
nor U2440 (N_2440,In_671,In_163);
and U2441 (N_2441,In_581,In_217);
and U2442 (N_2442,In_541,In_292);
nand U2443 (N_2443,In_608,In_689);
or U2444 (N_2444,In_395,In_415);
or U2445 (N_2445,In_656,In_984);
or U2446 (N_2446,In_960,In_380);
and U2447 (N_2447,In_745,In_854);
nand U2448 (N_2448,In_361,In_637);
and U2449 (N_2449,In_368,In_962);
nor U2450 (N_2450,In_840,In_668);
xnor U2451 (N_2451,In_808,In_959);
nand U2452 (N_2452,In_198,In_185);
or U2453 (N_2453,In_999,In_761);
nor U2454 (N_2454,In_314,In_22);
nor U2455 (N_2455,In_322,In_34);
nor U2456 (N_2456,In_935,In_535);
nand U2457 (N_2457,In_286,In_455);
and U2458 (N_2458,In_513,In_23);
nand U2459 (N_2459,In_275,In_157);
or U2460 (N_2460,In_149,In_878);
or U2461 (N_2461,In_133,In_30);
xor U2462 (N_2462,In_176,In_792);
and U2463 (N_2463,In_510,In_792);
or U2464 (N_2464,In_189,In_941);
and U2465 (N_2465,In_816,In_763);
or U2466 (N_2466,In_551,In_678);
and U2467 (N_2467,In_308,In_198);
nor U2468 (N_2468,In_765,In_597);
nand U2469 (N_2469,In_738,In_607);
and U2470 (N_2470,In_55,In_637);
xor U2471 (N_2471,In_514,In_358);
and U2472 (N_2472,In_218,In_650);
or U2473 (N_2473,In_910,In_360);
nor U2474 (N_2474,In_499,In_731);
nand U2475 (N_2475,In_105,In_493);
or U2476 (N_2476,In_105,In_996);
nor U2477 (N_2477,In_988,In_609);
nor U2478 (N_2478,In_585,In_71);
xor U2479 (N_2479,In_172,In_635);
nor U2480 (N_2480,In_692,In_361);
or U2481 (N_2481,In_734,In_749);
or U2482 (N_2482,In_364,In_887);
or U2483 (N_2483,In_752,In_742);
nor U2484 (N_2484,In_276,In_375);
nor U2485 (N_2485,In_470,In_619);
nand U2486 (N_2486,In_338,In_321);
xor U2487 (N_2487,In_186,In_341);
xor U2488 (N_2488,In_342,In_526);
nor U2489 (N_2489,In_290,In_157);
nor U2490 (N_2490,In_13,In_286);
or U2491 (N_2491,In_497,In_916);
and U2492 (N_2492,In_506,In_663);
or U2493 (N_2493,In_203,In_177);
or U2494 (N_2494,In_71,In_746);
nor U2495 (N_2495,In_526,In_404);
and U2496 (N_2496,In_869,In_549);
and U2497 (N_2497,In_73,In_474);
or U2498 (N_2498,In_762,In_473);
or U2499 (N_2499,In_405,In_821);
and U2500 (N_2500,In_862,In_276);
nor U2501 (N_2501,In_332,In_139);
and U2502 (N_2502,In_931,In_152);
and U2503 (N_2503,In_55,In_837);
xnor U2504 (N_2504,In_775,In_376);
and U2505 (N_2505,In_645,In_513);
nor U2506 (N_2506,In_424,In_570);
or U2507 (N_2507,In_812,In_528);
or U2508 (N_2508,In_727,In_700);
nand U2509 (N_2509,In_311,In_862);
or U2510 (N_2510,In_25,In_6);
and U2511 (N_2511,In_554,In_84);
and U2512 (N_2512,In_103,In_791);
and U2513 (N_2513,In_422,In_913);
xnor U2514 (N_2514,In_78,In_770);
nand U2515 (N_2515,In_389,In_511);
or U2516 (N_2516,In_834,In_185);
nand U2517 (N_2517,In_592,In_855);
nand U2518 (N_2518,In_175,In_191);
nor U2519 (N_2519,In_805,In_395);
or U2520 (N_2520,In_253,In_731);
nor U2521 (N_2521,In_988,In_799);
nor U2522 (N_2522,In_458,In_410);
and U2523 (N_2523,In_963,In_749);
nand U2524 (N_2524,In_463,In_310);
xnor U2525 (N_2525,In_309,In_487);
or U2526 (N_2526,In_146,In_644);
or U2527 (N_2527,In_306,In_785);
nand U2528 (N_2528,In_311,In_988);
nor U2529 (N_2529,In_611,In_38);
nor U2530 (N_2530,In_503,In_856);
or U2531 (N_2531,In_19,In_607);
nor U2532 (N_2532,In_935,In_294);
nor U2533 (N_2533,In_776,In_838);
nor U2534 (N_2534,In_576,In_951);
nand U2535 (N_2535,In_437,In_39);
nor U2536 (N_2536,In_758,In_518);
nor U2537 (N_2537,In_149,In_833);
nor U2538 (N_2538,In_109,In_400);
or U2539 (N_2539,In_675,In_708);
nand U2540 (N_2540,In_540,In_704);
nand U2541 (N_2541,In_399,In_875);
or U2542 (N_2542,In_300,In_366);
and U2543 (N_2543,In_84,In_381);
nor U2544 (N_2544,In_970,In_383);
or U2545 (N_2545,In_936,In_389);
and U2546 (N_2546,In_774,In_307);
or U2547 (N_2547,In_212,In_20);
or U2548 (N_2548,In_898,In_330);
nand U2549 (N_2549,In_852,In_70);
or U2550 (N_2550,In_197,In_427);
nand U2551 (N_2551,In_291,In_20);
nand U2552 (N_2552,In_548,In_530);
or U2553 (N_2553,In_395,In_15);
nor U2554 (N_2554,In_617,In_936);
nand U2555 (N_2555,In_868,In_331);
and U2556 (N_2556,In_862,In_2);
or U2557 (N_2557,In_37,In_640);
and U2558 (N_2558,In_901,In_48);
nand U2559 (N_2559,In_556,In_287);
nand U2560 (N_2560,In_439,In_176);
and U2561 (N_2561,In_212,In_278);
and U2562 (N_2562,In_795,In_123);
or U2563 (N_2563,In_438,In_640);
nand U2564 (N_2564,In_982,In_360);
and U2565 (N_2565,In_901,In_268);
and U2566 (N_2566,In_925,In_105);
and U2567 (N_2567,In_652,In_828);
nand U2568 (N_2568,In_796,In_703);
or U2569 (N_2569,In_566,In_433);
nor U2570 (N_2570,In_313,In_544);
nor U2571 (N_2571,In_641,In_559);
nor U2572 (N_2572,In_608,In_731);
nor U2573 (N_2573,In_643,In_446);
nor U2574 (N_2574,In_58,In_152);
or U2575 (N_2575,In_945,In_120);
nand U2576 (N_2576,In_139,In_216);
and U2577 (N_2577,In_180,In_328);
or U2578 (N_2578,In_157,In_521);
and U2579 (N_2579,In_522,In_512);
nor U2580 (N_2580,In_210,In_369);
or U2581 (N_2581,In_88,In_467);
or U2582 (N_2582,In_833,In_136);
or U2583 (N_2583,In_533,In_132);
nor U2584 (N_2584,In_784,In_226);
nand U2585 (N_2585,In_382,In_444);
and U2586 (N_2586,In_956,In_898);
nor U2587 (N_2587,In_980,In_307);
or U2588 (N_2588,In_31,In_57);
or U2589 (N_2589,In_290,In_762);
or U2590 (N_2590,In_96,In_972);
and U2591 (N_2591,In_66,In_713);
and U2592 (N_2592,In_482,In_623);
nor U2593 (N_2593,In_760,In_444);
or U2594 (N_2594,In_99,In_350);
nand U2595 (N_2595,In_606,In_374);
nor U2596 (N_2596,In_609,In_558);
nor U2597 (N_2597,In_177,In_151);
or U2598 (N_2598,In_140,In_461);
nor U2599 (N_2599,In_812,In_310);
nor U2600 (N_2600,In_323,In_283);
or U2601 (N_2601,In_287,In_677);
and U2602 (N_2602,In_598,In_934);
or U2603 (N_2603,In_960,In_596);
nor U2604 (N_2604,In_552,In_742);
xnor U2605 (N_2605,In_954,In_432);
or U2606 (N_2606,In_347,In_943);
or U2607 (N_2607,In_832,In_793);
nor U2608 (N_2608,In_928,In_657);
or U2609 (N_2609,In_924,In_605);
or U2610 (N_2610,In_876,In_647);
nor U2611 (N_2611,In_96,In_243);
or U2612 (N_2612,In_277,In_837);
or U2613 (N_2613,In_306,In_296);
nand U2614 (N_2614,In_981,In_110);
or U2615 (N_2615,In_368,In_353);
or U2616 (N_2616,In_711,In_90);
nor U2617 (N_2617,In_435,In_517);
nand U2618 (N_2618,In_151,In_737);
nor U2619 (N_2619,In_737,In_745);
and U2620 (N_2620,In_638,In_605);
nor U2621 (N_2621,In_954,In_243);
nor U2622 (N_2622,In_123,In_139);
or U2623 (N_2623,In_246,In_522);
nand U2624 (N_2624,In_209,In_926);
and U2625 (N_2625,In_440,In_29);
and U2626 (N_2626,In_515,In_335);
and U2627 (N_2627,In_642,In_612);
nand U2628 (N_2628,In_299,In_646);
and U2629 (N_2629,In_997,In_467);
nand U2630 (N_2630,In_642,In_487);
and U2631 (N_2631,In_105,In_116);
and U2632 (N_2632,In_872,In_759);
and U2633 (N_2633,In_158,In_658);
and U2634 (N_2634,In_0,In_836);
nand U2635 (N_2635,In_850,In_733);
xor U2636 (N_2636,In_425,In_227);
and U2637 (N_2637,In_902,In_528);
or U2638 (N_2638,In_532,In_419);
nand U2639 (N_2639,In_275,In_716);
or U2640 (N_2640,In_993,In_444);
or U2641 (N_2641,In_644,In_248);
nor U2642 (N_2642,In_962,In_697);
or U2643 (N_2643,In_400,In_498);
nor U2644 (N_2644,In_313,In_915);
or U2645 (N_2645,In_843,In_523);
nand U2646 (N_2646,In_4,In_77);
or U2647 (N_2647,In_169,In_141);
and U2648 (N_2648,In_542,In_737);
and U2649 (N_2649,In_771,In_229);
nand U2650 (N_2650,In_140,In_758);
nor U2651 (N_2651,In_11,In_414);
or U2652 (N_2652,In_624,In_808);
and U2653 (N_2653,In_291,In_200);
or U2654 (N_2654,In_773,In_200);
or U2655 (N_2655,In_566,In_824);
nand U2656 (N_2656,In_46,In_566);
nand U2657 (N_2657,In_768,In_868);
nand U2658 (N_2658,In_175,In_196);
nand U2659 (N_2659,In_710,In_163);
nor U2660 (N_2660,In_759,In_269);
nand U2661 (N_2661,In_44,In_560);
or U2662 (N_2662,In_394,In_848);
or U2663 (N_2663,In_201,In_867);
nand U2664 (N_2664,In_893,In_680);
nor U2665 (N_2665,In_465,In_740);
nor U2666 (N_2666,In_519,In_382);
or U2667 (N_2667,In_354,In_396);
and U2668 (N_2668,In_232,In_333);
or U2669 (N_2669,In_803,In_538);
or U2670 (N_2670,In_681,In_316);
or U2671 (N_2671,In_102,In_75);
or U2672 (N_2672,In_242,In_253);
and U2673 (N_2673,In_18,In_512);
nor U2674 (N_2674,In_829,In_127);
nand U2675 (N_2675,In_918,In_711);
and U2676 (N_2676,In_406,In_318);
and U2677 (N_2677,In_517,In_623);
nand U2678 (N_2678,In_581,In_87);
and U2679 (N_2679,In_594,In_123);
nand U2680 (N_2680,In_263,In_406);
or U2681 (N_2681,In_553,In_746);
or U2682 (N_2682,In_622,In_895);
xor U2683 (N_2683,In_487,In_683);
and U2684 (N_2684,In_522,In_528);
nand U2685 (N_2685,In_719,In_481);
and U2686 (N_2686,In_156,In_107);
or U2687 (N_2687,In_596,In_393);
nand U2688 (N_2688,In_490,In_83);
nor U2689 (N_2689,In_828,In_964);
and U2690 (N_2690,In_509,In_126);
nor U2691 (N_2691,In_540,In_966);
or U2692 (N_2692,In_692,In_608);
or U2693 (N_2693,In_173,In_214);
and U2694 (N_2694,In_72,In_799);
nand U2695 (N_2695,In_255,In_127);
or U2696 (N_2696,In_140,In_849);
and U2697 (N_2697,In_865,In_69);
nor U2698 (N_2698,In_660,In_884);
or U2699 (N_2699,In_122,In_590);
nand U2700 (N_2700,In_781,In_4);
nand U2701 (N_2701,In_250,In_365);
and U2702 (N_2702,In_476,In_543);
nand U2703 (N_2703,In_866,In_726);
nor U2704 (N_2704,In_54,In_244);
nand U2705 (N_2705,In_917,In_628);
nand U2706 (N_2706,In_602,In_638);
nand U2707 (N_2707,In_797,In_431);
nand U2708 (N_2708,In_179,In_774);
nor U2709 (N_2709,In_785,In_580);
nor U2710 (N_2710,In_77,In_71);
or U2711 (N_2711,In_382,In_464);
or U2712 (N_2712,In_637,In_820);
and U2713 (N_2713,In_647,In_934);
and U2714 (N_2714,In_877,In_778);
or U2715 (N_2715,In_150,In_285);
nand U2716 (N_2716,In_334,In_756);
and U2717 (N_2717,In_294,In_374);
and U2718 (N_2718,In_498,In_817);
nand U2719 (N_2719,In_192,In_805);
nor U2720 (N_2720,In_903,In_963);
and U2721 (N_2721,In_217,In_371);
nand U2722 (N_2722,In_737,In_992);
or U2723 (N_2723,In_8,In_636);
nand U2724 (N_2724,In_765,In_247);
nor U2725 (N_2725,In_419,In_817);
and U2726 (N_2726,In_658,In_214);
or U2727 (N_2727,In_203,In_97);
nand U2728 (N_2728,In_232,In_725);
nand U2729 (N_2729,In_459,In_538);
or U2730 (N_2730,In_429,In_948);
nand U2731 (N_2731,In_991,In_262);
nand U2732 (N_2732,In_507,In_104);
nor U2733 (N_2733,In_555,In_811);
nand U2734 (N_2734,In_133,In_597);
or U2735 (N_2735,In_255,In_570);
or U2736 (N_2736,In_884,In_832);
or U2737 (N_2737,In_218,In_548);
or U2738 (N_2738,In_903,In_482);
or U2739 (N_2739,In_754,In_618);
nand U2740 (N_2740,In_509,In_966);
or U2741 (N_2741,In_578,In_848);
and U2742 (N_2742,In_370,In_393);
and U2743 (N_2743,In_410,In_745);
nor U2744 (N_2744,In_209,In_169);
nand U2745 (N_2745,In_286,In_929);
or U2746 (N_2746,In_364,In_130);
and U2747 (N_2747,In_811,In_679);
or U2748 (N_2748,In_770,In_20);
nand U2749 (N_2749,In_105,In_109);
or U2750 (N_2750,In_366,In_502);
nand U2751 (N_2751,In_923,In_375);
nor U2752 (N_2752,In_177,In_450);
and U2753 (N_2753,In_116,In_611);
nor U2754 (N_2754,In_890,In_793);
nand U2755 (N_2755,In_7,In_916);
and U2756 (N_2756,In_255,In_728);
or U2757 (N_2757,In_994,In_802);
and U2758 (N_2758,In_604,In_711);
or U2759 (N_2759,In_602,In_388);
and U2760 (N_2760,In_268,In_927);
nand U2761 (N_2761,In_189,In_483);
or U2762 (N_2762,In_888,In_785);
or U2763 (N_2763,In_227,In_178);
or U2764 (N_2764,In_216,In_166);
and U2765 (N_2765,In_662,In_468);
xor U2766 (N_2766,In_99,In_108);
and U2767 (N_2767,In_452,In_611);
and U2768 (N_2768,In_768,In_746);
or U2769 (N_2769,In_427,In_247);
and U2770 (N_2770,In_67,In_630);
or U2771 (N_2771,In_4,In_393);
or U2772 (N_2772,In_456,In_204);
or U2773 (N_2773,In_342,In_181);
or U2774 (N_2774,In_408,In_170);
nand U2775 (N_2775,In_364,In_533);
nand U2776 (N_2776,In_649,In_625);
nor U2777 (N_2777,In_20,In_638);
xnor U2778 (N_2778,In_467,In_141);
nor U2779 (N_2779,In_530,In_748);
nor U2780 (N_2780,In_404,In_593);
nand U2781 (N_2781,In_582,In_916);
nor U2782 (N_2782,In_843,In_997);
nor U2783 (N_2783,In_836,In_516);
and U2784 (N_2784,In_353,In_32);
nand U2785 (N_2785,In_557,In_220);
or U2786 (N_2786,In_797,In_280);
nand U2787 (N_2787,In_814,In_304);
and U2788 (N_2788,In_18,In_712);
nor U2789 (N_2789,In_630,In_903);
and U2790 (N_2790,In_706,In_794);
and U2791 (N_2791,In_214,In_959);
and U2792 (N_2792,In_632,In_930);
or U2793 (N_2793,In_971,In_242);
nand U2794 (N_2794,In_335,In_212);
nand U2795 (N_2795,In_266,In_762);
nand U2796 (N_2796,In_756,In_626);
or U2797 (N_2797,In_557,In_534);
nand U2798 (N_2798,In_800,In_692);
and U2799 (N_2799,In_48,In_353);
and U2800 (N_2800,In_84,In_431);
and U2801 (N_2801,In_484,In_916);
nand U2802 (N_2802,In_906,In_69);
nand U2803 (N_2803,In_202,In_67);
and U2804 (N_2804,In_269,In_934);
nor U2805 (N_2805,In_223,In_315);
nand U2806 (N_2806,In_142,In_806);
and U2807 (N_2807,In_179,In_424);
nor U2808 (N_2808,In_655,In_902);
nor U2809 (N_2809,In_937,In_301);
nand U2810 (N_2810,In_287,In_228);
and U2811 (N_2811,In_339,In_36);
and U2812 (N_2812,In_572,In_890);
nand U2813 (N_2813,In_941,In_42);
and U2814 (N_2814,In_610,In_40);
or U2815 (N_2815,In_55,In_892);
or U2816 (N_2816,In_419,In_617);
and U2817 (N_2817,In_897,In_593);
nand U2818 (N_2818,In_221,In_781);
nand U2819 (N_2819,In_280,In_290);
nand U2820 (N_2820,In_527,In_567);
and U2821 (N_2821,In_274,In_63);
or U2822 (N_2822,In_304,In_997);
and U2823 (N_2823,In_221,In_346);
xor U2824 (N_2824,In_299,In_730);
nand U2825 (N_2825,In_524,In_55);
nand U2826 (N_2826,In_475,In_127);
and U2827 (N_2827,In_961,In_387);
nand U2828 (N_2828,In_106,In_150);
or U2829 (N_2829,In_480,In_666);
or U2830 (N_2830,In_70,In_391);
and U2831 (N_2831,In_413,In_805);
or U2832 (N_2832,In_431,In_739);
and U2833 (N_2833,In_705,In_279);
xor U2834 (N_2834,In_953,In_161);
nand U2835 (N_2835,In_358,In_190);
and U2836 (N_2836,In_262,In_333);
or U2837 (N_2837,In_375,In_210);
nand U2838 (N_2838,In_472,In_238);
and U2839 (N_2839,In_911,In_831);
nand U2840 (N_2840,In_783,In_252);
and U2841 (N_2841,In_203,In_347);
xor U2842 (N_2842,In_438,In_332);
and U2843 (N_2843,In_877,In_878);
nor U2844 (N_2844,In_374,In_476);
nand U2845 (N_2845,In_558,In_85);
nand U2846 (N_2846,In_720,In_766);
or U2847 (N_2847,In_690,In_950);
or U2848 (N_2848,In_856,In_222);
or U2849 (N_2849,In_377,In_248);
and U2850 (N_2850,In_574,In_567);
nand U2851 (N_2851,In_318,In_4);
nand U2852 (N_2852,In_659,In_254);
nand U2853 (N_2853,In_160,In_454);
nand U2854 (N_2854,In_883,In_880);
nand U2855 (N_2855,In_5,In_676);
nand U2856 (N_2856,In_865,In_241);
nand U2857 (N_2857,In_627,In_508);
or U2858 (N_2858,In_240,In_653);
and U2859 (N_2859,In_851,In_205);
nor U2860 (N_2860,In_975,In_656);
and U2861 (N_2861,In_781,In_819);
and U2862 (N_2862,In_534,In_976);
or U2863 (N_2863,In_939,In_586);
nor U2864 (N_2864,In_948,In_532);
or U2865 (N_2865,In_710,In_282);
and U2866 (N_2866,In_700,In_373);
and U2867 (N_2867,In_706,In_992);
nand U2868 (N_2868,In_659,In_580);
or U2869 (N_2869,In_710,In_191);
or U2870 (N_2870,In_749,In_375);
or U2871 (N_2871,In_779,In_370);
nor U2872 (N_2872,In_564,In_836);
nor U2873 (N_2873,In_765,In_916);
nand U2874 (N_2874,In_480,In_854);
and U2875 (N_2875,In_566,In_315);
and U2876 (N_2876,In_312,In_778);
nor U2877 (N_2877,In_919,In_447);
and U2878 (N_2878,In_321,In_208);
and U2879 (N_2879,In_189,In_57);
nor U2880 (N_2880,In_902,In_470);
xor U2881 (N_2881,In_269,In_72);
nand U2882 (N_2882,In_128,In_255);
nand U2883 (N_2883,In_503,In_30);
nand U2884 (N_2884,In_474,In_505);
nor U2885 (N_2885,In_926,In_456);
and U2886 (N_2886,In_449,In_84);
xor U2887 (N_2887,In_524,In_128);
nor U2888 (N_2888,In_658,In_648);
or U2889 (N_2889,In_596,In_54);
and U2890 (N_2890,In_562,In_37);
and U2891 (N_2891,In_703,In_422);
and U2892 (N_2892,In_36,In_327);
and U2893 (N_2893,In_776,In_610);
nand U2894 (N_2894,In_326,In_644);
nand U2895 (N_2895,In_260,In_889);
nand U2896 (N_2896,In_282,In_791);
nor U2897 (N_2897,In_360,In_313);
nand U2898 (N_2898,In_786,In_503);
or U2899 (N_2899,In_439,In_958);
nor U2900 (N_2900,In_120,In_583);
nand U2901 (N_2901,In_940,In_592);
or U2902 (N_2902,In_980,In_259);
nand U2903 (N_2903,In_361,In_971);
and U2904 (N_2904,In_981,In_511);
and U2905 (N_2905,In_782,In_212);
nor U2906 (N_2906,In_888,In_408);
and U2907 (N_2907,In_255,In_606);
nand U2908 (N_2908,In_378,In_207);
nor U2909 (N_2909,In_809,In_70);
and U2910 (N_2910,In_545,In_194);
nand U2911 (N_2911,In_931,In_861);
nand U2912 (N_2912,In_443,In_217);
and U2913 (N_2913,In_778,In_787);
or U2914 (N_2914,In_488,In_673);
nand U2915 (N_2915,In_592,In_406);
nor U2916 (N_2916,In_570,In_811);
nand U2917 (N_2917,In_807,In_227);
xnor U2918 (N_2918,In_693,In_252);
or U2919 (N_2919,In_439,In_171);
nand U2920 (N_2920,In_806,In_787);
or U2921 (N_2921,In_90,In_183);
or U2922 (N_2922,In_704,In_492);
and U2923 (N_2923,In_852,In_251);
nand U2924 (N_2924,In_808,In_815);
nor U2925 (N_2925,In_502,In_40);
and U2926 (N_2926,In_279,In_18);
nor U2927 (N_2927,In_298,In_369);
nor U2928 (N_2928,In_832,In_648);
or U2929 (N_2929,In_178,In_290);
nand U2930 (N_2930,In_975,In_986);
nor U2931 (N_2931,In_601,In_815);
or U2932 (N_2932,In_392,In_717);
and U2933 (N_2933,In_747,In_982);
nand U2934 (N_2934,In_272,In_124);
or U2935 (N_2935,In_947,In_733);
and U2936 (N_2936,In_377,In_360);
nor U2937 (N_2937,In_14,In_865);
nor U2938 (N_2938,In_937,In_879);
and U2939 (N_2939,In_239,In_359);
nand U2940 (N_2940,In_290,In_364);
nor U2941 (N_2941,In_759,In_595);
nor U2942 (N_2942,In_835,In_787);
nand U2943 (N_2943,In_254,In_26);
or U2944 (N_2944,In_731,In_819);
nand U2945 (N_2945,In_176,In_620);
or U2946 (N_2946,In_541,In_274);
nand U2947 (N_2947,In_602,In_372);
nor U2948 (N_2948,In_876,In_68);
or U2949 (N_2949,In_690,In_459);
or U2950 (N_2950,In_432,In_152);
nand U2951 (N_2951,In_100,In_188);
nor U2952 (N_2952,In_122,In_485);
nand U2953 (N_2953,In_851,In_565);
and U2954 (N_2954,In_186,In_830);
or U2955 (N_2955,In_105,In_460);
or U2956 (N_2956,In_328,In_232);
and U2957 (N_2957,In_184,In_913);
or U2958 (N_2958,In_577,In_62);
nor U2959 (N_2959,In_65,In_129);
and U2960 (N_2960,In_518,In_536);
and U2961 (N_2961,In_793,In_441);
and U2962 (N_2962,In_698,In_758);
nor U2963 (N_2963,In_895,In_676);
and U2964 (N_2964,In_763,In_151);
nor U2965 (N_2965,In_460,In_674);
and U2966 (N_2966,In_234,In_688);
nor U2967 (N_2967,In_171,In_133);
and U2968 (N_2968,In_468,In_887);
or U2969 (N_2969,In_176,In_618);
or U2970 (N_2970,In_335,In_874);
nand U2971 (N_2971,In_247,In_799);
or U2972 (N_2972,In_566,In_569);
nor U2973 (N_2973,In_401,In_583);
or U2974 (N_2974,In_875,In_941);
nor U2975 (N_2975,In_754,In_350);
or U2976 (N_2976,In_349,In_408);
nand U2977 (N_2977,In_747,In_907);
or U2978 (N_2978,In_13,In_845);
nand U2979 (N_2979,In_305,In_267);
xnor U2980 (N_2980,In_455,In_468);
or U2981 (N_2981,In_932,In_780);
and U2982 (N_2982,In_82,In_614);
and U2983 (N_2983,In_715,In_378);
or U2984 (N_2984,In_351,In_521);
and U2985 (N_2985,In_7,In_691);
or U2986 (N_2986,In_328,In_845);
and U2987 (N_2987,In_481,In_209);
nand U2988 (N_2988,In_451,In_405);
and U2989 (N_2989,In_990,In_269);
or U2990 (N_2990,In_338,In_552);
nand U2991 (N_2991,In_405,In_892);
nor U2992 (N_2992,In_373,In_188);
nor U2993 (N_2993,In_151,In_515);
nor U2994 (N_2994,In_721,In_745);
or U2995 (N_2995,In_884,In_500);
nor U2996 (N_2996,In_826,In_406);
nor U2997 (N_2997,In_924,In_358);
and U2998 (N_2998,In_484,In_657);
and U2999 (N_2999,In_421,In_58);
nand U3000 (N_3000,In_602,In_496);
nand U3001 (N_3001,In_834,In_585);
xor U3002 (N_3002,In_87,In_323);
or U3003 (N_3003,In_98,In_454);
or U3004 (N_3004,In_416,In_692);
and U3005 (N_3005,In_542,In_995);
and U3006 (N_3006,In_311,In_849);
and U3007 (N_3007,In_970,In_53);
nand U3008 (N_3008,In_427,In_701);
and U3009 (N_3009,In_889,In_511);
or U3010 (N_3010,In_167,In_402);
and U3011 (N_3011,In_938,In_365);
xor U3012 (N_3012,In_4,In_731);
nor U3013 (N_3013,In_761,In_779);
or U3014 (N_3014,In_21,In_883);
nand U3015 (N_3015,In_948,In_399);
nand U3016 (N_3016,In_861,In_621);
and U3017 (N_3017,In_908,In_415);
and U3018 (N_3018,In_36,In_228);
nor U3019 (N_3019,In_261,In_965);
nand U3020 (N_3020,In_806,In_301);
nand U3021 (N_3021,In_59,In_849);
and U3022 (N_3022,In_233,In_167);
and U3023 (N_3023,In_371,In_534);
and U3024 (N_3024,In_658,In_185);
and U3025 (N_3025,In_981,In_33);
nand U3026 (N_3026,In_867,In_906);
nor U3027 (N_3027,In_508,In_716);
and U3028 (N_3028,In_948,In_750);
or U3029 (N_3029,In_893,In_460);
nand U3030 (N_3030,In_290,In_807);
nor U3031 (N_3031,In_720,In_479);
nand U3032 (N_3032,In_80,In_432);
nor U3033 (N_3033,In_373,In_974);
nor U3034 (N_3034,In_11,In_989);
or U3035 (N_3035,In_254,In_114);
nand U3036 (N_3036,In_379,In_889);
nor U3037 (N_3037,In_823,In_996);
and U3038 (N_3038,In_729,In_205);
nor U3039 (N_3039,In_639,In_783);
and U3040 (N_3040,In_469,In_995);
and U3041 (N_3041,In_870,In_275);
or U3042 (N_3042,In_811,In_655);
and U3043 (N_3043,In_194,In_779);
nor U3044 (N_3044,In_463,In_841);
and U3045 (N_3045,In_493,In_350);
nor U3046 (N_3046,In_834,In_544);
and U3047 (N_3047,In_280,In_38);
and U3048 (N_3048,In_710,In_40);
nor U3049 (N_3049,In_129,In_147);
or U3050 (N_3050,In_621,In_378);
nand U3051 (N_3051,In_103,In_994);
nand U3052 (N_3052,In_766,In_852);
nand U3053 (N_3053,In_745,In_457);
or U3054 (N_3054,In_652,In_17);
and U3055 (N_3055,In_705,In_96);
nand U3056 (N_3056,In_810,In_632);
nand U3057 (N_3057,In_962,In_303);
or U3058 (N_3058,In_852,In_416);
nor U3059 (N_3059,In_731,In_895);
and U3060 (N_3060,In_177,In_221);
xnor U3061 (N_3061,In_920,In_149);
nand U3062 (N_3062,In_381,In_619);
or U3063 (N_3063,In_241,In_447);
nand U3064 (N_3064,In_212,In_16);
and U3065 (N_3065,In_321,In_677);
nand U3066 (N_3066,In_696,In_145);
and U3067 (N_3067,In_494,In_120);
nand U3068 (N_3068,In_243,In_573);
nand U3069 (N_3069,In_202,In_835);
nand U3070 (N_3070,In_331,In_725);
or U3071 (N_3071,In_167,In_987);
and U3072 (N_3072,In_760,In_423);
nand U3073 (N_3073,In_965,In_761);
nand U3074 (N_3074,In_844,In_38);
nand U3075 (N_3075,In_129,In_934);
or U3076 (N_3076,In_791,In_825);
or U3077 (N_3077,In_218,In_939);
or U3078 (N_3078,In_694,In_962);
and U3079 (N_3079,In_933,In_418);
nor U3080 (N_3080,In_72,In_397);
and U3081 (N_3081,In_68,In_987);
nand U3082 (N_3082,In_453,In_343);
or U3083 (N_3083,In_600,In_519);
and U3084 (N_3084,In_299,In_264);
xnor U3085 (N_3085,In_567,In_990);
and U3086 (N_3086,In_710,In_364);
nor U3087 (N_3087,In_181,In_672);
xor U3088 (N_3088,In_79,In_635);
xnor U3089 (N_3089,In_628,In_700);
and U3090 (N_3090,In_436,In_929);
nor U3091 (N_3091,In_381,In_812);
and U3092 (N_3092,In_343,In_160);
or U3093 (N_3093,In_612,In_985);
or U3094 (N_3094,In_971,In_325);
xnor U3095 (N_3095,In_130,In_943);
and U3096 (N_3096,In_668,In_889);
nand U3097 (N_3097,In_197,In_582);
nor U3098 (N_3098,In_524,In_75);
nand U3099 (N_3099,In_134,In_282);
or U3100 (N_3100,In_7,In_333);
or U3101 (N_3101,In_418,In_519);
nor U3102 (N_3102,In_824,In_467);
or U3103 (N_3103,In_284,In_386);
nand U3104 (N_3104,In_294,In_288);
or U3105 (N_3105,In_191,In_722);
and U3106 (N_3106,In_818,In_959);
and U3107 (N_3107,In_760,In_309);
and U3108 (N_3108,In_794,In_613);
nor U3109 (N_3109,In_516,In_534);
and U3110 (N_3110,In_529,In_899);
or U3111 (N_3111,In_111,In_896);
nor U3112 (N_3112,In_476,In_123);
nor U3113 (N_3113,In_776,In_641);
or U3114 (N_3114,In_347,In_718);
or U3115 (N_3115,In_786,In_142);
and U3116 (N_3116,In_279,In_171);
and U3117 (N_3117,In_350,In_70);
nor U3118 (N_3118,In_905,In_729);
nand U3119 (N_3119,In_912,In_822);
nand U3120 (N_3120,In_915,In_580);
nand U3121 (N_3121,In_571,In_837);
nand U3122 (N_3122,In_857,In_13);
or U3123 (N_3123,In_533,In_32);
nand U3124 (N_3124,In_655,In_222);
and U3125 (N_3125,In_805,In_460);
nor U3126 (N_3126,In_891,In_876);
and U3127 (N_3127,In_912,In_556);
or U3128 (N_3128,In_304,In_787);
or U3129 (N_3129,In_816,In_945);
nor U3130 (N_3130,In_466,In_624);
nand U3131 (N_3131,In_918,In_319);
or U3132 (N_3132,In_950,In_420);
nand U3133 (N_3133,In_625,In_321);
and U3134 (N_3134,In_518,In_983);
nor U3135 (N_3135,In_96,In_790);
or U3136 (N_3136,In_801,In_820);
nand U3137 (N_3137,In_139,In_114);
or U3138 (N_3138,In_712,In_417);
nand U3139 (N_3139,In_557,In_196);
and U3140 (N_3140,In_421,In_868);
and U3141 (N_3141,In_293,In_969);
nand U3142 (N_3142,In_637,In_988);
nor U3143 (N_3143,In_774,In_569);
nand U3144 (N_3144,In_797,In_937);
xnor U3145 (N_3145,In_737,In_305);
or U3146 (N_3146,In_147,In_818);
nor U3147 (N_3147,In_632,In_604);
nor U3148 (N_3148,In_909,In_438);
and U3149 (N_3149,In_575,In_933);
nor U3150 (N_3150,In_697,In_389);
nor U3151 (N_3151,In_552,In_655);
or U3152 (N_3152,In_790,In_944);
and U3153 (N_3153,In_193,In_409);
nand U3154 (N_3154,In_352,In_877);
nand U3155 (N_3155,In_994,In_287);
and U3156 (N_3156,In_748,In_493);
nand U3157 (N_3157,In_787,In_631);
and U3158 (N_3158,In_907,In_500);
and U3159 (N_3159,In_230,In_916);
nand U3160 (N_3160,In_700,In_832);
and U3161 (N_3161,In_153,In_711);
nand U3162 (N_3162,In_330,In_126);
and U3163 (N_3163,In_769,In_742);
and U3164 (N_3164,In_47,In_586);
nand U3165 (N_3165,In_168,In_728);
and U3166 (N_3166,In_243,In_946);
nand U3167 (N_3167,In_547,In_350);
nor U3168 (N_3168,In_891,In_747);
and U3169 (N_3169,In_113,In_337);
or U3170 (N_3170,In_148,In_653);
and U3171 (N_3171,In_20,In_236);
nand U3172 (N_3172,In_652,In_358);
and U3173 (N_3173,In_352,In_749);
or U3174 (N_3174,In_701,In_500);
nand U3175 (N_3175,In_233,In_208);
and U3176 (N_3176,In_641,In_259);
nand U3177 (N_3177,In_894,In_686);
nor U3178 (N_3178,In_663,In_552);
and U3179 (N_3179,In_200,In_114);
and U3180 (N_3180,In_568,In_624);
nor U3181 (N_3181,In_228,In_365);
nand U3182 (N_3182,In_770,In_558);
or U3183 (N_3183,In_576,In_66);
nand U3184 (N_3184,In_557,In_233);
nand U3185 (N_3185,In_431,In_907);
nor U3186 (N_3186,In_937,In_752);
and U3187 (N_3187,In_600,In_803);
nand U3188 (N_3188,In_275,In_512);
nand U3189 (N_3189,In_191,In_537);
or U3190 (N_3190,In_533,In_509);
nor U3191 (N_3191,In_13,In_245);
or U3192 (N_3192,In_540,In_437);
nor U3193 (N_3193,In_360,In_144);
and U3194 (N_3194,In_302,In_898);
or U3195 (N_3195,In_93,In_980);
nor U3196 (N_3196,In_582,In_566);
or U3197 (N_3197,In_433,In_645);
nand U3198 (N_3198,In_181,In_232);
nor U3199 (N_3199,In_877,In_40);
or U3200 (N_3200,In_674,In_104);
or U3201 (N_3201,In_444,In_103);
nor U3202 (N_3202,In_372,In_960);
and U3203 (N_3203,In_725,In_485);
nor U3204 (N_3204,In_77,In_768);
nand U3205 (N_3205,In_420,In_497);
nor U3206 (N_3206,In_576,In_865);
nand U3207 (N_3207,In_355,In_680);
and U3208 (N_3208,In_14,In_932);
or U3209 (N_3209,In_201,In_548);
or U3210 (N_3210,In_172,In_53);
or U3211 (N_3211,In_466,In_628);
nor U3212 (N_3212,In_59,In_346);
or U3213 (N_3213,In_750,In_202);
and U3214 (N_3214,In_190,In_539);
and U3215 (N_3215,In_563,In_216);
or U3216 (N_3216,In_85,In_522);
or U3217 (N_3217,In_578,In_661);
nor U3218 (N_3218,In_892,In_901);
nand U3219 (N_3219,In_452,In_315);
and U3220 (N_3220,In_529,In_187);
nand U3221 (N_3221,In_836,In_747);
nor U3222 (N_3222,In_646,In_803);
nand U3223 (N_3223,In_138,In_685);
and U3224 (N_3224,In_575,In_446);
nand U3225 (N_3225,In_640,In_870);
or U3226 (N_3226,In_196,In_24);
and U3227 (N_3227,In_432,In_477);
and U3228 (N_3228,In_549,In_233);
nor U3229 (N_3229,In_943,In_777);
xnor U3230 (N_3230,In_332,In_881);
and U3231 (N_3231,In_193,In_408);
nand U3232 (N_3232,In_495,In_575);
nor U3233 (N_3233,In_706,In_144);
nor U3234 (N_3234,In_989,In_885);
and U3235 (N_3235,In_767,In_196);
or U3236 (N_3236,In_48,In_871);
and U3237 (N_3237,In_633,In_26);
nand U3238 (N_3238,In_4,In_743);
and U3239 (N_3239,In_265,In_505);
and U3240 (N_3240,In_339,In_797);
or U3241 (N_3241,In_343,In_595);
nand U3242 (N_3242,In_191,In_405);
nor U3243 (N_3243,In_580,In_686);
nand U3244 (N_3244,In_9,In_972);
or U3245 (N_3245,In_435,In_610);
nor U3246 (N_3246,In_94,In_729);
xnor U3247 (N_3247,In_307,In_724);
nand U3248 (N_3248,In_205,In_506);
nor U3249 (N_3249,In_170,In_619);
nand U3250 (N_3250,In_338,In_438);
nand U3251 (N_3251,In_38,In_241);
and U3252 (N_3252,In_292,In_270);
or U3253 (N_3253,In_186,In_974);
nand U3254 (N_3254,In_303,In_805);
nand U3255 (N_3255,In_123,In_861);
and U3256 (N_3256,In_111,In_481);
and U3257 (N_3257,In_862,In_39);
nor U3258 (N_3258,In_28,In_907);
nand U3259 (N_3259,In_112,In_582);
nor U3260 (N_3260,In_140,In_276);
or U3261 (N_3261,In_337,In_301);
nor U3262 (N_3262,In_678,In_939);
and U3263 (N_3263,In_108,In_903);
nor U3264 (N_3264,In_396,In_738);
nand U3265 (N_3265,In_175,In_45);
or U3266 (N_3266,In_307,In_757);
nand U3267 (N_3267,In_722,In_502);
or U3268 (N_3268,In_65,In_716);
or U3269 (N_3269,In_108,In_832);
nand U3270 (N_3270,In_866,In_870);
and U3271 (N_3271,In_869,In_381);
nand U3272 (N_3272,In_34,In_33);
nor U3273 (N_3273,In_243,In_758);
nor U3274 (N_3274,In_693,In_156);
nand U3275 (N_3275,In_366,In_179);
and U3276 (N_3276,In_321,In_588);
or U3277 (N_3277,In_800,In_638);
and U3278 (N_3278,In_903,In_891);
nor U3279 (N_3279,In_517,In_94);
nand U3280 (N_3280,In_670,In_519);
nor U3281 (N_3281,In_752,In_717);
nand U3282 (N_3282,In_813,In_670);
or U3283 (N_3283,In_184,In_618);
or U3284 (N_3284,In_480,In_278);
or U3285 (N_3285,In_447,In_583);
nand U3286 (N_3286,In_945,In_641);
nand U3287 (N_3287,In_536,In_669);
and U3288 (N_3288,In_461,In_920);
nor U3289 (N_3289,In_957,In_207);
nor U3290 (N_3290,In_611,In_681);
nor U3291 (N_3291,In_107,In_877);
nor U3292 (N_3292,In_776,In_77);
nor U3293 (N_3293,In_13,In_780);
nor U3294 (N_3294,In_220,In_806);
nor U3295 (N_3295,In_691,In_829);
nor U3296 (N_3296,In_593,In_222);
nor U3297 (N_3297,In_934,In_304);
and U3298 (N_3298,In_71,In_203);
or U3299 (N_3299,In_718,In_215);
xor U3300 (N_3300,In_281,In_456);
and U3301 (N_3301,In_914,In_130);
and U3302 (N_3302,In_780,In_53);
and U3303 (N_3303,In_296,In_318);
or U3304 (N_3304,In_305,In_5);
and U3305 (N_3305,In_257,In_400);
or U3306 (N_3306,In_774,In_734);
or U3307 (N_3307,In_110,In_142);
nor U3308 (N_3308,In_544,In_973);
nor U3309 (N_3309,In_671,In_810);
and U3310 (N_3310,In_163,In_852);
or U3311 (N_3311,In_309,In_130);
or U3312 (N_3312,In_270,In_2);
or U3313 (N_3313,In_383,In_922);
or U3314 (N_3314,In_866,In_261);
nand U3315 (N_3315,In_797,In_698);
and U3316 (N_3316,In_398,In_366);
nand U3317 (N_3317,In_556,In_20);
nor U3318 (N_3318,In_124,In_515);
or U3319 (N_3319,In_756,In_643);
or U3320 (N_3320,In_186,In_154);
xor U3321 (N_3321,In_161,In_332);
nand U3322 (N_3322,In_490,In_689);
and U3323 (N_3323,In_628,In_985);
nand U3324 (N_3324,In_146,In_886);
nor U3325 (N_3325,In_595,In_513);
and U3326 (N_3326,In_136,In_224);
and U3327 (N_3327,In_114,In_609);
nor U3328 (N_3328,In_819,In_568);
nor U3329 (N_3329,In_926,In_580);
and U3330 (N_3330,In_896,In_304);
and U3331 (N_3331,In_586,In_903);
nand U3332 (N_3332,In_51,In_439);
or U3333 (N_3333,In_285,In_534);
nand U3334 (N_3334,In_677,In_523);
nor U3335 (N_3335,In_379,In_701);
or U3336 (N_3336,In_468,In_645);
or U3337 (N_3337,In_74,In_674);
nor U3338 (N_3338,In_984,In_603);
nand U3339 (N_3339,In_2,In_776);
nor U3340 (N_3340,In_349,In_851);
or U3341 (N_3341,In_790,In_467);
nand U3342 (N_3342,In_297,In_116);
and U3343 (N_3343,In_229,In_652);
and U3344 (N_3344,In_535,In_669);
or U3345 (N_3345,In_434,In_572);
and U3346 (N_3346,In_48,In_187);
nor U3347 (N_3347,In_76,In_946);
nand U3348 (N_3348,In_578,In_765);
nand U3349 (N_3349,In_823,In_260);
xor U3350 (N_3350,In_923,In_919);
and U3351 (N_3351,In_248,In_108);
nand U3352 (N_3352,In_593,In_867);
nor U3353 (N_3353,In_759,In_859);
and U3354 (N_3354,In_497,In_788);
nand U3355 (N_3355,In_305,In_798);
and U3356 (N_3356,In_943,In_752);
nand U3357 (N_3357,In_303,In_232);
and U3358 (N_3358,In_436,In_219);
nand U3359 (N_3359,In_35,In_201);
or U3360 (N_3360,In_947,In_718);
nand U3361 (N_3361,In_103,In_500);
nor U3362 (N_3362,In_369,In_474);
and U3363 (N_3363,In_522,In_357);
or U3364 (N_3364,In_926,In_539);
or U3365 (N_3365,In_738,In_610);
nor U3366 (N_3366,In_575,In_322);
nor U3367 (N_3367,In_297,In_207);
nand U3368 (N_3368,In_432,In_562);
or U3369 (N_3369,In_671,In_197);
nand U3370 (N_3370,In_948,In_499);
or U3371 (N_3371,In_938,In_187);
and U3372 (N_3372,In_328,In_819);
and U3373 (N_3373,In_71,In_387);
nand U3374 (N_3374,In_935,In_62);
nand U3375 (N_3375,In_735,In_672);
nand U3376 (N_3376,In_236,In_306);
or U3377 (N_3377,In_788,In_164);
or U3378 (N_3378,In_259,In_466);
nand U3379 (N_3379,In_793,In_138);
nand U3380 (N_3380,In_666,In_855);
nor U3381 (N_3381,In_853,In_786);
nor U3382 (N_3382,In_187,In_7);
xnor U3383 (N_3383,In_318,In_817);
nor U3384 (N_3384,In_309,In_537);
nor U3385 (N_3385,In_664,In_777);
nor U3386 (N_3386,In_406,In_473);
or U3387 (N_3387,In_922,In_625);
and U3388 (N_3388,In_523,In_793);
nor U3389 (N_3389,In_63,In_662);
and U3390 (N_3390,In_83,In_998);
nand U3391 (N_3391,In_47,In_773);
and U3392 (N_3392,In_372,In_699);
or U3393 (N_3393,In_675,In_941);
and U3394 (N_3394,In_885,In_100);
or U3395 (N_3395,In_640,In_586);
nand U3396 (N_3396,In_273,In_219);
nand U3397 (N_3397,In_282,In_232);
and U3398 (N_3398,In_272,In_699);
nor U3399 (N_3399,In_663,In_460);
and U3400 (N_3400,In_326,In_336);
nand U3401 (N_3401,In_276,In_128);
or U3402 (N_3402,In_459,In_677);
nor U3403 (N_3403,In_656,In_275);
and U3404 (N_3404,In_572,In_382);
and U3405 (N_3405,In_868,In_976);
or U3406 (N_3406,In_688,In_379);
nor U3407 (N_3407,In_343,In_745);
nor U3408 (N_3408,In_388,In_748);
nor U3409 (N_3409,In_395,In_310);
and U3410 (N_3410,In_715,In_987);
nor U3411 (N_3411,In_603,In_203);
or U3412 (N_3412,In_520,In_550);
or U3413 (N_3413,In_731,In_931);
nor U3414 (N_3414,In_118,In_339);
nor U3415 (N_3415,In_2,In_670);
and U3416 (N_3416,In_592,In_158);
nand U3417 (N_3417,In_258,In_190);
xnor U3418 (N_3418,In_250,In_880);
nand U3419 (N_3419,In_865,In_309);
xnor U3420 (N_3420,In_672,In_679);
nor U3421 (N_3421,In_237,In_823);
xnor U3422 (N_3422,In_338,In_40);
and U3423 (N_3423,In_310,In_567);
and U3424 (N_3424,In_845,In_324);
nor U3425 (N_3425,In_929,In_817);
or U3426 (N_3426,In_997,In_131);
or U3427 (N_3427,In_110,In_600);
and U3428 (N_3428,In_900,In_73);
nor U3429 (N_3429,In_39,In_883);
or U3430 (N_3430,In_633,In_988);
nand U3431 (N_3431,In_410,In_233);
nor U3432 (N_3432,In_28,In_83);
or U3433 (N_3433,In_889,In_291);
or U3434 (N_3434,In_891,In_631);
nor U3435 (N_3435,In_24,In_559);
nand U3436 (N_3436,In_279,In_34);
or U3437 (N_3437,In_30,In_238);
and U3438 (N_3438,In_608,In_730);
xor U3439 (N_3439,In_795,In_527);
and U3440 (N_3440,In_373,In_404);
nor U3441 (N_3441,In_637,In_25);
or U3442 (N_3442,In_486,In_914);
and U3443 (N_3443,In_187,In_50);
or U3444 (N_3444,In_865,In_664);
nor U3445 (N_3445,In_339,In_678);
nand U3446 (N_3446,In_963,In_645);
nand U3447 (N_3447,In_777,In_936);
xor U3448 (N_3448,In_154,In_655);
nor U3449 (N_3449,In_954,In_346);
nor U3450 (N_3450,In_59,In_738);
nor U3451 (N_3451,In_140,In_275);
or U3452 (N_3452,In_827,In_220);
xnor U3453 (N_3453,In_704,In_464);
nand U3454 (N_3454,In_159,In_706);
nor U3455 (N_3455,In_810,In_851);
nand U3456 (N_3456,In_348,In_434);
or U3457 (N_3457,In_875,In_600);
nand U3458 (N_3458,In_248,In_442);
or U3459 (N_3459,In_362,In_256);
nand U3460 (N_3460,In_64,In_551);
and U3461 (N_3461,In_432,In_538);
or U3462 (N_3462,In_202,In_191);
nor U3463 (N_3463,In_70,In_872);
and U3464 (N_3464,In_74,In_864);
and U3465 (N_3465,In_910,In_443);
or U3466 (N_3466,In_81,In_727);
nand U3467 (N_3467,In_391,In_805);
nand U3468 (N_3468,In_631,In_845);
nand U3469 (N_3469,In_470,In_632);
nand U3470 (N_3470,In_98,In_518);
nor U3471 (N_3471,In_792,In_491);
nand U3472 (N_3472,In_674,In_775);
nor U3473 (N_3473,In_686,In_524);
nand U3474 (N_3474,In_966,In_580);
nor U3475 (N_3475,In_345,In_608);
and U3476 (N_3476,In_962,In_530);
or U3477 (N_3477,In_983,In_556);
xnor U3478 (N_3478,In_879,In_373);
or U3479 (N_3479,In_562,In_42);
nand U3480 (N_3480,In_952,In_65);
nand U3481 (N_3481,In_479,In_615);
nand U3482 (N_3482,In_718,In_873);
nor U3483 (N_3483,In_844,In_486);
or U3484 (N_3484,In_183,In_1);
or U3485 (N_3485,In_56,In_235);
nand U3486 (N_3486,In_493,In_741);
or U3487 (N_3487,In_981,In_372);
nor U3488 (N_3488,In_823,In_879);
or U3489 (N_3489,In_644,In_224);
nor U3490 (N_3490,In_45,In_346);
or U3491 (N_3491,In_80,In_989);
nand U3492 (N_3492,In_319,In_880);
nand U3493 (N_3493,In_247,In_139);
and U3494 (N_3494,In_768,In_226);
or U3495 (N_3495,In_575,In_170);
or U3496 (N_3496,In_20,In_336);
and U3497 (N_3497,In_904,In_447);
and U3498 (N_3498,In_282,In_334);
nand U3499 (N_3499,In_159,In_17);
nor U3500 (N_3500,In_948,In_730);
nor U3501 (N_3501,In_816,In_568);
nor U3502 (N_3502,In_238,In_900);
and U3503 (N_3503,In_542,In_744);
nand U3504 (N_3504,In_383,In_279);
or U3505 (N_3505,In_13,In_505);
nor U3506 (N_3506,In_498,In_649);
and U3507 (N_3507,In_917,In_143);
and U3508 (N_3508,In_102,In_584);
and U3509 (N_3509,In_202,In_514);
nand U3510 (N_3510,In_84,In_775);
nor U3511 (N_3511,In_294,In_793);
or U3512 (N_3512,In_87,In_535);
nand U3513 (N_3513,In_251,In_188);
nor U3514 (N_3514,In_604,In_421);
nor U3515 (N_3515,In_364,In_745);
xnor U3516 (N_3516,In_103,In_804);
nor U3517 (N_3517,In_920,In_2);
and U3518 (N_3518,In_972,In_587);
and U3519 (N_3519,In_192,In_629);
nor U3520 (N_3520,In_583,In_796);
nand U3521 (N_3521,In_897,In_947);
nor U3522 (N_3522,In_975,In_700);
and U3523 (N_3523,In_799,In_240);
and U3524 (N_3524,In_946,In_530);
nand U3525 (N_3525,In_797,In_649);
nand U3526 (N_3526,In_740,In_295);
and U3527 (N_3527,In_763,In_426);
and U3528 (N_3528,In_580,In_943);
nand U3529 (N_3529,In_619,In_38);
nand U3530 (N_3530,In_145,In_567);
nand U3531 (N_3531,In_649,In_777);
or U3532 (N_3532,In_854,In_876);
or U3533 (N_3533,In_534,In_127);
and U3534 (N_3534,In_725,In_483);
or U3535 (N_3535,In_834,In_690);
nor U3536 (N_3536,In_637,In_549);
or U3537 (N_3537,In_478,In_571);
nor U3538 (N_3538,In_272,In_677);
nand U3539 (N_3539,In_31,In_507);
nor U3540 (N_3540,In_149,In_282);
nand U3541 (N_3541,In_541,In_697);
or U3542 (N_3542,In_820,In_497);
nand U3543 (N_3543,In_703,In_939);
or U3544 (N_3544,In_260,In_178);
or U3545 (N_3545,In_760,In_415);
or U3546 (N_3546,In_669,In_236);
xnor U3547 (N_3547,In_748,In_681);
or U3548 (N_3548,In_356,In_838);
nand U3549 (N_3549,In_302,In_691);
nor U3550 (N_3550,In_671,In_970);
xnor U3551 (N_3551,In_275,In_308);
or U3552 (N_3552,In_528,In_139);
and U3553 (N_3553,In_29,In_873);
or U3554 (N_3554,In_465,In_3);
nand U3555 (N_3555,In_706,In_67);
or U3556 (N_3556,In_994,In_760);
or U3557 (N_3557,In_991,In_574);
nor U3558 (N_3558,In_698,In_470);
nand U3559 (N_3559,In_76,In_416);
nand U3560 (N_3560,In_91,In_676);
or U3561 (N_3561,In_584,In_319);
nand U3562 (N_3562,In_979,In_973);
or U3563 (N_3563,In_339,In_410);
nor U3564 (N_3564,In_153,In_986);
nand U3565 (N_3565,In_658,In_99);
nand U3566 (N_3566,In_310,In_397);
nor U3567 (N_3567,In_405,In_693);
nor U3568 (N_3568,In_75,In_928);
nor U3569 (N_3569,In_366,In_807);
and U3570 (N_3570,In_178,In_429);
or U3571 (N_3571,In_571,In_489);
xor U3572 (N_3572,In_682,In_614);
or U3573 (N_3573,In_755,In_837);
or U3574 (N_3574,In_639,In_108);
and U3575 (N_3575,In_724,In_145);
or U3576 (N_3576,In_62,In_20);
nor U3577 (N_3577,In_393,In_150);
and U3578 (N_3578,In_404,In_647);
and U3579 (N_3579,In_895,In_534);
and U3580 (N_3580,In_38,In_357);
nand U3581 (N_3581,In_196,In_208);
nand U3582 (N_3582,In_1,In_148);
nand U3583 (N_3583,In_114,In_950);
and U3584 (N_3584,In_178,In_226);
and U3585 (N_3585,In_367,In_592);
and U3586 (N_3586,In_817,In_327);
or U3587 (N_3587,In_859,In_725);
and U3588 (N_3588,In_600,In_520);
nand U3589 (N_3589,In_878,In_711);
nor U3590 (N_3590,In_655,In_494);
nand U3591 (N_3591,In_710,In_560);
or U3592 (N_3592,In_599,In_694);
nor U3593 (N_3593,In_281,In_333);
nor U3594 (N_3594,In_629,In_516);
or U3595 (N_3595,In_571,In_410);
nor U3596 (N_3596,In_483,In_863);
or U3597 (N_3597,In_152,In_653);
nand U3598 (N_3598,In_735,In_463);
nor U3599 (N_3599,In_236,In_302);
nor U3600 (N_3600,In_146,In_964);
or U3601 (N_3601,In_514,In_392);
nand U3602 (N_3602,In_915,In_458);
nor U3603 (N_3603,In_420,In_263);
nor U3604 (N_3604,In_370,In_570);
and U3605 (N_3605,In_539,In_968);
nand U3606 (N_3606,In_337,In_679);
nand U3607 (N_3607,In_568,In_884);
nor U3608 (N_3608,In_131,In_578);
and U3609 (N_3609,In_62,In_29);
nor U3610 (N_3610,In_705,In_765);
or U3611 (N_3611,In_220,In_777);
xor U3612 (N_3612,In_893,In_807);
nand U3613 (N_3613,In_704,In_992);
and U3614 (N_3614,In_355,In_856);
nor U3615 (N_3615,In_545,In_527);
nand U3616 (N_3616,In_497,In_368);
nand U3617 (N_3617,In_775,In_766);
or U3618 (N_3618,In_648,In_785);
nand U3619 (N_3619,In_286,In_484);
or U3620 (N_3620,In_141,In_152);
nor U3621 (N_3621,In_879,In_771);
nand U3622 (N_3622,In_734,In_213);
nand U3623 (N_3623,In_456,In_642);
or U3624 (N_3624,In_569,In_536);
and U3625 (N_3625,In_314,In_323);
or U3626 (N_3626,In_781,In_62);
nor U3627 (N_3627,In_45,In_347);
xor U3628 (N_3628,In_305,In_903);
xnor U3629 (N_3629,In_900,In_134);
nor U3630 (N_3630,In_341,In_583);
and U3631 (N_3631,In_896,In_577);
nor U3632 (N_3632,In_533,In_165);
xnor U3633 (N_3633,In_443,In_680);
nand U3634 (N_3634,In_792,In_511);
xor U3635 (N_3635,In_953,In_447);
or U3636 (N_3636,In_180,In_960);
nand U3637 (N_3637,In_131,In_24);
nor U3638 (N_3638,In_351,In_219);
nor U3639 (N_3639,In_527,In_997);
nor U3640 (N_3640,In_443,In_663);
nor U3641 (N_3641,In_667,In_881);
nor U3642 (N_3642,In_573,In_323);
and U3643 (N_3643,In_211,In_124);
nor U3644 (N_3644,In_482,In_655);
or U3645 (N_3645,In_418,In_679);
and U3646 (N_3646,In_733,In_743);
nand U3647 (N_3647,In_944,In_634);
nor U3648 (N_3648,In_649,In_708);
nor U3649 (N_3649,In_88,In_596);
or U3650 (N_3650,In_873,In_310);
or U3651 (N_3651,In_37,In_941);
or U3652 (N_3652,In_456,In_188);
nor U3653 (N_3653,In_623,In_635);
nor U3654 (N_3654,In_767,In_72);
or U3655 (N_3655,In_707,In_981);
nor U3656 (N_3656,In_559,In_222);
and U3657 (N_3657,In_821,In_642);
and U3658 (N_3658,In_210,In_378);
and U3659 (N_3659,In_318,In_755);
nand U3660 (N_3660,In_445,In_908);
nor U3661 (N_3661,In_734,In_740);
nand U3662 (N_3662,In_753,In_759);
or U3663 (N_3663,In_487,In_720);
nor U3664 (N_3664,In_224,In_191);
or U3665 (N_3665,In_472,In_868);
nor U3666 (N_3666,In_100,In_112);
nor U3667 (N_3667,In_754,In_485);
xnor U3668 (N_3668,In_718,In_220);
or U3669 (N_3669,In_431,In_812);
or U3670 (N_3670,In_399,In_28);
nand U3671 (N_3671,In_351,In_504);
nor U3672 (N_3672,In_256,In_468);
nor U3673 (N_3673,In_38,In_3);
or U3674 (N_3674,In_130,In_901);
nor U3675 (N_3675,In_369,In_910);
xor U3676 (N_3676,In_84,In_41);
and U3677 (N_3677,In_69,In_87);
nor U3678 (N_3678,In_225,In_33);
and U3679 (N_3679,In_565,In_469);
nand U3680 (N_3680,In_95,In_871);
nand U3681 (N_3681,In_147,In_552);
nand U3682 (N_3682,In_279,In_55);
nor U3683 (N_3683,In_794,In_333);
and U3684 (N_3684,In_192,In_452);
nor U3685 (N_3685,In_472,In_422);
or U3686 (N_3686,In_317,In_274);
and U3687 (N_3687,In_767,In_40);
or U3688 (N_3688,In_609,In_457);
nand U3689 (N_3689,In_447,In_647);
or U3690 (N_3690,In_485,In_285);
nor U3691 (N_3691,In_968,In_170);
and U3692 (N_3692,In_21,In_969);
nand U3693 (N_3693,In_947,In_24);
nand U3694 (N_3694,In_842,In_507);
nand U3695 (N_3695,In_397,In_108);
or U3696 (N_3696,In_516,In_146);
nand U3697 (N_3697,In_414,In_898);
nand U3698 (N_3698,In_698,In_859);
or U3699 (N_3699,In_64,In_805);
nand U3700 (N_3700,In_976,In_580);
and U3701 (N_3701,In_161,In_891);
nand U3702 (N_3702,In_380,In_244);
nor U3703 (N_3703,In_58,In_922);
nor U3704 (N_3704,In_548,In_334);
nand U3705 (N_3705,In_563,In_955);
nand U3706 (N_3706,In_708,In_204);
nor U3707 (N_3707,In_308,In_929);
nor U3708 (N_3708,In_133,In_852);
or U3709 (N_3709,In_292,In_483);
nor U3710 (N_3710,In_926,In_125);
xor U3711 (N_3711,In_555,In_961);
or U3712 (N_3712,In_341,In_668);
or U3713 (N_3713,In_703,In_600);
or U3714 (N_3714,In_503,In_141);
nand U3715 (N_3715,In_693,In_591);
or U3716 (N_3716,In_754,In_772);
nor U3717 (N_3717,In_639,In_92);
and U3718 (N_3718,In_859,In_992);
or U3719 (N_3719,In_323,In_143);
nand U3720 (N_3720,In_675,In_826);
and U3721 (N_3721,In_372,In_492);
or U3722 (N_3722,In_605,In_676);
nand U3723 (N_3723,In_993,In_312);
and U3724 (N_3724,In_707,In_803);
nor U3725 (N_3725,In_333,In_426);
nor U3726 (N_3726,In_274,In_468);
or U3727 (N_3727,In_816,In_209);
nand U3728 (N_3728,In_39,In_713);
xnor U3729 (N_3729,In_369,In_161);
and U3730 (N_3730,In_528,In_625);
nand U3731 (N_3731,In_925,In_857);
nor U3732 (N_3732,In_286,In_292);
nor U3733 (N_3733,In_474,In_304);
and U3734 (N_3734,In_78,In_885);
xnor U3735 (N_3735,In_300,In_291);
nor U3736 (N_3736,In_360,In_477);
nor U3737 (N_3737,In_398,In_900);
nand U3738 (N_3738,In_497,In_456);
and U3739 (N_3739,In_433,In_801);
nor U3740 (N_3740,In_614,In_368);
nand U3741 (N_3741,In_986,In_345);
nand U3742 (N_3742,In_15,In_432);
or U3743 (N_3743,In_136,In_813);
nand U3744 (N_3744,In_309,In_885);
nand U3745 (N_3745,In_248,In_1);
nand U3746 (N_3746,In_335,In_915);
or U3747 (N_3747,In_11,In_63);
nor U3748 (N_3748,In_580,In_649);
nand U3749 (N_3749,In_968,In_567);
nand U3750 (N_3750,In_386,In_506);
or U3751 (N_3751,In_286,In_144);
nor U3752 (N_3752,In_878,In_321);
or U3753 (N_3753,In_502,In_838);
or U3754 (N_3754,In_776,In_682);
and U3755 (N_3755,In_6,In_855);
nor U3756 (N_3756,In_644,In_660);
and U3757 (N_3757,In_914,In_205);
and U3758 (N_3758,In_417,In_840);
and U3759 (N_3759,In_41,In_349);
and U3760 (N_3760,In_205,In_285);
nor U3761 (N_3761,In_855,In_203);
nand U3762 (N_3762,In_454,In_23);
and U3763 (N_3763,In_118,In_552);
nor U3764 (N_3764,In_40,In_98);
or U3765 (N_3765,In_221,In_706);
nand U3766 (N_3766,In_726,In_677);
nor U3767 (N_3767,In_299,In_623);
or U3768 (N_3768,In_258,In_486);
or U3769 (N_3769,In_964,In_235);
and U3770 (N_3770,In_319,In_205);
or U3771 (N_3771,In_879,In_313);
or U3772 (N_3772,In_529,In_95);
nand U3773 (N_3773,In_57,In_554);
or U3774 (N_3774,In_750,In_749);
xor U3775 (N_3775,In_660,In_575);
or U3776 (N_3776,In_449,In_640);
nor U3777 (N_3777,In_854,In_199);
and U3778 (N_3778,In_326,In_624);
nor U3779 (N_3779,In_658,In_193);
nor U3780 (N_3780,In_372,In_84);
and U3781 (N_3781,In_487,In_283);
nor U3782 (N_3782,In_534,In_638);
and U3783 (N_3783,In_531,In_556);
and U3784 (N_3784,In_243,In_227);
nand U3785 (N_3785,In_716,In_2);
nor U3786 (N_3786,In_858,In_699);
nand U3787 (N_3787,In_946,In_478);
nor U3788 (N_3788,In_197,In_972);
and U3789 (N_3789,In_267,In_228);
nand U3790 (N_3790,In_229,In_394);
nor U3791 (N_3791,In_794,In_746);
nor U3792 (N_3792,In_752,In_242);
and U3793 (N_3793,In_617,In_981);
and U3794 (N_3794,In_561,In_822);
nor U3795 (N_3795,In_260,In_870);
xor U3796 (N_3796,In_116,In_381);
nor U3797 (N_3797,In_537,In_869);
xor U3798 (N_3798,In_568,In_242);
nor U3799 (N_3799,In_777,In_136);
nor U3800 (N_3800,In_575,In_701);
or U3801 (N_3801,In_834,In_830);
nand U3802 (N_3802,In_908,In_889);
nor U3803 (N_3803,In_469,In_636);
or U3804 (N_3804,In_865,In_994);
nor U3805 (N_3805,In_620,In_4);
nand U3806 (N_3806,In_489,In_465);
nor U3807 (N_3807,In_128,In_279);
nand U3808 (N_3808,In_229,In_100);
or U3809 (N_3809,In_212,In_371);
nand U3810 (N_3810,In_156,In_646);
or U3811 (N_3811,In_731,In_481);
and U3812 (N_3812,In_840,In_983);
nand U3813 (N_3813,In_928,In_390);
nor U3814 (N_3814,In_586,In_882);
or U3815 (N_3815,In_174,In_353);
and U3816 (N_3816,In_606,In_492);
xnor U3817 (N_3817,In_633,In_160);
and U3818 (N_3818,In_493,In_717);
and U3819 (N_3819,In_195,In_165);
or U3820 (N_3820,In_349,In_821);
nand U3821 (N_3821,In_412,In_969);
or U3822 (N_3822,In_348,In_723);
and U3823 (N_3823,In_91,In_723);
and U3824 (N_3824,In_593,In_290);
nand U3825 (N_3825,In_221,In_925);
nand U3826 (N_3826,In_326,In_823);
nor U3827 (N_3827,In_789,In_649);
and U3828 (N_3828,In_277,In_750);
nand U3829 (N_3829,In_905,In_89);
or U3830 (N_3830,In_978,In_160);
or U3831 (N_3831,In_338,In_748);
and U3832 (N_3832,In_789,In_804);
or U3833 (N_3833,In_709,In_684);
and U3834 (N_3834,In_779,In_166);
and U3835 (N_3835,In_346,In_140);
and U3836 (N_3836,In_780,In_757);
nor U3837 (N_3837,In_579,In_435);
nor U3838 (N_3838,In_427,In_680);
and U3839 (N_3839,In_111,In_323);
nand U3840 (N_3840,In_538,In_479);
nand U3841 (N_3841,In_161,In_424);
nand U3842 (N_3842,In_409,In_853);
xnor U3843 (N_3843,In_715,In_236);
or U3844 (N_3844,In_945,In_239);
and U3845 (N_3845,In_267,In_275);
nand U3846 (N_3846,In_310,In_786);
nand U3847 (N_3847,In_717,In_704);
or U3848 (N_3848,In_495,In_161);
and U3849 (N_3849,In_677,In_641);
and U3850 (N_3850,In_116,In_554);
and U3851 (N_3851,In_266,In_26);
nand U3852 (N_3852,In_654,In_901);
or U3853 (N_3853,In_543,In_817);
nand U3854 (N_3854,In_674,In_837);
xor U3855 (N_3855,In_73,In_780);
nand U3856 (N_3856,In_504,In_401);
nor U3857 (N_3857,In_258,In_747);
and U3858 (N_3858,In_944,In_866);
and U3859 (N_3859,In_686,In_86);
nand U3860 (N_3860,In_241,In_147);
and U3861 (N_3861,In_516,In_699);
and U3862 (N_3862,In_946,In_369);
nor U3863 (N_3863,In_592,In_786);
nand U3864 (N_3864,In_0,In_308);
nor U3865 (N_3865,In_898,In_742);
nand U3866 (N_3866,In_158,In_414);
nor U3867 (N_3867,In_280,In_495);
nand U3868 (N_3868,In_139,In_914);
or U3869 (N_3869,In_370,In_432);
nor U3870 (N_3870,In_292,In_562);
or U3871 (N_3871,In_597,In_280);
and U3872 (N_3872,In_256,In_507);
and U3873 (N_3873,In_372,In_629);
xor U3874 (N_3874,In_97,In_517);
and U3875 (N_3875,In_235,In_461);
nor U3876 (N_3876,In_205,In_708);
and U3877 (N_3877,In_428,In_704);
or U3878 (N_3878,In_282,In_319);
nand U3879 (N_3879,In_206,In_203);
nor U3880 (N_3880,In_44,In_796);
nand U3881 (N_3881,In_200,In_99);
or U3882 (N_3882,In_190,In_946);
or U3883 (N_3883,In_907,In_375);
or U3884 (N_3884,In_716,In_778);
nor U3885 (N_3885,In_983,In_23);
and U3886 (N_3886,In_1,In_899);
and U3887 (N_3887,In_725,In_412);
and U3888 (N_3888,In_294,In_172);
or U3889 (N_3889,In_945,In_928);
or U3890 (N_3890,In_40,In_120);
xnor U3891 (N_3891,In_90,In_841);
nor U3892 (N_3892,In_830,In_448);
or U3893 (N_3893,In_453,In_661);
xor U3894 (N_3894,In_298,In_594);
and U3895 (N_3895,In_284,In_632);
nand U3896 (N_3896,In_225,In_671);
or U3897 (N_3897,In_511,In_931);
nand U3898 (N_3898,In_401,In_961);
or U3899 (N_3899,In_846,In_545);
or U3900 (N_3900,In_203,In_221);
nand U3901 (N_3901,In_843,In_284);
nor U3902 (N_3902,In_388,In_401);
nand U3903 (N_3903,In_235,In_441);
nor U3904 (N_3904,In_496,In_947);
and U3905 (N_3905,In_725,In_231);
or U3906 (N_3906,In_770,In_610);
and U3907 (N_3907,In_970,In_551);
and U3908 (N_3908,In_847,In_268);
nor U3909 (N_3909,In_562,In_617);
nor U3910 (N_3910,In_380,In_787);
nor U3911 (N_3911,In_334,In_67);
nand U3912 (N_3912,In_163,In_850);
nand U3913 (N_3913,In_500,In_212);
or U3914 (N_3914,In_676,In_210);
or U3915 (N_3915,In_755,In_461);
nand U3916 (N_3916,In_407,In_251);
and U3917 (N_3917,In_225,In_436);
nor U3918 (N_3918,In_250,In_84);
or U3919 (N_3919,In_344,In_882);
and U3920 (N_3920,In_905,In_151);
or U3921 (N_3921,In_496,In_285);
and U3922 (N_3922,In_887,In_218);
nand U3923 (N_3923,In_677,In_667);
nand U3924 (N_3924,In_730,In_258);
nand U3925 (N_3925,In_823,In_67);
and U3926 (N_3926,In_193,In_506);
and U3927 (N_3927,In_185,In_483);
or U3928 (N_3928,In_338,In_340);
or U3929 (N_3929,In_532,In_122);
or U3930 (N_3930,In_439,In_490);
nand U3931 (N_3931,In_275,In_738);
nor U3932 (N_3932,In_876,In_213);
nor U3933 (N_3933,In_795,In_936);
and U3934 (N_3934,In_697,In_200);
nand U3935 (N_3935,In_856,In_920);
or U3936 (N_3936,In_183,In_733);
and U3937 (N_3937,In_29,In_891);
nor U3938 (N_3938,In_573,In_132);
xor U3939 (N_3939,In_461,In_307);
nand U3940 (N_3940,In_996,In_490);
nand U3941 (N_3941,In_70,In_502);
or U3942 (N_3942,In_134,In_121);
nor U3943 (N_3943,In_791,In_362);
and U3944 (N_3944,In_540,In_922);
and U3945 (N_3945,In_642,In_625);
and U3946 (N_3946,In_533,In_908);
nand U3947 (N_3947,In_426,In_526);
and U3948 (N_3948,In_48,In_333);
and U3949 (N_3949,In_795,In_71);
nand U3950 (N_3950,In_385,In_498);
or U3951 (N_3951,In_69,In_717);
nand U3952 (N_3952,In_915,In_967);
nor U3953 (N_3953,In_839,In_78);
and U3954 (N_3954,In_354,In_630);
and U3955 (N_3955,In_987,In_666);
nand U3956 (N_3956,In_892,In_271);
nand U3957 (N_3957,In_778,In_450);
nor U3958 (N_3958,In_325,In_500);
nand U3959 (N_3959,In_621,In_194);
or U3960 (N_3960,In_243,In_639);
nor U3961 (N_3961,In_685,In_298);
nor U3962 (N_3962,In_377,In_529);
or U3963 (N_3963,In_560,In_810);
or U3964 (N_3964,In_785,In_107);
nor U3965 (N_3965,In_847,In_503);
nand U3966 (N_3966,In_853,In_892);
or U3967 (N_3967,In_842,In_459);
and U3968 (N_3968,In_915,In_845);
or U3969 (N_3969,In_332,In_87);
nor U3970 (N_3970,In_144,In_53);
nor U3971 (N_3971,In_362,In_471);
nand U3972 (N_3972,In_792,In_879);
or U3973 (N_3973,In_271,In_362);
or U3974 (N_3974,In_972,In_976);
nor U3975 (N_3975,In_636,In_617);
nor U3976 (N_3976,In_894,In_550);
and U3977 (N_3977,In_584,In_116);
nor U3978 (N_3978,In_913,In_447);
or U3979 (N_3979,In_197,In_27);
or U3980 (N_3980,In_356,In_503);
or U3981 (N_3981,In_146,In_765);
and U3982 (N_3982,In_209,In_591);
and U3983 (N_3983,In_971,In_275);
nand U3984 (N_3984,In_780,In_101);
xor U3985 (N_3985,In_648,In_678);
or U3986 (N_3986,In_357,In_920);
nand U3987 (N_3987,In_73,In_708);
or U3988 (N_3988,In_586,In_334);
or U3989 (N_3989,In_900,In_636);
nor U3990 (N_3990,In_821,In_438);
nand U3991 (N_3991,In_105,In_207);
or U3992 (N_3992,In_248,In_520);
nand U3993 (N_3993,In_827,In_512);
or U3994 (N_3994,In_200,In_117);
nand U3995 (N_3995,In_722,In_282);
and U3996 (N_3996,In_457,In_23);
nand U3997 (N_3997,In_10,In_194);
nor U3998 (N_3998,In_868,In_154);
or U3999 (N_3999,In_233,In_639);
and U4000 (N_4000,In_650,In_102);
nand U4001 (N_4001,In_459,In_294);
nand U4002 (N_4002,In_586,In_203);
nand U4003 (N_4003,In_259,In_42);
nor U4004 (N_4004,In_887,In_28);
or U4005 (N_4005,In_425,In_531);
nor U4006 (N_4006,In_165,In_89);
nand U4007 (N_4007,In_778,In_215);
xor U4008 (N_4008,In_877,In_176);
nand U4009 (N_4009,In_946,In_651);
or U4010 (N_4010,In_797,In_315);
nor U4011 (N_4011,In_526,In_953);
and U4012 (N_4012,In_478,In_244);
and U4013 (N_4013,In_18,In_193);
xor U4014 (N_4014,In_465,In_124);
nand U4015 (N_4015,In_249,In_996);
nand U4016 (N_4016,In_597,In_2);
or U4017 (N_4017,In_671,In_545);
or U4018 (N_4018,In_316,In_49);
and U4019 (N_4019,In_699,In_754);
and U4020 (N_4020,In_68,In_16);
or U4021 (N_4021,In_369,In_569);
or U4022 (N_4022,In_515,In_14);
or U4023 (N_4023,In_905,In_357);
nor U4024 (N_4024,In_214,In_554);
nand U4025 (N_4025,In_409,In_202);
nor U4026 (N_4026,In_517,In_447);
and U4027 (N_4027,In_628,In_849);
and U4028 (N_4028,In_867,In_21);
nand U4029 (N_4029,In_72,In_347);
xor U4030 (N_4030,In_791,In_295);
or U4031 (N_4031,In_116,In_396);
or U4032 (N_4032,In_168,In_582);
nor U4033 (N_4033,In_62,In_910);
nor U4034 (N_4034,In_843,In_868);
or U4035 (N_4035,In_43,In_934);
nor U4036 (N_4036,In_321,In_397);
nor U4037 (N_4037,In_431,In_818);
and U4038 (N_4038,In_658,In_825);
and U4039 (N_4039,In_503,In_322);
and U4040 (N_4040,In_151,In_519);
nor U4041 (N_4041,In_610,In_833);
nand U4042 (N_4042,In_219,In_119);
and U4043 (N_4043,In_123,In_383);
or U4044 (N_4044,In_539,In_211);
nand U4045 (N_4045,In_632,In_20);
nor U4046 (N_4046,In_918,In_240);
and U4047 (N_4047,In_931,In_229);
nand U4048 (N_4048,In_370,In_866);
nand U4049 (N_4049,In_984,In_933);
nand U4050 (N_4050,In_108,In_461);
nand U4051 (N_4051,In_877,In_183);
and U4052 (N_4052,In_465,In_137);
or U4053 (N_4053,In_985,In_720);
nor U4054 (N_4054,In_127,In_994);
or U4055 (N_4055,In_390,In_155);
and U4056 (N_4056,In_582,In_73);
nor U4057 (N_4057,In_141,In_878);
nand U4058 (N_4058,In_444,In_840);
and U4059 (N_4059,In_347,In_753);
or U4060 (N_4060,In_423,In_974);
nand U4061 (N_4061,In_206,In_744);
nor U4062 (N_4062,In_137,In_604);
nor U4063 (N_4063,In_643,In_111);
or U4064 (N_4064,In_500,In_919);
and U4065 (N_4065,In_177,In_988);
or U4066 (N_4066,In_387,In_554);
and U4067 (N_4067,In_152,In_667);
nand U4068 (N_4068,In_330,In_417);
or U4069 (N_4069,In_780,In_580);
nor U4070 (N_4070,In_526,In_211);
or U4071 (N_4071,In_422,In_11);
nor U4072 (N_4072,In_109,In_170);
and U4073 (N_4073,In_31,In_243);
or U4074 (N_4074,In_819,In_132);
or U4075 (N_4075,In_46,In_201);
nor U4076 (N_4076,In_791,In_461);
or U4077 (N_4077,In_562,In_566);
or U4078 (N_4078,In_539,In_448);
and U4079 (N_4079,In_43,In_402);
nor U4080 (N_4080,In_754,In_43);
nand U4081 (N_4081,In_881,In_723);
or U4082 (N_4082,In_458,In_844);
nor U4083 (N_4083,In_230,In_425);
nor U4084 (N_4084,In_156,In_262);
and U4085 (N_4085,In_179,In_770);
or U4086 (N_4086,In_69,In_651);
and U4087 (N_4087,In_608,In_361);
nand U4088 (N_4088,In_710,In_486);
and U4089 (N_4089,In_117,In_591);
or U4090 (N_4090,In_758,In_668);
nand U4091 (N_4091,In_181,In_99);
nand U4092 (N_4092,In_7,In_823);
nor U4093 (N_4093,In_759,In_550);
or U4094 (N_4094,In_361,In_940);
nor U4095 (N_4095,In_674,In_130);
and U4096 (N_4096,In_646,In_185);
or U4097 (N_4097,In_225,In_109);
nand U4098 (N_4098,In_574,In_396);
and U4099 (N_4099,In_383,In_228);
nor U4100 (N_4100,In_180,In_777);
nand U4101 (N_4101,In_706,In_725);
and U4102 (N_4102,In_101,In_382);
nor U4103 (N_4103,In_601,In_255);
nand U4104 (N_4104,In_406,In_614);
or U4105 (N_4105,In_477,In_274);
or U4106 (N_4106,In_652,In_24);
or U4107 (N_4107,In_551,In_144);
and U4108 (N_4108,In_230,In_650);
nand U4109 (N_4109,In_293,In_848);
or U4110 (N_4110,In_516,In_179);
or U4111 (N_4111,In_670,In_584);
or U4112 (N_4112,In_857,In_537);
nor U4113 (N_4113,In_466,In_417);
or U4114 (N_4114,In_304,In_315);
nand U4115 (N_4115,In_2,In_111);
nor U4116 (N_4116,In_368,In_60);
or U4117 (N_4117,In_181,In_849);
nand U4118 (N_4118,In_185,In_301);
and U4119 (N_4119,In_636,In_216);
or U4120 (N_4120,In_39,In_547);
nand U4121 (N_4121,In_207,In_815);
or U4122 (N_4122,In_566,In_161);
nor U4123 (N_4123,In_48,In_96);
or U4124 (N_4124,In_242,In_920);
nand U4125 (N_4125,In_544,In_200);
nand U4126 (N_4126,In_960,In_723);
nor U4127 (N_4127,In_932,In_269);
nand U4128 (N_4128,In_443,In_858);
and U4129 (N_4129,In_796,In_625);
or U4130 (N_4130,In_31,In_36);
or U4131 (N_4131,In_693,In_332);
nor U4132 (N_4132,In_851,In_662);
nand U4133 (N_4133,In_753,In_467);
and U4134 (N_4134,In_730,In_783);
and U4135 (N_4135,In_661,In_232);
nand U4136 (N_4136,In_394,In_231);
nand U4137 (N_4137,In_43,In_720);
nand U4138 (N_4138,In_95,In_960);
nand U4139 (N_4139,In_512,In_96);
and U4140 (N_4140,In_584,In_857);
or U4141 (N_4141,In_973,In_387);
xor U4142 (N_4142,In_909,In_981);
or U4143 (N_4143,In_592,In_29);
and U4144 (N_4144,In_376,In_576);
nand U4145 (N_4145,In_793,In_251);
nor U4146 (N_4146,In_222,In_259);
or U4147 (N_4147,In_202,In_714);
nand U4148 (N_4148,In_986,In_320);
nand U4149 (N_4149,In_371,In_892);
and U4150 (N_4150,In_556,In_724);
nor U4151 (N_4151,In_972,In_304);
or U4152 (N_4152,In_187,In_445);
and U4153 (N_4153,In_252,In_58);
and U4154 (N_4154,In_61,In_139);
nor U4155 (N_4155,In_685,In_177);
and U4156 (N_4156,In_241,In_949);
nand U4157 (N_4157,In_206,In_40);
nand U4158 (N_4158,In_46,In_283);
nand U4159 (N_4159,In_370,In_522);
and U4160 (N_4160,In_674,In_604);
or U4161 (N_4161,In_365,In_163);
nand U4162 (N_4162,In_277,In_964);
nor U4163 (N_4163,In_784,In_173);
nor U4164 (N_4164,In_996,In_186);
nand U4165 (N_4165,In_182,In_570);
nand U4166 (N_4166,In_786,In_45);
or U4167 (N_4167,In_931,In_944);
and U4168 (N_4168,In_558,In_998);
nor U4169 (N_4169,In_660,In_110);
nand U4170 (N_4170,In_998,In_577);
nand U4171 (N_4171,In_42,In_161);
and U4172 (N_4172,In_384,In_954);
or U4173 (N_4173,In_398,In_922);
and U4174 (N_4174,In_378,In_895);
nor U4175 (N_4175,In_180,In_143);
and U4176 (N_4176,In_390,In_242);
nand U4177 (N_4177,In_209,In_320);
nor U4178 (N_4178,In_512,In_626);
or U4179 (N_4179,In_299,In_52);
nor U4180 (N_4180,In_928,In_667);
and U4181 (N_4181,In_563,In_452);
xor U4182 (N_4182,In_762,In_150);
nor U4183 (N_4183,In_745,In_462);
nand U4184 (N_4184,In_593,In_941);
nand U4185 (N_4185,In_244,In_770);
nand U4186 (N_4186,In_168,In_794);
xnor U4187 (N_4187,In_444,In_44);
nand U4188 (N_4188,In_533,In_608);
nand U4189 (N_4189,In_329,In_73);
and U4190 (N_4190,In_450,In_378);
nand U4191 (N_4191,In_288,In_753);
nand U4192 (N_4192,In_382,In_832);
or U4193 (N_4193,In_476,In_417);
nor U4194 (N_4194,In_74,In_964);
nor U4195 (N_4195,In_670,In_223);
or U4196 (N_4196,In_417,In_155);
and U4197 (N_4197,In_414,In_658);
nor U4198 (N_4198,In_325,In_57);
or U4199 (N_4199,In_138,In_437);
or U4200 (N_4200,In_943,In_184);
and U4201 (N_4201,In_550,In_66);
and U4202 (N_4202,In_953,In_183);
and U4203 (N_4203,In_594,In_328);
or U4204 (N_4204,In_702,In_448);
or U4205 (N_4205,In_889,In_937);
and U4206 (N_4206,In_987,In_812);
nor U4207 (N_4207,In_463,In_174);
and U4208 (N_4208,In_211,In_859);
nand U4209 (N_4209,In_861,In_591);
nor U4210 (N_4210,In_115,In_482);
nor U4211 (N_4211,In_387,In_916);
xor U4212 (N_4212,In_848,In_0);
or U4213 (N_4213,In_246,In_559);
nor U4214 (N_4214,In_575,In_180);
nor U4215 (N_4215,In_136,In_489);
or U4216 (N_4216,In_616,In_364);
or U4217 (N_4217,In_513,In_564);
nor U4218 (N_4218,In_181,In_124);
nand U4219 (N_4219,In_591,In_826);
nor U4220 (N_4220,In_832,In_869);
and U4221 (N_4221,In_292,In_629);
nor U4222 (N_4222,In_159,In_142);
xor U4223 (N_4223,In_334,In_637);
and U4224 (N_4224,In_355,In_634);
and U4225 (N_4225,In_306,In_943);
and U4226 (N_4226,In_817,In_957);
or U4227 (N_4227,In_722,In_706);
nor U4228 (N_4228,In_866,In_946);
nor U4229 (N_4229,In_359,In_570);
and U4230 (N_4230,In_144,In_270);
or U4231 (N_4231,In_193,In_650);
and U4232 (N_4232,In_13,In_396);
nand U4233 (N_4233,In_937,In_637);
nor U4234 (N_4234,In_572,In_500);
nor U4235 (N_4235,In_932,In_503);
and U4236 (N_4236,In_11,In_647);
and U4237 (N_4237,In_656,In_219);
nor U4238 (N_4238,In_123,In_458);
nand U4239 (N_4239,In_81,In_687);
or U4240 (N_4240,In_871,In_697);
nand U4241 (N_4241,In_362,In_44);
nand U4242 (N_4242,In_76,In_792);
xor U4243 (N_4243,In_661,In_408);
nor U4244 (N_4244,In_175,In_715);
xnor U4245 (N_4245,In_948,In_547);
or U4246 (N_4246,In_330,In_324);
nand U4247 (N_4247,In_953,In_374);
nor U4248 (N_4248,In_464,In_179);
nor U4249 (N_4249,In_754,In_546);
and U4250 (N_4250,In_365,In_275);
nor U4251 (N_4251,In_571,In_713);
nor U4252 (N_4252,In_495,In_975);
or U4253 (N_4253,In_341,In_984);
nand U4254 (N_4254,In_731,In_119);
nor U4255 (N_4255,In_248,In_688);
nand U4256 (N_4256,In_908,In_770);
xnor U4257 (N_4257,In_63,In_890);
and U4258 (N_4258,In_444,In_569);
and U4259 (N_4259,In_103,In_270);
or U4260 (N_4260,In_536,In_610);
nor U4261 (N_4261,In_576,In_837);
nor U4262 (N_4262,In_753,In_787);
and U4263 (N_4263,In_329,In_777);
and U4264 (N_4264,In_295,In_371);
or U4265 (N_4265,In_910,In_501);
nand U4266 (N_4266,In_335,In_153);
nor U4267 (N_4267,In_598,In_805);
nand U4268 (N_4268,In_116,In_17);
xor U4269 (N_4269,In_958,In_199);
nor U4270 (N_4270,In_336,In_232);
or U4271 (N_4271,In_731,In_983);
or U4272 (N_4272,In_93,In_513);
or U4273 (N_4273,In_752,In_44);
nand U4274 (N_4274,In_190,In_343);
nand U4275 (N_4275,In_116,In_178);
nor U4276 (N_4276,In_658,In_710);
nor U4277 (N_4277,In_207,In_258);
and U4278 (N_4278,In_377,In_502);
nand U4279 (N_4279,In_304,In_413);
nor U4280 (N_4280,In_98,In_515);
and U4281 (N_4281,In_590,In_879);
or U4282 (N_4282,In_349,In_701);
or U4283 (N_4283,In_212,In_787);
nand U4284 (N_4284,In_123,In_687);
nor U4285 (N_4285,In_299,In_230);
nand U4286 (N_4286,In_178,In_958);
nand U4287 (N_4287,In_65,In_795);
nor U4288 (N_4288,In_721,In_430);
or U4289 (N_4289,In_910,In_714);
and U4290 (N_4290,In_759,In_234);
and U4291 (N_4291,In_713,In_860);
or U4292 (N_4292,In_207,In_873);
and U4293 (N_4293,In_279,In_105);
nand U4294 (N_4294,In_612,In_171);
nor U4295 (N_4295,In_218,In_657);
nor U4296 (N_4296,In_178,In_208);
nor U4297 (N_4297,In_489,In_892);
and U4298 (N_4298,In_633,In_13);
and U4299 (N_4299,In_895,In_439);
nand U4300 (N_4300,In_150,In_858);
or U4301 (N_4301,In_56,In_646);
and U4302 (N_4302,In_71,In_872);
and U4303 (N_4303,In_669,In_467);
nor U4304 (N_4304,In_181,In_885);
and U4305 (N_4305,In_799,In_859);
or U4306 (N_4306,In_316,In_621);
and U4307 (N_4307,In_665,In_775);
and U4308 (N_4308,In_877,In_587);
and U4309 (N_4309,In_843,In_897);
nand U4310 (N_4310,In_96,In_773);
and U4311 (N_4311,In_69,In_138);
nor U4312 (N_4312,In_321,In_478);
nor U4313 (N_4313,In_805,In_206);
nand U4314 (N_4314,In_170,In_877);
or U4315 (N_4315,In_428,In_690);
or U4316 (N_4316,In_551,In_176);
nand U4317 (N_4317,In_16,In_321);
nand U4318 (N_4318,In_330,In_744);
or U4319 (N_4319,In_249,In_50);
or U4320 (N_4320,In_361,In_916);
and U4321 (N_4321,In_680,In_960);
nor U4322 (N_4322,In_597,In_167);
or U4323 (N_4323,In_985,In_462);
nand U4324 (N_4324,In_189,In_45);
nor U4325 (N_4325,In_407,In_706);
nand U4326 (N_4326,In_96,In_38);
nor U4327 (N_4327,In_694,In_585);
nor U4328 (N_4328,In_163,In_489);
nand U4329 (N_4329,In_537,In_231);
and U4330 (N_4330,In_553,In_300);
nand U4331 (N_4331,In_998,In_832);
or U4332 (N_4332,In_683,In_794);
nand U4333 (N_4333,In_179,In_919);
or U4334 (N_4334,In_947,In_657);
and U4335 (N_4335,In_188,In_196);
and U4336 (N_4336,In_674,In_750);
nand U4337 (N_4337,In_729,In_116);
or U4338 (N_4338,In_370,In_386);
nand U4339 (N_4339,In_64,In_683);
nand U4340 (N_4340,In_606,In_21);
nand U4341 (N_4341,In_996,In_193);
or U4342 (N_4342,In_997,In_177);
nand U4343 (N_4343,In_373,In_895);
nor U4344 (N_4344,In_928,In_466);
nand U4345 (N_4345,In_552,In_789);
xnor U4346 (N_4346,In_327,In_410);
nand U4347 (N_4347,In_821,In_371);
nor U4348 (N_4348,In_752,In_963);
and U4349 (N_4349,In_217,In_398);
xor U4350 (N_4350,In_136,In_418);
and U4351 (N_4351,In_410,In_435);
or U4352 (N_4352,In_359,In_161);
or U4353 (N_4353,In_831,In_285);
and U4354 (N_4354,In_633,In_278);
or U4355 (N_4355,In_697,In_887);
xnor U4356 (N_4356,In_924,In_844);
nor U4357 (N_4357,In_478,In_618);
nor U4358 (N_4358,In_261,In_973);
nand U4359 (N_4359,In_71,In_915);
nand U4360 (N_4360,In_767,In_540);
nand U4361 (N_4361,In_579,In_137);
nor U4362 (N_4362,In_379,In_757);
nor U4363 (N_4363,In_95,In_67);
nand U4364 (N_4364,In_520,In_900);
nand U4365 (N_4365,In_916,In_305);
nor U4366 (N_4366,In_706,In_95);
or U4367 (N_4367,In_661,In_998);
nand U4368 (N_4368,In_311,In_286);
nor U4369 (N_4369,In_991,In_731);
nand U4370 (N_4370,In_860,In_132);
nand U4371 (N_4371,In_58,In_165);
nor U4372 (N_4372,In_619,In_809);
nor U4373 (N_4373,In_117,In_555);
nand U4374 (N_4374,In_751,In_861);
nor U4375 (N_4375,In_326,In_581);
and U4376 (N_4376,In_711,In_979);
nor U4377 (N_4377,In_918,In_29);
or U4378 (N_4378,In_604,In_285);
nor U4379 (N_4379,In_671,In_737);
nand U4380 (N_4380,In_402,In_530);
nor U4381 (N_4381,In_255,In_199);
nand U4382 (N_4382,In_838,In_818);
nand U4383 (N_4383,In_351,In_994);
or U4384 (N_4384,In_747,In_248);
or U4385 (N_4385,In_947,In_62);
nand U4386 (N_4386,In_862,In_472);
nor U4387 (N_4387,In_866,In_844);
or U4388 (N_4388,In_497,In_863);
or U4389 (N_4389,In_124,In_610);
or U4390 (N_4390,In_212,In_505);
nor U4391 (N_4391,In_235,In_712);
nand U4392 (N_4392,In_716,In_735);
nor U4393 (N_4393,In_250,In_72);
nor U4394 (N_4394,In_172,In_566);
nand U4395 (N_4395,In_662,In_936);
nor U4396 (N_4396,In_429,In_641);
or U4397 (N_4397,In_919,In_67);
nand U4398 (N_4398,In_925,In_269);
nand U4399 (N_4399,In_528,In_259);
or U4400 (N_4400,In_656,In_425);
nand U4401 (N_4401,In_202,In_504);
and U4402 (N_4402,In_416,In_301);
nand U4403 (N_4403,In_716,In_411);
nand U4404 (N_4404,In_422,In_989);
and U4405 (N_4405,In_913,In_7);
and U4406 (N_4406,In_15,In_928);
or U4407 (N_4407,In_281,In_390);
nand U4408 (N_4408,In_424,In_340);
nor U4409 (N_4409,In_575,In_458);
nand U4410 (N_4410,In_854,In_397);
or U4411 (N_4411,In_391,In_516);
nor U4412 (N_4412,In_225,In_309);
or U4413 (N_4413,In_842,In_711);
or U4414 (N_4414,In_110,In_583);
or U4415 (N_4415,In_914,In_500);
or U4416 (N_4416,In_328,In_606);
or U4417 (N_4417,In_651,In_297);
or U4418 (N_4418,In_723,In_374);
nand U4419 (N_4419,In_489,In_894);
nand U4420 (N_4420,In_869,In_168);
or U4421 (N_4421,In_597,In_825);
nor U4422 (N_4422,In_50,In_11);
and U4423 (N_4423,In_683,In_874);
or U4424 (N_4424,In_823,In_249);
nand U4425 (N_4425,In_933,In_127);
xor U4426 (N_4426,In_650,In_767);
nand U4427 (N_4427,In_238,In_917);
nand U4428 (N_4428,In_580,In_817);
nand U4429 (N_4429,In_271,In_894);
xor U4430 (N_4430,In_846,In_779);
and U4431 (N_4431,In_454,In_151);
nand U4432 (N_4432,In_271,In_336);
and U4433 (N_4433,In_829,In_572);
and U4434 (N_4434,In_650,In_365);
nand U4435 (N_4435,In_992,In_208);
nand U4436 (N_4436,In_336,In_365);
nor U4437 (N_4437,In_407,In_220);
nor U4438 (N_4438,In_584,In_987);
nand U4439 (N_4439,In_679,In_796);
nor U4440 (N_4440,In_753,In_657);
nor U4441 (N_4441,In_806,In_970);
xnor U4442 (N_4442,In_641,In_824);
nor U4443 (N_4443,In_641,In_925);
nand U4444 (N_4444,In_17,In_795);
xor U4445 (N_4445,In_808,In_698);
nand U4446 (N_4446,In_862,In_35);
or U4447 (N_4447,In_343,In_668);
or U4448 (N_4448,In_533,In_783);
and U4449 (N_4449,In_913,In_992);
nand U4450 (N_4450,In_392,In_200);
xor U4451 (N_4451,In_929,In_404);
nand U4452 (N_4452,In_315,In_21);
nand U4453 (N_4453,In_770,In_786);
nor U4454 (N_4454,In_919,In_613);
and U4455 (N_4455,In_490,In_75);
nand U4456 (N_4456,In_378,In_926);
and U4457 (N_4457,In_14,In_414);
nand U4458 (N_4458,In_976,In_502);
nor U4459 (N_4459,In_182,In_272);
nand U4460 (N_4460,In_885,In_16);
nand U4461 (N_4461,In_371,In_592);
nand U4462 (N_4462,In_143,In_793);
or U4463 (N_4463,In_394,In_424);
nand U4464 (N_4464,In_159,In_580);
and U4465 (N_4465,In_582,In_756);
nand U4466 (N_4466,In_748,In_303);
and U4467 (N_4467,In_797,In_242);
or U4468 (N_4468,In_273,In_986);
nor U4469 (N_4469,In_786,In_933);
and U4470 (N_4470,In_282,In_887);
nand U4471 (N_4471,In_125,In_534);
nor U4472 (N_4472,In_536,In_705);
or U4473 (N_4473,In_675,In_745);
nand U4474 (N_4474,In_572,In_796);
or U4475 (N_4475,In_164,In_387);
nand U4476 (N_4476,In_173,In_512);
nor U4477 (N_4477,In_222,In_805);
and U4478 (N_4478,In_515,In_921);
nand U4479 (N_4479,In_675,In_394);
nor U4480 (N_4480,In_537,In_560);
nand U4481 (N_4481,In_888,In_134);
or U4482 (N_4482,In_349,In_63);
or U4483 (N_4483,In_285,In_138);
or U4484 (N_4484,In_631,In_909);
or U4485 (N_4485,In_642,In_118);
nor U4486 (N_4486,In_633,In_755);
nor U4487 (N_4487,In_494,In_592);
nor U4488 (N_4488,In_759,In_539);
nand U4489 (N_4489,In_349,In_424);
and U4490 (N_4490,In_61,In_726);
nor U4491 (N_4491,In_850,In_312);
nor U4492 (N_4492,In_505,In_869);
and U4493 (N_4493,In_932,In_307);
or U4494 (N_4494,In_158,In_7);
and U4495 (N_4495,In_305,In_39);
and U4496 (N_4496,In_144,In_627);
xor U4497 (N_4497,In_11,In_879);
nor U4498 (N_4498,In_285,In_317);
or U4499 (N_4499,In_210,In_181);
nand U4500 (N_4500,In_88,In_825);
nand U4501 (N_4501,In_234,In_318);
nand U4502 (N_4502,In_444,In_283);
or U4503 (N_4503,In_153,In_851);
nor U4504 (N_4504,In_837,In_247);
and U4505 (N_4505,In_421,In_961);
nand U4506 (N_4506,In_729,In_554);
nor U4507 (N_4507,In_734,In_558);
or U4508 (N_4508,In_980,In_103);
or U4509 (N_4509,In_659,In_884);
nand U4510 (N_4510,In_861,In_196);
nor U4511 (N_4511,In_457,In_756);
nand U4512 (N_4512,In_54,In_956);
nor U4513 (N_4513,In_872,In_799);
or U4514 (N_4514,In_928,In_109);
and U4515 (N_4515,In_367,In_730);
nor U4516 (N_4516,In_917,In_196);
and U4517 (N_4517,In_483,In_45);
nor U4518 (N_4518,In_453,In_540);
and U4519 (N_4519,In_120,In_253);
nor U4520 (N_4520,In_570,In_729);
nand U4521 (N_4521,In_436,In_47);
nor U4522 (N_4522,In_462,In_987);
or U4523 (N_4523,In_522,In_343);
nand U4524 (N_4524,In_936,In_523);
nand U4525 (N_4525,In_3,In_928);
and U4526 (N_4526,In_546,In_651);
or U4527 (N_4527,In_981,In_267);
or U4528 (N_4528,In_922,In_255);
nor U4529 (N_4529,In_176,In_542);
or U4530 (N_4530,In_193,In_331);
nor U4531 (N_4531,In_68,In_648);
and U4532 (N_4532,In_37,In_547);
and U4533 (N_4533,In_620,In_491);
nand U4534 (N_4534,In_590,In_829);
xor U4535 (N_4535,In_578,In_741);
or U4536 (N_4536,In_362,In_687);
nor U4537 (N_4537,In_265,In_342);
nor U4538 (N_4538,In_674,In_32);
or U4539 (N_4539,In_581,In_123);
or U4540 (N_4540,In_957,In_434);
nor U4541 (N_4541,In_330,In_357);
and U4542 (N_4542,In_359,In_382);
nor U4543 (N_4543,In_556,In_270);
or U4544 (N_4544,In_155,In_151);
and U4545 (N_4545,In_555,In_389);
nor U4546 (N_4546,In_639,In_672);
nor U4547 (N_4547,In_705,In_530);
or U4548 (N_4548,In_457,In_138);
or U4549 (N_4549,In_816,In_774);
nand U4550 (N_4550,In_913,In_612);
nand U4551 (N_4551,In_927,In_199);
nand U4552 (N_4552,In_399,In_77);
nand U4553 (N_4553,In_843,In_681);
and U4554 (N_4554,In_874,In_816);
or U4555 (N_4555,In_40,In_485);
nand U4556 (N_4556,In_439,In_652);
nor U4557 (N_4557,In_45,In_911);
or U4558 (N_4558,In_555,In_741);
or U4559 (N_4559,In_55,In_681);
and U4560 (N_4560,In_145,In_768);
or U4561 (N_4561,In_713,In_31);
xor U4562 (N_4562,In_20,In_918);
nand U4563 (N_4563,In_425,In_988);
nand U4564 (N_4564,In_812,In_33);
nor U4565 (N_4565,In_133,In_624);
or U4566 (N_4566,In_420,In_444);
and U4567 (N_4567,In_353,In_677);
nand U4568 (N_4568,In_882,In_621);
or U4569 (N_4569,In_329,In_843);
and U4570 (N_4570,In_234,In_975);
nor U4571 (N_4571,In_199,In_245);
nor U4572 (N_4572,In_890,In_761);
and U4573 (N_4573,In_25,In_662);
and U4574 (N_4574,In_229,In_50);
nor U4575 (N_4575,In_612,In_370);
and U4576 (N_4576,In_371,In_666);
nand U4577 (N_4577,In_65,In_462);
or U4578 (N_4578,In_653,In_749);
or U4579 (N_4579,In_78,In_602);
or U4580 (N_4580,In_356,In_670);
or U4581 (N_4581,In_775,In_253);
or U4582 (N_4582,In_747,In_887);
or U4583 (N_4583,In_699,In_823);
nor U4584 (N_4584,In_175,In_917);
nor U4585 (N_4585,In_537,In_199);
nor U4586 (N_4586,In_646,In_545);
or U4587 (N_4587,In_503,In_713);
nor U4588 (N_4588,In_97,In_924);
nor U4589 (N_4589,In_539,In_872);
nor U4590 (N_4590,In_296,In_528);
and U4591 (N_4591,In_658,In_327);
or U4592 (N_4592,In_264,In_507);
nor U4593 (N_4593,In_670,In_94);
nand U4594 (N_4594,In_668,In_933);
or U4595 (N_4595,In_258,In_13);
and U4596 (N_4596,In_957,In_368);
nand U4597 (N_4597,In_316,In_717);
nand U4598 (N_4598,In_550,In_354);
nand U4599 (N_4599,In_974,In_716);
nand U4600 (N_4600,In_925,In_597);
nand U4601 (N_4601,In_289,In_610);
or U4602 (N_4602,In_755,In_395);
nor U4603 (N_4603,In_85,In_74);
nor U4604 (N_4604,In_50,In_242);
and U4605 (N_4605,In_648,In_417);
and U4606 (N_4606,In_617,In_800);
nor U4607 (N_4607,In_586,In_919);
or U4608 (N_4608,In_805,In_798);
or U4609 (N_4609,In_35,In_27);
and U4610 (N_4610,In_118,In_313);
and U4611 (N_4611,In_759,In_34);
nor U4612 (N_4612,In_555,In_94);
nor U4613 (N_4613,In_745,In_782);
nor U4614 (N_4614,In_868,In_560);
or U4615 (N_4615,In_957,In_650);
xor U4616 (N_4616,In_812,In_397);
or U4617 (N_4617,In_138,In_638);
and U4618 (N_4618,In_541,In_722);
nand U4619 (N_4619,In_643,In_908);
nand U4620 (N_4620,In_384,In_288);
nor U4621 (N_4621,In_576,In_457);
or U4622 (N_4622,In_526,In_896);
nor U4623 (N_4623,In_82,In_489);
or U4624 (N_4624,In_164,In_947);
nand U4625 (N_4625,In_801,In_167);
and U4626 (N_4626,In_902,In_805);
nand U4627 (N_4627,In_735,In_225);
and U4628 (N_4628,In_85,In_604);
nor U4629 (N_4629,In_760,In_722);
xor U4630 (N_4630,In_97,In_608);
nand U4631 (N_4631,In_574,In_421);
nand U4632 (N_4632,In_571,In_737);
and U4633 (N_4633,In_947,In_874);
nand U4634 (N_4634,In_196,In_435);
and U4635 (N_4635,In_183,In_436);
or U4636 (N_4636,In_961,In_283);
and U4637 (N_4637,In_38,In_25);
and U4638 (N_4638,In_257,In_278);
nor U4639 (N_4639,In_470,In_770);
nand U4640 (N_4640,In_356,In_431);
nand U4641 (N_4641,In_346,In_359);
and U4642 (N_4642,In_167,In_635);
or U4643 (N_4643,In_32,In_365);
or U4644 (N_4644,In_175,In_14);
nor U4645 (N_4645,In_541,In_36);
nand U4646 (N_4646,In_874,In_669);
or U4647 (N_4647,In_398,In_56);
nand U4648 (N_4648,In_840,In_878);
or U4649 (N_4649,In_96,In_133);
or U4650 (N_4650,In_542,In_79);
nand U4651 (N_4651,In_587,In_414);
nand U4652 (N_4652,In_620,In_167);
or U4653 (N_4653,In_699,In_525);
or U4654 (N_4654,In_643,In_152);
nor U4655 (N_4655,In_826,In_44);
nor U4656 (N_4656,In_921,In_690);
or U4657 (N_4657,In_341,In_865);
and U4658 (N_4658,In_314,In_394);
nor U4659 (N_4659,In_686,In_964);
xnor U4660 (N_4660,In_6,In_22);
nand U4661 (N_4661,In_285,In_159);
or U4662 (N_4662,In_318,In_537);
nand U4663 (N_4663,In_505,In_134);
or U4664 (N_4664,In_611,In_409);
and U4665 (N_4665,In_430,In_428);
nor U4666 (N_4666,In_325,In_749);
nand U4667 (N_4667,In_326,In_484);
nor U4668 (N_4668,In_938,In_742);
or U4669 (N_4669,In_284,In_727);
nand U4670 (N_4670,In_789,In_876);
nor U4671 (N_4671,In_424,In_280);
nor U4672 (N_4672,In_558,In_835);
or U4673 (N_4673,In_143,In_255);
or U4674 (N_4674,In_878,In_637);
nor U4675 (N_4675,In_118,In_122);
nand U4676 (N_4676,In_600,In_334);
nor U4677 (N_4677,In_737,In_416);
nor U4678 (N_4678,In_219,In_247);
nor U4679 (N_4679,In_135,In_219);
or U4680 (N_4680,In_819,In_964);
and U4681 (N_4681,In_539,In_603);
and U4682 (N_4682,In_867,In_983);
or U4683 (N_4683,In_133,In_121);
nor U4684 (N_4684,In_725,In_341);
and U4685 (N_4685,In_129,In_790);
nand U4686 (N_4686,In_175,In_844);
or U4687 (N_4687,In_552,In_222);
and U4688 (N_4688,In_249,In_190);
nand U4689 (N_4689,In_505,In_161);
nor U4690 (N_4690,In_924,In_969);
and U4691 (N_4691,In_84,In_38);
and U4692 (N_4692,In_19,In_49);
nand U4693 (N_4693,In_258,In_525);
and U4694 (N_4694,In_813,In_495);
or U4695 (N_4695,In_731,In_726);
nor U4696 (N_4696,In_931,In_578);
nand U4697 (N_4697,In_951,In_661);
nor U4698 (N_4698,In_478,In_509);
or U4699 (N_4699,In_837,In_752);
nor U4700 (N_4700,In_584,In_200);
nand U4701 (N_4701,In_53,In_431);
and U4702 (N_4702,In_273,In_378);
nor U4703 (N_4703,In_814,In_732);
nor U4704 (N_4704,In_295,In_464);
nand U4705 (N_4705,In_874,In_803);
or U4706 (N_4706,In_162,In_20);
nand U4707 (N_4707,In_215,In_310);
and U4708 (N_4708,In_181,In_56);
and U4709 (N_4709,In_936,In_759);
or U4710 (N_4710,In_222,In_533);
or U4711 (N_4711,In_381,In_773);
nand U4712 (N_4712,In_634,In_997);
or U4713 (N_4713,In_665,In_235);
and U4714 (N_4714,In_708,In_509);
nor U4715 (N_4715,In_474,In_472);
and U4716 (N_4716,In_76,In_147);
nand U4717 (N_4717,In_651,In_844);
nor U4718 (N_4718,In_265,In_354);
nor U4719 (N_4719,In_386,In_752);
nor U4720 (N_4720,In_771,In_736);
or U4721 (N_4721,In_358,In_108);
or U4722 (N_4722,In_187,In_982);
nand U4723 (N_4723,In_733,In_31);
nor U4724 (N_4724,In_837,In_811);
or U4725 (N_4725,In_968,In_640);
or U4726 (N_4726,In_64,In_170);
and U4727 (N_4727,In_723,In_315);
nor U4728 (N_4728,In_371,In_144);
nand U4729 (N_4729,In_853,In_718);
and U4730 (N_4730,In_531,In_852);
nand U4731 (N_4731,In_59,In_149);
or U4732 (N_4732,In_763,In_121);
and U4733 (N_4733,In_351,In_996);
or U4734 (N_4734,In_318,In_781);
nand U4735 (N_4735,In_884,In_104);
and U4736 (N_4736,In_250,In_355);
or U4737 (N_4737,In_194,In_584);
and U4738 (N_4738,In_853,In_458);
nor U4739 (N_4739,In_849,In_657);
or U4740 (N_4740,In_861,In_840);
or U4741 (N_4741,In_303,In_956);
nand U4742 (N_4742,In_465,In_719);
or U4743 (N_4743,In_126,In_495);
or U4744 (N_4744,In_561,In_473);
nor U4745 (N_4745,In_213,In_791);
or U4746 (N_4746,In_912,In_946);
nor U4747 (N_4747,In_256,In_451);
xnor U4748 (N_4748,In_289,In_314);
and U4749 (N_4749,In_724,In_321);
or U4750 (N_4750,In_494,In_125);
and U4751 (N_4751,In_760,In_329);
and U4752 (N_4752,In_343,In_174);
nor U4753 (N_4753,In_354,In_139);
nand U4754 (N_4754,In_273,In_177);
and U4755 (N_4755,In_852,In_445);
nor U4756 (N_4756,In_21,In_562);
and U4757 (N_4757,In_611,In_904);
and U4758 (N_4758,In_360,In_549);
nand U4759 (N_4759,In_84,In_417);
and U4760 (N_4760,In_490,In_755);
nand U4761 (N_4761,In_840,In_339);
nand U4762 (N_4762,In_590,In_923);
or U4763 (N_4763,In_483,In_205);
nor U4764 (N_4764,In_377,In_878);
nand U4765 (N_4765,In_9,In_770);
nor U4766 (N_4766,In_953,In_236);
nand U4767 (N_4767,In_793,In_601);
nor U4768 (N_4768,In_810,In_711);
or U4769 (N_4769,In_472,In_943);
and U4770 (N_4770,In_484,In_509);
or U4771 (N_4771,In_633,In_64);
nand U4772 (N_4772,In_813,In_463);
or U4773 (N_4773,In_452,In_437);
nor U4774 (N_4774,In_144,In_863);
nand U4775 (N_4775,In_185,In_284);
and U4776 (N_4776,In_731,In_673);
nand U4777 (N_4777,In_742,In_5);
nor U4778 (N_4778,In_84,In_835);
or U4779 (N_4779,In_733,In_176);
nor U4780 (N_4780,In_128,In_126);
and U4781 (N_4781,In_466,In_270);
nand U4782 (N_4782,In_999,In_852);
nand U4783 (N_4783,In_114,In_853);
and U4784 (N_4784,In_64,In_780);
or U4785 (N_4785,In_660,In_865);
and U4786 (N_4786,In_383,In_130);
nor U4787 (N_4787,In_313,In_65);
nand U4788 (N_4788,In_246,In_463);
and U4789 (N_4789,In_367,In_958);
nand U4790 (N_4790,In_519,In_200);
nor U4791 (N_4791,In_48,In_797);
or U4792 (N_4792,In_958,In_826);
or U4793 (N_4793,In_55,In_496);
and U4794 (N_4794,In_921,In_133);
or U4795 (N_4795,In_76,In_643);
nand U4796 (N_4796,In_883,In_860);
and U4797 (N_4797,In_517,In_782);
nor U4798 (N_4798,In_144,In_684);
or U4799 (N_4799,In_652,In_367);
nor U4800 (N_4800,In_85,In_909);
nand U4801 (N_4801,In_521,In_594);
nand U4802 (N_4802,In_243,In_803);
and U4803 (N_4803,In_714,In_489);
and U4804 (N_4804,In_552,In_0);
or U4805 (N_4805,In_115,In_160);
nand U4806 (N_4806,In_432,In_391);
nand U4807 (N_4807,In_343,In_585);
or U4808 (N_4808,In_645,In_330);
and U4809 (N_4809,In_683,In_722);
and U4810 (N_4810,In_889,In_708);
nor U4811 (N_4811,In_462,In_732);
nand U4812 (N_4812,In_830,In_336);
nor U4813 (N_4813,In_918,In_805);
or U4814 (N_4814,In_888,In_855);
nand U4815 (N_4815,In_828,In_762);
and U4816 (N_4816,In_207,In_843);
nand U4817 (N_4817,In_445,In_985);
nor U4818 (N_4818,In_886,In_517);
and U4819 (N_4819,In_83,In_635);
nor U4820 (N_4820,In_936,In_548);
and U4821 (N_4821,In_872,In_221);
nand U4822 (N_4822,In_370,In_73);
or U4823 (N_4823,In_436,In_198);
and U4824 (N_4824,In_353,In_550);
xnor U4825 (N_4825,In_617,In_113);
nand U4826 (N_4826,In_68,In_166);
and U4827 (N_4827,In_680,In_45);
and U4828 (N_4828,In_465,In_831);
and U4829 (N_4829,In_920,In_354);
and U4830 (N_4830,In_74,In_754);
nor U4831 (N_4831,In_338,In_294);
and U4832 (N_4832,In_120,In_367);
nor U4833 (N_4833,In_651,In_957);
or U4834 (N_4834,In_78,In_677);
nor U4835 (N_4835,In_730,In_687);
and U4836 (N_4836,In_755,In_939);
nor U4837 (N_4837,In_801,In_516);
or U4838 (N_4838,In_395,In_668);
nand U4839 (N_4839,In_638,In_456);
nand U4840 (N_4840,In_405,In_16);
or U4841 (N_4841,In_368,In_505);
nand U4842 (N_4842,In_85,In_480);
and U4843 (N_4843,In_878,In_384);
or U4844 (N_4844,In_658,In_767);
and U4845 (N_4845,In_162,In_489);
nor U4846 (N_4846,In_143,In_717);
or U4847 (N_4847,In_821,In_154);
and U4848 (N_4848,In_156,In_79);
nor U4849 (N_4849,In_968,In_218);
nand U4850 (N_4850,In_999,In_241);
and U4851 (N_4851,In_57,In_118);
nand U4852 (N_4852,In_98,In_854);
nand U4853 (N_4853,In_702,In_209);
or U4854 (N_4854,In_25,In_181);
nand U4855 (N_4855,In_769,In_630);
xnor U4856 (N_4856,In_312,In_954);
or U4857 (N_4857,In_417,In_26);
nand U4858 (N_4858,In_500,In_95);
and U4859 (N_4859,In_661,In_533);
nor U4860 (N_4860,In_407,In_342);
nor U4861 (N_4861,In_375,In_656);
and U4862 (N_4862,In_208,In_43);
and U4863 (N_4863,In_95,In_411);
nor U4864 (N_4864,In_685,In_646);
nand U4865 (N_4865,In_746,In_475);
and U4866 (N_4866,In_836,In_157);
nor U4867 (N_4867,In_670,In_382);
nor U4868 (N_4868,In_672,In_183);
or U4869 (N_4869,In_598,In_326);
or U4870 (N_4870,In_81,In_472);
or U4871 (N_4871,In_243,In_711);
and U4872 (N_4872,In_369,In_299);
nand U4873 (N_4873,In_584,In_418);
or U4874 (N_4874,In_237,In_503);
nand U4875 (N_4875,In_468,In_961);
nand U4876 (N_4876,In_566,In_155);
and U4877 (N_4877,In_346,In_892);
nor U4878 (N_4878,In_519,In_963);
or U4879 (N_4879,In_16,In_695);
nor U4880 (N_4880,In_940,In_20);
or U4881 (N_4881,In_507,In_514);
nand U4882 (N_4882,In_748,In_17);
or U4883 (N_4883,In_102,In_553);
xnor U4884 (N_4884,In_543,In_162);
and U4885 (N_4885,In_857,In_837);
or U4886 (N_4886,In_494,In_346);
nor U4887 (N_4887,In_610,In_36);
nand U4888 (N_4888,In_877,In_953);
nand U4889 (N_4889,In_63,In_592);
nand U4890 (N_4890,In_29,In_36);
and U4891 (N_4891,In_127,In_21);
and U4892 (N_4892,In_2,In_182);
or U4893 (N_4893,In_95,In_10);
nand U4894 (N_4894,In_101,In_256);
nand U4895 (N_4895,In_791,In_778);
or U4896 (N_4896,In_657,In_205);
nand U4897 (N_4897,In_838,In_947);
nand U4898 (N_4898,In_120,In_564);
and U4899 (N_4899,In_924,In_428);
nand U4900 (N_4900,In_789,In_277);
and U4901 (N_4901,In_94,In_875);
nor U4902 (N_4902,In_772,In_933);
and U4903 (N_4903,In_159,In_567);
nand U4904 (N_4904,In_400,In_668);
or U4905 (N_4905,In_762,In_676);
nand U4906 (N_4906,In_572,In_127);
and U4907 (N_4907,In_196,In_559);
and U4908 (N_4908,In_725,In_73);
and U4909 (N_4909,In_137,In_0);
or U4910 (N_4910,In_395,In_514);
nand U4911 (N_4911,In_753,In_140);
and U4912 (N_4912,In_20,In_159);
or U4913 (N_4913,In_813,In_462);
or U4914 (N_4914,In_800,In_60);
and U4915 (N_4915,In_394,In_732);
or U4916 (N_4916,In_887,In_369);
nand U4917 (N_4917,In_180,In_47);
nand U4918 (N_4918,In_467,In_511);
and U4919 (N_4919,In_17,In_183);
nand U4920 (N_4920,In_891,In_442);
and U4921 (N_4921,In_571,In_369);
nand U4922 (N_4922,In_104,In_592);
and U4923 (N_4923,In_892,In_195);
and U4924 (N_4924,In_920,In_772);
and U4925 (N_4925,In_930,In_944);
nor U4926 (N_4926,In_342,In_371);
or U4927 (N_4927,In_323,In_782);
and U4928 (N_4928,In_559,In_157);
nand U4929 (N_4929,In_754,In_728);
nor U4930 (N_4930,In_743,In_897);
and U4931 (N_4931,In_415,In_574);
or U4932 (N_4932,In_193,In_518);
and U4933 (N_4933,In_259,In_683);
nor U4934 (N_4934,In_801,In_862);
xnor U4935 (N_4935,In_565,In_372);
or U4936 (N_4936,In_195,In_828);
nand U4937 (N_4937,In_588,In_899);
nand U4938 (N_4938,In_924,In_625);
and U4939 (N_4939,In_972,In_646);
nand U4940 (N_4940,In_624,In_293);
nor U4941 (N_4941,In_736,In_171);
nor U4942 (N_4942,In_779,In_21);
nor U4943 (N_4943,In_270,In_952);
or U4944 (N_4944,In_759,In_83);
and U4945 (N_4945,In_911,In_332);
and U4946 (N_4946,In_454,In_433);
nor U4947 (N_4947,In_985,In_923);
nor U4948 (N_4948,In_13,In_579);
or U4949 (N_4949,In_222,In_458);
nand U4950 (N_4950,In_732,In_123);
or U4951 (N_4951,In_788,In_554);
or U4952 (N_4952,In_501,In_887);
nand U4953 (N_4953,In_148,In_660);
or U4954 (N_4954,In_256,In_422);
nand U4955 (N_4955,In_50,In_634);
nand U4956 (N_4956,In_33,In_88);
or U4957 (N_4957,In_970,In_988);
nand U4958 (N_4958,In_5,In_883);
nand U4959 (N_4959,In_936,In_855);
nand U4960 (N_4960,In_782,In_409);
xor U4961 (N_4961,In_863,In_436);
or U4962 (N_4962,In_396,In_587);
or U4963 (N_4963,In_567,In_911);
or U4964 (N_4964,In_482,In_74);
and U4965 (N_4965,In_869,In_476);
and U4966 (N_4966,In_319,In_464);
or U4967 (N_4967,In_982,In_422);
xnor U4968 (N_4968,In_976,In_681);
nor U4969 (N_4969,In_505,In_835);
nand U4970 (N_4970,In_946,In_733);
and U4971 (N_4971,In_259,In_622);
nor U4972 (N_4972,In_16,In_557);
xor U4973 (N_4973,In_0,In_170);
nor U4974 (N_4974,In_155,In_367);
and U4975 (N_4975,In_203,In_488);
nor U4976 (N_4976,In_49,In_446);
nand U4977 (N_4977,In_804,In_743);
or U4978 (N_4978,In_548,In_217);
nand U4979 (N_4979,In_565,In_513);
or U4980 (N_4980,In_532,In_328);
and U4981 (N_4981,In_801,In_72);
or U4982 (N_4982,In_777,In_947);
nand U4983 (N_4983,In_521,In_150);
nor U4984 (N_4984,In_475,In_77);
or U4985 (N_4985,In_579,In_3);
and U4986 (N_4986,In_840,In_440);
nor U4987 (N_4987,In_324,In_113);
xnor U4988 (N_4988,In_944,In_700);
nand U4989 (N_4989,In_874,In_290);
or U4990 (N_4990,In_148,In_395);
and U4991 (N_4991,In_334,In_58);
nor U4992 (N_4992,In_768,In_220);
nand U4993 (N_4993,In_25,In_95);
nand U4994 (N_4994,In_900,In_421);
nor U4995 (N_4995,In_636,In_481);
nand U4996 (N_4996,In_315,In_985);
nand U4997 (N_4997,In_678,In_872);
nor U4998 (N_4998,In_778,In_150);
or U4999 (N_4999,In_994,In_505);
nand U5000 (N_5000,N_364,N_3388);
or U5001 (N_5001,N_2364,N_4765);
and U5002 (N_5002,N_2140,N_3083);
nor U5003 (N_5003,N_1766,N_4709);
nor U5004 (N_5004,N_1900,N_1392);
or U5005 (N_5005,N_185,N_1922);
nor U5006 (N_5006,N_1435,N_4979);
nand U5007 (N_5007,N_2860,N_3853);
or U5008 (N_5008,N_3005,N_2622);
and U5009 (N_5009,N_2348,N_3706);
and U5010 (N_5010,N_1996,N_4872);
or U5011 (N_5011,N_4427,N_2529);
or U5012 (N_5012,N_2009,N_3798);
or U5013 (N_5013,N_3828,N_1528);
nor U5014 (N_5014,N_51,N_721);
nand U5015 (N_5015,N_3529,N_3666);
xnor U5016 (N_5016,N_2427,N_4155);
or U5017 (N_5017,N_309,N_752);
and U5018 (N_5018,N_3258,N_1880);
nand U5019 (N_5019,N_2807,N_1669);
and U5020 (N_5020,N_4624,N_4336);
and U5021 (N_5021,N_1445,N_4177);
and U5022 (N_5022,N_32,N_4033);
or U5023 (N_5023,N_1191,N_1491);
nand U5024 (N_5024,N_546,N_3033);
nor U5025 (N_5025,N_2127,N_1493);
and U5026 (N_5026,N_1373,N_4063);
nor U5027 (N_5027,N_3653,N_4272);
nor U5028 (N_5028,N_523,N_4157);
nor U5029 (N_5029,N_2870,N_2318);
or U5030 (N_5030,N_235,N_3262);
or U5031 (N_5031,N_1647,N_306);
or U5032 (N_5032,N_307,N_4262);
nor U5033 (N_5033,N_1292,N_2800);
or U5034 (N_5034,N_535,N_2926);
nor U5035 (N_5035,N_520,N_2459);
nand U5036 (N_5036,N_4524,N_2243);
and U5037 (N_5037,N_1122,N_1472);
nor U5038 (N_5038,N_1141,N_694);
and U5039 (N_5039,N_3581,N_2681);
nand U5040 (N_5040,N_237,N_2828);
nand U5041 (N_5041,N_3183,N_3990);
and U5042 (N_5042,N_4257,N_3191);
and U5043 (N_5043,N_2306,N_2324);
or U5044 (N_5044,N_3310,N_275);
xnor U5045 (N_5045,N_4736,N_945);
or U5046 (N_5046,N_3435,N_1116);
and U5047 (N_5047,N_3279,N_4369);
or U5048 (N_5048,N_2830,N_4808);
and U5049 (N_5049,N_1350,N_3969);
and U5050 (N_5050,N_1746,N_1813);
nand U5051 (N_5051,N_1225,N_4946);
or U5052 (N_5052,N_3359,N_2301);
and U5053 (N_5053,N_1474,N_4529);
nor U5054 (N_5054,N_2871,N_4040);
and U5055 (N_5055,N_4732,N_1836);
or U5056 (N_5056,N_2637,N_2510);
and U5057 (N_5057,N_1312,N_3655);
and U5058 (N_5058,N_1018,N_2541);
or U5059 (N_5059,N_4647,N_3958);
or U5060 (N_5060,N_638,N_1561);
and U5061 (N_5061,N_565,N_1741);
nor U5062 (N_5062,N_4803,N_3139);
and U5063 (N_5063,N_4539,N_1728);
and U5064 (N_5064,N_4756,N_3902);
and U5065 (N_5065,N_1654,N_696);
and U5066 (N_5066,N_1261,N_545);
or U5067 (N_5067,N_1840,N_3142);
nand U5068 (N_5068,N_4982,N_2157);
and U5069 (N_5069,N_2922,N_3304);
nand U5070 (N_5070,N_796,N_4285);
nand U5071 (N_5071,N_2073,N_314);
and U5072 (N_5072,N_1533,N_3732);
and U5073 (N_5073,N_238,N_4408);
or U5074 (N_5074,N_1989,N_422);
or U5075 (N_5075,N_1040,N_4201);
or U5076 (N_5076,N_849,N_2381);
and U5077 (N_5077,N_1185,N_2469);
and U5078 (N_5078,N_706,N_947);
nand U5079 (N_5079,N_2095,N_4772);
and U5080 (N_5080,N_398,N_155);
nor U5081 (N_5081,N_1558,N_3146);
nor U5082 (N_5082,N_2258,N_3463);
or U5083 (N_5083,N_2919,N_1685);
nand U5084 (N_5084,N_2936,N_2868);
and U5085 (N_5085,N_4282,N_3194);
or U5086 (N_5086,N_3626,N_551);
nor U5087 (N_5087,N_190,N_1497);
nand U5088 (N_5088,N_1991,N_3839);
or U5089 (N_5089,N_2528,N_1012);
nor U5090 (N_5090,N_4092,N_588);
or U5091 (N_5091,N_47,N_279);
nand U5092 (N_5092,N_4221,N_3862);
and U5093 (N_5093,N_3547,N_2779);
and U5094 (N_5094,N_1452,N_746);
and U5095 (N_5095,N_1406,N_338);
nor U5096 (N_5096,N_2651,N_1219);
and U5097 (N_5097,N_1213,N_2012);
xor U5098 (N_5098,N_3078,N_3336);
or U5099 (N_5099,N_3992,N_278);
and U5100 (N_5100,N_1448,N_1438);
and U5101 (N_5101,N_4975,N_1439);
or U5102 (N_5102,N_2222,N_1340);
nand U5103 (N_5103,N_438,N_2092);
or U5104 (N_5104,N_3170,N_3491);
nor U5105 (N_5105,N_4650,N_99);
nand U5106 (N_5106,N_1961,N_4217);
nand U5107 (N_5107,N_4036,N_1098);
or U5108 (N_5108,N_879,N_1341);
xnor U5109 (N_5109,N_3343,N_378);
and U5110 (N_5110,N_1658,N_641);
or U5111 (N_5111,N_997,N_4591);
or U5112 (N_5112,N_2424,N_3207);
nor U5113 (N_5113,N_905,N_825);
and U5114 (N_5114,N_3891,N_649);
nor U5115 (N_5115,N_3549,N_2239);
or U5116 (N_5116,N_4853,N_4673);
nand U5117 (N_5117,N_1987,N_2975);
or U5118 (N_5118,N_2123,N_90);
and U5119 (N_5119,N_762,N_2718);
and U5120 (N_5120,N_1867,N_487);
and U5121 (N_5121,N_2696,N_2250);
nor U5122 (N_5122,N_1982,N_1364);
or U5123 (N_5123,N_4125,N_3273);
or U5124 (N_5124,N_3895,N_1200);
nand U5125 (N_5125,N_4963,N_3120);
nand U5126 (N_5126,N_3269,N_4644);
nor U5127 (N_5127,N_1894,N_2313);
nor U5128 (N_5128,N_2628,N_2767);
and U5129 (N_5129,N_428,N_4315);
or U5130 (N_5130,N_2988,N_1168);
nor U5131 (N_5131,N_3582,N_4542);
nor U5132 (N_5132,N_4555,N_3180);
or U5133 (N_5133,N_1875,N_2168);
nand U5134 (N_5134,N_3603,N_1333);
nor U5135 (N_5135,N_679,N_4120);
nor U5136 (N_5136,N_4871,N_2395);
nor U5137 (N_5137,N_1915,N_351);
and U5138 (N_5138,N_4466,N_4099);
and U5139 (N_5139,N_2846,N_2064);
nor U5140 (N_5140,N_1120,N_4609);
or U5141 (N_5141,N_882,N_1831);
nor U5142 (N_5142,N_1635,N_3757);
nor U5143 (N_5143,N_4997,N_1864);
and U5144 (N_5144,N_1718,N_2575);
nand U5145 (N_5145,N_2247,N_2474);
or U5146 (N_5146,N_1810,N_2037);
or U5147 (N_5147,N_807,N_2107);
or U5148 (N_5148,N_2795,N_3540);
nand U5149 (N_5149,N_2408,N_2264);
nand U5150 (N_5150,N_1837,N_3222);
and U5151 (N_5151,N_800,N_2791);
nor U5152 (N_5152,N_4925,N_2697);
or U5153 (N_5153,N_2773,N_153);
nand U5154 (N_5154,N_3617,N_4522);
or U5155 (N_5155,N_4265,N_2735);
and U5156 (N_5156,N_30,N_4324);
and U5157 (N_5157,N_108,N_1890);
nor U5158 (N_5158,N_967,N_3885);
nand U5159 (N_5159,N_3133,N_4737);
nand U5160 (N_5160,N_683,N_748);
nor U5161 (N_5161,N_836,N_3487);
and U5162 (N_5162,N_3389,N_3206);
nand U5163 (N_5163,N_1304,N_171);
and U5164 (N_5164,N_2151,N_2670);
and U5165 (N_5165,N_1357,N_4258);
xor U5166 (N_5166,N_3478,N_2603);
nand U5167 (N_5167,N_3884,N_2928);
nand U5168 (N_5168,N_4064,N_1817);
or U5169 (N_5169,N_615,N_1955);
or U5170 (N_5170,N_1115,N_397);
or U5171 (N_5171,N_4831,N_2385);
xor U5172 (N_5172,N_2553,N_990);
nor U5173 (N_5173,N_3574,N_1949);
nand U5174 (N_5174,N_1471,N_3450);
nand U5175 (N_5175,N_3668,N_212);
or U5176 (N_5176,N_2354,N_3621);
nand U5177 (N_5177,N_3227,N_1787);
nor U5178 (N_5178,N_3234,N_3496);
or U5179 (N_5179,N_2196,N_4194);
nand U5180 (N_5180,N_335,N_3260);
or U5181 (N_5181,N_1503,N_1740);
or U5182 (N_5182,N_2625,N_4735);
and U5183 (N_5183,N_1873,N_579);
or U5184 (N_5184,N_2024,N_1593);
and U5185 (N_5185,N_2366,N_4405);
or U5186 (N_5186,N_702,N_3953);
nor U5187 (N_5187,N_4047,N_45);
or U5188 (N_5188,N_3531,N_4031);
or U5189 (N_5189,N_3254,N_3879);
or U5190 (N_5190,N_1466,N_2129);
nand U5191 (N_5191,N_4478,N_1101);
nand U5192 (N_5192,N_1090,N_2624);
or U5193 (N_5193,N_722,N_1268);
nand U5194 (N_5194,N_341,N_1110);
nor U5195 (N_5195,N_1283,N_2498);
nand U5196 (N_5196,N_270,N_2524);
or U5197 (N_5197,N_1904,N_43);
or U5198 (N_5198,N_1693,N_1828);
nor U5199 (N_5199,N_2494,N_65);
nand U5200 (N_5200,N_1723,N_1286);
xnor U5201 (N_5201,N_3930,N_24);
or U5202 (N_5202,N_2439,N_1086);
nor U5203 (N_5203,N_2475,N_3831);
or U5204 (N_5204,N_2406,N_1396);
or U5205 (N_5205,N_2193,N_3345);
and U5206 (N_5206,N_699,N_4331);
and U5207 (N_5207,N_861,N_1580);
nand U5208 (N_5208,N_3964,N_2048);
or U5209 (N_5209,N_713,N_1211);
and U5210 (N_5210,N_4788,N_1829);
nand U5211 (N_5211,N_3319,N_2608);
nand U5212 (N_5212,N_2332,N_1198);
or U5213 (N_5213,N_4606,N_3316);
nand U5214 (N_5214,N_4384,N_2956);
or U5215 (N_5215,N_1737,N_3098);
and U5216 (N_5216,N_3019,N_4206);
nand U5217 (N_5217,N_223,N_4859);
nor U5218 (N_5218,N_466,N_2461);
nand U5219 (N_5219,N_2465,N_3628);
nor U5220 (N_5220,N_3469,N_926);
xor U5221 (N_5221,N_105,N_2714);
xor U5222 (N_5222,N_1372,N_2421);
nand U5223 (N_5223,N_2104,N_431);
and U5224 (N_5224,N_2191,N_1260);
and U5225 (N_5225,N_3759,N_899);
and U5226 (N_5226,N_39,N_1517);
nand U5227 (N_5227,N_2548,N_1711);
nor U5228 (N_5228,N_4549,N_4464);
nand U5229 (N_5229,N_712,N_3820);
nand U5230 (N_5230,N_3165,N_3625);
nor U5231 (N_5231,N_2485,N_433);
or U5232 (N_5232,N_350,N_4860);
nand U5233 (N_5233,N_1221,N_2817);
or U5234 (N_5234,N_4132,N_4573);
and U5235 (N_5235,N_1006,N_4163);
or U5236 (N_5236,N_3767,N_1031);
or U5237 (N_5237,N_2454,N_4188);
and U5238 (N_5238,N_1699,N_2547);
nor U5239 (N_5239,N_2317,N_424);
nor U5240 (N_5240,N_86,N_1182);
and U5241 (N_5241,N_3132,N_3486);
nand U5242 (N_5242,N_4538,N_1251);
or U5243 (N_5243,N_1770,N_2911);
and U5244 (N_5244,N_1055,N_4355);
and U5245 (N_5245,N_2458,N_4800);
nor U5246 (N_5246,N_4560,N_3093);
nor U5247 (N_5247,N_818,N_3114);
nand U5248 (N_5248,N_2434,N_710);
nor U5249 (N_5249,N_297,N_1725);
nand U5250 (N_5250,N_4008,N_4395);
or U5251 (N_5251,N_4114,N_685);
and U5252 (N_5252,N_4920,N_4247);
and U5253 (N_5253,N_4884,N_1639);
or U5254 (N_5254,N_2367,N_4564);
nand U5255 (N_5255,N_291,N_21);
nand U5256 (N_5256,N_46,N_4865);
nor U5257 (N_5257,N_2550,N_4356);
or U5258 (N_5258,N_3334,N_4182);
and U5259 (N_5259,N_1895,N_4806);
xnor U5260 (N_5260,N_4172,N_1087);
xnor U5261 (N_5261,N_3701,N_290);
nor U5262 (N_5262,N_4437,N_4081);
nand U5263 (N_5263,N_91,N_289);
nor U5264 (N_5264,N_4143,N_3841);
and U5265 (N_5265,N_4722,N_3330);
nor U5266 (N_5266,N_126,N_1719);
nor U5267 (N_5267,N_3850,N_3144);
or U5268 (N_5268,N_4419,N_3810);
nor U5269 (N_5269,N_1908,N_4096);
nor U5270 (N_5270,N_3804,N_2754);
and U5271 (N_5271,N_1407,N_4115);
nand U5272 (N_5272,N_1710,N_742);
xnor U5273 (N_5273,N_964,N_3278);
nand U5274 (N_5274,N_2588,N_4377);
nor U5275 (N_5275,N_4433,N_4705);
and U5276 (N_5276,N_2610,N_4232);
nor U5277 (N_5277,N_2057,N_654);
nor U5278 (N_5278,N_3061,N_3023);
nor U5279 (N_5279,N_2780,N_3638);
nand U5280 (N_5280,N_3454,N_4986);
or U5281 (N_5281,N_3792,N_3899);
and U5282 (N_5282,N_2914,N_3312);
nor U5283 (N_5283,N_788,N_1415);
and U5284 (N_5284,N_4202,N_1887);
or U5285 (N_5285,N_224,N_4826);
nor U5286 (N_5286,N_4747,N_2045);
or U5287 (N_5287,N_2294,N_3199);
or U5288 (N_5288,N_1431,N_2199);
or U5289 (N_5289,N_1679,N_3569);
nand U5290 (N_5290,N_3918,N_409);
or U5291 (N_5291,N_4291,N_591);
nor U5292 (N_5292,N_4415,N_3699);
and U5293 (N_5293,N_1671,N_4337);
xor U5294 (N_5294,N_3838,N_4868);
and U5295 (N_5295,N_3662,N_1072);
and U5296 (N_5296,N_2020,N_2314);
and U5297 (N_5297,N_548,N_1147);
nor U5298 (N_5298,N_4128,N_2738);
nor U5299 (N_5299,N_1347,N_301);
nand U5300 (N_5300,N_1868,N_1180);
or U5301 (N_5301,N_4948,N_328);
or U5302 (N_5302,N_347,N_2197);
or U5303 (N_5303,N_1194,N_2563);
nor U5304 (N_5304,N_1481,N_3054);
or U5305 (N_5305,N_3016,N_1743);
or U5306 (N_5306,N_2874,N_2456);
and U5307 (N_5307,N_1485,N_4334);
nor U5308 (N_5308,N_4242,N_2235);
and U5309 (N_5309,N_1425,N_1351);
nand U5310 (N_5310,N_3597,N_2600);
nand U5311 (N_5311,N_196,N_3137);
or U5312 (N_5312,N_3742,N_4526);
and U5313 (N_5313,N_2182,N_4276);
and U5314 (N_5314,N_4267,N_2666);
and U5315 (N_5315,N_4319,N_1564);
or U5316 (N_5316,N_4245,N_3242);
nand U5317 (N_5317,N_3538,N_4911);
or U5318 (N_5318,N_2504,N_1729);
nand U5319 (N_5319,N_2983,N_3426);
nand U5320 (N_5320,N_559,N_3399);
nor U5321 (N_5321,N_1322,N_1834);
and U5322 (N_5322,N_4779,N_456);
nand U5323 (N_5323,N_3593,N_2296);
and U5324 (N_5324,N_906,N_2763);
and U5325 (N_5325,N_3657,N_4583);
nand U5326 (N_5326,N_2288,N_310);
nor U5327 (N_5327,N_2941,N_2816);
and U5328 (N_5328,N_1751,N_3360);
and U5329 (N_5329,N_630,N_1660);
and U5330 (N_5330,N_3664,N_1239);
nor U5331 (N_5331,N_31,N_2668);
or U5332 (N_5332,N_4210,N_2977);
or U5333 (N_5333,N_3072,N_1331);
nand U5334 (N_5334,N_1557,N_4670);
nor U5335 (N_5335,N_2841,N_3716);
nor U5336 (N_5336,N_1428,N_1796);
and U5337 (N_5337,N_2530,N_3419);
and U5338 (N_5338,N_3353,N_2915);
nor U5339 (N_5339,N_3289,N_2233);
and U5340 (N_5340,N_3494,N_2108);
and U5341 (N_5341,N_2279,N_1325);
nor U5342 (N_5342,N_4281,N_56);
nor U5343 (N_5343,N_3746,N_3173);
nand U5344 (N_5344,N_2230,N_736);
nor U5345 (N_5345,N_440,N_2620);
nand U5346 (N_5346,N_1627,N_3584);
or U5347 (N_5347,N_3843,N_3980);
and U5348 (N_5348,N_4418,N_553);
and U5349 (N_5349,N_4869,N_603);
or U5350 (N_5350,N_4049,N_4898);
and U5351 (N_5351,N_3109,N_140);
and U5352 (N_5352,N_236,N_2353);
and U5353 (N_5353,N_1231,N_690);
nand U5354 (N_5354,N_3298,N_1019);
and U5355 (N_5355,N_4776,N_589);
and U5356 (N_5356,N_3246,N_110);
nand U5357 (N_5357,N_427,N_3718);
nand U5358 (N_5358,N_525,N_360);
nor U5359 (N_5359,N_640,N_544);
or U5360 (N_5360,N_1427,N_4752);
or U5361 (N_5361,N_131,N_2591);
nor U5362 (N_5362,N_1551,N_910);
nand U5363 (N_5363,N_3158,N_3393);
nand U5364 (N_5364,N_1927,N_4508);
or U5365 (N_5365,N_222,N_542);
and U5366 (N_5366,N_3119,N_4795);
xnor U5367 (N_5367,N_453,N_819);
and U5368 (N_5368,N_4461,N_1600);
nand U5369 (N_5369,N_2452,N_2244);
xor U5370 (N_5370,N_1010,N_1637);
or U5371 (N_5371,N_1898,N_2555);
nand U5372 (N_5372,N_3602,N_3669);
nor U5373 (N_5373,N_3274,N_2007);
and U5374 (N_5374,N_3167,N_2274);
nand U5375 (N_5375,N_883,N_1818);
or U5376 (N_5376,N_856,N_4373);
nand U5377 (N_5377,N_1986,N_1527);
nor U5378 (N_5378,N_2811,N_4026);
nand U5379 (N_5379,N_1222,N_2105);
nand U5380 (N_5380,N_1608,N_2695);
nor U5381 (N_5381,N_4957,N_4828);
and U5382 (N_5382,N_1575,N_759);
and U5383 (N_5383,N_1158,N_2721);
nand U5384 (N_5384,N_614,N_1423);
nor U5385 (N_5385,N_1815,N_3760);
nor U5386 (N_5386,N_4711,N_3526);
or U5387 (N_5387,N_4003,N_4055);
nor U5388 (N_5388,N_4045,N_2984);
and U5389 (N_5389,N_519,N_4578);
nor U5390 (N_5390,N_4955,N_3338);
nand U5391 (N_5391,N_2925,N_1977);
xnor U5392 (N_5392,N_3643,N_2303);
nand U5393 (N_5393,N_3615,N_3413);
nand U5394 (N_5394,N_2166,N_4745);
or U5395 (N_5395,N_2701,N_560);
and U5396 (N_5396,N_3741,N_2505);
nor U5397 (N_5397,N_570,N_1562);
and U5398 (N_5398,N_3344,N_3280);
nor U5399 (N_5399,N_75,N_3103);
nor U5400 (N_5400,N_4543,N_4509);
nor U5401 (N_5401,N_3204,N_2599);
nor U5402 (N_5402,N_2497,N_4556);
and U5403 (N_5403,N_1084,N_2609);
and U5404 (N_5404,N_3765,N_953);
nor U5405 (N_5405,N_1498,N_1936);
and U5406 (N_5406,N_2124,N_1852);
or U5407 (N_5407,N_709,N_4175);
and U5408 (N_5408,N_2520,N_3160);
nor U5409 (N_5409,N_593,N_2938);
nor U5410 (N_5410,N_87,N_831);
or U5411 (N_5411,N_4615,N_2295);
nand U5412 (N_5412,N_353,N_2085);
and U5413 (N_5413,N_4195,N_1444);
nor U5414 (N_5414,N_4004,N_207);
or U5415 (N_5415,N_2590,N_1583);
and U5416 (N_5416,N_3386,N_1342);
nor U5417 (N_5417,N_1210,N_1826);
xor U5418 (N_5418,N_2831,N_4619);
or U5419 (N_5419,N_1385,N_4900);
nor U5420 (N_5420,N_3445,N_1789);
and U5421 (N_5421,N_1310,N_2453);
nor U5422 (N_5422,N_4738,N_1942);
nor U5423 (N_5423,N_4571,N_4687);
or U5424 (N_5424,N_2745,N_1588);
or U5425 (N_5425,N_2298,N_2902);
or U5426 (N_5426,N_3202,N_4791);
or U5427 (N_5427,N_4138,N_2908);
nand U5428 (N_5428,N_4360,N_4332);
nor U5429 (N_5429,N_4296,N_2826);
or U5430 (N_5430,N_3795,N_605);
nor U5431 (N_5431,N_2570,N_4443);
or U5432 (N_5432,N_3975,N_326);
and U5433 (N_5433,N_4910,N_3397);
nor U5434 (N_5434,N_1749,N_1937);
or U5435 (N_5435,N_3239,N_3789);
nand U5436 (N_5436,N_3794,N_650);
or U5437 (N_5437,N_760,N_3863);
nor U5438 (N_5438,N_2751,N_3064);
nor U5439 (N_5439,N_4390,N_3402);
nor U5440 (N_5440,N_135,N_3115);
nor U5441 (N_5441,N_3238,N_1553);
nand U5442 (N_5442,N_4940,N_2357);
nand U5443 (N_5443,N_28,N_922);
nand U5444 (N_5444,N_2214,N_2210);
or U5445 (N_5445,N_239,N_599);
nand U5446 (N_5446,N_3288,N_2885);
and U5447 (N_5447,N_3307,N_859);
and U5448 (N_5448,N_4545,N_3368);
or U5449 (N_5449,N_1519,N_4027);
and U5450 (N_5450,N_1756,N_4180);
nand U5451 (N_5451,N_2046,N_2972);
nand U5452 (N_5452,N_4584,N_4783);
nor U5453 (N_5453,N_4227,N_4482);
nand U5454 (N_5454,N_935,N_1531);
or U5455 (N_5455,N_3906,N_1550);
or U5456 (N_5456,N_1138,N_1112);
and U5457 (N_5457,N_1137,N_2187);
and U5458 (N_5458,N_2596,N_4156);
nand U5459 (N_5459,N_1514,N_2835);
nand U5460 (N_5460,N_3162,N_804);
nor U5461 (N_5461,N_1689,N_4926);
or U5462 (N_5462,N_2909,N_4632);
or U5463 (N_5463,N_119,N_2967);
nand U5464 (N_5464,N_1494,N_3986);
nand U5465 (N_5465,N_485,N_2999);
nand U5466 (N_5466,N_1629,N_1577);
nand U5467 (N_5467,N_160,N_1074);
or U5468 (N_5468,N_123,N_3882);
xor U5469 (N_5469,N_4069,N_1193);
nand U5470 (N_5470,N_4091,N_1957);
nand U5471 (N_5471,N_107,N_3650);
nand U5472 (N_5472,N_3230,N_1050);
or U5473 (N_5473,N_3708,N_4347);
nand U5474 (N_5474,N_266,N_2825);
xor U5475 (N_5475,N_3504,N_1166);
and U5476 (N_5476,N_2019,N_4611);
and U5477 (N_5477,N_3104,N_2708);
or U5478 (N_5478,N_914,N_4107);
and U5479 (N_5479,N_758,N_3237);
xor U5480 (N_5480,N_2989,N_1784);
nand U5481 (N_5481,N_2158,N_1457);
and U5482 (N_5482,N_122,N_3177);
or U5483 (N_5483,N_3367,N_611);
or U5484 (N_5484,N_2694,N_3846);
or U5485 (N_5485,N_4000,N_1167);
and U5486 (N_5486,N_4567,N_120);
nand U5487 (N_5487,N_186,N_1504);
nor U5488 (N_5488,N_3020,N_776);
and U5489 (N_5489,N_661,N_3516);
nor U5490 (N_5490,N_705,N_4973);
and U5491 (N_5491,N_2473,N_2093);
nor U5492 (N_5492,N_568,N_4789);
nand U5493 (N_5493,N_533,N_4741);
and U5494 (N_5494,N_381,N_2812);
nand U5495 (N_5495,N_1139,N_3335);
or U5496 (N_5496,N_867,N_4794);
or U5497 (N_5497,N_3609,N_4896);
xnor U5498 (N_5498,N_3284,N_2358);
and U5499 (N_5499,N_4820,N_3646);
or U5500 (N_5500,N_1204,N_566);
and U5501 (N_5501,N_2809,N_3339);
nor U5502 (N_5502,N_3954,N_4454);
nor U5503 (N_5503,N_3872,N_4116);
nor U5504 (N_5504,N_233,N_4974);
nand U5505 (N_5505,N_4527,N_2781);
nor U5506 (N_5506,N_952,N_3126);
nand U5507 (N_5507,N_3658,N_4046);
or U5508 (N_5508,N_1638,N_4448);
nor U5509 (N_5509,N_2951,N_4024);
nor U5510 (N_5510,N_3156,N_2815);
nor U5511 (N_5511,N_3989,N_2516);
nand U5512 (N_5512,N_3155,N_384);
nand U5513 (N_5513,N_383,N_3743);
nor U5514 (N_5514,N_731,N_4661);
or U5515 (N_5515,N_2058,N_4029);
or U5516 (N_5516,N_3927,N_4495);
nor U5517 (N_5517,N_4298,N_2645);
and U5518 (N_5518,N_4187,N_1052);
and U5519 (N_5519,N_3729,N_170);
or U5520 (N_5520,N_2177,N_4459);
nand U5521 (N_5521,N_1911,N_3976);
nand U5522 (N_5522,N_2017,N_2282);
and U5523 (N_5523,N_2029,N_4421);
nor U5524 (N_5524,N_3580,N_3942);
and U5525 (N_5525,N_2380,N_2665);
and U5526 (N_5526,N_2750,N_3123);
nor U5527 (N_5527,N_2878,N_2340);
or U5528 (N_5528,N_1590,N_1603);
or U5529 (N_5529,N_3713,N_1739);
nand U5530 (N_5530,N_4858,N_4981);
and U5531 (N_5531,N_142,N_794);
nor U5532 (N_5532,N_4013,N_3755);
nand U5533 (N_5533,N_4700,N_4060);
or U5534 (N_5534,N_1237,N_2884);
nand U5535 (N_5535,N_4876,N_4304);
or U5536 (N_5536,N_154,N_1604);
xor U5537 (N_5537,N_2960,N_747);
nand U5538 (N_5538,N_627,N_4707);
or U5539 (N_5539,N_4716,N_1107);
or U5540 (N_5540,N_4639,N_1378);
or U5541 (N_5541,N_2521,N_320);
and U5542 (N_5542,N_3842,N_1480);
nor U5543 (N_5543,N_2040,N_1633);
nand U5544 (N_5544,N_816,N_444);
nor U5545 (N_5545,N_1674,N_569);
or U5546 (N_5546,N_3176,N_1832);
nor U5547 (N_5547,N_4229,N_943);
nand U5548 (N_5548,N_4111,N_3203);
nand U5549 (N_5549,N_248,N_1458);
or U5550 (N_5550,N_837,N_567);
nand U5551 (N_5551,N_4603,N_3875);
nor U5552 (N_5552,N_4553,N_2713);
or U5553 (N_5553,N_4637,N_1259);
or U5554 (N_5554,N_2111,N_4152);
nor U5555 (N_5555,N_3205,N_4271);
and U5556 (N_5556,N_1142,N_4622);
or U5557 (N_5557,N_2478,N_2818);
nor U5558 (N_5558,N_4368,N_4617);
nand U5559 (N_5559,N_3816,N_48);
and U5560 (N_5560,N_4598,N_978);
nand U5561 (N_5561,N_4387,N_2221);
nor U5562 (N_5562,N_2267,N_3805);
nand U5563 (N_5563,N_4016,N_4321);
nor U5564 (N_5564,N_3769,N_2141);
xor U5565 (N_5565,N_4062,N_2854);
nand U5566 (N_5566,N_1702,N_3350);
nor U5567 (N_5567,N_136,N_2717);
or U5568 (N_5568,N_3225,N_1652);
nor U5569 (N_5569,N_2643,N_561);
nor U5570 (N_5570,N_284,N_241);
and U5571 (N_5571,N_4328,N_3545);
and U5572 (N_5572,N_4083,N_4226);
or U5573 (N_5573,N_2576,N_3629);
nor U5574 (N_5574,N_4102,N_3517);
or U5575 (N_5575,N_2171,N_4058);
nor U5576 (N_5576,N_4780,N_1215);
nor U5577 (N_5577,N_3575,N_4947);
xnor U5578 (N_5578,N_232,N_4101);
or U5579 (N_5579,N_813,N_3346);
nor U5580 (N_5580,N_1290,N_1666);
nor U5581 (N_5581,N_3524,N_4557);
nand U5582 (N_5582,N_1368,N_3086);
nor U5583 (N_5583,N_4365,N_125);
nand U5584 (N_5584,N_1806,N_152);
nand U5585 (N_5585,N_729,N_3901);
nand U5586 (N_5586,N_4778,N_3196);
nor U5587 (N_5587,N_625,N_1014);
xor U5588 (N_5588,N_3553,N_4667);
or U5589 (N_5589,N_4873,N_1404);
or U5590 (N_5590,N_1667,N_754);
or U5591 (N_5591,N_821,N_2627);
nor U5592 (N_5592,N_667,N_1684);
and U5593 (N_5593,N_3101,N_1998);
nand U5594 (N_5594,N_669,N_2175);
or U5595 (N_5595,N_4176,N_4525);
nor U5596 (N_5596,N_2752,N_2648);
and U5597 (N_5597,N_3017,N_2047);
and U5598 (N_5598,N_473,N_592);
nand U5599 (N_5599,N_3438,N_783);
or U5600 (N_5600,N_4412,N_426);
and U5601 (N_5601,N_2195,N_1397);
nand U5602 (N_5602,N_1620,N_2772);
nor U5603 (N_5603,N_2476,N_2100);
or U5604 (N_5604,N_3187,N_2998);
or U5605 (N_5605,N_4541,N_1302);
nand U5606 (N_5606,N_2011,N_3704);
nand U5607 (N_5607,N_1266,N_3200);
and U5608 (N_5608,N_4523,N_707);
or U5609 (N_5609,N_571,N_2667);
and U5610 (N_5610,N_1676,N_367);
and U5611 (N_5611,N_3147,N_2066);
nand U5612 (N_5612,N_3159,N_4654);
nor U5613 (N_5613,N_1569,N_2152);
nand U5614 (N_5614,N_4239,N_157);
xor U5615 (N_5615,N_247,N_4394);
nor U5616 (N_5616,N_2996,N_2139);
nor U5617 (N_5617,N_1119,N_1064);
and U5618 (N_5618,N_2392,N_1117);
xnor U5619 (N_5619,N_4253,N_1063);
nor U5620 (N_5620,N_3489,N_4462);
xnor U5621 (N_5621,N_3380,N_3936);
nor U5622 (N_5622,N_2273,N_373);
xnor U5623 (N_5623,N_4279,N_4894);
nand U5624 (N_5624,N_4372,N_1136);
nand U5625 (N_5625,N_1103,N_4839);
nand U5626 (N_5626,N_1812,N_3153);
nand U5627 (N_5627,N_1413,N_3472);
nor U5628 (N_5628,N_2704,N_2004);
and U5629 (N_5629,N_2272,N_1057);
nand U5630 (N_5630,N_4350,N_2562);
nand U5631 (N_5631,N_2448,N_2654);
and U5632 (N_5632,N_3400,N_2442);
nor U5633 (N_5633,N_4912,N_3324);
or U5634 (N_5634,N_1020,N_4883);
nand U5635 (N_5635,N_4701,N_4781);
nor U5636 (N_5636,N_4287,N_1499);
or U5637 (N_5637,N_1054,N_4230);
and U5638 (N_5638,N_2265,N_3698);
or U5639 (N_5639,N_1091,N_2142);
nand U5640 (N_5640,N_1980,N_3886);
and U5641 (N_5641,N_4958,N_838);
nand U5642 (N_5642,N_3856,N_1143);
and U5643 (N_5643,N_1863,N_1856);
and U5644 (N_5644,N_321,N_2837);
or U5645 (N_5645,N_4113,N_3859);
nand U5646 (N_5646,N_2343,N_3548);
and U5647 (N_5647,N_4616,N_3610);
and U5648 (N_5648,N_1849,N_3654);
nor U5649 (N_5649,N_3305,N_97);
nand U5650 (N_5650,N_4725,N_116);
nand U5651 (N_5651,N_1907,N_483);
nand U5652 (N_5652,N_1162,N_79);
nand U5653 (N_5653,N_4546,N_4108);
and U5654 (N_5654,N_4944,N_738);
nor U5655 (N_5655,N_1327,N_789);
nor U5656 (N_5656,N_4097,N_1944);
nor U5657 (N_5657,N_1509,N_3788);
or U5658 (N_5658,N_761,N_2774);
and U5659 (N_5659,N_1105,N_988);
and U5660 (N_5660,N_2137,N_3431);
or U5661 (N_5661,N_1346,N_3661);
nor U5662 (N_5662,N_4225,N_1616);
nand U5663 (N_5663,N_4706,N_3045);
and U5664 (N_5664,N_792,N_4693);
or U5665 (N_5665,N_3773,N_1555);
or U5666 (N_5666,N_4733,N_3908);
nor U5667 (N_5667,N_3753,N_396);
nand U5668 (N_5668,N_1681,N_4335);
and U5669 (N_5669,N_296,N_3189);
nor U5670 (N_5670,N_2790,N_2067);
and U5671 (N_5671,N_2194,N_733);
xor U5672 (N_5672,N_1314,N_3691);
or U5673 (N_5673,N_1628,N_1264);
and U5674 (N_5674,N_4893,N_887);
xor U5675 (N_5675,N_3572,N_1447);
nor U5676 (N_5676,N_972,N_797);
or U5677 (N_5677,N_4648,N_4048);
nor U5678 (N_5678,N_4274,N_2444);
nand U5679 (N_5679,N_4362,N_4145);
and U5680 (N_5680,N_4255,N_317);
or U5681 (N_5681,N_3263,N_4011);
nand U5682 (N_5682,N_658,N_3074);
nor U5683 (N_5683,N_1988,N_2634);
or U5684 (N_5684,N_2827,N_1518);
nand U5685 (N_5685,N_3848,N_4079);
nor U5686 (N_5686,N_2077,N_1173);
and U5687 (N_5687,N_3174,N_4140);
nand U5688 (N_5688,N_2991,N_2394);
and U5689 (N_5689,N_714,N_3300);
nand U5690 (N_5690,N_2937,N_4570);
and U5691 (N_5691,N_245,N_2890);
nand U5692 (N_5692,N_4683,N_213);
or U5693 (N_5693,N_2121,N_2892);
and U5694 (N_5694,N_940,N_2167);
or U5695 (N_5695,N_1421,N_3069);
nand U5696 (N_5696,N_1078,N_2180);
or U5697 (N_5697,N_3408,N_1296);
nand U5698 (N_5698,N_1178,N_3904);
or U5699 (N_5699,N_419,N_1701);
and U5700 (N_5700,N_1767,N_675);
or U5701 (N_5701,N_1934,N_4734);
nor U5702 (N_5702,N_3692,N_753);
nand U5703 (N_5703,N_527,N_955);
nor U5704 (N_5704,N_973,N_1794);
and U5705 (N_5705,N_2601,N_2234);
and U5706 (N_5706,N_4708,N_459);
or U5707 (N_5707,N_4497,N_2944);
or U5708 (N_5708,N_2644,N_891);
nor U5709 (N_5709,N_4753,N_1241);
and U5710 (N_5710,N_356,N_3981);
or U5711 (N_5711,N_4450,N_1974);
and U5712 (N_5712,N_55,N_2323);
or U5713 (N_5713,N_210,N_4014);
or U5714 (N_5714,N_872,N_2271);
nand U5715 (N_5715,N_2690,N_4769);
nand U5716 (N_5716,N_2917,N_711);
nor U5717 (N_5717,N_4098,N_4379);
or U5718 (N_5718,N_4671,N_2005);
nor U5719 (N_5719,N_2090,N_3303);
and U5720 (N_5720,N_1707,N_3152);
or U5721 (N_5721,N_3800,N_2087);
or U5722 (N_5722,N_2990,N_2312);
nor U5723 (N_5723,N_1981,N_4843);
or U5724 (N_5724,N_775,N_975);
and U5725 (N_5725,N_3608,N_3649);
and U5726 (N_5726,N_4740,N_1263);
nand U5727 (N_5727,N_323,N_1807);
nor U5728 (N_5728,N_3959,N_73);
or U5729 (N_5729,N_3720,N_1475);
and U5730 (N_5730,N_2684,N_750);
nor U5731 (N_5731,N_612,N_1434);
and U5732 (N_5732,N_3213,N_2316);
nor U5733 (N_5733,N_2675,N_1926);
nand U5734 (N_5734,N_745,N_4203);
and U5735 (N_5735,N_2880,N_3733);
nor U5736 (N_5736,N_1747,N_2613);
nor U5737 (N_5737,N_3209,N_2889);
nand U5738 (N_5738,N_44,N_1626);
nand U5739 (N_5739,N_3833,N_2577);
and U5740 (N_5740,N_2852,N_4434);
nor U5741 (N_5741,N_1104,N_898);
and U5742 (N_5742,N_4561,N_2933);
or U5743 (N_5743,N_2331,N_3821);
or U5744 (N_5744,N_267,N_3966);
nand U5745 (N_5745,N_4847,N_3080);
or U5746 (N_5746,N_4403,N_4193);
nand U5747 (N_5747,N_989,N_893);
or U5748 (N_5748,N_1526,N_172);
xor U5749 (N_5749,N_3880,N_2023);
and U5750 (N_5750,N_4095,N_3724);
nand U5751 (N_5751,N_4532,N_3326);
and U5752 (N_5752,N_2181,N_3049);
or U5753 (N_5753,N_4886,N_1370);
nand U5754 (N_5754,N_205,N_549);
and U5755 (N_5755,N_115,N_2404);
nand U5756 (N_5756,N_3216,N_639);
or U5757 (N_5757,N_2184,N_194);
xnor U5758 (N_5758,N_4939,N_1155);
or U5759 (N_5759,N_2631,N_2640);
xor U5760 (N_5760,N_3606,N_2039);
nor U5761 (N_5761,N_2050,N_3541);
nor U5762 (N_5762,N_2224,N_1933);
nand U5763 (N_5763,N_4146,N_4492);
or U5764 (N_5764,N_4676,N_3145);
nand U5765 (N_5765,N_4961,N_3261);
or U5766 (N_5766,N_1830,N_1262);
nand U5767 (N_5767,N_1203,N_2251);
nand U5768 (N_5768,N_2156,N_4645);
nor U5769 (N_5769,N_1939,N_3476);
and U5770 (N_5770,N_4825,N_4134);
nand U5771 (N_5771,N_524,N_176);
xnor U5772 (N_5772,N_1309,N_3221);
and U5773 (N_5773,N_790,N_2436);
nand U5774 (N_5774,N_261,N_3982);
nor U5775 (N_5775,N_2071,N_4782);
nor U5776 (N_5776,N_3432,N_1329);
and U5777 (N_5777,N_3534,N_1058);
nand U5778 (N_5778,N_1878,N_1151);
or U5779 (N_5779,N_877,N_942);
or U5780 (N_5780,N_4792,N_4656);
and U5781 (N_5781,N_2947,N_3715);
nor U5782 (N_5782,N_934,N_2200);
nor U5783 (N_5783,N_3240,N_749);
or U5784 (N_5784,N_3611,N_283);
and U5785 (N_5785,N_3392,N_1275);
nand U5786 (N_5786,N_1594,N_4684);
nor U5787 (N_5787,N_2897,N_1556);
or U5788 (N_5788,N_2567,N_672);
nand U5789 (N_5789,N_2607,N_2389);
nor U5790 (N_5790,N_62,N_3091);
or U5791 (N_5791,N_2001,N_2390);
nand U5792 (N_5792,N_4829,N_1113);
nand U5793 (N_5793,N_2270,N_3542);
or U5794 (N_5794,N_1967,N_4921);
nor U5795 (N_5795,N_3968,N_322);
and U5796 (N_5796,N_109,N_3802);
or U5797 (N_5797,N_2053,N_1479);
nand U5798 (N_5798,N_59,N_3328);
nand U5799 (N_5799,N_1170,N_1909);
nor U5800 (N_5800,N_2240,N_4118);
nand U5801 (N_5801,N_2535,N_585);
nand U5802 (N_5802,N_2653,N_4236);
nand U5803 (N_5803,N_1672,N_2307);
or U5804 (N_5804,N_3854,N_2397);
nand U5805 (N_5805,N_3488,N_1641);
and U5806 (N_5806,N_3296,N_3645);
and U5807 (N_5807,N_980,N_1048);
nor U5808 (N_5808,N_3223,N_3815);
and U5809 (N_5809,N_3825,N_2144);
or U5810 (N_5810,N_1636,N_552);
nand U5811 (N_5811,N_2076,N_4763);
or U5812 (N_5812,N_3051,N_1492);
nand U5813 (N_5813,N_1883,N_1884);
nor U5814 (N_5814,N_1768,N_265);
nand U5815 (N_5815,N_1319,N_269);
nand U5816 (N_5816,N_19,N_1469);
nand U5817 (N_5817,N_2810,N_4582);
nor U5818 (N_5818,N_303,N_4343);
nor U5819 (N_5819,N_3150,N_4754);
and U5820 (N_5820,N_619,N_4878);
nand U5821 (N_5821,N_3294,N_4980);
and U5822 (N_5822,N_474,N_164);
nand U5823 (N_5823,N_3616,N_1030);
or U5824 (N_5824,N_1081,N_252);
nor U5825 (N_5825,N_3149,N_1578);
nand U5826 (N_5826,N_3779,N_4080);
nor U5827 (N_5827,N_1935,N_1510);
or U5828 (N_5828,N_580,N_255);
nor U5829 (N_5829,N_2993,N_3363);
nand U5830 (N_5830,N_476,N_4363);
nand U5831 (N_5831,N_3317,N_1634);
nor U5832 (N_5832,N_4340,N_1866);
nand U5833 (N_5833,N_3070,N_1176);
nor U5834 (N_5834,N_631,N_256);
and U5835 (N_5835,N_3283,N_4838);
nor U5836 (N_5836,N_408,N_1405);
nor U5837 (N_5837,N_1083,N_2082);
xnor U5838 (N_5838,N_2446,N_451);
or U5839 (N_5839,N_4685,N_1696);
nor U5840 (N_5840,N_4550,N_217);
nand U5841 (N_5841,N_3201,N_3447);
and U5842 (N_5842,N_3869,N_4768);
nor U5843 (N_5843,N_3554,N_1038);
or U5844 (N_5844,N_101,N_3318);
nor U5845 (N_5845,N_3694,N_1242);
or U5846 (N_5846,N_3987,N_1360);
nand U5847 (N_5847,N_2382,N_1482);
nand U5848 (N_5848,N_2062,N_3040);
nand U5849 (N_5849,N_2413,N_616);
nor U5850 (N_5850,N_3903,N_2982);
and U5851 (N_5851,N_2322,N_2349);
nor U5852 (N_5852,N_2981,N_4042);
or U5853 (N_5853,N_2146,N_2162);
or U5854 (N_5854,N_581,N_4534);
or U5855 (N_5855,N_3604,N_3436);
nand U5856 (N_5856,N_912,N_4923);
or U5857 (N_5857,N_4811,N_2220);
and U5858 (N_5858,N_2787,N_4275);
nand U5859 (N_5859,N_2396,N_1963);
nor U5860 (N_5860,N_1384,N_928);
nor U5861 (N_5861,N_1848,N_1465);
nand U5862 (N_5862,N_1245,N_4446);
or U5863 (N_5863,N_1025,N_2471);
and U5864 (N_5864,N_4793,N_594);
and U5865 (N_5865,N_4655,N_2881);
or U5866 (N_5866,N_995,N_156);
nor U5867 (N_5867,N_695,N_858);
nand U5868 (N_5868,N_4802,N_1330);
or U5869 (N_5869,N_655,N_1665);
nor U5870 (N_5870,N_1271,N_4919);
or U5871 (N_5871,N_4841,N_1515);
nand U5872 (N_5872,N_4866,N_2549);
or U5873 (N_5873,N_1822,N_4660);
and U5874 (N_5874,N_4480,N_2561);
or U5875 (N_5875,N_4669,N_3797);
nand U5876 (N_5876,N_159,N_4404);
nand U5877 (N_5877,N_298,N_246);
and U5878 (N_5878,N_4721,N_226);
and U5879 (N_5879,N_1648,N_4771);
or U5880 (N_5880,N_2769,N_1153);
nor U5881 (N_5881,N_2583,N_3844);
nand U5882 (N_5882,N_1412,N_3920);
nand U5883 (N_5883,N_4476,N_4299);
and U5884 (N_5884,N_917,N_169);
nor U5885 (N_5885,N_1541,N_2398);
nand U5886 (N_5886,N_932,N_3315);
and U5887 (N_5887,N_1144,N_182);
nor U5888 (N_5888,N_3532,N_3679);
or U5889 (N_5889,N_4686,N_1670);
nor U5890 (N_5890,N_3163,N_1700);
nor U5891 (N_5891,N_4823,N_1946);
nand U5892 (N_5892,N_4854,N_63);
nor U5893 (N_5893,N_1069,N_4213);
and U5894 (N_5894,N_2115,N_1073);
nor U5895 (N_5895,N_852,N_3323);
or U5896 (N_5896,N_2297,N_313);
and U5897 (N_5897,N_1973,N_2776);
nor U5898 (N_5898,N_4490,N_671);
or U5899 (N_5899,N_4519,N_3847);
nor U5900 (N_5900,N_1146,N_437);
or U5901 (N_5901,N_4790,N_2018);
nand U5902 (N_5902,N_1745,N_4065);
and U5903 (N_5903,N_2308,N_3468);
or U5904 (N_5904,N_4717,N_4652);
and U5905 (N_5905,N_539,N_1714);
and U5906 (N_5906,N_3299,N_930);
nand U5907 (N_5907,N_4413,N_1708);
nand U5908 (N_5908,N_1095,N_2598);
nand U5909 (N_5909,N_4220,N_4512);
or U5910 (N_5910,N_998,N_3985);
nor U5911 (N_5911,N_148,N_502);
and U5912 (N_5912,N_9,N_406);
nor U5913 (N_5913,N_595,N_96);
nor U5914 (N_5914,N_1993,N_312);
nand U5915 (N_5915,N_3465,N_4219);
or U5916 (N_5916,N_1243,N_70);
nand U5917 (N_5917,N_723,N_2832);
nor U5918 (N_5918,N_5,N_1532);
and U5919 (N_5919,N_4770,N_1779);
nand U5920 (N_5920,N_3464,N_1971);
and U5921 (N_5921,N_2733,N_277);
or U5922 (N_5922,N_4153,N_3639);
and U5923 (N_5923,N_1776,N_178);
nor U5924 (N_5924,N_2113,N_4518);
and U5925 (N_5925,N_522,N_3689);
nand U5926 (N_5926,N_3217,N_4238);
or U5927 (N_5927,N_2056,N_2179);
or U5928 (N_5928,N_3898,N_2517);
or U5929 (N_5929,N_4592,N_1254);
and U5930 (N_5930,N_2440,N_302);
and U5931 (N_5931,N_4662,N_4484);
xor U5932 (N_5932,N_4383,N_8);
nand U5933 (N_5933,N_330,N_3446);
nand U5934 (N_5934,N_218,N_2231);
and U5935 (N_5935,N_4241,N_2183);
and U5936 (N_5936,N_3306,N_3808);
and U5937 (N_5937,N_3796,N_2883);
xor U5938 (N_5938,N_2482,N_2748);
nand U5939 (N_5939,N_1359,N_3267);
nor U5940 (N_5940,N_3484,N_4468);
nand U5941 (N_5941,N_144,N_4688);
and U5942 (N_5942,N_3974,N_1456);
nand U5943 (N_5943,N_4349,N_1282);
nor U5944 (N_5944,N_2163,N_467);
nor U5945 (N_5945,N_4589,N_4041);
nor U5946 (N_5946,N_577,N_4178);
and U5947 (N_5947,N_3440,N_2002);
and U5948 (N_5948,N_3111,N_2965);
and U5949 (N_5949,N_3787,N_728);
or U5950 (N_5950,N_3220,N_4757);
or U5951 (N_5951,N_3241,N_4710);
nand U5952 (N_5952,N_4414,N_1206);
nand U5953 (N_5953,N_4621,N_1567);
nand U5954 (N_5954,N_3893,N_3697);
nand U5955 (N_5955,N_2484,N_2642);
nor U5956 (N_5956,N_3416,N_2145);
or U5957 (N_5957,N_2778,N_3881);
or U5958 (N_5958,N_2963,N_1495);
and U5959 (N_5959,N_469,N_951);
or U5960 (N_5960,N_366,N_400);
nand U5961 (N_5961,N_1443,N_4727);
and U5962 (N_5962,N_878,N_3618);
or U5963 (N_5963,N_3770,N_3357);
nor U5964 (N_5964,N_2110,N_1649);
and U5965 (N_5965,N_780,N_1644);
nor U5966 (N_5966,N_907,N_3919);
xor U5967 (N_5967,N_3539,N_1218);
and U5968 (N_5968,N_4593,N_4076);
or U5969 (N_5969,N_1181,N_1507);
nor U5970 (N_5970,N_4481,N_449);
or U5971 (N_5971,N_2829,N_2378);
or U5972 (N_5972,N_2333,N_486);
nand U5973 (N_5973,N_2997,N_497);
or U5974 (N_5974,N_4266,N_2882);
or U5975 (N_5975,N_4273,N_3559);
nand U5976 (N_5976,N_3006,N_834);
and U5977 (N_5977,N_1258,N_2824);
nand U5978 (N_5978,N_333,N_1984);
xnor U5979 (N_5979,N_1529,N_2804);
or U5980 (N_5980,N_2743,N_2797);
nand U5981 (N_5981,N_949,N_1952);
or U5982 (N_5982,N_1906,N_653);
nand U5983 (N_5983,N_1896,N_1301);
nand U5984 (N_5984,N_993,N_610);
and U5985 (N_5985,N_4005,N_4154);
or U5986 (N_5986,N_1559,N_4536);
nand U5987 (N_5987,N_3750,N_1389);
or U5988 (N_5988,N_242,N_1028);
nor U5989 (N_5989,N_1838,N_2499);
nand U5990 (N_5990,N_1717,N_4174);
nor U5991 (N_5991,N_94,N_2650);
and U5992 (N_5992,N_4640,N_2310);
and U5993 (N_5993,N_4445,N_2572);
or U5994 (N_5994,N_2334,N_41);
nand U5995 (N_5995,N_4856,N_3928);
or U5996 (N_5996,N_971,N_1335);
nand U5997 (N_5997,N_4001,N_4169);
or U5998 (N_5998,N_3915,N_1317);
and U5999 (N_5999,N_425,N_2946);
nand U6000 (N_6000,N_1149,N_4067);
nand U6001 (N_6001,N_555,N_2212);
nor U6002 (N_6002,N_939,N_2784);
nand U6003 (N_6003,N_1584,N_4417);
nand U6004 (N_6004,N_2971,N_1668);
nand U6005 (N_6005,N_4903,N_1249);
and U6006 (N_6006,N_287,N_886);
or U6007 (N_6007,N_2245,N_505);
and U6008 (N_6008,N_3910,N_4326);
and U6009 (N_6009,N_4375,N_1630);
or U6010 (N_6010,N_2261,N_3332);
nand U6011 (N_6011,N_4474,N_1380);
nand U6012 (N_6012,N_4586,N_677);
nand U6013 (N_6013,N_410,N_795);
or U6014 (N_6014,N_1805,N_2786);
nor U6015 (N_6015,N_1617,N_4943);
or U6016 (N_6016,N_4059,N_3874);
nand U6017 (N_6017,N_1589,N_657);
or U6018 (N_6018,N_4953,N_4032);
nor U6019 (N_6019,N_3533,N_3229);
or U6020 (N_6020,N_1614,N_687);
or U6021 (N_6021,N_1854,N_3022);
and U6022 (N_6022,N_3952,N_3635);
nor U6023 (N_6023,N_1041,N_634);
or U6024 (N_6024,N_4380,N_1978);
nor U6025 (N_6025,N_3995,N_174);
nand U6026 (N_6026,N_2792,N_4692);
and U6027 (N_6027,N_3523,N_3731);
or U6028 (N_6028,N_3190,N_1992);
or U6029 (N_6029,N_941,N_337);
or U6030 (N_6030,N_876,N_3511);
nand U6031 (N_6031,N_865,N_2958);
nor U6032 (N_6032,N_4964,N_3424);
and U6033 (N_6033,N_1197,N_3943);
nor U6034 (N_6034,N_4346,N_3727);
and U6035 (N_6035,N_2078,N_1726);
nor U6036 (N_6036,N_2211,N_1941);
and U6037 (N_6037,N_4449,N_2566);
nand U6038 (N_6038,N_1650,N_3577);
nand U6039 (N_6039,N_4424,N_1678);
and U6040 (N_6040,N_1348,N_167);
nand U6041 (N_6041,N_3827,N_4641);
or U6042 (N_6042,N_983,N_3378);
nand U6043 (N_6043,N_501,N_225);
nand U6044 (N_6044,N_4924,N_1677);
or U6045 (N_6045,N_3751,N_3799);
or U6046 (N_6046,N_418,N_1764);
or U6047 (N_6047,N_3557,N_4499);
nor U6048 (N_6048,N_281,N_880);
or U6049 (N_6049,N_2621,N_915);
or U6050 (N_6050,N_1289,N_1913);
and U6051 (N_6051,N_1673,N_3502);
and U6052 (N_6052,N_4294,N_3370);
xnor U6053 (N_6053,N_3448,N_4243);
or U6054 (N_6054,N_4168,N_1111);
nor U6055 (N_6055,N_4848,N_4165);
or U6056 (N_6056,N_4506,N_3970);
or U6057 (N_6057,N_3871,N_511);
nor U6058 (N_6058,N_2867,N_779);
and U6059 (N_6059,N_3337,N_243);
nor U6060 (N_6060,N_3481,N_2161);
nand U6061 (N_6061,N_7,N_4455);
or U6062 (N_6062,N_1801,N_3188);
and U6063 (N_6063,N_4085,N_3624);
xor U6064 (N_6064,N_541,N_4931);
or U6065 (N_6065,N_1736,N_2165);
nand U6066 (N_6066,N_2291,N_4159);
nand U6067 (N_6067,N_2770,N_3087);
or U6068 (N_6068,N_3428,N_1053);
nor U6069 (N_6069,N_4714,N_999);
and U6070 (N_6070,N_3113,N_1821);
or U6071 (N_6071,N_240,N_2749);
nand U6072 (N_6072,N_3665,N_2302);
or U6073 (N_6073,N_985,N_1381);
nor U6074 (N_6074,N_2920,N_832);
nor U6075 (N_6075,N_1851,N_260);
nor U6076 (N_6076,N_4628,N_3556);
nor U6077 (N_6077,N_507,N_766);
nand U6078 (N_6078,N_2513,N_2707);
nor U6079 (N_6079,N_4927,N_1294);
or U6080 (N_6080,N_452,N_1819);
and U6081 (N_6081,N_3977,N_4633);
nor U6082 (N_6082,N_4695,N_4426);
nor U6083 (N_6083,N_2685,N_4942);
nor U6084 (N_6084,N_2061,N_2022);
or U6085 (N_6085,N_2514,N_1201);
nand U6086 (N_6086,N_2702,N_4167);
nor U6087 (N_6087,N_4082,N_3521);
nor U6088 (N_6088,N_3387,N_1442);
nand U6089 (N_6089,N_4500,N_1663);
nor U6090 (N_6090,N_2580,N_4882);
and U6091 (N_6091,N_4447,N_1953);
nor U6092 (N_6092,N_968,N_1205);
nand U6093 (N_6093,N_2619,N_1780);
nand U6094 (N_6094,N_4237,N_2327);
nand U6095 (N_6095,N_1459,N_3672);
nand U6096 (N_6096,N_149,N_643);
or U6097 (N_6097,N_2252,N_4398);
nand U6098 (N_6098,N_3961,N_773);
nor U6099 (N_6099,N_2573,N_1855);
nand U6100 (N_6100,N_963,N_3677);
nand U6101 (N_6101,N_3998,N_3712);
or U6102 (N_6102,N_2594,N_2679);
and U6103 (N_6103,N_1080,N_2386);
nor U6104 (N_6104,N_4286,N_4899);
nor U6105 (N_6105,N_3197,N_448);
or U6106 (N_6106,N_4467,N_1755);
or U6107 (N_6107,N_1862,N_3095);
nand U6108 (N_6108,N_1716,N_2545);
nor U6109 (N_6109,N_1371,N_2460);
or U6110 (N_6110,N_3937,N_3932);
or U6111 (N_6111,N_822,N_315);
xnor U6112 (N_6112,N_4562,N_976);
and U6113 (N_6113,N_805,N_257);
and U6114 (N_6114,N_1893,N_4472);
or U6115 (N_6115,N_4330,N_2449);
nand U6116 (N_6116,N_1297,N_2351);
and U6117 (N_6117,N_3433,N_4822);
nor U6118 (N_6118,N_1664,N_1748);
and U6119 (N_6119,N_4751,N_168);
nand U6120 (N_6120,N_2041,N_2387);
nand U6121 (N_6121,N_2268,N_2669);
nand U6122 (N_6122,N_3374,N_4767);
and U6123 (N_6123,N_2203,N_2391);
nand U6124 (N_6124,N_564,N_355);
nand U6125 (N_6125,N_2321,N_1436);
nor U6126 (N_6126,N_3551,N_4867);
and U6127 (N_6127,N_3466,N_2403);
nand U6128 (N_6128,N_4658,N_4361);
and U6129 (N_6129,N_801,N_4775);
and U6130 (N_6130,N_2285,N_785);
and U6131 (N_6131,N_2741,N_4610);
or U6132 (N_6132,N_2164,N_3011);
or U6133 (N_6133,N_609,N_2737);
nand U6134 (N_6134,N_4681,N_496);
and U6135 (N_6135,N_2907,N_4635);
nor U6136 (N_6136,N_1769,N_1592);
or U6137 (N_6137,N_4471,N_1538);
and U6138 (N_6138,N_150,N_3764);
nor U6139 (N_6139,N_4030,N_191);
nor U6140 (N_6140,N_2170,N_4849);
and U6141 (N_6141,N_3801,N_4517);
xnor U6142 (N_6142,N_1874,N_4690);
nor U6143 (N_6143,N_4240,N_403);
nand U6144 (N_6144,N_3866,N_477);
and U6145 (N_6145,N_2636,N_4345);
and U6146 (N_6146,N_1256,N_1089);
nand U6147 (N_6147,N_3709,N_2564);
nor U6148 (N_6148,N_2441,N_1643);
nand U6149 (N_6149,N_4728,N_4936);
and U6150 (N_6150,N_1537,N_715);
nand U6151 (N_6151,N_40,N_4590);
nand U6152 (N_6152,N_2355,N_3973);
nand U6153 (N_6153,N_2225,N_3371);
or U6154 (N_6154,N_1524,N_229);
or U6155 (N_6155,N_1468,N_4630);
or U6156 (N_6156,N_1972,N_4905);
and U6157 (N_6157,N_2489,N_3128);
nand U6158 (N_6158,N_3544,N_902);
or U6159 (N_6159,N_4149,N_1549);
nand U6160 (N_6160,N_4025,N_3041);
or U6161 (N_6161,N_4998,N_4540);
nor U6162 (N_6162,N_3140,N_2190);
nand U6163 (N_6163,N_4653,N_2205);
nand U6164 (N_6164,N_3329,N_4694);
or U6165 (N_6165,N_1662,N_4493);
nor U6166 (N_6166,N_2808,N_3427);
or U6167 (N_6167,N_1713,N_4914);
xor U6168 (N_6168,N_4010,N_2970);
or U6169 (N_6169,N_2924,N_2821);
and U6170 (N_6170,N_2916,N_897);
or U6171 (N_6171,N_3470,N_986);
nor U6172 (N_6172,N_2994,N_2072);
or U6173 (N_6173,N_1273,N_4314);
and U6174 (N_6174,N_4935,N_4932);
and U6175 (N_6175,N_793,N_1774);
nor U6176 (N_6176,N_2698,N_618);
nand U6177 (N_6177,N_4548,N_4148);
or U6178 (N_6178,N_2674,N_4376);
nor U6179 (N_6179,N_992,N_4056);
and U6180 (N_6180,N_1394,N_2886);
nor U6181 (N_6181,N_4595,N_4411);
nor U6182 (N_6182,N_3819,N_1920);
and U6183 (N_6183,N_354,N_66);
nand U6184 (N_6184,N_938,N_888);
and U6185 (N_6185,N_2758,N_1597);
nand U6186 (N_6186,N_1945,N_15);
nor U6187 (N_6187,N_1065,N_1408);
or U6188 (N_6188,N_2094,N_786);
nor U6189 (N_6189,N_1839,N_1697);
or U6190 (N_6190,N_3252,N_2683);
nand U6191 (N_6191,N_4977,N_468);
nand U6192 (N_6192,N_4724,N_1827);
nor U6193 (N_6193,N_862,N_219);
nand U6194 (N_6194,N_4845,N_211);
nor U6195 (N_6195,N_379,N_3705);
and U6196 (N_6196,N_584,N_1721);
nand U6197 (N_6197,N_1501,N_4039);
nor U6198 (N_6198,N_2626,N_3993);
nor U6199 (N_6199,N_1114,N_2246);
nand U6200 (N_6200,N_1383,N_3430);
nand U6201 (N_6201,N_3314,N_4988);
nand U6202 (N_6202,N_1374,N_2515);
nor U6203 (N_6203,N_133,N_4313);
or U6204 (N_6204,N_2794,N_2560);
and U6205 (N_6205,N_2673,N_3457);
nor U6206 (N_6206,N_2617,N_1744);
or U6207 (N_6207,N_2602,N_2260);
nand U6208 (N_6208,N_987,N_3594);
or U6209 (N_6209,N_4123,N_4162);
nand U6210 (N_6210,N_1586,N_3056);
and U6211 (N_6211,N_4216,N_4978);
nor U6212 (N_6212,N_208,N_2501);
or U6213 (N_6213,N_3458,N_3062);
xnor U6214 (N_6214,N_4028,N_4960);
or U6215 (N_6215,N_4017,N_2589);
and U6216 (N_6216,N_3690,N_3860);
and U6217 (N_6217,N_4840,N_72);
and U6218 (N_6218,N_1688,N_2143);
or U6219 (N_6219,N_4870,N_3714);
and U6220 (N_6220,N_4009,N_1293);
xor U6221 (N_6221,N_2857,N_4094);
and U6222 (N_6222,N_3587,N_4300);
nor U6223 (N_6223,N_2635,N_472);
nor U6224 (N_6224,N_3780,N_924);
nor U6225 (N_6225,N_3642,N_622);
nor U6226 (N_6226,N_840,N_4520);
nor U6227 (N_6227,N_770,N_362);
or U6228 (N_6228,N_1189,N_1106);
nor U6229 (N_6229,N_3215,N_3612);
nand U6230 (N_6230,N_3829,N_1250);
nor U6231 (N_6231,N_2227,N_2217);
or U6232 (N_6232,N_1765,N_3493);
nand U6233 (N_6233,N_1621,N_1393);
nor U6234 (N_6234,N_1865,N_1344);
nand U6235 (N_6235,N_4874,N_1530);
nor U6236 (N_6236,N_598,N_12);
nand U6237 (N_6237,N_777,N_4552);
nand U6238 (N_6238,N_2877,N_602);
nor U6239 (N_6239,N_2263,N_4325);
nand U6240 (N_6240,N_3967,N_4836);
nor U6241 (N_6241,N_1440,N_2894);
and U6242 (N_6242,N_2228,N_3375);
xnor U6243 (N_6243,N_673,N_3068);
nor U6244 (N_6244,N_2026,N_1999);
nand U6245 (N_6245,N_2518,N_727);
or U6246 (N_6246,N_4348,N_4505);
and U6247 (N_6247,N_3354,N_4863);
nand U6248 (N_6248,N_3883,N_3175);
and U6249 (N_6249,N_4697,N_4303);
nand U6250 (N_6250,N_583,N_1097);
nor U6251 (N_6251,N_221,N_2419);
nor U6252 (N_6252,N_4535,N_1931);
nand U6253 (N_6253,N_3681,N_2987);
nand U6254 (N_6254,N_1613,N_2661);
and U6255 (N_6255,N_913,N_143);
or U6256 (N_6256,N_2136,N_3686);
or U6257 (N_6257,N_665,N_1291);
and U6258 (N_6258,N_4212,N_503);
nand U6259 (N_6259,N_3394,N_1568);
and U6260 (N_6260,N_3601,N_959);
or U6261 (N_6261,N_4453,N_3437);
and U6262 (N_6262,N_530,N_1618);
or U6263 (N_6263,N_33,N_787);
nor U6264 (N_6264,N_2950,N_2823);
or U6265 (N_6265,N_2546,N_970);
and U6266 (N_6266,N_2388,N_693);
nand U6267 (N_6267,N_4833,N_4929);
and U6268 (N_6268,N_1131,N_2025);
nor U6269 (N_6269,N_3761,N_128);
and U6270 (N_6270,N_3031,N_540);
nand U6271 (N_6271,N_1606,N_1624);
nor U6272 (N_6272,N_1277,N_2122);
xor U6273 (N_6273,N_2507,N_3777);
nand U6274 (N_6274,N_2309,N_919);
nor U6275 (N_6275,N_817,N_4588);
and U6276 (N_6276,N_3364,N_2953);
nand U6277 (N_6277,N_4293,N_1535);
and U6278 (N_6278,N_4704,N_2487);
nand U6279 (N_6279,N_3482,N_1026);
nor U6280 (N_6280,N_1782,N_376);
or U6281 (N_6281,N_4503,N_1489);
xor U6282 (N_6282,N_1735,N_4126);
and U6283 (N_6283,N_4659,N_1338);
or U6284 (N_6284,N_1554,N_2765);
nand U6285 (N_6285,N_1727,N_848);
nand U6286 (N_6286,N_3425,N_1240);
and U6287 (N_6287,N_249,N_4183);
nor U6288 (N_6288,N_336,N_3473);
nand U6289 (N_6289,N_2031,N_3395);
or U6290 (N_6290,N_1108,N_2000);
and U6291 (N_6291,N_2379,N_4196);
nor U6292 (N_6292,N_3811,N_4626);
and U6293 (N_6293,N_2257,N_4594);
nor U6294 (N_6294,N_2534,N_36);
nor U6295 (N_6295,N_3124,N_490);
and U6296 (N_6296,N_3034,N_1966);
or U6297 (N_6297,N_295,N_20);
nand U6298 (N_6298,N_2503,N_415);
nor U6299 (N_6299,N_4995,N_4342);
nor U6300 (N_6300,N_3562,N_996);
or U6301 (N_6301,N_4050,N_484);
or U6302 (N_6302,N_4970,N_1337);
or U6303 (N_6303,N_2223,N_826);
xnor U6304 (N_6304,N_1602,N_102);
nor U6305 (N_6305,N_3758,N_3046);
and U6306 (N_6306,N_2557,N_1079);
nand U6307 (N_6307,N_2796,N_1477);
and U6308 (N_6308,N_3313,N_1733);
or U6309 (N_6309,N_3084,N_429);
or U6310 (N_6310,N_1943,N_575);
or U6311 (N_6311,N_4817,N_1376);
and U6312 (N_6312,N_628,N_3896);
or U6313 (N_6313,N_4127,N_2033);
and U6314 (N_6314,N_363,N_1916);
nor U6315 (N_6315,N_509,N_4389);
or U6316 (N_6316,N_1228,N_4318);
nand U6317 (N_6317,N_3983,N_1857);
nand U6318 (N_6318,N_4402,N_4664);
nor U6319 (N_6319,N_578,N_908);
or U6320 (N_6320,N_2593,N_806);
xor U6321 (N_6321,N_1033,N_3782);
nand U6322 (N_6322,N_193,N_244);
or U6323 (N_6323,N_2905,N_2838);
or U6324 (N_6324,N_528,N_2973);
and U6325 (N_6325,N_417,N_2060);
nor U6326 (N_6326,N_4604,N_3129);
nor U6327 (N_6327,N_2006,N_81);
and U6328 (N_6328,N_2116,N_529);
and U6329 (N_6329,N_3412,N_23);
nand U6330 (N_6330,N_2592,N_2898);
and U6331 (N_6331,N_3079,N_391);
or U6332 (N_6332,N_2401,N_2490);
nand U6333 (N_6333,N_1305,N_1847);
nor U6334 (N_6334,N_2138,N_4425);
or U6335 (N_6335,N_1071,N_127);
nor U6336 (N_6336,N_1049,N_2262);
nor U6337 (N_6337,N_751,N_3627);
and U6338 (N_6338,N_765,N_1914);
and U6339 (N_6339,N_3824,N_1135);
and U6340 (N_6340,N_1752,N_1750);
and U6341 (N_6341,N_4713,N_3707);
nor U6342 (N_6342,N_4199,N_4442);
or U6343 (N_6343,N_292,N_432);
nor U6344 (N_6344,N_2361,N_1566);
nor U6345 (N_6345,N_2569,N_294);
and U6346 (N_6346,N_841,N_2581);
or U6347 (N_6347,N_489,N_2106);
or U6348 (N_6348,N_4915,N_514);
or U6349 (N_6349,N_2682,N_1099);
and U6350 (N_6350,N_2542,N_4844);
nand U6351 (N_6351,N_2102,N_4223);
or U6352 (N_6352,N_2584,N_772);
and U6353 (N_6353,N_76,N_2462);
and U6354 (N_6354,N_4784,N_3208);
nor U6355 (N_6355,N_380,N_2923);
nand U6356 (N_6356,N_3342,N_4385);
nand U6357 (N_6357,N_547,N_4197);
and U6358 (N_6358,N_3730,N_3684);
or U6359 (N_6359,N_3295,N_132);
nor U6360 (N_6360,N_3957,N_3277);
or U6361 (N_6361,N_4702,N_209);
nand U6362 (N_6362,N_3460,N_799);
and U6363 (N_6363,N_183,N_1129);
and U6364 (N_6364,N_4723,N_1734);
and U6365 (N_6365,N_735,N_319);
and U6366 (N_6366,N_1199,N_4105);
or U6367 (N_6367,N_4665,N_4818);
nand U6368 (N_6368,N_4989,N_3442);
and U6369 (N_6369,N_2125,N_2755);
nand U6370 (N_6370,N_214,N_77);
xor U6371 (N_6371,N_4486,N_4139);
or U6372 (N_6372,N_4451,N_4575);
or U6373 (N_6373,N_2539,N_1623);
nand U6374 (N_6374,N_446,N_3271);
nand U6375 (N_6375,N_2693,N_3102);
or U6376 (N_6376,N_1411,N_4516);
or U6377 (N_6377,N_1910,N_2839);
nor U6378 (N_6378,N_4066,N_4881);
nand U6379 (N_6379,N_2376,N_2);
nor U6380 (N_6380,N_3409,N_504);
nor U6381 (N_6381,N_3505,N_3118);
or U6382 (N_6382,N_4618,N_1724);
nor U6383 (N_6383,N_1171,N_4214);
nand U6384 (N_6384,N_1133,N_2209);
and U6385 (N_6385,N_2248,N_526);
or U6386 (N_6386,N_2893,N_342);
or U6387 (N_6387,N_3290,N_4715);
nor U6388 (N_6388,N_1148,N_4755);
nand U6389 (N_6389,N_4309,N_2502);
and U6390 (N_6390,N_1007,N_3591);
and U6391 (N_6391,N_1437,N_2842);
and U6392 (N_6392,N_2074,N_515);
and U6393 (N_6393,N_4629,N_2383);
nand U6394 (N_6394,N_3774,N_3099);
or U6395 (N_6395,N_3373,N_2544);
nand U6396 (N_6396,N_3785,N_1761);
nor U6397 (N_6397,N_4551,N_2496);
and U6398 (N_6398,N_60,N_1046);
nand U6399 (N_6399,N_1172,N_2068);
or U6400 (N_6400,N_4407,N_2834);
or U6401 (N_6401,N_1255,N_3287);
or U6402 (N_6402,N_562,N_3592);
nor U6403 (N_6403,N_1281,N_4006);
nand U6404 (N_6404,N_113,N_4945);
nor U6405 (N_6405,N_1130,N_1247);
nand U6406 (N_6406,N_3411,N_3453);
and U6407 (N_6407,N_3055,N_4444);
nor U6408 (N_6408,N_4289,N_4278);
nor U6409 (N_6409,N_3135,N_4805);
and U6410 (N_6410,N_744,N_3182);
or U6411 (N_6411,N_2402,N_1924);
and U6412 (N_6412,N_1772,N_2904);
and U6413 (N_6413,N_1102,N_4086);
xor U6414 (N_6414,N_234,N_2435);
or U6415 (N_6415,N_1540,N_3685);
and U6416 (N_6416,N_4381,N_2130);
and U6417 (N_6417,N_4037,N_4110);
or U6418 (N_6418,N_4386,N_3979);
or U6419 (N_6419,N_4435,N_1388);
nand U6420 (N_6420,N_1345,N_3858);
nor U6421 (N_6421,N_1361,N_4950);
xnor U6422 (N_6422,N_1352,N_1092);
and U6423 (N_6423,N_2571,N_3583);
nor U6424 (N_6424,N_1424,N_1803);
or U6425 (N_6425,N_4209,N_82);
and U6426 (N_6426,N_2732,N_216);
and U6427 (N_6427,N_659,N_2178);
and U6428 (N_6428,N_4720,N_4906);
nor U6429 (N_6429,N_3032,N_4441);
nor U6430 (N_6430,N_2336,N_2945);
nand U6431 (N_6431,N_3571,N_4574);
nand U6432 (N_6432,N_3749,N_4816);
nand U6433 (N_6433,N_3671,N_3590);
or U6434 (N_6434,N_35,N_720);
nand U6435 (N_6435,N_678,N_4057);
and U6436 (N_6436,N_1661,N_1226);
nor U6437 (N_6437,N_2604,N_4133);
and U6438 (N_6438,N_4129,N_3510);
and U6439 (N_6439,N_2238,N_3561);
or U6440 (N_6440,N_2719,N_4812);
nor U6441 (N_6441,N_2931,N_4358);
and U6442 (N_6442,N_129,N_2979);
or U6443 (N_6443,N_3752,N_4674);
nand U6444 (N_6444,N_2506,N_1496);
or U6445 (N_6445,N_2753,N_2552);
nand U6446 (N_6446,N_743,N_2255);
nand U6447 (N_6447,N_994,N_4344);
nand U6448 (N_6448,N_2417,N_4759);
nor U6449 (N_6449,N_2216,N_2595);
and U6450 (N_6450,N_1797,N_1021);
nor U6451 (N_6451,N_3623,N_4366);
nor U6452 (N_6452,N_1682,N_3396);
nor U6453 (N_6453,N_586,N_1013);
nor U6454 (N_6454,N_1591,N_2533);
or U6455 (N_6455,N_2638,N_2639);
nand U6456 (N_6456,N_620,N_4739);
xnor U6457 (N_6457,N_4430,N_2647);
nor U6458 (N_6458,N_3390,N_1284);
or U6459 (N_6459,N_1534,N_4181);
and U6460 (N_6460,N_2226,N_4699);
nand U6461 (N_6461,N_681,N_4638);
nor U6462 (N_6462,N_3495,N_1609);
nor U6463 (N_6463,N_1962,N_1954);
or U6464 (N_6464,N_2065,N_1209);
or U6465 (N_6465,N_1321,N_3589);
nor U6466 (N_6466,N_3013,N_2840);
or U6467 (N_6467,N_3452,N_4392);
and U6468 (N_6468,N_3127,N_830);
and U6469 (N_6469,N_2370,N_1326);
nand U6470 (N_6470,N_2659,N_3599);
and U6471 (N_6471,N_846,N_3047);
or U6472 (N_6472,N_3297,N_844);
nand U6473 (N_6473,N_202,N_3900);
nand U6474 (N_6474,N_2277,N_29);
or U6475 (N_6475,N_868,N_4473);
nor U6476 (N_6476,N_1581,N_2605);
nor U6477 (N_6477,N_414,N_3648);
nor U6478 (N_6478,N_2445,N_1246);
or U6479 (N_6479,N_2612,N_2207);
nand U6480 (N_6480,N_3406,N_3852);
xnor U6481 (N_6481,N_1450,N_3812);
nor U6482 (N_6482,N_4891,N_3747);
nor U6483 (N_6483,N_1076,N_3226);
and U6484 (N_6484,N_1016,N_2287);
and U6485 (N_6485,N_2672,N_2088);
and U6486 (N_6486,N_177,N_3231);
nand U6487 (N_6487,N_491,N_1161);
or U6488 (N_6488,N_1683,N_2833);
or U6489 (N_6489,N_2418,N_1785);
and U6490 (N_6490,N_78,N_1646);
nand U6491 (N_6491,N_2455,N_3007);
nor U6492 (N_6492,N_3057,N_3676);
and U6493 (N_6493,N_1179,N_2662);
or U6494 (N_6494,N_2479,N_3211);
or U6495 (N_6495,N_1022,N_2236);
and U6496 (N_6496,N_471,N_725);
nor U6497 (N_6497,N_2049,N_4357);
and U6498 (N_6498,N_1186,N_875);
or U6499 (N_6499,N_2760,N_2457);
and U6500 (N_6500,N_2952,N_815);
and U6501 (N_6501,N_4200,N_4600);
and U6502 (N_6502,N_617,N_2280);
and U6503 (N_6503,N_4815,N_4634);
nor U6504 (N_6504,N_11,N_1227);
nor U6505 (N_6505,N_3641,N_2806);
nand U6506 (N_6506,N_2428,N_3912);
and U6507 (N_6507,N_1969,N_4320);
nor U6508 (N_6508,N_4773,N_784);
or U6509 (N_6509,N_2495,N_2275);
nand U6510 (N_6510,N_1045,N_1003);
and U6511 (N_6511,N_929,N_1576);
nand U6512 (N_6512,N_4071,N_684);
nor U6513 (N_6513,N_4222,N_732);
nor U6514 (N_6514,N_4643,N_4996);
nand U6515 (N_6515,N_4749,N_500);
and U6516 (N_6516,N_664,N_470);
or U6517 (N_6517,N_3651,N_1574);
and U6518 (N_6518,N_18,N_2188);
or U6519 (N_6519,N_2253,N_1002);
or U6520 (N_6520,N_3867,N_4034);
and U6521 (N_6521,N_651,N_421);
or U6522 (N_6522,N_769,N_304);
nand U6523 (N_6523,N_4719,N_2939);
nor U6524 (N_6524,N_1008,N_3688);
and U6525 (N_6525,N_3471,N_4607);
and U6526 (N_6526,N_37,N_3563);
xor U6527 (N_6527,N_3341,N_4290);
or U6528 (N_6528,N_3377,N_574);
nor U6529 (N_6529,N_3255,N_3245);
and U6530 (N_6530,N_982,N_1808);
nor U6531 (N_6531,N_582,N_3889);
xnor U6532 (N_6532,N_1274,N_3520);
or U6533 (N_6533,N_4131,N_1788);
xnor U6534 (N_6534,N_1005,N_42);
nand U6535 (N_6535,N_1029,N_4930);
and U6536 (N_6536,N_1706,N_4608);
nor U6537 (N_6537,N_3232,N_4164);
or U6538 (N_6538,N_1196,N_3151);
nor U6539 (N_6539,N_2728,N_1506);
and U6540 (N_6540,N_2756,N_1877);
and U6541 (N_6541,N_3634,N_4796);
and U6542 (N_6542,N_2888,N_179);
or U6543 (N_6543,N_2112,N_1841);
and U6544 (N_6544,N_4311,N_3793);
nand U6545 (N_6545,N_2101,N_1269);
or U6546 (N_6546,N_2293,N_3285);
nor U6547 (N_6547,N_280,N_4317);
nand U6548 (N_6548,N_2254,N_2992);
or U6549 (N_6549,N_1454,N_407);
and U6550 (N_6550,N_931,N_67);
nand U6551 (N_6551,N_299,N_3933);
nand U6552 (N_6552,N_3039,N_4880);
or U6553 (N_6553,N_4249,N_3195);
nand U6554 (N_6554,N_2036,N_1001);
nand U6555 (N_6555,N_4758,N_2114);
nand U6556 (N_6556,N_2218,N_458);
nand U6557 (N_6557,N_2198,N_3633);
nand U6558 (N_6558,N_2734,N_4696);
or U6559 (N_6559,N_1229,N_3512);
and U6560 (N_6560,N_2836,N_2706);
nand U6561 (N_6561,N_495,N_600);
nor U6562 (N_6562,N_2360,N_2699);
or U6563 (N_6563,N_264,N_3971);
nor U6564 (N_6564,N_739,N_4585);
xnor U6565 (N_6565,N_1353,N_1187);
xnor U6566 (N_6566,N_2174,N_3348);
nor U6567 (N_6567,N_3090,N_2284);
nand U6568 (N_6568,N_1881,N_3663);
nand U6569 (N_6569,N_192,N_1252);
nand U6570 (N_6570,N_2961,N_2845);
nor U6571 (N_6571,N_1513,N_111);
nor U6572 (N_6572,N_163,N_3855);
and U6573 (N_6573,N_534,N_3925);
nor U6574 (N_6574,N_2739,N_4339);
nand U6575 (N_6575,N_368,N_3897);
nor U6576 (N_6576,N_1446,N_1157);
or U6577 (N_6577,N_3736,N_724);
xor U6578 (N_6578,N_623,N_4173);
nor U6579 (N_6579,N_3660,N_636);
nor U6580 (N_6580,N_3949,N_1096);
and U6581 (N_6581,N_4742,N_4897);
or U6582 (N_6582,N_2117,N_52);
and U6583 (N_6583,N_2901,N_2438);
nand U6584 (N_6584,N_3000,N_4969);
nor U6585 (N_6585,N_1313,N_3784);
and U6586 (N_6586,N_2126,N_3024);
or U6587 (N_6587,N_3125,N_3576);
or U6588 (N_6588,N_4510,N_4044);
nand U6589 (N_6589,N_2204,N_2729);
and U6590 (N_6590,N_4457,N_2320);
nor U6591 (N_6591,N_2470,N_4612);
or U6592 (N_6592,N_1478,N_4678);
nand U6593 (N_6593,N_3439,N_85);
and U6594 (N_6594,N_2464,N_4198);
or U6595 (N_6595,N_173,N_812);
nand U6596 (N_6596,N_1024,N_405);
nor U6597 (N_6597,N_1552,N_4916);
nand U6598 (N_6598,N_3052,N_3365);
nor U6599 (N_6599,N_2538,N_2433);
or U6600 (N_6600,N_2913,N_4577);
and U6601 (N_6601,N_647,N_1522);
nand U6602 (N_6602,N_305,N_3786);
nand U6603 (N_6603,N_4284,N_1656);
nor U6604 (N_6604,N_4875,N_3951);
nor U6605 (N_6605,N_1595,N_1901);
and U6606 (N_6606,N_2844,N_1429);
nand U6607 (N_6607,N_4809,N_1872);
and U6608 (N_6608,N_3479,N_2798);
nor U6609 (N_6609,N_4054,N_1267);
and U6610 (N_6610,N_4537,N_3567);
and U6611 (N_6611,N_2512,N_3122);
nor U6612 (N_6612,N_1902,N_4807);
or U6613 (N_6613,N_423,N_3018);
or U6614 (N_6614,N_3894,N_2686);
or U6615 (N_6615,N_2895,N_3745);
and U6616 (N_6616,N_1467,N_4682);
nand U6617 (N_6617,N_1521,N_606);
nand U6618 (N_6618,N_2432,N_4179);
and U6619 (N_6619,N_4649,N_3619);
and U6620 (N_6620,N_3934,N_1299);
nor U6621 (N_6621,N_1164,N_2711);
or U6622 (N_6622,N_3652,N_1);
xnor U6623 (N_6623,N_2481,N_4879);
nor U6624 (N_6624,N_390,N_1520);
and U6625 (N_6625,N_2736,N_1691);
nor U6626 (N_6626,N_756,N_1109);
nor U6627 (N_6627,N_2652,N_4465);
nor U6628 (N_6628,N_1462,N_950);
or U6629 (N_6629,N_4141,N_2954);
or U6630 (N_6630,N_3281,N_3775);
nand U6631 (N_6631,N_1059,N_198);
nor U6632 (N_6632,N_2900,N_1391);
nor U6633 (N_6633,N_450,N_262);
or U6634 (N_6634,N_4821,N_1375);
and U6635 (N_6635,N_4569,N_1000);
and U6636 (N_6636,N_3352,N_2775);
nor U6637 (N_6637,N_1402,N_4485);
nor U6638 (N_6638,N_137,N_1127);
or U6639 (N_6639,N_4625,N_2633);
and U6640 (N_6640,N_3148,N_1571);
or U6641 (N_6641,N_1612,N_4189);
or U6642 (N_6642,N_3293,N_4675);
or U6643 (N_6643,N_365,N_2887);
nand U6644 (N_6644,N_158,N_4);
and U6645 (N_6645,N_4308,N_2208);
nand U6646 (N_6646,N_3421,N_2726);
nor U6647 (N_6647,N_1253,N_4786);
nand U6648 (N_6648,N_4718,N_3929);
or U6649 (N_6649,N_2703,N_4117);
or U6650 (N_6650,N_1833,N_1487);
or U6651 (N_6651,N_1367,N_2027);
and U6652 (N_6652,N_3210,N_798);
nand U6653 (N_6653,N_1027,N_4698);
or U6654 (N_6654,N_4135,N_4205);
and U6655 (N_6655,N_3236,N_4301);
or U6656 (N_6656,N_1238,N_4984);
or U6657 (N_6657,N_1844,N_1339);
nand U6658 (N_6658,N_1233,N_4703);
nand U6659 (N_6659,N_435,N_3276);
nand U6660 (N_6660,N_4231,N_1354);
nand U6661 (N_6661,N_4952,N_662);
nor U6662 (N_6662,N_824,N_2147);
nand U6663 (N_6663,N_3498,N_357);
and U6664 (N_6664,N_58,N_4666);
nor U6665 (N_6665,N_498,N_3807);
nor U6666 (N_6666,N_2611,N_2630);
nand U6667 (N_6667,N_2109,N_2300);
and U6668 (N_6668,N_1473,N_3762);
nor U6669 (N_6669,N_2957,N_1791);
and U6670 (N_6670,N_1453,N_741);
or U6671 (N_6671,N_3813,N_103);
xor U6672 (N_6672,N_1410,N_2290);
nor U6673 (N_6673,N_4312,N_4295);
xor U6674 (N_6674,N_2289,N_2044);
or U6675 (N_6675,N_4077,N_1760);
and U6676 (N_6676,N_1853,N_3916);
and U6677 (N_6677,N_1287,N_394);
nor U6678 (N_6678,N_2731,N_2853);
nand U6679 (N_6679,N_1888,N_2641);
nor U6680 (N_6680,N_1809,N_343);
and U6681 (N_6681,N_512,N_1975);
nand U6682 (N_6682,N_3038,N_2864);
and U6683 (N_6683,N_3422,N_372);
nor U6684 (N_6684,N_3094,N_3996);
nor U6685 (N_6685,N_1451,N_811);
and U6686 (N_6686,N_2866,N_3266);
nand U6687 (N_6687,N_1034,N_3161);
xor U6688 (N_6688,N_2764,N_1645);
and U6689 (N_6689,N_141,N_2491);
and U6690 (N_6690,N_2523,N_1948);
nand U6691 (N_6691,N_764,N_4053);
or U6692 (N_6692,N_2632,N_4934);
nand U6693 (N_6693,N_4248,N_385);
nor U6694 (N_6694,N_4100,N_1270);
or U6695 (N_6695,N_166,N_2623);
nor U6696 (N_6696,N_53,N_3878);
nor U6697 (N_6697,N_4297,N_3739);
nand U6698 (N_6698,N_1997,N_708);
and U6699 (N_6699,N_960,N_1653);
nor U6700 (N_6700,N_632,N_2414);
or U6701 (N_6701,N_573,N_3636);
nand U6702 (N_6702,N_1921,N_3381);
nor U6703 (N_6703,N_4019,N_3256);
or U6704 (N_6704,N_3631,N_3026);
nor U6705 (N_6705,N_2788,N_4460);
and U6706 (N_6706,N_4580,N_3429);
nor U6707 (N_6707,N_2783,N_4494);
or U6708 (N_6708,N_4023,N_1846);
and U6709 (N_6709,N_1709,N_2614);
or U6710 (N_6710,N_1811,N_100);
and U6711 (N_6711,N_340,N_2430);
or U6712 (N_6712,N_1965,N_2789);
nand U6713 (N_6713,N_401,N_1680);
or U6714 (N_6714,N_607,N_2335);
or U6715 (N_6715,N_4835,N_3112);
nor U6716 (N_6716,N_462,N_3243);
or U6717 (N_6717,N_1230,N_718);
nor U6718 (N_6718,N_393,N_4502);
nor U6719 (N_6719,N_2079,N_3972);
or U6720 (N_6720,N_4954,N_4972);
nand U6721 (N_6721,N_2149,N_3492);
and U6722 (N_6722,N_2927,N_698);
or U6723 (N_6723,N_2962,N_272);
nand U6724 (N_6724,N_3253,N_601);
nor U6725 (N_6725,N_3907,N_936);
nor U6726 (N_6726,N_4819,N_2929);
and U6727 (N_6727,N_3535,N_3887);
nand U6728 (N_6728,N_189,N_2671);
nor U6729 (N_6729,N_3391,N_339);
and U6730 (N_6730,N_3558,N_2959);
nand U6731 (N_6731,N_864,N_3404);
and U6732 (N_6732,N_4093,N_4416);
nor U6733 (N_6733,N_3963,N_1035);
nor U6734 (N_6734,N_4088,N_510);
nand U6735 (N_6735,N_2799,N_1563);
or U6736 (N_6736,N_1587,N_854);
nor U6737 (N_6737,N_3010,N_1958);
nor U6738 (N_6738,N_4458,N_1994);
or U6739 (N_6739,N_2375,N_1234);
or U6740 (N_6740,N_4158,N_4160);
or U6741 (N_6741,N_3723,N_1655);
or U6742 (N_6742,N_3272,N_4581);
and U6743 (N_6743,N_1043,N_3405);
nor U6744 (N_6744,N_604,N_1152);
and U6745 (N_6745,N_4976,N_1823);
and U6746 (N_6746,N_1486,N_3459);
and U6747 (N_6747,N_1379,N_4579);
nor U6748 (N_6748,N_4074,N_4837);
xnor U6749 (N_6749,N_2906,N_4679);
and U6750 (N_6750,N_1596,N_98);
and U6751 (N_6751,N_2266,N_2802);
nor U6752 (N_6752,N_4566,N_2213);
nor U6753 (N_6753,N_1835,N_1715);
or U6754 (N_6754,N_1704,N_3361);
nor U6755 (N_6755,N_3456,N_855);
or U6756 (N_6756,N_478,N_26);
nand U6757 (N_6757,N_2851,N_3092);
or U6758 (N_6758,N_3322,N_1960);
and U6759 (N_6759,N_3913,N_4922);
nor U6760 (N_6760,N_1642,N_1640);
nand U6761 (N_6761,N_2813,N_3550);
nor U6762 (N_6762,N_1232,N_1047);
and U6763 (N_6763,N_1288,N_2863);
nor U6764 (N_6764,N_1542,N_4746);
and U6765 (N_6765,N_4400,N_2032);
xnor U6766 (N_6766,N_2805,N_3940);
or U6767 (N_6767,N_3224,N_554);
or U6768 (N_6768,N_3347,N_3809);
xor U6769 (N_6769,N_274,N_4035);
nand U6770 (N_6770,N_2879,N_195);
and U6771 (N_6771,N_1599,N_331);
and U6772 (N_6772,N_4949,N_4367);
nor U6773 (N_6773,N_4268,N_4994);
or U6774 (N_6774,N_2949,N_2678);
or U6775 (N_6775,N_1695,N_1925);
nor U6776 (N_6776,N_1605,N_2096);
or U6777 (N_6777,N_1918,N_2762);
nor U6778 (N_6778,N_536,N_399);
nor U6779 (N_6779,N_215,N_1349);
and U6780 (N_6780,N_1800,N_4810);
or U6781 (N_6781,N_2415,N_2876);
or U6782 (N_6782,N_4798,N_1919);
or U6783 (N_6783,N_4475,N_1307);
nor U6784 (N_6784,N_896,N_4269);
nor U6785 (N_6785,N_2384,N_2010);
nor U6786 (N_6786,N_4185,N_3923);
or U6787 (N_6787,N_3921,N_2328);
nand U6788 (N_6788,N_228,N_4112);
nor U6789 (N_6789,N_4572,N_387);
or U6790 (N_6790,N_4672,N_325);
nand U6791 (N_6791,N_1938,N_4887);
nor U6792 (N_6792,N_1470,N_645);
or U6793 (N_6793,N_884,N_3822);
and U6794 (N_6794,N_3321,N_1870);
or U6795 (N_6795,N_2649,N_2347);
nor U6796 (N_6796,N_3768,N_1929);
or U6797 (N_6797,N_4438,N_4489);
or U6798 (N_6798,N_3076,N_3564);
xor U6799 (N_6799,N_4889,N_2118);
and U6800 (N_6800,N_2759,N_2771);
nand U6801 (N_6801,N_4613,N_1369);
or U6802 (N_6802,N_1536,N_250);
and U6803 (N_6803,N_3513,N_4351);
nand U6804 (N_6804,N_1611,N_1156);
nand U6805 (N_6805,N_3938,N_220);
nor U6806 (N_6806,N_642,N_1892);
nand U6807 (N_6807,N_2299,N_3962);
or U6808 (N_6808,N_4965,N_901);
nor U6809 (N_6809,N_1401,N_1039);
and U6810 (N_6810,N_2861,N_3890);
nand U6811 (N_6811,N_1490,N_1009);
nor U6812 (N_6812,N_1502,N_1891);
nand U6813 (N_6813,N_188,N_251);
or U6814 (N_6814,N_737,N_563);
or U6815 (N_6815,N_2042,N_4431);
nand U6816 (N_6816,N_4130,N_3265);
nor U6817 (N_6817,N_1060,N_2664);
and U6818 (N_6818,N_371,N_1483);
or U6819 (N_6819,N_4904,N_1516);
and U6820 (N_6820,N_4022,N_4370);
or U6821 (N_6821,N_3218,N_4862);
nand U6822 (N_6822,N_3214,N_121);
or U6823 (N_6823,N_3965,N_2903);
and U6824 (N_6824,N_1414,N_629);
nand U6825 (N_6825,N_3462,N_3555);
nor U6826 (N_6826,N_2940,N_843);
and U6827 (N_6827,N_4726,N_2527);
and U6828 (N_6828,N_2872,N_621);
and U6829 (N_6829,N_2431,N_857);
nor U6830 (N_6830,N_4021,N_3014);
nor U6831 (N_6831,N_374,N_3154);
nand U6832 (N_6832,N_4353,N_2131);
or U6833 (N_6833,N_4307,N_4283);
nor U6834 (N_6834,N_130,N_1793);
and U6835 (N_6835,N_4762,N_2477);
or U6836 (N_6836,N_4983,N_259);
nor U6837 (N_6837,N_2995,N_3081);
nor U6838 (N_6838,N_2059,N_3008);
and U6839 (N_6839,N_4885,N_4993);
nor U6840 (N_6840,N_2028,N_4170);
and U6841 (N_6841,N_927,N_4316);
or U6842 (N_6842,N_2450,N_4211);
nand U6843 (N_6843,N_4280,N_1426);
or U6844 (N_6844,N_3121,N_1159);
nand U6845 (N_6845,N_258,N_1285);
nor U6846 (N_6846,N_3754,N_3116);
xnor U6847 (N_6847,N_4852,N_2070);
nor U6848 (N_6848,N_3687,N_2525);
or U6849 (N_6849,N_1441,N_3702);
and U6850 (N_6850,N_3192,N_3461);
nor U6851 (N_6851,N_3259,N_3106);
or U6852 (N_6852,N_2865,N_2723);
nor U6853 (N_6853,N_543,N_14);
and U6854 (N_6854,N_187,N_1732);
and U6855 (N_6855,N_2935,N_1085);
and U6856 (N_6856,N_3100,N_558);
nand U6857 (N_6857,N_4636,N_1118);
nor U6858 (N_6858,N_3522,N_2412);
nor U6859 (N_6859,N_1279,N_3131);
or U6860 (N_6860,N_3065,N_2429);
or U6861 (N_6861,N_2091,N_4877);
nor U6862 (N_6862,N_2405,N_4106);
and U6863 (N_6863,N_4764,N_3803);
or U6864 (N_6864,N_124,N_2859);
or U6865 (N_6865,N_1976,N_1601);
or U6866 (N_6866,N_3418,N_1382);
and U6867 (N_6867,N_4888,N_370);
nor U6868 (N_6868,N_1657,N_3984);
and U6869 (N_6869,N_3444,N_2486);
nand U6870 (N_6870,N_803,N_871);
nor U6871 (N_6871,N_626,N_719);
nand U6872 (N_6872,N_3501,N_1970);
and U6873 (N_6873,N_3474,N_4310);
nor U6874 (N_6874,N_2700,N_344);
or U6875 (N_6875,N_288,N_1332);
and U6876 (N_6876,N_2055,N_2522);
or U6877 (N_6877,N_2155,N_83);
nand U6878 (N_6878,N_3763,N_2132);
nor U6879 (N_6879,N_2326,N_308);
nor U6880 (N_6880,N_1165,N_4051);
xnor U6881 (N_6881,N_833,N_3721);
and U6882 (N_6882,N_2932,N_2304);
nor U6883 (N_6883,N_276,N_1804);
nand U6884 (N_6884,N_3674,N_2766);
nand U6885 (N_6885,N_2526,N_1484);
and U6886 (N_6886,N_2119,N_4171);
nand U6887 (N_6887,N_2912,N_4846);
nor U6888 (N_6888,N_2283,N_2980);
and U6889 (N_6889,N_3292,N_895);
nand U6890 (N_6890,N_2014,N_3673);
nand U6891 (N_6891,N_3327,N_2083);
nor U6892 (N_6892,N_4748,N_3579);
nand U6893 (N_6893,N_4382,N_1460);
and U6894 (N_6894,N_1651,N_921);
and U6895 (N_6895,N_2918,N_969);
nor U6896 (N_6896,N_1917,N_441);
or U6897 (N_6897,N_3369,N_4563);
xnor U6898 (N_6898,N_4627,N_389);
or U6899 (N_6899,N_92,N_3955);
nor U6900 (N_6900,N_2281,N_2374);
nand U6901 (N_6901,N_2030,N_4554);
and U6902 (N_6902,N_4689,N_2377);
nor U6903 (N_6903,N_1758,N_2891);
or U6904 (N_6904,N_4470,N_4834);
or U6905 (N_6905,N_2447,N_3888);
and U6906 (N_6906,N_3696,N_2185);
nand U6907 (N_6907,N_3490,N_2103);
nand U6908 (N_6908,N_3067,N_1932);
or U6909 (N_6909,N_1825,N_4260);
and U6910 (N_6910,N_1500,N_2176);
and U6911 (N_6911,N_4264,N_3423);
or U6912 (N_6912,N_3449,N_443);
nor U6913 (N_6913,N_3647,N_4576);
or U6914 (N_6914,N_10,N_1280);
nor U6915 (N_6915,N_3097,N_1850);
or U6916 (N_6916,N_4399,N_3117);
and U6917 (N_6917,N_916,N_676);
nand U6918 (N_6918,N_3876,N_2519);
nor U6919 (N_6919,N_2038,N_587);
nand U6920 (N_6920,N_1257,N_358);
and U6921 (N_6921,N_1543,N_1738);
or U6922 (N_6922,N_2352,N_1066);
or U6923 (N_6923,N_2359,N_4895);
and U6924 (N_6924,N_3948,N_3656);
and U6925 (N_6925,N_1011,N_767);
nand U6926 (N_6926,N_1463,N_4144);
xnor U6927 (N_6927,N_2249,N_3185);
nand U6928 (N_6928,N_227,N_3978);
and U6929 (N_6929,N_637,N_3003);
nor U6930 (N_6930,N_2493,N_1950);
and U6931 (N_6931,N_4992,N_3735);
and U6932 (N_6932,N_652,N_3379);
nor U6933 (N_6933,N_781,N_2848);
nor U6934 (N_6934,N_1123,N_1223);
nand U6935 (N_6935,N_2715,N_3946);
or U6936 (N_6936,N_3861,N_4533);
nand U6937 (N_6937,N_3917,N_2311);
nor U6938 (N_6938,N_3870,N_3415);
nand U6939 (N_6939,N_3414,N_2423);
nor U6940 (N_6940,N_1042,N_1077);
nor U6941 (N_6941,N_1420,N_2399);
nand U6942 (N_6942,N_4528,N_4832);
nor U6943 (N_6943,N_4104,N_2554);
or U6944 (N_6944,N_4292,N_670);
xnor U6945 (N_6945,N_4729,N_1216);
nand U6946 (N_6946,N_1169,N_1798);
nor U6947 (N_6947,N_3164,N_686);
nand U6948 (N_6948,N_3857,N_2843);
nor U6949 (N_6949,N_118,N_2086);
and U6950 (N_6950,N_3172,N_2722);
or U6951 (N_6951,N_442,N_853);
or U6952 (N_6952,N_3568,N_3939);
and U6953 (N_6953,N_54,N_1037);
nor U6954 (N_6954,N_850,N_2016);
nor U6955 (N_6955,N_4483,N_3527);
and U6956 (N_6956,N_3443,N_3659);
nand U6957 (N_6957,N_404,N_3228);
and U6958 (N_6958,N_4750,N_4151);
or U6959 (N_6959,N_909,N_2768);
or U6960 (N_6960,N_3719,N_4513);
and U6961 (N_6961,N_2587,N_203);
nor U6962 (N_6962,N_4966,N_4215);
nor U6963 (N_6963,N_206,N_4043);
or U6964 (N_6964,N_3250,N_2618);
nand U6965 (N_6965,N_3009,N_656);
or U6966 (N_6966,N_2451,N_3999);
or U6967 (N_6967,N_2579,N_1207);
nor U6968 (N_6968,N_4463,N_3141);
or U6969 (N_6969,N_4744,N_4990);
or U6970 (N_6970,N_3783,N_2921);
or U6971 (N_6971,N_359,N_3835);
nor U6972 (N_6972,N_4109,N_1220);
nand U6973 (N_6973,N_3905,N_1771);
nor U6974 (N_6974,N_4422,N_4121);
nor U6975 (N_6975,N_2043,N_981);
and U6976 (N_6976,N_4491,N_2411);
and U6977 (N_6977,N_2337,N_2013);
and U6978 (N_6978,N_1731,N_2615);
nor U6979 (N_6979,N_3082,N_4620);
nand U6980 (N_6980,N_1390,N_2873);
or U6981 (N_6981,N_1795,N_1968);
and U6982 (N_6982,N_2015,N_4233);
xnor U6983 (N_6983,N_3622,N_4452);
nor U6984 (N_6984,N_84,N_1607);
nor U6985 (N_6985,N_1082,N_230);
and U6986 (N_6986,N_2969,N_4785);
and U6987 (N_6987,N_2676,N_991);
and U6988 (N_6988,N_4073,N_3157);
nand U6989 (N_6989,N_34,N_311);
or U6990 (N_6990,N_984,N_465);
nand U6991 (N_6991,N_1202,N_1759);
and U6992 (N_6992,N_3790,N_2169);
or U6993 (N_6993,N_1124,N_2063);
or U6994 (N_6994,N_2687,N_2680);
nand U6995 (N_6995,N_889,N_3358);
nand U6996 (N_6996,N_646,N_2556);
nand U6997 (N_6997,N_3043,N_4761);
nor U6998 (N_6998,N_4305,N_2350);
and U6999 (N_6999,N_2325,N_740);
nor U7000 (N_7000,N_1177,N_4252);
and U7001 (N_7001,N_481,N_3499);
and U7002 (N_7002,N_4406,N_851);
or U7003 (N_7003,N_2089,N_3868);
or U7004 (N_7004,N_4530,N_416);
xnor U7005 (N_7005,N_1236,N_3291);
and U7006 (N_7006,N_161,N_700);
nor U7007 (N_7007,N_1355,N_332);
or U7008 (N_7008,N_3826,N_3042);
and U7009 (N_7009,N_4208,N_4623);
nand U7010 (N_7010,N_1188,N_1343);
nand U7011 (N_7011,N_644,N_730);
or U7012 (N_7012,N_4830,N_590);
and U7013 (N_7013,N_962,N_1278);
nand U7014 (N_7014,N_64,N_3107);
or U7015 (N_7015,N_494,N_2822);
or U7016 (N_7016,N_3744,N_4901);
and U7017 (N_7017,N_2319,N_3640);
nand U7018 (N_7018,N_3944,N_1272);
nor U7019 (N_7019,N_4354,N_4323);
nand U7020 (N_7020,N_2582,N_388);
nor U7021 (N_7021,N_2269,N_1783);
nand U7022 (N_7022,N_829,N_1100);
nand U7023 (N_7023,N_1897,N_4333);
nor U7024 (N_7024,N_682,N_3607);
nor U7025 (N_7025,N_1720,N_1061);
and U7026 (N_7026,N_499,N_4052);
and U7027 (N_7027,N_3325,N_197);
or U7028 (N_7028,N_482,N_2286);
or U7029 (N_7029,N_1377,N_324);
nand U7030 (N_7030,N_2278,N_3355);
and U7031 (N_7031,N_3028,N_516);
nand U7032 (N_7032,N_4469,N_3960);
or U7033 (N_7033,N_4864,N_820);
nand U7034 (N_7034,N_3085,N_3683);
nand U7035 (N_7035,N_3036,N_3372);
nand U7036 (N_7036,N_4797,N_329);
nor U7037 (N_7037,N_2585,N_3166);
or U7038 (N_7038,N_755,N_4327);
and U7039 (N_7039,N_4501,N_3130);
and U7040 (N_7040,N_1432,N_4256);
and U7041 (N_7041,N_145,N_2508);
and U7042 (N_7042,N_3037,N_4224);
xnor U7043 (N_7043,N_1160,N_4015);
xor U7044 (N_7044,N_61,N_1753);
or U7045 (N_7045,N_1859,N_4498);
nor U7046 (N_7046,N_633,N_680);
and U7047 (N_7047,N_2688,N_3994);
nand U7048 (N_7048,N_1861,N_1395);
and U7049 (N_7049,N_4436,N_4075);
nor U7050 (N_7050,N_2492,N_1195);
nor U7051 (N_7051,N_1398,N_3356);
or U7052 (N_7052,N_538,N_2069);
nand U7053 (N_7053,N_4259,N_1964);
nand U7054 (N_7054,N_1422,N_954);
nand U7055 (N_7055,N_2206,N_2716);
or U7056 (N_7056,N_1525,N_3235);
or U7057 (N_7057,N_3048,N_4207);
or U7058 (N_7058,N_2052,N_3417);
xor U7059 (N_7059,N_1032,N_885);
and U7060 (N_7060,N_608,N_2862);
nand U7061 (N_7061,N_1068,N_823);
or U7062 (N_7062,N_2942,N_1730);
nor U7063 (N_7063,N_488,N_430);
nand U7064 (N_7064,N_763,N_1570);
nand U7065 (N_7065,N_517,N_3025);
nor U7066 (N_7066,N_3515,N_2691);
nand U7067 (N_7067,N_4306,N_1622);
or U7068 (N_7068,N_253,N_1951);
and U7069 (N_7069,N_38,N_4559);
nand U7070 (N_7070,N_2586,N_1334);
nand U7071 (N_7071,N_1959,N_2955);
or U7072 (N_7072,N_1134,N_4359);
nand U7073 (N_7073,N_757,N_2339);
nand U7074 (N_7074,N_4322,N_4396);
and U7075 (N_7075,N_4605,N_3849);
and U7076 (N_7076,N_1316,N_3585);
nand U7077 (N_7077,N_863,N_1356);
xnor U7078 (N_7078,N_918,N_572);
nor U7079 (N_7079,N_4020,N_2656);
nor U7080 (N_7080,N_2869,N_3877);
nor U7081 (N_7081,N_3,N_3546);
nand U7082 (N_7082,N_842,N_2466);
and U7083 (N_7083,N_1295,N_4089);
nand U7084 (N_7084,N_791,N_460);
nand U7085 (N_7085,N_920,N_2856);
nor U7086 (N_7086,N_2154,N_4558);
or U7087 (N_7087,N_3286,N_2416);
nor U7088 (N_7088,N_2849,N_2488);
xor U7089 (N_7089,N_2710,N_3644);
and U7090 (N_7090,N_3588,N_2964);
xnor U7091 (N_7091,N_2597,N_814);
nand U7092 (N_7092,N_4338,N_2803);
or U7093 (N_7093,N_1912,N_1183);
and U7094 (N_7094,N_734,N_181);
and U7095 (N_7095,N_1610,N_869);
nand U7096 (N_7096,N_1882,N_2054);
and U7097 (N_7097,N_4968,N_1573);
nand U7098 (N_7098,N_4743,N_3506);
and U7099 (N_7099,N_1775,N_703);
nor U7100 (N_7100,N_1416,N_1418);
or U7101 (N_7101,N_93,N_2342);
nor U7102 (N_7102,N_2153,N_2934);
or U7103 (N_7103,N_3134,N_436);
nor U7104 (N_7104,N_881,N_2858);
nor U7105 (N_7105,N_802,N_2855);
and U7106 (N_7106,N_4691,N_3044);
nand U7107 (N_7107,N_1615,N_3004);
or U7108 (N_7108,N_933,N_1244);
nor U7109 (N_7109,N_1192,N_3063);
or U7110 (N_7110,N_199,N_1505);
or U7111 (N_7111,N_3002,N_4850);
nand U7112 (N_7112,N_4228,N_810);
or U7113 (N_7113,N_3845,N_4456);
nand U7114 (N_7114,N_2242,N_1928);
nand U7115 (N_7115,N_293,N_3050);
xnor U7116 (N_7116,N_4250,N_4244);
xor U7117 (N_7117,N_2658,N_114);
xnor U7118 (N_7118,N_597,N_3168);
nand U7119 (N_7119,N_1778,N_3105);
and U7120 (N_7120,N_104,N_268);
nor U7121 (N_7121,N_3475,N_2189);
and U7122 (N_7122,N_3600,N_4251);
nand U7123 (N_7123,N_2329,N_3331);
nand U7124 (N_7124,N_2657,N_4191);
and U7125 (N_7125,N_273,N_3695);
nor U7126 (N_7126,N_112,N_146);
nand U7127 (N_7127,N_1879,N_3403);
and U7128 (N_7128,N_1692,N_1508);
nor U7129 (N_7129,N_3911,N_2134);
nand U7130 (N_7130,N_475,N_3376);
nor U7131 (N_7131,N_3012,N_1208);
or U7132 (N_7132,N_3725,N_1094);
nand U7133 (N_7133,N_1686,N_937);
and U7134 (N_7134,N_3950,N_1126);
nand U7135 (N_7135,N_4813,N_2574);
nor U7136 (N_7136,N_2099,N_4488);
nand U7137 (N_7137,N_4186,N_3514);
nor U7138 (N_7138,N_845,N_3264);
nand U7139 (N_7139,N_4614,N_3941);
and U7140 (N_7140,N_3830,N_1214);
nand U7141 (N_7141,N_2730,N_1845);
nor U7142 (N_7142,N_2160,N_4090);
and U7143 (N_7143,N_106,N_3525);
nor U7144 (N_7144,N_1276,N_782);
nor U7145 (N_7145,N_4599,N_3333);
or U7146 (N_7146,N_2393,N_464);
or U7147 (N_7147,N_3734,N_1869);
and U7148 (N_7148,N_692,N_2305);
nor U7149 (N_7149,N_2974,N_3184);
and U7150 (N_7150,N_3248,N_2150);
nand U7151 (N_7151,N_1036,N_1757);
and U7152 (N_7152,N_3351,N_2660);
nand U7153 (N_7153,N_2135,N_550);
nand U7154 (N_7154,N_71,N_1387);
xnor U7155 (N_7155,N_3771,N_4991);
or U7156 (N_7156,N_413,N_420);
nand U7157 (N_7157,N_2034,N_1318);
nand U7158 (N_7158,N_557,N_2646);
nand U7159 (N_7159,N_1386,N_3477);
or U7160 (N_7160,N_3947,N_3311);
nor U7161 (N_7161,N_1184,N_69);
nand U7162 (N_7162,N_1140,N_2186);
nor U7163 (N_7163,N_3682,N_349);
xnor U7164 (N_7164,N_958,N_2565);
and U7165 (N_7165,N_22,N_3560);
nor U7166 (N_7166,N_3700,N_4951);
nor U7167 (N_7167,N_2677,N_2744);
or U7168 (N_7168,N_1790,N_2338);
nand U7169 (N_7169,N_3536,N_300);
xor U7170 (N_7170,N_2850,N_701);
and U7171 (N_7171,N_3748,N_334);
or U7172 (N_7172,N_3552,N_2930);
or U7173 (N_7173,N_4119,N_4007);
nand U7174 (N_7174,N_3073,N_4907);
or U7175 (N_7175,N_1145,N_1248);
and U7176 (N_7176,N_2985,N_402);
or U7177 (N_7177,N_532,N_2777);
nor U7178 (N_7178,N_4787,N_3837);
and U7179 (N_7179,N_392,N_3832);
nor U7180 (N_7180,N_4521,N_979);
nor U7181 (N_7181,N_4827,N_965);
nand U7182 (N_7182,N_827,N_4677);
nand U7183 (N_7183,N_4909,N_4642);
nor U7184 (N_7184,N_4288,N_716);
nand U7185 (N_7185,N_4774,N_556);
and U7186 (N_7186,N_3778,N_2720);
xnor U7187 (N_7187,N_2709,N_1093);
nor U7188 (N_7188,N_3171,N_13);
nor U7189 (N_7189,N_2021,N_3717);
nor U7190 (N_7190,N_513,N_6);
nand U7191 (N_7191,N_1712,N_1814);
xnor U7192 (N_7192,N_3071,N_3362);
xnor U7193 (N_7193,N_1886,N_1995);
nand U7194 (N_7194,N_1224,N_4150);
nor U7195 (N_7195,N_1548,N_3922);
and U7196 (N_7196,N_2173,N_1754);
nor U7197 (N_7197,N_2968,N_2035);
xnor U7198 (N_7198,N_2536,N_3614);
nor U7199 (N_7199,N_966,N_2172);
nand U7200 (N_7200,N_2943,N_808);
and U7201 (N_7201,N_2543,N_1150);
xor U7202 (N_7202,N_2537,N_2578);
nand U7203 (N_7203,N_4890,N_386);
or U7204 (N_7204,N_3186,N_3791);
and U7205 (N_7205,N_3349,N_873);
nor U7206 (N_7206,N_4277,N_1579);
or U7207 (N_7207,N_4428,N_4597);
and U7208 (N_7208,N_2705,N_3181);
nor U7209 (N_7209,N_180,N_3401);
and U7210 (N_7210,N_3275,N_1461);
nor U7211 (N_7211,N_2420,N_1056);
or U7212 (N_7212,N_923,N_894);
or U7213 (N_7213,N_4908,N_1298);
and U7214 (N_7214,N_3818,N_3366);
nand U7215 (N_7215,N_89,N_2896);
and U7216 (N_7216,N_2346,N_771);
nor U7217 (N_7217,N_2782,N_1174);
and U7218 (N_7218,N_866,N_4018);
nand U7219 (N_7219,N_668,N_1512);
nor U7220 (N_7220,N_4420,N_2655);
or U7221 (N_7221,N_147,N_80);
or U7222 (N_7222,N_1858,N_3578);
nor U7223 (N_7223,N_3451,N_4479);
nand U7224 (N_7224,N_1004,N_3956);
or U7225 (N_7225,N_3935,N_4235);
nor U7226 (N_7226,N_2629,N_1163);
or U7227 (N_7227,N_2080,N_2232);
and U7228 (N_7228,N_3212,N_1632);
and U7229 (N_7229,N_3497,N_3909);
nand U7230 (N_7230,N_3756,N_2568);
nor U7231 (N_7231,N_2373,N_847);
nand U7232 (N_7232,N_2345,N_2847);
and U7233 (N_7233,N_892,N_139);
and U7234 (N_7234,N_835,N_3667);
and U7235 (N_7235,N_3302,N_1572);
or U7236 (N_7236,N_1799,N_3053);
nand U7237 (N_7237,N_3924,N_2426);
nand U7238 (N_7238,N_4842,N_1659);
nor U7239 (N_7239,N_138,N_1983);
nor U7240 (N_7240,N_4103,N_613);
and U7241 (N_7241,N_4142,N_4061);
nor U7242 (N_7242,N_2757,N_1762);
or U7243 (N_7243,N_2008,N_1990);
or U7244 (N_7244,N_948,N_663);
and U7245 (N_7245,N_839,N_2371);
and U7246 (N_7246,N_3407,N_1889);
and U7247 (N_7247,N_506,N_4352);
and U7248 (N_7248,N_4204,N_2120);
or U7249 (N_7249,N_874,N_2133);
nor U7250 (N_7250,N_2532,N_1128);
nand U7251 (N_7251,N_2372,N_3637);
nor U7252 (N_7252,N_1303,N_2966);
nand U7253 (N_7253,N_2201,N_493);
and U7254 (N_7254,N_828,N_4432);
nor U7255 (N_7255,N_1544,N_1539);
nor U7256 (N_7256,N_492,N_2075);
nor U7257 (N_7257,N_3179,N_3077);
or U7258 (N_7258,N_3528,N_3219);
and U7259 (N_7259,N_4544,N_1781);
and U7260 (N_7260,N_3198,N_3088);
and U7261 (N_7261,N_1075,N_1308);
nand U7262 (N_7262,N_1905,N_2540);
nand U7263 (N_7263,N_4254,N_1366);
nor U7264 (N_7264,N_624,N_1930);
xor U7265 (N_7265,N_4038,N_2437);
nand U7266 (N_7266,N_1212,N_2237);
or U7267 (N_7267,N_4596,N_2480);
or U7268 (N_7268,N_4712,N_3096);
nand U7269 (N_7269,N_3509,N_596);
nand U7270 (N_7270,N_1336,N_4651);
nand U7271 (N_7271,N_3143,N_1476);
xnor U7272 (N_7272,N_445,N_2215);
nor U7273 (N_7273,N_3519,N_2409);
nand U7274 (N_7274,N_3931,N_3001);
nand U7275 (N_7275,N_1625,N_4855);
nand U7276 (N_7276,N_27,N_2229);
nand U7277 (N_7277,N_2192,N_95);
xnor U7278 (N_7278,N_2219,N_4364);
nor U7279 (N_7279,N_348,N_25);
or U7280 (N_7280,N_454,N_3500);
nand U7281 (N_7281,N_361,N_4122);
and U7282 (N_7282,N_1763,N_1235);
and U7283 (N_7283,N_1947,N_3434);
and U7284 (N_7284,N_1842,N_3030);
and U7285 (N_7285,N_1430,N_2801);
and U7286 (N_7286,N_1324,N_977);
xor U7287 (N_7287,N_184,N_3817);
nand U7288 (N_7288,N_3518,N_1545);
nor U7289 (N_7289,N_4568,N_3029);
and U7290 (N_7290,N_1694,N_1690);
nand U7291 (N_7291,N_4391,N_635);
nor U7292 (N_7292,N_395,N_4913);
nand U7293 (N_7293,N_3728,N_4184);
or U7294 (N_7294,N_57,N_1675);
and U7295 (N_7295,N_4263,N_1323);
nand U7296 (N_7296,N_1824,N_1121);
nor U7297 (N_7297,N_434,N_4511);
or U7298 (N_7298,N_1876,N_3710);
nor U7299 (N_7299,N_1044,N_3455);
nand U7300 (N_7300,N_0,N_2820);
and U7301 (N_7301,N_648,N_3340);
and U7302 (N_7302,N_2793,N_1154);
or U7303 (N_7303,N_4515,N_3543);
nand U7304 (N_7304,N_4070,N_778);
nand U7305 (N_7305,N_4801,N_2724);
nand U7306 (N_7306,N_4270,N_674);
nor U7307 (N_7307,N_3410,N_3089);
nor U7308 (N_7308,N_3722,N_2363);
and U7309 (N_7309,N_2472,N_4565);
nand U7310 (N_7310,N_4147,N_4137);
or U7311 (N_7311,N_3711,N_4917);
nand U7312 (N_7312,N_68,N_3693);
nand U7313 (N_7313,N_3892,N_4371);
nor U7314 (N_7314,N_521,N_4680);
nor U7315 (N_7315,N_2356,N_2689);
and U7316 (N_7316,N_3613,N_537);
or U7317 (N_7317,N_2330,N_1125);
xnor U7318 (N_7318,N_809,N_900);
nor U7319 (N_7319,N_411,N_2468);
and U7320 (N_7320,N_4218,N_4959);
nor U7321 (N_7321,N_2097,N_4477);
nand U7322 (N_7322,N_412,N_4302);
nor U7323 (N_7323,N_4601,N_3244);
or U7324 (N_7324,N_4487,N_2368);
nor U7325 (N_7325,N_691,N_4393);
and U7326 (N_7326,N_3865,N_1217);
nor U7327 (N_7327,N_1067,N_1792);
nand U7328 (N_7328,N_1598,N_3573);
and U7329 (N_7329,N_3320,N_4967);
and U7330 (N_7330,N_2551,N_4124);
or U7331 (N_7331,N_1300,N_4192);
nor U7332 (N_7332,N_3851,N_1860);
or U7333 (N_7333,N_3301,N_1488);
or U7334 (N_7334,N_870,N_3249);
nand U7335 (N_7335,N_1940,N_3632);
nor U7336 (N_7336,N_1190,N_3630);
and U7337 (N_7337,N_461,N_4531);
and U7338 (N_7338,N_1899,N_4547);
or U7339 (N_7339,N_1363,N_3781);
nor U7340 (N_7340,N_3997,N_956);
nand U7341 (N_7341,N_2500,N_2910);
or U7342 (N_7342,N_74,N_2128);
xnor U7343 (N_7343,N_1409,N_4985);
or U7344 (N_7344,N_162,N_4804);
nand U7345 (N_7345,N_904,N_49);
nand U7346 (N_7346,N_4440,N_3485);
or U7347 (N_7347,N_4851,N_375);
or U7348 (N_7348,N_2483,N_4012);
nor U7349 (N_7349,N_1023,N_2692);
and U7350 (N_7350,N_903,N_1820);
or U7351 (N_7351,N_2785,N_3383);
and U7352 (N_7352,N_4663,N_3678);
and U7353 (N_7353,N_2712,N_1705);
and U7354 (N_7354,N_2511,N_346);
or U7355 (N_7355,N_4824,N_4971);
or U7356 (N_7356,N_2202,N_1051);
nor U7357 (N_7357,N_1328,N_1786);
or U7358 (N_7358,N_3586,N_2742);
or U7359 (N_7359,N_345,N_1358);
nand U7360 (N_7360,N_2899,N_2292);
xor U7361 (N_7361,N_4246,N_3670);
xor U7362 (N_7362,N_3480,N_1582);
and U7363 (N_7363,N_4423,N_4507);
nor U7364 (N_7364,N_2410,N_3703);
or U7365 (N_7365,N_3060,N_3066);
nand U7366 (N_7366,N_508,N_4657);
nand U7367 (N_7367,N_377,N_3257);
and U7368 (N_7368,N_3680,N_3840);
and U7369 (N_7369,N_1777,N_3059);
nor U7370 (N_7370,N_2400,N_4374);
nor U7371 (N_7371,N_88,N_2463);
and U7372 (N_7372,N_151,N_531);
nor U7373 (N_7373,N_957,N_3058);
nor U7374 (N_7374,N_2740,N_1017);
or U7375 (N_7375,N_4514,N_2084);
nor U7376 (N_7376,N_1956,N_3110);
nand U7377 (N_7377,N_4631,N_2276);
or U7378 (N_7378,N_1315,N_3914);
nor U7379 (N_7379,N_3138,N_3270);
or U7380 (N_7380,N_3169,N_1985);
or U7381 (N_7381,N_1449,N_3441);
nor U7382 (N_7382,N_4388,N_1362);
and U7383 (N_7383,N_457,N_1619);
nand U7384 (N_7384,N_4799,N_1132);
nand U7385 (N_7385,N_1546,N_1417);
and U7386 (N_7386,N_447,N_1088);
or U7387 (N_7387,N_4429,N_2875);
nand U7388 (N_7388,N_4401,N_3507);
nand U7389 (N_7389,N_717,N_1464);
and U7390 (N_7390,N_1885,N_4190);
and U7391 (N_7391,N_518,N_1816);
or U7392 (N_7392,N_2559,N_1703);
nand U7393 (N_7393,N_1175,N_2003);
nand U7394 (N_7394,N_455,N_4409);
nand U7395 (N_7395,N_3864,N_282);
nand U7396 (N_7396,N_4938,N_439);
nand U7397 (N_7397,N_704,N_1585);
nor U7398 (N_7398,N_944,N_3384);
and U7399 (N_7399,N_17,N_3740);
or U7400 (N_7400,N_4002,N_4941);
nand U7401 (N_7401,N_318,N_1560);
or U7402 (N_7402,N_175,N_2259);
or U7403 (N_7403,N_2531,N_1311);
xor U7404 (N_7404,N_3776,N_688);
nand U7405 (N_7405,N_4730,N_254);
and U7406 (N_7406,N_2341,N_3015);
nand U7407 (N_7407,N_3467,N_4410);
nand U7408 (N_7408,N_1923,N_3988);
nand U7409 (N_7409,N_4504,N_4378);
nand U7410 (N_7410,N_689,N_4234);
nor U7411 (N_7411,N_3035,N_271);
nand U7412 (N_7412,N_2986,N_3926);
nand U7413 (N_7413,N_117,N_1742);
nor U7414 (N_7414,N_697,N_3398);
xor U7415 (N_7415,N_2051,N_3382);
nand U7416 (N_7416,N_3530,N_3738);
or U7417 (N_7417,N_2814,N_3620);
and U7418 (N_7418,N_4892,N_2747);
and U7419 (N_7419,N_4857,N_285);
nand U7420 (N_7420,N_1698,N_2425);
nand U7421 (N_7421,N_3737,N_2976);
or U7422 (N_7422,N_3836,N_3247);
or U7423 (N_7423,N_1455,N_3308);
or U7424 (N_7424,N_3823,N_286);
or U7425 (N_7425,N_2558,N_3570);
and U7426 (N_7426,N_2315,N_2727);
or U7427 (N_7427,N_2443,N_576);
or U7428 (N_7428,N_3605,N_4731);
nor U7429 (N_7429,N_4861,N_4902);
nand U7430 (N_7430,N_3178,N_1400);
nor U7431 (N_7431,N_660,N_2606);
nand U7432 (N_7432,N_2159,N_3420);
and U7433 (N_7433,N_2467,N_2256);
or U7434 (N_7434,N_911,N_726);
nand U7435 (N_7435,N_1306,N_3766);
nor U7436 (N_7436,N_4161,N_3136);
nand U7437 (N_7437,N_946,N_3772);
and U7438 (N_7438,N_4646,N_2746);
nand U7439 (N_7439,N_3251,N_3566);
xor U7440 (N_7440,N_4962,N_1843);
xor U7441 (N_7441,N_200,N_4587);
or U7442 (N_7442,N_4439,N_134);
and U7443 (N_7443,N_382,N_3193);
nand U7444 (N_7444,N_480,N_327);
or U7445 (N_7445,N_4918,N_2148);
or U7446 (N_7446,N_3508,N_1062);
or U7447 (N_7447,N_1687,N_3814);
and U7448 (N_7448,N_1419,N_2098);
and U7449 (N_7449,N_2407,N_4777);
or U7450 (N_7450,N_2819,N_3873);
or U7451 (N_7451,N_2344,N_2616);
or U7452 (N_7452,N_4078,N_50);
nand U7453 (N_7453,N_2362,N_3503);
and U7454 (N_7454,N_1979,N_316);
nand U7455 (N_7455,N_1722,N_4668);
and U7456 (N_7456,N_890,N_3282);
nor U7457 (N_7457,N_1773,N_860);
or U7458 (N_7458,N_1320,N_3945);
nand U7459 (N_7459,N_4602,N_204);
and U7460 (N_7460,N_3309,N_1015);
nand U7461 (N_7461,N_1070,N_4068);
nand U7462 (N_7462,N_2948,N_4814);
nor U7463 (N_7463,N_2422,N_4928);
nand U7464 (N_7464,N_3537,N_3108);
nand U7465 (N_7465,N_3595,N_3021);
nand U7466 (N_7466,N_4496,N_231);
nand U7467 (N_7467,N_974,N_16);
and U7468 (N_7468,N_2081,N_479);
or U7469 (N_7469,N_4136,N_352);
and U7470 (N_7470,N_4072,N_2509);
or U7471 (N_7471,N_4766,N_4956);
nand U7472 (N_7472,N_961,N_263);
or U7473 (N_7473,N_1565,N_2663);
nor U7474 (N_7474,N_2369,N_4087);
nor U7475 (N_7475,N_3385,N_3806);
and U7476 (N_7476,N_4329,N_1399);
or U7477 (N_7477,N_3075,N_4987);
or U7478 (N_7478,N_4760,N_1365);
nor U7479 (N_7479,N_2978,N_201);
xnor U7480 (N_7480,N_1903,N_3834);
or U7481 (N_7481,N_666,N_1631);
nand U7482 (N_7482,N_4341,N_4937);
nor U7483 (N_7483,N_768,N_463);
nand U7484 (N_7484,N_3027,N_1433);
nor U7485 (N_7485,N_4933,N_3991);
nand U7486 (N_7486,N_2241,N_3233);
and U7487 (N_7487,N_1523,N_3598);
and U7488 (N_7488,N_4397,N_2725);
or U7489 (N_7489,N_1547,N_3726);
or U7490 (N_7490,N_774,N_1511);
nor U7491 (N_7491,N_3483,N_925);
and U7492 (N_7492,N_3675,N_1403);
and U7493 (N_7493,N_2761,N_1871);
and U7494 (N_7494,N_3565,N_4999);
nand U7495 (N_7495,N_165,N_369);
and U7496 (N_7496,N_4166,N_3268);
or U7497 (N_7497,N_1802,N_4084);
or U7498 (N_7498,N_4261,N_1265);
or U7499 (N_7499,N_3596,N_2365);
nor U7500 (N_7500,N_4063,N_1041);
nand U7501 (N_7501,N_1570,N_3276);
and U7502 (N_7502,N_3224,N_1068);
nand U7503 (N_7503,N_960,N_4313);
and U7504 (N_7504,N_3851,N_2023);
or U7505 (N_7505,N_332,N_3183);
nor U7506 (N_7506,N_1006,N_4387);
or U7507 (N_7507,N_1968,N_4698);
and U7508 (N_7508,N_167,N_2562);
or U7509 (N_7509,N_3109,N_2772);
or U7510 (N_7510,N_872,N_325);
nand U7511 (N_7511,N_132,N_1194);
nand U7512 (N_7512,N_3344,N_4611);
nand U7513 (N_7513,N_2910,N_3564);
or U7514 (N_7514,N_3659,N_4737);
or U7515 (N_7515,N_4422,N_568);
nor U7516 (N_7516,N_1489,N_4061);
nand U7517 (N_7517,N_195,N_4596);
and U7518 (N_7518,N_2504,N_3972);
nand U7519 (N_7519,N_2173,N_3855);
and U7520 (N_7520,N_4103,N_1487);
or U7521 (N_7521,N_3370,N_2252);
nand U7522 (N_7522,N_2985,N_4849);
nand U7523 (N_7523,N_4871,N_4354);
nor U7524 (N_7524,N_841,N_3344);
nand U7525 (N_7525,N_4548,N_1447);
or U7526 (N_7526,N_1849,N_3803);
nand U7527 (N_7527,N_3920,N_208);
nand U7528 (N_7528,N_480,N_1058);
nand U7529 (N_7529,N_586,N_3012);
or U7530 (N_7530,N_1275,N_2818);
nor U7531 (N_7531,N_635,N_2759);
nor U7532 (N_7532,N_1493,N_1772);
and U7533 (N_7533,N_1961,N_325);
xor U7534 (N_7534,N_4776,N_3367);
nand U7535 (N_7535,N_3571,N_1496);
and U7536 (N_7536,N_1697,N_2443);
nor U7537 (N_7537,N_4481,N_630);
nor U7538 (N_7538,N_1248,N_3394);
xnor U7539 (N_7539,N_3617,N_367);
nand U7540 (N_7540,N_4193,N_4256);
nor U7541 (N_7541,N_209,N_4251);
xnor U7542 (N_7542,N_2204,N_2313);
and U7543 (N_7543,N_1354,N_365);
and U7544 (N_7544,N_3622,N_743);
and U7545 (N_7545,N_4868,N_881);
nand U7546 (N_7546,N_1009,N_4361);
and U7547 (N_7547,N_1727,N_4707);
nor U7548 (N_7548,N_3450,N_3053);
nand U7549 (N_7549,N_3144,N_66);
and U7550 (N_7550,N_262,N_3820);
or U7551 (N_7551,N_4739,N_4965);
nand U7552 (N_7552,N_1108,N_4966);
nand U7553 (N_7553,N_2033,N_2914);
and U7554 (N_7554,N_2653,N_2391);
nor U7555 (N_7555,N_274,N_4270);
nand U7556 (N_7556,N_261,N_2824);
xnor U7557 (N_7557,N_1439,N_4680);
or U7558 (N_7558,N_1085,N_4418);
nor U7559 (N_7559,N_1693,N_240);
nand U7560 (N_7560,N_728,N_2078);
nand U7561 (N_7561,N_4039,N_2429);
nor U7562 (N_7562,N_607,N_2510);
nand U7563 (N_7563,N_2511,N_1258);
nor U7564 (N_7564,N_851,N_2107);
or U7565 (N_7565,N_1006,N_1852);
xor U7566 (N_7566,N_4454,N_4277);
nor U7567 (N_7567,N_2899,N_3898);
and U7568 (N_7568,N_3699,N_1718);
or U7569 (N_7569,N_1552,N_2739);
and U7570 (N_7570,N_510,N_2665);
and U7571 (N_7571,N_4507,N_3947);
and U7572 (N_7572,N_3047,N_1538);
or U7573 (N_7573,N_2478,N_4);
and U7574 (N_7574,N_1651,N_3450);
or U7575 (N_7575,N_2837,N_2443);
or U7576 (N_7576,N_1156,N_2534);
or U7577 (N_7577,N_3971,N_1434);
nor U7578 (N_7578,N_3450,N_3492);
nor U7579 (N_7579,N_648,N_2700);
nand U7580 (N_7580,N_1183,N_1098);
nor U7581 (N_7581,N_887,N_2998);
nand U7582 (N_7582,N_3530,N_210);
nand U7583 (N_7583,N_4119,N_4013);
nand U7584 (N_7584,N_2393,N_2922);
or U7585 (N_7585,N_13,N_2238);
nor U7586 (N_7586,N_289,N_4508);
xnor U7587 (N_7587,N_185,N_2510);
nor U7588 (N_7588,N_3200,N_378);
or U7589 (N_7589,N_4839,N_1454);
and U7590 (N_7590,N_3777,N_4899);
nand U7591 (N_7591,N_2818,N_3269);
nor U7592 (N_7592,N_4653,N_209);
nor U7593 (N_7593,N_4648,N_4862);
xnor U7594 (N_7594,N_863,N_1237);
and U7595 (N_7595,N_3136,N_1064);
and U7596 (N_7596,N_1774,N_3792);
and U7597 (N_7597,N_2674,N_3957);
nor U7598 (N_7598,N_3071,N_931);
nand U7599 (N_7599,N_23,N_3335);
and U7600 (N_7600,N_143,N_4196);
nand U7601 (N_7601,N_4987,N_1840);
or U7602 (N_7602,N_23,N_4060);
nand U7603 (N_7603,N_3550,N_4383);
nor U7604 (N_7604,N_1983,N_4299);
and U7605 (N_7605,N_1439,N_1864);
or U7606 (N_7606,N_2073,N_4783);
nand U7607 (N_7607,N_852,N_165);
and U7608 (N_7608,N_3995,N_3296);
nand U7609 (N_7609,N_1228,N_2329);
nor U7610 (N_7610,N_1696,N_4688);
and U7611 (N_7611,N_479,N_3638);
xor U7612 (N_7612,N_3505,N_2389);
and U7613 (N_7613,N_2094,N_4364);
nand U7614 (N_7614,N_1504,N_150);
xnor U7615 (N_7615,N_4523,N_769);
and U7616 (N_7616,N_761,N_3809);
nand U7617 (N_7617,N_3233,N_2308);
nand U7618 (N_7618,N_1403,N_2532);
and U7619 (N_7619,N_3827,N_1119);
nand U7620 (N_7620,N_1220,N_3651);
nor U7621 (N_7621,N_4119,N_3334);
nand U7622 (N_7622,N_750,N_3835);
or U7623 (N_7623,N_310,N_3996);
nor U7624 (N_7624,N_1243,N_179);
nand U7625 (N_7625,N_616,N_4657);
or U7626 (N_7626,N_4481,N_3032);
and U7627 (N_7627,N_1547,N_2473);
and U7628 (N_7628,N_920,N_2437);
and U7629 (N_7629,N_1279,N_64);
nor U7630 (N_7630,N_1344,N_2840);
or U7631 (N_7631,N_2581,N_1026);
and U7632 (N_7632,N_1556,N_3556);
nand U7633 (N_7633,N_4727,N_2403);
nor U7634 (N_7634,N_1444,N_1519);
and U7635 (N_7635,N_1659,N_1740);
or U7636 (N_7636,N_1124,N_4487);
and U7637 (N_7637,N_1838,N_4758);
or U7638 (N_7638,N_2256,N_3970);
xor U7639 (N_7639,N_2213,N_1101);
and U7640 (N_7640,N_89,N_2394);
nand U7641 (N_7641,N_4563,N_2658);
and U7642 (N_7642,N_2794,N_4134);
or U7643 (N_7643,N_1995,N_4042);
or U7644 (N_7644,N_4134,N_1400);
nor U7645 (N_7645,N_856,N_2090);
nor U7646 (N_7646,N_1558,N_2359);
and U7647 (N_7647,N_1932,N_1972);
or U7648 (N_7648,N_331,N_4781);
nor U7649 (N_7649,N_2521,N_3535);
and U7650 (N_7650,N_1610,N_2439);
and U7651 (N_7651,N_2625,N_3886);
and U7652 (N_7652,N_3115,N_2334);
or U7653 (N_7653,N_344,N_570);
xnor U7654 (N_7654,N_389,N_4750);
nand U7655 (N_7655,N_4566,N_1532);
xor U7656 (N_7656,N_3257,N_4978);
nand U7657 (N_7657,N_4902,N_4834);
nand U7658 (N_7658,N_3771,N_4418);
nand U7659 (N_7659,N_4019,N_2083);
nor U7660 (N_7660,N_2880,N_1104);
or U7661 (N_7661,N_68,N_270);
and U7662 (N_7662,N_1288,N_1928);
and U7663 (N_7663,N_1679,N_3602);
nand U7664 (N_7664,N_828,N_2464);
nand U7665 (N_7665,N_2540,N_3393);
or U7666 (N_7666,N_4984,N_1791);
nor U7667 (N_7667,N_1225,N_4490);
nand U7668 (N_7668,N_4645,N_3021);
or U7669 (N_7669,N_3052,N_1018);
nand U7670 (N_7670,N_3041,N_1187);
nand U7671 (N_7671,N_1745,N_4776);
nand U7672 (N_7672,N_498,N_4363);
and U7673 (N_7673,N_4023,N_4380);
and U7674 (N_7674,N_1035,N_117);
nor U7675 (N_7675,N_4167,N_4514);
or U7676 (N_7676,N_1466,N_177);
and U7677 (N_7677,N_1767,N_4633);
nor U7678 (N_7678,N_2745,N_463);
nand U7679 (N_7679,N_2988,N_3990);
or U7680 (N_7680,N_3369,N_1768);
or U7681 (N_7681,N_355,N_3753);
and U7682 (N_7682,N_4660,N_3732);
nand U7683 (N_7683,N_2162,N_1142);
nand U7684 (N_7684,N_2535,N_2293);
nor U7685 (N_7685,N_564,N_924);
or U7686 (N_7686,N_3954,N_3065);
or U7687 (N_7687,N_2545,N_3768);
nor U7688 (N_7688,N_2580,N_413);
nand U7689 (N_7689,N_907,N_2019);
nor U7690 (N_7690,N_3039,N_3132);
nor U7691 (N_7691,N_1685,N_2915);
nand U7692 (N_7692,N_3945,N_1879);
or U7693 (N_7693,N_2263,N_535);
nand U7694 (N_7694,N_3257,N_1351);
and U7695 (N_7695,N_2769,N_2172);
or U7696 (N_7696,N_1487,N_2445);
nand U7697 (N_7697,N_3458,N_2496);
nor U7698 (N_7698,N_1145,N_1348);
and U7699 (N_7699,N_600,N_3023);
or U7700 (N_7700,N_4746,N_4387);
and U7701 (N_7701,N_3653,N_189);
nand U7702 (N_7702,N_2595,N_3925);
or U7703 (N_7703,N_4411,N_4050);
or U7704 (N_7704,N_4695,N_685);
and U7705 (N_7705,N_2074,N_4641);
and U7706 (N_7706,N_1195,N_2724);
nand U7707 (N_7707,N_2522,N_1924);
nor U7708 (N_7708,N_861,N_2350);
nand U7709 (N_7709,N_934,N_589);
or U7710 (N_7710,N_2999,N_2886);
nand U7711 (N_7711,N_952,N_1179);
nor U7712 (N_7712,N_4080,N_1474);
and U7713 (N_7713,N_2235,N_4830);
and U7714 (N_7714,N_558,N_505);
nand U7715 (N_7715,N_2843,N_3560);
nand U7716 (N_7716,N_101,N_79);
nor U7717 (N_7717,N_2374,N_2532);
or U7718 (N_7718,N_4274,N_3773);
nand U7719 (N_7719,N_3777,N_3210);
or U7720 (N_7720,N_4179,N_1096);
nor U7721 (N_7721,N_1481,N_4102);
nor U7722 (N_7722,N_3316,N_1198);
nor U7723 (N_7723,N_3543,N_1170);
nor U7724 (N_7724,N_1237,N_2599);
nor U7725 (N_7725,N_4794,N_976);
and U7726 (N_7726,N_1357,N_3211);
nor U7727 (N_7727,N_1491,N_1383);
nand U7728 (N_7728,N_3190,N_4019);
or U7729 (N_7729,N_4236,N_1206);
nor U7730 (N_7730,N_3330,N_3726);
nand U7731 (N_7731,N_2142,N_1750);
or U7732 (N_7732,N_953,N_3582);
nor U7733 (N_7733,N_690,N_426);
nand U7734 (N_7734,N_3783,N_1288);
and U7735 (N_7735,N_133,N_4293);
or U7736 (N_7736,N_3698,N_1586);
nor U7737 (N_7737,N_4384,N_1371);
and U7738 (N_7738,N_389,N_3624);
nor U7739 (N_7739,N_4980,N_37);
and U7740 (N_7740,N_3767,N_4401);
nand U7741 (N_7741,N_1838,N_2578);
nand U7742 (N_7742,N_2330,N_1567);
and U7743 (N_7743,N_1758,N_1563);
nand U7744 (N_7744,N_2083,N_3623);
nand U7745 (N_7745,N_4582,N_3043);
nand U7746 (N_7746,N_4731,N_584);
nand U7747 (N_7747,N_1060,N_3225);
nor U7748 (N_7748,N_1532,N_4518);
nor U7749 (N_7749,N_3158,N_2942);
or U7750 (N_7750,N_993,N_1196);
nand U7751 (N_7751,N_4368,N_3529);
and U7752 (N_7752,N_2951,N_1000);
nand U7753 (N_7753,N_1070,N_542);
nand U7754 (N_7754,N_1800,N_4182);
and U7755 (N_7755,N_3144,N_328);
nand U7756 (N_7756,N_896,N_3592);
nor U7757 (N_7757,N_1472,N_4327);
and U7758 (N_7758,N_3460,N_4376);
or U7759 (N_7759,N_15,N_3741);
nor U7760 (N_7760,N_2955,N_3719);
and U7761 (N_7761,N_3018,N_2900);
nor U7762 (N_7762,N_4236,N_3300);
or U7763 (N_7763,N_1296,N_2413);
nor U7764 (N_7764,N_3052,N_4955);
xor U7765 (N_7765,N_4058,N_1625);
nor U7766 (N_7766,N_2282,N_1682);
nor U7767 (N_7767,N_2084,N_855);
nand U7768 (N_7768,N_1254,N_4700);
nor U7769 (N_7769,N_2541,N_2506);
nand U7770 (N_7770,N_4461,N_3644);
nor U7771 (N_7771,N_3031,N_1174);
nand U7772 (N_7772,N_834,N_4507);
xnor U7773 (N_7773,N_1044,N_807);
nor U7774 (N_7774,N_1572,N_877);
or U7775 (N_7775,N_3181,N_2395);
or U7776 (N_7776,N_2253,N_2928);
nand U7777 (N_7777,N_1362,N_81);
or U7778 (N_7778,N_3970,N_4542);
nand U7779 (N_7779,N_750,N_522);
nand U7780 (N_7780,N_2665,N_338);
nand U7781 (N_7781,N_454,N_4659);
and U7782 (N_7782,N_229,N_2468);
nand U7783 (N_7783,N_861,N_3471);
or U7784 (N_7784,N_2251,N_3820);
or U7785 (N_7785,N_1749,N_2561);
and U7786 (N_7786,N_3369,N_1293);
xnor U7787 (N_7787,N_4466,N_2659);
and U7788 (N_7788,N_1873,N_1854);
or U7789 (N_7789,N_1564,N_4841);
nand U7790 (N_7790,N_3334,N_3787);
and U7791 (N_7791,N_4754,N_4013);
and U7792 (N_7792,N_2553,N_2820);
nand U7793 (N_7793,N_2865,N_525);
xnor U7794 (N_7794,N_3502,N_1523);
or U7795 (N_7795,N_4024,N_474);
and U7796 (N_7796,N_1847,N_3478);
nand U7797 (N_7797,N_1452,N_3216);
nor U7798 (N_7798,N_4971,N_3388);
nand U7799 (N_7799,N_4599,N_4198);
nor U7800 (N_7800,N_2391,N_2752);
or U7801 (N_7801,N_63,N_2738);
nor U7802 (N_7802,N_2228,N_2439);
nand U7803 (N_7803,N_135,N_3908);
and U7804 (N_7804,N_1228,N_4105);
nor U7805 (N_7805,N_4660,N_3181);
xor U7806 (N_7806,N_4177,N_1699);
and U7807 (N_7807,N_1974,N_2067);
or U7808 (N_7808,N_4193,N_1315);
or U7809 (N_7809,N_1033,N_1363);
and U7810 (N_7810,N_1522,N_3059);
or U7811 (N_7811,N_4250,N_1863);
nand U7812 (N_7812,N_3913,N_1369);
or U7813 (N_7813,N_4372,N_125);
or U7814 (N_7814,N_3165,N_2730);
nand U7815 (N_7815,N_4382,N_40);
and U7816 (N_7816,N_2653,N_1596);
and U7817 (N_7817,N_4979,N_1603);
xnor U7818 (N_7818,N_523,N_1870);
nor U7819 (N_7819,N_1336,N_4952);
nand U7820 (N_7820,N_14,N_279);
nor U7821 (N_7821,N_4037,N_1804);
and U7822 (N_7822,N_330,N_2411);
nand U7823 (N_7823,N_477,N_3969);
and U7824 (N_7824,N_4968,N_3417);
or U7825 (N_7825,N_2499,N_368);
nand U7826 (N_7826,N_3470,N_4157);
nand U7827 (N_7827,N_4482,N_2052);
or U7828 (N_7828,N_3650,N_4408);
nand U7829 (N_7829,N_3500,N_1575);
nand U7830 (N_7830,N_3189,N_2638);
and U7831 (N_7831,N_2557,N_4775);
nand U7832 (N_7832,N_2123,N_4142);
and U7833 (N_7833,N_634,N_384);
and U7834 (N_7834,N_4026,N_692);
and U7835 (N_7835,N_3772,N_2446);
and U7836 (N_7836,N_1801,N_3686);
and U7837 (N_7837,N_2577,N_4817);
and U7838 (N_7838,N_3096,N_382);
nor U7839 (N_7839,N_42,N_2561);
nand U7840 (N_7840,N_4245,N_2391);
or U7841 (N_7841,N_3857,N_3500);
and U7842 (N_7842,N_1317,N_221);
and U7843 (N_7843,N_1160,N_963);
or U7844 (N_7844,N_812,N_4548);
nor U7845 (N_7845,N_3201,N_374);
or U7846 (N_7846,N_2828,N_1897);
or U7847 (N_7847,N_2075,N_2457);
or U7848 (N_7848,N_2964,N_2364);
nor U7849 (N_7849,N_4764,N_277);
and U7850 (N_7850,N_4237,N_3932);
nand U7851 (N_7851,N_4915,N_4223);
nor U7852 (N_7852,N_330,N_4626);
nand U7853 (N_7853,N_3678,N_697);
nand U7854 (N_7854,N_895,N_4331);
and U7855 (N_7855,N_3296,N_253);
nand U7856 (N_7856,N_1390,N_1205);
nor U7857 (N_7857,N_4002,N_4237);
nor U7858 (N_7858,N_295,N_4695);
or U7859 (N_7859,N_3441,N_4152);
and U7860 (N_7860,N_1125,N_764);
and U7861 (N_7861,N_3597,N_2431);
nand U7862 (N_7862,N_2008,N_2682);
nor U7863 (N_7863,N_4055,N_495);
and U7864 (N_7864,N_718,N_1651);
or U7865 (N_7865,N_348,N_4977);
nand U7866 (N_7866,N_543,N_4939);
or U7867 (N_7867,N_3909,N_3057);
nand U7868 (N_7868,N_4337,N_1807);
nand U7869 (N_7869,N_3160,N_1687);
or U7870 (N_7870,N_1213,N_4304);
and U7871 (N_7871,N_1763,N_3411);
and U7872 (N_7872,N_4666,N_1234);
or U7873 (N_7873,N_852,N_4278);
and U7874 (N_7874,N_3535,N_2112);
nor U7875 (N_7875,N_2470,N_4674);
and U7876 (N_7876,N_3432,N_3214);
nand U7877 (N_7877,N_4069,N_1933);
nand U7878 (N_7878,N_2360,N_2659);
nand U7879 (N_7879,N_2595,N_132);
nand U7880 (N_7880,N_1751,N_2141);
and U7881 (N_7881,N_4636,N_2899);
nand U7882 (N_7882,N_3293,N_3510);
or U7883 (N_7883,N_2366,N_3918);
nand U7884 (N_7884,N_696,N_4389);
xnor U7885 (N_7885,N_1605,N_4637);
nor U7886 (N_7886,N_3153,N_3648);
nor U7887 (N_7887,N_1583,N_2535);
nand U7888 (N_7888,N_1354,N_4816);
xnor U7889 (N_7889,N_23,N_3266);
nor U7890 (N_7890,N_4829,N_3883);
or U7891 (N_7891,N_1370,N_3496);
nor U7892 (N_7892,N_634,N_3202);
or U7893 (N_7893,N_4156,N_3025);
nand U7894 (N_7894,N_4206,N_1549);
nor U7895 (N_7895,N_1216,N_2853);
nand U7896 (N_7896,N_2152,N_1862);
or U7897 (N_7897,N_483,N_4899);
and U7898 (N_7898,N_3137,N_4803);
and U7899 (N_7899,N_551,N_3591);
and U7900 (N_7900,N_3888,N_1377);
nor U7901 (N_7901,N_4347,N_1429);
and U7902 (N_7902,N_4956,N_4858);
xor U7903 (N_7903,N_1627,N_4093);
nor U7904 (N_7904,N_1758,N_4787);
and U7905 (N_7905,N_1744,N_4250);
and U7906 (N_7906,N_1989,N_2685);
nand U7907 (N_7907,N_1086,N_2122);
nand U7908 (N_7908,N_2468,N_4893);
nand U7909 (N_7909,N_3623,N_1590);
and U7910 (N_7910,N_2079,N_56);
nor U7911 (N_7911,N_3103,N_496);
or U7912 (N_7912,N_144,N_2013);
xnor U7913 (N_7913,N_1558,N_313);
nor U7914 (N_7914,N_2826,N_3189);
and U7915 (N_7915,N_2466,N_47);
and U7916 (N_7916,N_1327,N_4540);
and U7917 (N_7917,N_334,N_1559);
or U7918 (N_7918,N_4635,N_4205);
nand U7919 (N_7919,N_2522,N_3666);
and U7920 (N_7920,N_247,N_4500);
and U7921 (N_7921,N_86,N_2579);
nand U7922 (N_7922,N_4197,N_2256);
and U7923 (N_7923,N_3955,N_420);
nor U7924 (N_7924,N_3996,N_4364);
and U7925 (N_7925,N_417,N_4115);
or U7926 (N_7926,N_3173,N_760);
or U7927 (N_7927,N_2571,N_4852);
or U7928 (N_7928,N_2303,N_1492);
or U7929 (N_7929,N_4955,N_3990);
and U7930 (N_7930,N_1696,N_507);
nand U7931 (N_7931,N_1941,N_2511);
or U7932 (N_7932,N_3826,N_2743);
nor U7933 (N_7933,N_1588,N_3313);
nor U7934 (N_7934,N_4104,N_287);
nor U7935 (N_7935,N_3304,N_4350);
or U7936 (N_7936,N_1949,N_885);
nand U7937 (N_7937,N_4389,N_3063);
nor U7938 (N_7938,N_4921,N_100);
and U7939 (N_7939,N_1207,N_1684);
nor U7940 (N_7940,N_1560,N_4223);
nor U7941 (N_7941,N_3415,N_1940);
nor U7942 (N_7942,N_3374,N_2650);
or U7943 (N_7943,N_644,N_1933);
and U7944 (N_7944,N_211,N_1416);
nor U7945 (N_7945,N_3916,N_2922);
or U7946 (N_7946,N_826,N_201);
or U7947 (N_7947,N_4263,N_670);
or U7948 (N_7948,N_1972,N_657);
or U7949 (N_7949,N_601,N_4134);
or U7950 (N_7950,N_3935,N_139);
nand U7951 (N_7951,N_1857,N_4389);
and U7952 (N_7952,N_4409,N_4183);
or U7953 (N_7953,N_1180,N_1849);
or U7954 (N_7954,N_4652,N_3095);
and U7955 (N_7955,N_2727,N_3143);
and U7956 (N_7956,N_3356,N_3753);
nand U7957 (N_7957,N_2406,N_1229);
nand U7958 (N_7958,N_188,N_1256);
or U7959 (N_7959,N_321,N_3127);
nand U7960 (N_7960,N_668,N_4964);
nor U7961 (N_7961,N_2449,N_4574);
nor U7962 (N_7962,N_43,N_2507);
and U7963 (N_7963,N_1004,N_2187);
and U7964 (N_7964,N_3180,N_1440);
or U7965 (N_7965,N_2668,N_1114);
nand U7966 (N_7966,N_4705,N_4718);
and U7967 (N_7967,N_3704,N_1433);
nor U7968 (N_7968,N_3584,N_4795);
or U7969 (N_7969,N_4927,N_4575);
and U7970 (N_7970,N_3766,N_4076);
xnor U7971 (N_7971,N_2468,N_4797);
xnor U7972 (N_7972,N_3764,N_2972);
and U7973 (N_7973,N_2628,N_4742);
nor U7974 (N_7974,N_3433,N_2133);
and U7975 (N_7975,N_583,N_1583);
or U7976 (N_7976,N_2560,N_3016);
and U7977 (N_7977,N_13,N_1371);
and U7978 (N_7978,N_4909,N_110);
or U7979 (N_7979,N_3580,N_3411);
or U7980 (N_7980,N_3096,N_399);
nand U7981 (N_7981,N_3355,N_1060);
nand U7982 (N_7982,N_4625,N_2760);
or U7983 (N_7983,N_4239,N_4697);
or U7984 (N_7984,N_232,N_4973);
nand U7985 (N_7985,N_3228,N_1704);
and U7986 (N_7986,N_3320,N_2516);
nor U7987 (N_7987,N_4124,N_1115);
nor U7988 (N_7988,N_3206,N_770);
and U7989 (N_7989,N_943,N_3982);
nor U7990 (N_7990,N_464,N_1983);
nor U7991 (N_7991,N_2500,N_4932);
and U7992 (N_7992,N_2427,N_195);
nor U7993 (N_7993,N_3616,N_3990);
or U7994 (N_7994,N_3330,N_3749);
and U7995 (N_7995,N_4596,N_2040);
nand U7996 (N_7996,N_1276,N_2823);
nor U7997 (N_7997,N_1318,N_3528);
nand U7998 (N_7998,N_3113,N_1361);
or U7999 (N_7999,N_1089,N_1751);
nor U8000 (N_8000,N_2638,N_1260);
and U8001 (N_8001,N_4809,N_1218);
nand U8002 (N_8002,N_214,N_4084);
or U8003 (N_8003,N_3347,N_2525);
or U8004 (N_8004,N_3619,N_4605);
or U8005 (N_8005,N_3432,N_858);
xnor U8006 (N_8006,N_1218,N_4011);
and U8007 (N_8007,N_1567,N_3863);
or U8008 (N_8008,N_92,N_2108);
and U8009 (N_8009,N_415,N_2885);
nand U8010 (N_8010,N_3161,N_630);
nand U8011 (N_8011,N_3274,N_3362);
nand U8012 (N_8012,N_400,N_2405);
and U8013 (N_8013,N_4904,N_2323);
and U8014 (N_8014,N_3242,N_118);
nand U8015 (N_8015,N_798,N_1151);
or U8016 (N_8016,N_3614,N_3949);
nor U8017 (N_8017,N_3269,N_4285);
and U8018 (N_8018,N_1100,N_3205);
nor U8019 (N_8019,N_3214,N_2685);
nand U8020 (N_8020,N_833,N_3505);
and U8021 (N_8021,N_4488,N_3575);
or U8022 (N_8022,N_3294,N_1929);
nor U8023 (N_8023,N_1816,N_1793);
nor U8024 (N_8024,N_3269,N_2195);
nor U8025 (N_8025,N_4286,N_3298);
nor U8026 (N_8026,N_4781,N_3570);
and U8027 (N_8027,N_3352,N_2403);
and U8028 (N_8028,N_866,N_984);
nand U8029 (N_8029,N_1857,N_3655);
nor U8030 (N_8030,N_4771,N_3726);
nor U8031 (N_8031,N_4244,N_940);
nor U8032 (N_8032,N_1825,N_4914);
nor U8033 (N_8033,N_1796,N_1391);
and U8034 (N_8034,N_8,N_2789);
nor U8035 (N_8035,N_3184,N_2171);
or U8036 (N_8036,N_2079,N_2475);
and U8037 (N_8037,N_4636,N_1773);
and U8038 (N_8038,N_324,N_4329);
nand U8039 (N_8039,N_1788,N_132);
nor U8040 (N_8040,N_1363,N_4467);
or U8041 (N_8041,N_3960,N_3613);
nor U8042 (N_8042,N_2070,N_2816);
nor U8043 (N_8043,N_1268,N_3159);
and U8044 (N_8044,N_4018,N_830);
nand U8045 (N_8045,N_2673,N_3720);
or U8046 (N_8046,N_2479,N_3558);
nor U8047 (N_8047,N_4484,N_1465);
nor U8048 (N_8048,N_2445,N_3504);
and U8049 (N_8049,N_2751,N_1086);
nand U8050 (N_8050,N_1596,N_642);
or U8051 (N_8051,N_386,N_2932);
nor U8052 (N_8052,N_994,N_4051);
nand U8053 (N_8053,N_2731,N_3857);
or U8054 (N_8054,N_2270,N_4830);
or U8055 (N_8055,N_9,N_3825);
or U8056 (N_8056,N_1427,N_4429);
or U8057 (N_8057,N_491,N_3313);
nand U8058 (N_8058,N_1228,N_3437);
and U8059 (N_8059,N_966,N_3126);
and U8060 (N_8060,N_3640,N_2040);
or U8061 (N_8061,N_965,N_1327);
or U8062 (N_8062,N_3652,N_3530);
or U8063 (N_8063,N_2998,N_2967);
nand U8064 (N_8064,N_4386,N_3927);
nor U8065 (N_8065,N_4774,N_2418);
and U8066 (N_8066,N_1913,N_102);
nor U8067 (N_8067,N_1055,N_1843);
and U8068 (N_8068,N_370,N_859);
and U8069 (N_8069,N_3527,N_1378);
nand U8070 (N_8070,N_4450,N_3874);
and U8071 (N_8071,N_3576,N_1191);
nor U8072 (N_8072,N_2062,N_4898);
or U8073 (N_8073,N_3996,N_2729);
and U8074 (N_8074,N_4192,N_4837);
and U8075 (N_8075,N_2929,N_2058);
nand U8076 (N_8076,N_4036,N_2758);
nand U8077 (N_8077,N_1775,N_1638);
and U8078 (N_8078,N_1344,N_4218);
nand U8079 (N_8079,N_3319,N_313);
or U8080 (N_8080,N_2294,N_1717);
or U8081 (N_8081,N_4523,N_4060);
nand U8082 (N_8082,N_4987,N_102);
or U8083 (N_8083,N_3105,N_160);
nand U8084 (N_8084,N_280,N_2343);
or U8085 (N_8085,N_4367,N_1794);
nand U8086 (N_8086,N_3772,N_423);
or U8087 (N_8087,N_212,N_1829);
or U8088 (N_8088,N_2435,N_4425);
and U8089 (N_8089,N_3947,N_228);
or U8090 (N_8090,N_2242,N_3671);
and U8091 (N_8091,N_1866,N_3025);
or U8092 (N_8092,N_3400,N_2270);
xnor U8093 (N_8093,N_1105,N_3815);
and U8094 (N_8094,N_1494,N_3497);
and U8095 (N_8095,N_17,N_4445);
or U8096 (N_8096,N_4924,N_4950);
nor U8097 (N_8097,N_4345,N_3170);
or U8098 (N_8098,N_4022,N_470);
or U8099 (N_8099,N_2996,N_2027);
and U8100 (N_8100,N_4500,N_2549);
nor U8101 (N_8101,N_4029,N_890);
and U8102 (N_8102,N_3315,N_2822);
nand U8103 (N_8103,N_1337,N_524);
nor U8104 (N_8104,N_973,N_1294);
or U8105 (N_8105,N_1410,N_3090);
and U8106 (N_8106,N_101,N_755);
and U8107 (N_8107,N_3371,N_3220);
or U8108 (N_8108,N_1574,N_2682);
or U8109 (N_8109,N_2278,N_3464);
or U8110 (N_8110,N_531,N_635);
or U8111 (N_8111,N_3778,N_1413);
xor U8112 (N_8112,N_3151,N_1905);
nand U8113 (N_8113,N_269,N_278);
or U8114 (N_8114,N_707,N_3729);
nand U8115 (N_8115,N_4743,N_4963);
nor U8116 (N_8116,N_1175,N_4879);
or U8117 (N_8117,N_2219,N_3387);
xnor U8118 (N_8118,N_2518,N_1209);
nand U8119 (N_8119,N_801,N_87);
nand U8120 (N_8120,N_833,N_2933);
nor U8121 (N_8121,N_4190,N_187);
or U8122 (N_8122,N_916,N_2440);
nor U8123 (N_8123,N_3277,N_2123);
nand U8124 (N_8124,N_2001,N_1864);
nor U8125 (N_8125,N_655,N_2819);
or U8126 (N_8126,N_4516,N_2441);
or U8127 (N_8127,N_4307,N_3509);
or U8128 (N_8128,N_1537,N_1476);
xor U8129 (N_8129,N_1267,N_4385);
or U8130 (N_8130,N_510,N_3085);
or U8131 (N_8131,N_3416,N_3809);
nand U8132 (N_8132,N_2809,N_2862);
xor U8133 (N_8133,N_59,N_626);
and U8134 (N_8134,N_1150,N_2634);
nand U8135 (N_8135,N_116,N_4845);
nand U8136 (N_8136,N_856,N_4430);
xor U8137 (N_8137,N_277,N_2088);
nand U8138 (N_8138,N_4324,N_2036);
nand U8139 (N_8139,N_3646,N_1622);
or U8140 (N_8140,N_4031,N_1600);
or U8141 (N_8141,N_2713,N_1845);
and U8142 (N_8142,N_1742,N_23);
nand U8143 (N_8143,N_2321,N_563);
nand U8144 (N_8144,N_2339,N_3135);
nor U8145 (N_8145,N_2432,N_3179);
nand U8146 (N_8146,N_1165,N_3790);
nor U8147 (N_8147,N_1661,N_2667);
nor U8148 (N_8148,N_1058,N_4042);
or U8149 (N_8149,N_2918,N_3918);
and U8150 (N_8150,N_1161,N_1821);
and U8151 (N_8151,N_473,N_1259);
nand U8152 (N_8152,N_3588,N_3265);
nand U8153 (N_8153,N_3297,N_4523);
nor U8154 (N_8154,N_764,N_4755);
nand U8155 (N_8155,N_3595,N_4667);
nor U8156 (N_8156,N_174,N_4139);
nand U8157 (N_8157,N_3264,N_4577);
and U8158 (N_8158,N_404,N_1828);
nand U8159 (N_8159,N_936,N_728);
nand U8160 (N_8160,N_2516,N_947);
and U8161 (N_8161,N_2876,N_4770);
or U8162 (N_8162,N_4690,N_3069);
nor U8163 (N_8163,N_1170,N_729);
or U8164 (N_8164,N_2170,N_4156);
or U8165 (N_8165,N_3491,N_1819);
or U8166 (N_8166,N_4158,N_243);
nor U8167 (N_8167,N_4329,N_101);
or U8168 (N_8168,N_1821,N_570);
nand U8169 (N_8169,N_1078,N_1350);
nand U8170 (N_8170,N_3485,N_2217);
or U8171 (N_8171,N_3832,N_4747);
and U8172 (N_8172,N_725,N_831);
and U8173 (N_8173,N_2472,N_1066);
nand U8174 (N_8174,N_4110,N_1299);
and U8175 (N_8175,N_3747,N_1358);
or U8176 (N_8176,N_2093,N_3746);
or U8177 (N_8177,N_1856,N_1411);
nand U8178 (N_8178,N_1510,N_1058);
nand U8179 (N_8179,N_4658,N_208);
or U8180 (N_8180,N_4582,N_2177);
or U8181 (N_8181,N_699,N_2136);
and U8182 (N_8182,N_1358,N_1137);
xnor U8183 (N_8183,N_1693,N_4049);
nand U8184 (N_8184,N_1643,N_346);
or U8185 (N_8185,N_4579,N_1461);
nand U8186 (N_8186,N_4495,N_2800);
nor U8187 (N_8187,N_4888,N_4401);
nor U8188 (N_8188,N_4541,N_1340);
or U8189 (N_8189,N_3659,N_821);
nand U8190 (N_8190,N_2696,N_4595);
nor U8191 (N_8191,N_356,N_0);
nor U8192 (N_8192,N_4828,N_4924);
nor U8193 (N_8193,N_1975,N_1395);
nand U8194 (N_8194,N_2956,N_4170);
and U8195 (N_8195,N_112,N_870);
nand U8196 (N_8196,N_1452,N_1054);
nor U8197 (N_8197,N_1676,N_3260);
nor U8198 (N_8198,N_2808,N_1565);
nor U8199 (N_8199,N_1162,N_1021);
or U8200 (N_8200,N_2858,N_4001);
and U8201 (N_8201,N_3594,N_814);
nor U8202 (N_8202,N_4808,N_1804);
nor U8203 (N_8203,N_154,N_754);
nand U8204 (N_8204,N_3203,N_3755);
nor U8205 (N_8205,N_2853,N_1091);
or U8206 (N_8206,N_2434,N_3273);
or U8207 (N_8207,N_4628,N_4704);
or U8208 (N_8208,N_2849,N_2337);
and U8209 (N_8209,N_3877,N_4934);
or U8210 (N_8210,N_933,N_4858);
nor U8211 (N_8211,N_3148,N_3043);
nor U8212 (N_8212,N_2131,N_3440);
or U8213 (N_8213,N_3400,N_712);
nand U8214 (N_8214,N_332,N_483);
and U8215 (N_8215,N_2810,N_458);
nor U8216 (N_8216,N_2317,N_2519);
or U8217 (N_8217,N_4015,N_4109);
nand U8218 (N_8218,N_1756,N_1826);
and U8219 (N_8219,N_1109,N_2844);
nand U8220 (N_8220,N_4066,N_2845);
nor U8221 (N_8221,N_1191,N_3391);
nor U8222 (N_8222,N_4882,N_3575);
xor U8223 (N_8223,N_2278,N_4310);
nand U8224 (N_8224,N_1427,N_4282);
or U8225 (N_8225,N_4565,N_2147);
and U8226 (N_8226,N_439,N_1846);
nand U8227 (N_8227,N_4236,N_2090);
and U8228 (N_8228,N_3735,N_3508);
nand U8229 (N_8229,N_3159,N_310);
nand U8230 (N_8230,N_3590,N_467);
and U8231 (N_8231,N_2505,N_409);
or U8232 (N_8232,N_3328,N_1504);
or U8233 (N_8233,N_113,N_4348);
or U8234 (N_8234,N_3888,N_4647);
nand U8235 (N_8235,N_2637,N_1465);
or U8236 (N_8236,N_3913,N_2095);
nand U8237 (N_8237,N_4236,N_3635);
nand U8238 (N_8238,N_1921,N_2145);
and U8239 (N_8239,N_4575,N_3508);
or U8240 (N_8240,N_3276,N_3357);
nand U8241 (N_8241,N_1589,N_4531);
nor U8242 (N_8242,N_950,N_554);
and U8243 (N_8243,N_2045,N_524);
or U8244 (N_8244,N_145,N_1680);
and U8245 (N_8245,N_1907,N_3763);
and U8246 (N_8246,N_3399,N_4931);
and U8247 (N_8247,N_2920,N_1968);
or U8248 (N_8248,N_2396,N_4864);
nand U8249 (N_8249,N_1660,N_1944);
or U8250 (N_8250,N_988,N_523);
nand U8251 (N_8251,N_4964,N_4032);
and U8252 (N_8252,N_166,N_3919);
and U8253 (N_8253,N_4433,N_1120);
nor U8254 (N_8254,N_2828,N_4356);
or U8255 (N_8255,N_1653,N_2866);
or U8256 (N_8256,N_3849,N_4094);
nor U8257 (N_8257,N_4113,N_2188);
or U8258 (N_8258,N_2158,N_4791);
or U8259 (N_8259,N_3067,N_4786);
or U8260 (N_8260,N_4513,N_4107);
and U8261 (N_8261,N_1219,N_1491);
and U8262 (N_8262,N_4833,N_4518);
nor U8263 (N_8263,N_916,N_1628);
and U8264 (N_8264,N_4526,N_3441);
and U8265 (N_8265,N_279,N_784);
or U8266 (N_8266,N_4431,N_4803);
nor U8267 (N_8267,N_457,N_2759);
nand U8268 (N_8268,N_605,N_4724);
nand U8269 (N_8269,N_2699,N_1279);
nand U8270 (N_8270,N_1408,N_3362);
nor U8271 (N_8271,N_1397,N_1861);
and U8272 (N_8272,N_1593,N_4498);
nor U8273 (N_8273,N_4649,N_335);
nand U8274 (N_8274,N_4676,N_3713);
nor U8275 (N_8275,N_2564,N_4284);
nor U8276 (N_8276,N_3505,N_2283);
nor U8277 (N_8277,N_4439,N_1961);
or U8278 (N_8278,N_4456,N_3040);
nor U8279 (N_8279,N_617,N_2791);
or U8280 (N_8280,N_2051,N_1519);
xnor U8281 (N_8281,N_313,N_2823);
xnor U8282 (N_8282,N_1925,N_3716);
and U8283 (N_8283,N_1144,N_722);
nand U8284 (N_8284,N_4251,N_149);
and U8285 (N_8285,N_2081,N_2709);
or U8286 (N_8286,N_482,N_2140);
or U8287 (N_8287,N_1873,N_668);
and U8288 (N_8288,N_718,N_2631);
or U8289 (N_8289,N_3081,N_1471);
and U8290 (N_8290,N_2022,N_4016);
nand U8291 (N_8291,N_2454,N_4568);
or U8292 (N_8292,N_4425,N_1911);
nand U8293 (N_8293,N_387,N_4723);
nor U8294 (N_8294,N_2407,N_4941);
nand U8295 (N_8295,N_611,N_2264);
or U8296 (N_8296,N_4687,N_3247);
and U8297 (N_8297,N_650,N_193);
nor U8298 (N_8298,N_846,N_4270);
nor U8299 (N_8299,N_1550,N_2798);
or U8300 (N_8300,N_4285,N_458);
or U8301 (N_8301,N_603,N_4989);
and U8302 (N_8302,N_4898,N_1555);
or U8303 (N_8303,N_2667,N_3039);
and U8304 (N_8304,N_1718,N_1124);
nand U8305 (N_8305,N_4823,N_2541);
nand U8306 (N_8306,N_3215,N_3206);
nand U8307 (N_8307,N_2499,N_1364);
or U8308 (N_8308,N_3505,N_73);
nor U8309 (N_8309,N_4441,N_585);
nor U8310 (N_8310,N_3879,N_579);
nand U8311 (N_8311,N_1587,N_4962);
nor U8312 (N_8312,N_552,N_3468);
nor U8313 (N_8313,N_2232,N_509);
and U8314 (N_8314,N_4326,N_2580);
and U8315 (N_8315,N_4239,N_1037);
or U8316 (N_8316,N_1687,N_505);
or U8317 (N_8317,N_3406,N_3065);
and U8318 (N_8318,N_4163,N_571);
nand U8319 (N_8319,N_2399,N_956);
and U8320 (N_8320,N_784,N_2303);
and U8321 (N_8321,N_1350,N_2383);
nor U8322 (N_8322,N_3968,N_4876);
and U8323 (N_8323,N_1331,N_2697);
nor U8324 (N_8324,N_4385,N_4390);
nand U8325 (N_8325,N_2677,N_4001);
and U8326 (N_8326,N_608,N_1350);
nand U8327 (N_8327,N_1879,N_1513);
or U8328 (N_8328,N_4772,N_1493);
or U8329 (N_8329,N_4525,N_4081);
or U8330 (N_8330,N_3971,N_1821);
nand U8331 (N_8331,N_2469,N_4212);
or U8332 (N_8332,N_4092,N_3447);
or U8333 (N_8333,N_648,N_4609);
and U8334 (N_8334,N_2583,N_3065);
or U8335 (N_8335,N_3124,N_2392);
or U8336 (N_8336,N_70,N_2025);
and U8337 (N_8337,N_2936,N_2097);
nor U8338 (N_8338,N_437,N_3993);
nor U8339 (N_8339,N_469,N_1175);
nand U8340 (N_8340,N_4097,N_2341);
nor U8341 (N_8341,N_137,N_1896);
or U8342 (N_8342,N_648,N_2913);
nor U8343 (N_8343,N_1318,N_1426);
nand U8344 (N_8344,N_3057,N_2484);
nand U8345 (N_8345,N_4440,N_711);
nor U8346 (N_8346,N_1570,N_3801);
nor U8347 (N_8347,N_3245,N_4257);
nor U8348 (N_8348,N_887,N_359);
and U8349 (N_8349,N_3220,N_708);
nor U8350 (N_8350,N_2614,N_3166);
nand U8351 (N_8351,N_309,N_6);
nand U8352 (N_8352,N_91,N_214);
nand U8353 (N_8353,N_2278,N_4601);
and U8354 (N_8354,N_1418,N_541);
and U8355 (N_8355,N_2975,N_3967);
nand U8356 (N_8356,N_4081,N_1721);
nand U8357 (N_8357,N_2099,N_822);
nor U8358 (N_8358,N_2765,N_4036);
nor U8359 (N_8359,N_1086,N_1706);
nand U8360 (N_8360,N_659,N_723);
or U8361 (N_8361,N_3006,N_3092);
nand U8362 (N_8362,N_3339,N_4694);
and U8363 (N_8363,N_1865,N_4691);
nor U8364 (N_8364,N_546,N_4291);
or U8365 (N_8365,N_1330,N_367);
or U8366 (N_8366,N_1300,N_2317);
or U8367 (N_8367,N_2356,N_2096);
nor U8368 (N_8368,N_409,N_2969);
or U8369 (N_8369,N_3200,N_548);
or U8370 (N_8370,N_1187,N_1555);
nor U8371 (N_8371,N_3697,N_1544);
nand U8372 (N_8372,N_2214,N_1690);
xnor U8373 (N_8373,N_367,N_72);
and U8374 (N_8374,N_3984,N_3490);
and U8375 (N_8375,N_4378,N_4372);
or U8376 (N_8376,N_1745,N_1255);
or U8377 (N_8377,N_4681,N_2104);
nand U8378 (N_8378,N_988,N_4305);
and U8379 (N_8379,N_4952,N_2245);
nand U8380 (N_8380,N_2717,N_1994);
nand U8381 (N_8381,N_4861,N_3726);
xnor U8382 (N_8382,N_3439,N_4917);
and U8383 (N_8383,N_555,N_3757);
nand U8384 (N_8384,N_4142,N_1468);
xnor U8385 (N_8385,N_3117,N_3514);
or U8386 (N_8386,N_944,N_1146);
or U8387 (N_8387,N_1590,N_1705);
nor U8388 (N_8388,N_351,N_1641);
and U8389 (N_8389,N_4129,N_3178);
or U8390 (N_8390,N_2529,N_3694);
and U8391 (N_8391,N_2569,N_1428);
nor U8392 (N_8392,N_3221,N_4600);
nor U8393 (N_8393,N_2120,N_833);
nor U8394 (N_8394,N_2333,N_350);
nor U8395 (N_8395,N_1617,N_4835);
and U8396 (N_8396,N_802,N_3904);
nand U8397 (N_8397,N_1607,N_2374);
nand U8398 (N_8398,N_4667,N_3813);
nor U8399 (N_8399,N_3727,N_4994);
and U8400 (N_8400,N_4341,N_3324);
nor U8401 (N_8401,N_2655,N_3529);
nand U8402 (N_8402,N_4382,N_1652);
and U8403 (N_8403,N_2482,N_2030);
nor U8404 (N_8404,N_3864,N_983);
or U8405 (N_8405,N_37,N_4247);
nand U8406 (N_8406,N_2796,N_3377);
and U8407 (N_8407,N_983,N_1722);
nand U8408 (N_8408,N_1171,N_4725);
nor U8409 (N_8409,N_2055,N_531);
and U8410 (N_8410,N_4099,N_3892);
or U8411 (N_8411,N_4259,N_2257);
nor U8412 (N_8412,N_1265,N_4676);
or U8413 (N_8413,N_859,N_2649);
or U8414 (N_8414,N_3527,N_1197);
and U8415 (N_8415,N_2581,N_1040);
nor U8416 (N_8416,N_1290,N_2057);
and U8417 (N_8417,N_1521,N_946);
xnor U8418 (N_8418,N_1317,N_3169);
nand U8419 (N_8419,N_2287,N_4519);
nor U8420 (N_8420,N_2792,N_1906);
or U8421 (N_8421,N_454,N_198);
nor U8422 (N_8422,N_3246,N_4502);
or U8423 (N_8423,N_4644,N_1638);
nand U8424 (N_8424,N_3964,N_4855);
nor U8425 (N_8425,N_2932,N_26);
nor U8426 (N_8426,N_2760,N_1373);
or U8427 (N_8427,N_1388,N_427);
or U8428 (N_8428,N_4823,N_3855);
nand U8429 (N_8429,N_2049,N_4667);
or U8430 (N_8430,N_1130,N_7);
nor U8431 (N_8431,N_2416,N_4331);
and U8432 (N_8432,N_278,N_1303);
nand U8433 (N_8433,N_2502,N_723);
nand U8434 (N_8434,N_1531,N_3856);
or U8435 (N_8435,N_1301,N_3337);
and U8436 (N_8436,N_2401,N_2441);
nand U8437 (N_8437,N_493,N_1428);
and U8438 (N_8438,N_2475,N_2426);
and U8439 (N_8439,N_4250,N_434);
nand U8440 (N_8440,N_4940,N_4708);
nor U8441 (N_8441,N_1136,N_1893);
and U8442 (N_8442,N_3634,N_777);
nor U8443 (N_8443,N_2044,N_4074);
nand U8444 (N_8444,N_1911,N_128);
nand U8445 (N_8445,N_3198,N_2853);
nand U8446 (N_8446,N_2281,N_2169);
xor U8447 (N_8447,N_1607,N_4161);
nand U8448 (N_8448,N_2898,N_3622);
and U8449 (N_8449,N_4282,N_836);
and U8450 (N_8450,N_2261,N_2227);
nor U8451 (N_8451,N_1090,N_4485);
or U8452 (N_8452,N_2472,N_3441);
nand U8453 (N_8453,N_2487,N_1619);
and U8454 (N_8454,N_3314,N_1672);
or U8455 (N_8455,N_322,N_2190);
nor U8456 (N_8456,N_2582,N_1711);
and U8457 (N_8457,N_292,N_2198);
and U8458 (N_8458,N_69,N_2739);
or U8459 (N_8459,N_3420,N_443);
or U8460 (N_8460,N_704,N_4316);
and U8461 (N_8461,N_1188,N_2493);
nor U8462 (N_8462,N_4094,N_11);
nor U8463 (N_8463,N_4574,N_1734);
and U8464 (N_8464,N_4134,N_2439);
nand U8465 (N_8465,N_954,N_1402);
nor U8466 (N_8466,N_3768,N_2131);
and U8467 (N_8467,N_2085,N_110);
nor U8468 (N_8468,N_1237,N_3943);
or U8469 (N_8469,N_1160,N_1635);
nor U8470 (N_8470,N_3049,N_998);
nor U8471 (N_8471,N_2286,N_2190);
nand U8472 (N_8472,N_4837,N_20);
nand U8473 (N_8473,N_3860,N_1937);
and U8474 (N_8474,N_4111,N_2559);
or U8475 (N_8475,N_2733,N_1369);
nor U8476 (N_8476,N_3740,N_78);
xor U8477 (N_8477,N_1893,N_4355);
and U8478 (N_8478,N_4640,N_523);
or U8479 (N_8479,N_4861,N_1723);
nor U8480 (N_8480,N_4371,N_337);
and U8481 (N_8481,N_3779,N_1938);
nand U8482 (N_8482,N_3440,N_4333);
or U8483 (N_8483,N_4120,N_4261);
nand U8484 (N_8484,N_3819,N_1648);
nand U8485 (N_8485,N_3813,N_3398);
or U8486 (N_8486,N_4421,N_3526);
or U8487 (N_8487,N_702,N_376);
nand U8488 (N_8488,N_3904,N_4334);
nor U8489 (N_8489,N_2234,N_245);
or U8490 (N_8490,N_2550,N_2426);
and U8491 (N_8491,N_4598,N_1144);
and U8492 (N_8492,N_3329,N_1502);
and U8493 (N_8493,N_3214,N_252);
and U8494 (N_8494,N_3294,N_1685);
and U8495 (N_8495,N_387,N_1838);
nand U8496 (N_8496,N_3549,N_4509);
or U8497 (N_8497,N_3459,N_3664);
and U8498 (N_8498,N_4963,N_4937);
nand U8499 (N_8499,N_1493,N_1567);
and U8500 (N_8500,N_2820,N_3451);
and U8501 (N_8501,N_951,N_3880);
nand U8502 (N_8502,N_461,N_1358);
and U8503 (N_8503,N_4077,N_2950);
nor U8504 (N_8504,N_22,N_4373);
and U8505 (N_8505,N_370,N_879);
nand U8506 (N_8506,N_330,N_4813);
nand U8507 (N_8507,N_4530,N_4932);
or U8508 (N_8508,N_3850,N_2868);
nand U8509 (N_8509,N_3021,N_1387);
and U8510 (N_8510,N_3520,N_1562);
nor U8511 (N_8511,N_3956,N_4197);
nand U8512 (N_8512,N_3047,N_2051);
and U8513 (N_8513,N_4541,N_711);
nor U8514 (N_8514,N_2684,N_852);
nand U8515 (N_8515,N_2355,N_2935);
nand U8516 (N_8516,N_151,N_1043);
and U8517 (N_8517,N_998,N_840);
nand U8518 (N_8518,N_4689,N_4584);
and U8519 (N_8519,N_1273,N_4551);
nand U8520 (N_8520,N_4298,N_3774);
nand U8521 (N_8521,N_220,N_1177);
or U8522 (N_8522,N_3195,N_1015);
and U8523 (N_8523,N_4834,N_3884);
or U8524 (N_8524,N_2744,N_1740);
and U8525 (N_8525,N_2000,N_577);
nand U8526 (N_8526,N_4456,N_3249);
nor U8527 (N_8527,N_2995,N_2945);
or U8528 (N_8528,N_4111,N_3497);
nand U8529 (N_8529,N_3981,N_2117);
and U8530 (N_8530,N_2992,N_3264);
nor U8531 (N_8531,N_62,N_913);
or U8532 (N_8532,N_4444,N_998);
nor U8533 (N_8533,N_590,N_739);
nor U8534 (N_8534,N_3075,N_1560);
nor U8535 (N_8535,N_4351,N_257);
nand U8536 (N_8536,N_2553,N_3665);
or U8537 (N_8537,N_2626,N_388);
or U8538 (N_8538,N_4160,N_2384);
and U8539 (N_8539,N_3546,N_1831);
or U8540 (N_8540,N_2714,N_924);
nand U8541 (N_8541,N_3225,N_4887);
nor U8542 (N_8542,N_3336,N_570);
xor U8543 (N_8543,N_1931,N_3576);
nor U8544 (N_8544,N_345,N_2502);
or U8545 (N_8545,N_314,N_4537);
or U8546 (N_8546,N_782,N_3296);
and U8547 (N_8547,N_599,N_2577);
nor U8548 (N_8548,N_2807,N_459);
or U8549 (N_8549,N_3016,N_2321);
and U8550 (N_8550,N_37,N_2756);
or U8551 (N_8551,N_3455,N_2411);
nand U8552 (N_8552,N_1477,N_4197);
and U8553 (N_8553,N_4845,N_4267);
or U8554 (N_8554,N_872,N_4895);
or U8555 (N_8555,N_289,N_599);
or U8556 (N_8556,N_3526,N_3029);
and U8557 (N_8557,N_777,N_4547);
or U8558 (N_8558,N_49,N_458);
nor U8559 (N_8559,N_2022,N_13);
nor U8560 (N_8560,N_2212,N_1911);
or U8561 (N_8561,N_2879,N_3418);
and U8562 (N_8562,N_2677,N_4254);
or U8563 (N_8563,N_1487,N_4817);
and U8564 (N_8564,N_3991,N_2322);
nor U8565 (N_8565,N_2277,N_3140);
nand U8566 (N_8566,N_3986,N_3230);
nor U8567 (N_8567,N_2920,N_4037);
nand U8568 (N_8568,N_4622,N_4530);
or U8569 (N_8569,N_4089,N_1599);
and U8570 (N_8570,N_1452,N_3210);
and U8571 (N_8571,N_1526,N_1574);
and U8572 (N_8572,N_520,N_1220);
nor U8573 (N_8573,N_2976,N_2263);
nand U8574 (N_8574,N_2676,N_4930);
or U8575 (N_8575,N_3360,N_2696);
nand U8576 (N_8576,N_2448,N_3420);
nor U8577 (N_8577,N_2003,N_228);
or U8578 (N_8578,N_4517,N_1250);
nand U8579 (N_8579,N_3167,N_3275);
and U8580 (N_8580,N_1749,N_2984);
or U8581 (N_8581,N_1599,N_429);
nand U8582 (N_8582,N_1440,N_1314);
nor U8583 (N_8583,N_862,N_638);
or U8584 (N_8584,N_61,N_4650);
or U8585 (N_8585,N_1173,N_1439);
and U8586 (N_8586,N_3411,N_3373);
nand U8587 (N_8587,N_3509,N_786);
or U8588 (N_8588,N_1558,N_4059);
and U8589 (N_8589,N_2622,N_4151);
and U8590 (N_8590,N_2472,N_4813);
and U8591 (N_8591,N_3410,N_2148);
nor U8592 (N_8592,N_4937,N_4379);
nor U8593 (N_8593,N_1357,N_3840);
nor U8594 (N_8594,N_3893,N_3340);
nand U8595 (N_8595,N_3675,N_2104);
nand U8596 (N_8596,N_4102,N_1336);
nand U8597 (N_8597,N_2331,N_4783);
or U8598 (N_8598,N_222,N_4031);
nor U8599 (N_8599,N_2458,N_2131);
nand U8600 (N_8600,N_2085,N_4777);
or U8601 (N_8601,N_3309,N_343);
xnor U8602 (N_8602,N_2514,N_496);
nand U8603 (N_8603,N_1409,N_4063);
or U8604 (N_8604,N_3042,N_3149);
or U8605 (N_8605,N_3473,N_3847);
nand U8606 (N_8606,N_3986,N_3924);
nor U8607 (N_8607,N_2526,N_4251);
or U8608 (N_8608,N_1551,N_2937);
nor U8609 (N_8609,N_1907,N_2181);
nand U8610 (N_8610,N_4717,N_1452);
nand U8611 (N_8611,N_2087,N_3566);
or U8612 (N_8612,N_2082,N_3918);
xnor U8613 (N_8613,N_1007,N_4661);
nor U8614 (N_8614,N_997,N_3403);
and U8615 (N_8615,N_1300,N_3803);
xor U8616 (N_8616,N_1414,N_1988);
nor U8617 (N_8617,N_2693,N_1058);
nand U8618 (N_8618,N_4709,N_912);
nor U8619 (N_8619,N_2808,N_4793);
or U8620 (N_8620,N_1668,N_4458);
xnor U8621 (N_8621,N_3076,N_2503);
nand U8622 (N_8622,N_1844,N_1037);
and U8623 (N_8623,N_1637,N_485);
and U8624 (N_8624,N_2204,N_3076);
nor U8625 (N_8625,N_142,N_2664);
nand U8626 (N_8626,N_4322,N_1145);
or U8627 (N_8627,N_2467,N_3231);
nand U8628 (N_8628,N_615,N_3025);
and U8629 (N_8629,N_2751,N_2576);
or U8630 (N_8630,N_4671,N_564);
or U8631 (N_8631,N_4000,N_4640);
nor U8632 (N_8632,N_1982,N_3793);
nor U8633 (N_8633,N_4013,N_4545);
or U8634 (N_8634,N_2388,N_2727);
or U8635 (N_8635,N_4343,N_3181);
nor U8636 (N_8636,N_177,N_3501);
nand U8637 (N_8637,N_1708,N_3934);
and U8638 (N_8638,N_3148,N_2289);
or U8639 (N_8639,N_3558,N_390);
and U8640 (N_8640,N_3560,N_343);
nand U8641 (N_8641,N_339,N_354);
and U8642 (N_8642,N_1582,N_55);
nand U8643 (N_8643,N_2771,N_2736);
or U8644 (N_8644,N_886,N_1892);
and U8645 (N_8645,N_1546,N_514);
nor U8646 (N_8646,N_3467,N_2681);
nand U8647 (N_8647,N_1720,N_1634);
nor U8648 (N_8648,N_3904,N_3096);
nor U8649 (N_8649,N_2952,N_774);
nand U8650 (N_8650,N_2430,N_1284);
or U8651 (N_8651,N_3084,N_4951);
and U8652 (N_8652,N_2848,N_4575);
xnor U8653 (N_8653,N_4890,N_2904);
or U8654 (N_8654,N_3924,N_1269);
and U8655 (N_8655,N_4194,N_1926);
nor U8656 (N_8656,N_1686,N_3827);
and U8657 (N_8657,N_3038,N_2745);
nor U8658 (N_8658,N_471,N_891);
and U8659 (N_8659,N_1022,N_2329);
nand U8660 (N_8660,N_4498,N_1221);
nand U8661 (N_8661,N_1623,N_1985);
nor U8662 (N_8662,N_1673,N_1558);
and U8663 (N_8663,N_3298,N_3806);
or U8664 (N_8664,N_997,N_1234);
nor U8665 (N_8665,N_3901,N_1269);
or U8666 (N_8666,N_2571,N_507);
or U8667 (N_8667,N_75,N_1553);
nand U8668 (N_8668,N_2671,N_635);
nand U8669 (N_8669,N_2023,N_3795);
or U8670 (N_8670,N_4487,N_3905);
nor U8671 (N_8671,N_2559,N_4691);
and U8672 (N_8672,N_4240,N_3445);
and U8673 (N_8673,N_2752,N_4742);
nor U8674 (N_8674,N_489,N_4310);
or U8675 (N_8675,N_4067,N_1101);
nand U8676 (N_8676,N_514,N_709);
or U8677 (N_8677,N_2317,N_3732);
or U8678 (N_8678,N_3049,N_2779);
nand U8679 (N_8679,N_2243,N_1916);
xor U8680 (N_8680,N_2799,N_4249);
nor U8681 (N_8681,N_2217,N_3431);
nand U8682 (N_8682,N_4343,N_2370);
nor U8683 (N_8683,N_4190,N_1662);
nand U8684 (N_8684,N_2581,N_4525);
or U8685 (N_8685,N_2381,N_3301);
or U8686 (N_8686,N_1795,N_4677);
or U8687 (N_8687,N_678,N_2750);
xor U8688 (N_8688,N_1448,N_3285);
or U8689 (N_8689,N_1992,N_2177);
nand U8690 (N_8690,N_2918,N_2702);
and U8691 (N_8691,N_3912,N_172);
xnor U8692 (N_8692,N_4722,N_3939);
nand U8693 (N_8693,N_4372,N_3895);
nor U8694 (N_8694,N_1752,N_2952);
or U8695 (N_8695,N_3376,N_563);
nor U8696 (N_8696,N_3657,N_4110);
or U8697 (N_8697,N_795,N_3926);
nand U8698 (N_8698,N_3926,N_1392);
nor U8699 (N_8699,N_3931,N_4794);
nand U8700 (N_8700,N_1999,N_1160);
nand U8701 (N_8701,N_3932,N_4250);
and U8702 (N_8702,N_4346,N_4247);
nor U8703 (N_8703,N_2852,N_52);
or U8704 (N_8704,N_2231,N_2909);
or U8705 (N_8705,N_2810,N_2232);
and U8706 (N_8706,N_734,N_2567);
or U8707 (N_8707,N_2150,N_2823);
and U8708 (N_8708,N_2191,N_4846);
nor U8709 (N_8709,N_3689,N_4589);
nand U8710 (N_8710,N_2765,N_1155);
nand U8711 (N_8711,N_3950,N_4632);
xor U8712 (N_8712,N_2278,N_1304);
nor U8713 (N_8713,N_1551,N_1982);
nor U8714 (N_8714,N_3061,N_169);
nand U8715 (N_8715,N_2496,N_3353);
nor U8716 (N_8716,N_2670,N_1480);
nor U8717 (N_8717,N_2436,N_4196);
nor U8718 (N_8718,N_3278,N_4586);
or U8719 (N_8719,N_1823,N_3593);
nor U8720 (N_8720,N_2507,N_724);
or U8721 (N_8721,N_542,N_2539);
nand U8722 (N_8722,N_1168,N_3253);
nand U8723 (N_8723,N_1800,N_2358);
nand U8724 (N_8724,N_818,N_3222);
nor U8725 (N_8725,N_3399,N_2341);
nor U8726 (N_8726,N_1323,N_1494);
nor U8727 (N_8727,N_4361,N_4946);
or U8728 (N_8728,N_3830,N_2526);
nand U8729 (N_8729,N_3935,N_655);
nand U8730 (N_8730,N_4875,N_1510);
nand U8731 (N_8731,N_3901,N_2729);
or U8732 (N_8732,N_3543,N_2727);
and U8733 (N_8733,N_1003,N_4562);
nor U8734 (N_8734,N_840,N_2632);
nor U8735 (N_8735,N_1377,N_2968);
or U8736 (N_8736,N_2769,N_3428);
or U8737 (N_8737,N_44,N_4280);
nand U8738 (N_8738,N_944,N_1917);
nand U8739 (N_8739,N_448,N_3538);
nor U8740 (N_8740,N_3960,N_964);
nor U8741 (N_8741,N_3719,N_4880);
or U8742 (N_8742,N_3987,N_4182);
nor U8743 (N_8743,N_919,N_3653);
or U8744 (N_8744,N_1005,N_1163);
nand U8745 (N_8745,N_2609,N_889);
or U8746 (N_8746,N_581,N_2157);
or U8747 (N_8747,N_4828,N_2585);
nand U8748 (N_8748,N_4625,N_4150);
nor U8749 (N_8749,N_713,N_2927);
or U8750 (N_8750,N_4823,N_882);
and U8751 (N_8751,N_4120,N_2881);
xor U8752 (N_8752,N_4921,N_703);
and U8753 (N_8753,N_3939,N_4738);
or U8754 (N_8754,N_163,N_3719);
or U8755 (N_8755,N_4207,N_1543);
nand U8756 (N_8756,N_3311,N_2179);
or U8757 (N_8757,N_4659,N_367);
and U8758 (N_8758,N_4927,N_1301);
nor U8759 (N_8759,N_1963,N_197);
nand U8760 (N_8760,N_76,N_3605);
and U8761 (N_8761,N_3866,N_4804);
nand U8762 (N_8762,N_4519,N_1611);
or U8763 (N_8763,N_840,N_2067);
xor U8764 (N_8764,N_4214,N_3518);
or U8765 (N_8765,N_120,N_4484);
nor U8766 (N_8766,N_572,N_4242);
nor U8767 (N_8767,N_2532,N_4259);
nor U8768 (N_8768,N_2243,N_4454);
or U8769 (N_8769,N_82,N_3541);
and U8770 (N_8770,N_540,N_4945);
nand U8771 (N_8771,N_804,N_1290);
or U8772 (N_8772,N_406,N_2672);
and U8773 (N_8773,N_680,N_140);
nand U8774 (N_8774,N_4432,N_550);
nor U8775 (N_8775,N_4574,N_2034);
nor U8776 (N_8776,N_2434,N_2021);
or U8777 (N_8777,N_3460,N_918);
or U8778 (N_8778,N_635,N_2462);
nand U8779 (N_8779,N_4809,N_4211);
nand U8780 (N_8780,N_4903,N_489);
or U8781 (N_8781,N_55,N_4980);
nor U8782 (N_8782,N_683,N_785);
or U8783 (N_8783,N_1845,N_3347);
and U8784 (N_8784,N_2607,N_1730);
and U8785 (N_8785,N_1462,N_1124);
or U8786 (N_8786,N_893,N_1472);
or U8787 (N_8787,N_70,N_447);
nor U8788 (N_8788,N_1187,N_4156);
nor U8789 (N_8789,N_1520,N_1585);
nand U8790 (N_8790,N_4491,N_1971);
nor U8791 (N_8791,N_1798,N_700);
xor U8792 (N_8792,N_2755,N_3030);
nor U8793 (N_8793,N_2027,N_4876);
and U8794 (N_8794,N_1266,N_4352);
nor U8795 (N_8795,N_1126,N_2548);
nor U8796 (N_8796,N_4027,N_3499);
nor U8797 (N_8797,N_3264,N_3141);
nor U8798 (N_8798,N_1803,N_619);
nand U8799 (N_8799,N_830,N_4655);
or U8800 (N_8800,N_609,N_4256);
and U8801 (N_8801,N_2863,N_2927);
or U8802 (N_8802,N_3778,N_43);
and U8803 (N_8803,N_1050,N_2976);
nand U8804 (N_8804,N_1330,N_1871);
nor U8805 (N_8805,N_662,N_3784);
and U8806 (N_8806,N_564,N_3877);
and U8807 (N_8807,N_1719,N_4927);
and U8808 (N_8808,N_224,N_382);
nor U8809 (N_8809,N_2414,N_459);
nand U8810 (N_8810,N_4623,N_2809);
nor U8811 (N_8811,N_483,N_1605);
nand U8812 (N_8812,N_3236,N_1205);
and U8813 (N_8813,N_665,N_3951);
or U8814 (N_8814,N_3576,N_976);
nor U8815 (N_8815,N_462,N_1402);
nor U8816 (N_8816,N_1677,N_3843);
nand U8817 (N_8817,N_148,N_58);
nor U8818 (N_8818,N_2345,N_2729);
and U8819 (N_8819,N_384,N_1291);
nor U8820 (N_8820,N_1369,N_1948);
and U8821 (N_8821,N_2726,N_256);
nor U8822 (N_8822,N_2662,N_1942);
nand U8823 (N_8823,N_3986,N_3242);
nand U8824 (N_8824,N_2728,N_3262);
or U8825 (N_8825,N_511,N_1776);
nor U8826 (N_8826,N_4594,N_2262);
or U8827 (N_8827,N_1987,N_2417);
or U8828 (N_8828,N_182,N_1251);
and U8829 (N_8829,N_1530,N_3999);
and U8830 (N_8830,N_1115,N_2578);
nor U8831 (N_8831,N_3983,N_1206);
nand U8832 (N_8832,N_3100,N_1034);
nor U8833 (N_8833,N_2192,N_1087);
nor U8834 (N_8834,N_4337,N_3867);
nor U8835 (N_8835,N_1062,N_4182);
nand U8836 (N_8836,N_38,N_2889);
nand U8837 (N_8837,N_3780,N_4899);
nand U8838 (N_8838,N_648,N_2530);
or U8839 (N_8839,N_254,N_409);
and U8840 (N_8840,N_963,N_3405);
nor U8841 (N_8841,N_2906,N_1592);
and U8842 (N_8842,N_834,N_192);
nand U8843 (N_8843,N_3796,N_3827);
and U8844 (N_8844,N_4061,N_4089);
or U8845 (N_8845,N_1731,N_1073);
nor U8846 (N_8846,N_1773,N_1561);
nand U8847 (N_8847,N_4065,N_1291);
nand U8848 (N_8848,N_97,N_1067);
nand U8849 (N_8849,N_2356,N_1593);
or U8850 (N_8850,N_3741,N_3093);
nor U8851 (N_8851,N_3025,N_2289);
and U8852 (N_8852,N_1618,N_1747);
nor U8853 (N_8853,N_3136,N_3414);
nand U8854 (N_8854,N_4560,N_3274);
or U8855 (N_8855,N_3015,N_2875);
or U8856 (N_8856,N_2559,N_3875);
or U8857 (N_8857,N_2736,N_2861);
and U8858 (N_8858,N_1061,N_4181);
or U8859 (N_8859,N_1979,N_985);
nor U8860 (N_8860,N_696,N_3955);
nor U8861 (N_8861,N_3846,N_3865);
and U8862 (N_8862,N_2756,N_2645);
nor U8863 (N_8863,N_1129,N_1364);
nor U8864 (N_8864,N_1384,N_2813);
and U8865 (N_8865,N_2691,N_4934);
or U8866 (N_8866,N_4563,N_1226);
xnor U8867 (N_8867,N_3863,N_3638);
nand U8868 (N_8868,N_1632,N_4014);
nor U8869 (N_8869,N_1534,N_4642);
or U8870 (N_8870,N_4190,N_3136);
nand U8871 (N_8871,N_3333,N_3438);
nor U8872 (N_8872,N_1147,N_2203);
or U8873 (N_8873,N_2841,N_3605);
or U8874 (N_8874,N_910,N_1187);
nand U8875 (N_8875,N_4855,N_2241);
or U8876 (N_8876,N_3688,N_2381);
nor U8877 (N_8877,N_1358,N_738);
or U8878 (N_8878,N_38,N_2119);
or U8879 (N_8879,N_1730,N_347);
and U8880 (N_8880,N_4563,N_4935);
nand U8881 (N_8881,N_2679,N_3078);
and U8882 (N_8882,N_2319,N_796);
nor U8883 (N_8883,N_2560,N_3703);
and U8884 (N_8884,N_1582,N_848);
and U8885 (N_8885,N_3826,N_1059);
or U8886 (N_8886,N_673,N_1074);
or U8887 (N_8887,N_1940,N_289);
xor U8888 (N_8888,N_1550,N_157);
nor U8889 (N_8889,N_2548,N_2807);
nor U8890 (N_8890,N_4710,N_3260);
or U8891 (N_8891,N_4507,N_3944);
nor U8892 (N_8892,N_4918,N_3539);
xnor U8893 (N_8893,N_3088,N_678);
or U8894 (N_8894,N_260,N_795);
nand U8895 (N_8895,N_588,N_2533);
xor U8896 (N_8896,N_567,N_864);
nand U8897 (N_8897,N_1003,N_513);
xnor U8898 (N_8898,N_3972,N_1344);
nand U8899 (N_8899,N_3827,N_3752);
nor U8900 (N_8900,N_4289,N_4140);
and U8901 (N_8901,N_735,N_439);
nor U8902 (N_8902,N_1008,N_84);
or U8903 (N_8903,N_4247,N_352);
nand U8904 (N_8904,N_3346,N_582);
or U8905 (N_8905,N_4112,N_3762);
and U8906 (N_8906,N_2576,N_1378);
nor U8907 (N_8907,N_1398,N_3024);
or U8908 (N_8908,N_160,N_4491);
nor U8909 (N_8909,N_2468,N_739);
and U8910 (N_8910,N_507,N_2141);
and U8911 (N_8911,N_4030,N_4920);
nor U8912 (N_8912,N_1903,N_2571);
or U8913 (N_8913,N_2794,N_4148);
nand U8914 (N_8914,N_284,N_2001);
nor U8915 (N_8915,N_2136,N_491);
nor U8916 (N_8916,N_4608,N_1177);
nand U8917 (N_8917,N_2233,N_3714);
and U8918 (N_8918,N_1053,N_4150);
nor U8919 (N_8919,N_1345,N_3308);
or U8920 (N_8920,N_2285,N_2458);
and U8921 (N_8921,N_2879,N_602);
nor U8922 (N_8922,N_2774,N_903);
nor U8923 (N_8923,N_4033,N_1369);
and U8924 (N_8924,N_3940,N_3796);
nor U8925 (N_8925,N_22,N_4489);
nand U8926 (N_8926,N_1032,N_1731);
nor U8927 (N_8927,N_2266,N_820);
nand U8928 (N_8928,N_1938,N_3689);
nand U8929 (N_8929,N_2951,N_3364);
and U8930 (N_8930,N_4086,N_2335);
nand U8931 (N_8931,N_1639,N_2597);
or U8932 (N_8932,N_4802,N_920);
nor U8933 (N_8933,N_4592,N_579);
and U8934 (N_8934,N_4782,N_475);
xor U8935 (N_8935,N_2718,N_2130);
nor U8936 (N_8936,N_4365,N_246);
nand U8937 (N_8937,N_3063,N_4436);
or U8938 (N_8938,N_4847,N_1521);
nand U8939 (N_8939,N_2481,N_1382);
and U8940 (N_8940,N_4767,N_187);
nand U8941 (N_8941,N_3272,N_4555);
nor U8942 (N_8942,N_2017,N_4501);
or U8943 (N_8943,N_3118,N_3430);
nand U8944 (N_8944,N_2662,N_723);
nand U8945 (N_8945,N_3294,N_1074);
nor U8946 (N_8946,N_4506,N_1945);
nor U8947 (N_8947,N_3480,N_3014);
or U8948 (N_8948,N_4096,N_3904);
nand U8949 (N_8949,N_4807,N_1806);
nand U8950 (N_8950,N_2318,N_150);
nor U8951 (N_8951,N_132,N_3822);
and U8952 (N_8952,N_1568,N_2243);
xnor U8953 (N_8953,N_3817,N_1584);
nor U8954 (N_8954,N_1926,N_4901);
or U8955 (N_8955,N_3680,N_3736);
and U8956 (N_8956,N_3864,N_2222);
or U8957 (N_8957,N_3315,N_4106);
and U8958 (N_8958,N_1422,N_3044);
or U8959 (N_8959,N_4849,N_4772);
nor U8960 (N_8960,N_3370,N_2756);
and U8961 (N_8961,N_238,N_4565);
nor U8962 (N_8962,N_1158,N_4680);
or U8963 (N_8963,N_459,N_1626);
nor U8964 (N_8964,N_683,N_585);
or U8965 (N_8965,N_4680,N_4983);
and U8966 (N_8966,N_209,N_1925);
or U8967 (N_8967,N_4006,N_3247);
nand U8968 (N_8968,N_752,N_4307);
nor U8969 (N_8969,N_4556,N_4858);
xor U8970 (N_8970,N_876,N_1207);
xor U8971 (N_8971,N_1564,N_1602);
and U8972 (N_8972,N_1176,N_2672);
or U8973 (N_8973,N_107,N_309);
or U8974 (N_8974,N_4605,N_151);
nor U8975 (N_8975,N_1789,N_3644);
nor U8976 (N_8976,N_3904,N_2460);
nor U8977 (N_8977,N_3360,N_2968);
nor U8978 (N_8978,N_861,N_2273);
or U8979 (N_8979,N_3494,N_1904);
nand U8980 (N_8980,N_423,N_2055);
nor U8981 (N_8981,N_3021,N_1614);
or U8982 (N_8982,N_219,N_954);
and U8983 (N_8983,N_1546,N_577);
nand U8984 (N_8984,N_570,N_2225);
nand U8985 (N_8985,N_2366,N_2257);
nand U8986 (N_8986,N_3902,N_2860);
nand U8987 (N_8987,N_4789,N_1623);
and U8988 (N_8988,N_2074,N_3733);
nand U8989 (N_8989,N_881,N_3619);
nor U8990 (N_8990,N_2650,N_1414);
nor U8991 (N_8991,N_138,N_489);
or U8992 (N_8992,N_1218,N_2592);
and U8993 (N_8993,N_3212,N_1096);
nand U8994 (N_8994,N_1521,N_2457);
or U8995 (N_8995,N_3498,N_70);
nand U8996 (N_8996,N_4039,N_2595);
and U8997 (N_8997,N_2885,N_445);
and U8998 (N_8998,N_3018,N_3168);
nor U8999 (N_8999,N_4238,N_4961);
nor U9000 (N_9000,N_2875,N_374);
nand U9001 (N_9001,N_4137,N_1623);
xnor U9002 (N_9002,N_1945,N_2974);
nand U9003 (N_9003,N_3637,N_778);
nor U9004 (N_9004,N_1794,N_615);
xnor U9005 (N_9005,N_3114,N_2924);
or U9006 (N_9006,N_3074,N_317);
and U9007 (N_9007,N_1235,N_1386);
nor U9008 (N_9008,N_344,N_412);
nor U9009 (N_9009,N_707,N_4757);
nor U9010 (N_9010,N_1615,N_4312);
and U9011 (N_9011,N_3439,N_2847);
nand U9012 (N_9012,N_272,N_172);
or U9013 (N_9013,N_452,N_2371);
nand U9014 (N_9014,N_4270,N_1340);
and U9015 (N_9015,N_2512,N_1977);
nand U9016 (N_9016,N_4546,N_3582);
nand U9017 (N_9017,N_4508,N_232);
nand U9018 (N_9018,N_629,N_2358);
and U9019 (N_9019,N_514,N_147);
and U9020 (N_9020,N_4732,N_3229);
or U9021 (N_9021,N_4320,N_3092);
or U9022 (N_9022,N_1680,N_4749);
xnor U9023 (N_9023,N_3217,N_2461);
and U9024 (N_9024,N_3919,N_58);
nand U9025 (N_9025,N_2980,N_3224);
nor U9026 (N_9026,N_3102,N_1332);
nand U9027 (N_9027,N_1106,N_3518);
or U9028 (N_9028,N_2668,N_4400);
and U9029 (N_9029,N_709,N_2647);
nand U9030 (N_9030,N_3341,N_2444);
nand U9031 (N_9031,N_3609,N_1231);
nor U9032 (N_9032,N_794,N_1500);
xnor U9033 (N_9033,N_4726,N_4849);
nor U9034 (N_9034,N_3856,N_1370);
or U9035 (N_9035,N_2161,N_146);
or U9036 (N_9036,N_3371,N_4456);
and U9037 (N_9037,N_2428,N_4202);
nand U9038 (N_9038,N_3864,N_2834);
and U9039 (N_9039,N_2938,N_2117);
or U9040 (N_9040,N_256,N_849);
and U9041 (N_9041,N_2933,N_4385);
nand U9042 (N_9042,N_4297,N_535);
nand U9043 (N_9043,N_266,N_4178);
nor U9044 (N_9044,N_4209,N_3099);
and U9045 (N_9045,N_4362,N_45);
nor U9046 (N_9046,N_3635,N_174);
or U9047 (N_9047,N_2991,N_1266);
or U9048 (N_9048,N_818,N_1313);
nand U9049 (N_9049,N_4928,N_4862);
or U9050 (N_9050,N_3490,N_4973);
and U9051 (N_9051,N_4386,N_3740);
and U9052 (N_9052,N_2899,N_3169);
nand U9053 (N_9053,N_2153,N_1213);
and U9054 (N_9054,N_563,N_3159);
nor U9055 (N_9055,N_3528,N_1027);
nand U9056 (N_9056,N_4167,N_2893);
and U9057 (N_9057,N_688,N_3799);
or U9058 (N_9058,N_3226,N_2415);
and U9059 (N_9059,N_1741,N_3270);
nor U9060 (N_9060,N_3120,N_1161);
nand U9061 (N_9061,N_2889,N_2510);
or U9062 (N_9062,N_3593,N_3304);
nand U9063 (N_9063,N_3491,N_1065);
or U9064 (N_9064,N_1859,N_2514);
and U9065 (N_9065,N_3565,N_2843);
or U9066 (N_9066,N_4681,N_1356);
and U9067 (N_9067,N_4180,N_24);
nand U9068 (N_9068,N_4289,N_1402);
or U9069 (N_9069,N_1922,N_1714);
nor U9070 (N_9070,N_3237,N_2283);
and U9071 (N_9071,N_1064,N_3688);
nor U9072 (N_9072,N_1365,N_3914);
xnor U9073 (N_9073,N_725,N_2875);
nor U9074 (N_9074,N_3427,N_1746);
nand U9075 (N_9075,N_3010,N_3128);
and U9076 (N_9076,N_3582,N_529);
or U9077 (N_9077,N_2989,N_2949);
nand U9078 (N_9078,N_3705,N_3224);
nand U9079 (N_9079,N_460,N_946);
or U9080 (N_9080,N_974,N_2596);
nor U9081 (N_9081,N_1829,N_3336);
nand U9082 (N_9082,N_3882,N_2145);
and U9083 (N_9083,N_528,N_3317);
or U9084 (N_9084,N_967,N_2731);
nand U9085 (N_9085,N_2002,N_1470);
and U9086 (N_9086,N_1215,N_2931);
nor U9087 (N_9087,N_3106,N_135);
and U9088 (N_9088,N_249,N_1160);
nand U9089 (N_9089,N_549,N_2083);
or U9090 (N_9090,N_2501,N_98);
or U9091 (N_9091,N_2655,N_976);
nor U9092 (N_9092,N_381,N_782);
nor U9093 (N_9093,N_1693,N_510);
nand U9094 (N_9094,N_4971,N_2902);
nand U9095 (N_9095,N_4447,N_301);
and U9096 (N_9096,N_3520,N_851);
nor U9097 (N_9097,N_179,N_1991);
or U9098 (N_9098,N_2372,N_719);
and U9099 (N_9099,N_1078,N_1594);
nor U9100 (N_9100,N_1780,N_4544);
and U9101 (N_9101,N_2951,N_3379);
nand U9102 (N_9102,N_139,N_2245);
nor U9103 (N_9103,N_1088,N_737);
nand U9104 (N_9104,N_856,N_3232);
nand U9105 (N_9105,N_2024,N_2114);
nor U9106 (N_9106,N_3553,N_2471);
nor U9107 (N_9107,N_3839,N_1528);
nor U9108 (N_9108,N_1482,N_4863);
and U9109 (N_9109,N_2460,N_3494);
nor U9110 (N_9110,N_4087,N_3033);
or U9111 (N_9111,N_295,N_4580);
or U9112 (N_9112,N_3616,N_2411);
nor U9113 (N_9113,N_449,N_4115);
and U9114 (N_9114,N_4345,N_4497);
nand U9115 (N_9115,N_4250,N_3337);
or U9116 (N_9116,N_2277,N_3745);
or U9117 (N_9117,N_2730,N_264);
or U9118 (N_9118,N_1325,N_4133);
and U9119 (N_9119,N_3849,N_1698);
nand U9120 (N_9120,N_22,N_247);
nand U9121 (N_9121,N_1504,N_1487);
nor U9122 (N_9122,N_2193,N_2742);
and U9123 (N_9123,N_4528,N_2809);
nand U9124 (N_9124,N_998,N_913);
or U9125 (N_9125,N_1852,N_2900);
nor U9126 (N_9126,N_1232,N_880);
nand U9127 (N_9127,N_4483,N_3006);
or U9128 (N_9128,N_4654,N_3253);
and U9129 (N_9129,N_69,N_4281);
or U9130 (N_9130,N_4197,N_2771);
and U9131 (N_9131,N_34,N_2232);
nor U9132 (N_9132,N_3776,N_4034);
xnor U9133 (N_9133,N_3752,N_160);
nor U9134 (N_9134,N_4126,N_389);
or U9135 (N_9135,N_4895,N_1131);
nor U9136 (N_9136,N_3296,N_4184);
and U9137 (N_9137,N_983,N_2144);
nor U9138 (N_9138,N_1361,N_2923);
nor U9139 (N_9139,N_189,N_1429);
and U9140 (N_9140,N_953,N_236);
nor U9141 (N_9141,N_4329,N_3501);
nand U9142 (N_9142,N_3405,N_512);
or U9143 (N_9143,N_4976,N_2079);
nor U9144 (N_9144,N_1225,N_1679);
and U9145 (N_9145,N_558,N_483);
nor U9146 (N_9146,N_3612,N_223);
nor U9147 (N_9147,N_2441,N_734);
nand U9148 (N_9148,N_1687,N_3743);
nand U9149 (N_9149,N_498,N_2744);
nand U9150 (N_9150,N_320,N_3437);
nand U9151 (N_9151,N_839,N_456);
and U9152 (N_9152,N_4336,N_2301);
nor U9153 (N_9153,N_4958,N_296);
and U9154 (N_9154,N_2065,N_2977);
nand U9155 (N_9155,N_1178,N_3921);
nand U9156 (N_9156,N_2087,N_1078);
or U9157 (N_9157,N_2036,N_4032);
and U9158 (N_9158,N_1907,N_3830);
nand U9159 (N_9159,N_4272,N_4221);
nor U9160 (N_9160,N_2028,N_2322);
or U9161 (N_9161,N_1661,N_3863);
nand U9162 (N_9162,N_4475,N_334);
nand U9163 (N_9163,N_577,N_4885);
and U9164 (N_9164,N_3542,N_120);
nor U9165 (N_9165,N_587,N_4162);
nand U9166 (N_9166,N_1165,N_1101);
nand U9167 (N_9167,N_3142,N_454);
and U9168 (N_9168,N_1222,N_957);
nand U9169 (N_9169,N_934,N_4284);
and U9170 (N_9170,N_2382,N_3423);
nor U9171 (N_9171,N_4973,N_2714);
or U9172 (N_9172,N_4327,N_3481);
or U9173 (N_9173,N_2335,N_2886);
and U9174 (N_9174,N_4147,N_4452);
and U9175 (N_9175,N_2807,N_2801);
nand U9176 (N_9176,N_4714,N_3819);
nor U9177 (N_9177,N_2073,N_1135);
nand U9178 (N_9178,N_549,N_1616);
nor U9179 (N_9179,N_2721,N_3704);
or U9180 (N_9180,N_4071,N_616);
nand U9181 (N_9181,N_2682,N_1128);
nand U9182 (N_9182,N_4209,N_647);
nand U9183 (N_9183,N_1174,N_3175);
and U9184 (N_9184,N_2655,N_1648);
nor U9185 (N_9185,N_3783,N_3532);
nor U9186 (N_9186,N_4829,N_4410);
nand U9187 (N_9187,N_706,N_665);
or U9188 (N_9188,N_4465,N_3611);
nand U9189 (N_9189,N_1751,N_4948);
and U9190 (N_9190,N_4091,N_1020);
nand U9191 (N_9191,N_3726,N_1477);
nand U9192 (N_9192,N_2699,N_4191);
or U9193 (N_9193,N_4108,N_3711);
or U9194 (N_9194,N_1418,N_1821);
or U9195 (N_9195,N_3938,N_2096);
nor U9196 (N_9196,N_2120,N_2367);
and U9197 (N_9197,N_2227,N_692);
and U9198 (N_9198,N_148,N_504);
and U9199 (N_9199,N_4442,N_2594);
and U9200 (N_9200,N_3844,N_4998);
or U9201 (N_9201,N_1480,N_2647);
and U9202 (N_9202,N_1810,N_2462);
and U9203 (N_9203,N_3404,N_3607);
nor U9204 (N_9204,N_4978,N_3994);
nor U9205 (N_9205,N_2500,N_2541);
nor U9206 (N_9206,N_1505,N_3270);
and U9207 (N_9207,N_4017,N_3581);
and U9208 (N_9208,N_4049,N_4376);
and U9209 (N_9209,N_870,N_428);
or U9210 (N_9210,N_2076,N_680);
nand U9211 (N_9211,N_620,N_2302);
and U9212 (N_9212,N_1824,N_1122);
or U9213 (N_9213,N_2496,N_2699);
nand U9214 (N_9214,N_4868,N_3811);
or U9215 (N_9215,N_4767,N_616);
nand U9216 (N_9216,N_1578,N_254);
nand U9217 (N_9217,N_1138,N_4180);
nand U9218 (N_9218,N_974,N_2898);
or U9219 (N_9219,N_4555,N_1655);
nor U9220 (N_9220,N_3185,N_3324);
nor U9221 (N_9221,N_1605,N_3438);
or U9222 (N_9222,N_1361,N_1262);
or U9223 (N_9223,N_2638,N_956);
or U9224 (N_9224,N_4530,N_1975);
or U9225 (N_9225,N_1024,N_2803);
or U9226 (N_9226,N_2216,N_1058);
or U9227 (N_9227,N_1622,N_19);
nor U9228 (N_9228,N_1346,N_963);
or U9229 (N_9229,N_3605,N_364);
and U9230 (N_9230,N_998,N_4762);
and U9231 (N_9231,N_732,N_1431);
nand U9232 (N_9232,N_2218,N_1470);
nor U9233 (N_9233,N_159,N_4991);
and U9234 (N_9234,N_2115,N_3945);
or U9235 (N_9235,N_4361,N_2277);
or U9236 (N_9236,N_1210,N_2338);
nor U9237 (N_9237,N_1487,N_2400);
nand U9238 (N_9238,N_3928,N_4241);
nand U9239 (N_9239,N_1832,N_2228);
nor U9240 (N_9240,N_3756,N_3965);
or U9241 (N_9241,N_2195,N_3464);
nor U9242 (N_9242,N_1946,N_2466);
nand U9243 (N_9243,N_4073,N_4414);
or U9244 (N_9244,N_3690,N_4145);
or U9245 (N_9245,N_1505,N_1365);
nor U9246 (N_9246,N_1752,N_518);
and U9247 (N_9247,N_1889,N_1636);
nor U9248 (N_9248,N_351,N_399);
or U9249 (N_9249,N_914,N_487);
and U9250 (N_9250,N_2055,N_3742);
nand U9251 (N_9251,N_4702,N_4429);
and U9252 (N_9252,N_2474,N_3903);
and U9253 (N_9253,N_3561,N_1624);
nand U9254 (N_9254,N_2743,N_4159);
or U9255 (N_9255,N_4718,N_4347);
nor U9256 (N_9256,N_2209,N_2633);
nand U9257 (N_9257,N_901,N_4715);
nand U9258 (N_9258,N_1507,N_1207);
or U9259 (N_9259,N_1982,N_137);
and U9260 (N_9260,N_637,N_2542);
or U9261 (N_9261,N_1879,N_1118);
nand U9262 (N_9262,N_2826,N_198);
nor U9263 (N_9263,N_3191,N_437);
nand U9264 (N_9264,N_4210,N_2387);
nand U9265 (N_9265,N_2336,N_1119);
or U9266 (N_9266,N_2687,N_2593);
and U9267 (N_9267,N_4762,N_1518);
or U9268 (N_9268,N_3714,N_3238);
or U9269 (N_9269,N_2095,N_3547);
or U9270 (N_9270,N_469,N_1235);
nand U9271 (N_9271,N_1241,N_3729);
xor U9272 (N_9272,N_48,N_4017);
nor U9273 (N_9273,N_2154,N_1766);
or U9274 (N_9274,N_4036,N_3709);
or U9275 (N_9275,N_3577,N_4367);
and U9276 (N_9276,N_4129,N_4928);
or U9277 (N_9277,N_1941,N_2324);
and U9278 (N_9278,N_564,N_3797);
and U9279 (N_9279,N_3211,N_1079);
nand U9280 (N_9280,N_2400,N_3253);
nor U9281 (N_9281,N_4353,N_1034);
nor U9282 (N_9282,N_2843,N_3450);
nor U9283 (N_9283,N_4034,N_3079);
nor U9284 (N_9284,N_893,N_3987);
and U9285 (N_9285,N_4982,N_617);
and U9286 (N_9286,N_2727,N_730);
or U9287 (N_9287,N_2037,N_4414);
nor U9288 (N_9288,N_3644,N_3657);
or U9289 (N_9289,N_1664,N_2778);
nor U9290 (N_9290,N_1421,N_3715);
nand U9291 (N_9291,N_1980,N_1608);
nand U9292 (N_9292,N_2194,N_3789);
and U9293 (N_9293,N_612,N_4847);
or U9294 (N_9294,N_498,N_289);
nand U9295 (N_9295,N_4107,N_4281);
or U9296 (N_9296,N_2749,N_962);
and U9297 (N_9297,N_1700,N_2732);
nor U9298 (N_9298,N_2349,N_3021);
or U9299 (N_9299,N_1056,N_784);
nand U9300 (N_9300,N_2648,N_2383);
or U9301 (N_9301,N_4441,N_2915);
nand U9302 (N_9302,N_2702,N_663);
nor U9303 (N_9303,N_2719,N_3932);
and U9304 (N_9304,N_1436,N_4636);
and U9305 (N_9305,N_164,N_4259);
and U9306 (N_9306,N_2893,N_1446);
nor U9307 (N_9307,N_806,N_4407);
nor U9308 (N_9308,N_3231,N_2574);
nor U9309 (N_9309,N_489,N_1116);
nor U9310 (N_9310,N_3905,N_656);
or U9311 (N_9311,N_2844,N_1384);
nor U9312 (N_9312,N_259,N_3342);
or U9313 (N_9313,N_2671,N_4869);
or U9314 (N_9314,N_2349,N_3793);
and U9315 (N_9315,N_4833,N_876);
or U9316 (N_9316,N_4972,N_2737);
and U9317 (N_9317,N_861,N_4886);
nand U9318 (N_9318,N_2519,N_2235);
or U9319 (N_9319,N_3043,N_671);
or U9320 (N_9320,N_1690,N_3465);
and U9321 (N_9321,N_4283,N_1842);
or U9322 (N_9322,N_320,N_3797);
or U9323 (N_9323,N_1580,N_1961);
and U9324 (N_9324,N_3178,N_1388);
or U9325 (N_9325,N_293,N_3386);
or U9326 (N_9326,N_1446,N_3682);
and U9327 (N_9327,N_1765,N_4977);
nor U9328 (N_9328,N_1414,N_4550);
nand U9329 (N_9329,N_4796,N_1326);
or U9330 (N_9330,N_2687,N_2101);
nor U9331 (N_9331,N_2954,N_811);
and U9332 (N_9332,N_1715,N_3066);
or U9333 (N_9333,N_4891,N_3583);
nor U9334 (N_9334,N_2075,N_3607);
nand U9335 (N_9335,N_3767,N_1685);
and U9336 (N_9336,N_243,N_3473);
or U9337 (N_9337,N_2946,N_2026);
or U9338 (N_9338,N_2941,N_2517);
and U9339 (N_9339,N_1333,N_3844);
nor U9340 (N_9340,N_3202,N_4857);
or U9341 (N_9341,N_4728,N_3324);
nor U9342 (N_9342,N_3962,N_3687);
nand U9343 (N_9343,N_3921,N_4940);
or U9344 (N_9344,N_4811,N_2528);
and U9345 (N_9345,N_2260,N_1870);
nand U9346 (N_9346,N_1381,N_4737);
or U9347 (N_9347,N_4916,N_2821);
and U9348 (N_9348,N_2684,N_2603);
nand U9349 (N_9349,N_4137,N_4823);
nand U9350 (N_9350,N_1805,N_3239);
nand U9351 (N_9351,N_3314,N_3602);
and U9352 (N_9352,N_4290,N_1311);
or U9353 (N_9353,N_1215,N_138);
or U9354 (N_9354,N_3280,N_4080);
nand U9355 (N_9355,N_1537,N_4003);
or U9356 (N_9356,N_3955,N_91);
nand U9357 (N_9357,N_60,N_2922);
and U9358 (N_9358,N_3681,N_1566);
and U9359 (N_9359,N_405,N_845);
nand U9360 (N_9360,N_611,N_2440);
nor U9361 (N_9361,N_665,N_2240);
nand U9362 (N_9362,N_2111,N_2004);
and U9363 (N_9363,N_1380,N_1974);
and U9364 (N_9364,N_3775,N_1022);
nor U9365 (N_9365,N_2364,N_1276);
and U9366 (N_9366,N_3765,N_418);
nand U9367 (N_9367,N_481,N_1137);
or U9368 (N_9368,N_2550,N_2283);
nor U9369 (N_9369,N_1910,N_1457);
nand U9370 (N_9370,N_3277,N_2376);
or U9371 (N_9371,N_1730,N_4888);
or U9372 (N_9372,N_4244,N_4930);
nor U9373 (N_9373,N_4072,N_2768);
and U9374 (N_9374,N_4210,N_434);
nand U9375 (N_9375,N_4648,N_3517);
or U9376 (N_9376,N_1758,N_2976);
or U9377 (N_9377,N_4584,N_4325);
and U9378 (N_9378,N_1742,N_483);
or U9379 (N_9379,N_536,N_4909);
or U9380 (N_9380,N_3235,N_149);
nand U9381 (N_9381,N_1057,N_3813);
or U9382 (N_9382,N_3206,N_2544);
or U9383 (N_9383,N_4103,N_143);
nand U9384 (N_9384,N_842,N_1360);
and U9385 (N_9385,N_2286,N_3811);
nand U9386 (N_9386,N_146,N_147);
nand U9387 (N_9387,N_1577,N_4317);
nand U9388 (N_9388,N_2338,N_2721);
nand U9389 (N_9389,N_365,N_3619);
nand U9390 (N_9390,N_1844,N_660);
nor U9391 (N_9391,N_3967,N_395);
or U9392 (N_9392,N_214,N_17);
and U9393 (N_9393,N_1984,N_2528);
and U9394 (N_9394,N_3608,N_3222);
xor U9395 (N_9395,N_3654,N_1479);
and U9396 (N_9396,N_3309,N_2261);
nand U9397 (N_9397,N_4004,N_3572);
and U9398 (N_9398,N_2781,N_4182);
nand U9399 (N_9399,N_2877,N_2240);
and U9400 (N_9400,N_2865,N_2575);
or U9401 (N_9401,N_2507,N_4054);
or U9402 (N_9402,N_1917,N_3901);
and U9403 (N_9403,N_4259,N_3723);
or U9404 (N_9404,N_1676,N_3995);
or U9405 (N_9405,N_3633,N_240);
nor U9406 (N_9406,N_2372,N_2112);
or U9407 (N_9407,N_573,N_4662);
and U9408 (N_9408,N_3546,N_3122);
or U9409 (N_9409,N_4258,N_991);
nor U9410 (N_9410,N_2086,N_1804);
and U9411 (N_9411,N_4505,N_2620);
nor U9412 (N_9412,N_4668,N_1801);
xor U9413 (N_9413,N_3477,N_2209);
and U9414 (N_9414,N_3063,N_2262);
nand U9415 (N_9415,N_2718,N_779);
xnor U9416 (N_9416,N_2179,N_3345);
nor U9417 (N_9417,N_2347,N_2586);
nand U9418 (N_9418,N_1444,N_1601);
and U9419 (N_9419,N_4158,N_1178);
and U9420 (N_9420,N_3839,N_328);
or U9421 (N_9421,N_997,N_2097);
or U9422 (N_9422,N_1046,N_4084);
or U9423 (N_9423,N_416,N_3477);
nor U9424 (N_9424,N_726,N_1540);
or U9425 (N_9425,N_232,N_2335);
nor U9426 (N_9426,N_4438,N_1829);
nand U9427 (N_9427,N_1017,N_3774);
nor U9428 (N_9428,N_4397,N_1456);
or U9429 (N_9429,N_3841,N_1675);
and U9430 (N_9430,N_2056,N_1055);
and U9431 (N_9431,N_2453,N_1987);
or U9432 (N_9432,N_2759,N_1732);
xnor U9433 (N_9433,N_633,N_3862);
xnor U9434 (N_9434,N_3818,N_2616);
or U9435 (N_9435,N_4562,N_3308);
nand U9436 (N_9436,N_4685,N_1277);
and U9437 (N_9437,N_4522,N_3851);
nor U9438 (N_9438,N_1805,N_412);
nor U9439 (N_9439,N_4793,N_2913);
nor U9440 (N_9440,N_2224,N_2168);
nor U9441 (N_9441,N_4974,N_4653);
or U9442 (N_9442,N_2515,N_2843);
and U9443 (N_9443,N_2294,N_2857);
nor U9444 (N_9444,N_2108,N_2195);
or U9445 (N_9445,N_4396,N_1991);
nor U9446 (N_9446,N_4412,N_4884);
or U9447 (N_9447,N_4446,N_1585);
or U9448 (N_9448,N_1141,N_1552);
nand U9449 (N_9449,N_1475,N_2768);
nor U9450 (N_9450,N_2053,N_4347);
and U9451 (N_9451,N_3396,N_54);
nor U9452 (N_9452,N_1486,N_1799);
nand U9453 (N_9453,N_1476,N_248);
nand U9454 (N_9454,N_3717,N_2934);
nand U9455 (N_9455,N_4251,N_4137);
or U9456 (N_9456,N_3316,N_1185);
and U9457 (N_9457,N_445,N_1574);
and U9458 (N_9458,N_2887,N_712);
nor U9459 (N_9459,N_4834,N_4406);
nor U9460 (N_9460,N_4673,N_3769);
or U9461 (N_9461,N_3616,N_2332);
nand U9462 (N_9462,N_1497,N_329);
xnor U9463 (N_9463,N_1400,N_3454);
nor U9464 (N_9464,N_4994,N_3652);
nor U9465 (N_9465,N_4128,N_871);
and U9466 (N_9466,N_2370,N_3851);
nand U9467 (N_9467,N_2063,N_599);
nand U9468 (N_9468,N_1256,N_2956);
and U9469 (N_9469,N_3879,N_877);
or U9470 (N_9470,N_282,N_877);
and U9471 (N_9471,N_2501,N_298);
and U9472 (N_9472,N_908,N_1218);
and U9473 (N_9473,N_3321,N_4490);
and U9474 (N_9474,N_3434,N_1492);
nand U9475 (N_9475,N_2619,N_981);
or U9476 (N_9476,N_1082,N_4961);
and U9477 (N_9477,N_1868,N_4371);
nand U9478 (N_9478,N_2857,N_4705);
nand U9479 (N_9479,N_216,N_702);
or U9480 (N_9480,N_3522,N_1092);
nor U9481 (N_9481,N_2394,N_4965);
or U9482 (N_9482,N_3459,N_505);
nor U9483 (N_9483,N_3597,N_2601);
nor U9484 (N_9484,N_4698,N_3411);
nand U9485 (N_9485,N_113,N_2664);
and U9486 (N_9486,N_4714,N_202);
or U9487 (N_9487,N_1376,N_4385);
nand U9488 (N_9488,N_4500,N_3357);
or U9489 (N_9489,N_4812,N_2100);
nand U9490 (N_9490,N_2181,N_637);
or U9491 (N_9491,N_2981,N_626);
or U9492 (N_9492,N_869,N_807);
nor U9493 (N_9493,N_4825,N_2534);
and U9494 (N_9494,N_38,N_126);
and U9495 (N_9495,N_4806,N_3215);
or U9496 (N_9496,N_224,N_1236);
nand U9497 (N_9497,N_2336,N_3486);
nand U9498 (N_9498,N_776,N_2758);
and U9499 (N_9499,N_2398,N_755);
or U9500 (N_9500,N_4661,N_1250);
nor U9501 (N_9501,N_3470,N_1831);
nand U9502 (N_9502,N_4651,N_3705);
nand U9503 (N_9503,N_3769,N_4742);
nand U9504 (N_9504,N_127,N_759);
nor U9505 (N_9505,N_1584,N_1631);
or U9506 (N_9506,N_2047,N_3928);
nor U9507 (N_9507,N_4029,N_1103);
nand U9508 (N_9508,N_4926,N_3338);
nand U9509 (N_9509,N_720,N_1582);
or U9510 (N_9510,N_3361,N_2298);
nand U9511 (N_9511,N_430,N_121);
nor U9512 (N_9512,N_2816,N_3698);
nor U9513 (N_9513,N_3574,N_2574);
nand U9514 (N_9514,N_2460,N_2728);
nor U9515 (N_9515,N_77,N_3509);
nor U9516 (N_9516,N_853,N_4906);
and U9517 (N_9517,N_1795,N_1967);
nand U9518 (N_9518,N_3393,N_4498);
and U9519 (N_9519,N_3288,N_2450);
nand U9520 (N_9520,N_3595,N_3351);
and U9521 (N_9521,N_2812,N_1432);
nor U9522 (N_9522,N_4908,N_2724);
nor U9523 (N_9523,N_4302,N_4937);
nand U9524 (N_9524,N_2428,N_3732);
or U9525 (N_9525,N_647,N_317);
or U9526 (N_9526,N_4218,N_3382);
nor U9527 (N_9527,N_3730,N_4220);
or U9528 (N_9528,N_3801,N_1966);
nand U9529 (N_9529,N_2983,N_4460);
or U9530 (N_9530,N_4853,N_1980);
nor U9531 (N_9531,N_1510,N_3940);
nand U9532 (N_9532,N_3972,N_628);
nor U9533 (N_9533,N_546,N_1531);
nand U9534 (N_9534,N_1970,N_2723);
and U9535 (N_9535,N_1695,N_1026);
nand U9536 (N_9536,N_1421,N_4335);
and U9537 (N_9537,N_4593,N_4774);
nor U9538 (N_9538,N_186,N_3028);
nor U9539 (N_9539,N_4331,N_3889);
or U9540 (N_9540,N_4968,N_295);
or U9541 (N_9541,N_3971,N_4331);
nor U9542 (N_9542,N_779,N_3596);
or U9543 (N_9543,N_4416,N_3260);
nor U9544 (N_9544,N_2407,N_3738);
or U9545 (N_9545,N_1837,N_1021);
or U9546 (N_9546,N_4500,N_4104);
and U9547 (N_9547,N_4960,N_2596);
or U9548 (N_9548,N_4293,N_1749);
and U9549 (N_9549,N_24,N_1054);
and U9550 (N_9550,N_120,N_4543);
nor U9551 (N_9551,N_3294,N_504);
or U9552 (N_9552,N_3831,N_3464);
or U9553 (N_9553,N_2455,N_3371);
nor U9554 (N_9554,N_4761,N_1147);
nor U9555 (N_9555,N_1397,N_2023);
nor U9556 (N_9556,N_889,N_3258);
nor U9557 (N_9557,N_371,N_3043);
nor U9558 (N_9558,N_2341,N_1852);
nand U9559 (N_9559,N_3985,N_56);
or U9560 (N_9560,N_3238,N_298);
and U9561 (N_9561,N_4247,N_1880);
nand U9562 (N_9562,N_1363,N_555);
nor U9563 (N_9563,N_3167,N_294);
or U9564 (N_9564,N_4201,N_1711);
nand U9565 (N_9565,N_484,N_4926);
or U9566 (N_9566,N_846,N_3771);
and U9567 (N_9567,N_2738,N_1233);
nor U9568 (N_9568,N_371,N_4773);
or U9569 (N_9569,N_2581,N_987);
nand U9570 (N_9570,N_4967,N_4433);
nor U9571 (N_9571,N_3235,N_4352);
and U9572 (N_9572,N_1383,N_4864);
nor U9573 (N_9573,N_822,N_707);
and U9574 (N_9574,N_1813,N_4679);
nor U9575 (N_9575,N_1720,N_2488);
and U9576 (N_9576,N_4728,N_3939);
nand U9577 (N_9577,N_3283,N_2309);
nand U9578 (N_9578,N_1522,N_814);
and U9579 (N_9579,N_138,N_3185);
nor U9580 (N_9580,N_1488,N_1457);
and U9581 (N_9581,N_649,N_4043);
nand U9582 (N_9582,N_1391,N_2107);
and U9583 (N_9583,N_1354,N_4800);
xnor U9584 (N_9584,N_2291,N_3634);
nor U9585 (N_9585,N_2426,N_183);
and U9586 (N_9586,N_3619,N_93);
and U9587 (N_9587,N_2644,N_492);
nor U9588 (N_9588,N_1530,N_788);
or U9589 (N_9589,N_2391,N_1461);
nand U9590 (N_9590,N_1428,N_2188);
or U9591 (N_9591,N_3633,N_2437);
or U9592 (N_9592,N_2066,N_1564);
nand U9593 (N_9593,N_4340,N_2182);
or U9594 (N_9594,N_931,N_318);
nand U9595 (N_9595,N_2362,N_2364);
nor U9596 (N_9596,N_4888,N_2773);
and U9597 (N_9597,N_403,N_812);
or U9598 (N_9598,N_447,N_214);
nor U9599 (N_9599,N_1020,N_1646);
or U9600 (N_9600,N_848,N_2535);
and U9601 (N_9601,N_137,N_4355);
and U9602 (N_9602,N_607,N_2575);
or U9603 (N_9603,N_3022,N_688);
nor U9604 (N_9604,N_3600,N_150);
and U9605 (N_9605,N_2361,N_1359);
and U9606 (N_9606,N_1247,N_2208);
nor U9607 (N_9607,N_1151,N_3170);
and U9608 (N_9608,N_3053,N_1425);
nor U9609 (N_9609,N_78,N_3650);
or U9610 (N_9610,N_3738,N_562);
or U9611 (N_9611,N_910,N_3731);
and U9612 (N_9612,N_3559,N_4388);
or U9613 (N_9613,N_1503,N_3918);
nor U9614 (N_9614,N_3318,N_4216);
or U9615 (N_9615,N_3483,N_4777);
and U9616 (N_9616,N_2080,N_758);
nor U9617 (N_9617,N_2441,N_4025);
or U9618 (N_9618,N_815,N_4786);
nand U9619 (N_9619,N_4925,N_300);
and U9620 (N_9620,N_3396,N_182);
nand U9621 (N_9621,N_343,N_2136);
nor U9622 (N_9622,N_4084,N_2719);
nand U9623 (N_9623,N_3130,N_2347);
and U9624 (N_9624,N_3641,N_2603);
nand U9625 (N_9625,N_3769,N_3690);
nand U9626 (N_9626,N_4129,N_755);
nand U9627 (N_9627,N_4334,N_1886);
nor U9628 (N_9628,N_4394,N_3272);
nor U9629 (N_9629,N_2705,N_1971);
xor U9630 (N_9630,N_2816,N_2613);
or U9631 (N_9631,N_1321,N_1206);
nand U9632 (N_9632,N_3260,N_4791);
or U9633 (N_9633,N_1244,N_4291);
nor U9634 (N_9634,N_785,N_4591);
and U9635 (N_9635,N_1165,N_1448);
and U9636 (N_9636,N_3866,N_1807);
nor U9637 (N_9637,N_4700,N_61);
or U9638 (N_9638,N_334,N_2332);
nor U9639 (N_9639,N_3060,N_4737);
or U9640 (N_9640,N_2238,N_643);
nor U9641 (N_9641,N_1146,N_3275);
or U9642 (N_9642,N_3459,N_654);
nor U9643 (N_9643,N_3596,N_923);
nand U9644 (N_9644,N_3482,N_166);
nor U9645 (N_9645,N_3072,N_2288);
or U9646 (N_9646,N_416,N_4644);
nor U9647 (N_9647,N_4505,N_1308);
and U9648 (N_9648,N_1693,N_748);
xnor U9649 (N_9649,N_363,N_3681);
and U9650 (N_9650,N_3212,N_368);
nor U9651 (N_9651,N_980,N_3215);
and U9652 (N_9652,N_398,N_3256);
nand U9653 (N_9653,N_3507,N_4537);
nor U9654 (N_9654,N_3336,N_2324);
and U9655 (N_9655,N_4557,N_648);
nor U9656 (N_9656,N_732,N_727);
nor U9657 (N_9657,N_4421,N_4419);
and U9658 (N_9658,N_1258,N_768);
or U9659 (N_9659,N_4468,N_1466);
xnor U9660 (N_9660,N_4741,N_1241);
or U9661 (N_9661,N_98,N_192);
or U9662 (N_9662,N_3679,N_3748);
nor U9663 (N_9663,N_1527,N_366);
and U9664 (N_9664,N_4318,N_4059);
nand U9665 (N_9665,N_4825,N_1950);
and U9666 (N_9666,N_3213,N_4654);
nor U9667 (N_9667,N_1229,N_3613);
nand U9668 (N_9668,N_3848,N_132);
nand U9669 (N_9669,N_4704,N_809);
nand U9670 (N_9670,N_131,N_2627);
nand U9671 (N_9671,N_4389,N_2231);
nor U9672 (N_9672,N_2909,N_1591);
and U9673 (N_9673,N_2589,N_277);
or U9674 (N_9674,N_4636,N_4427);
or U9675 (N_9675,N_3643,N_2199);
nor U9676 (N_9676,N_2582,N_1442);
nand U9677 (N_9677,N_1542,N_4980);
and U9678 (N_9678,N_507,N_100);
or U9679 (N_9679,N_384,N_1520);
nand U9680 (N_9680,N_882,N_186);
nor U9681 (N_9681,N_222,N_2633);
or U9682 (N_9682,N_136,N_2254);
nor U9683 (N_9683,N_308,N_226);
nand U9684 (N_9684,N_3873,N_1597);
or U9685 (N_9685,N_2675,N_389);
and U9686 (N_9686,N_3596,N_2270);
or U9687 (N_9687,N_4078,N_4281);
nand U9688 (N_9688,N_2341,N_3453);
nand U9689 (N_9689,N_2065,N_41);
nand U9690 (N_9690,N_1246,N_2324);
nand U9691 (N_9691,N_2395,N_558);
nand U9692 (N_9692,N_4312,N_4003);
and U9693 (N_9693,N_1374,N_1940);
nand U9694 (N_9694,N_269,N_121);
or U9695 (N_9695,N_4954,N_591);
xnor U9696 (N_9696,N_2848,N_3904);
nand U9697 (N_9697,N_1786,N_3459);
and U9698 (N_9698,N_4177,N_3728);
nor U9699 (N_9699,N_2628,N_4986);
and U9700 (N_9700,N_1006,N_889);
nor U9701 (N_9701,N_928,N_2365);
nand U9702 (N_9702,N_991,N_2187);
and U9703 (N_9703,N_1806,N_1034);
nand U9704 (N_9704,N_4461,N_2342);
and U9705 (N_9705,N_1809,N_478);
nor U9706 (N_9706,N_808,N_373);
and U9707 (N_9707,N_1160,N_1486);
nand U9708 (N_9708,N_4442,N_825);
or U9709 (N_9709,N_3551,N_338);
nor U9710 (N_9710,N_4540,N_1353);
nor U9711 (N_9711,N_278,N_100);
xnor U9712 (N_9712,N_2144,N_310);
nand U9713 (N_9713,N_1320,N_3685);
nor U9714 (N_9714,N_3735,N_2309);
and U9715 (N_9715,N_367,N_3351);
nor U9716 (N_9716,N_4181,N_108);
nand U9717 (N_9717,N_940,N_4453);
nor U9718 (N_9718,N_2180,N_3210);
nor U9719 (N_9719,N_1590,N_3253);
nand U9720 (N_9720,N_1652,N_612);
xor U9721 (N_9721,N_2345,N_4802);
and U9722 (N_9722,N_3594,N_4918);
and U9723 (N_9723,N_623,N_2741);
and U9724 (N_9724,N_4310,N_4382);
or U9725 (N_9725,N_1295,N_3234);
and U9726 (N_9726,N_3197,N_1144);
and U9727 (N_9727,N_1391,N_3410);
and U9728 (N_9728,N_4165,N_1900);
nor U9729 (N_9729,N_2902,N_202);
and U9730 (N_9730,N_1092,N_4341);
or U9731 (N_9731,N_2085,N_1101);
or U9732 (N_9732,N_2982,N_926);
nor U9733 (N_9733,N_3299,N_236);
nand U9734 (N_9734,N_1309,N_1264);
nand U9735 (N_9735,N_1405,N_3642);
nor U9736 (N_9736,N_3745,N_2200);
nand U9737 (N_9737,N_2493,N_2350);
nand U9738 (N_9738,N_4488,N_3832);
and U9739 (N_9739,N_4559,N_2314);
or U9740 (N_9740,N_2970,N_1941);
or U9741 (N_9741,N_623,N_4698);
and U9742 (N_9742,N_417,N_3034);
or U9743 (N_9743,N_4716,N_1091);
nor U9744 (N_9744,N_4302,N_1898);
nor U9745 (N_9745,N_2788,N_163);
nor U9746 (N_9746,N_1717,N_3975);
nor U9747 (N_9747,N_4902,N_1625);
or U9748 (N_9748,N_2074,N_4872);
nand U9749 (N_9749,N_1691,N_4243);
or U9750 (N_9750,N_1947,N_368);
and U9751 (N_9751,N_2895,N_339);
nor U9752 (N_9752,N_2693,N_3658);
nand U9753 (N_9753,N_831,N_4735);
or U9754 (N_9754,N_660,N_2296);
nor U9755 (N_9755,N_4787,N_2241);
or U9756 (N_9756,N_1126,N_3520);
nand U9757 (N_9757,N_892,N_4125);
nor U9758 (N_9758,N_4631,N_293);
and U9759 (N_9759,N_3569,N_1847);
or U9760 (N_9760,N_2747,N_3334);
xor U9761 (N_9761,N_1630,N_1421);
or U9762 (N_9762,N_899,N_1678);
or U9763 (N_9763,N_4701,N_4306);
or U9764 (N_9764,N_2694,N_1133);
and U9765 (N_9765,N_2179,N_2584);
nor U9766 (N_9766,N_1280,N_1220);
nand U9767 (N_9767,N_1382,N_2092);
nor U9768 (N_9768,N_2550,N_1249);
nor U9769 (N_9769,N_353,N_2213);
or U9770 (N_9770,N_2949,N_578);
or U9771 (N_9771,N_227,N_11);
and U9772 (N_9772,N_1545,N_4063);
nor U9773 (N_9773,N_1640,N_2322);
nand U9774 (N_9774,N_1069,N_2087);
nand U9775 (N_9775,N_431,N_211);
and U9776 (N_9776,N_3816,N_2724);
nand U9777 (N_9777,N_566,N_4644);
nor U9778 (N_9778,N_170,N_51);
xor U9779 (N_9779,N_1070,N_3813);
nor U9780 (N_9780,N_3929,N_4678);
and U9781 (N_9781,N_449,N_3420);
nor U9782 (N_9782,N_4947,N_840);
nor U9783 (N_9783,N_3336,N_263);
and U9784 (N_9784,N_963,N_1427);
or U9785 (N_9785,N_4316,N_1215);
xor U9786 (N_9786,N_3976,N_4164);
nor U9787 (N_9787,N_44,N_1329);
nand U9788 (N_9788,N_1352,N_1371);
or U9789 (N_9789,N_878,N_4118);
nand U9790 (N_9790,N_2308,N_1476);
or U9791 (N_9791,N_3676,N_2087);
nor U9792 (N_9792,N_3641,N_1646);
nand U9793 (N_9793,N_4576,N_7);
or U9794 (N_9794,N_4917,N_2586);
or U9795 (N_9795,N_4511,N_4877);
or U9796 (N_9796,N_2577,N_4614);
nand U9797 (N_9797,N_5,N_3164);
or U9798 (N_9798,N_4274,N_573);
and U9799 (N_9799,N_2147,N_1665);
or U9800 (N_9800,N_4894,N_2938);
and U9801 (N_9801,N_3423,N_3365);
nand U9802 (N_9802,N_2867,N_1029);
nor U9803 (N_9803,N_1045,N_4221);
and U9804 (N_9804,N_2996,N_1047);
nand U9805 (N_9805,N_1750,N_2759);
and U9806 (N_9806,N_3237,N_3765);
nand U9807 (N_9807,N_4808,N_3250);
nor U9808 (N_9808,N_4645,N_3045);
and U9809 (N_9809,N_2159,N_982);
and U9810 (N_9810,N_1119,N_4370);
and U9811 (N_9811,N_3710,N_358);
or U9812 (N_9812,N_3379,N_2315);
or U9813 (N_9813,N_3932,N_3139);
nand U9814 (N_9814,N_2759,N_1443);
and U9815 (N_9815,N_2434,N_3978);
nand U9816 (N_9816,N_4428,N_258);
or U9817 (N_9817,N_3916,N_2447);
nor U9818 (N_9818,N_681,N_2790);
or U9819 (N_9819,N_291,N_491);
or U9820 (N_9820,N_115,N_2840);
nand U9821 (N_9821,N_170,N_1810);
nand U9822 (N_9822,N_4848,N_4341);
or U9823 (N_9823,N_1863,N_182);
nand U9824 (N_9824,N_4181,N_4172);
nand U9825 (N_9825,N_2145,N_4186);
nand U9826 (N_9826,N_1429,N_816);
nor U9827 (N_9827,N_1385,N_1079);
or U9828 (N_9828,N_4339,N_1671);
and U9829 (N_9829,N_3076,N_1716);
xor U9830 (N_9830,N_2710,N_2545);
nor U9831 (N_9831,N_2970,N_4418);
and U9832 (N_9832,N_1537,N_122);
nor U9833 (N_9833,N_1128,N_2408);
xor U9834 (N_9834,N_4860,N_1445);
or U9835 (N_9835,N_3366,N_461);
and U9836 (N_9836,N_3880,N_4691);
nor U9837 (N_9837,N_3806,N_4203);
or U9838 (N_9838,N_3310,N_1790);
or U9839 (N_9839,N_4784,N_2232);
nor U9840 (N_9840,N_2754,N_2609);
nand U9841 (N_9841,N_1176,N_3721);
nor U9842 (N_9842,N_431,N_1952);
or U9843 (N_9843,N_566,N_4203);
or U9844 (N_9844,N_3971,N_458);
or U9845 (N_9845,N_1381,N_2611);
nor U9846 (N_9846,N_3450,N_2738);
or U9847 (N_9847,N_2071,N_24);
nand U9848 (N_9848,N_2850,N_1360);
nor U9849 (N_9849,N_3217,N_2911);
or U9850 (N_9850,N_412,N_4208);
nand U9851 (N_9851,N_548,N_295);
nor U9852 (N_9852,N_4157,N_3099);
and U9853 (N_9853,N_4455,N_3541);
nor U9854 (N_9854,N_2516,N_47);
and U9855 (N_9855,N_489,N_4240);
and U9856 (N_9856,N_666,N_515);
nor U9857 (N_9857,N_2231,N_4011);
and U9858 (N_9858,N_4506,N_1129);
or U9859 (N_9859,N_1579,N_4904);
and U9860 (N_9860,N_4843,N_4752);
nor U9861 (N_9861,N_4216,N_3445);
nor U9862 (N_9862,N_4396,N_2649);
or U9863 (N_9863,N_1701,N_3493);
and U9864 (N_9864,N_4375,N_2779);
nand U9865 (N_9865,N_2949,N_4068);
nor U9866 (N_9866,N_1465,N_4197);
and U9867 (N_9867,N_3069,N_4310);
nor U9868 (N_9868,N_1619,N_2422);
and U9869 (N_9869,N_1890,N_4863);
and U9870 (N_9870,N_1303,N_2809);
nand U9871 (N_9871,N_1991,N_2650);
nand U9872 (N_9872,N_4556,N_1512);
and U9873 (N_9873,N_3244,N_1302);
and U9874 (N_9874,N_179,N_2991);
or U9875 (N_9875,N_801,N_1520);
or U9876 (N_9876,N_4950,N_2948);
nand U9877 (N_9877,N_17,N_1199);
nor U9878 (N_9878,N_3706,N_981);
or U9879 (N_9879,N_776,N_3792);
nand U9880 (N_9880,N_2799,N_2406);
nand U9881 (N_9881,N_4216,N_1490);
nor U9882 (N_9882,N_4621,N_135);
and U9883 (N_9883,N_2961,N_804);
nor U9884 (N_9884,N_3567,N_2784);
nor U9885 (N_9885,N_2172,N_3930);
nor U9886 (N_9886,N_1771,N_3985);
nor U9887 (N_9887,N_4534,N_4890);
nor U9888 (N_9888,N_1065,N_146);
nor U9889 (N_9889,N_3908,N_4990);
or U9890 (N_9890,N_3616,N_508);
nand U9891 (N_9891,N_504,N_926);
nor U9892 (N_9892,N_2829,N_2780);
and U9893 (N_9893,N_4436,N_1389);
nor U9894 (N_9894,N_2541,N_1629);
nor U9895 (N_9895,N_1482,N_2231);
and U9896 (N_9896,N_381,N_3281);
and U9897 (N_9897,N_739,N_1842);
nor U9898 (N_9898,N_704,N_4130);
and U9899 (N_9899,N_718,N_893);
or U9900 (N_9900,N_342,N_244);
or U9901 (N_9901,N_2379,N_3546);
and U9902 (N_9902,N_2527,N_4985);
nor U9903 (N_9903,N_2281,N_4215);
nand U9904 (N_9904,N_53,N_3544);
and U9905 (N_9905,N_3390,N_381);
or U9906 (N_9906,N_3424,N_2861);
or U9907 (N_9907,N_1008,N_4637);
nor U9908 (N_9908,N_742,N_1064);
or U9909 (N_9909,N_363,N_3556);
and U9910 (N_9910,N_2089,N_1642);
and U9911 (N_9911,N_3294,N_4637);
or U9912 (N_9912,N_2832,N_1054);
and U9913 (N_9913,N_4795,N_1110);
nand U9914 (N_9914,N_4624,N_4947);
and U9915 (N_9915,N_211,N_2216);
nor U9916 (N_9916,N_4995,N_3394);
nor U9917 (N_9917,N_390,N_3262);
and U9918 (N_9918,N_891,N_2531);
or U9919 (N_9919,N_3053,N_423);
nand U9920 (N_9920,N_2489,N_4969);
nand U9921 (N_9921,N_4708,N_3986);
and U9922 (N_9922,N_2411,N_2435);
or U9923 (N_9923,N_1531,N_4875);
and U9924 (N_9924,N_4033,N_2967);
nor U9925 (N_9925,N_3788,N_2879);
nand U9926 (N_9926,N_500,N_4471);
nor U9927 (N_9927,N_2190,N_4160);
and U9928 (N_9928,N_2741,N_971);
or U9929 (N_9929,N_4817,N_3174);
nor U9930 (N_9930,N_3846,N_4148);
nand U9931 (N_9931,N_2798,N_2064);
nor U9932 (N_9932,N_2405,N_3847);
xor U9933 (N_9933,N_811,N_1385);
or U9934 (N_9934,N_851,N_2292);
or U9935 (N_9935,N_599,N_965);
nor U9936 (N_9936,N_2764,N_702);
nand U9937 (N_9937,N_4699,N_4353);
nor U9938 (N_9938,N_3849,N_4863);
nor U9939 (N_9939,N_3548,N_1702);
or U9940 (N_9940,N_1953,N_648);
nand U9941 (N_9941,N_2175,N_1435);
and U9942 (N_9942,N_426,N_4317);
nand U9943 (N_9943,N_4157,N_1571);
nand U9944 (N_9944,N_917,N_591);
nand U9945 (N_9945,N_2524,N_606);
and U9946 (N_9946,N_770,N_4138);
nand U9947 (N_9947,N_1074,N_1260);
nand U9948 (N_9948,N_3569,N_3883);
nand U9949 (N_9949,N_0,N_4942);
and U9950 (N_9950,N_911,N_3559);
nor U9951 (N_9951,N_3159,N_3061);
nand U9952 (N_9952,N_714,N_940);
nand U9953 (N_9953,N_3981,N_4623);
nand U9954 (N_9954,N_2916,N_2321);
and U9955 (N_9955,N_1050,N_1735);
and U9956 (N_9956,N_3315,N_2976);
or U9957 (N_9957,N_4032,N_2709);
or U9958 (N_9958,N_2308,N_4446);
or U9959 (N_9959,N_3049,N_233);
or U9960 (N_9960,N_4486,N_2151);
or U9961 (N_9961,N_2444,N_34);
and U9962 (N_9962,N_4770,N_2808);
xor U9963 (N_9963,N_1485,N_754);
nor U9964 (N_9964,N_4116,N_1836);
and U9965 (N_9965,N_1270,N_1251);
nor U9966 (N_9966,N_4226,N_3114);
or U9967 (N_9967,N_132,N_3368);
or U9968 (N_9968,N_496,N_257);
nand U9969 (N_9969,N_3313,N_3171);
nand U9970 (N_9970,N_2646,N_1142);
and U9971 (N_9971,N_1939,N_2835);
or U9972 (N_9972,N_4086,N_902);
and U9973 (N_9973,N_1848,N_3080);
nor U9974 (N_9974,N_1580,N_4008);
or U9975 (N_9975,N_46,N_2727);
nor U9976 (N_9976,N_1399,N_3288);
nand U9977 (N_9977,N_4371,N_2144);
nand U9978 (N_9978,N_4552,N_900);
or U9979 (N_9979,N_2439,N_651);
nand U9980 (N_9980,N_4032,N_1403);
or U9981 (N_9981,N_198,N_4623);
and U9982 (N_9982,N_80,N_506);
nor U9983 (N_9983,N_1307,N_1787);
or U9984 (N_9984,N_204,N_2185);
and U9985 (N_9985,N_1110,N_2313);
nor U9986 (N_9986,N_3306,N_3417);
or U9987 (N_9987,N_1752,N_77);
and U9988 (N_9988,N_16,N_2547);
nand U9989 (N_9989,N_2151,N_3279);
nor U9990 (N_9990,N_4858,N_2790);
or U9991 (N_9991,N_1726,N_2419);
and U9992 (N_9992,N_2208,N_1242);
nand U9993 (N_9993,N_2578,N_3073);
nor U9994 (N_9994,N_1637,N_2006);
nor U9995 (N_9995,N_976,N_2379);
nor U9996 (N_9996,N_273,N_3505);
nor U9997 (N_9997,N_1501,N_4132);
nor U9998 (N_9998,N_3938,N_1260);
or U9999 (N_9999,N_4488,N_4110);
and UO_0 (O_0,N_7756,N_5635);
nor UO_1 (O_1,N_8023,N_8721);
nor UO_2 (O_2,N_9352,N_5641);
or UO_3 (O_3,N_6037,N_9084);
or UO_4 (O_4,N_6354,N_7893);
or UO_5 (O_5,N_7225,N_7002);
nand UO_6 (O_6,N_5404,N_7717);
or UO_7 (O_7,N_7882,N_7352);
or UO_8 (O_8,N_7759,N_6079);
nand UO_9 (O_9,N_7190,N_9452);
nand UO_10 (O_10,N_5540,N_8936);
and UO_11 (O_11,N_7184,N_6592);
nor UO_12 (O_12,N_5391,N_9299);
and UO_13 (O_13,N_9247,N_9919);
nand UO_14 (O_14,N_8793,N_8674);
nor UO_15 (O_15,N_5973,N_6909);
or UO_16 (O_16,N_7192,N_5501);
or UO_17 (O_17,N_6426,N_7417);
nor UO_18 (O_18,N_7622,N_5523);
nand UO_19 (O_19,N_9342,N_7782);
and UO_20 (O_20,N_7284,N_5985);
nor UO_21 (O_21,N_9599,N_7525);
and UO_22 (O_22,N_6882,N_6436);
and UO_23 (O_23,N_9478,N_5430);
nor UO_24 (O_24,N_5765,N_7143);
nand UO_25 (O_25,N_5812,N_7557);
nor UO_26 (O_26,N_9748,N_7397);
nand UO_27 (O_27,N_8537,N_5190);
and UO_28 (O_28,N_5151,N_8574);
nor UO_29 (O_29,N_6424,N_5322);
and UO_30 (O_30,N_8947,N_9311);
nand UO_31 (O_31,N_7711,N_6522);
nor UO_32 (O_32,N_5869,N_9784);
or UO_33 (O_33,N_8461,N_8206);
xnor UO_34 (O_34,N_6264,N_7987);
and UO_35 (O_35,N_6686,N_9976);
nand UO_36 (O_36,N_9064,N_6525);
or UO_37 (O_37,N_8358,N_6348);
nand UO_38 (O_38,N_6473,N_7850);
or UO_39 (O_39,N_5307,N_8983);
nand UO_40 (O_40,N_8715,N_9281);
or UO_41 (O_41,N_8694,N_5166);
and UO_42 (O_42,N_5539,N_6123);
nor UO_43 (O_43,N_9155,N_6710);
or UO_44 (O_44,N_7999,N_8436);
nand UO_45 (O_45,N_7678,N_6230);
or UO_46 (O_46,N_7962,N_9592);
nor UO_47 (O_47,N_6487,N_5184);
or UO_48 (O_48,N_9612,N_7776);
or UO_49 (O_49,N_6517,N_8089);
nand UO_50 (O_50,N_5308,N_6973);
and UO_51 (O_51,N_7285,N_5572);
nor UO_52 (O_52,N_6219,N_6607);
or UO_53 (O_53,N_7670,N_9934);
or UO_54 (O_54,N_7356,N_9657);
or UO_55 (O_55,N_8034,N_9940);
and UO_56 (O_56,N_6548,N_5874);
nor UO_57 (O_57,N_7728,N_7599);
or UO_58 (O_58,N_5024,N_6901);
nor UO_59 (O_59,N_8748,N_6139);
or UO_60 (O_60,N_6254,N_8512);
and UO_61 (O_61,N_9979,N_7402);
nand UO_62 (O_62,N_9947,N_5662);
and UO_63 (O_63,N_8705,N_7532);
xnor UO_64 (O_64,N_8796,N_8202);
nor UO_65 (O_65,N_7445,N_9914);
and UO_66 (O_66,N_5928,N_5750);
nand UO_67 (O_67,N_6477,N_5037);
nor UO_68 (O_68,N_5624,N_9754);
nand UO_69 (O_69,N_6338,N_5000);
nor UO_70 (O_70,N_8524,N_9893);
nand UO_71 (O_71,N_6930,N_7818);
or UO_72 (O_72,N_7311,N_5556);
nor UO_73 (O_73,N_6696,N_8801);
or UO_74 (O_74,N_7546,N_9369);
nor UO_75 (O_75,N_9750,N_8119);
nand UO_76 (O_76,N_9703,N_7039);
nand UO_77 (O_77,N_5981,N_5658);
and UO_78 (O_78,N_6545,N_5642);
and UO_79 (O_79,N_9404,N_8451);
and UO_80 (O_80,N_6620,N_7709);
nor UO_81 (O_81,N_9395,N_8097);
nand UO_82 (O_82,N_6115,N_8808);
and UO_83 (O_83,N_5086,N_6834);
xnor UO_84 (O_84,N_6726,N_8906);
or UO_85 (O_85,N_6020,N_9805);
nand UO_86 (O_86,N_8734,N_6077);
nor UO_87 (O_87,N_8256,N_6113);
and UO_88 (O_88,N_8806,N_7376);
nor UO_89 (O_89,N_6950,N_6032);
nand UO_90 (O_90,N_9324,N_9020);
or UO_91 (O_91,N_7792,N_5186);
nand UO_92 (O_92,N_6107,N_7297);
or UO_93 (O_93,N_7841,N_6804);
and UO_94 (O_94,N_5916,N_5757);
nor UO_95 (O_95,N_8786,N_8121);
or UO_96 (O_96,N_9670,N_8586);
or UO_97 (O_97,N_9686,N_6287);
or UO_98 (O_98,N_7357,N_7022);
and UO_99 (O_99,N_5801,N_8720);
nand UO_100 (O_100,N_5761,N_9560);
or UO_101 (O_101,N_5449,N_5313);
and UO_102 (O_102,N_9231,N_8476);
and UO_103 (O_103,N_8094,N_8951);
nor UO_104 (O_104,N_6389,N_6922);
nor UO_105 (O_105,N_5866,N_5298);
nor UO_106 (O_106,N_8261,N_7720);
and UO_107 (O_107,N_9021,N_6168);
nor UO_108 (O_108,N_5249,N_5517);
or UO_109 (O_109,N_9114,N_6279);
nand UO_110 (O_110,N_6866,N_8170);
nor UO_111 (O_111,N_5768,N_7423);
nor UO_112 (O_112,N_7049,N_9801);
and UO_113 (O_113,N_8509,N_5390);
xnor UO_114 (O_114,N_5243,N_9116);
or UO_115 (O_115,N_9946,N_8057);
nand UO_116 (O_116,N_7632,N_9425);
nor UO_117 (O_117,N_6434,N_5117);
nand UO_118 (O_118,N_6797,N_8555);
or UO_119 (O_119,N_8063,N_8559);
and UO_120 (O_120,N_9485,N_8904);
or UO_121 (O_121,N_8542,N_8083);
nor UO_122 (O_122,N_8124,N_9582);
or UO_123 (O_123,N_7136,N_8523);
nor UO_124 (O_124,N_8493,N_5235);
nand UO_125 (O_125,N_7770,N_7306);
nor UO_126 (O_126,N_6421,N_6148);
nor UO_127 (O_127,N_8249,N_8272);
nand UO_128 (O_128,N_8031,N_6367);
nand UO_129 (O_129,N_7856,N_6376);
xnor UO_130 (O_130,N_5018,N_5553);
or UO_131 (O_131,N_7147,N_7953);
and UO_132 (O_132,N_7411,N_5969);
or UO_133 (O_133,N_7517,N_9809);
nor UO_134 (O_134,N_7263,N_6406);
nand UO_135 (O_135,N_6236,N_5378);
nor UO_136 (O_136,N_8688,N_5785);
and UO_137 (O_137,N_9306,N_6857);
or UO_138 (O_138,N_7388,N_7361);
nand UO_139 (O_139,N_8357,N_8139);
nor UO_140 (O_140,N_6842,N_9908);
nor UO_141 (O_141,N_6641,N_8622);
or UO_142 (O_142,N_7071,N_5464);
nor UO_143 (O_143,N_9529,N_9069);
nand UO_144 (O_144,N_9567,N_5477);
or UO_145 (O_145,N_5337,N_8086);
nor UO_146 (O_146,N_9506,N_7122);
nand UO_147 (O_147,N_5542,N_7401);
nor UO_148 (O_148,N_9651,N_5864);
nor UO_149 (O_149,N_5722,N_6189);
or UO_150 (O_150,N_9985,N_5351);
xor UO_151 (O_151,N_8407,N_7735);
nand UO_152 (O_152,N_7377,N_8778);
xor UO_153 (O_153,N_5780,N_7198);
nand UO_154 (O_154,N_5104,N_8861);
xnor UO_155 (O_155,N_8142,N_7613);
nor UO_156 (O_156,N_5718,N_8000);
and UO_157 (O_157,N_8532,N_8913);
or UO_158 (O_158,N_8540,N_5708);
nor UO_159 (O_159,N_5452,N_5361);
nor UO_160 (O_160,N_9671,N_9099);
nand UO_161 (O_161,N_6578,N_9065);
or UO_162 (O_162,N_6727,N_9337);
nand UO_163 (O_163,N_7333,N_8550);
or UO_164 (O_164,N_6295,N_9165);
nand UO_165 (O_165,N_8342,N_5080);
nand UO_166 (O_166,N_9285,N_5283);
and UO_167 (O_167,N_8247,N_7798);
and UO_168 (O_168,N_6396,N_5046);
nand UO_169 (O_169,N_7319,N_7574);
or UO_170 (O_170,N_9212,N_9093);
nand UO_171 (O_171,N_5357,N_8197);
or UO_172 (O_172,N_5027,N_7021);
nor UO_173 (O_173,N_7324,N_9848);
nor UO_174 (O_174,N_7310,N_7468);
or UO_175 (O_175,N_7030,N_9615);
nor UO_176 (O_176,N_8629,N_5224);
nand UO_177 (O_177,N_5794,N_8177);
nor UO_178 (O_178,N_9439,N_8218);
or UO_179 (O_179,N_6657,N_8371);
and UO_180 (O_180,N_9140,N_6012);
and UO_181 (O_181,N_6746,N_9504);
nand UO_182 (O_182,N_5050,N_6374);
xor UO_183 (O_183,N_8771,N_7371);
and UO_184 (O_184,N_8307,N_9361);
nand UO_185 (O_185,N_6556,N_9983);
and UO_186 (O_186,N_5116,N_6170);
nand UO_187 (O_187,N_8812,N_7304);
nand UO_188 (O_188,N_5389,N_6399);
and UO_189 (O_189,N_6554,N_5279);
or UO_190 (O_190,N_7428,N_9334);
nand UO_191 (O_191,N_6888,N_8908);
or UO_192 (O_192,N_9917,N_8743);
nor UO_193 (O_193,N_7437,N_7339);
nand UO_194 (O_194,N_5113,N_8832);
and UO_195 (O_195,N_8620,N_5316);
nor UO_196 (O_196,N_5557,N_6387);
or UO_197 (O_197,N_8345,N_5787);
or UO_198 (O_198,N_5558,N_7249);
nor UO_199 (O_199,N_7515,N_7913);
nor UO_200 (O_200,N_6262,N_9963);
and UO_201 (O_201,N_9343,N_6778);
nand UO_202 (O_202,N_5788,N_8687);
or UO_203 (O_203,N_5863,N_7653);
and UO_204 (O_204,N_7392,N_9625);
and UO_205 (O_205,N_6504,N_7539);
nand UO_206 (O_206,N_9468,N_6716);
nor UO_207 (O_207,N_5480,N_9060);
nor UO_208 (O_208,N_8462,N_6428);
nor UO_209 (O_209,N_8581,N_6536);
nor UO_210 (O_210,N_9139,N_9974);
or UO_211 (O_211,N_6272,N_5686);
and UO_212 (O_212,N_6796,N_8732);
and UO_213 (O_213,N_6081,N_5133);
xor UO_214 (O_214,N_5296,N_7692);
and UO_215 (O_215,N_6783,N_7159);
nor UO_216 (O_216,N_6198,N_6082);
nand UO_217 (O_217,N_6823,N_6397);
and UO_218 (O_218,N_7119,N_5892);
or UO_219 (O_219,N_6099,N_5995);
xor UO_220 (O_220,N_6575,N_6526);
and UO_221 (O_221,N_9847,N_7942);
nand UO_222 (O_222,N_6415,N_9328);
and UO_223 (O_223,N_6535,N_8315);
and UO_224 (O_224,N_6280,N_9941);
and UO_225 (O_225,N_8038,N_7323);
nor UO_226 (O_226,N_9696,N_7098);
or UO_227 (O_227,N_7037,N_7124);
and UO_228 (O_228,N_8836,N_6157);
nand UO_229 (O_229,N_6178,N_5295);
nor UO_230 (O_230,N_8783,N_7421);
or UO_231 (O_231,N_9735,N_9017);
and UO_232 (O_232,N_8353,N_6046);
nor UO_233 (O_233,N_8431,N_6179);
or UO_234 (O_234,N_9283,N_7876);
or UO_235 (O_235,N_5216,N_8069);
nand UO_236 (O_236,N_9547,N_9172);
nor UO_237 (O_237,N_8131,N_8169);
or UO_238 (O_238,N_6597,N_7418);
xor UO_239 (O_239,N_6734,N_9533);
and UO_240 (O_240,N_5803,N_8652);
nand UO_241 (O_241,N_5840,N_9229);
and UO_242 (O_242,N_8394,N_9879);
or UO_243 (O_243,N_5450,N_7463);
or UO_244 (O_244,N_5244,N_5330);
nor UO_245 (O_245,N_9119,N_9505);
and UO_246 (O_246,N_7181,N_5977);
and UO_247 (O_247,N_8330,N_9429);
and UO_248 (O_248,N_9571,N_5880);
nand UO_249 (O_249,N_7171,N_7887);
nor UO_250 (O_250,N_9300,N_8376);
or UO_251 (O_251,N_5957,N_9907);
nand UO_252 (O_252,N_7559,N_7328);
and UO_253 (O_253,N_5314,N_7658);
and UO_254 (O_254,N_6065,N_8616);
or UO_255 (O_255,N_8722,N_7248);
nand UO_256 (O_256,N_5564,N_9428);
nor UO_257 (O_257,N_6963,N_7257);
nor UO_258 (O_258,N_5022,N_5693);
and UO_259 (O_259,N_7127,N_8595);
nand UO_260 (O_260,N_7812,N_6119);
or UO_261 (O_261,N_9549,N_5029);
nand UO_262 (O_262,N_5365,N_6688);
or UO_263 (O_263,N_5201,N_5689);
nand UO_264 (O_264,N_9978,N_7830);
or UO_265 (O_265,N_8813,N_8157);
nand UO_266 (O_266,N_9777,N_8979);
or UO_267 (O_267,N_9487,N_9824);
or UO_268 (O_268,N_8564,N_6450);
nor UO_269 (O_269,N_8424,N_9975);
or UO_270 (O_270,N_5559,N_6066);
or UO_271 (O_271,N_8103,N_5836);
nor UO_272 (O_272,N_6579,N_6190);
nand UO_273 (O_273,N_9245,N_8106);
and UO_274 (O_274,N_9660,N_7811);
and UO_275 (O_275,N_7983,N_5073);
nor UO_276 (O_276,N_6323,N_9164);
and UO_277 (O_277,N_8676,N_5070);
or UO_278 (O_278,N_8530,N_9909);
nor UO_279 (O_279,N_6429,N_7829);
nand UO_280 (O_280,N_6890,N_6978);
nand UO_281 (O_281,N_9108,N_9776);
nor UO_282 (O_282,N_7980,N_8740);
or UO_283 (O_283,N_5344,N_9349);
or UO_284 (O_284,N_8229,N_8145);
nand UO_285 (O_285,N_6912,N_7836);
and UO_286 (O_286,N_7964,N_6829);
or UO_287 (O_287,N_7084,N_7817);
nor UO_288 (O_288,N_8526,N_9682);
nand UO_289 (O_289,N_7020,N_9626);
and UO_290 (O_290,N_8890,N_5930);
nand UO_291 (O_291,N_9161,N_6084);
nor UO_292 (O_292,N_8677,N_6223);
nand UO_293 (O_293,N_9684,N_8830);
nor UO_294 (O_294,N_9787,N_5301);
and UO_295 (O_295,N_6988,N_7760);
nor UO_296 (O_296,N_7746,N_9702);
or UO_297 (O_297,N_5488,N_6530);
and UO_298 (O_298,N_7738,N_5047);
nor UO_299 (O_299,N_8961,N_5397);
nor UO_300 (O_300,N_9236,N_7381);
and UO_301 (O_301,N_6411,N_9856);
nand UO_302 (O_302,N_8848,N_8084);
and UO_303 (O_303,N_6673,N_8624);
and UO_304 (O_304,N_9162,N_9182);
and UO_305 (O_305,N_8309,N_8772);
or UO_306 (O_306,N_6229,N_9620);
or UO_307 (O_307,N_5161,N_9650);
or UO_308 (O_308,N_9143,N_5877);
or UO_309 (O_309,N_9348,N_6814);
nand UO_310 (O_310,N_9135,N_7360);
and UO_311 (O_311,N_9159,N_8338);
and UO_312 (O_312,N_8443,N_7082);
nand UO_313 (O_313,N_8588,N_6033);
and UO_314 (O_314,N_6701,N_9261);
or UO_315 (O_315,N_8865,N_7890);
or UO_316 (O_316,N_5229,N_7605);
nand UO_317 (O_317,N_7771,N_7314);
nand UO_318 (O_318,N_6160,N_6040);
and UO_319 (O_319,N_9636,N_8067);
nand UO_320 (O_320,N_9779,N_7837);
and UO_321 (O_321,N_7601,N_9604);
nand UO_322 (O_322,N_9480,N_9719);
and UO_323 (O_323,N_6770,N_6413);
nand UO_324 (O_324,N_8448,N_6102);
and UO_325 (O_325,N_6699,N_6671);
or UO_326 (O_326,N_9724,N_8188);
nor UO_327 (O_327,N_9818,N_5723);
nand UO_328 (O_328,N_7644,N_7734);
nor UO_329 (O_329,N_5158,N_6968);
nor UO_330 (O_330,N_8450,N_6570);
and UO_331 (O_331,N_9826,N_7307);
nor UO_332 (O_332,N_9964,N_7897);
nor UO_333 (O_333,N_8579,N_7679);
nor UO_334 (O_334,N_5382,N_8754);
and UO_335 (O_335,N_7224,N_7351);
or UO_336 (O_336,N_6966,N_5119);
nand UO_337 (O_337,N_8318,N_9386);
or UO_338 (O_338,N_6547,N_8976);
or UO_339 (O_339,N_5440,N_6290);
nor UO_340 (O_340,N_5850,N_9396);
or UO_341 (O_341,N_8617,N_5797);
or UO_342 (O_342,N_7172,N_7461);
nor UO_343 (O_343,N_6317,N_5500);
or UO_344 (O_344,N_9123,N_5436);
and UO_345 (O_345,N_7444,N_6754);
xor UO_346 (O_346,N_8880,N_8416);
nand UO_347 (O_347,N_9572,N_6691);
or UO_348 (O_348,N_6712,N_8187);
nor UO_349 (O_349,N_5808,N_6334);
and UO_350 (O_350,N_8520,N_8355);
nor UO_351 (O_351,N_8986,N_6861);
or UO_352 (O_352,N_7067,N_5293);
or UO_353 (O_353,N_9448,N_6409);
nand UO_354 (O_354,N_8876,N_8502);
and UO_355 (O_355,N_6445,N_6121);
nand UO_356 (O_356,N_8459,N_9296);
and UO_357 (O_357,N_5493,N_6337);
and UO_358 (O_358,N_6386,N_8105);
nor UO_359 (O_359,N_8236,N_7597);
nand UO_360 (O_360,N_9117,N_6837);
nor UO_361 (O_361,N_8874,N_9688);
nand UO_362 (O_362,N_6195,N_6430);
or UO_363 (O_363,N_7460,N_8974);
or UO_364 (O_364,N_6956,N_9738);
nor UO_365 (O_365,N_7174,N_5530);
and UO_366 (O_366,N_8418,N_7009);
and UO_367 (O_367,N_7979,N_9575);
nor UO_368 (O_368,N_9055,N_5105);
nor UO_369 (O_369,N_6439,N_7179);
and UO_370 (O_370,N_6478,N_8078);
or UO_371 (O_371,N_8938,N_5174);
nand UO_372 (O_372,N_5813,N_9500);
or UO_373 (O_373,N_9633,N_7277);
nand UO_374 (O_374,N_9874,N_5885);
nand UO_375 (O_375,N_5144,N_7784);
nor UO_376 (O_376,N_8774,N_6497);
or UO_377 (O_377,N_7167,N_6466);
xor UO_378 (O_378,N_8109,N_6293);
and UO_379 (O_379,N_6967,N_8005);
nand UO_380 (O_380,N_6053,N_9998);
or UO_381 (O_381,N_9725,N_8634);
nand UO_382 (O_382,N_8920,N_9276);
xnor UO_383 (O_383,N_9622,N_5745);
nand UO_384 (O_384,N_9196,N_9648);
nor UO_385 (O_385,N_9273,N_9493);
nand UO_386 (O_386,N_9319,N_8580);
or UO_387 (O_387,N_7218,N_7270);
or UO_388 (O_388,N_8499,N_5846);
and UO_389 (O_389,N_6362,N_7593);
and UO_390 (O_390,N_5453,N_5095);
and UO_391 (O_391,N_7034,N_7010);
or UO_392 (O_392,N_8958,N_6586);
or UO_393 (O_393,N_6867,N_9409);
and UO_394 (O_394,N_5830,N_5189);
nand UO_395 (O_395,N_8007,N_9808);
and UO_396 (O_396,N_5967,N_7937);
or UO_397 (O_397,N_8985,N_6222);
nand UO_398 (O_398,N_7778,N_5349);
nor UO_399 (O_399,N_7240,N_6731);
or UO_400 (O_400,N_5373,N_8685);
or UO_401 (O_401,N_6714,N_7241);
and UO_402 (O_402,N_8434,N_6088);
nand UO_403 (O_403,N_7620,N_9745);
and UO_404 (O_404,N_9061,N_5792);
nor UO_405 (O_405,N_5381,N_6392);
nor UO_406 (O_406,N_8563,N_7335);
and UO_407 (O_407,N_8326,N_6924);
nand UO_408 (O_408,N_8288,N_9837);
nand UO_409 (O_409,N_9095,N_9982);
or UO_410 (O_410,N_8587,N_6241);
nor UO_411 (O_411,N_9372,N_9652);
nand UO_412 (O_412,N_7814,N_5601);
or UO_413 (O_413,N_9792,N_9010);
or UO_414 (O_414,N_5690,N_8381);
nor UO_415 (O_415,N_8669,N_6540);
or UO_416 (O_416,N_7434,N_6140);
or UO_417 (O_417,N_5310,N_8973);
or UO_418 (O_418,N_9871,N_8544);
nor UO_419 (O_419,N_9566,N_9552);
or UO_420 (O_420,N_8811,N_9027);
or UO_421 (O_421,N_6931,N_9758);
nand UO_422 (O_422,N_6418,N_5007);
or UO_423 (O_423,N_7946,N_6339);
nor UO_424 (O_424,N_5081,N_8691);
nor UO_425 (O_425,N_5188,N_5683);
nor UO_426 (O_426,N_8183,N_6156);
nor UO_427 (O_427,N_7666,N_5076);
and UO_428 (O_428,N_9953,N_7378);
nand UO_429 (O_429,N_5560,N_8398);
nand UO_430 (O_430,N_9811,N_6758);
or UO_431 (O_431,N_8590,N_8648);
nand UO_432 (O_432,N_8348,N_7029);
or UO_433 (O_433,N_8368,N_7816);
or UO_434 (O_434,N_7772,N_8382);
nand UO_435 (O_435,N_8966,N_6732);
nand UO_436 (O_436,N_6192,N_6690);
and UO_437 (O_437,N_8210,N_8932);
nand UO_438 (O_438,N_8356,N_9867);
nand UO_439 (O_439,N_7853,N_8768);
or UO_440 (O_440,N_8599,N_5747);
or UO_441 (O_441,N_5739,N_9038);
and UO_442 (O_442,N_5783,N_5700);
nand UO_443 (O_443,N_7112,N_5255);
nor UO_444 (O_444,N_6382,N_6945);
nand UO_445 (O_445,N_7289,N_7226);
and UO_446 (O_446,N_9388,N_5992);
or UO_447 (O_447,N_9384,N_8004);
nor UO_448 (O_448,N_8181,N_6709);
nor UO_449 (O_449,N_7849,N_5842);
nand UO_450 (O_450,N_5715,N_8467);
and UO_451 (O_451,N_5066,N_6555);
nand UO_452 (O_452,N_6289,N_8668);
and UO_453 (O_453,N_7788,N_8301);
and UO_454 (O_454,N_8383,N_6344);
or UO_455 (O_455,N_6191,N_7316);
and UO_456 (O_456,N_5417,N_6373);
nor UO_457 (O_457,N_9325,N_8070);
nor UO_458 (O_458,N_7042,N_5471);
nor UO_459 (O_459,N_9841,N_9621);
nand UO_460 (O_460,N_8441,N_9025);
or UO_461 (O_461,N_7057,N_6166);
and UO_462 (O_462,N_7366,N_6454);
or UO_463 (O_463,N_9708,N_5385);
and UO_464 (O_464,N_7242,N_6388);
nor UO_465 (O_465,N_7509,N_8928);
and UO_466 (O_466,N_7178,N_6314);
nor UO_467 (O_467,N_5807,N_5388);
and UO_468 (O_468,N_9473,N_9205);
nand UO_469 (O_469,N_5320,N_9986);
nor UO_470 (O_470,N_7901,N_7394);
or UO_471 (O_471,N_8905,N_7116);
and UO_472 (O_472,N_8859,N_7683);
nand UO_473 (O_473,N_6992,N_8130);
nor UO_474 (O_474,N_8637,N_8548);
and UO_475 (O_475,N_7967,N_8175);
or UO_476 (O_476,N_8295,N_8763);
nor UO_477 (O_477,N_7611,N_7825);
and UO_478 (O_478,N_7985,N_9743);
and UO_479 (O_479,N_9062,N_8377);
xnor UO_480 (O_480,N_9214,N_5267);
or UO_481 (O_481,N_5582,N_5795);
nand UO_482 (O_482,N_7504,N_5525);
or UO_483 (O_483,N_9374,N_8346);
or UO_484 (O_484,N_6826,N_5644);
and UO_485 (O_485,N_8207,N_9227);
nor UO_486 (O_486,N_8366,N_9459);
nor UO_487 (O_487,N_5634,N_7820);
nor UO_488 (O_488,N_9812,N_6664);
xor UO_489 (O_489,N_8308,N_5231);
and UO_490 (O_490,N_7861,N_7221);
nand UO_491 (O_491,N_5094,N_7631);
and UO_492 (O_492,N_8283,N_5526);
or UO_493 (O_493,N_6868,N_8887);
nand UO_494 (O_494,N_6475,N_9959);
and UO_495 (O_495,N_8931,N_9440);
or UO_496 (O_496,N_6562,N_8090);
or UO_497 (O_497,N_7672,N_6258);
nand UO_498 (O_498,N_5882,N_8079);
nor UO_499 (O_499,N_6713,N_6298);
nor UO_500 (O_500,N_8625,N_6126);
nor UO_501 (O_501,N_7469,N_5649);
nor UO_502 (O_502,N_5975,N_7899);
nand UO_503 (O_503,N_9729,N_5872);
nor UO_504 (O_504,N_6364,N_7975);
or UO_505 (O_505,N_6326,N_7779);
and UO_506 (O_506,N_8760,N_7194);
and UO_507 (O_507,N_7888,N_5124);
or UO_508 (O_508,N_8320,N_5261);
nand UO_509 (O_509,N_9085,N_7900);
nor UO_510 (O_510,N_5049,N_5306);
nand UO_511 (O_511,N_9160,N_7303);
and UO_512 (O_512,N_9731,N_8826);
nand UO_513 (O_513,N_6325,N_9316);
and UO_514 (O_514,N_6790,N_6644);
and UO_515 (O_515,N_9426,N_5544);
xnor UO_516 (O_516,N_5653,N_7005);
nand UO_517 (O_517,N_9435,N_5988);
or UO_518 (O_518,N_9375,N_8927);
or UO_519 (O_519,N_9855,N_6989);
xnor UO_520 (O_520,N_6933,N_9966);
nand UO_521 (O_521,N_8445,N_6542);
nand UO_522 (O_522,N_5110,N_9376);
xor UO_523 (O_523,N_7134,N_8902);
or UO_524 (O_524,N_7639,N_5533);
nand UO_525 (O_525,N_9427,N_6895);
or UO_526 (O_526,N_7364,N_9835);
nor UO_527 (O_527,N_6075,N_7222);
or UO_528 (O_528,N_9206,N_5139);
and UO_529 (O_529,N_6167,N_9023);
nand UO_530 (O_530,N_9888,N_6076);
or UO_531 (O_531,N_6549,N_8263);
and UO_532 (O_532,N_7527,N_7600);
nor UO_533 (O_533,N_7462,N_6899);
or UO_534 (O_534,N_6932,N_9070);
nand UO_535 (O_535,N_6464,N_7199);
and UO_536 (O_536,N_6960,N_9987);
and UO_537 (O_537,N_6648,N_6271);
and UO_538 (O_538,N_9067,N_7781);
and UO_539 (O_539,N_5638,N_9443);
or UO_540 (O_540,N_7299,N_6089);
and UO_541 (O_541,N_7802,N_6383);
and UO_542 (O_542,N_9994,N_7928);
and UO_543 (O_543,N_6771,N_9786);
or UO_544 (O_544,N_5604,N_8017);
or UO_545 (O_545,N_6164,N_9484);
and UO_546 (O_546,N_5984,N_5387);
nor UO_547 (O_547,N_9332,N_9329);
nand UO_548 (O_548,N_8592,N_7996);
and UO_549 (O_549,N_9613,N_5876);
nor UO_550 (O_550,N_9931,N_8200);
nor UO_551 (O_551,N_6427,N_7748);
or UO_552 (O_552,N_8765,N_8511);
nor UO_553 (O_553,N_8259,N_7884);
nand UO_554 (O_554,N_6043,N_7024);
nand UO_555 (O_555,N_6090,N_8650);
nand UO_556 (O_556,N_6990,N_5669);
xor UO_557 (O_557,N_8148,N_6291);
nor UO_558 (O_558,N_9167,N_6986);
nor UO_559 (O_559,N_5630,N_9659);
and UO_560 (O_560,N_5481,N_6035);
nand UO_561 (O_561,N_5346,N_9903);
nor UO_562 (O_562,N_7585,N_9488);
or UO_563 (O_563,N_5777,N_7558);
and UO_564 (O_564,N_9886,N_7384);
nor UO_565 (O_565,N_6557,N_9104);
nor UO_566 (O_566,N_5259,N_9420);
nand UO_567 (O_567,N_9532,N_5991);
nand UO_568 (O_568,N_9118,N_6467);
nor UO_569 (O_569,N_9795,N_6629);
nand UO_570 (O_570,N_5776,N_5097);
nand UO_571 (O_571,N_8882,N_8313);
or UO_572 (O_572,N_5575,N_7219);
nand UO_573 (O_573,N_8680,N_7729);
nor UO_574 (O_574,N_8739,N_8195);
and UO_575 (O_575,N_6896,N_8710);
and UO_576 (O_576,N_9312,N_5672);
or UO_577 (O_577,N_6403,N_5045);
nor UO_578 (O_578,N_6071,N_7810);
nand UO_579 (O_579,N_7195,N_5976);
or UO_580 (O_580,N_7997,N_5228);
nor UO_581 (O_581,N_6692,N_7821);
and UO_582 (O_582,N_7208,N_5516);
or UO_583 (O_583,N_9260,N_7245);
and UO_584 (O_584,N_7091,N_5288);
and UO_585 (O_585,N_9149,N_6889);
and UO_586 (O_586,N_5455,N_5405);
nand UO_587 (O_587,N_9692,N_9073);
nand UO_588 (O_588,N_7808,N_9494);
nor UO_589 (O_589,N_8745,N_8846);
nand UO_590 (O_590,N_6275,N_8693);
nand UO_591 (O_591,N_6571,N_9145);
and UO_592 (O_592,N_7768,N_9098);
nand UO_593 (O_593,N_9230,N_7133);
nand UO_594 (O_594,N_7447,N_6036);
nand UO_595 (O_595,N_5590,N_7571);
and UO_596 (O_596,N_5937,N_8002);
or UO_597 (O_597,N_7851,N_6821);
nand UO_598 (O_598,N_5875,N_9658);
and UO_599 (O_599,N_6352,N_7896);
nand UO_600 (O_600,N_7976,N_9407);
nand UO_601 (O_601,N_5676,N_6022);
and UO_602 (O_602,N_5246,N_9127);
nand UO_603 (O_603,N_7362,N_7511);
and UO_604 (O_604,N_6761,N_6728);
nand UO_605 (O_605,N_8065,N_7846);
and UO_606 (O_606,N_9289,N_6108);
nor UO_607 (O_607,N_9339,N_7169);
nor UO_608 (O_608,N_8567,N_6026);
and UO_609 (O_609,N_5328,N_9510);
or UO_610 (O_610,N_7992,N_8948);
and UO_611 (O_611,N_9585,N_8964);
xnor UO_612 (O_612,N_7243,N_5614);
nor UO_613 (O_613,N_9347,N_5867);
nand UO_614 (O_614,N_8699,N_8611);
xnor UO_615 (O_615,N_6904,N_9195);
or UO_616 (O_616,N_6566,N_7457);
xnor UO_617 (O_617,N_8930,N_5716);
and UO_618 (O_618,N_6885,N_7950);
nor UO_619 (O_619,N_5593,N_6221);
nand UO_620 (O_620,N_6580,N_9244);
or UO_621 (O_621,N_9665,N_5814);
nand UO_622 (O_622,N_9796,N_8606);
or UO_623 (O_623,N_5861,N_7652);
or UO_624 (O_624,N_6602,N_5239);
nand UO_625 (O_625,N_8369,N_5462);
or UO_626 (O_626,N_8191,N_8967);
nand UO_627 (O_627,N_8239,N_5423);
nor UO_628 (O_628,N_5832,N_6928);
and UO_629 (O_629,N_6651,N_8665);
nand UO_630 (O_630,N_5323,N_6112);
or UO_631 (O_631,N_8490,N_5497);
or UO_632 (O_632,N_8437,N_9255);
nor UO_633 (O_633,N_5865,N_7630);
xor UO_634 (O_634,N_6524,N_9223);
or UO_635 (O_635,N_7787,N_9181);
or UO_636 (O_636,N_8432,N_6433);
xnor UO_637 (O_637,N_5458,N_6753);
nor UO_638 (O_638,N_6110,N_7287);
nand UO_639 (O_639,N_5643,N_7018);
and UO_640 (O_640,N_8303,N_5862);
and UO_641 (O_641,N_5652,N_7891);
nor UO_642 (O_642,N_8149,N_7547);
and UO_643 (O_643,N_6196,N_5537);
or UO_644 (O_644,N_8998,N_8790);
xnor UO_645 (O_645,N_9358,N_5063);
and UO_646 (O_646,N_5541,N_7908);
or UO_647 (O_647,N_9579,N_9521);
or UO_648 (O_648,N_7485,N_9377);
and UO_649 (O_649,N_8276,N_6134);
nand UO_650 (O_650,N_6836,N_9716);
nand UO_651 (O_651,N_6656,N_9142);
or UO_652 (O_652,N_9870,N_7988);
nor UO_653 (O_653,N_8286,N_5569);
and UO_654 (O_654,N_7340,N_7094);
xnor UO_655 (O_655,N_5147,N_5921);
and UO_656 (O_656,N_5784,N_7706);
nor UO_657 (O_657,N_7562,N_6902);
nor UO_658 (O_658,N_6500,N_5146);
nand UO_659 (O_659,N_6689,N_7390);
and UO_660 (O_660,N_5412,N_7142);
nor UO_661 (O_661,N_8658,N_7530);
nor UO_662 (O_662,N_7845,N_8267);
or UO_663 (O_663,N_7696,N_5127);
or UO_664 (O_664,N_9894,N_9690);
nor UO_665 (O_665,N_8248,N_9737);
or UO_666 (O_666,N_6985,N_7046);
nand UO_667 (O_667,N_5810,N_8655);
nand UO_668 (O_668,N_5510,N_6784);
or UO_669 (O_669,N_7905,N_7583);
or UO_670 (O_670,N_8212,N_8531);
nor UO_671 (O_671,N_9454,N_6316);
or UO_672 (O_672,N_5543,N_7490);
nor UO_673 (O_673,N_7535,N_5730);
nor UO_674 (O_674,N_9596,N_8776);
or UO_675 (O_675,N_5741,N_7635);
or UO_676 (O_676,N_5499,N_6938);
or UO_677 (O_677,N_8799,N_7623);
nor UO_678 (O_678,N_9744,N_9077);
or UO_679 (O_679,N_5535,N_9460);
nand UO_680 (O_680,N_5496,N_5233);
or UO_681 (O_681,N_5627,N_8934);
nor UO_682 (O_682,N_5947,N_5278);
nor UO_683 (O_683,N_6582,N_5353);
or UO_684 (O_684,N_9989,N_5790);
nand UO_685 (O_685,N_5230,N_5399);
nand UO_686 (O_686,N_5696,N_8695);
nor UO_687 (O_687,N_6583,N_8896);
nor UO_688 (O_688,N_8037,N_8654);
and UO_689 (O_689,N_5732,N_6158);
or UO_690 (O_690,N_9518,N_5631);
and UO_691 (O_691,N_5178,N_8147);
nand UO_692 (O_692,N_8909,N_6006);
or UO_693 (O_693,N_6060,N_5737);
or UO_694 (O_694,N_5597,N_6054);
and UO_695 (O_695,N_7684,N_5042);
and UO_696 (O_696,N_6563,N_6748);
nand UO_697 (O_697,N_7336,N_5195);
nor UO_698 (O_698,N_7141,N_8155);
and UO_699 (O_699,N_5245,N_7725);
or UO_700 (O_700,N_9057,N_5704);
nor UO_701 (O_701,N_6407,N_8226);
and UO_702 (O_702,N_7294,N_6735);
nor UO_703 (O_703,N_8995,N_8088);
and UO_704 (O_704,N_6993,N_9187);
and UO_705 (O_705,N_9045,N_8682);
nand UO_706 (O_706,N_9634,N_7028);
or UO_707 (O_707,N_5668,N_5052);
nor UO_708 (O_708,N_5023,N_7196);
nor UO_709 (O_709,N_9043,N_6007);
or UO_710 (O_710,N_7262,N_6419);
or UO_711 (O_711,N_9565,N_6064);
or UO_712 (O_712,N_5857,N_5610);
or UO_713 (O_713,N_6087,N_5828);
or UO_714 (O_714,N_8649,N_8657);
nand UO_715 (O_715,N_7582,N_6080);
nand UO_716 (O_716,N_9563,N_8250);
or UO_717 (O_717,N_6702,N_7508);
nor UO_718 (O_718,N_5657,N_8129);
nand UO_719 (O_719,N_9993,N_9185);
nor UO_720 (O_720,N_8980,N_6341);
or UO_721 (O_721,N_5871,N_8297);
and UO_722 (O_722,N_5152,N_5319);
and UO_723 (O_723,N_6462,N_5096);
nor UO_724 (O_724,N_5305,N_5411);
and UO_725 (O_725,N_8294,N_8942);
or UO_726 (O_726,N_7286,N_9655);
nor UO_727 (O_727,N_5036,N_7948);
and UO_728 (O_728,N_5251,N_9417);
or UO_729 (O_729,N_7592,N_5160);
nor UO_730 (O_730,N_7676,N_5756);
or UO_731 (O_731,N_5519,N_5384);
or UO_732 (O_732,N_8408,N_7602);
or UO_733 (O_733,N_5343,N_5617);
nor UO_734 (O_734,N_7528,N_9803);
xnor UO_735 (O_735,N_8917,N_9669);
nand UO_736 (O_736,N_8870,N_7393);
or UO_737 (O_737,N_6502,N_5987);
nor UO_738 (O_738,N_8469,N_7331);
nand UO_739 (O_739,N_7726,N_7086);
nand UO_740 (O_740,N_9810,N_5075);
and UO_741 (O_741,N_7634,N_6908);
and UO_742 (O_742,N_9208,N_9216);
nand UO_743 (O_743,N_8957,N_5368);
nand UO_744 (O_744,N_7298,N_8275);
and UO_745 (O_745,N_7070,N_9389);
nor UO_746 (O_746,N_5299,N_8008);
and UO_747 (O_747,N_5200,N_9200);
nor UO_748 (O_748,N_5887,N_8798);
or UO_749 (O_749,N_6977,N_7283);
or UO_750 (O_750,N_9307,N_7715);
or UO_751 (O_751,N_9106,N_6655);
nor UO_752 (O_752,N_5895,N_6017);
xor UO_753 (O_753,N_8252,N_9556);
and UO_754 (O_754,N_7664,N_6704);
nor UO_755 (O_755,N_8350,N_7341);
or UO_756 (O_756,N_6560,N_8324);
or UO_757 (O_757,N_7795,N_8971);
nand UO_758 (O_758,N_7835,N_6417);
nand UO_759 (O_759,N_7939,N_6883);
nor UO_760 (O_760,N_6971,N_5182);
and UO_761 (O_761,N_7907,N_7158);
or UO_762 (O_762,N_5153,N_5179);
and UO_763 (O_763,N_9477,N_7281);
or UO_764 (O_764,N_7682,N_8711);
nand UO_765 (O_765,N_8752,N_5933);
and UO_766 (O_766,N_7480,N_7809);
nand UO_767 (O_767,N_7702,N_9971);
and UO_768 (O_768,N_8113,N_7302);
nor UO_769 (O_769,N_9103,N_9110);
or UO_770 (O_770,N_8857,N_6009);
xnor UO_771 (O_771,N_8429,N_6514);
and UO_772 (O_772,N_9387,N_9806);
and UO_773 (O_773,N_6870,N_9400);
or UO_774 (O_774,N_6706,N_5505);
nor UO_775 (O_775,N_9015,N_9561);
or UO_776 (O_776,N_7747,N_9595);
nor UO_777 (O_777,N_5469,N_8897);
or UO_778 (O_778,N_5433,N_9201);
nor UO_779 (O_779,N_9872,N_8568);
nor UO_780 (O_780,N_8795,N_7823);
nand UO_781 (O_781,N_7618,N_5621);
or UO_782 (O_782,N_7165,N_8881);
nor UO_783 (O_783,N_7864,N_8015);
nor UO_784 (O_784,N_7560,N_7410);
and UO_785 (O_785,N_8347,N_9270);
or UO_786 (O_786,N_8314,N_9829);
or UO_787 (O_787,N_8910,N_7176);
nor UO_788 (O_788,N_5072,N_7207);
and UO_789 (O_789,N_8955,N_7625);
nand UO_790 (O_790,N_6328,N_6869);
nand UO_791 (O_791,N_7163,N_5061);
and UO_792 (O_792,N_6983,N_6068);
nand UO_793 (O_793,N_8554,N_9345);
nand UO_794 (O_794,N_8725,N_8602);
nand UO_795 (O_795,N_7521,N_6744);
and UO_796 (O_796,N_9791,N_9969);
and UO_797 (O_797,N_6234,N_7854);
or UO_798 (O_798,N_6810,N_9988);
and UO_799 (O_799,N_6646,N_9537);
nor UO_800 (O_800,N_8993,N_6276);
or UO_801 (O_801,N_6146,N_6529);
xor UO_802 (O_802,N_5694,N_6833);
or UO_803 (O_803,N_5931,N_5017);
or UO_804 (O_804,N_6911,N_5609);
or UO_805 (O_805,N_8605,N_7466);
or UO_806 (O_806,N_5905,N_8290);
nand UO_807 (O_807,N_7677,N_5107);
or UO_808 (O_808,N_7069,N_9709);
nor UO_809 (O_809,N_5837,N_7429);
or UO_810 (O_810,N_5013,N_8061);
nand UO_811 (O_811,N_8481,N_5376);
and UO_812 (O_812,N_7292,N_5983);
or UO_813 (O_813,N_6456,N_5623);
nor UO_814 (O_814,N_5005,N_7741);
or UO_815 (O_815,N_8989,N_7933);
xor UO_816 (O_816,N_5587,N_6347);
and UO_817 (O_817,N_9609,N_6197);
nand UO_818 (O_818,N_5434,N_8742);
nand UO_819 (O_819,N_7761,N_7416);
or UO_820 (O_820,N_6097,N_6366);
nor UO_821 (O_821,N_6852,N_7633);
nor UO_822 (O_822,N_6543,N_7235);
nand UO_823 (O_823,N_8736,N_5102);
nor UO_824 (O_824,N_8464,N_8273);
or UO_825 (O_825,N_9156,N_5521);
or UO_826 (O_826,N_5130,N_9335);
and UO_827 (O_827,N_7470,N_8255);
nand UO_828 (O_828,N_6740,N_7713);
nor UO_829 (O_829,N_5035,N_9834);
or UO_830 (O_830,N_6848,N_7016);
nand UO_831 (O_831,N_7865,N_6131);
or UO_832 (O_832,N_5125,N_6098);
nor UO_833 (O_833,N_6016,N_5596);
nand UO_834 (O_834,N_7822,N_5898);
or UO_835 (O_835,N_7140,N_9036);
nand UO_836 (O_836,N_8335,N_8517);
nor UO_837 (O_837,N_7205,N_6957);
nor UO_838 (O_838,N_8058,N_6375);
and UO_839 (O_839,N_5264,N_5819);
or UO_840 (O_840,N_5742,N_6311);
nor UO_841 (O_841,N_6019,N_7902);
nor UO_842 (O_842,N_8340,N_8954);
xor UO_843 (O_843,N_5083,N_6052);
or UO_844 (O_844,N_7088,N_8102);
and UO_845 (O_845,N_7960,N_6920);
or UO_846 (O_846,N_8547,N_8364);
or UO_847 (O_847,N_8496,N_8686);
or UO_848 (O_848,N_5034,N_6550);
nand UO_849 (O_849,N_8044,N_8101);
xor UO_850 (O_850,N_9775,N_9930);
or UO_851 (O_851,N_6384,N_6807);
and UO_852 (O_852,N_7234,N_8052);
or UO_853 (O_853,N_8287,N_7342);
nor UO_854 (O_854,N_6935,N_6752);
nor UO_855 (O_855,N_7923,N_6939);
or UO_856 (O_856,N_6892,N_5284);
or UO_857 (O_857,N_6370,N_9763);
or UO_858 (O_858,N_6654,N_8641);
or UO_859 (O_859,N_5974,N_9752);
nor UO_860 (O_860,N_7089,N_9188);
and UO_861 (O_861,N_5079,N_8251);
or UO_862 (O_862,N_5547,N_9321);
or UO_863 (O_863,N_8104,N_8878);
or UO_864 (O_864,N_9132,N_7931);
and UO_865 (O_865,N_7995,N_6569);
nor UO_866 (O_866,N_9483,N_5752);
nand UO_867 (O_867,N_5600,N_5329);
and UO_868 (O_868,N_5912,N_8316);
nor UO_869 (O_869,N_7125,N_7796);
and UO_870 (O_870,N_6256,N_8405);
or UO_871 (O_871,N_8844,N_9006);
nand UO_872 (O_872,N_9839,N_5549);
nor UO_873 (O_873,N_9174,N_7524);
nor UO_874 (O_874,N_8991,N_6995);
and UO_875 (O_875,N_9075,N_5806);
nor UO_876 (O_876,N_6991,N_9574);
nor UO_877 (O_877,N_9148,N_9924);
and UO_878 (O_878,N_5919,N_7744);
nor UO_879 (O_879,N_6395,N_6002);
and UO_880 (O_880,N_9495,N_6819);
nor UO_881 (O_881,N_9177,N_9915);
nor UO_882 (O_882,N_6521,N_6446);
and UO_883 (O_883,N_5581,N_5907);
or UO_884 (O_884,N_8521,N_6136);
or UO_885 (O_885,N_8003,N_7038);
nor UO_886 (O_886,N_8533,N_9683);
and UO_887 (O_887,N_6503,N_8724);
or UO_888 (O_888,N_8562,N_5173);
nor UO_889 (O_889,N_6161,N_8926);
nor UO_890 (O_890,N_9814,N_7044);
nor UO_891 (O_891,N_9653,N_7595);
or UO_892 (O_892,N_7252,N_7727);
nor UO_893 (O_893,N_9904,N_7433);
or UO_894 (O_894,N_8321,N_9865);
and UO_895 (O_895,N_8825,N_6340);
nor UO_896 (O_896,N_8842,N_9646);
and UO_897 (O_897,N_9782,N_5953);
nor UO_898 (O_898,N_9525,N_9415);
or UO_899 (O_899,N_5618,N_6608);
and UO_900 (O_900,N_8427,N_6058);
nor UO_901 (O_901,N_8504,N_8898);
nand UO_902 (O_902,N_7432,N_8838);
or UO_903 (O_903,N_9406,N_6211);
and UO_904 (O_904,N_9024,N_8225);
nand UO_905 (O_905,N_8161,N_5767);
nand UO_906 (O_906,N_9594,N_6185);
nand UO_907 (O_907,N_5685,N_7993);
and UO_908 (O_908,N_7250,N_8636);
nand UO_909 (O_909,N_7565,N_9961);
nand UO_910 (O_910,N_7649,N_6801);
nor UO_911 (O_911,N_5199,N_6520);
and UO_912 (O_912,N_5735,N_9718);
nand UO_913 (O_913,N_8675,N_5936);
nand UO_914 (O_914,N_6305,N_5755);
or UO_915 (O_915,N_8862,N_5055);
xnor UO_916 (O_916,N_7671,N_6114);
or UO_917 (O_917,N_5691,N_8945);
xnor UO_918 (O_918,N_8497,N_9326);
or UO_919 (O_919,N_9364,N_6169);
nand UO_920 (O_920,N_9661,N_6494);
nor UO_921 (O_921,N_7472,N_9863);
and UO_922 (O_922,N_5266,N_8758);
nand UO_923 (O_923,N_5498,N_5175);
nor UO_924 (O_924,N_8679,N_8091);
xnor UO_925 (O_925,N_9338,N_9717);
xor UO_926 (O_926,N_6679,N_6335);
nor UO_927 (O_927,N_9922,N_7386);
nand UO_928 (O_928,N_8108,N_6313);
and UO_929 (O_929,N_8486,N_9889);
nand UO_930 (O_930,N_6152,N_6231);
nor UO_931 (O_931,N_9150,N_9662);
nor UO_932 (O_932,N_6061,N_7152);
nor UO_933 (O_933,N_9864,N_7007);
or UO_934 (O_934,N_6532,N_8831);
and UO_935 (O_935,N_6303,N_7452);
nand UO_936 (O_936,N_7420,N_5044);
or UO_937 (O_937,N_8343,N_8500);
nand UO_938 (O_938,N_8264,N_8096);
nor UO_939 (O_939,N_5269,N_5941);
or UO_940 (O_940,N_8277,N_9960);
or UO_941 (O_941,N_9990,N_5647);
nand UO_942 (O_942,N_5646,N_5068);
and UO_943 (O_943,N_7769,N_9721);
and UO_944 (O_944,N_5402,N_6910);
or UO_945 (O_945,N_7448,N_6561);
and UO_946 (O_946,N_6719,N_5951);
or UO_947 (O_947,N_6310,N_6610);
or UO_948 (O_948,N_6511,N_6820);
or UO_949 (O_949,N_9751,N_5911);
nor UO_950 (O_950,N_5217,N_9047);
nand UO_951 (O_951,N_5071,N_7577);
nand UO_952 (O_952,N_6951,N_6492);
and UO_953 (O_953,N_7719,N_8262);
or UO_954 (O_954,N_9044,N_8626);
and UO_955 (O_955,N_7126,N_5506);
and UO_956 (O_956,N_9447,N_8570);
nor UO_957 (O_957,N_5746,N_5502);
or UO_958 (O_958,N_8222,N_6270);
or UO_959 (O_959,N_6934,N_8428);
xnor UO_960 (O_960,N_5731,N_7819);
nor UO_961 (O_961,N_5972,N_6105);
nor UO_962 (O_962,N_8516,N_7797);
nor UO_963 (O_963,N_7843,N_6903);
or UO_964 (O_964,N_6668,N_8189);
nor UO_965 (O_965,N_9040,N_8135);
nor UO_966 (O_966,N_5802,N_6943);
and UO_967 (O_967,N_6422,N_7483);
nor UO_968 (O_968,N_9292,N_6906);
nand UO_969 (O_969,N_5854,N_9471);
nand UO_970 (O_970,N_7743,N_5532);
nor UO_971 (O_971,N_6459,N_9355);
nor UO_972 (O_972,N_6138,N_6587);
or UO_973 (O_973,N_6001,N_5720);
nand UO_974 (O_974,N_8393,N_9336);
or UO_975 (O_975,N_9654,N_5403);
nand UO_976 (O_976,N_8156,N_5773);
and UO_977 (O_977,N_8618,N_6632);
or UO_978 (O_978,N_5311,N_7587);
or UO_979 (O_979,N_7703,N_7523);
nand UO_980 (O_980,N_6078,N_5352);
nand UO_981 (O_981,N_8701,N_6442);
nand UO_982 (O_982,N_8228,N_6285);
nor UO_983 (O_983,N_6013,N_8172);
nor UO_984 (O_984,N_6369,N_5913);
and UO_985 (O_985,N_8999,N_6441);
nor UO_986 (O_986,N_8397,N_6787);
nor UO_987 (O_987,N_8460,N_6470);
xor UO_988 (O_988,N_7233,N_6723);
and UO_989 (O_989,N_8940,N_7764);
or UO_990 (O_990,N_7246,N_9972);
and UO_991 (O_991,N_8193,N_6327);
nor UO_992 (O_992,N_5663,N_6259);
and UO_993 (O_993,N_9753,N_8048);
or UO_994 (O_994,N_9869,N_6321);
and UO_995 (O_995,N_5292,N_6021);
or UO_996 (O_996,N_8788,N_8583);
and UO_997 (O_997,N_7309,N_5467);
or UO_998 (O_998,N_8209,N_5815);
nor UO_999 (O_999,N_5226,N_5552);
and UO_1000 (O_1000,N_6453,N_5563);
and UO_1001 (O_1001,N_7408,N_9825);
and UO_1002 (O_1002,N_7166,N_9936);
or UO_1003 (O_1003,N_6962,N_8981);
nor UO_1004 (O_1004,N_8982,N_9918);
nor UO_1005 (O_1005,N_8747,N_7000);
and UO_1006 (O_1006,N_5655,N_5565);
nand UO_1007 (O_1007,N_9189,N_6508);
nand UO_1008 (O_1008,N_9833,N_5089);
nor UO_1009 (O_1009,N_8205,N_8615);
nor UO_1010 (O_1010,N_8704,N_5286);
or UO_1011 (O_1011,N_7102,N_8391);
nand UO_1012 (O_1012,N_6278,N_5414);
nor UO_1013 (O_1013,N_7612,N_9305);
and UO_1014 (O_1014,N_7971,N_6483);
or UO_1015 (O_1015,N_7708,N_5128);
or UO_1016 (O_1016,N_5041,N_8133);
nor UO_1017 (O_1017,N_9628,N_9144);
nand UO_1018 (O_1018,N_7237,N_8173);
nor UO_1019 (O_1019,N_9938,N_5774);
or UO_1020 (O_1020,N_9049,N_7954);
and UO_1021 (O_1021,N_7427,N_8871);
or UO_1022 (O_1022,N_6964,N_5078);
nand UO_1023 (O_1023,N_8243,N_6795);
or UO_1024 (O_1024,N_6631,N_9790);
nand UO_1025 (O_1025,N_8950,N_6639);
nand UO_1026 (O_1026,N_9284,N_6914);
nor UO_1027 (O_1027,N_8514,N_8835);
nand UO_1028 (O_1028,N_8107,N_5721);
nand UO_1029 (O_1029,N_9707,N_6391);
or UO_1030 (O_1030,N_9382,N_7146);
or UO_1031 (O_1031,N_9588,N_7330);
nand UO_1032 (O_1032,N_5207,N_9598);
nor UO_1033 (O_1033,N_5062,N_6636);
and UO_1034 (O_1034,N_9220,N_7934);
and UO_1035 (O_1035,N_6858,N_6248);
and UO_1036 (O_1036,N_9513,N_8696);
nand UO_1037 (O_1037,N_9516,N_5594);
nand UO_1038 (O_1038,N_5366,N_7721);
or UO_1039 (O_1039,N_9211,N_5324);
or UO_1040 (O_1040,N_6048,N_9082);
or UO_1041 (O_1041,N_6025,N_7150);
and UO_1042 (O_1042,N_8400,N_9294);
or UO_1043 (O_1043,N_7615,N_9304);
and UO_1044 (O_1044,N_9266,N_7261);
nand UO_1045 (O_1045,N_7927,N_5345);
and UO_1046 (O_1046,N_6283,N_5507);
nand UO_1047 (O_1047,N_5446,N_8663);
nor UO_1048 (O_1048,N_8387,N_6918);
and UO_1049 (O_1049,N_5332,N_7687);
nor UO_1050 (O_1050,N_7092,N_5100);
and UO_1051 (O_1051,N_7075,N_7862);
and UO_1052 (O_1052,N_8116,N_5379);
nor UO_1053 (O_1053,N_9842,N_5122);
or UO_1054 (O_1054,N_7391,N_8232);
nand UO_1055 (O_1055,N_7757,N_9000);
and UO_1056 (O_1056,N_7940,N_9462);
nor UO_1057 (O_1057,N_5626,N_8671);
and UO_1058 (O_1058,N_8203,N_9687);
nor UO_1059 (O_1059,N_9178,N_9507);
or UO_1060 (O_1060,N_5008,N_8578);
nand UO_1061 (O_1061,N_8843,N_9515);
nor UO_1062 (O_1062,N_6447,N_8442);
nor UO_1063 (O_1063,N_7449,N_7347);
nand UO_1064 (O_1064,N_7765,N_5736);
or UO_1065 (O_1065,N_6643,N_6175);
nor UO_1066 (O_1066,N_5438,N_8026);
nand UO_1067 (O_1067,N_7930,N_7526);
xnor UO_1068 (O_1068,N_9056,N_5847);
and UO_1069 (O_1069,N_9706,N_7828);
or UO_1070 (O_1070,N_5183,N_6135);
nand UO_1071 (O_1071,N_5336,N_7128);
and UO_1072 (O_1072,N_7129,N_6182);
xnor UO_1073 (O_1073,N_6484,N_5335);
and UO_1074 (O_1074,N_9771,N_9068);
or UO_1075 (O_1075,N_8414,N_9222);
and UO_1076 (O_1076,N_5702,N_6847);
or UO_1077 (O_1077,N_6125,N_7518);
or UO_1078 (O_1078,N_5561,N_8138);
and UO_1079 (O_1079,N_6351,N_5291);
and UO_1080 (O_1080,N_8194,N_9949);
nor UO_1081 (O_1081,N_6940,N_6150);
nand UO_1082 (O_1082,N_6501,N_5567);
or UO_1083 (O_1083,N_5670,N_7870);
or UO_1084 (O_1084,N_7004,N_7686);
nor UO_1085 (O_1085,N_9739,N_8244);
nand UO_1086 (O_1086,N_5294,N_6739);
and UO_1087 (O_1087,N_5297,N_6479);
nand UO_1088 (O_1088,N_6537,N_8339);
nand UO_1089 (O_1089,N_5010,N_9955);
or UO_1090 (O_1090,N_9410,N_7534);
nor UO_1091 (O_1091,N_9243,N_6916);
nand UO_1092 (O_1092,N_9880,N_6558);
nor UO_1093 (O_1093,N_6301,N_8723);
and UO_1094 (O_1094,N_9367,N_9623);
nor UO_1095 (O_1095,N_9458,N_7701);
or UO_1096 (O_1096,N_7651,N_8093);
nand UO_1097 (O_1097,N_7343,N_8190);
nor UO_1098 (O_1098,N_9933,N_8589);
and UO_1099 (O_1099,N_6871,N_6785);
nand UO_1100 (O_1100,N_6779,N_8328);
and UO_1101 (O_1101,N_5131,N_9416);
or UO_1102 (O_1102,N_6880,N_7355);
nor UO_1103 (O_1103,N_5589,N_9293);
and UO_1104 (O_1104,N_7584,N_5562);
or UO_1105 (O_1105,N_9821,N_7380);
nand UO_1106 (O_1106,N_8012,N_6350);
nor UO_1107 (O_1107,N_5408,N_5529);
nand UO_1108 (O_1108,N_9631,N_7570);
and UO_1109 (O_1109,N_5851,N_8735);
and UO_1110 (O_1110,N_8341,N_9906);
or UO_1111 (O_1111,N_6063,N_7162);
nand UO_1112 (O_1112,N_5628,N_6047);
nor UO_1113 (O_1113,N_7621,N_8660);
or UO_1114 (O_1114,N_5666,N_7399);
and UO_1115 (O_1115,N_8850,N_7935);
or UO_1116 (O_1116,N_9126,N_8215);
nor UO_1117 (O_1117,N_9340,N_9380);
or UO_1118 (O_1118,N_7061,N_9090);
and UO_1119 (O_1119,N_9910,N_9578);
nor UO_1120 (O_1120,N_5823,N_7395);
or UO_1121 (O_1121,N_9942,N_6124);
nand UO_1122 (O_1122,N_9072,N_9469);
or UO_1123 (O_1123,N_8047,N_6461);
nor UO_1124 (O_1124,N_5461,N_8018);
nor UO_1125 (O_1125,N_7767,N_7451);
and UO_1126 (O_1126,N_6506,N_7068);
nor UO_1127 (O_1127,N_8417,N_9939);
or UO_1128 (O_1128,N_7272,N_9968);
and UO_1129 (O_1129,N_9733,N_6365);
or UO_1130 (O_1130,N_5949,N_9597);
nand UO_1131 (O_1131,N_5883,N_5074);
nand UO_1132 (O_1132,N_7027,N_8852);
nor UO_1133 (O_1133,N_5422,N_9330);
or UO_1134 (O_1134,N_8608,N_5622);
and UO_1135 (O_1135,N_8488,N_5914);
nor UO_1136 (O_1136,N_7680,N_8901);
nand UO_1137 (O_1137,N_7264,N_9762);
nand UO_1138 (O_1138,N_8238,N_9861);
and UO_1139 (O_1139,N_5383,N_5354);
or UO_1140 (O_1140,N_6905,N_5943);
or UO_1141 (O_1141,N_5415,N_6917);
and UO_1142 (O_1142,N_9385,N_7952);
nor UO_1143 (O_1143,N_5342,N_9446);
nand UO_1144 (O_1144,N_7847,N_8501);
or UO_1145 (O_1145,N_8363,N_9011);
and UO_1146 (O_1146,N_8392,N_9052);
nor UO_1147 (O_1147,N_7573,N_6855);
and UO_1148 (O_1148,N_6813,N_9005);
and UO_1149 (O_1149,N_5274,N_8136);
nand UO_1150 (O_1150,N_8575,N_9531);
or UO_1151 (O_1151,N_6941,N_6539);
or UO_1152 (O_1152,N_5524,N_5809);
nor UO_1153 (O_1153,N_5348,N_7989);
nand UO_1154 (O_1154,N_6872,N_8918);
nor UO_1155 (O_1155,N_8604,N_9042);
nor UO_1156 (O_1156,N_6594,N_7636);
nand UO_1157 (O_1157,N_7453,N_5156);
nor UO_1158 (O_1158,N_6854,N_5019);
or UO_1159 (O_1159,N_7581,N_5833);
nor UO_1160 (O_1160,N_6412,N_7911);
nand UO_1161 (O_1161,N_8118,N_8153);
and UO_1162 (O_1162,N_8716,N_8666);
or UO_1163 (O_1163,N_8171,N_9503);
or UO_1164 (O_1164,N_5109,N_5154);
or UO_1165 (O_1165,N_5359,N_6118);
nand UO_1166 (O_1166,N_9722,N_6997);
and UO_1167 (O_1167,N_6923,N_7740);
nor UO_1168 (O_1168,N_8071,N_9180);
or UO_1169 (O_1169,N_6206,N_5327);
nor UO_1170 (O_1170,N_6685,N_6318);
and UO_1171 (O_1171,N_6385,N_8401);
nand UO_1172 (O_1172,N_8095,N_6024);
nor UO_1173 (O_1173,N_6677,N_6319);
or UO_1174 (O_1174,N_8184,N_6846);
or UO_1175 (O_1175,N_7938,N_7153);
or UO_1176 (O_1176,N_9028,N_8479);
or UO_1177 (O_1177,N_8123,N_7054);
and UO_1178 (O_1178,N_7803,N_6589);
or UO_1179 (O_1179,N_9766,N_5315);
or UO_1180 (O_1180,N_5375,N_5303);
and UO_1181 (O_1181,N_9134,N_8681);
or UO_1182 (O_1182,N_7647,N_9301);
or UO_1183 (O_1183,N_8291,N_8576);
nor UO_1184 (O_1184,N_7922,N_8024);
nand UO_1185 (O_1185,N_6645,N_5258);
or UO_1186 (O_1186,N_8060,N_6612);
nand UO_1187 (O_1187,N_8329,N_6463);
nor UO_1188 (O_1188,N_5660,N_6684);
or UO_1189 (O_1189,N_5744,N_7213);
or UO_1190 (O_1190,N_5724,N_5571);
or UO_1191 (O_1191,N_6232,N_8762);
or UO_1192 (O_1192,N_8332,N_6282);
or UO_1193 (O_1193,N_5509,N_9616);
xor UO_1194 (O_1194,N_9878,N_5990);
and UO_1195 (O_1195,N_9951,N_7970);
nand UO_1196 (O_1196,N_8528,N_8182);
and UO_1197 (O_1197,N_6162,N_9170);
nand UO_1198 (O_1198,N_6982,N_9715);
and UO_1199 (O_1199,N_8351,N_5699);
nor UO_1200 (O_1200,N_6155,N_6205);
nand UO_1201 (O_1201,N_5712,N_5270);
nand UO_1202 (O_1202,N_8433,N_9433);
nand UO_1203 (O_1203,N_6062,N_8869);
or UO_1204 (O_1204,N_6623,N_8534);
and UO_1205 (O_1205,N_9666,N_6884);
nand UO_1206 (O_1206,N_8389,N_6621);
nor UO_1207 (O_1207,N_7430,N_6830);
or UO_1208 (O_1208,N_8062,N_5753);
nor UO_1209 (O_1209,N_9215,N_7439);
and UO_1210 (O_1210,N_7863,N_8610);
or UO_1211 (O_1211,N_5038,N_8465);
nor UO_1212 (O_1212,N_5858,N_5416);
and UO_1213 (O_1213,N_9538,N_9642);
and UO_1214 (O_1214,N_6666,N_6667);
or UO_1215 (O_1215,N_7419,N_5845);
nand UO_1216 (O_1216,N_8922,N_8556);
nand UO_1217 (O_1217,N_6177,N_9760);
nand UO_1218 (O_1218,N_6838,N_9249);
nand UO_1219 (O_1219,N_7512,N_8727);
and UO_1220 (O_1220,N_6817,N_9274);
nand UO_1221 (O_1221,N_9600,N_6972);
nand UO_1222 (O_1222,N_9287,N_5138);
or UO_1223 (O_1223,N_7731,N_5554);
or UO_1224 (O_1224,N_5701,N_9183);
nor UO_1225 (O_1225,N_7137,N_7051);
or UO_1226 (O_1226,N_6320,N_7957);
or UO_1227 (O_1227,N_7614,N_9109);
nor UO_1228 (O_1228,N_7267,N_5799);
nand UO_1229 (O_1229,N_5595,N_6193);
nand UO_1230 (O_1230,N_6181,N_5016);
nor UO_1231 (O_1231,N_8423,N_5751);
nand UO_1232 (O_1232,N_5599,N_6083);
and UO_1233 (O_1233,N_7596,N_5629);
and UO_1234 (O_1234,N_8227,N_8787);
and UO_1235 (O_1235,N_6831,N_9158);
and UO_1236 (O_1236,N_7694,N_8403);
and UO_1237 (O_1237,N_8741,N_5103);
nand UO_1238 (O_1238,N_5922,N_6457);
or UO_1239 (O_1239,N_8992,N_7608);
nor UO_1240 (O_1240,N_5678,N_8372);
nor UO_1241 (O_1241,N_7714,N_9602);
and UO_1242 (O_1242,N_8935,N_9558);
and UO_1243 (O_1243,N_9481,N_6669);
or UO_1244 (O_1244,N_5486,N_9232);
nand UO_1245 (O_1245,N_5162,N_6086);
nor UO_1246 (O_1246,N_5796,N_7450);
or UO_1247 (O_1247,N_8325,N_8282);
nor UO_1248 (O_1248,N_7737,N_7185);
nand UO_1249 (O_1249,N_7003,N_7598);
nand UO_1250 (O_1250,N_5640,N_9524);
or UO_1251 (O_1251,N_7561,N_5221);
nand UO_1252 (O_1252,N_9772,N_6210);
or UO_1253 (O_1253,N_8847,N_6242);
nand UO_1254 (O_1254,N_8028,N_9441);
nor UO_1255 (O_1255,N_5213,N_9219);
or UO_1256 (O_1256,N_5468,N_7465);
nand UO_1257 (O_1257,N_9318,N_6425);
or UO_1258 (O_1258,N_7403,N_8883);
nand UO_1259 (O_1259,N_7145,N_7332);
and UO_1260 (O_1260,N_8492,N_8804);
nor UO_1261 (O_1261,N_6800,N_8770);
nand UO_1262 (O_1262,N_7223,N_5998);
and UO_1263 (O_1263,N_7852,N_6094);
nand UO_1264 (O_1264,N_6769,N_5252);
nor UO_1265 (O_1265,N_7925,N_6402);
or UO_1266 (O_1266,N_9370,N_6309);
or UO_1267 (O_1267,N_8965,N_5084);
nor UO_1268 (O_1268,N_7074,N_7346);
nand UO_1269 (O_1269,N_9202,N_8025);
nand UO_1270 (O_1270,N_7079,N_8779);
or UO_1271 (O_1271,N_8885,N_9606);
nor UO_1272 (O_1272,N_5275,N_9550);
nand UO_1273 (O_1273,N_6372,N_5856);
and UO_1274 (O_1274,N_9333,N_5282);
and UO_1275 (O_1275,N_5860,N_9290);
nand UO_1276 (O_1276,N_8098,N_6224);
nor UO_1277 (O_1277,N_7972,N_9553);
nor UO_1278 (O_1278,N_7063,N_6815);
nor UO_1279 (O_1279,N_9852,N_9858);
or UO_1280 (O_1280,N_6519,N_6183);
or UO_1281 (O_1281,N_9875,N_9365);
xnor UO_1282 (O_1282,N_9768,N_5419);
nor UO_1283 (O_1283,N_9499,N_5069);
and UO_1284 (O_1284,N_5115,N_7259);
or UO_1285 (O_1285,N_7880,N_7698);
nand UO_1286 (O_1286,N_7555,N_7023);
and UO_1287 (O_1287,N_6864,N_7032);
xor UO_1288 (O_1288,N_6130,N_6715);
xnor UO_1289 (O_1289,N_7442,N_8551);
and UO_1290 (O_1290,N_7986,N_8737);
nor UO_1291 (O_1291,N_6465,N_8164);
or UO_1292 (O_1292,N_9136,N_6851);
or UO_1293 (O_1293,N_8706,N_9204);
nand UO_1294 (O_1294,N_8767,N_6634);
nand UO_1295 (O_1295,N_9950,N_5959);
nor UO_1296 (O_1296,N_8162,N_9601);
nor UO_1297 (O_1297,N_8056,N_9562);
nand UO_1298 (O_1298,N_6828,N_5778);
nand UO_1299 (O_1299,N_9071,N_8246);
or UO_1300 (O_1300,N_9381,N_9793);
nand UO_1301 (O_1301,N_7372,N_5180);
xnor UO_1302 (O_1302,N_6665,N_5762);
nand UO_1303 (O_1303,N_5980,N_7373);
and UO_1304 (O_1304,N_9418,N_5606);
nor UO_1305 (O_1305,N_7106,N_8174);
nand UO_1306 (O_1306,N_9252,N_7860);
nor UO_1307 (O_1307,N_7288,N_5350);
and UO_1308 (O_1308,N_6947,N_8794);
nor UO_1309 (O_1309,N_6472,N_7327);
nand UO_1310 (O_1310,N_8659,N_6405);
nor UO_1311 (O_1311,N_6533,N_8027);
nor UO_1312 (O_1312,N_5576,N_6239);
and UO_1313 (O_1313,N_9080,N_5485);
and UO_1314 (O_1314,N_5651,N_9436);
or UO_1315 (O_1315,N_6774,N_7085);
nor UO_1316 (O_1316,N_5059,N_6738);
nand UO_1317 (O_1317,N_5859,N_9397);
nand UO_1318 (O_1318,N_7790,N_9836);
xnor UO_1319 (O_1319,N_5548,N_7750);
or UO_1320 (O_1320,N_5968,N_8046);
nor UO_1321 (O_1321,N_9944,N_7657);
and UO_1322 (O_1322,N_6050,N_7920);
or UO_1323 (O_1323,N_5738,N_8344);
or UO_1324 (O_1324,N_7188,N_5060);
nor UO_1325 (O_1325,N_6762,N_8254);
or UO_1326 (O_1326,N_5664,N_5934);
nand UO_1327 (O_1327,N_6929,N_8081);
nand UO_1328 (O_1328,N_8756,N_6876);
nand UO_1329 (O_1329,N_5944,N_7446);
nand UO_1330 (O_1330,N_8125,N_9122);
and UO_1331 (O_1331,N_8970,N_8311);
or UO_1332 (O_1332,N_9542,N_6100);
nor UO_1333 (O_1333,N_6252,N_5771);
and UO_1334 (O_1334,N_9645,N_7275);
nor UO_1335 (O_1335,N_6984,N_5926);
or UO_1336 (O_1336,N_8010,N_9742);
nand UO_1337 (O_1337,N_9007,N_8508);
or UO_1338 (O_1338,N_6306,N_7398);
nand UO_1339 (O_1339,N_5902,N_5087);
nand UO_1340 (O_1340,N_9357,N_8543);
or UO_1341 (O_1341,N_9590,N_5592);
nor UO_1342 (O_1342,N_9569,N_5527);
nand UO_1343 (O_1343,N_7350,N_5026);
nand UO_1344 (O_1344,N_8087,N_7161);
or UO_1345 (O_1345,N_8435,N_9587);
nand UO_1346 (O_1346,N_8444,N_6615);
and UO_1347 (O_1347,N_5811,N_7033);
nor UO_1348 (O_1348,N_7123,N_5025);
nor UO_1349 (O_1349,N_8378,N_6055);
nor UO_1350 (O_1350,N_8839,N_7961);
nor UO_1351 (O_1351,N_5717,N_7732);
nand UO_1352 (O_1352,N_9253,N_8092);
and UO_1353 (O_1353,N_5454,N_6622);
or UO_1354 (O_1354,N_5012,N_6998);
nor UO_1355 (O_1355,N_6286,N_7542);
and UO_1356 (O_1356,N_9536,N_8352);
or UO_1357 (O_1357,N_7906,N_7369);
nor UO_1358 (O_1358,N_5789,N_8717);
or UO_1359 (O_1359,N_5897,N_5169);
and UO_1360 (O_1360,N_7047,N_7282);
nor UO_1361 (O_1361,N_8390,N_6773);
nand UO_1362 (O_1362,N_8030,N_9854);
nand UO_1363 (O_1363,N_7320,N_7855);
or UO_1364 (O_1364,N_7675,N_8258);
and UO_1365 (O_1365,N_7312,N_6788);
nand UO_1366 (O_1366,N_7793,N_7197);
nor UO_1367 (O_1367,N_7318,N_5271);
or UO_1368 (O_1368,N_6245,N_8411);
or UO_1369 (O_1369,N_7697,N_8996);
nand UO_1370 (O_1370,N_6944,N_8969);
and UO_1371 (O_1371,N_6137,N_9391);
and UO_1372 (O_1372,N_7055,N_8016);
xor UO_1373 (O_1373,N_7498,N_9911);
or UO_1374 (O_1374,N_6371,N_9125);
nand UO_1375 (O_1375,N_8596,N_7209);
nand UO_1376 (O_1376,N_7139,N_8134);
nor UO_1377 (O_1377,N_9734,N_9618);
nand UO_1378 (O_1378,N_5954,N_5441);
nor UO_1379 (O_1379,N_9476,N_5491);
and UO_1380 (O_1380,N_6777,N_9539);
nand UO_1381 (O_1381,N_9474,N_7104);
and UO_1382 (O_1382,N_7156,N_5393);
nor UO_1383 (O_1383,N_5684,N_5302);
and UO_1384 (O_1384,N_7755,N_8815);
and UO_1385 (O_1385,N_8841,N_9614);
nor UO_1386 (O_1386,N_6129,N_8296);
or UO_1387 (O_1387,N_7646,N_8073);
xnor UO_1388 (O_1388,N_7689,N_9627);
and UO_1389 (O_1389,N_9091,N_7754);
or UO_1390 (O_1390,N_7097,N_6014);
nand UO_1391 (O_1391,N_5518,N_9054);
nor UO_1392 (O_1392,N_6721,N_7567);
nor UO_1393 (O_1393,N_6505,N_5665);
xnor UO_1394 (O_1394,N_9203,N_5157);
nand UO_1395 (O_1395,N_7187,N_9778);
xnor UO_1396 (O_1396,N_5205,N_5171);
and UO_1397 (O_1397,N_9128,N_6693);
nand UO_1398 (O_1398,N_8638,N_6925);
and UO_1399 (O_1399,N_7643,N_6151);
or UO_1400 (O_1400,N_9896,N_9413);
and UO_1401 (O_1401,N_5935,N_9551);
and UO_1402 (O_1402,N_7497,N_9438);
or UO_1403 (O_1403,N_6538,N_5479);
or UO_1404 (O_1404,N_8614,N_7254);
nand UO_1405 (O_1405,N_6541,N_6452);
nor UO_1406 (O_1406,N_7025,N_8466);
nor UO_1407 (O_1407,N_7968,N_9408);
nor UO_1408 (O_1408,N_7580,N_9850);
and UO_1409 (O_1409,N_5698,N_5321);
and UO_1410 (O_1410,N_5650,N_8719);
nand UO_1411 (O_1411,N_5826,N_8984);
nor UO_1412 (O_1412,N_9213,N_6499);
or UO_1413 (O_1413,N_8535,N_6675);
xnor UO_1414 (O_1414,N_7723,N_6128);
and UO_1415 (O_1415,N_6886,N_6041);
nand UO_1416 (O_1416,N_7081,N_8994);
nor UO_1417 (O_1417,N_5611,N_6353);
nand UO_1418 (O_1418,N_8854,N_8698);
or UO_1419 (O_1419,N_7295,N_6603);
nor UO_1420 (O_1420,N_5996,N_6741);
or UO_1421 (O_1421,N_8440,N_6638);
nand UO_1422 (O_1422,N_7875,N_7238);
or UO_1423 (O_1423,N_9251,N_5248);
and UO_1424 (O_1424,N_7707,N_7578);
nand UO_1425 (O_1425,N_7916,N_5040);
and UO_1426 (O_1426,N_9859,N_9714);
nor UO_1427 (O_1427,N_6841,N_5225);
and UO_1428 (O_1428,N_7078,N_8600);
nor UO_1429 (O_1429,N_6768,N_5487);
nand UO_1430 (O_1430,N_7918,N_9797);
or UO_1431 (O_1431,N_7591,N_7160);
nand UO_1432 (O_1432,N_5456,N_9298);
nand UO_1433 (O_1433,N_6284,N_7266);
nand UO_1434 (O_1434,N_8829,N_7990);
nand UO_1435 (O_1435,N_6737,N_5822);
and UO_1436 (O_1436,N_6432,N_5713);
nand UO_1437 (O_1437,N_5939,N_9761);
and UO_1438 (O_1438,N_9121,N_9663);
and UO_1439 (O_1439,N_7762,N_8785);
or UO_1440 (O_1440,N_6042,N_6824);
nand UO_1441 (O_1441,N_7505,N_8281);
nor UO_1442 (O_1442,N_5636,N_5360);
or UO_1443 (O_1443,N_6249,N_6618);
or UO_1444 (O_1444,N_9916,N_6596);
or UO_1445 (O_1445,N_8415,N_7663);
and UO_1446 (O_1446,N_7441,N_8302);
and UO_1447 (O_1447,N_7783,N_7859);
nor UO_1448 (O_1448,N_8128,N_6736);
or UO_1449 (O_1449,N_9378,N_9309);
nor UO_1450 (O_1450,N_7624,N_9467);
nor UO_1451 (O_1451,N_6605,N_7915);
and UO_1452 (O_1452,N_8630,N_7440);
and UO_1453 (O_1453,N_7536,N_9780);
and UO_1454 (O_1454,N_5613,N_9713);
nor UO_1455 (O_1455,N_6187,N_5938);
nor UO_1456 (O_1456,N_6515,N_9945);
and UO_1457 (O_1457,N_8111,N_8802);
and UO_1458 (O_1458,N_9923,N_7955);
and UO_1459 (O_1459,N_8260,N_5743);
nor UO_1460 (O_1460,N_9548,N_5966);
nor UO_1461 (O_1461,N_5483,N_5276);
nor UO_1462 (O_1462,N_5263,N_7353);
and UO_1463 (O_1463,N_6390,N_9295);
or UO_1464 (O_1464,N_6616,N_8198);
and UO_1465 (O_1465,N_6101,N_9929);
and UO_1466 (O_1466,N_5839,N_9900);
or UO_1467 (O_1467,N_5878,N_5793);
nor UO_1468 (O_1468,N_7035,N_8234);
nand UO_1469 (O_1469,N_7118,N_6297);
and UO_1470 (O_1470,N_5431,N_9184);
nand UO_1471 (O_1471,N_8268,N_9063);
and UO_1472 (O_1472,N_6207,N_7186);
or UO_1473 (O_1473,N_7045,N_9101);
nand UO_1474 (O_1474,N_9235,N_5304);
or UO_1475 (O_1475,N_9535,N_5272);
and UO_1476 (O_1476,N_9689,N_5340);
nor UO_1477 (O_1477,N_5903,N_6805);
and UO_1478 (O_1478,N_8925,N_7766);
nor UO_1479 (O_1479,N_7753,N_8990);
nand UO_1480 (O_1480,N_9699,N_8085);
and UO_1481 (O_1481,N_8879,N_5203);
xor UO_1482 (O_1482,N_6875,N_7638);
nand UO_1483 (O_1483,N_5504,N_7367);
and UO_1484 (O_1484,N_6059,N_8653);
nand UO_1485 (O_1485,N_6711,N_9492);
and UO_1486 (O_1486,N_8042,N_7269);
and UO_1487 (O_1487,N_5247,N_8455);
and UO_1488 (O_1488,N_6468,N_6144);
nand UO_1489 (O_1489,N_6775,N_5172);
and UO_1490 (O_1490,N_7858,N_6717);
nor UO_1491 (O_1491,N_8895,N_9895);
or UO_1492 (O_1492,N_7872,N_5002);
or UO_1493 (O_1493,N_5448,N_7244);
or UO_1494 (O_1494,N_5827,N_7645);
or UO_1495 (O_1495,N_6626,N_5918);
nor UO_1496 (O_1496,N_6363,N_8020);
or UO_1497 (O_1497,N_7239,N_6444);
and UO_1498 (O_1498,N_6845,N_6919);
or UO_1499 (O_1499,N_7958,N_6897);
endmodule