module basic_3000_30000_3500_15_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_1736,In_2978);
or U1 (N_1,In_1616,In_533);
xor U2 (N_2,In_1200,In_813);
or U3 (N_3,In_2129,In_858);
nand U4 (N_4,In_783,In_2728);
xor U5 (N_5,In_728,In_1256);
xor U6 (N_6,In_2551,In_970);
nor U7 (N_7,In_1229,In_653);
or U8 (N_8,In_1781,In_1040);
and U9 (N_9,In_560,In_1545);
xnor U10 (N_10,In_878,In_2482);
xnor U11 (N_11,In_1336,In_1236);
nand U12 (N_12,In_850,In_932);
and U13 (N_13,In_2508,In_1377);
or U14 (N_14,In_790,In_677);
nand U15 (N_15,In_1885,In_111);
nand U16 (N_16,In_629,In_2647);
or U17 (N_17,In_2128,In_1217);
xnor U18 (N_18,In_2297,In_191);
nor U19 (N_19,In_1532,In_639);
and U20 (N_20,In_1536,In_2102);
or U21 (N_21,In_325,In_1913);
or U22 (N_22,In_458,In_730);
nor U23 (N_23,In_2154,In_2717);
xnor U24 (N_24,In_206,In_1013);
nor U25 (N_25,In_1588,In_2502);
xnor U26 (N_26,In_1655,In_1467);
xnor U27 (N_27,In_1740,In_269);
or U28 (N_28,In_1441,In_364);
xnor U29 (N_29,In_1832,In_358);
nand U30 (N_30,In_2181,In_2877);
nor U31 (N_31,In_2976,In_225);
and U32 (N_32,In_2490,In_354);
or U33 (N_33,In_1291,In_1857);
nor U34 (N_34,In_2776,In_2320);
nor U35 (N_35,In_809,In_1366);
nor U36 (N_36,In_1898,In_1714);
nor U37 (N_37,In_2291,In_2783);
nor U38 (N_38,In_1828,In_2930);
nand U39 (N_39,In_1850,In_507);
nor U40 (N_40,In_2423,In_285);
nand U41 (N_41,In_2131,In_2959);
nor U42 (N_42,In_2414,In_769);
and U43 (N_43,In_1841,In_2180);
nor U44 (N_44,In_1919,In_2556);
nor U45 (N_45,In_2521,In_569);
and U46 (N_46,In_1868,In_1665);
nor U47 (N_47,In_2351,In_2277);
or U48 (N_48,In_663,In_1255);
and U49 (N_49,In_1439,In_2324);
xnor U50 (N_50,In_415,In_870);
nor U51 (N_51,In_1424,In_1604);
xor U52 (N_52,In_365,In_71);
nor U53 (N_53,In_295,In_319);
or U54 (N_54,In_1263,In_2357);
or U55 (N_55,In_497,In_1786);
nand U56 (N_56,In_1936,In_2732);
xnor U57 (N_57,In_1835,In_2239);
and U58 (N_58,In_2662,In_385);
and U59 (N_59,In_774,In_2344);
nor U60 (N_60,In_2446,In_1825);
nand U61 (N_61,In_2268,In_2924);
or U62 (N_62,In_955,In_69);
xnor U63 (N_63,In_2720,In_1071);
or U64 (N_64,In_1007,In_1614);
xnor U65 (N_65,In_2619,In_1711);
xor U66 (N_66,In_2273,In_456);
nor U67 (N_67,In_1091,In_2472);
or U68 (N_68,In_380,In_1098);
nor U69 (N_69,In_1262,In_2553);
nor U70 (N_70,In_707,In_438);
and U71 (N_71,In_2910,In_2917);
and U72 (N_72,In_95,In_2745);
nor U73 (N_73,In_644,In_2455);
xnor U74 (N_74,In_698,In_1659);
and U75 (N_75,In_2396,In_2219);
xor U76 (N_76,In_1598,In_1726);
nor U77 (N_77,In_2404,In_820);
xor U78 (N_78,In_2987,In_1183);
nor U79 (N_79,In_2633,In_1904);
or U80 (N_80,In_938,In_1710);
nand U81 (N_81,In_2321,In_660);
and U82 (N_82,In_514,In_1402);
or U83 (N_83,In_2083,In_2729);
xor U84 (N_84,In_788,In_374);
nand U85 (N_85,In_572,In_1385);
xor U86 (N_86,In_722,In_690);
xnor U87 (N_87,In_1586,In_25);
nand U88 (N_88,In_1952,In_1221);
nand U89 (N_89,In_185,In_1663);
nand U90 (N_90,In_162,In_123);
nand U91 (N_91,In_895,In_510);
or U92 (N_92,In_410,In_404);
nand U93 (N_93,In_1693,In_742);
or U94 (N_94,In_2886,In_57);
or U95 (N_95,In_2018,In_837);
xor U96 (N_96,In_1957,In_2356);
xnor U97 (N_97,In_2421,In_2862);
xnor U98 (N_98,In_135,In_2054);
or U99 (N_99,In_695,In_1188);
nor U100 (N_100,In_454,In_2806);
nor U101 (N_101,In_2780,In_149);
xor U102 (N_102,In_1486,In_763);
or U103 (N_103,In_1466,In_1430);
or U104 (N_104,In_1184,In_1353);
and U105 (N_105,In_2889,In_2123);
nor U106 (N_106,In_817,In_2919);
nor U107 (N_107,In_2042,In_1228);
xor U108 (N_108,In_2907,In_203);
or U109 (N_109,In_964,In_2163);
nand U110 (N_110,In_1802,In_1414);
nor U111 (N_111,In_948,In_592);
or U112 (N_112,In_2080,In_2270);
or U113 (N_113,In_1016,In_2021);
xor U114 (N_114,In_2640,In_1053);
nor U115 (N_115,In_1133,In_2452);
nand U116 (N_116,In_360,In_1761);
xnor U117 (N_117,In_2703,In_388);
and U118 (N_118,In_1943,In_2781);
nor U119 (N_119,In_1312,In_2686);
nand U120 (N_120,In_2069,In_897);
nand U121 (N_121,In_708,In_2705);
nand U122 (N_122,In_737,In_1516);
nand U123 (N_123,In_2736,In_19);
and U124 (N_124,In_248,In_1167);
or U125 (N_125,In_1288,In_2503);
and U126 (N_126,In_810,In_2861);
and U127 (N_127,In_1622,In_848);
nand U128 (N_128,In_2192,In_2989);
or U129 (N_129,In_428,In_1840);
and U130 (N_130,In_1771,In_1784);
and U131 (N_131,In_2485,In_1941);
nand U132 (N_132,In_831,In_2601);
xor U133 (N_133,In_2460,In_596);
nor U134 (N_134,In_1956,In_315);
nor U135 (N_135,In_1028,In_367);
nand U136 (N_136,In_1005,In_2487);
nor U137 (N_137,In_198,In_1477);
or U138 (N_138,In_2464,In_1880);
and U139 (N_139,In_1820,In_1314);
xor U140 (N_140,In_2994,In_1011);
xor U141 (N_141,In_842,In_1719);
and U142 (N_142,In_92,In_1803);
xnor U143 (N_143,In_2272,In_102);
and U144 (N_144,In_449,In_1589);
and U145 (N_145,In_987,In_1045);
xnor U146 (N_146,In_1155,In_1605);
nor U147 (N_147,In_614,In_1310);
and U148 (N_148,In_72,In_1476);
nand U149 (N_149,In_1980,In_1550);
nor U150 (N_150,In_2644,In_642);
or U151 (N_151,In_2873,In_2355);
nand U152 (N_152,In_1753,In_2880);
or U153 (N_153,In_2349,In_2738);
xor U154 (N_154,In_140,In_2721);
or U155 (N_155,In_390,In_53);
nand U156 (N_156,In_392,In_2865);
xnor U157 (N_157,In_2658,In_224);
nor U158 (N_158,In_652,In_1756);
nand U159 (N_159,In_1082,In_2588);
nand U160 (N_160,In_2326,In_1089);
nand U161 (N_161,In_62,In_1357);
xnor U162 (N_162,In_1688,In_2055);
or U163 (N_163,In_2758,In_2819);
and U164 (N_164,In_1842,In_1282);
or U165 (N_165,In_594,In_631);
and U166 (N_166,In_2832,In_2342);
nand U167 (N_167,In_2554,In_227);
or U168 (N_168,In_951,In_1940);
xor U169 (N_169,In_1576,In_2584);
xnor U170 (N_170,In_2656,In_2169);
or U171 (N_171,In_662,In_2657);
or U172 (N_172,In_38,In_1638);
or U173 (N_173,In_762,In_2578);
nand U174 (N_174,In_1555,In_575);
and U175 (N_175,In_362,In_1390);
and U176 (N_176,In_1884,In_734);
or U177 (N_177,In_2231,In_1853);
nand U178 (N_178,In_2453,In_2391);
nand U179 (N_179,In_233,In_1408);
or U180 (N_180,In_509,In_2100);
nor U181 (N_181,In_2835,In_2791);
nor U182 (N_182,In_2848,In_1295);
or U183 (N_183,In_2950,In_473);
nand U184 (N_184,In_1066,In_1539);
nand U185 (N_185,In_245,In_1524);
nor U186 (N_186,In_1100,In_582);
xor U187 (N_187,In_2111,In_1325);
nand U188 (N_188,In_1656,In_214);
or U189 (N_189,In_996,In_241);
nor U190 (N_190,In_1149,In_1725);
nor U191 (N_191,In_923,In_267);
or U192 (N_192,In_587,In_440);
nand U193 (N_193,In_451,In_1800);
nor U194 (N_194,In_2847,In_1674);
nor U195 (N_195,In_1728,In_2969);
nand U196 (N_196,In_780,In_1602);
xor U197 (N_197,In_376,In_1739);
xor U198 (N_198,In_2067,In_2401);
nor U199 (N_199,In_2682,In_2918);
nor U200 (N_200,In_610,In_1685);
and U201 (N_201,In_1925,In_158);
xnor U202 (N_202,In_1902,In_787);
nand U203 (N_203,In_2577,In_1404);
nand U204 (N_204,In_2755,In_798);
and U205 (N_205,In_2084,In_1501);
nand U206 (N_206,In_1552,In_975);
or U207 (N_207,In_1698,In_2434);
nand U208 (N_208,In_670,In_2432);
nand U209 (N_209,In_2618,In_931);
or U210 (N_210,In_1488,In_1933);
and U211 (N_211,In_2540,In_234);
and U212 (N_212,In_1345,In_1384);
and U213 (N_213,In_1206,In_993);
nor U214 (N_214,In_257,In_1497);
xor U215 (N_215,In_2766,In_579);
nor U216 (N_216,In_1680,In_2032);
nand U217 (N_217,In_395,In_1316);
nor U218 (N_218,In_768,In_2844);
and U219 (N_219,In_1966,In_398);
nand U220 (N_220,In_1067,In_998);
and U221 (N_221,In_34,In_301);
xor U222 (N_222,In_2768,In_1244);
xnor U223 (N_223,In_2591,In_2264);
nand U224 (N_224,In_1117,In_1724);
xor U225 (N_225,In_676,In_2991);
and U226 (N_226,In_2742,In_2428);
nand U227 (N_227,In_2778,In_2127);
xor U228 (N_228,In_283,In_2827);
xor U229 (N_229,In_2648,In_1442);
or U230 (N_230,In_2375,In_1762);
and U231 (N_231,In_1352,In_58);
xnor U232 (N_232,In_2267,In_2757);
xor U233 (N_233,In_402,In_2626);
and U234 (N_234,In_985,In_699);
or U235 (N_235,In_103,In_944);
nand U236 (N_236,In_2541,In_1290);
or U237 (N_237,In_1116,In_2805);
nor U238 (N_238,In_389,In_1759);
or U239 (N_239,In_1746,In_2348);
nor U240 (N_240,In_2718,In_814);
or U241 (N_241,In_2345,In_661);
xor U242 (N_242,In_546,In_99);
xnor U243 (N_243,In_2395,In_523);
and U244 (N_244,In_2585,In_442);
and U245 (N_245,In_694,In_1745);
or U246 (N_246,In_683,In_1729);
and U247 (N_247,In_1618,In_2869);
xnor U248 (N_248,In_1349,In_1839);
nor U249 (N_249,In_119,In_1174);
nand U250 (N_250,In_2872,In_1348);
nand U251 (N_251,In_2966,In_1964);
and U252 (N_252,In_521,In_1881);
nand U253 (N_253,In_1858,In_2816);
nand U254 (N_254,In_720,In_323);
and U255 (N_255,In_2689,In_351);
or U256 (N_256,In_1766,In_1062);
nand U257 (N_257,In_356,In_2539);
nor U258 (N_258,In_108,In_2458);
nand U259 (N_259,In_2437,In_217);
or U260 (N_260,In_835,In_2088);
xnor U261 (N_261,In_1138,In_87);
xnor U262 (N_262,In_2676,In_531);
or U263 (N_263,In_960,In_2614);
or U264 (N_264,In_2826,In_636);
and U265 (N_265,In_2990,In_256);
nor U266 (N_266,In_1838,In_142);
nand U267 (N_267,In_2660,In_483);
xnor U268 (N_268,In_1976,In_335);
nor U269 (N_269,In_1675,In_2311);
or U270 (N_270,In_1854,In_375);
or U271 (N_271,In_1626,In_423);
and U272 (N_272,In_1096,In_1879);
nand U273 (N_273,In_1735,In_2363);
and U274 (N_274,In_89,In_2140);
nor U275 (N_275,In_1392,In_1456);
or U276 (N_276,In_548,In_254);
and U277 (N_277,In_2794,In_43);
and U278 (N_278,In_1742,In_2062);
and U279 (N_279,In_173,In_1585);
xnor U280 (N_280,In_2424,In_1483);
or U281 (N_281,In_745,In_526);
nor U282 (N_282,In_45,In_51);
or U283 (N_283,In_1261,In_2975);
xor U284 (N_284,In_2152,In_1246);
xor U285 (N_285,In_1387,In_2125);
xnor U286 (N_286,In_859,In_2668);
xor U287 (N_287,In_1448,In_1421);
and U288 (N_288,In_2217,In_1632);
or U289 (N_289,In_1051,In_1105);
nand U290 (N_290,In_2531,In_2024);
nor U291 (N_291,In_2714,In_779);
and U292 (N_292,In_1446,In_2493);
xor U293 (N_293,In_247,In_1526);
nor U294 (N_294,In_2229,In_1667);
and U295 (N_295,In_2513,In_131);
or U296 (N_296,In_2678,In_2769);
nand U297 (N_297,In_175,In_1621);
and U298 (N_298,In_718,In_1977);
or U299 (N_299,In_2572,In_566);
xnor U300 (N_300,In_2912,In_1205);
xor U301 (N_301,In_105,In_2764);
and U302 (N_302,In_12,In_66);
xor U303 (N_303,In_28,In_971);
or U304 (N_304,In_1641,In_1300);
or U305 (N_305,In_252,In_1415);
xor U306 (N_306,In_2606,In_2936);
or U307 (N_307,In_891,In_2761);
and U308 (N_308,In_50,In_263);
nand U309 (N_309,In_528,In_1715);
or U310 (N_310,In_129,In_1059);
nor U311 (N_311,In_188,In_876);
or U312 (N_312,In_1308,In_2571);
xor U313 (N_313,In_11,In_2596);
or U314 (N_314,In_2358,In_1048);
xnor U315 (N_315,In_2305,In_840);
nand U316 (N_316,In_2979,In_1106);
or U317 (N_317,In_2426,In_1189);
and U318 (N_318,In_1620,In_2120);
and U319 (N_319,In_597,In_1723);
nor U320 (N_320,In_1033,In_2174);
nor U321 (N_321,In_168,In_327);
and U322 (N_322,In_834,In_802);
xor U323 (N_323,In_1574,In_1831);
xnor U324 (N_324,In_1423,In_2535);
nor U325 (N_325,In_761,In_239);
nand U326 (N_326,In_264,In_2447);
xor U327 (N_327,In_2227,In_2599);
and U328 (N_328,In_1085,In_101);
or U329 (N_329,In_1642,In_682);
xor U330 (N_330,In_2688,In_2722);
or U331 (N_331,In_2313,In_1333);
nand U332 (N_332,In_30,In_669);
and U333 (N_333,In_2151,In_477);
xor U334 (N_334,In_2538,In_472);
or U335 (N_335,In_621,In_1939);
or U336 (N_336,In_10,In_532);
nor U337 (N_337,In_1773,In_1578);
xnor U338 (N_338,In_296,In_1145);
nand U339 (N_339,In_892,In_2477);
nor U340 (N_340,In_94,In_287);
nor U341 (N_341,In_2103,In_1027);
nand U342 (N_342,In_2028,In_2370);
and U343 (N_343,In_202,In_2293);
nor U344 (N_344,In_446,In_2759);
nor U345 (N_345,In_1917,In_736);
or U346 (N_346,In_1363,In_2840);
xor U347 (N_347,In_6,In_2507);
nor U348 (N_348,In_9,In_700);
and U349 (N_349,In_703,In_867);
xnor U350 (N_350,In_1379,In_2050);
and U351 (N_351,In_1700,In_950);
nand U352 (N_352,In_2863,In_41);
nand U353 (N_353,In_384,In_2779);
xnor U354 (N_354,In_1457,In_1407);
nand U355 (N_355,In_222,In_693);
xnor U356 (N_356,In_2383,In_1485);
nand U357 (N_357,In_2394,In_641);
nand U358 (N_358,In_275,In_489);
xnor U359 (N_359,In_2871,In_591);
and U360 (N_360,In_2854,In_986);
nand U361 (N_361,In_2518,In_167);
nand U362 (N_362,In_1861,In_2203);
xnor U363 (N_363,In_2929,In_1744);
xnor U364 (N_364,In_941,In_265);
nand U365 (N_365,In_416,In_1912);
nand U366 (N_366,In_1903,In_2725);
and U367 (N_367,In_1613,In_2998);
or U368 (N_368,In_453,In_2124);
and U369 (N_369,In_2684,In_618);
xnor U370 (N_370,In_1367,In_1592);
nand U371 (N_371,In_2033,In_1788);
nor U372 (N_372,In_1703,In_1808);
and U373 (N_373,In_545,In_2726);
and U374 (N_374,In_434,In_2712);
nand U375 (N_375,In_1818,In_1266);
and U376 (N_376,In_1230,In_1185);
and U377 (N_377,In_2860,In_1533);
or U378 (N_378,In_866,In_620);
nand U379 (N_379,In_1630,In_349);
nor U380 (N_380,In_113,In_1326);
and U381 (N_381,In_2488,In_1169);
or U382 (N_382,In_2536,In_2971);
nand U383 (N_383,In_1410,In_795);
or U384 (N_384,In_529,In_2956);
nor U385 (N_385,In_1,In_1389);
xor U386 (N_386,In_1990,In_148);
nor U387 (N_387,In_485,In_1609);
xor U388 (N_388,In_1697,In_432);
nor U389 (N_389,In_2182,In_1572);
xnor U390 (N_390,In_2548,In_2636);
xnor U391 (N_391,In_554,In_231);
nor U392 (N_392,In_1296,In_2948);
or U393 (N_393,In_789,In_794);
nor U394 (N_394,In_2234,In_2456);
nand U395 (N_395,In_2749,In_291);
and U396 (N_396,In_139,In_611);
nor U397 (N_397,In_2164,In_1900);
or U398 (N_398,In_2312,In_1458);
xor U399 (N_399,In_1021,In_2592);
nand U400 (N_400,In_2261,In_2091);
and U401 (N_401,In_2200,In_1770);
and U402 (N_402,In_2193,In_2795);
or U403 (N_403,In_1420,In_7);
nand U404 (N_404,In_1931,In_486);
or U405 (N_405,In_862,In_1358);
nand U406 (N_406,In_1231,In_875);
nor U407 (N_407,In_1264,In_300);
or U408 (N_408,In_2798,In_1660);
and U409 (N_409,In_1567,In_2337);
nand U410 (N_410,In_1170,In_178);
xor U411 (N_411,In_2559,In_612);
nor U412 (N_412,In_1401,In_967);
nor U413 (N_413,In_674,In_1961);
nor U414 (N_414,In_154,In_1809);
nand U415 (N_415,In_2038,In_901);
xnor U416 (N_416,In_2409,In_2566);
nand U417 (N_417,In_2122,In_2499);
xnor U418 (N_418,In_1052,In_2988);
nor U419 (N_419,In_276,In_1346);
nand U420 (N_420,In_826,In_1676);
nand U421 (N_421,In_2800,In_1544);
nand U422 (N_422,In_1671,In_2951);
nand U423 (N_423,In_1055,In_1472);
xor U424 (N_424,In_2006,In_973);
xor U425 (N_425,In_1019,In_746);
nor U426 (N_426,In_633,In_161);
xor U427 (N_427,In_0,In_2010);
nor U428 (N_428,In_1259,In_2244);
and U429 (N_429,In_1751,In_598);
xor U430 (N_430,In_1543,In_2222);
xor U431 (N_431,In_2824,In_2374);
nand U432 (N_432,In_2365,In_1225);
xnor U433 (N_433,In_1899,In_1210);
and U434 (N_434,In_60,In_2465);
nor U435 (N_435,In_2065,In_1851);
or U436 (N_436,In_2281,In_2237);
or U437 (N_437,In_854,In_2802);
or U438 (N_438,In_2292,In_1874);
nor U439 (N_439,In_2878,In_2590);
nor U440 (N_440,In_304,In_2014);
nor U441 (N_441,In_286,In_1426);
and U442 (N_442,In_2296,In_1435);
or U443 (N_443,In_2341,In_2307);
xnor U444 (N_444,In_1923,In_339);
and U445 (N_445,In_1650,In_520);
nor U446 (N_446,In_2224,In_1548);
nor U447 (N_447,In_1168,In_2699);
nor U448 (N_448,In_1252,In_2467);
nand U449 (N_449,In_1554,In_1972);
or U450 (N_450,In_1627,In_1148);
or U451 (N_451,In_2254,In_580);
or U452 (N_452,In_2271,In_297);
and U453 (N_453,In_1565,In_1294);
or U454 (N_454,In_83,In_492);
and U455 (N_455,In_916,In_1954);
or U456 (N_456,In_864,In_1720);
and U457 (N_457,In_2378,In_371);
xnor U458 (N_458,In_536,In_617);
nand U459 (N_459,In_583,In_2524);
or U460 (N_460,In_56,In_136);
and U461 (N_461,In_49,In_86);
nor U462 (N_462,In_147,In_2072);
and U463 (N_463,In_1505,In_1517);
nor U464 (N_464,In_2459,In_1651);
nand U465 (N_465,In_885,In_2146);
xnor U466 (N_466,In_1304,In_2997);
nor U467 (N_467,In_650,In_2765);
nor U468 (N_468,In_1672,In_2955);
xor U469 (N_469,In_2533,In_731);
nor U470 (N_470,In_1635,In_1783);
or U471 (N_471,In_2753,In_459);
nand U472 (N_472,In_2331,In_2439);
or U473 (N_473,In_90,In_2719);
nand U474 (N_474,In_553,In_689);
and U475 (N_475,In_100,In_1232);
nand U476 (N_476,In_1186,In_461);
and U477 (N_477,In_715,In_2973);
nand U478 (N_478,In_898,In_1372);
or U479 (N_479,In_420,In_1559);
or U480 (N_480,In_2744,In_2444);
nand U481 (N_481,In_1000,In_1750);
nand U482 (N_482,In_1530,In_872);
and U483 (N_483,In_1437,In_204);
and U484 (N_484,In_293,In_1918);
xnor U485 (N_485,In_116,In_1837);
and U486 (N_486,In_749,In_220);
xnor U487 (N_487,In_1580,In_2534);
nor U488 (N_488,In_455,In_1193);
nor U489 (N_489,In_226,In_2046);
and U490 (N_490,In_1286,In_366);
nor U491 (N_491,In_2667,In_2519);
xnor U492 (N_492,In_500,In_1342);
xor U493 (N_493,In_1141,In_2977);
or U494 (N_494,In_2515,In_1950);
xnor U495 (N_495,In_2334,In_2265);
and U496 (N_496,In_2905,In_236);
xnor U497 (N_497,In_2594,In_2457);
or U498 (N_498,In_2438,In_1041);
or U499 (N_499,In_751,In_2299);
nor U500 (N_500,In_482,In_2491);
xor U501 (N_501,In_2801,In_2500);
and U502 (N_502,In_2278,In_357);
and U503 (N_503,In_2788,In_574);
nand U504 (N_504,In_851,In_855);
and U505 (N_505,In_1238,In_1425);
nor U506 (N_506,In_2256,In_31);
and U507 (N_507,In_1191,In_2213);
and U508 (N_508,In_608,In_180);
and U509 (N_509,In_13,In_1562);
or U510 (N_510,In_112,In_691);
and U511 (N_511,In_2450,In_1558);
and U512 (N_512,In_2484,In_2115);
and U513 (N_513,In_284,In_905);
or U514 (N_514,In_1937,In_2389);
nor U515 (N_515,In_2544,In_1391);
xor U516 (N_516,In_251,In_1927);
xnor U517 (N_517,In_1269,In_1134);
nand U518 (N_518,In_1330,In_1568);
xnor U519 (N_519,In_1004,In_1577);
nor U520 (N_520,In_1097,In_818);
and U521 (N_521,In_2413,In_664);
or U522 (N_522,In_668,In_1633);
nor U523 (N_523,In_1160,In_2909);
nand U524 (N_524,In_64,In_1699);
xnor U525 (N_525,In_2037,In_444);
or U526 (N_526,In_525,In_1668);
or U527 (N_527,In_1107,In_1684);
and U528 (N_528,In_671,In_2157);
and U529 (N_529,In_2760,In_1867);
and U530 (N_530,In_2690,In_277);
and U531 (N_531,In_1465,In_2492);
nor U532 (N_532,In_109,In_2167);
and U533 (N_533,In_2627,In_1515);
or U534 (N_534,In_1844,In_1212);
nor U535 (N_535,In_706,In_2246);
xnor U536 (N_536,In_150,In_839);
nand U537 (N_537,In_2144,In_67);
xor U538 (N_538,In_2258,In_606);
nor U539 (N_539,In_1126,In_2509);
nand U540 (N_540,In_273,In_823);
xor U541 (N_541,In_2945,In_2251);
nand U542 (N_542,In_1382,In_2853);
nand U543 (N_543,In_607,In_2992);
nand U544 (N_544,In_1712,In_2552);
nor U545 (N_545,In_2646,In_2443);
and U546 (N_546,In_2922,In_121);
xor U547 (N_547,In_2332,In_408);
xor U548 (N_548,In_1022,In_2023);
or U549 (N_549,In_915,In_1359);
and U550 (N_550,In_1776,In_318);
xor U551 (N_551,In_1988,In_2173);
nand U552 (N_552,In_551,In_2250);
or U553 (N_553,In_796,In_1427);
nor U554 (N_554,In_513,In_2575);
or U555 (N_555,In_2215,In_1508);
xnor U556 (N_556,In_1780,In_448);
xnor U557 (N_557,In_752,In_2665);
and U558 (N_558,In_781,In_1157);
nand U559 (N_559,In_1090,In_2784);
and U560 (N_560,In_1194,In_21);
or U561 (N_561,In_1519,In_2223);
nand U562 (N_562,In_666,In_1587);
or U563 (N_563,In_2856,In_2821);
xor U564 (N_564,In_1969,In_1953);
and U565 (N_565,In_2454,In_2762);
nor U566 (N_566,In_2527,In_760);
nand U567 (N_567,In_2284,In_1795);
xnor U568 (N_568,In_2191,In_902);
xnor U569 (N_569,In_1755,In_2498);
xor U570 (N_570,In_1332,In_1491);
nor U571 (N_571,In_2388,In_2304);
nor U572 (N_572,In_2117,In_1540);
nor U573 (N_573,In_2053,In_2479);
and U574 (N_574,In_2399,In_55);
nand U575 (N_575,In_115,In_98);
and U576 (N_576,In_1997,In_2036);
or U577 (N_577,In_2846,In_2266);
or U578 (N_578,In_1075,In_1566);
nor U579 (N_579,In_1637,In_1002);
xor U580 (N_580,In_1434,In_649);
nor U581 (N_581,In_330,In_2445);
and U582 (N_582,In_1118,In_238);
and U583 (N_583,In_399,In_462);
nand U584 (N_584,In_2198,In_2177);
nor U585 (N_585,In_2700,In_894);
or U586 (N_586,In_174,In_383);
xnor U587 (N_587,In_2804,In_888);
and U588 (N_588,In_2078,In_2851);
xor U589 (N_589,In_1876,In_1769);
nand U590 (N_590,In_1624,In_1905);
nand U591 (N_591,In_2184,In_712);
nor U592 (N_592,In_963,In_1845);
nand U593 (N_593,In_1871,In_1509);
or U594 (N_594,In_160,In_2419);
xnor U595 (N_595,In_2210,In_1691);
and U596 (N_596,In_1653,In_2661);
and U597 (N_597,In_2005,In_2262);
or U598 (N_598,In_2077,In_2563);
or U599 (N_599,In_1073,In_1570);
and U600 (N_600,In_2674,In_1805);
and U601 (N_601,In_1500,In_305);
or U602 (N_602,In_1599,In_2775);
and U603 (N_603,In_1843,In_1086);
nand U604 (N_604,In_341,In_1920);
nor U605 (N_605,In_2063,In_2397);
nor U606 (N_606,In_2451,In_1317);
nor U607 (N_607,In_68,In_1049);
nand U608 (N_608,In_2407,In_733);
and U609 (N_609,In_2654,In_679);
nand U610 (N_610,In_84,In_1452);
or U611 (N_611,In_1657,In_1275);
nor U612 (N_612,In_1137,In_2695);
or U613 (N_613,In_1087,In_2114);
xor U614 (N_614,In_637,In_1738);
or U615 (N_615,In_2135,In_1865);
nand U616 (N_616,In_4,In_983);
and U617 (N_617,In_565,In_1794);
nor U618 (N_618,In_2132,In_1419);
or U619 (N_619,In_1971,In_2603);
nor U620 (N_620,In_705,In_588);
xnor U621 (N_621,In_2473,In_1181);
xnor U622 (N_622,In_1202,In_995);
and U623 (N_623,In_1730,In_2449);
or U624 (N_624,In_1076,In_2743);
and U625 (N_625,In_2842,In_1666);
xor U626 (N_626,In_1763,In_1373);
nand U627 (N_627,In_2208,In_336);
nor U628 (N_628,In_2166,In_2435);
and U629 (N_629,In_1084,In_2952);
or U630 (N_630,In_2330,In_1257);
nand U631 (N_631,In_2073,In_1528);
xor U632 (N_632,In_2980,In_1192);
nand U633 (N_633,In_278,In_704);
xnor U634 (N_634,In_726,In_982);
nor U635 (N_635,In_1271,In_2070);
and U636 (N_636,In_2625,In_393);
nor U637 (N_637,In_2583,In_1433);
nor U638 (N_638,In_2673,In_39);
and U639 (N_639,In_1152,In_54);
or U640 (N_640,In_1161,In_907);
and U641 (N_641,In_804,In_564);
and U642 (N_642,In_2579,In_2859);
xnor U643 (N_643,In_1224,In_1686);
or U644 (N_644,In_710,In_1339);
nor U645 (N_645,In_558,In_1147);
nand U646 (N_646,In_2734,In_2694);
or U647 (N_647,In_179,In_1878);
and U648 (N_648,In_1721,In_1409);
nand U649 (N_649,In_2346,In_2221);
xor U650 (N_650,In_2843,In_2663);
or U651 (N_651,In_1462,In_2338);
nand U652 (N_652,In_966,In_2620);
or U653 (N_653,In_2303,In_2172);
xor U654 (N_654,In_1764,In_1872);
nand U655 (N_655,In_845,In_1896);
or U656 (N_656,In_246,In_2171);
nor U657 (N_657,In_1661,In_499);
xnor U658 (N_658,In_2422,In_1222);
nor U659 (N_659,In_2000,In_2380);
xor U660 (N_660,In_2876,In_1982);
and U661 (N_661,In_1983,In_2106);
and U662 (N_662,In_1495,In_2286);
nand U663 (N_663,In_1281,In_811);
xnor U664 (N_664,In_1108,In_945);
nor U665 (N_665,In_126,In_882);
and U666 (N_666,In_1777,In_2677);
nand U667 (N_667,In_2890,In_1234);
nor U668 (N_668,In_2022,In_2186);
nor U669 (N_669,In_1461,In_1305);
xor U670 (N_670,In_927,In_877);
xnor U671 (N_671,In_271,In_2982);
and U672 (N_672,In_76,In_1819);
xor U673 (N_673,In_1612,In_2112);
nand U674 (N_674,In_904,In_460);
nand U675 (N_675,In_437,In_208);
and U676 (N_676,In_1199,In_166);
or U677 (N_677,In_1381,In_1834);
or U678 (N_678,In_346,In_524);
nand U679 (N_679,In_1219,In_1591);
nand U680 (N_680,In_1717,In_1468);
nor U681 (N_681,In_1877,In_1413);
or U682 (N_682,In_1386,In_329);
xor U683 (N_683,In_2683,In_1890);
and U684 (N_684,In_1179,In_141);
xnor U685 (N_685,In_2562,In_1113);
xnor U686 (N_686,In_378,In_2225);
or U687 (N_687,In_425,In_2252);
and U688 (N_688,In_469,In_1215);
and U689 (N_689,In_1362,In_1006);
or U690 (N_690,In_2108,In_1365);
and U691 (N_691,In_793,In_2328);
nor U692 (N_692,In_1573,In_195);
nor U693 (N_693,In_1506,In_1600);
and U694 (N_694,In_658,In_2373);
xor U695 (N_695,In_871,In_601);
xnor U696 (N_696,In_2894,In_1647);
xnor U697 (N_697,In_869,In_559);
and U698 (N_698,In_1343,In_2480);
nor U699 (N_699,In_186,In_1277);
or U700 (N_700,In_2589,In_3);
or U701 (N_701,In_2642,In_2561);
nand U702 (N_702,In_1998,In_2336);
nor U703 (N_703,In_673,In_427);
and U704 (N_704,In_576,In_2368);
nand U705 (N_705,In_934,In_2274);
nand U706 (N_706,In_1187,In_2938);
nor U707 (N_707,In_2961,In_1492);
or U708 (N_708,In_2698,In_1388);
nand U709 (N_709,In_2605,In_2384);
and U710 (N_710,In_343,In_1046);
nand U711 (N_711,In_1512,In_2);
xnor U712 (N_712,In_2367,In_303);
xnor U713 (N_713,In_1397,In_1180);
and U714 (N_714,In_1243,In_316);
xnor U715 (N_715,In_1038,In_822);
xor U716 (N_716,In_2099,In_2162);
xor U717 (N_717,In_2771,In_1454);
and U718 (N_718,In_1560,In_1124);
xnor U719 (N_719,In_1814,In_1993);
xor U720 (N_720,In_2130,In_1163);
or U721 (N_721,In_2302,In_1173);
nand U722 (N_722,In_604,In_860);
and U723 (N_723,In_1584,In_2850);
xnor U724 (N_724,In_2020,In_171);
and U725 (N_725,In_250,In_2786);
and U726 (N_726,In_441,In_2400);
nand U727 (N_727,In_2474,In_1687);
and U728 (N_728,In_2685,In_480);
and U729 (N_729,In_2985,In_2483);
xor U730 (N_730,In_1396,In_2420);
nand U731 (N_731,In_1328,In_218);
nor U732 (N_732,In_600,In_1907);
xnor U733 (N_733,In_372,In_800);
or U734 (N_734,In_2034,In_1929);
or U735 (N_735,In_2041,In_1816);
nand U736 (N_736,In_18,In_2796);
and U737 (N_737,In_1223,In_2899);
nor U738 (N_738,In_1996,In_2838);
and U739 (N_739,In_1159,In_1144);
and U740 (N_740,In_2962,In_1088);
and U741 (N_741,In_1617,In_1035);
or U742 (N_742,In_556,In_1894);
nor U743 (N_743,In_189,In_1799);
or U744 (N_744,In_651,In_542);
or U745 (N_745,In_2650,In_1371);
and U746 (N_746,In_1429,In_37);
nor U747 (N_747,In_799,In_2094);
xor U748 (N_748,In_82,In_1321);
nand U749 (N_749,In_159,In_2188);
and U750 (N_750,In_2471,In_2604);
xor U751 (N_751,In_956,In_2406);
nor U752 (N_752,In_156,In_1121);
xnor U753 (N_753,In_2196,In_1658);
xor U754 (N_754,In_959,In_1025);
nor U755 (N_755,In_832,In_990);
and U756 (N_756,In_29,In_52);
nand U757 (N_757,In_2574,In_2290);
or U758 (N_758,In_2681,In_2891);
nand U759 (N_759,In_1449,In_2137);
nand U760 (N_760,In_502,In_1758);
nor U761 (N_761,In_1455,In_1399);
xnor U762 (N_762,In_2039,In_2008);
xnor U763 (N_763,In_386,In_1061);
nand U764 (N_764,In_1398,In_1986);
and U765 (N_765,In_2923,In_567);
xnor U766 (N_766,In_1796,In_1648);
or U767 (N_767,In_1708,In_1860);
nand U768 (N_768,In_2415,In_2481);
and U769 (N_769,In_2999,In_954);
nor U770 (N_770,In_96,In_2965);
or U771 (N_771,In_1253,In_1280);
xnor U772 (N_772,In_2582,In_2076);
xor U773 (N_773,In_2666,In_1475);
nor U774 (N_774,In_2153,In_957);
and U775 (N_775,In_170,In_2044);
and U776 (N_776,In_47,In_2505);
nand U777 (N_777,In_1833,In_917);
xor U778 (N_778,In_397,In_1012);
xor U779 (N_779,In_1852,In_2026);
or U780 (N_780,In_1115,In_874);
or U781 (N_781,In_2622,In_883);
or U782 (N_782,In_881,In_450);
xnor U783 (N_783,In_613,In_2052);
nor U784 (N_784,In_1298,In_240);
or U785 (N_785,In_1810,In_235);
nor U786 (N_786,In_757,In_2741);
and U787 (N_787,In_2611,In_2178);
and U788 (N_788,In_2361,In_439);
nand U789 (N_789,In_1018,In_413);
or U790 (N_790,In_2398,In_1636);
and U791 (N_791,In_2354,In_2968);
and U792 (N_792,In_324,In_2623);
nand U793 (N_793,In_602,In_2327);
nor U794 (N_794,In_646,In_1162);
nor U795 (N_795,In_1177,In_1518);
or U796 (N_796,In_581,In_2727);
nand U797 (N_797,In_1068,In_2340);
and U798 (N_798,In_1494,In_114);
or U799 (N_799,In_2081,In_772);
nor U800 (N_800,In_211,In_310);
xnor U801 (N_801,In_2697,In_541);
nand U802 (N_802,In_672,In_1132);
or U803 (N_803,In_2972,In_2830);
nand U804 (N_804,In_223,In_829);
xnor U805 (N_805,In_833,In_1251);
or U806 (N_806,In_1779,In_503);
xnor U807 (N_807,In_759,In_2911);
and U808 (N_808,In_110,In_727);
xor U809 (N_809,In_1276,In_1502);
nor U810 (N_810,In_2436,In_685);
and U811 (N_811,In_1122,In_258);
or U812 (N_812,In_230,In_738);
xor U813 (N_813,In_2953,In_2543);
nor U814 (N_814,In_2836,In_207);
and U815 (N_815,In_2248,In_2680);
nand U816 (N_816,In_2269,In_2609);
and U817 (N_817,In_1639,In_2820);
nor U818 (N_818,In_16,In_15);
xnor U819 (N_819,In_1054,In_2294);
nand U820 (N_820,In_1888,In_2933);
and U821 (N_821,In_282,In_79);
nand U822 (N_822,In_127,In_1696);
nor U823 (N_823,In_1610,In_302);
and U824 (N_824,In_1037,In_2110);
and U825 (N_825,In_1741,In_557);
nand U826 (N_826,In_73,In_1198);
and U827 (N_827,In_816,In_1376);
nand U828 (N_828,In_825,In_1503);
and U829 (N_829,In_2101,In_2525);
or U830 (N_830,In_2318,In_999);
and U831 (N_831,In_1704,In_93);
xor U832 (N_832,In_1313,In_1026);
or U833 (N_833,In_547,In_2385);
nor U834 (N_834,In_2206,In_299);
and U835 (N_835,In_430,In_2560);
xnor U836 (N_836,In_2118,In_1023);
and U837 (N_837,In_2870,In_643);
nand U838 (N_838,In_2285,In_1125);
xnor U839 (N_839,In_2275,In_2866);
nand U840 (N_840,In_379,In_382);
nand U841 (N_841,In_599,In_1947);
xor U842 (N_842,In_2353,In_192);
xnor U843 (N_843,In_2185,In_2932);
xor U844 (N_844,In_2003,In_1327);
and U845 (N_845,In_2071,In_2993);
nand U846 (N_846,In_1216,In_2212);
nor U847 (N_847,In_2119,In_1318);
and U848 (N_848,In_479,In_925);
nor U849 (N_849,In_619,In_464);
nor U850 (N_850,In_355,In_1942);
xor U851 (N_851,In_2226,In_2747);
xnor U852 (N_852,In_1237,In_1975);
nand U853 (N_853,In_426,In_2696);
or U854 (N_854,In_537,In_2064);
and U855 (N_855,In_792,In_1203);
nand U856 (N_856,In_194,In_122);
nand U857 (N_857,In_819,In_2194);
nand U858 (N_858,In_2298,In_595);
nand U859 (N_859,In_1864,In_2496);
nand U860 (N_860,In_2004,In_716);
nor U861 (N_861,In_471,In_2881);
xnor U862 (N_862,In_1070,In_585);
nand U863 (N_863,In_1099,In_632);
nor U864 (N_864,In_974,In_1496);
or U865 (N_865,In_2517,In_2187);
or U866 (N_866,In_2837,In_1959);
and U867 (N_867,In_2995,In_125);
xor U868 (N_868,In_298,In_1207);
or U869 (N_869,In_721,In_1767);
xor U870 (N_870,In_2511,In_132);
and U871 (N_871,In_2238,In_155);
xor U872 (N_872,In_221,In_2126);
nand U873 (N_873,In_1393,In_2797);
and U874 (N_874,In_1922,In_91);
and U875 (N_875,In_1889,In_2209);
nor U876 (N_876,In_2136,In_1970);
and U877 (N_877,In_2691,In_2621);
xor U878 (N_878,In_1140,In_2201);
xnor U879 (N_879,In_433,In_1247);
nor U880 (N_880,In_1875,In_1863);
nor U881 (N_881,In_70,In_778);
or U882 (N_882,In_713,In_1513);
xnor U883 (N_883,In_1722,In_2925);
xor U884 (N_884,In_1204,In_1406);
nand U885 (N_885,In_2082,In_2913);
nor U886 (N_886,In_1211,In_843);
and U887 (N_887,In_1438,In_1460);
nand U888 (N_888,In_2545,In_1102);
nor U889 (N_889,In_2339,In_527);
nand U890 (N_890,In_910,In_2532);
nand U891 (N_891,In_2839,In_2598);
nand U892 (N_892,In_830,In_1267);
nor U893 (N_893,In_1522,In_196);
or U894 (N_894,In_1058,In_1760);
and U895 (N_895,In_1866,In_656);
or U896 (N_896,In_228,In_177);
or U897 (N_897,In_1590,In_1553);
xor U898 (N_898,In_1171,In_2875);
nor U899 (N_899,In_2263,In_2109);
or U900 (N_900,In_812,In_1279);
nand U901 (N_901,In_2462,In_391);
nor U902 (N_902,In_1369,In_447);
or U903 (N_903,In_2568,In_2715);
nand U904 (N_904,In_2143,In_782);
and U905 (N_905,In_1095,In_1596);
xor U906 (N_906,In_624,In_1047);
nor U907 (N_907,In_1412,In_1527);
and U908 (N_908,In_684,In_868);
and U909 (N_909,In_1994,In_487);
xor U910 (N_910,In_255,In_1582);
and U911 (N_911,In_861,In_2904);
xnor U912 (N_912,In_1248,In_2074);
nor U913 (N_913,In_1153,In_36);
xnor U914 (N_914,In_755,In_1707);
or U915 (N_915,In_518,In_1702);
xor U916 (N_916,In_80,In_2205);
xnor U917 (N_917,In_281,In_949);
or U918 (N_918,In_2043,In_1445);
or U919 (N_919,In_1176,In_2031);
or U920 (N_920,In_2651,In_1938);
nand U921 (N_921,In_815,In_1351);
nor U922 (N_922,In_2523,In_2506);
and U923 (N_923,In_1921,In_1417);
xor U924 (N_924,In_765,In_2898);
or U925 (N_925,In_2692,In_1306);
xor U926 (N_926,In_2629,In_120);
and U927 (N_927,In_2895,In_2638);
or U928 (N_928,In_961,In_803);
xor U929 (N_929,In_1951,In_770);
xor U930 (N_930,In_2183,In_2770);
xnor U931 (N_931,In_2570,In_667);
nand U932 (N_932,In_616,In_306);
nor U933 (N_933,In_984,In_272);
nor U934 (N_934,In_827,In_1344);
nand U935 (N_935,In_786,In_400);
nor U936 (N_936,In_1114,In_2879);
and U937 (N_937,In_1538,In_981);
or U938 (N_938,In_2300,In_919);
nor U939 (N_939,In_143,In_2207);
nor U940 (N_940,In_2664,In_2659);
nand U941 (N_941,In_937,In_331);
or U942 (N_942,In_2597,In_1083);
or U943 (N_943,In_926,In_1713);
or U944 (N_944,In_725,In_797);
nand U945 (N_945,In_2016,In_506);
xnor U946 (N_946,In_776,In_61);
or U947 (N_947,In_165,In_1329);
nor U948 (N_948,In_630,In_1443);
xor U949 (N_949,In_654,In_732);
xnor U950 (N_950,In_1213,In_348);
nand U951 (N_951,In_2731,In_2649);
and U952 (N_952,In_2086,In_2075);
xor U953 (N_953,In_2983,In_2735);
and U954 (N_954,In_2740,In_2792);
or U955 (N_955,In_1649,In_85);
and U956 (N_956,In_290,In_1292);
nand U957 (N_957,In_2610,In_2236);
or U958 (N_958,In_1142,In_1556);
xnor U959 (N_959,In_146,In_2928);
and U960 (N_960,In_1010,In_436);
xnor U961 (N_961,In_289,In_1916);
or U962 (N_962,In_2061,In_2874);
and U963 (N_963,In_841,In_2259);
or U964 (N_964,In_2967,In_2138);
nand U965 (N_965,In_468,In_2670);
nand U966 (N_966,In_753,In_2814);
or U967 (N_967,In_20,In_1064);
xnor U968 (N_968,In_1209,In_187);
or U969 (N_969,In_107,In_63);
nand U970 (N_970,In_1042,In_422);
or U971 (N_971,In_1749,In_2372);
and U972 (N_972,In_1380,In_2701);
nand U973 (N_973,In_261,In_1790);
xor U974 (N_974,In_2165,In_976);
nand U975 (N_975,In_2808,In_74);
nor U976 (N_976,In_476,In_735);
nand U977 (N_977,In_1891,In_387);
nor U978 (N_978,In_863,In_2547);
nor U979 (N_979,In_229,In_190);
nand U980 (N_980,In_1727,In_2752);
nand U981 (N_981,In_1440,In_1849);
nand U982 (N_982,In_2011,In_687);
or U983 (N_983,In_2573,In_2569);
or U984 (N_984,In_2613,In_1337);
xor U985 (N_985,In_962,In_1734);
nand U986 (N_986,In_1806,In_2974);
nand U987 (N_987,In_952,In_1201);
and U988 (N_988,In_2371,In_2405);
nand U989 (N_989,In_979,In_2092);
and U990 (N_990,In_2335,In_322);
or U991 (N_991,In_2807,In_909);
nor U992 (N_992,In_1249,In_65);
nand U993 (N_993,In_342,In_1895);
nand U994 (N_994,In_1166,In_628);
or U995 (N_995,In_1341,In_2204);
or U996 (N_996,In_1254,In_2494);
and U997 (N_997,In_2617,In_1525);
or U998 (N_998,In_2679,In_543);
xnor U999 (N_999,In_2325,In_723);
and U1000 (N_1000,In_1069,In_163);
xnor U1001 (N_1001,In_1214,In_2637);
or U1002 (N_1002,In_1057,In_1705);
xor U1003 (N_1003,In_1594,In_1689);
nor U1004 (N_1004,In_1017,In_2220);
or U1005 (N_1005,In_1932,In_2903);
and U1006 (N_1006,In_573,In_2448);
xor U1007 (N_1007,In_2416,In_2602);
nor U1008 (N_1008,In_1473,In_1074);
or U1009 (N_1009,In_692,In_517);
nand U1010 (N_1010,In_1274,In_1120);
xor U1011 (N_1011,In_791,In_1374);
nor U1012 (N_1012,In_1625,In_1507);
nor U1013 (N_1013,In_1930,In_1030);
nor U1014 (N_1014,In_2555,In_714);
nand U1015 (N_1015,In_2653,In_1182);
nand U1016 (N_1016,In_920,In_1774);
nand U1017 (N_1017,In_1985,In_2476);
nand U1018 (N_1018,In_2809,In_2934);
xor U1019 (N_1019,In_2366,In_2655);
and U1020 (N_1020,In_484,In_2049);
or U1021 (N_1021,In_2159,In_1909);
nand U1022 (N_1022,In_133,In_117);
or U1023 (N_1023,In_1463,In_615);
and U1024 (N_1024,In_199,In_151);
or U1025 (N_1025,In_665,In_2687);
xor U1026 (N_1026,In_2858,In_478);
nor U1027 (N_1027,In_1436,In_512);
or U1028 (N_1028,In_1615,In_2564);
nand U1029 (N_1029,In_2410,In_1239);
nor U1030 (N_1030,In_2986,In_2546);
nand U1031 (N_1031,In_1887,In_2964);
nor U1032 (N_1032,In_1178,In_181);
nor U1033 (N_1033,In_1471,In_27);
nand U1034 (N_1034,In_2295,In_908);
or U1035 (N_1035,In_1601,In_2772);
and U1036 (N_1036,In_590,In_2773);
nand U1037 (N_1037,In_2565,In_911);
and U1038 (N_1038,In_2035,In_394);
and U1039 (N_1039,In_2516,In_2461);
nand U1040 (N_1040,In_1459,In_539);
nand U1041 (N_1041,In_488,In_2645);
or U1042 (N_1042,In_740,In_1265);
and U1043 (N_1043,In_2628,In_1158);
xor U1044 (N_1044,In_994,In_405);
nand U1045 (N_1045,In_773,In_1934);
nor U1046 (N_1046,In_1606,In_2202);
nand U1047 (N_1047,In_739,In_138);
or U1048 (N_1048,In_78,In_879);
xor U1049 (N_1049,In_2333,In_1375);
or U1050 (N_1050,In_1801,In_1464);
nor U1051 (N_1051,In_1883,In_2669);
xor U1052 (N_1052,In_2803,In_516);
nor U1053 (N_1053,In_1112,In_340);
xor U1054 (N_1054,In_2142,In_369);
nand U1055 (N_1055,In_1646,In_1826);
and U1056 (N_1056,In_1856,In_2567);
or U1057 (N_1057,In_431,In_1043);
or U1058 (N_1058,In_2116,In_370);
or U1059 (N_1059,In_634,In_2711);
nor U1060 (N_1060,In_1289,In_2260);
xnor U1061 (N_1061,In_930,In_466);
nand U1062 (N_1062,In_307,In_2240);
or U1063 (N_1063,In_942,In_729);
nor U1064 (N_1064,In_2739,In_2093);
nor U1065 (N_1065,In_1489,In_1694);
and U1066 (N_1066,In_1164,In_1360);
nor U1067 (N_1067,In_2047,In_2892);
and U1068 (N_1068,In_77,In_184);
xor U1069 (N_1069,In_1273,In_2897);
xnor U1070 (N_1070,In_1682,In_2520);
and U1071 (N_1071,In_1060,In_2350);
nand U1072 (N_1072,In_2440,In_2377);
xor U1073 (N_1073,In_2782,In_2241);
nand U1074 (N_1074,In_2056,In_2530);
nor U1075 (N_1075,In_2643,In_1498);
nor U1076 (N_1076,In_893,In_530);
xor U1077 (N_1077,In_1817,In_1323);
and U1078 (N_1078,In_2301,In_1772);
nand U1079 (N_1079,In_213,In_172);
nor U1080 (N_1080,In_2381,In_128);
or U1081 (N_1081,In_562,In_1945);
or U1082 (N_1082,In_1383,In_2015);
nand U1083 (N_1083,In_1422,In_1283);
nand U1084 (N_1084,In_969,In_972);
or U1085 (N_1085,In_2382,In_2707);
nor U1086 (N_1086,In_1511,In_2408);
nor U1087 (N_1087,In_1901,In_627);
and U1088 (N_1088,In_1611,In_435);
or U1089 (N_1089,In_2831,In_134);
nor U1090 (N_1090,In_2002,In_182);
nor U1091 (N_1091,In_2510,In_640);
or U1092 (N_1092,In_577,In_1631);
or U1093 (N_1093,In_81,In_2417);
and U1094 (N_1094,In_2051,In_709);
and U1095 (N_1095,In_403,In_1989);
xnor U1096 (N_1096,In_2287,In_1015);
or U1097 (N_1097,In_2096,In_2133);
xnor U1098 (N_1098,In_2528,In_1451);
nand U1099 (N_1099,In_2001,In_452);
nand U1100 (N_1100,In_724,In_1299);
xnor U1101 (N_1101,In_197,In_1196);
and U1102 (N_1102,In_748,In_2013);
and U1103 (N_1103,In_1172,In_2218);
nor U1104 (N_1104,In_1886,In_2045);
or U1105 (N_1105,In_750,In_2068);
nor U1106 (N_1106,In_2121,In_853);
nand U1107 (N_1107,In_609,In_805);
xnor U1108 (N_1108,In_1319,In_743);
and U1109 (N_1109,In_2902,In_2105);
and U1110 (N_1110,In_2901,In_2789);
and U1111 (N_1111,In_807,In_2774);
or U1112 (N_1112,In_1241,In_2817);
nor U1113 (N_1113,In_1848,In_953);
or U1114 (N_1114,In_2139,In_2504);
nand U1115 (N_1115,In_1079,In_1474);
and U1116 (N_1116,In_766,In_1987);
or U1117 (N_1117,In_2433,In_1129);
nor U1118 (N_1118,In_1979,In_921);
and U1119 (N_1119,In_345,In_906);
nand U1120 (N_1120,In_635,In_1645);
and U1121 (N_1121,In_1354,In_2672);
nor U1122 (N_1122,In_880,In_2896);
and U1123 (N_1123,In_1250,In_1546);
xor U1124 (N_1124,In_1733,In_1765);
xnor U1125 (N_1125,In_2322,In_625);
and U1126 (N_1126,In_1418,In_1958);
and U1127 (N_1127,In_1768,In_42);
and U1128 (N_1128,In_549,In_317);
nor U1129 (N_1129,In_2825,In_1747);
nand U1130 (N_1130,In_645,In_1242);
xor U1131 (N_1131,In_2616,In_2529);
xor U1132 (N_1132,In_2040,In_767);
and U1133 (N_1133,In_2724,In_785);
xnor U1134 (N_1134,In_1478,In_2087);
and U1135 (N_1135,In_1670,In_2750);
xor U1136 (N_1136,In_570,In_2017);
nand U1137 (N_1137,In_1233,In_26);
xor U1138 (N_1138,In_1807,In_1830);
nand U1139 (N_1139,In_2019,In_2329);
and U1140 (N_1140,In_1870,In_2737);
nor U1141 (N_1141,In_1394,In_46);
nor U1142 (N_1142,In_2716,In_1775);
nand U1143 (N_1143,In_2463,In_1690);
or U1144 (N_1144,In_344,In_1240);
xor U1145 (N_1145,In_2748,In_1999);
xnor U1146 (N_1146,In_474,In_1563);
xnor U1147 (N_1147,In_2702,In_2352);
or U1148 (N_1148,In_2403,In_1995);
nor U1149 (N_1149,In_1128,In_1285);
xor U1150 (N_1150,In_992,In_1123);
or U1151 (N_1151,In_200,In_1103);
or U1152 (N_1152,In_1403,In_1811);
and U1153 (N_1153,In_2671,In_1195);
xnor U1154 (N_1154,In_481,In_2442);
and U1155 (N_1155,In_1301,In_771);
xnor U1156 (N_1156,In_421,In_1411);
and U1157 (N_1157,In_104,In_2392);
or U1158 (N_1158,In_2887,In_8);
nor U1159 (N_1159,In_1297,In_118);
or U1160 (N_1160,In_2427,In_1284);
nand U1161 (N_1161,In_1960,In_2309);
nor U1162 (N_1162,In_44,In_1356);
or U1163 (N_1163,In_946,In_2158);
or U1164 (N_1164,In_169,In_544);
or U1165 (N_1165,In_688,In_1322);
nor U1166 (N_1166,In_445,In_1859);
nor U1167 (N_1167,In_1479,In_1797);
and U1168 (N_1168,In_1469,In_2495);
nor U1169 (N_1169,In_678,In_913);
or U1170 (N_1170,In_1320,In_2190);
nand U1171 (N_1171,In_1718,In_2709);
or U1172 (N_1172,In_475,In_997);
xor U1173 (N_1173,In_933,In_1136);
nor U1174 (N_1174,In_1514,In_2822);
or U1175 (N_1175,In_2704,In_2257);
nor U1176 (N_1176,In_2155,In_1855);
xor U1177 (N_1177,In_1752,In_2468);
or U1178 (N_1178,In_2706,In_1962);
nor U1179 (N_1179,In_2027,In_1034);
nor U1180 (N_1180,In_2387,In_2970);
nand U1181 (N_1181,In_1220,In_1190);
or U1182 (N_1182,In_991,In_259);
or U1183 (N_1183,In_1662,In_965);
nand U1184 (N_1184,In_1824,In_1032);
nor U1185 (N_1185,In_2549,In_1673);
xnor U1186 (N_1186,In_157,In_2957);
and U1187 (N_1187,In_1991,In_2486);
nor U1188 (N_1188,In_2841,In_2113);
or U1189 (N_1189,In_381,In_988);
nor U1190 (N_1190,In_847,In_2558);
or U1191 (N_1191,In_924,In_1643);
xor U1192 (N_1192,In_429,In_2362);
xnor U1193 (N_1193,In_1197,In_1523);
xor U1194 (N_1194,In_2425,In_747);
or U1195 (N_1195,In_2915,In_2057);
nand U1196 (N_1196,In_1127,In_2787);
nor U1197 (N_1197,In_311,In_237);
xor U1198 (N_1198,In_1003,In_1303);
nand U1199 (N_1199,In_1307,In_2926);
or U1200 (N_1200,In_2441,In_209);
nor U1201 (N_1201,In_1529,In_396);
or U1202 (N_1202,In_1581,In_2723);
xnor U1203 (N_1203,In_417,In_1135);
nor U1204 (N_1204,In_24,In_106);
xnor U1205 (N_1205,In_2756,In_1227);
or U1206 (N_1206,In_1571,In_744);
xor U1207 (N_1207,In_1293,In_2939);
and U1208 (N_1208,In_1315,In_2214);
xor U1209 (N_1209,In_470,In_2280);
xnor U1210 (N_1210,In_1654,In_309);
or U1211 (N_1211,In_719,In_337);
nand U1212 (N_1212,In_1009,In_1955);
nand U1213 (N_1213,In_2942,In_552);
nand U1214 (N_1214,In_193,In_2315);
or U1215 (N_1215,In_2288,In_1370);
or U1216 (N_1216,In_655,In_215);
or U1217 (N_1217,In_1892,In_409);
or U1218 (N_1218,In_1681,In_947);
nand U1219 (N_1219,In_2066,In_242);
nor U1220 (N_1220,In_1143,In_2943);
nand U1221 (N_1221,In_1652,In_253);
or U1222 (N_1222,In_754,In_1716);
nor U1223 (N_1223,In_1504,In_1992);
and U1224 (N_1224,In_232,In_2754);
xor U1225 (N_1225,In_884,In_424);
or U1226 (N_1226,In_1493,In_2882);
and U1227 (N_1227,In_2639,In_1311);
xnor U1228 (N_1228,In_1965,In_1823);
or U1229 (N_1229,In_359,In_1911);
and U1230 (N_1230,In_75,In_2211);
or U1231 (N_1231,In_1793,In_647);
xor U1232 (N_1232,In_1541,In_48);
nand U1233 (N_1233,In_2813,In_522);
nor U1234 (N_1234,In_1480,In_2418);
and U1235 (N_1235,In_137,In_2811);
nor U1236 (N_1236,In_373,In_313);
nor U1237 (N_1237,In_347,In_1827);
nand U1238 (N_1238,In_2360,In_2829);
nor U1239 (N_1239,In_443,In_1535);
nor U1240 (N_1240,In_2030,In_2431);
and U1241 (N_1241,In_270,In_702);
nor U1242 (N_1242,In_1081,In_1050);
or U1243 (N_1243,In_1968,In_1072);
nor U1244 (N_1244,In_2514,In_17);
xnor U1245 (N_1245,In_1981,In_1165);
or U1246 (N_1246,In_2799,In_686);
xor U1247 (N_1247,In_294,In_2029);
xnor U1248 (N_1248,In_406,In_821);
nor U1249 (N_1249,In_1549,In_1092);
and U1250 (N_1250,In_2233,In_2466);
nor U1251 (N_1251,In_1355,In_2379);
nor U1252 (N_1252,In_1619,In_1104);
nor U1253 (N_1253,In_1629,In_2940);
nor U1254 (N_1254,In_1350,In_1557);
nand U1255 (N_1255,In_2624,In_1340);
xnor U1256 (N_1256,In_540,In_1175);
xor U1257 (N_1257,In_838,In_2812);
nand U1258 (N_1258,In_2833,In_279);
and U1259 (N_1259,In_977,In_2580);
xnor U1260 (N_1260,In_2104,In_1278);
nand U1261 (N_1261,In_1334,In_2607);
nor U1262 (N_1262,In_2310,In_2810);
and U1263 (N_1263,In_1287,In_2927);
and U1264 (N_1264,In_2242,In_97);
xor U1265 (N_1265,In_1405,In_697);
or U1266 (N_1266,In_1924,In_2884);
nor U1267 (N_1267,In_1804,In_2161);
nand U1268 (N_1268,In_216,In_2941);
nor U1269 (N_1269,In_2888,In_2308);
or U1270 (N_1270,In_292,In_846);
nor U1271 (N_1271,In_515,In_1065);
xnor U1272 (N_1272,In_1908,In_2085);
nor U1273 (N_1273,In_1748,In_201);
xnor U1274 (N_1274,In_943,In_2512);
nor U1275 (N_1275,In_1094,In_320);
or U1276 (N_1276,In_2316,In_1111);
or U1277 (N_1277,In_1683,In_210);
xnor U1278 (N_1278,In_1335,In_2058);
nand U1279 (N_1279,In_1869,In_1893);
nor U1280 (N_1280,In_1324,In_1583);
or U1281 (N_1281,In_176,In_1731);
or U1282 (N_1282,In_183,In_2098);
nand U1283 (N_1283,In_519,In_2949);
and U1284 (N_1284,In_2478,In_2059);
or U1285 (N_1285,In_1347,In_377);
and U1286 (N_1286,In_2920,In_467);
or U1287 (N_1287,In_2733,In_968);
nor U1288 (N_1288,In_59,In_2652);
and U1289 (N_1289,In_980,In_1915);
nand U1290 (N_1290,In_929,In_1732);
or U1291 (N_1291,In_1595,In_1547);
xnor U1292 (N_1292,In_491,In_1948);
or U1293 (N_1293,In_1815,In_1709);
xnor U1294 (N_1294,In_2849,In_701);
nand U1295 (N_1295,In_887,In_334);
and U1296 (N_1296,In_903,In_1973);
xor U1297 (N_1297,In_1531,In_2089);
or U1298 (N_1298,In_2635,In_2168);
or U1299 (N_1299,In_756,In_2247);
or U1300 (N_1300,In_1080,In_260);
or U1301 (N_1301,In_2931,In_1813);
nor U1302 (N_1302,In_2557,In_2883);
and U1303 (N_1303,In_2981,In_508);
nor U1304 (N_1304,In_2746,In_900);
or U1305 (N_1305,In_696,In_563);
nand U1306 (N_1306,In_1534,In_280);
nor U1307 (N_1307,In_836,In_2245);
nor U1308 (N_1308,In_936,In_584);
nand U1309 (N_1309,In_2230,In_1608);
or U1310 (N_1310,In_2900,In_2009);
nor U1311 (N_1311,In_958,In_2777);
nand U1312 (N_1312,In_1520,In_1692);
nand U1313 (N_1313,In_2469,In_2323);
xor U1314 (N_1314,In_1906,In_1754);
xor U1315 (N_1315,In_1395,In_1226);
nand U1316 (N_1316,In_332,In_2197);
xnor U1317 (N_1317,In_333,In_2947);
nand U1318 (N_1318,In_419,In_1935);
xor U1319 (N_1319,In_498,In_312);
nor U1320 (N_1320,In_2828,In_1101);
and U1321 (N_1321,In_2608,In_130);
or U1322 (N_1322,In_764,In_496);
nand U1323 (N_1323,In_1778,In_2675);
nand U1324 (N_1324,In_899,In_1757);
or U1325 (N_1325,In_2963,In_1678);
nand U1326 (N_1326,In_338,In_1258);
nor U1327 (N_1327,In_321,In_1695);
and U1328 (N_1328,In_824,In_2282);
nor U1329 (N_1329,In_1482,In_1782);
nand U1330 (N_1330,In_1677,In_1008);
nand U1331 (N_1331,In_1151,In_2475);
or U1332 (N_1332,In_511,In_326);
and U1333 (N_1333,In_2189,In_350);
or U1334 (N_1334,In_741,In_828);
xnor U1335 (N_1335,In_1847,In_2908);
nor U1336 (N_1336,In_555,In_586);
nor U1337 (N_1337,In_2935,In_493);
and U1338 (N_1338,In_856,In_353);
or U1339 (N_1339,In_2937,In_561);
nor U1340 (N_1340,In_2946,In_1791);
nor U1341 (N_1341,In_288,In_638);
xnor U1342 (N_1342,In_2079,In_852);
and U1343 (N_1343,In_2893,In_849);
xor U1344 (N_1344,In_1787,In_490);
xnor U1345 (N_1345,In_2600,In_717);
and U1346 (N_1346,In_412,In_1593);
or U1347 (N_1347,In_1270,In_2713);
or U1348 (N_1348,In_2631,In_1078);
nand U1349 (N_1349,In_1944,In_2576);
nand U1350 (N_1350,In_1208,In_2012);
and U1351 (N_1351,In_2359,In_2612);
and U1352 (N_1352,In_1873,In_889);
xnor U1353 (N_1353,In_1897,In_2790);
nor U1354 (N_1354,In_1487,In_243);
nand U1355 (N_1355,In_2025,In_249);
or U1356 (N_1356,In_1364,In_1154);
or U1357 (N_1357,In_1792,In_2542);
nand U1358 (N_1358,In_1812,In_935);
and U1359 (N_1359,In_2763,In_2411);
xor U1360 (N_1360,In_914,In_1701);
or U1361 (N_1361,In_896,In_144);
xor U1362 (N_1362,In_659,In_2550);
nand U1363 (N_1363,In_2632,In_411);
xnor U1364 (N_1364,In_2818,In_465);
or U1365 (N_1365,In_2730,In_32);
xor U1366 (N_1366,In_2823,In_1926);
xor U1367 (N_1367,In_1020,In_928);
and U1368 (N_1368,In_2855,In_363);
or U1369 (N_1369,In_2587,In_2148);
nand U1370 (N_1370,In_501,In_14);
nor U1371 (N_1371,In_368,In_124);
xor U1372 (N_1372,In_1110,In_40);
nand U1373 (N_1373,In_2693,In_2793);
or U1374 (N_1374,In_1822,In_2347);
and U1375 (N_1375,In_1946,In_1862);
nor U1376 (N_1376,In_2314,In_2369);
xor U1377 (N_1377,In_2253,In_1447);
or U1378 (N_1378,In_2412,In_940);
nand U1379 (N_1379,In_2156,In_2586);
nand U1380 (N_1380,In_622,In_1109);
nor U1381 (N_1381,In_922,In_5);
nor U1382 (N_1382,In_1963,In_989);
nand U1383 (N_1383,In_2522,In_2048);
nor U1384 (N_1384,In_1139,In_2147);
nor U1385 (N_1385,In_589,In_939);
xor U1386 (N_1386,In_2845,In_2867);
nand U1387 (N_1387,In_2984,In_1338);
and U1388 (N_1388,In_1302,In_758);
nor U1389 (N_1389,In_801,In_1131);
or U1390 (N_1390,In_2615,In_414);
nand U1391 (N_1391,In_1789,In_2179);
xnor U1392 (N_1392,In_2195,In_1119);
nor U1393 (N_1393,In_1235,In_2857);
xor U1394 (N_1394,In_1910,In_2007);
nand U1395 (N_1395,In_2402,In_2885);
xnor U1396 (N_1396,In_1031,In_164);
xor U1397 (N_1397,In_2906,In_1798);
nor U1398 (N_1398,In_1453,In_1470);
nand U1399 (N_1399,In_890,In_1150);
and U1400 (N_1400,In_1428,In_205);
or U1401 (N_1401,In_1679,In_1967);
and U1402 (N_1402,In_2289,In_23);
or U1403 (N_1403,In_2916,In_2852);
nor U1404 (N_1404,In_2489,In_2921);
nand U1405 (N_1405,In_2176,In_2914);
and U1406 (N_1406,In_1928,In_1510);
or U1407 (N_1407,In_1669,In_2276);
xor U1408 (N_1408,In_2319,In_2634);
xor U1409 (N_1409,In_1036,In_1484);
or U1410 (N_1410,In_308,In_1490);
nand U1411 (N_1411,In_2243,In_535);
or U1412 (N_1412,In_2317,In_2060);
nor U1413 (N_1413,In_1737,In_2996);
and U1414 (N_1414,In_1914,In_1450);
and U1415 (N_1415,In_1623,In_568);
xnor U1416 (N_1416,In_1644,In_457);
nor U1417 (N_1417,In_1821,In_534);
nand U1418 (N_1418,In_2630,In_2160);
and U1419 (N_1419,In_1579,In_1056);
nor U1420 (N_1420,In_1093,In_1077);
and U1421 (N_1421,In_1245,In_1024);
and U1422 (N_1422,In_274,In_711);
nor U1423 (N_1423,In_2429,In_2708);
and U1424 (N_1424,In_145,In_219);
xor U1425 (N_1425,In_1551,In_1416);
nand U1426 (N_1426,In_886,In_2095);
xor U1427 (N_1427,In_2864,In_1218);
nor U1428 (N_1428,In_657,In_2430);
xor U1429 (N_1429,In_1836,In_873);
and U1430 (N_1430,In_1039,In_978);
and U1431 (N_1431,In_2537,In_2090);
and U1432 (N_1432,In_2141,In_494);
xnor U1433 (N_1433,In_1444,In_495);
nor U1434 (N_1434,In_2255,In_1569);
nand U1435 (N_1435,In_571,In_2710);
and U1436 (N_1436,In_777,In_2595);
and U1437 (N_1437,In_1260,In_2526);
xnor U1438 (N_1438,In_623,In_1537);
nand U1439 (N_1439,In_1628,In_775);
nand U1440 (N_1440,In_857,In_152);
xnor U1441 (N_1441,In_1361,In_1607);
and U1442 (N_1442,In_33,In_262);
nand U1443 (N_1443,In_1561,In_681);
and U1444 (N_1444,In_1014,In_1331);
and U1445 (N_1445,In_1974,In_1564);
nor U1446 (N_1446,In_2944,In_22);
nor U1447 (N_1447,In_2641,In_912);
nand U1448 (N_1448,In_352,In_918);
and U1449 (N_1449,In_2170,In_593);
nand U1450 (N_1450,In_328,In_1640);
nor U1451 (N_1451,In_2785,In_2279);
nand U1452 (N_1452,In_2501,In_844);
and U1453 (N_1453,In_1978,In_1063);
nor U1454 (N_1454,In_2283,In_361);
or U1455 (N_1455,In_2960,In_1542);
nand U1456 (N_1456,In_1029,In_550);
nor U1457 (N_1457,In_2235,In_2145);
nor U1458 (N_1458,In_1272,In_88);
nor U1459 (N_1459,In_418,In_2834);
xor U1460 (N_1460,In_2497,In_1146);
or U1461 (N_1461,In_1001,In_1400);
nand U1462 (N_1462,In_2149,In_2954);
xor U1463 (N_1463,In_1432,In_266);
and U1464 (N_1464,In_1575,In_1268);
nor U1465 (N_1465,In_2232,In_2097);
nor U1466 (N_1466,In_1785,In_578);
nor U1467 (N_1467,In_1743,In_680);
and U1468 (N_1468,In_2249,In_2815);
xor U1469 (N_1469,In_784,In_603);
or U1470 (N_1470,In_314,In_2581);
and U1471 (N_1471,In_808,In_1706);
nor U1472 (N_1472,In_463,In_244);
xor U1473 (N_1473,In_675,In_2767);
or U1474 (N_1474,In_212,In_2134);
nor U1475 (N_1475,In_626,In_504);
xor U1476 (N_1476,In_2751,In_1984);
xor U1477 (N_1477,In_2306,In_2868);
nor U1478 (N_1478,In_1431,In_2593);
or U1479 (N_1479,In_2390,In_1634);
or U1480 (N_1480,In_35,In_2958);
nor U1481 (N_1481,In_1378,In_648);
or U1482 (N_1482,In_2228,In_538);
nand U1483 (N_1483,In_605,In_2216);
and U1484 (N_1484,In_1368,In_1829);
nand U1485 (N_1485,In_2107,In_2175);
xor U1486 (N_1486,In_1846,In_1949);
nand U1487 (N_1487,In_2150,In_268);
nor U1488 (N_1488,In_1481,In_153);
or U1489 (N_1489,In_1882,In_2393);
or U1490 (N_1490,In_2470,In_1044);
and U1491 (N_1491,In_2343,In_1664);
or U1492 (N_1492,In_865,In_806);
or U1493 (N_1493,In_505,In_1156);
xor U1494 (N_1494,In_2199,In_401);
or U1495 (N_1495,In_1130,In_1499);
nand U1496 (N_1496,In_2376,In_1309);
or U1497 (N_1497,In_407,In_1597);
nor U1498 (N_1498,In_2386,In_1603);
nor U1499 (N_1499,In_1521,In_2364);
nand U1500 (N_1500,In_1782,In_1369);
or U1501 (N_1501,In_941,In_1774);
xnor U1502 (N_1502,In_2672,In_2403);
or U1503 (N_1503,In_2635,In_1645);
xor U1504 (N_1504,In_2895,In_690);
nor U1505 (N_1505,In_25,In_786);
and U1506 (N_1506,In_2730,In_1175);
xor U1507 (N_1507,In_532,In_1530);
nand U1508 (N_1508,In_109,In_1389);
nor U1509 (N_1509,In_1386,In_405);
or U1510 (N_1510,In_1199,In_2949);
xor U1511 (N_1511,In_1682,In_1014);
nand U1512 (N_1512,In_823,In_1240);
and U1513 (N_1513,In_2769,In_280);
nor U1514 (N_1514,In_1474,In_2177);
nor U1515 (N_1515,In_2696,In_702);
or U1516 (N_1516,In_1099,In_676);
nor U1517 (N_1517,In_2650,In_1249);
xor U1518 (N_1518,In_1510,In_576);
or U1519 (N_1519,In_2558,In_365);
and U1520 (N_1520,In_2500,In_1018);
or U1521 (N_1521,In_334,In_583);
xnor U1522 (N_1522,In_1151,In_2229);
nor U1523 (N_1523,In_675,In_1783);
and U1524 (N_1524,In_1848,In_1024);
xnor U1525 (N_1525,In_1973,In_1685);
and U1526 (N_1526,In_1341,In_811);
nor U1527 (N_1527,In_2901,In_2288);
nor U1528 (N_1528,In_671,In_2232);
or U1529 (N_1529,In_2896,In_2726);
and U1530 (N_1530,In_88,In_2705);
xnor U1531 (N_1531,In_1805,In_363);
and U1532 (N_1532,In_883,In_865);
nand U1533 (N_1533,In_846,In_388);
and U1534 (N_1534,In_995,In_2665);
xor U1535 (N_1535,In_277,In_2521);
and U1536 (N_1536,In_479,In_1140);
nor U1537 (N_1537,In_1692,In_1958);
nand U1538 (N_1538,In_718,In_916);
or U1539 (N_1539,In_1699,In_625);
and U1540 (N_1540,In_1961,In_1436);
or U1541 (N_1541,In_2815,In_1345);
nand U1542 (N_1542,In_2981,In_2461);
and U1543 (N_1543,In_1130,In_1375);
or U1544 (N_1544,In_2371,In_2349);
nor U1545 (N_1545,In_2464,In_1959);
or U1546 (N_1546,In_2112,In_1232);
or U1547 (N_1547,In_1532,In_2418);
and U1548 (N_1548,In_2336,In_2619);
or U1549 (N_1549,In_1391,In_1939);
xnor U1550 (N_1550,In_448,In_1001);
and U1551 (N_1551,In_2486,In_2625);
nand U1552 (N_1552,In_2760,In_2634);
nand U1553 (N_1553,In_792,In_780);
xor U1554 (N_1554,In_866,In_1182);
nand U1555 (N_1555,In_1405,In_1925);
nand U1556 (N_1556,In_1704,In_1342);
xor U1557 (N_1557,In_411,In_1662);
nand U1558 (N_1558,In_1097,In_449);
xor U1559 (N_1559,In_1938,In_121);
xnor U1560 (N_1560,In_1770,In_863);
or U1561 (N_1561,In_1225,In_2795);
or U1562 (N_1562,In_2737,In_995);
and U1563 (N_1563,In_1865,In_2516);
xnor U1564 (N_1564,In_1091,In_1423);
or U1565 (N_1565,In_239,In_754);
and U1566 (N_1566,In_2669,In_470);
nor U1567 (N_1567,In_1321,In_2423);
nand U1568 (N_1568,In_2713,In_2896);
nor U1569 (N_1569,In_1394,In_1338);
nand U1570 (N_1570,In_420,In_1088);
nand U1571 (N_1571,In_1553,In_288);
and U1572 (N_1572,In_1116,In_2463);
xnor U1573 (N_1573,In_1858,In_267);
and U1574 (N_1574,In_1687,In_685);
nor U1575 (N_1575,In_2699,In_297);
xor U1576 (N_1576,In_209,In_470);
xnor U1577 (N_1577,In_1074,In_677);
and U1578 (N_1578,In_1711,In_2760);
nor U1579 (N_1579,In_2012,In_2972);
xor U1580 (N_1580,In_2557,In_2684);
and U1581 (N_1581,In_2724,In_1069);
nor U1582 (N_1582,In_2295,In_972);
and U1583 (N_1583,In_1396,In_454);
or U1584 (N_1584,In_646,In_935);
nand U1585 (N_1585,In_1212,In_2512);
or U1586 (N_1586,In_437,In_566);
or U1587 (N_1587,In_735,In_1774);
nand U1588 (N_1588,In_2086,In_1612);
or U1589 (N_1589,In_1814,In_54);
xor U1590 (N_1590,In_1489,In_2038);
xor U1591 (N_1591,In_2308,In_969);
xnor U1592 (N_1592,In_1941,In_580);
nand U1593 (N_1593,In_84,In_2684);
or U1594 (N_1594,In_2635,In_1398);
or U1595 (N_1595,In_1018,In_1292);
nand U1596 (N_1596,In_1465,In_2061);
nor U1597 (N_1597,In_2210,In_1007);
nand U1598 (N_1598,In_607,In_2225);
and U1599 (N_1599,In_275,In_2633);
nand U1600 (N_1600,In_360,In_11);
or U1601 (N_1601,In_1958,In_732);
xor U1602 (N_1602,In_1858,In_1719);
nor U1603 (N_1603,In_1473,In_2374);
and U1604 (N_1604,In_778,In_1808);
nor U1605 (N_1605,In_1039,In_1299);
and U1606 (N_1606,In_863,In_1121);
nor U1607 (N_1607,In_2151,In_2405);
xnor U1608 (N_1608,In_1136,In_1232);
xor U1609 (N_1609,In_2242,In_1480);
and U1610 (N_1610,In_1373,In_953);
or U1611 (N_1611,In_2695,In_195);
or U1612 (N_1612,In_2052,In_340);
xor U1613 (N_1613,In_1917,In_2947);
or U1614 (N_1614,In_569,In_1639);
or U1615 (N_1615,In_2779,In_1818);
nor U1616 (N_1616,In_2125,In_675);
or U1617 (N_1617,In_1718,In_275);
or U1618 (N_1618,In_439,In_1554);
xnor U1619 (N_1619,In_1969,In_145);
nor U1620 (N_1620,In_570,In_473);
or U1621 (N_1621,In_467,In_2504);
nor U1622 (N_1622,In_311,In_1257);
or U1623 (N_1623,In_1772,In_2950);
xnor U1624 (N_1624,In_1157,In_1383);
xor U1625 (N_1625,In_2751,In_59);
nor U1626 (N_1626,In_2215,In_2834);
nor U1627 (N_1627,In_1025,In_1042);
and U1628 (N_1628,In_1632,In_173);
nand U1629 (N_1629,In_2353,In_720);
nand U1630 (N_1630,In_321,In_1795);
nor U1631 (N_1631,In_549,In_60);
xnor U1632 (N_1632,In_1579,In_1163);
nand U1633 (N_1633,In_1717,In_199);
or U1634 (N_1634,In_2266,In_2766);
nor U1635 (N_1635,In_1131,In_2034);
nand U1636 (N_1636,In_1601,In_2329);
xor U1637 (N_1637,In_2934,In_2183);
and U1638 (N_1638,In_1323,In_2978);
nand U1639 (N_1639,In_858,In_627);
nor U1640 (N_1640,In_1323,In_2289);
or U1641 (N_1641,In_2555,In_760);
nor U1642 (N_1642,In_2408,In_17);
xor U1643 (N_1643,In_467,In_2555);
nor U1644 (N_1644,In_1321,In_140);
xor U1645 (N_1645,In_381,In_1741);
and U1646 (N_1646,In_2338,In_1269);
or U1647 (N_1647,In_1805,In_1166);
or U1648 (N_1648,In_1104,In_2136);
nor U1649 (N_1649,In_1875,In_1871);
nor U1650 (N_1650,In_482,In_2282);
or U1651 (N_1651,In_585,In_1897);
and U1652 (N_1652,In_1455,In_558);
nor U1653 (N_1653,In_1485,In_2194);
or U1654 (N_1654,In_2294,In_2050);
nor U1655 (N_1655,In_424,In_265);
xor U1656 (N_1656,In_29,In_26);
or U1657 (N_1657,In_988,In_497);
nor U1658 (N_1658,In_554,In_2219);
and U1659 (N_1659,In_151,In_1380);
nor U1660 (N_1660,In_2526,In_1941);
nand U1661 (N_1661,In_1754,In_1648);
xnor U1662 (N_1662,In_2897,In_1433);
nand U1663 (N_1663,In_1995,In_38);
and U1664 (N_1664,In_688,In_1773);
nand U1665 (N_1665,In_28,In_1186);
nand U1666 (N_1666,In_577,In_958);
nor U1667 (N_1667,In_1596,In_2684);
xor U1668 (N_1668,In_790,In_6);
or U1669 (N_1669,In_2657,In_1376);
or U1670 (N_1670,In_334,In_2587);
or U1671 (N_1671,In_758,In_2587);
and U1672 (N_1672,In_2788,In_1612);
nand U1673 (N_1673,In_1446,In_1805);
or U1674 (N_1674,In_1737,In_2961);
nand U1675 (N_1675,In_204,In_1025);
and U1676 (N_1676,In_706,In_879);
and U1677 (N_1677,In_165,In_423);
and U1678 (N_1678,In_1907,In_2312);
nand U1679 (N_1679,In_1010,In_1880);
and U1680 (N_1680,In_1839,In_874);
xnor U1681 (N_1681,In_172,In_2763);
nor U1682 (N_1682,In_1955,In_2044);
nand U1683 (N_1683,In_2797,In_1673);
nor U1684 (N_1684,In_1204,In_281);
xor U1685 (N_1685,In_100,In_1909);
or U1686 (N_1686,In_557,In_731);
or U1687 (N_1687,In_697,In_2603);
nor U1688 (N_1688,In_2648,In_1202);
and U1689 (N_1689,In_1634,In_1690);
and U1690 (N_1690,In_1122,In_2567);
nor U1691 (N_1691,In_2590,In_1976);
or U1692 (N_1692,In_1893,In_2431);
nand U1693 (N_1693,In_238,In_2654);
and U1694 (N_1694,In_2991,In_245);
nor U1695 (N_1695,In_2256,In_1497);
or U1696 (N_1696,In_120,In_429);
or U1697 (N_1697,In_2912,In_2429);
nand U1698 (N_1698,In_1868,In_2476);
and U1699 (N_1699,In_2863,In_569);
nand U1700 (N_1700,In_2149,In_508);
nand U1701 (N_1701,In_499,In_2232);
and U1702 (N_1702,In_2422,In_2830);
nand U1703 (N_1703,In_2116,In_2066);
nor U1704 (N_1704,In_1385,In_1823);
and U1705 (N_1705,In_266,In_629);
nor U1706 (N_1706,In_2450,In_2368);
or U1707 (N_1707,In_1237,In_827);
xnor U1708 (N_1708,In_1421,In_174);
or U1709 (N_1709,In_31,In_1219);
xnor U1710 (N_1710,In_1052,In_1401);
xnor U1711 (N_1711,In_1954,In_1335);
or U1712 (N_1712,In_1446,In_2528);
or U1713 (N_1713,In_685,In_2636);
xor U1714 (N_1714,In_2329,In_1244);
nor U1715 (N_1715,In_732,In_1178);
and U1716 (N_1716,In_457,In_44);
and U1717 (N_1717,In_78,In_343);
nand U1718 (N_1718,In_976,In_1650);
nand U1719 (N_1719,In_444,In_1678);
nand U1720 (N_1720,In_883,In_2338);
nor U1721 (N_1721,In_2355,In_2177);
xor U1722 (N_1722,In_979,In_1104);
xnor U1723 (N_1723,In_2136,In_1572);
xor U1724 (N_1724,In_879,In_1348);
xor U1725 (N_1725,In_2597,In_913);
or U1726 (N_1726,In_991,In_1818);
nand U1727 (N_1727,In_961,In_2983);
and U1728 (N_1728,In_1750,In_2374);
or U1729 (N_1729,In_673,In_1875);
nor U1730 (N_1730,In_2324,In_1562);
and U1731 (N_1731,In_2390,In_514);
xnor U1732 (N_1732,In_411,In_632);
nor U1733 (N_1733,In_1384,In_2127);
or U1734 (N_1734,In_593,In_1233);
xor U1735 (N_1735,In_678,In_1521);
xor U1736 (N_1736,In_1615,In_2726);
or U1737 (N_1737,In_2518,In_1976);
nand U1738 (N_1738,In_2626,In_2366);
xor U1739 (N_1739,In_388,In_1101);
and U1740 (N_1740,In_178,In_1173);
and U1741 (N_1741,In_1950,In_2475);
xor U1742 (N_1742,In_174,In_766);
xnor U1743 (N_1743,In_1706,In_585);
nor U1744 (N_1744,In_2330,In_2784);
and U1745 (N_1745,In_1748,In_1710);
xnor U1746 (N_1746,In_1304,In_2866);
and U1747 (N_1747,In_1493,In_2451);
nand U1748 (N_1748,In_2687,In_2646);
nand U1749 (N_1749,In_1684,In_2941);
xor U1750 (N_1750,In_2077,In_1984);
nor U1751 (N_1751,In_996,In_1912);
nor U1752 (N_1752,In_2440,In_567);
nand U1753 (N_1753,In_2103,In_212);
xnor U1754 (N_1754,In_23,In_319);
nor U1755 (N_1755,In_2410,In_919);
or U1756 (N_1756,In_2847,In_2624);
nor U1757 (N_1757,In_1058,In_809);
xor U1758 (N_1758,In_1678,In_157);
or U1759 (N_1759,In_2243,In_64);
nor U1760 (N_1760,In_844,In_560);
or U1761 (N_1761,In_110,In_1135);
xnor U1762 (N_1762,In_1852,In_1053);
nand U1763 (N_1763,In_2073,In_1243);
nor U1764 (N_1764,In_2059,In_360);
nand U1765 (N_1765,In_614,In_1932);
xnor U1766 (N_1766,In_798,In_2291);
xnor U1767 (N_1767,In_310,In_1129);
and U1768 (N_1768,In_1300,In_1592);
xor U1769 (N_1769,In_1198,In_676);
nor U1770 (N_1770,In_2893,In_561);
nor U1771 (N_1771,In_2841,In_2131);
nor U1772 (N_1772,In_2662,In_1959);
or U1773 (N_1773,In_1030,In_894);
and U1774 (N_1774,In_17,In_405);
and U1775 (N_1775,In_2739,In_1905);
and U1776 (N_1776,In_2445,In_2222);
xor U1777 (N_1777,In_785,In_1550);
and U1778 (N_1778,In_393,In_1923);
nand U1779 (N_1779,In_89,In_43);
and U1780 (N_1780,In_1733,In_296);
nor U1781 (N_1781,In_2938,In_1341);
or U1782 (N_1782,In_1138,In_2402);
nor U1783 (N_1783,In_934,In_2591);
and U1784 (N_1784,In_465,In_1905);
xnor U1785 (N_1785,In_1624,In_1672);
or U1786 (N_1786,In_40,In_1287);
xnor U1787 (N_1787,In_292,In_2887);
xnor U1788 (N_1788,In_821,In_1638);
or U1789 (N_1789,In_142,In_2207);
nor U1790 (N_1790,In_1418,In_2887);
nand U1791 (N_1791,In_2200,In_501);
or U1792 (N_1792,In_2304,In_839);
xnor U1793 (N_1793,In_2627,In_398);
and U1794 (N_1794,In_2476,In_1896);
xor U1795 (N_1795,In_820,In_869);
and U1796 (N_1796,In_860,In_2499);
and U1797 (N_1797,In_2322,In_1963);
xor U1798 (N_1798,In_202,In_2281);
xor U1799 (N_1799,In_542,In_1483);
and U1800 (N_1800,In_2867,In_1096);
xnor U1801 (N_1801,In_1990,In_2788);
xnor U1802 (N_1802,In_2287,In_1138);
nor U1803 (N_1803,In_1358,In_1338);
xnor U1804 (N_1804,In_2775,In_743);
and U1805 (N_1805,In_1393,In_2276);
xor U1806 (N_1806,In_2332,In_1690);
nand U1807 (N_1807,In_2303,In_2086);
nor U1808 (N_1808,In_1293,In_579);
nor U1809 (N_1809,In_379,In_1481);
nand U1810 (N_1810,In_1709,In_1888);
nand U1811 (N_1811,In_1856,In_2942);
and U1812 (N_1812,In_577,In_791);
nor U1813 (N_1813,In_2148,In_2216);
and U1814 (N_1814,In_1860,In_1840);
xor U1815 (N_1815,In_55,In_81);
and U1816 (N_1816,In_1409,In_1018);
or U1817 (N_1817,In_1021,In_2251);
xnor U1818 (N_1818,In_1755,In_2220);
nand U1819 (N_1819,In_372,In_2885);
nand U1820 (N_1820,In_2315,In_2375);
or U1821 (N_1821,In_1148,In_2894);
nand U1822 (N_1822,In_1051,In_2128);
nor U1823 (N_1823,In_2011,In_2630);
or U1824 (N_1824,In_410,In_822);
xnor U1825 (N_1825,In_1879,In_1937);
and U1826 (N_1826,In_808,In_2998);
or U1827 (N_1827,In_2810,In_1947);
or U1828 (N_1828,In_1179,In_2294);
or U1829 (N_1829,In_848,In_1665);
nand U1830 (N_1830,In_1081,In_1744);
or U1831 (N_1831,In_1853,In_688);
and U1832 (N_1832,In_38,In_739);
or U1833 (N_1833,In_1925,In_2652);
or U1834 (N_1834,In_2236,In_2426);
xnor U1835 (N_1835,In_1074,In_1514);
or U1836 (N_1836,In_2779,In_1522);
nor U1837 (N_1837,In_2830,In_2444);
or U1838 (N_1838,In_2369,In_1483);
and U1839 (N_1839,In_1285,In_549);
xnor U1840 (N_1840,In_432,In_2785);
nand U1841 (N_1841,In_144,In_2693);
or U1842 (N_1842,In_2009,In_517);
xnor U1843 (N_1843,In_2493,In_471);
nor U1844 (N_1844,In_332,In_215);
or U1845 (N_1845,In_470,In_613);
nor U1846 (N_1846,In_2947,In_699);
xnor U1847 (N_1847,In_1629,In_2667);
nand U1848 (N_1848,In_1028,In_759);
or U1849 (N_1849,In_2428,In_25);
xnor U1850 (N_1850,In_306,In_1446);
and U1851 (N_1851,In_885,In_2395);
nand U1852 (N_1852,In_1958,In_537);
nor U1853 (N_1853,In_1591,In_867);
nand U1854 (N_1854,In_2064,In_2086);
or U1855 (N_1855,In_202,In_265);
or U1856 (N_1856,In_2820,In_716);
or U1857 (N_1857,In_1562,In_2932);
nand U1858 (N_1858,In_2521,In_392);
and U1859 (N_1859,In_54,In_100);
xnor U1860 (N_1860,In_1582,In_2259);
or U1861 (N_1861,In_1481,In_989);
nand U1862 (N_1862,In_2347,In_47);
and U1863 (N_1863,In_1118,In_868);
nor U1864 (N_1864,In_923,In_1172);
nand U1865 (N_1865,In_224,In_263);
and U1866 (N_1866,In_1400,In_31);
xor U1867 (N_1867,In_2212,In_1792);
xor U1868 (N_1868,In_1838,In_1580);
nand U1869 (N_1869,In_395,In_793);
xnor U1870 (N_1870,In_59,In_860);
or U1871 (N_1871,In_2434,In_14);
and U1872 (N_1872,In_2834,In_1496);
and U1873 (N_1873,In_1183,In_163);
or U1874 (N_1874,In_450,In_647);
and U1875 (N_1875,In_500,In_2467);
and U1876 (N_1876,In_1023,In_414);
xor U1877 (N_1877,In_1475,In_2438);
nor U1878 (N_1878,In_2676,In_2223);
or U1879 (N_1879,In_774,In_2339);
nor U1880 (N_1880,In_701,In_1240);
xor U1881 (N_1881,In_11,In_399);
nand U1882 (N_1882,In_2540,In_692);
nor U1883 (N_1883,In_1004,In_432);
and U1884 (N_1884,In_1459,In_1818);
or U1885 (N_1885,In_2464,In_894);
or U1886 (N_1886,In_82,In_241);
nand U1887 (N_1887,In_2775,In_2763);
and U1888 (N_1888,In_2942,In_233);
xnor U1889 (N_1889,In_1279,In_2341);
nor U1890 (N_1890,In_228,In_413);
and U1891 (N_1891,In_854,In_1502);
nand U1892 (N_1892,In_2325,In_1641);
nand U1893 (N_1893,In_2095,In_1338);
and U1894 (N_1894,In_279,In_909);
and U1895 (N_1895,In_595,In_682);
xnor U1896 (N_1896,In_2728,In_2362);
nand U1897 (N_1897,In_891,In_1242);
and U1898 (N_1898,In_1027,In_2990);
xor U1899 (N_1899,In_1017,In_2299);
nand U1900 (N_1900,In_2152,In_226);
xnor U1901 (N_1901,In_1432,In_1699);
xor U1902 (N_1902,In_2978,In_123);
nor U1903 (N_1903,In_2687,In_2071);
and U1904 (N_1904,In_265,In_2540);
or U1905 (N_1905,In_1158,In_1776);
or U1906 (N_1906,In_43,In_470);
nor U1907 (N_1907,In_422,In_336);
nand U1908 (N_1908,In_1250,In_2356);
nand U1909 (N_1909,In_1495,In_411);
or U1910 (N_1910,In_1177,In_2272);
xnor U1911 (N_1911,In_2920,In_2613);
nor U1912 (N_1912,In_1370,In_53);
or U1913 (N_1913,In_254,In_2851);
nand U1914 (N_1914,In_1318,In_2212);
nand U1915 (N_1915,In_1069,In_535);
nand U1916 (N_1916,In_949,In_2400);
nand U1917 (N_1917,In_875,In_547);
or U1918 (N_1918,In_1976,In_84);
nor U1919 (N_1919,In_1749,In_952);
or U1920 (N_1920,In_1684,In_289);
or U1921 (N_1921,In_2434,In_2331);
xor U1922 (N_1922,In_1167,In_76);
xnor U1923 (N_1923,In_2759,In_2050);
nor U1924 (N_1924,In_422,In_2717);
nor U1925 (N_1925,In_283,In_27);
or U1926 (N_1926,In_883,In_1670);
nor U1927 (N_1927,In_2851,In_1570);
xor U1928 (N_1928,In_2392,In_2615);
xnor U1929 (N_1929,In_116,In_2376);
nor U1930 (N_1930,In_1253,In_1539);
and U1931 (N_1931,In_695,In_467);
xnor U1932 (N_1932,In_1227,In_1711);
nor U1933 (N_1933,In_1471,In_253);
xor U1934 (N_1934,In_241,In_1956);
nor U1935 (N_1935,In_2306,In_648);
or U1936 (N_1936,In_317,In_2183);
or U1937 (N_1937,In_765,In_2919);
or U1938 (N_1938,In_1340,In_207);
nor U1939 (N_1939,In_1768,In_1794);
and U1940 (N_1940,In_1174,In_63);
and U1941 (N_1941,In_1866,In_675);
or U1942 (N_1942,In_161,In_418);
and U1943 (N_1943,In_1192,In_1637);
or U1944 (N_1944,In_787,In_1164);
nand U1945 (N_1945,In_457,In_298);
or U1946 (N_1946,In_957,In_1072);
xor U1947 (N_1947,In_260,In_2121);
or U1948 (N_1948,In_2233,In_1902);
nor U1949 (N_1949,In_1810,In_901);
nor U1950 (N_1950,In_2364,In_67);
nor U1951 (N_1951,In_2734,In_1948);
xor U1952 (N_1952,In_2505,In_2933);
and U1953 (N_1953,In_1331,In_1006);
xnor U1954 (N_1954,In_1089,In_394);
nor U1955 (N_1955,In_30,In_2359);
and U1956 (N_1956,In_962,In_543);
nand U1957 (N_1957,In_2933,In_1655);
and U1958 (N_1958,In_1109,In_1285);
and U1959 (N_1959,In_1140,In_824);
and U1960 (N_1960,In_219,In_2069);
nor U1961 (N_1961,In_2139,In_2144);
nor U1962 (N_1962,In_297,In_2492);
and U1963 (N_1963,In_140,In_2732);
nor U1964 (N_1964,In_32,In_87);
and U1965 (N_1965,In_1140,In_284);
nand U1966 (N_1966,In_2243,In_1106);
xor U1967 (N_1967,In_2352,In_103);
nor U1968 (N_1968,In_2181,In_2660);
nand U1969 (N_1969,In_775,In_2253);
and U1970 (N_1970,In_1271,In_2617);
or U1971 (N_1971,In_2903,In_786);
xnor U1972 (N_1972,In_832,In_737);
or U1973 (N_1973,In_626,In_1945);
xnor U1974 (N_1974,In_2416,In_1200);
or U1975 (N_1975,In_264,In_39);
xor U1976 (N_1976,In_2938,In_1822);
xnor U1977 (N_1977,In_1082,In_2317);
nand U1978 (N_1978,In_385,In_2470);
nor U1979 (N_1979,In_1769,In_2314);
or U1980 (N_1980,In_2484,In_2986);
nor U1981 (N_1981,In_9,In_1246);
and U1982 (N_1982,In_2784,In_2648);
or U1983 (N_1983,In_1242,In_2360);
xor U1984 (N_1984,In_1935,In_1386);
xnor U1985 (N_1985,In_1314,In_165);
xor U1986 (N_1986,In_1895,In_1426);
and U1987 (N_1987,In_989,In_124);
nor U1988 (N_1988,In_2927,In_561);
or U1989 (N_1989,In_746,In_2063);
nand U1990 (N_1990,In_1287,In_2387);
nand U1991 (N_1991,In_1117,In_749);
and U1992 (N_1992,In_80,In_1717);
nor U1993 (N_1993,In_164,In_2897);
nand U1994 (N_1994,In_569,In_1230);
or U1995 (N_1995,In_489,In_916);
nand U1996 (N_1996,In_426,In_1214);
xor U1997 (N_1997,In_1367,In_2977);
nand U1998 (N_1998,In_2108,In_2408);
xnor U1999 (N_1999,In_835,In_2490);
xor U2000 (N_2000,N_641,N_1655);
nor U2001 (N_2001,N_1596,N_1196);
xor U2002 (N_2002,N_1700,N_1769);
nor U2003 (N_2003,N_297,N_809);
nand U2004 (N_2004,N_598,N_1846);
nor U2005 (N_2005,N_1699,N_697);
or U2006 (N_2006,N_1938,N_211);
or U2007 (N_2007,N_862,N_249);
or U2008 (N_2008,N_535,N_1042);
xnor U2009 (N_2009,N_1189,N_1997);
nand U2010 (N_2010,N_1979,N_780);
xor U2011 (N_2011,N_1236,N_1133);
or U2012 (N_2012,N_715,N_658);
nand U2013 (N_2013,N_1030,N_247);
or U2014 (N_2014,N_1705,N_1487);
nand U2015 (N_2015,N_37,N_123);
nor U2016 (N_2016,N_986,N_511);
or U2017 (N_2017,N_1695,N_1607);
xor U2018 (N_2018,N_1973,N_1474);
and U2019 (N_2019,N_976,N_1867);
or U2020 (N_2020,N_806,N_1527);
or U2021 (N_2021,N_1721,N_1959);
and U2022 (N_2022,N_1424,N_1711);
nand U2023 (N_2023,N_837,N_280);
nor U2024 (N_2024,N_1730,N_1896);
nand U2025 (N_2025,N_1082,N_712);
nor U2026 (N_2026,N_1638,N_64);
or U2027 (N_2027,N_753,N_1334);
nand U2028 (N_2028,N_790,N_952);
or U2029 (N_2029,N_1281,N_133);
nand U2030 (N_2030,N_201,N_492);
nand U2031 (N_2031,N_782,N_1900);
nor U2032 (N_2032,N_531,N_510);
nor U2033 (N_2033,N_1104,N_361);
nor U2034 (N_2034,N_198,N_626);
xnor U2035 (N_2035,N_538,N_437);
or U2036 (N_2036,N_1963,N_1460);
nand U2037 (N_2037,N_1007,N_891);
xor U2038 (N_2038,N_1983,N_1112);
or U2039 (N_2039,N_518,N_1568);
xor U2040 (N_2040,N_1839,N_1817);
and U2041 (N_2041,N_1138,N_487);
or U2042 (N_2042,N_663,N_1593);
and U2043 (N_2043,N_1388,N_1457);
nand U2044 (N_2044,N_1767,N_1078);
and U2045 (N_2045,N_1520,N_1032);
nand U2046 (N_2046,N_1562,N_26);
or U2047 (N_2047,N_114,N_1701);
and U2048 (N_2048,N_334,N_764);
nand U2049 (N_2049,N_1167,N_371);
xor U2050 (N_2050,N_556,N_1110);
or U2051 (N_2051,N_1759,N_1871);
nor U2052 (N_2052,N_1360,N_1355);
or U2053 (N_2053,N_345,N_1768);
nand U2054 (N_2054,N_86,N_933);
xor U2055 (N_2055,N_1774,N_398);
xor U2056 (N_2056,N_1116,N_257);
nand U2057 (N_2057,N_634,N_1830);
xnor U2058 (N_2058,N_1845,N_1234);
nor U2059 (N_2059,N_754,N_1881);
and U2060 (N_2060,N_909,N_328);
and U2061 (N_2061,N_1416,N_668);
nor U2062 (N_2062,N_1047,N_102);
and U2063 (N_2063,N_536,N_1375);
nor U2064 (N_2064,N_530,N_585);
or U2065 (N_2065,N_901,N_1980);
xnor U2066 (N_2066,N_935,N_1976);
nor U2067 (N_2067,N_84,N_1913);
xor U2068 (N_2068,N_1089,N_1788);
nor U2069 (N_2069,N_713,N_1930);
or U2070 (N_2070,N_1405,N_252);
nand U2071 (N_2071,N_1569,N_1223);
and U2072 (N_2072,N_1164,N_843);
nor U2073 (N_2073,N_1456,N_880);
nand U2074 (N_2074,N_1458,N_691);
nor U2075 (N_2075,N_919,N_484);
or U2076 (N_2076,N_745,N_1296);
or U2077 (N_2077,N_1622,N_1159);
nand U2078 (N_2078,N_564,N_1381);
nor U2079 (N_2079,N_240,N_409);
nor U2080 (N_2080,N_1464,N_647);
and U2081 (N_2081,N_1273,N_1378);
nand U2082 (N_2082,N_509,N_1827);
nor U2083 (N_2083,N_840,N_268);
nand U2084 (N_2084,N_769,N_228);
and U2085 (N_2085,N_229,N_1544);
or U2086 (N_2086,N_1861,N_597);
or U2087 (N_2087,N_338,N_418);
and U2088 (N_2088,N_822,N_78);
nor U2089 (N_2089,N_905,N_747);
or U2090 (N_2090,N_273,N_1433);
nor U2091 (N_2091,N_355,N_205);
nor U2092 (N_2092,N_548,N_230);
nand U2093 (N_2093,N_1,N_1087);
and U2094 (N_2094,N_354,N_650);
or U2095 (N_2095,N_1175,N_360);
xnor U2096 (N_2096,N_235,N_233);
nand U2097 (N_2097,N_636,N_1821);
and U2098 (N_2098,N_161,N_1735);
nand U2099 (N_2099,N_1123,N_1937);
nand U2100 (N_2100,N_287,N_471);
and U2101 (N_2101,N_956,N_1782);
and U2102 (N_2102,N_1750,N_1960);
or U2103 (N_2103,N_802,N_794);
nand U2104 (N_2104,N_1998,N_1688);
nand U2105 (N_2105,N_1583,N_1842);
nand U2106 (N_2106,N_610,N_278);
or U2107 (N_2107,N_567,N_512);
nand U2108 (N_2108,N_1518,N_1214);
xor U2109 (N_2109,N_299,N_1131);
nor U2110 (N_2110,N_523,N_1329);
or U2111 (N_2111,N_1323,N_993);
nor U2112 (N_2112,N_340,N_662);
and U2113 (N_2113,N_20,N_1805);
nand U2114 (N_2114,N_1801,N_13);
and U2115 (N_2115,N_1708,N_62);
and U2116 (N_2116,N_131,N_7);
xor U2117 (N_2117,N_331,N_61);
xnor U2118 (N_2118,N_476,N_803);
xor U2119 (N_2119,N_683,N_1027);
nand U2120 (N_2120,N_1964,N_1529);
and U2121 (N_2121,N_1256,N_871);
or U2122 (N_2122,N_1485,N_1860);
nand U2123 (N_2123,N_458,N_337);
nand U2124 (N_2124,N_895,N_736);
nor U2125 (N_2125,N_1102,N_1080);
nor U2126 (N_2126,N_1865,N_1417);
or U2127 (N_2127,N_56,N_990);
xor U2128 (N_2128,N_357,N_1951);
nand U2129 (N_2129,N_1363,N_1336);
nor U2130 (N_2130,N_846,N_1307);
or U2131 (N_2131,N_1247,N_391);
and U2132 (N_2132,N_1429,N_282);
xor U2133 (N_2133,N_1859,N_1357);
or U2134 (N_2134,N_1362,N_1193);
and U2135 (N_2135,N_559,N_711);
and U2136 (N_2136,N_592,N_1057);
nor U2137 (N_2137,N_1269,N_1358);
xor U2138 (N_2138,N_529,N_1887);
or U2139 (N_2139,N_8,N_1035);
xnor U2140 (N_2140,N_1898,N_1576);
nor U2141 (N_2141,N_1286,N_1284);
nand U2142 (N_2142,N_914,N_600);
and U2143 (N_2143,N_1134,N_607);
or U2144 (N_2144,N_1864,N_1412);
or U2145 (N_2145,N_687,N_916);
or U2146 (N_2146,N_1119,N_1466);
and U2147 (N_2147,N_1475,N_321);
xnor U2148 (N_2148,N_425,N_581);
and U2149 (N_2149,N_242,N_175);
or U2150 (N_2150,N_136,N_1609);
xor U2151 (N_2151,N_1868,N_128);
nor U2152 (N_2152,N_107,N_1046);
xor U2153 (N_2153,N_1333,N_1761);
and U2154 (N_2154,N_1213,N_1091);
nor U2155 (N_2155,N_859,N_152);
nor U2156 (N_2156,N_540,N_838);
and U2157 (N_2157,N_1055,N_1858);
nand U2158 (N_2158,N_72,N_1771);
nor U2159 (N_2159,N_1679,N_1002);
xnor U2160 (N_2160,N_542,N_1293);
nor U2161 (N_2161,N_1848,N_311);
nor U2162 (N_2162,N_502,N_664);
nor U2163 (N_2163,N_1807,N_1813);
nand U2164 (N_2164,N_1071,N_1115);
nand U2165 (N_2165,N_1984,N_1943);
or U2166 (N_2166,N_975,N_1103);
or U2167 (N_2167,N_200,N_524);
nand U2168 (N_2168,N_587,N_979);
nor U2169 (N_2169,N_1694,N_959);
or U2170 (N_2170,N_1832,N_1634);
xor U2171 (N_2171,N_1932,N_725);
xnor U2172 (N_2172,N_1816,N_1681);
and U2173 (N_2173,N_1044,N_1471);
nor U2174 (N_2174,N_1888,N_1169);
nand U2175 (N_2175,N_1312,N_1461);
and U2176 (N_2176,N_36,N_857);
nand U2177 (N_2177,N_285,N_861);
nor U2178 (N_2178,N_1208,N_545);
xor U2179 (N_2179,N_44,N_1776);
and U2180 (N_2180,N_738,N_468);
xnor U2181 (N_2181,N_1674,N_69);
and U2182 (N_2182,N_1770,N_267);
nand U2183 (N_2183,N_187,N_1833);
or U2184 (N_2184,N_106,N_1928);
nand U2185 (N_2185,N_804,N_964);
nand U2186 (N_2186,N_73,N_485);
xor U2187 (N_2187,N_479,N_1652);
nor U2188 (N_2188,N_430,N_130);
or U2189 (N_2189,N_138,N_1492);
or U2190 (N_2190,N_723,N_1248);
xor U2191 (N_2191,N_1716,N_1737);
xor U2192 (N_2192,N_42,N_788);
xnor U2193 (N_2193,N_1958,N_785);
or U2194 (N_2194,N_923,N_1083);
nand U2195 (N_2195,N_1498,N_659);
nand U2196 (N_2196,N_601,N_98);
nand U2197 (N_2197,N_1483,N_870);
nand U2198 (N_2198,N_1374,N_1715);
nand U2199 (N_2199,N_558,N_258);
xnor U2200 (N_2200,N_1250,N_183);
and U2201 (N_2201,N_1573,N_238);
nand U2202 (N_2202,N_1946,N_833);
nand U2203 (N_2203,N_34,N_1878);
nand U2204 (N_2204,N_917,N_1379);
or U2205 (N_2205,N_265,N_1905);
nor U2206 (N_2206,N_1361,N_446);
xor U2207 (N_2207,N_1194,N_1394);
nand U2208 (N_2208,N_832,N_765);
xor U2209 (N_2209,N_519,N_1459);
nor U2210 (N_2210,N_59,N_1100);
xor U2211 (N_2211,N_1017,N_1228);
xor U2212 (N_2212,N_649,N_1717);
and U2213 (N_2213,N_1356,N_619);
nand U2214 (N_2214,N_1844,N_149);
xnor U2215 (N_2215,N_1918,N_1903);
nand U2216 (N_2216,N_1525,N_1441);
or U2217 (N_2217,N_1703,N_611);
xor U2218 (N_2218,N_892,N_1722);
or U2219 (N_2219,N_218,N_1682);
nand U2220 (N_2220,N_1987,N_1101);
and U2221 (N_2221,N_1551,N_879);
nand U2222 (N_2222,N_716,N_1560);
nand U2223 (N_2223,N_170,N_65);
xor U2224 (N_2224,N_1920,N_33);
and U2225 (N_2225,N_874,N_1264);
xor U2226 (N_2226,N_435,N_1040);
nand U2227 (N_2227,N_223,N_427);
or U2228 (N_2228,N_1230,N_450);
or U2229 (N_2229,N_546,N_466);
or U2230 (N_2230,N_316,N_169);
xnor U2231 (N_2231,N_1023,N_461);
or U2232 (N_2232,N_147,N_277);
or U2233 (N_2233,N_405,N_1073);
nor U2234 (N_2234,N_1022,N_689);
nand U2235 (N_2235,N_731,N_815);
or U2236 (N_2236,N_55,N_1020);
xor U2237 (N_2237,N_1337,N_1786);
or U2238 (N_2238,N_982,N_196);
nor U2239 (N_2239,N_643,N_653);
or U2240 (N_2240,N_23,N_1014);
or U2241 (N_2241,N_795,N_1742);
xor U2242 (N_2242,N_332,N_625);
or U2243 (N_2243,N_836,N_721);
and U2244 (N_2244,N_1066,N_801);
xnor U2245 (N_2245,N_352,N_347);
nand U2246 (N_2246,N_1237,N_561);
nor U2247 (N_2247,N_1015,N_317);
xnor U2248 (N_2248,N_186,N_876);
xor U2249 (N_2249,N_399,N_1636);
or U2250 (N_2250,N_259,N_928);
nand U2251 (N_2251,N_602,N_1524);
nor U2252 (N_2252,N_1052,N_48);
nor U2253 (N_2253,N_1693,N_225);
and U2254 (N_2254,N_1400,N_1241);
xnor U2255 (N_2255,N_818,N_1117);
xnor U2256 (N_2256,N_1808,N_1425);
nor U2257 (N_2257,N_944,N_1926);
xor U2258 (N_2258,N_1760,N_1874);
and U2259 (N_2259,N_1390,N_1132);
and U2260 (N_2260,N_1539,N_307);
nand U2261 (N_2261,N_1974,N_410);
nor U2262 (N_2262,N_47,N_1319);
xor U2263 (N_2263,N_491,N_1646);
and U2264 (N_2264,N_436,N_29);
and U2265 (N_2265,N_657,N_1811);
nand U2266 (N_2266,N_528,N_253);
xnor U2267 (N_2267,N_274,N_1442);
xnor U2268 (N_2268,N_1377,N_1989);
nor U2269 (N_2269,N_1592,N_1885);
xnor U2270 (N_2270,N_1702,N_670);
nor U2271 (N_2271,N_516,N_1720);
xor U2272 (N_2272,N_1187,N_1673);
nor U2273 (N_2273,N_1950,N_1272);
nand U2274 (N_2274,N_555,N_1599);
xor U2275 (N_2275,N_620,N_622);
nor U2276 (N_2276,N_1528,N_527);
and U2277 (N_2277,N_671,N_1155);
xnor U2278 (N_2278,N_1426,N_981);
and U2279 (N_2279,N_1641,N_1407);
xor U2280 (N_2280,N_557,N_178);
xor U2281 (N_2281,N_447,N_1111);
and U2282 (N_2282,N_1108,N_1684);
nand U2283 (N_2283,N_388,N_148);
or U2284 (N_2284,N_1724,N_1509);
nor U2285 (N_2285,N_1260,N_214);
and U2286 (N_2286,N_88,N_57);
or U2287 (N_2287,N_629,N_1516);
or U2288 (N_2288,N_448,N_1163);
xnor U2289 (N_2289,N_908,N_883);
and U2290 (N_2290,N_1156,N_1077);
nor U2291 (N_2291,N_762,N_881);
xor U2292 (N_2292,N_496,N_967);
and U2293 (N_2293,N_251,N_889);
xor U2294 (N_2294,N_1661,N_1150);
nand U2295 (N_2295,N_735,N_1178);
or U2296 (N_2296,N_1439,N_925);
nor U2297 (N_2297,N_828,N_1467);
or U2298 (N_2298,N_1389,N_1581);
xor U2299 (N_2299,N_699,N_313);
nand U2300 (N_2300,N_550,N_453);
nor U2301 (N_2301,N_493,N_244);
or U2302 (N_2302,N_1588,N_797);
or U2303 (N_2303,N_1519,N_1727);
and U2304 (N_2304,N_1359,N_1220);
xor U2305 (N_2305,N_972,N_1606);
nand U2306 (N_2306,N_1654,N_1049);
xor U2307 (N_2307,N_656,N_1262);
nand U2308 (N_2308,N_547,N_640);
and U2309 (N_2309,N_324,N_1207);
or U2310 (N_2310,N_193,N_1346);
nor U2311 (N_2311,N_953,N_31);
nor U2312 (N_2312,N_93,N_1602);
nand U2313 (N_2313,N_1386,N_1303);
xnor U2314 (N_2314,N_1050,N_1500);
nor U2315 (N_2315,N_1675,N_526);
and U2316 (N_2316,N_1470,N_685);
and U2317 (N_2317,N_1243,N_963);
or U2318 (N_2318,N_490,N_1153);
or U2319 (N_2319,N_568,N_841);
xnor U2320 (N_2320,N_467,N_566);
or U2321 (N_2321,N_1183,N_1697);
xor U2322 (N_2322,N_1021,N_684);
nor U2323 (N_2323,N_284,N_269);
and U2324 (N_2324,N_191,N_1170);
and U2325 (N_2325,N_1719,N_146);
nand U2326 (N_2326,N_1124,N_1095);
and U2327 (N_2327,N_30,N_932);
and U2328 (N_2328,N_829,N_965);
and U2329 (N_2329,N_488,N_1372);
and U2330 (N_2330,N_1503,N_693);
nand U2331 (N_2331,N_291,N_350);
nor U2332 (N_2332,N_748,N_369);
xor U2333 (N_2333,N_1841,N_1924);
and U2334 (N_2334,N_1904,N_1755);
and U2335 (N_2335,N_434,N_1076);
xor U2336 (N_2336,N_184,N_991);
nand U2337 (N_2337,N_1199,N_698);
nand U2338 (N_2338,N_318,N_344);
nand U2339 (N_2339,N_514,N_1476);
and U2340 (N_2340,N_503,N_115);
nand U2341 (N_2341,N_1909,N_1849);
nor U2342 (N_2342,N_577,N_1037);
nand U2343 (N_2343,N_1743,N_887);
or U2344 (N_2344,N_1738,N_1799);
and U2345 (N_2345,N_947,N_1773);
nand U2346 (N_2346,N_1211,N_1570);
or U2347 (N_2347,N_432,N_771);
and U2348 (N_2348,N_1517,N_996);
xnor U2349 (N_2349,N_1666,N_1752);
or U2350 (N_2350,N_1565,N_260);
nor U2351 (N_2351,N_216,N_43);
or U2352 (N_2352,N_1283,N_770);
xor U2353 (N_2353,N_117,N_929);
and U2354 (N_2354,N_759,N_203);
or U2355 (N_2355,N_1942,N_1907);
xor U2356 (N_2356,N_1270,N_1753);
and U2357 (N_2357,N_1473,N_173);
nand U2358 (N_2358,N_1826,N_1512);
and U2359 (N_2359,N_732,N_532);
or U2360 (N_2360,N_740,N_256);
and U2361 (N_2361,N_623,N_382);
xor U2362 (N_2362,N_1791,N_384);
or U2363 (N_2363,N_116,N_408);
xnor U2364 (N_2364,N_808,N_295);
xnor U2365 (N_2365,N_465,N_1129);
xor U2366 (N_2366,N_411,N_704);
or U2367 (N_2367,N_380,N_275);
or U2368 (N_2368,N_1869,N_749);
and U2369 (N_2369,N_153,N_896);
nor U2370 (N_2370,N_246,N_1616);
nor U2371 (N_2371,N_521,N_1756);
xor U2372 (N_2372,N_1741,N_1623);
and U2373 (N_2373,N_1061,N_579);
xnor U2374 (N_2374,N_1709,N_5);
and U2375 (N_2375,N_415,N_21);
nor U2376 (N_2376,N_1469,N_834);
xor U2377 (N_2377,N_938,N_915);
nor U2378 (N_2378,N_1162,N_94);
xnor U2379 (N_2379,N_376,N_639);
or U2380 (N_2380,N_1521,N_426);
nor U2381 (N_2381,N_1835,N_1484);
nor U2382 (N_2382,N_615,N_755);
xnor U2383 (N_2383,N_1886,N_945);
and U2384 (N_2384,N_574,N_652);
nand U2385 (N_2385,N_144,N_1026);
xor U2386 (N_2386,N_1838,N_1508);
nand U2387 (N_2387,N_1547,N_359);
nor U2388 (N_2388,N_1301,N_660);
nand U2389 (N_2389,N_76,N_142);
nand U2390 (N_2390,N_1582,N_91);
or U2391 (N_2391,N_1889,N_777);
or U2392 (N_2392,N_1068,N_1149);
and U2393 (N_2393,N_968,N_160);
nor U2394 (N_2394,N_912,N_682);
or U2395 (N_2395,N_1955,N_1004);
nand U2396 (N_2396,N_1142,N_97);
or U2397 (N_2397,N_1444,N_495);
nand U2398 (N_2398,N_609,N_1060);
nand U2399 (N_2399,N_1449,N_1605);
nand U2400 (N_2400,N_444,N_604);
nand U2401 (N_2401,N_41,N_407);
nor U2402 (N_2402,N_1128,N_1923);
nand U2403 (N_2403,N_882,N_1902);
or U2404 (N_2404,N_35,N_1563);
nor U2405 (N_2405,N_875,N_543);
nand U2406 (N_2406,N_286,N_27);
or U2407 (N_2407,N_1880,N_1733);
nand U2408 (N_2408,N_541,N_758);
xor U2409 (N_2409,N_1914,N_417);
and U2410 (N_2410,N_821,N_50);
xnor U2411 (N_2411,N_279,N_1710);
nor U2412 (N_2412,N_1534,N_884);
xor U2413 (N_2413,N_1815,N_1310);
xnor U2414 (N_2414,N_1870,N_1919);
nor U2415 (N_2415,N_1854,N_994);
xor U2416 (N_2416,N_1268,N_1550);
nand U2417 (N_2417,N_1659,N_1277);
xor U2418 (N_2418,N_922,N_520);
or U2419 (N_2419,N_1670,N_81);
nor U2420 (N_2420,N_603,N_1225);
or U2421 (N_2421,N_624,N_962);
or U2422 (N_2422,N_853,N_1952);
or U2423 (N_2423,N_1726,N_353);
nand U2424 (N_2424,N_374,N_1018);
xnor U2425 (N_2425,N_686,N_1411);
xnor U2426 (N_2426,N_1478,N_737);
nand U2427 (N_2427,N_941,N_1341);
or U2428 (N_2428,N_414,N_1413);
nand U2429 (N_2429,N_366,N_1011);
nand U2430 (N_2430,N_995,N_378);
and U2431 (N_2431,N_1836,N_1488);
and U2432 (N_2432,N_1744,N_1687);
xor U2433 (N_2433,N_1445,N_264);
and U2434 (N_2434,N_954,N_1266);
xnor U2435 (N_2435,N_165,N_302);
and U2436 (N_2436,N_1348,N_1240);
and U2437 (N_2437,N_209,N_1893);
nand U2438 (N_2438,N_696,N_690);
nor U2439 (N_2439,N_594,N_1222);
and U2440 (N_2440,N_1613,N_87);
and U2441 (N_2441,N_1038,N_1448);
and U2442 (N_2442,N_606,N_825);
nor U2443 (N_2443,N_113,N_1586);
and U2444 (N_2444,N_984,N_381);
and U2445 (N_2445,N_507,N_1961);
and U2446 (N_2446,N_534,N_1174);
and U2447 (N_2447,N_301,N_406);
nor U2448 (N_2448,N_124,N_1642);
nor U2449 (N_2449,N_1604,N_1526);
nor U2450 (N_2450,N_1940,N_1567);
xnor U2451 (N_2451,N_1890,N_1347);
nor U2452 (N_2452,N_1351,N_851);
nand U2453 (N_2453,N_22,N_1287);
nand U2454 (N_2454,N_60,N_1438);
or U2455 (N_2455,N_1855,N_1649);
xor U2456 (N_2456,N_1707,N_1382);
or U2457 (N_2457,N_127,N_283);
xnor U2458 (N_2458,N_539,N_1653);
and U2459 (N_2459,N_1818,N_1280);
or U2460 (N_2460,N_1179,N_750);
xnor U2461 (N_2461,N_1549,N_1778);
nor U2462 (N_2462,N_1594,N_1891);
and U2463 (N_2463,N_1892,N_501);
xnor U2464 (N_2464,N_100,N_1392);
nor U2465 (N_2465,N_1276,N_787);
and U2466 (N_2466,N_1572,N_1010);
or U2467 (N_2467,N_1685,N_1857);
nor U2468 (N_2468,N_1354,N_395);
nand U2469 (N_2469,N_1899,N_1415);
and U2470 (N_2470,N_1949,N_1691);
or U2471 (N_2471,N_429,N_383);
or U2472 (N_2472,N_1418,N_918);
nor U2473 (N_2473,N_1837,N_1894);
nand U2474 (N_2474,N_1757,N_1840);
or U2475 (N_2475,N_1340,N_961);
nor U2476 (N_2476,N_1575,N_1219);
nor U2477 (N_2477,N_373,N_1479);
and U2478 (N_2478,N_10,N_586);
nor U2479 (N_2479,N_1054,N_680);
and U2480 (N_2480,N_1094,N_1645);
or U2481 (N_2481,N_631,N_776);
and U2482 (N_2482,N_1056,N_1154);
xor U2483 (N_2483,N_452,N_237);
or U2484 (N_2484,N_103,N_955);
and U2485 (N_2485,N_1239,N_1221);
and U2486 (N_2486,N_305,N_129);
nor U2487 (N_2487,N_1828,N_1081);
and U2488 (N_2488,N_143,N_1819);
or U2489 (N_2489,N_927,N_1802);
nor U2490 (N_2490,N_122,N_1427);
nand U2491 (N_2491,N_1431,N_1005);
xnor U2492 (N_2492,N_157,N_370);
or U2493 (N_2493,N_1099,N_2);
xnor U2494 (N_2494,N_617,N_70);
nor U2495 (N_2495,N_814,N_1764);
and U2496 (N_2496,N_621,N_997);
nor U2497 (N_2497,N_1862,N_569);
nand U2498 (N_2498,N_379,N_1798);
xor U2499 (N_2499,N_1165,N_971);
and U2500 (N_2500,N_1957,N_1352);
nand U2501 (N_2501,N_1734,N_319);
or U2502 (N_2502,N_1330,N_773);
nor U2503 (N_2503,N_1065,N_1618);
or U2504 (N_2504,N_613,N_1713);
nor U2505 (N_2505,N_3,N_958);
xnor U2506 (N_2506,N_270,N_351);
or U2507 (N_2507,N_1925,N_1295);
or U2508 (N_2508,N_811,N_1897);
xor U2509 (N_2509,N_562,N_1422);
and U2510 (N_2510,N_707,N_1140);
xor U2511 (N_2511,N_1784,N_1365);
or U2512 (N_2512,N_936,N_1587);
and U2513 (N_2513,N_1665,N_1024);
xor U2514 (N_2514,N_1406,N_1579);
and U2515 (N_2515,N_700,N_126);
xnor U2516 (N_2516,N_4,N_877);
and U2517 (N_2517,N_865,N_970);
or U2518 (N_2518,N_810,N_672);
or U2519 (N_2519,N_897,N_584);
or U2520 (N_2520,N_177,N_182);
xnor U2521 (N_2521,N_1553,N_241);
nand U2522 (N_2522,N_1589,N_1298);
and U2523 (N_2523,N_326,N_12);
and U2524 (N_2524,N_1809,N_1872);
nor U2525 (N_2525,N_25,N_1451);
or U2526 (N_2526,N_9,N_1396);
nand U2527 (N_2527,N_250,N_775);
or U2528 (N_2528,N_375,N_440);
or U2529 (N_2529,N_112,N_1197);
and U2530 (N_2530,N_688,N_768);
or U2531 (N_2531,N_1216,N_1177);
nor U2532 (N_2532,N_1215,N_1632);
and U2533 (N_2533,N_219,N_1663);
xnor U2534 (N_2534,N_1513,N_1751);
and U2535 (N_2535,N_389,N_800);
xor U2536 (N_2536,N_290,N_987);
or U2537 (N_2537,N_327,N_243);
nand U2538 (N_2538,N_1847,N_786);
xor U2539 (N_2539,N_1625,N_312);
nor U2540 (N_2540,N_1093,N_709);
nor U2541 (N_2541,N_717,N_1085);
nor U2542 (N_2542,N_1267,N_1097);
or U2543 (N_2543,N_403,N_1912);
nand U2544 (N_2544,N_197,N_1344);
xnor U2545 (N_2545,N_481,N_931);
xnor U2546 (N_2546,N_482,N_1789);
or U2547 (N_2547,N_1297,N_1496);
and U2548 (N_2548,N_204,N_66);
xor U2549 (N_2549,N_580,N_1088);
or U2550 (N_2550,N_220,N_1580);
and U2551 (N_2551,N_852,N_63);
xor U2552 (N_2552,N_141,N_571);
and U2553 (N_2553,N_343,N_1075);
nor U2554 (N_2554,N_1668,N_1986);
xor U2555 (N_2555,N_1992,N_767);
and U2556 (N_2556,N_1227,N_1689);
xnor U2557 (N_2557,N_1690,N_140);
nand U2558 (N_2558,N_839,N_743);
nand U2559 (N_2559,N_1045,N_729);
or U2560 (N_2560,N_207,N_948);
and U2561 (N_2561,N_635,N_120);
or U2562 (N_2562,N_1574,N_842);
xnor U2563 (N_2563,N_1332,N_505);
or U2564 (N_2564,N_590,N_869);
nand U2565 (N_2565,N_744,N_1324);
nor U2566 (N_2566,N_1245,N_1540);
or U2567 (N_2567,N_730,N_1188);
xor U2568 (N_2568,N_1936,N_1548);
nand U2569 (N_2569,N_424,N_651);
and U2570 (N_2570,N_486,N_1028);
xor U2571 (N_2571,N_504,N_1612);
or U2572 (N_2572,N_582,N_576);
or U2573 (N_2573,N_570,N_575);
xnor U2574 (N_2574,N_1704,N_1105);
xnor U2575 (N_2575,N_1403,N_525);
nand U2576 (N_2576,N_1195,N_537);
and U2577 (N_2577,N_413,N_392);
nand U2578 (N_2578,N_1235,N_386);
and U2579 (N_2579,N_346,N_92);
nor U2580 (N_2580,N_1048,N_1125);
or U2581 (N_2581,N_1723,N_900);
or U2582 (N_2582,N_1577,N_1146);
and U2583 (N_2583,N_1908,N_1996);
and U2584 (N_2584,N_1954,N_1883);
nor U2585 (N_2585,N_1285,N_1033);
nor U2586 (N_2586,N_1856,N_1274);
xnor U2587 (N_2587,N_1658,N_1258);
and U2588 (N_2588,N_32,N_1289);
nand U2589 (N_2589,N_1626,N_645);
and U2590 (N_2590,N_1008,N_816);
or U2591 (N_2591,N_1941,N_1985);
nor U2592 (N_2592,N_1536,N_1732);
and U2593 (N_2593,N_799,N_1916);
nor U2594 (N_2594,N_1793,N_1311);
nor U2595 (N_2595,N_506,N_1515);
or U2596 (N_2596,N_1931,N_1640);
xnor U2597 (N_2597,N_1135,N_1064);
nand U2598 (N_2598,N_630,N_533);
nand U2599 (N_2599,N_1031,N_137);
and U2600 (N_2600,N_1657,N_1939);
and U2601 (N_2601,N_805,N_1692);
xor U2602 (N_2602,N_80,N_1785);
nor U2603 (N_2603,N_1982,N_966);
or U2604 (N_2604,N_1895,N_1502);
and U2605 (N_2605,N_1205,N_210);
or U2606 (N_2606,N_1749,N_1631);
or U2607 (N_2607,N_1532,N_921);
xor U2608 (N_2608,N_1754,N_104);
nand U2609 (N_2609,N_194,N_1610);
or U2610 (N_2610,N_1316,N_1271);
nand U2611 (N_2611,N_798,N_1428);
and U2612 (N_2612,N_1109,N_1660);
nand U2613 (N_2613,N_53,N_589);
and U2614 (N_2614,N_306,N_1910);
nor U2615 (N_2615,N_367,N_470);
nor U2616 (N_2616,N_1058,N_368);
and U2617 (N_2617,N_423,N_320);
nor U2618 (N_2618,N_1810,N_1338);
or U2619 (N_2619,N_402,N_1877);
or U2620 (N_2620,N_431,N_1935);
or U2621 (N_2621,N_212,N_677);
xnor U2622 (N_2622,N_1564,N_1118);
nor U2623 (N_2623,N_1514,N_784);
or U2624 (N_2624,N_1971,N_474);
nor U2625 (N_2625,N_162,N_940);
xnor U2626 (N_2626,N_702,N_998);
xnor U2627 (N_2627,N_1462,N_1650);
and U2628 (N_2628,N_867,N_1615);
or U2629 (N_2629,N_1395,N_1947);
xor U2630 (N_2630,N_637,N_1299);
or U2631 (N_2631,N_276,N_692);
nor U2632 (N_2632,N_1401,N_812);
and U2633 (N_2633,N_325,N_412);
and U2634 (N_2634,N_1127,N_999);
xnor U2635 (N_2635,N_796,N_793);
nand U2636 (N_2636,N_1725,N_49);
nand U2637 (N_2637,N_293,N_159);
nand U2638 (N_2638,N_1440,N_1369);
nor U2639 (N_2639,N_185,N_1676);
or U2640 (N_2640,N_1794,N_1130);
or U2641 (N_2641,N_1434,N_1173);
nor U2642 (N_2642,N_1792,N_1968);
or U2643 (N_2643,N_83,N_1226);
or U2644 (N_2644,N_950,N_756);
nor U2645 (N_2645,N_1090,N_1139);
xnor U2646 (N_2646,N_1465,N_681);
nor U2647 (N_2647,N_96,N_1331);
and U2648 (N_2648,N_1036,N_74);
or U2649 (N_2649,N_633,N_980);
nand U2650 (N_2650,N_433,N_1988);
nand U2651 (N_2651,N_1309,N_1597);
xor U2652 (N_2652,N_1353,N_1543);
nand U2653 (N_2653,N_401,N_390);
nand U2654 (N_2654,N_1092,N_1677);
nand U2655 (N_2655,N_1911,N_1554);
xnor U2656 (N_2656,N_1621,N_217);
and U2657 (N_2657,N_983,N_150);
and U2658 (N_2658,N_1432,N_1797);
nor U2659 (N_2659,N_1399,N_1261);
nor U2660 (N_2660,N_1945,N_1366);
and U2661 (N_2661,N_1098,N_1729);
xor U2662 (N_2662,N_1647,N_858);
or U2663 (N_2663,N_674,N_1292);
or U2664 (N_2664,N_1318,N_1371);
and U2665 (N_2665,N_1160,N_583);
xor U2666 (N_2666,N_480,N_913);
or U2667 (N_2667,N_1062,N_232);
or U2668 (N_2668,N_1962,N_1039);
or U2669 (N_2669,N_46,N_1203);
nor U2670 (N_2670,N_573,N_722);
and U2671 (N_2671,N_1994,N_992);
xnor U2672 (N_2672,N_1545,N_695);
or U2673 (N_2673,N_937,N_844);
nand U2674 (N_2674,N_907,N_763);
nor U2675 (N_2675,N_1555,N_239);
and U2676 (N_2676,N_1494,N_885);
or U2677 (N_2677,N_315,N_1350);
nand U2678 (N_2678,N_778,N_1384);
or U2679 (N_2679,N_263,N_920);
xor U2680 (N_2680,N_648,N_939);
nand U2681 (N_2681,N_1879,N_16);
or U2682 (N_2682,N_1495,N_1566);
or U2683 (N_2683,N_1558,N_18);
xor U2684 (N_2684,N_308,N_309);
xor U2685 (N_2685,N_348,N_1468);
and U2686 (N_2686,N_1161,N_1067);
xnor U2687 (N_2687,N_701,N_271);
nand U2688 (N_2688,N_878,N_1137);
or U2689 (N_2689,N_362,N_614);
or U2690 (N_2690,N_1387,N_1531);
xor U2691 (N_2691,N_1447,N_1746);
xor U2692 (N_2692,N_105,N_298);
nand U2693 (N_2693,N_1965,N_760);
nand U2694 (N_2694,N_303,N_719);
and U2695 (N_2695,N_1882,N_1779);
and U2696 (N_2696,N_1113,N_1680);
nand U2697 (N_2697,N_281,N_1232);
or U2698 (N_2698,N_960,N_171);
nor U2699 (N_2699,N_1210,N_262);
and U2700 (N_2700,N_1414,N_428);
or U2701 (N_2701,N_416,N_957);
xnor U2702 (N_2702,N_1678,N_199);
nor U2703 (N_2703,N_441,N_632);
xnor U2704 (N_2704,N_400,N_1380);
nand U2705 (N_2705,N_294,N_942);
or U2706 (N_2706,N_1455,N_1079);
nor U2707 (N_2707,N_1559,N_1775);
and U2708 (N_2708,N_1107,N_1120);
or U2709 (N_2709,N_387,N_1635);
nor U2710 (N_2710,N_1504,N_1834);
xor U2711 (N_2711,N_245,N_823);
and U2712 (N_2712,N_898,N_1627);
nor U2713 (N_2713,N_419,N_1176);
xor U2714 (N_2714,N_1053,N_1385);
nand U2715 (N_2715,N_385,N_1373);
and U2716 (N_2716,N_202,N_1063);
or U2717 (N_2717,N_1765,N_1901);
nand U2718 (N_2718,N_304,N_1209);
nor U2719 (N_2719,N_1143,N_522);
xor U2720 (N_2720,N_1783,N_675);
nand U2721 (N_2721,N_830,N_1302);
xnor U2722 (N_2722,N_132,N_227);
xnor U2723 (N_2723,N_708,N_1148);
or U2724 (N_2724,N_1611,N_845);
xnor U2725 (N_2725,N_1736,N_456);
nand U2726 (N_2726,N_679,N_1740);
nor U2727 (N_2727,N_761,N_1288);
nand U2728 (N_2728,N_678,N_1185);
and U2729 (N_2729,N_167,N_1198);
xnor U2730 (N_2730,N_924,N_807);
or U2731 (N_2731,N_1001,N_563);
xnor U2732 (N_2732,N_1557,N_903);
nor U2733 (N_2733,N_1364,N_255);
nor U2734 (N_2734,N_1168,N_1242);
xor U2735 (N_2735,N_449,N_781);
nor U2736 (N_2736,N_422,N_248);
and U2737 (N_2737,N_1501,N_1806);
or U2738 (N_2738,N_254,N_339);
or U2739 (N_2739,N_1201,N_1383);
xnor U2740 (N_2740,N_1121,N_642);
and U2741 (N_2741,N_1922,N_421);
nor U2742 (N_2742,N_1978,N_236);
and U2743 (N_2743,N_71,N_135);
xnor U2744 (N_2744,N_864,N_101);
xnor U2745 (N_2745,N_1944,N_19);
nor U2746 (N_2746,N_1041,N_1698);
nor U2747 (N_2747,N_1421,N_1463);
or U2748 (N_2748,N_1546,N_572);
nor U2749 (N_2749,N_779,N_565);
nand U2750 (N_2750,N_1731,N_868);
and U2751 (N_2751,N_1999,N_1639);
xor U2752 (N_2752,N_1003,N_1917);
nand U2753 (N_2753,N_1667,N_1327);
xor U2754 (N_2754,N_110,N_1591);
and U2755 (N_2755,N_1419,N_1511);
nand U2756 (N_2756,N_1712,N_79);
nand U2757 (N_2757,N_1571,N_1070);
nand U2758 (N_2758,N_1278,N_1151);
xnor U2759 (N_2759,N_472,N_1990);
nand U2760 (N_2760,N_1643,N_1122);
or U2761 (N_2761,N_179,N_1368);
or U2762 (N_2762,N_1929,N_1795);
and U2763 (N_2763,N_1796,N_1051);
or U2764 (N_2764,N_1291,N_1206);
or U2765 (N_2765,N_1254,N_1158);
and U2766 (N_2766,N_1706,N_1934);
or U2767 (N_2767,N_904,N_145);
xnor U2768 (N_2768,N_1664,N_742);
and U2769 (N_2769,N_1304,N_1263);
and U2770 (N_2770,N_1029,N_644);
xnor U2771 (N_2771,N_58,N_1072);
or U2772 (N_2772,N_190,N_1480);
or U2773 (N_2773,N_1147,N_1530);
or U2774 (N_2774,N_1184,N_364);
or U2775 (N_2775,N_1402,N_310);
nor U2776 (N_2776,N_1763,N_1339);
or U2777 (N_2777,N_1969,N_323);
nand U2778 (N_2778,N_1043,N_1556);
or U2779 (N_2779,N_1322,N_1824);
or U2780 (N_2780,N_1000,N_508);
or U2781 (N_2781,N_500,N_1086);
xnor U2782 (N_2782,N_363,N_67);
nor U2783 (N_2783,N_1326,N_1186);
nand U2784 (N_2784,N_17,N_757);
xor U2785 (N_2785,N_1696,N_82);
xor U2786 (N_2786,N_1182,N_1967);
or U2787 (N_2787,N_1497,N_826);
or U2788 (N_2788,N_906,N_266);
and U2789 (N_2789,N_28,N_443);
nor U2790 (N_2790,N_1212,N_792);
or U2791 (N_2791,N_1656,N_694);
xnor U2792 (N_2792,N_1863,N_439);
or U2793 (N_2793,N_1410,N_498);
xor U2794 (N_2794,N_1648,N_213);
xor U2795 (N_2795,N_1921,N_654);
and U2796 (N_2796,N_934,N_726);
nand U2797 (N_2797,N_52,N_1489);
and U2798 (N_2798,N_1172,N_1523);
nor U2799 (N_2799,N_1800,N_1437);
nand U2800 (N_2800,N_638,N_899);
xor U2801 (N_2801,N_813,N_894);
and U2802 (N_2802,N_1747,N_341);
nor U2803 (N_2803,N_1204,N_1453);
and U2804 (N_2804,N_1981,N_372);
nor U2805 (N_2805,N_158,N_1252);
or U2806 (N_2806,N_1420,N_288);
or U2807 (N_2807,N_1306,N_1009);
nor U2808 (N_2808,N_734,N_1535);
nand U2809 (N_2809,N_1308,N_1608);
nand U2810 (N_2810,N_774,N_1181);
nand U2811 (N_2811,N_154,N_949);
xnor U2812 (N_2812,N_1450,N_1669);
xnor U2813 (N_2813,N_1533,N_599);
nor U2814 (N_2814,N_676,N_1012);
and U2815 (N_2815,N_1342,N_40);
xnor U2816 (N_2816,N_206,N_605);
nor U2817 (N_2817,N_224,N_1481);
and U2818 (N_2818,N_77,N_1454);
or U2819 (N_2819,N_499,N_616);
nor U2820 (N_2820,N_1482,N_1251);
or U2821 (N_2821,N_1144,N_221);
or U2822 (N_2822,N_24,N_930);
nor U2823 (N_2823,N_872,N_727);
xnor U2824 (N_2824,N_90,N_1233);
and U2825 (N_2825,N_835,N_710);
or U2826 (N_2826,N_1820,N_296);
xnor U2827 (N_2827,N_1180,N_1522);
nor U2828 (N_2828,N_1614,N_168);
nor U2829 (N_2829,N_1804,N_1404);
or U2830 (N_2830,N_1781,N_741);
or U2831 (N_2831,N_1443,N_554);
and U2832 (N_2832,N_478,N_1265);
nand U2833 (N_2833,N_910,N_349);
nand U2834 (N_2834,N_1777,N_85);
and U2835 (N_2835,N_1603,N_1822);
or U2836 (N_2836,N_1096,N_497);
nand U2837 (N_2837,N_1472,N_791);
nand U2838 (N_2838,N_1975,N_926);
nand U2839 (N_2839,N_1538,N_15);
nor U2840 (N_2840,N_1595,N_1537);
nand U2841 (N_2841,N_1505,N_1294);
nand U2842 (N_2842,N_549,N_1506);
and U2843 (N_2843,N_292,N_1409);
nand U2844 (N_2844,N_974,N_1850);
nand U2845 (N_2845,N_1259,N_300);
nand U2846 (N_2846,N_463,N_819);
and U2847 (N_2847,N_180,N_588);
nand U2848 (N_2848,N_1875,N_1948);
and U2849 (N_2849,N_1600,N_751);
or U2850 (N_2850,N_1430,N_1398);
nand U2851 (N_2851,N_1851,N_469);
and U2852 (N_2852,N_99,N_1257);
and U2853 (N_2853,N_578,N_1313);
xor U2854 (N_2854,N_1662,N_1282);
nand U2855 (N_2855,N_1803,N_1772);
or U2856 (N_2856,N_314,N_1672);
nand U2857 (N_2857,N_718,N_703);
nand U2858 (N_2858,N_1328,N_1074);
or U2859 (N_2859,N_393,N_1349);
and U2860 (N_2860,N_831,N_1671);
or U2861 (N_2861,N_628,N_1253);
nand U2862 (N_2862,N_1446,N_1541);
and U2863 (N_2863,N_1814,N_1728);
xnor U2864 (N_2864,N_1758,N_330);
xnor U2865 (N_2865,N_1637,N_11);
nand U2866 (N_2866,N_673,N_335);
or U2867 (N_2867,N_849,N_397);
and U2868 (N_2868,N_720,N_163);
and U2869 (N_2869,N_475,N_329);
nor U2870 (N_2870,N_226,N_336);
and U2871 (N_2871,N_553,N_817);
nor U2872 (N_2872,N_951,N_1218);
and U2873 (N_2873,N_95,N_1852);
xor U2874 (N_2874,N_1584,N_978);
and U2875 (N_2875,N_1873,N_1790);
and U2876 (N_2876,N_1493,N_1255);
or U2877 (N_2877,N_1853,N_1370);
nand U2878 (N_2878,N_1718,N_655);
nor U2879 (N_2879,N_1006,N_1831);
and U2880 (N_2880,N_1305,N_1617);
xor U2881 (N_2881,N_856,N_1972);
xnor U2882 (N_2882,N_850,N_1628);
nand U2883 (N_2883,N_1552,N_552);
xnor U2884 (N_2884,N_739,N_1585);
xor U2885 (N_2885,N_459,N_119);
xnor U2886 (N_2886,N_669,N_1300);
xor U2887 (N_2887,N_985,N_156);
nor U2888 (N_2888,N_705,N_396);
and U2889 (N_2889,N_873,N_125);
or U2890 (N_2890,N_1486,N_783);
and U2891 (N_2891,N_342,N_1510);
xnor U2892 (N_2892,N_1166,N_164);
xor U2893 (N_2893,N_890,N_1345);
nor U2894 (N_2894,N_866,N_121);
nor U2895 (N_2895,N_1315,N_1069);
xor U2896 (N_2896,N_438,N_1598);
xnor U2897 (N_2897,N_1279,N_38);
nor U2898 (N_2898,N_706,N_1238);
nor U2899 (N_2899,N_943,N_1966);
nor U2900 (N_2900,N_111,N_551);
or U2901 (N_2901,N_1766,N_1686);
or U2902 (N_2902,N_728,N_1970);
or U2903 (N_2903,N_1823,N_1876);
nor U2904 (N_2904,N_544,N_1224);
and U2905 (N_2905,N_1633,N_661);
nor U2906 (N_2906,N_1812,N_989);
nand U2907 (N_2907,N_322,N_789);
or U2908 (N_2908,N_517,N_1843);
and U2909 (N_2909,N_1025,N_1745);
nand U2910 (N_2910,N_1953,N_333);
or U2911 (N_2911,N_404,N_445);
or U2912 (N_2912,N_1106,N_473);
or U2913 (N_2913,N_1629,N_746);
and U2914 (N_2914,N_772,N_513);
or U2915 (N_2915,N_1244,N_192);
and U2916 (N_2916,N_1829,N_1927);
nand U2917 (N_2917,N_442,N_977);
and U2918 (N_2918,N_1192,N_394);
xor U2919 (N_2919,N_1084,N_365);
and U2920 (N_2920,N_1739,N_1780);
nor U2921 (N_2921,N_1630,N_1956);
nand U2922 (N_2922,N_1991,N_1590);
nor U2923 (N_2923,N_1490,N_1491);
nor U2924 (N_2924,N_1200,N_1367);
and U2925 (N_2925,N_6,N_195);
or U2926 (N_2926,N_1059,N_1249);
or U2927 (N_2927,N_1126,N_820);
nand U2928 (N_2928,N_176,N_1477);
xor U2929 (N_2929,N_358,N_860);
and U2930 (N_2930,N_724,N_1507);
nor U2931 (N_2931,N_1884,N_1993);
and U2932 (N_2932,N_714,N_595);
xnor U2933 (N_2933,N_174,N_455);
xor U2934 (N_2934,N_1217,N_1016);
or U2935 (N_2935,N_946,N_1436);
xor U2936 (N_2936,N_827,N_1320);
xor U2937 (N_2937,N_14,N_1620);
and U2938 (N_2938,N_1397,N_1748);
nand U2939 (N_2939,N_1435,N_1141);
nand U2940 (N_2940,N_666,N_1275);
nand U2941 (N_2941,N_457,N_1202);
and U2942 (N_2942,N_289,N_593);
nor U2943 (N_2943,N_1624,N_1325);
xnor U2944 (N_2944,N_231,N_854);
nand U2945 (N_2945,N_1391,N_118);
or U2946 (N_2946,N_272,N_181);
or U2947 (N_2947,N_1995,N_1762);
or U2948 (N_2948,N_139,N_646);
or U2949 (N_2949,N_1190,N_1321);
and U2950 (N_2950,N_888,N_1229);
nand U2951 (N_2951,N_1231,N_766);
nor U2952 (N_2952,N_108,N_665);
nor U2953 (N_2953,N_451,N_1019);
xnor U2954 (N_2954,N_109,N_51);
and U2955 (N_2955,N_377,N_627);
or U2956 (N_2956,N_863,N_1714);
nand U2957 (N_2957,N_560,N_618);
and U2958 (N_2958,N_1314,N_1825);
xor U2959 (N_2959,N_166,N_1393);
or U2960 (N_2960,N_1866,N_356);
and U2961 (N_2961,N_733,N_1317);
xnor U2962 (N_2962,N_1013,N_215);
nand U2963 (N_2963,N_1915,N_596);
nor U2964 (N_2964,N_1651,N_1561);
nor U2965 (N_2965,N_973,N_464);
nand U2966 (N_2966,N_1578,N_1683);
nor U2967 (N_2967,N_1034,N_75);
and U2968 (N_2968,N_1171,N_1619);
and U2969 (N_2969,N_969,N_45);
or U2970 (N_2970,N_667,N_1191);
nor U2971 (N_2971,N_454,N_988);
nor U2972 (N_2972,N_893,N_1452);
and U2973 (N_2973,N_902,N_151);
nand U2974 (N_2974,N_612,N_68);
xnor U2975 (N_2975,N_855,N_1933);
and U2976 (N_2976,N_172,N_189);
xnor U2977 (N_2977,N_1246,N_234);
nand U2978 (N_2978,N_208,N_1977);
xor U2979 (N_2979,N_483,N_54);
nand U2980 (N_2980,N_911,N_39);
xor U2981 (N_2981,N_188,N_89);
xor U2982 (N_2982,N_494,N_515);
nor U2983 (N_2983,N_1423,N_1376);
or U2984 (N_2984,N_1499,N_1290);
xor U2985 (N_2985,N_886,N_155);
xor U2986 (N_2986,N_420,N_1601);
nor U2987 (N_2987,N_608,N_1787);
xor U2988 (N_2988,N_1343,N_477);
or U2989 (N_2989,N_752,N_489);
xnor U2990 (N_2990,N_460,N_134);
and U2991 (N_2991,N_1157,N_1136);
nor U2992 (N_2992,N_462,N_847);
and U2993 (N_2993,N_1542,N_1152);
or U2994 (N_2994,N_591,N_1644);
nor U2995 (N_2995,N_1145,N_1114);
xor U2996 (N_2996,N_0,N_824);
nor U2997 (N_2997,N_1906,N_1408);
nand U2998 (N_2998,N_222,N_848);
xor U2999 (N_2999,N_1335,N_261);
nor U3000 (N_3000,N_1657,N_1994);
nand U3001 (N_3001,N_17,N_1024);
and U3002 (N_3002,N_1828,N_47);
nor U3003 (N_3003,N_1432,N_1085);
nand U3004 (N_3004,N_4,N_1457);
xnor U3005 (N_3005,N_166,N_621);
nand U3006 (N_3006,N_1345,N_486);
or U3007 (N_3007,N_1901,N_403);
nand U3008 (N_3008,N_1907,N_1649);
and U3009 (N_3009,N_1768,N_1772);
and U3010 (N_3010,N_1625,N_726);
nor U3011 (N_3011,N_1687,N_1332);
and U3012 (N_3012,N_47,N_247);
or U3013 (N_3013,N_416,N_1524);
or U3014 (N_3014,N_376,N_1640);
or U3015 (N_3015,N_940,N_1842);
and U3016 (N_3016,N_635,N_1380);
nand U3017 (N_3017,N_1334,N_285);
or U3018 (N_3018,N_1023,N_1071);
xor U3019 (N_3019,N_1527,N_625);
and U3020 (N_3020,N_594,N_534);
nor U3021 (N_3021,N_721,N_904);
and U3022 (N_3022,N_1206,N_1578);
nand U3023 (N_3023,N_447,N_274);
nand U3024 (N_3024,N_1650,N_1946);
and U3025 (N_3025,N_207,N_1873);
or U3026 (N_3026,N_24,N_1619);
nand U3027 (N_3027,N_856,N_251);
nand U3028 (N_3028,N_859,N_366);
or U3029 (N_3029,N_907,N_512);
xor U3030 (N_3030,N_1914,N_1932);
xnor U3031 (N_3031,N_1238,N_167);
nand U3032 (N_3032,N_1068,N_1837);
nor U3033 (N_3033,N_1845,N_1349);
nor U3034 (N_3034,N_221,N_1788);
nor U3035 (N_3035,N_26,N_1723);
nand U3036 (N_3036,N_27,N_1435);
or U3037 (N_3037,N_962,N_1541);
and U3038 (N_3038,N_1922,N_15);
nand U3039 (N_3039,N_29,N_918);
nor U3040 (N_3040,N_1499,N_1410);
nor U3041 (N_3041,N_1789,N_171);
and U3042 (N_3042,N_1376,N_354);
nand U3043 (N_3043,N_297,N_789);
nor U3044 (N_3044,N_365,N_1411);
nor U3045 (N_3045,N_972,N_1435);
or U3046 (N_3046,N_1439,N_377);
or U3047 (N_3047,N_1796,N_1889);
nand U3048 (N_3048,N_1434,N_385);
and U3049 (N_3049,N_1789,N_974);
xor U3050 (N_3050,N_718,N_752);
nand U3051 (N_3051,N_991,N_1003);
nor U3052 (N_3052,N_1256,N_150);
nand U3053 (N_3053,N_1322,N_1044);
nor U3054 (N_3054,N_777,N_1699);
xor U3055 (N_3055,N_1229,N_1440);
xnor U3056 (N_3056,N_1789,N_699);
nor U3057 (N_3057,N_54,N_768);
nor U3058 (N_3058,N_314,N_80);
nand U3059 (N_3059,N_1048,N_1945);
or U3060 (N_3060,N_480,N_1407);
or U3061 (N_3061,N_1430,N_30);
or U3062 (N_3062,N_1524,N_398);
or U3063 (N_3063,N_131,N_1262);
and U3064 (N_3064,N_1119,N_1830);
or U3065 (N_3065,N_762,N_1279);
and U3066 (N_3066,N_707,N_1296);
or U3067 (N_3067,N_61,N_493);
and U3068 (N_3068,N_246,N_823);
or U3069 (N_3069,N_134,N_262);
and U3070 (N_3070,N_1641,N_476);
nand U3071 (N_3071,N_523,N_1617);
nor U3072 (N_3072,N_1435,N_1644);
and U3073 (N_3073,N_1260,N_363);
and U3074 (N_3074,N_723,N_14);
xor U3075 (N_3075,N_230,N_333);
nand U3076 (N_3076,N_1288,N_1521);
nand U3077 (N_3077,N_1564,N_315);
xor U3078 (N_3078,N_1885,N_517);
and U3079 (N_3079,N_684,N_823);
or U3080 (N_3080,N_1197,N_1816);
xnor U3081 (N_3081,N_883,N_919);
and U3082 (N_3082,N_188,N_1114);
and U3083 (N_3083,N_798,N_1960);
xnor U3084 (N_3084,N_551,N_749);
and U3085 (N_3085,N_730,N_1580);
nor U3086 (N_3086,N_654,N_392);
nand U3087 (N_3087,N_1739,N_678);
and U3088 (N_3088,N_688,N_1721);
or U3089 (N_3089,N_380,N_924);
and U3090 (N_3090,N_322,N_621);
xnor U3091 (N_3091,N_62,N_418);
xnor U3092 (N_3092,N_895,N_1008);
nand U3093 (N_3093,N_527,N_1680);
xor U3094 (N_3094,N_15,N_583);
nor U3095 (N_3095,N_675,N_612);
xnor U3096 (N_3096,N_658,N_81);
nand U3097 (N_3097,N_342,N_321);
nand U3098 (N_3098,N_1395,N_713);
xnor U3099 (N_3099,N_952,N_449);
xor U3100 (N_3100,N_1692,N_450);
nor U3101 (N_3101,N_841,N_623);
xor U3102 (N_3102,N_1946,N_1980);
xor U3103 (N_3103,N_1548,N_12);
nor U3104 (N_3104,N_1671,N_1150);
nor U3105 (N_3105,N_1338,N_1001);
nor U3106 (N_3106,N_6,N_1092);
nor U3107 (N_3107,N_1713,N_527);
and U3108 (N_3108,N_909,N_218);
and U3109 (N_3109,N_1188,N_574);
nor U3110 (N_3110,N_269,N_31);
nor U3111 (N_3111,N_1284,N_44);
and U3112 (N_3112,N_648,N_1307);
nor U3113 (N_3113,N_1519,N_1779);
or U3114 (N_3114,N_1233,N_1619);
and U3115 (N_3115,N_1723,N_304);
nand U3116 (N_3116,N_1548,N_1094);
xor U3117 (N_3117,N_461,N_1411);
nand U3118 (N_3118,N_1325,N_1925);
and U3119 (N_3119,N_982,N_124);
nand U3120 (N_3120,N_1932,N_977);
or U3121 (N_3121,N_1659,N_1604);
or U3122 (N_3122,N_405,N_756);
xnor U3123 (N_3123,N_968,N_381);
nand U3124 (N_3124,N_1814,N_756);
or U3125 (N_3125,N_1472,N_785);
nor U3126 (N_3126,N_714,N_905);
nor U3127 (N_3127,N_1414,N_517);
xor U3128 (N_3128,N_240,N_141);
nand U3129 (N_3129,N_1040,N_151);
or U3130 (N_3130,N_1958,N_691);
nor U3131 (N_3131,N_1860,N_1197);
nand U3132 (N_3132,N_1106,N_348);
or U3133 (N_3133,N_1475,N_1403);
xnor U3134 (N_3134,N_1838,N_1668);
xnor U3135 (N_3135,N_1139,N_1202);
or U3136 (N_3136,N_1372,N_1894);
and U3137 (N_3137,N_1528,N_639);
or U3138 (N_3138,N_30,N_608);
and U3139 (N_3139,N_258,N_733);
nor U3140 (N_3140,N_1256,N_184);
or U3141 (N_3141,N_1808,N_624);
or U3142 (N_3142,N_682,N_1032);
and U3143 (N_3143,N_450,N_659);
xor U3144 (N_3144,N_1455,N_644);
nor U3145 (N_3145,N_1393,N_1873);
xnor U3146 (N_3146,N_1185,N_1482);
nor U3147 (N_3147,N_1965,N_250);
nand U3148 (N_3148,N_710,N_1508);
xnor U3149 (N_3149,N_1256,N_1108);
or U3150 (N_3150,N_164,N_335);
nand U3151 (N_3151,N_203,N_1680);
nand U3152 (N_3152,N_835,N_239);
xor U3153 (N_3153,N_409,N_1059);
or U3154 (N_3154,N_1662,N_1542);
nor U3155 (N_3155,N_445,N_1634);
xnor U3156 (N_3156,N_1961,N_1809);
nor U3157 (N_3157,N_500,N_1833);
nor U3158 (N_3158,N_607,N_79);
nor U3159 (N_3159,N_1185,N_1188);
and U3160 (N_3160,N_1158,N_176);
xnor U3161 (N_3161,N_54,N_1172);
and U3162 (N_3162,N_1798,N_244);
xnor U3163 (N_3163,N_713,N_26);
xor U3164 (N_3164,N_1568,N_1286);
xnor U3165 (N_3165,N_1382,N_244);
or U3166 (N_3166,N_973,N_1782);
and U3167 (N_3167,N_1906,N_1920);
and U3168 (N_3168,N_107,N_1825);
xnor U3169 (N_3169,N_1652,N_607);
xnor U3170 (N_3170,N_506,N_1388);
or U3171 (N_3171,N_388,N_607);
xor U3172 (N_3172,N_1757,N_841);
nor U3173 (N_3173,N_1642,N_1773);
nand U3174 (N_3174,N_166,N_865);
or U3175 (N_3175,N_906,N_1810);
xor U3176 (N_3176,N_1959,N_286);
nand U3177 (N_3177,N_1279,N_1633);
nor U3178 (N_3178,N_1749,N_504);
nand U3179 (N_3179,N_1040,N_816);
and U3180 (N_3180,N_494,N_782);
xnor U3181 (N_3181,N_1875,N_404);
and U3182 (N_3182,N_1758,N_1130);
nand U3183 (N_3183,N_1815,N_1309);
and U3184 (N_3184,N_1705,N_709);
and U3185 (N_3185,N_1352,N_70);
nor U3186 (N_3186,N_919,N_655);
or U3187 (N_3187,N_781,N_1199);
nand U3188 (N_3188,N_1956,N_499);
and U3189 (N_3189,N_976,N_1016);
nor U3190 (N_3190,N_836,N_45);
and U3191 (N_3191,N_1003,N_1123);
xor U3192 (N_3192,N_943,N_1013);
xnor U3193 (N_3193,N_1085,N_1384);
nand U3194 (N_3194,N_422,N_1917);
nand U3195 (N_3195,N_231,N_1073);
xnor U3196 (N_3196,N_982,N_1528);
nor U3197 (N_3197,N_260,N_537);
or U3198 (N_3198,N_219,N_1547);
nor U3199 (N_3199,N_1049,N_728);
xnor U3200 (N_3200,N_240,N_1034);
xnor U3201 (N_3201,N_748,N_982);
nand U3202 (N_3202,N_1609,N_902);
or U3203 (N_3203,N_1024,N_773);
nor U3204 (N_3204,N_340,N_1252);
nand U3205 (N_3205,N_455,N_1323);
nand U3206 (N_3206,N_1237,N_960);
and U3207 (N_3207,N_1823,N_750);
and U3208 (N_3208,N_1086,N_440);
and U3209 (N_3209,N_413,N_989);
and U3210 (N_3210,N_1274,N_1478);
nor U3211 (N_3211,N_122,N_1101);
nor U3212 (N_3212,N_1625,N_118);
xor U3213 (N_3213,N_1805,N_515);
xor U3214 (N_3214,N_434,N_1913);
or U3215 (N_3215,N_564,N_257);
or U3216 (N_3216,N_1275,N_150);
nand U3217 (N_3217,N_910,N_1021);
xnor U3218 (N_3218,N_210,N_795);
nor U3219 (N_3219,N_807,N_1623);
xnor U3220 (N_3220,N_49,N_234);
and U3221 (N_3221,N_550,N_723);
xnor U3222 (N_3222,N_638,N_1065);
or U3223 (N_3223,N_1710,N_1129);
nand U3224 (N_3224,N_302,N_995);
nor U3225 (N_3225,N_1675,N_162);
or U3226 (N_3226,N_908,N_1569);
xor U3227 (N_3227,N_1265,N_1239);
and U3228 (N_3228,N_875,N_1912);
xor U3229 (N_3229,N_1069,N_629);
or U3230 (N_3230,N_459,N_1686);
nor U3231 (N_3231,N_1173,N_1274);
nor U3232 (N_3232,N_1382,N_1862);
nand U3233 (N_3233,N_1780,N_344);
nor U3234 (N_3234,N_1154,N_1540);
nand U3235 (N_3235,N_68,N_1387);
nor U3236 (N_3236,N_1526,N_1309);
or U3237 (N_3237,N_1977,N_1355);
nor U3238 (N_3238,N_1723,N_51);
and U3239 (N_3239,N_821,N_897);
nor U3240 (N_3240,N_971,N_873);
nor U3241 (N_3241,N_294,N_63);
nand U3242 (N_3242,N_1757,N_1143);
nor U3243 (N_3243,N_448,N_655);
or U3244 (N_3244,N_1173,N_1296);
nor U3245 (N_3245,N_1482,N_694);
nand U3246 (N_3246,N_897,N_404);
xnor U3247 (N_3247,N_667,N_1796);
xnor U3248 (N_3248,N_123,N_718);
and U3249 (N_3249,N_656,N_1623);
xnor U3250 (N_3250,N_1957,N_1602);
nor U3251 (N_3251,N_950,N_1624);
xor U3252 (N_3252,N_1083,N_277);
and U3253 (N_3253,N_1962,N_757);
nor U3254 (N_3254,N_1809,N_86);
xor U3255 (N_3255,N_549,N_528);
and U3256 (N_3256,N_248,N_1196);
nor U3257 (N_3257,N_844,N_1304);
xnor U3258 (N_3258,N_1590,N_702);
nor U3259 (N_3259,N_533,N_1924);
xnor U3260 (N_3260,N_1146,N_191);
nor U3261 (N_3261,N_1925,N_828);
and U3262 (N_3262,N_1739,N_394);
xnor U3263 (N_3263,N_1084,N_934);
nor U3264 (N_3264,N_1074,N_117);
or U3265 (N_3265,N_1954,N_612);
and U3266 (N_3266,N_1289,N_1058);
nor U3267 (N_3267,N_1305,N_1152);
nor U3268 (N_3268,N_1305,N_1521);
or U3269 (N_3269,N_1446,N_913);
or U3270 (N_3270,N_1432,N_1096);
and U3271 (N_3271,N_1412,N_972);
xor U3272 (N_3272,N_635,N_796);
xor U3273 (N_3273,N_519,N_613);
nand U3274 (N_3274,N_1952,N_211);
nor U3275 (N_3275,N_354,N_245);
or U3276 (N_3276,N_1541,N_198);
and U3277 (N_3277,N_1278,N_525);
and U3278 (N_3278,N_1920,N_1276);
and U3279 (N_3279,N_540,N_1852);
nor U3280 (N_3280,N_631,N_106);
and U3281 (N_3281,N_345,N_1839);
and U3282 (N_3282,N_626,N_1490);
or U3283 (N_3283,N_1349,N_640);
nand U3284 (N_3284,N_408,N_1543);
or U3285 (N_3285,N_1141,N_1212);
nand U3286 (N_3286,N_1115,N_1645);
nand U3287 (N_3287,N_4,N_660);
nand U3288 (N_3288,N_1626,N_1801);
nor U3289 (N_3289,N_1330,N_193);
xor U3290 (N_3290,N_666,N_1635);
or U3291 (N_3291,N_1804,N_853);
nor U3292 (N_3292,N_1362,N_897);
and U3293 (N_3293,N_37,N_338);
nor U3294 (N_3294,N_1100,N_1408);
and U3295 (N_3295,N_1691,N_413);
or U3296 (N_3296,N_491,N_344);
nor U3297 (N_3297,N_733,N_1016);
or U3298 (N_3298,N_957,N_60);
and U3299 (N_3299,N_925,N_174);
nand U3300 (N_3300,N_981,N_1349);
xor U3301 (N_3301,N_221,N_889);
or U3302 (N_3302,N_1127,N_666);
xnor U3303 (N_3303,N_1259,N_1083);
or U3304 (N_3304,N_267,N_1288);
nand U3305 (N_3305,N_1039,N_939);
nand U3306 (N_3306,N_1868,N_764);
or U3307 (N_3307,N_350,N_1365);
or U3308 (N_3308,N_976,N_1622);
xor U3309 (N_3309,N_1211,N_36);
xnor U3310 (N_3310,N_100,N_80);
nor U3311 (N_3311,N_102,N_1216);
or U3312 (N_3312,N_547,N_1897);
xor U3313 (N_3313,N_1212,N_1578);
and U3314 (N_3314,N_1825,N_490);
or U3315 (N_3315,N_1441,N_455);
and U3316 (N_3316,N_1868,N_1112);
nand U3317 (N_3317,N_51,N_44);
or U3318 (N_3318,N_417,N_943);
nand U3319 (N_3319,N_1652,N_739);
nor U3320 (N_3320,N_1834,N_227);
xnor U3321 (N_3321,N_1655,N_780);
nand U3322 (N_3322,N_118,N_1419);
nor U3323 (N_3323,N_1599,N_946);
nand U3324 (N_3324,N_1799,N_1141);
nor U3325 (N_3325,N_830,N_1739);
and U3326 (N_3326,N_107,N_263);
xnor U3327 (N_3327,N_1511,N_1350);
xor U3328 (N_3328,N_125,N_413);
nor U3329 (N_3329,N_1233,N_1643);
nor U3330 (N_3330,N_1680,N_1754);
nand U3331 (N_3331,N_665,N_1354);
nand U3332 (N_3332,N_411,N_1332);
xnor U3333 (N_3333,N_1455,N_1891);
or U3334 (N_3334,N_670,N_1423);
nand U3335 (N_3335,N_1438,N_824);
xnor U3336 (N_3336,N_246,N_1346);
nor U3337 (N_3337,N_992,N_931);
xor U3338 (N_3338,N_1613,N_1271);
nand U3339 (N_3339,N_619,N_844);
nand U3340 (N_3340,N_195,N_927);
or U3341 (N_3341,N_1756,N_1326);
xnor U3342 (N_3342,N_96,N_1926);
nor U3343 (N_3343,N_1604,N_346);
or U3344 (N_3344,N_1679,N_1048);
nand U3345 (N_3345,N_1309,N_774);
and U3346 (N_3346,N_1770,N_1793);
xnor U3347 (N_3347,N_1006,N_231);
or U3348 (N_3348,N_568,N_481);
or U3349 (N_3349,N_620,N_1590);
xor U3350 (N_3350,N_232,N_1252);
and U3351 (N_3351,N_1213,N_70);
and U3352 (N_3352,N_91,N_552);
nand U3353 (N_3353,N_1210,N_421);
and U3354 (N_3354,N_1538,N_1379);
and U3355 (N_3355,N_1464,N_1773);
and U3356 (N_3356,N_366,N_1717);
and U3357 (N_3357,N_982,N_881);
or U3358 (N_3358,N_882,N_1671);
or U3359 (N_3359,N_1625,N_729);
and U3360 (N_3360,N_1968,N_560);
nand U3361 (N_3361,N_231,N_1680);
or U3362 (N_3362,N_1313,N_260);
nand U3363 (N_3363,N_378,N_322);
and U3364 (N_3364,N_1334,N_903);
and U3365 (N_3365,N_1793,N_557);
nor U3366 (N_3366,N_835,N_1180);
nor U3367 (N_3367,N_1725,N_1673);
and U3368 (N_3368,N_981,N_729);
and U3369 (N_3369,N_1411,N_1426);
and U3370 (N_3370,N_755,N_224);
nand U3371 (N_3371,N_1867,N_958);
and U3372 (N_3372,N_1053,N_1187);
and U3373 (N_3373,N_1652,N_1392);
or U3374 (N_3374,N_1576,N_1004);
or U3375 (N_3375,N_1402,N_797);
nand U3376 (N_3376,N_1759,N_1417);
xnor U3377 (N_3377,N_1082,N_315);
nand U3378 (N_3378,N_1582,N_1883);
or U3379 (N_3379,N_435,N_1192);
nand U3380 (N_3380,N_347,N_302);
nor U3381 (N_3381,N_527,N_1118);
or U3382 (N_3382,N_1843,N_281);
or U3383 (N_3383,N_1621,N_1145);
xnor U3384 (N_3384,N_748,N_1484);
and U3385 (N_3385,N_1067,N_949);
xnor U3386 (N_3386,N_1760,N_582);
nor U3387 (N_3387,N_1498,N_892);
and U3388 (N_3388,N_1161,N_1275);
nand U3389 (N_3389,N_977,N_794);
and U3390 (N_3390,N_56,N_1094);
or U3391 (N_3391,N_523,N_1030);
xor U3392 (N_3392,N_1333,N_1090);
or U3393 (N_3393,N_1060,N_1137);
nand U3394 (N_3394,N_409,N_273);
nor U3395 (N_3395,N_770,N_299);
or U3396 (N_3396,N_375,N_280);
and U3397 (N_3397,N_1753,N_965);
and U3398 (N_3398,N_1103,N_756);
nor U3399 (N_3399,N_1699,N_1703);
nand U3400 (N_3400,N_883,N_1239);
xnor U3401 (N_3401,N_1397,N_834);
nand U3402 (N_3402,N_1109,N_1676);
or U3403 (N_3403,N_1691,N_1899);
nand U3404 (N_3404,N_1502,N_1400);
or U3405 (N_3405,N_1805,N_1216);
and U3406 (N_3406,N_58,N_304);
and U3407 (N_3407,N_598,N_1265);
nand U3408 (N_3408,N_1232,N_1481);
and U3409 (N_3409,N_1221,N_1691);
xor U3410 (N_3410,N_485,N_826);
nor U3411 (N_3411,N_1115,N_863);
nor U3412 (N_3412,N_870,N_1060);
nor U3413 (N_3413,N_1007,N_268);
nand U3414 (N_3414,N_1745,N_40);
and U3415 (N_3415,N_1872,N_72);
nand U3416 (N_3416,N_1726,N_731);
xor U3417 (N_3417,N_1724,N_1263);
or U3418 (N_3418,N_1327,N_211);
xor U3419 (N_3419,N_1318,N_1617);
nand U3420 (N_3420,N_1282,N_1331);
xnor U3421 (N_3421,N_1012,N_1752);
nor U3422 (N_3422,N_487,N_357);
nand U3423 (N_3423,N_1941,N_959);
nor U3424 (N_3424,N_887,N_152);
nand U3425 (N_3425,N_264,N_79);
or U3426 (N_3426,N_525,N_78);
and U3427 (N_3427,N_454,N_1489);
nand U3428 (N_3428,N_1296,N_1461);
xor U3429 (N_3429,N_1817,N_1585);
nor U3430 (N_3430,N_941,N_1707);
nand U3431 (N_3431,N_989,N_1385);
or U3432 (N_3432,N_59,N_910);
nand U3433 (N_3433,N_572,N_1032);
and U3434 (N_3434,N_336,N_1240);
or U3435 (N_3435,N_1000,N_537);
nand U3436 (N_3436,N_1002,N_308);
and U3437 (N_3437,N_1950,N_1265);
nand U3438 (N_3438,N_962,N_356);
or U3439 (N_3439,N_1227,N_1139);
or U3440 (N_3440,N_697,N_1004);
nand U3441 (N_3441,N_168,N_1845);
xnor U3442 (N_3442,N_1672,N_284);
or U3443 (N_3443,N_770,N_1525);
and U3444 (N_3444,N_1843,N_1948);
and U3445 (N_3445,N_716,N_435);
nor U3446 (N_3446,N_647,N_402);
xor U3447 (N_3447,N_987,N_47);
and U3448 (N_3448,N_1646,N_1440);
xor U3449 (N_3449,N_1409,N_6);
nand U3450 (N_3450,N_932,N_256);
nor U3451 (N_3451,N_971,N_1892);
or U3452 (N_3452,N_1147,N_434);
and U3453 (N_3453,N_1323,N_1081);
and U3454 (N_3454,N_240,N_1214);
and U3455 (N_3455,N_715,N_515);
xnor U3456 (N_3456,N_746,N_996);
nand U3457 (N_3457,N_1415,N_1149);
or U3458 (N_3458,N_1300,N_1475);
nor U3459 (N_3459,N_1241,N_1379);
xor U3460 (N_3460,N_1640,N_1139);
nor U3461 (N_3461,N_1857,N_1666);
xnor U3462 (N_3462,N_1722,N_224);
nor U3463 (N_3463,N_1978,N_1241);
xnor U3464 (N_3464,N_1002,N_426);
or U3465 (N_3465,N_502,N_100);
xor U3466 (N_3466,N_711,N_765);
nand U3467 (N_3467,N_319,N_661);
nand U3468 (N_3468,N_1230,N_1939);
or U3469 (N_3469,N_541,N_1231);
or U3470 (N_3470,N_114,N_681);
or U3471 (N_3471,N_678,N_1354);
xor U3472 (N_3472,N_1832,N_1833);
nand U3473 (N_3473,N_1527,N_1024);
nor U3474 (N_3474,N_1774,N_633);
or U3475 (N_3475,N_148,N_1770);
nor U3476 (N_3476,N_564,N_994);
nor U3477 (N_3477,N_910,N_1816);
nor U3478 (N_3478,N_709,N_381);
nand U3479 (N_3479,N_1271,N_245);
xor U3480 (N_3480,N_1121,N_978);
xnor U3481 (N_3481,N_190,N_287);
nor U3482 (N_3482,N_997,N_243);
or U3483 (N_3483,N_332,N_1138);
and U3484 (N_3484,N_1969,N_306);
or U3485 (N_3485,N_1013,N_187);
or U3486 (N_3486,N_1490,N_1703);
and U3487 (N_3487,N_1049,N_42);
or U3488 (N_3488,N_1997,N_745);
or U3489 (N_3489,N_486,N_788);
xnor U3490 (N_3490,N_251,N_1131);
nand U3491 (N_3491,N_615,N_1489);
nand U3492 (N_3492,N_440,N_1053);
nand U3493 (N_3493,N_323,N_826);
nor U3494 (N_3494,N_988,N_709);
and U3495 (N_3495,N_324,N_1214);
or U3496 (N_3496,N_1833,N_808);
and U3497 (N_3497,N_1298,N_1357);
xnor U3498 (N_3498,N_918,N_1681);
nor U3499 (N_3499,N_1808,N_1516);
nand U3500 (N_3500,N_928,N_38);
or U3501 (N_3501,N_1615,N_1819);
nor U3502 (N_3502,N_1713,N_824);
and U3503 (N_3503,N_1242,N_1503);
xnor U3504 (N_3504,N_1748,N_1173);
nand U3505 (N_3505,N_1265,N_1518);
and U3506 (N_3506,N_1513,N_872);
nor U3507 (N_3507,N_1054,N_484);
or U3508 (N_3508,N_692,N_1794);
nand U3509 (N_3509,N_805,N_712);
nand U3510 (N_3510,N_1289,N_911);
nand U3511 (N_3511,N_862,N_1555);
nor U3512 (N_3512,N_693,N_200);
or U3513 (N_3513,N_241,N_1259);
or U3514 (N_3514,N_1358,N_363);
nor U3515 (N_3515,N_1427,N_1302);
and U3516 (N_3516,N_511,N_1231);
or U3517 (N_3517,N_1094,N_428);
and U3518 (N_3518,N_1369,N_864);
and U3519 (N_3519,N_680,N_1206);
xnor U3520 (N_3520,N_51,N_1681);
nor U3521 (N_3521,N_725,N_1051);
or U3522 (N_3522,N_200,N_860);
or U3523 (N_3523,N_1131,N_882);
or U3524 (N_3524,N_1766,N_1938);
xor U3525 (N_3525,N_27,N_1963);
nand U3526 (N_3526,N_266,N_1561);
nor U3527 (N_3527,N_1503,N_71);
nor U3528 (N_3528,N_56,N_802);
nand U3529 (N_3529,N_1144,N_947);
and U3530 (N_3530,N_1713,N_1902);
nor U3531 (N_3531,N_949,N_1700);
nand U3532 (N_3532,N_991,N_1484);
or U3533 (N_3533,N_1021,N_524);
and U3534 (N_3534,N_452,N_1000);
or U3535 (N_3535,N_1459,N_1623);
or U3536 (N_3536,N_463,N_1205);
nor U3537 (N_3537,N_106,N_1628);
or U3538 (N_3538,N_780,N_1000);
xnor U3539 (N_3539,N_396,N_1148);
and U3540 (N_3540,N_1639,N_933);
nand U3541 (N_3541,N_841,N_1571);
and U3542 (N_3542,N_1749,N_1683);
xor U3543 (N_3543,N_156,N_1566);
nor U3544 (N_3544,N_199,N_1312);
nor U3545 (N_3545,N_172,N_550);
nand U3546 (N_3546,N_103,N_1214);
nand U3547 (N_3547,N_109,N_1502);
nand U3548 (N_3548,N_350,N_386);
xor U3549 (N_3549,N_1852,N_1382);
nand U3550 (N_3550,N_1312,N_627);
nand U3551 (N_3551,N_1891,N_1678);
xnor U3552 (N_3552,N_343,N_1211);
nand U3553 (N_3553,N_1757,N_242);
nor U3554 (N_3554,N_801,N_152);
nor U3555 (N_3555,N_1343,N_1321);
and U3556 (N_3556,N_1016,N_1234);
and U3557 (N_3557,N_948,N_166);
xnor U3558 (N_3558,N_1433,N_1703);
or U3559 (N_3559,N_501,N_1072);
or U3560 (N_3560,N_508,N_385);
nor U3561 (N_3561,N_1889,N_160);
nor U3562 (N_3562,N_1442,N_52);
nand U3563 (N_3563,N_182,N_1580);
nand U3564 (N_3564,N_289,N_1988);
xnor U3565 (N_3565,N_1002,N_427);
nand U3566 (N_3566,N_35,N_1353);
and U3567 (N_3567,N_1362,N_1271);
nor U3568 (N_3568,N_815,N_1733);
nand U3569 (N_3569,N_1117,N_676);
nor U3570 (N_3570,N_1961,N_588);
nand U3571 (N_3571,N_1847,N_1629);
nand U3572 (N_3572,N_1595,N_1381);
xnor U3573 (N_3573,N_1919,N_1811);
or U3574 (N_3574,N_867,N_1345);
nor U3575 (N_3575,N_1757,N_414);
or U3576 (N_3576,N_482,N_98);
or U3577 (N_3577,N_883,N_421);
nand U3578 (N_3578,N_1767,N_434);
nor U3579 (N_3579,N_1514,N_1374);
and U3580 (N_3580,N_1470,N_439);
nand U3581 (N_3581,N_965,N_449);
and U3582 (N_3582,N_1491,N_1039);
nor U3583 (N_3583,N_1847,N_1475);
or U3584 (N_3584,N_1429,N_1157);
and U3585 (N_3585,N_656,N_214);
or U3586 (N_3586,N_1930,N_1243);
nand U3587 (N_3587,N_1629,N_1682);
xnor U3588 (N_3588,N_296,N_207);
nor U3589 (N_3589,N_353,N_1067);
nand U3590 (N_3590,N_1917,N_1893);
and U3591 (N_3591,N_630,N_1265);
and U3592 (N_3592,N_1106,N_1067);
or U3593 (N_3593,N_1918,N_1776);
nand U3594 (N_3594,N_1013,N_1361);
nand U3595 (N_3595,N_1044,N_1809);
or U3596 (N_3596,N_430,N_901);
nor U3597 (N_3597,N_1101,N_1197);
nand U3598 (N_3598,N_1685,N_563);
and U3599 (N_3599,N_351,N_832);
and U3600 (N_3600,N_807,N_113);
and U3601 (N_3601,N_1299,N_802);
or U3602 (N_3602,N_1456,N_146);
xor U3603 (N_3603,N_18,N_698);
nand U3604 (N_3604,N_1917,N_983);
nand U3605 (N_3605,N_257,N_1135);
and U3606 (N_3606,N_1823,N_975);
nand U3607 (N_3607,N_1432,N_960);
nor U3608 (N_3608,N_163,N_548);
or U3609 (N_3609,N_170,N_487);
nand U3610 (N_3610,N_1587,N_692);
nor U3611 (N_3611,N_1759,N_1586);
or U3612 (N_3612,N_548,N_1404);
xor U3613 (N_3613,N_263,N_1946);
and U3614 (N_3614,N_207,N_1281);
nand U3615 (N_3615,N_1226,N_863);
or U3616 (N_3616,N_318,N_1656);
nand U3617 (N_3617,N_851,N_1972);
or U3618 (N_3618,N_57,N_373);
nor U3619 (N_3619,N_389,N_1891);
nor U3620 (N_3620,N_1243,N_1628);
and U3621 (N_3621,N_778,N_807);
nor U3622 (N_3622,N_654,N_1689);
nor U3623 (N_3623,N_1637,N_1148);
or U3624 (N_3624,N_1023,N_1902);
and U3625 (N_3625,N_1664,N_710);
and U3626 (N_3626,N_1489,N_358);
or U3627 (N_3627,N_1347,N_1560);
and U3628 (N_3628,N_1168,N_1968);
nand U3629 (N_3629,N_1272,N_1275);
or U3630 (N_3630,N_1857,N_1751);
or U3631 (N_3631,N_446,N_1803);
xor U3632 (N_3632,N_1656,N_680);
and U3633 (N_3633,N_1612,N_26);
nor U3634 (N_3634,N_20,N_1145);
or U3635 (N_3635,N_169,N_1485);
or U3636 (N_3636,N_16,N_1683);
nor U3637 (N_3637,N_452,N_509);
nor U3638 (N_3638,N_1845,N_1499);
nor U3639 (N_3639,N_399,N_1069);
or U3640 (N_3640,N_504,N_1458);
and U3641 (N_3641,N_914,N_481);
nand U3642 (N_3642,N_1065,N_1485);
and U3643 (N_3643,N_816,N_271);
or U3644 (N_3644,N_1580,N_1485);
xnor U3645 (N_3645,N_1826,N_331);
nor U3646 (N_3646,N_1137,N_982);
or U3647 (N_3647,N_1330,N_1143);
or U3648 (N_3648,N_280,N_1222);
or U3649 (N_3649,N_1940,N_928);
nor U3650 (N_3650,N_104,N_1694);
nand U3651 (N_3651,N_1929,N_683);
xor U3652 (N_3652,N_1265,N_523);
or U3653 (N_3653,N_1175,N_1629);
nand U3654 (N_3654,N_1505,N_459);
xor U3655 (N_3655,N_1959,N_39);
nand U3656 (N_3656,N_140,N_419);
and U3657 (N_3657,N_986,N_853);
nand U3658 (N_3658,N_1177,N_786);
nor U3659 (N_3659,N_804,N_1454);
nor U3660 (N_3660,N_230,N_1466);
xnor U3661 (N_3661,N_1097,N_446);
or U3662 (N_3662,N_269,N_527);
or U3663 (N_3663,N_936,N_434);
nor U3664 (N_3664,N_358,N_1717);
xor U3665 (N_3665,N_1432,N_1157);
or U3666 (N_3666,N_33,N_161);
nor U3667 (N_3667,N_442,N_1129);
nand U3668 (N_3668,N_1050,N_1083);
and U3669 (N_3669,N_562,N_566);
nand U3670 (N_3670,N_106,N_1839);
or U3671 (N_3671,N_733,N_1427);
or U3672 (N_3672,N_1766,N_762);
xnor U3673 (N_3673,N_1499,N_504);
and U3674 (N_3674,N_1305,N_1528);
nor U3675 (N_3675,N_1535,N_1736);
nor U3676 (N_3676,N_1242,N_1400);
nor U3677 (N_3677,N_1687,N_1185);
nand U3678 (N_3678,N_606,N_1337);
nand U3679 (N_3679,N_628,N_1370);
nor U3680 (N_3680,N_23,N_350);
nand U3681 (N_3681,N_152,N_751);
nor U3682 (N_3682,N_997,N_1821);
and U3683 (N_3683,N_257,N_549);
nand U3684 (N_3684,N_945,N_1066);
nand U3685 (N_3685,N_772,N_1974);
xor U3686 (N_3686,N_737,N_1950);
xnor U3687 (N_3687,N_1839,N_927);
xor U3688 (N_3688,N_1068,N_1859);
xnor U3689 (N_3689,N_1006,N_801);
or U3690 (N_3690,N_1057,N_1503);
xor U3691 (N_3691,N_143,N_1290);
nand U3692 (N_3692,N_534,N_369);
nand U3693 (N_3693,N_959,N_927);
nand U3694 (N_3694,N_620,N_1751);
nand U3695 (N_3695,N_350,N_1085);
and U3696 (N_3696,N_718,N_1346);
xor U3697 (N_3697,N_477,N_214);
and U3698 (N_3698,N_1006,N_905);
nand U3699 (N_3699,N_1362,N_1349);
or U3700 (N_3700,N_455,N_899);
nor U3701 (N_3701,N_625,N_1956);
xor U3702 (N_3702,N_220,N_1404);
xor U3703 (N_3703,N_695,N_487);
and U3704 (N_3704,N_1840,N_543);
nor U3705 (N_3705,N_1583,N_1617);
and U3706 (N_3706,N_1267,N_479);
or U3707 (N_3707,N_379,N_162);
and U3708 (N_3708,N_1230,N_513);
or U3709 (N_3709,N_401,N_555);
and U3710 (N_3710,N_204,N_1931);
or U3711 (N_3711,N_1951,N_932);
and U3712 (N_3712,N_380,N_930);
xor U3713 (N_3713,N_196,N_953);
and U3714 (N_3714,N_1193,N_668);
nand U3715 (N_3715,N_6,N_1528);
nand U3716 (N_3716,N_641,N_1287);
and U3717 (N_3717,N_773,N_1559);
nand U3718 (N_3718,N_1018,N_1047);
xnor U3719 (N_3719,N_274,N_474);
and U3720 (N_3720,N_463,N_1520);
xnor U3721 (N_3721,N_980,N_1743);
nand U3722 (N_3722,N_672,N_1755);
nand U3723 (N_3723,N_309,N_958);
nand U3724 (N_3724,N_1814,N_1196);
nor U3725 (N_3725,N_321,N_322);
nor U3726 (N_3726,N_1097,N_835);
xor U3727 (N_3727,N_617,N_191);
or U3728 (N_3728,N_582,N_732);
nor U3729 (N_3729,N_812,N_1446);
nor U3730 (N_3730,N_1285,N_325);
nor U3731 (N_3731,N_1662,N_102);
nand U3732 (N_3732,N_1604,N_1684);
or U3733 (N_3733,N_558,N_1788);
nor U3734 (N_3734,N_466,N_789);
and U3735 (N_3735,N_1904,N_823);
and U3736 (N_3736,N_1628,N_1693);
xnor U3737 (N_3737,N_1952,N_1203);
nor U3738 (N_3738,N_1418,N_1479);
nand U3739 (N_3739,N_1156,N_1280);
xor U3740 (N_3740,N_1502,N_1822);
and U3741 (N_3741,N_1971,N_1846);
nand U3742 (N_3742,N_1142,N_1199);
xnor U3743 (N_3743,N_1819,N_1480);
nor U3744 (N_3744,N_1589,N_1547);
or U3745 (N_3745,N_424,N_392);
nand U3746 (N_3746,N_1471,N_477);
or U3747 (N_3747,N_1300,N_1173);
nand U3748 (N_3748,N_1257,N_1374);
or U3749 (N_3749,N_211,N_445);
xnor U3750 (N_3750,N_445,N_332);
xor U3751 (N_3751,N_573,N_1894);
nor U3752 (N_3752,N_65,N_1168);
or U3753 (N_3753,N_870,N_1320);
xnor U3754 (N_3754,N_326,N_827);
and U3755 (N_3755,N_1271,N_1056);
and U3756 (N_3756,N_1461,N_1928);
xor U3757 (N_3757,N_1676,N_965);
nor U3758 (N_3758,N_1248,N_1670);
nand U3759 (N_3759,N_917,N_1180);
or U3760 (N_3760,N_1365,N_572);
nor U3761 (N_3761,N_1371,N_98);
nor U3762 (N_3762,N_1957,N_1014);
nor U3763 (N_3763,N_1258,N_692);
xnor U3764 (N_3764,N_799,N_711);
nand U3765 (N_3765,N_474,N_954);
and U3766 (N_3766,N_130,N_1653);
or U3767 (N_3767,N_37,N_182);
or U3768 (N_3768,N_1042,N_1809);
nand U3769 (N_3769,N_838,N_1024);
nand U3770 (N_3770,N_561,N_1825);
nor U3771 (N_3771,N_70,N_1865);
xor U3772 (N_3772,N_737,N_1932);
nor U3773 (N_3773,N_524,N_512);
and U3774 (N_3774,N_1058,N_1852);
and U3775 (N_3775,N_631,N_300);
xnor U3776 (N_3776,N_1034,N_220);
xnor U3777 (N_3777,N_158,N_1050);
nand U3778 (N_3778,N_1330,N_1050);
and U3779 (N_3779,N_1429,N_1796);
and U3780 (N_3780,N_175,N_1559);
or U3781 (N_3781,N_661,N_440);
and U3782 (N_3782,N_547,N_1304);
nor U3783 (N_3783,N_1208,N_1318);
xor U3784 (N_3784,N_193,N_1498);
nand U3785 (N_3785,N_1037,N_1861);
or U3786 (N_3786,N_1797,N_1014);
nand U3787 (N_3787,N_1069,N_1470);
or U3788 (N_3788,N_133,N_843);
nand U3789 (N_3789,N_415,N_1464);
or U3790 (N_3790,N_231,N_436);
xor U3791 (N_3791,N_260,N_993);
nand U3792 (N_3792,N_54,N_1326);
and U3793 (N_3793,N_724,N_508);
xnor U3794 (N_3794,N_1645,N_473);
xnor U3795 (N_3795,N_818,N_26);
nor U3796 (N_3796,N_1373,N_1642);
nand U3797 (N_3797,N_1645,N_1131);
or U3798 (N_3798,N_853,N_1486);
or U3799 (N_3799,N_1067,N_499);
nand U3800 (N_3800,N_444,N_965);
nor U3801 (N_3801,N_1943,N_1112);
xor U3802 (N_3802,N_731,N_1493);
or U3803 (N_3803,N_1519,N_7);
or U3804 (N_3804,N_1867,N_878);
nand U3805 (N_3805,N_476,N_1832);
or U3806 (N_3806,N_121,N_178);
nor U3807 (N_3807,N_1775,N_1793);
and U3808 (N_3808,N_1168,N_1767);
or U3809 (N_3809,N_749,N_1245);
or U3810 (N_3810,N_663,N_1585);
or U3811 (N_3811,N_1885,N_1663);
nor U3812 (N_3812,N_191,N_1523);
xnor U3813 (N_3813,N_1238,N_531);
and U3814 (N_3814,N_996,N_766);
xor U3815 (N_3815,N_714,N_1463);
and U3816 (N_3816,N_359,N_350);
nor U3817 (N_3817,N_387,N_1369);
nor U3818 (N_3818,N_631,N_1335);
xnor U3819 (N_3819,N_1496,N_1794);
or U3820 (N_3820,N_1772,N_1727);
and U3821 (N_3821,N_1607,N_1182);
nand U3822 (N_3822,N_1827,N_817);
xnor U3823 (N_3823,N_836,N_771);
and U3824 (N_3824,N_1326,N_1433);
xnor U3825 (N_3825,N_155,N_735);
xnor U3826 (N_3826,N_1133,N_1967);
xnor U3827 (N_3827,N_1379,N_386);
nor U3828 (N_3828,N_1926,N_883);
and U3829 (N_3829,N_1163,N_46);
and U3830 (N_3830,N_980,N_1877);
and U3831 (N_3831,N_1239,N_740);
nand U3832 (N_3832,N_353,N_495);
nand U3833 (N_3833,N_1332,N_1856);
and U3834 (N_3834,N_1586,N_651);
nor U3835 (N_3835,N_1794,N_1841);
nand U3836 (N_3836,N_441,N_1539);
or U3837 (N_3837,N_1715,N_430);
or U3838 (N_3838,N_1229,N_272);
and U3839 (N_3839,N_931,N_1991);
nor U3840 (N_3840,N_191,N_1014);
nor U3841 (N_3841,N_1733,N_772);
nor U3842 (N_3842,N_584,N_393);
xor U3843 (N_3843,N_911,N_291);
or U3844 (N_3844,N_1494,N_1470);
and U3845 (N_3845,N_208,N_395);
and U3846 (N_3846,N_82,N_420);
or U3847 (N_3847,N_1495,N_158);
and U3848 (N_3848,N_1493,N_696);
or U3849 (N_3849,N_1918,N_1439);
nand U3850 (N_3850,N_1973,N_1434);
or U3851 (N_3851,N_627,N_1536);
or U3852 (N_3852,N_1718,N_1668);
and U3853 (N_3853,N_1201,N_1368);
and U3854 (N_3854,N_1727,N_1067);
nor U3855 (N_3855,N_620,N_534);
nor U3856 (N_3856,N_394,N_1782);
nand U3857 (N_3857,N_202,N_468);
nor U3858 (N_3858,N_629,N_612);
or U3859 (N_3859,N_0,N_757);
xor U3860 (N_3860,N_1654,N_1016);
nor U3861 (N_3861,N_603,N_245);
nand U3862 (N_3862,N_634,N_1352);
or U3863 (N_3863,N_561,N_1902);
nor U3864 (N_3864,N_1247,N_1533);
nand U3865 (N_3865,N_367,N_1295);
or U3866 (N_3866,N_1259,N_1692);
and U3867 (N_3867,N_284,N_1663);
nand U3868 (N_3868,N_771,N_1057);
or U3869 (N_3869,N_39,N_989);
or U3870 (N_3870,N_517,N_1892);
xnor U3871 (N_3871,N_455,N_341);
xnor U3872 (N_3872,N_1036,N_145);
or U3873 (N_3873,N_1470,N_884);
or U3874 (N_3874,N_1905,N_1847);
nand U3875 (N_3875,N_87,N_712);
nand U3876 (N_3876,N_1162,N_151);
nor U3877 (N_3877,N_430,N_1695);
xor U3878 (N_3878,N_232,N_921);
or U3879 (N_3879,N_1861,N_940);
xnor U3880 (N_3880,N_955,N_223);
nand U3881 (N_3881,N_605,N_1381);
xor U3882 (N_3882,N_147,N_1876);
and U3883 (N_3883,N_1070,N_1142);
xnor U3884 (N_3884,N_1192,N_55);
nor U3885 (N_3885,N_1910,N_405);
nand U3886 (N_3886,N_12,N_1827);
nand U3887 (N_3887,N_1815,N_1461);
or U3888 (N_3888,N_1093,N_820);
nand U3889 (N_3889,N_1060,N_1007);
nand U3890 (N_3890,N_243,N_607);
nand U3891 (N_3891,N_820,N_1531);
xor U3892 (N_3892,N_38,N_1589);
xnor U3893 (N_3893,N_1633,N_713);
and U3894 (N_3894,N_1553,N_105);
and U3895 (N_3895,N_788,N_1944);
nor U3896 (N_3896,N_1413,N_415);
xor U3897 (N_3897,N_617,N_228);
nor U3898 (N_3898,N_1750,N_229);
or U3899 (N_3899,N_136,N_530);
nor U3900 (N_3900,N_1267,N_1660);
nor U3901 (N_3901,N_17,N_517);
or U3902 (N_3902,N_1234,N_1003);
xor U3903 (N_3903,N_547,N_435);
or U3904 (N_3904,N_1798,N_1226);
nand U3905 (N_3905,N_1922,N_1339);
nand U3906 (N_3906,N_1893,N_220);
or U3907 (N_3907,N_1500,N_1613);
and U3908 (N_3908,N_243,N_699);
or U3909 (N_3909,N_997,N_831);
nor U3910 (N_3910,N_498,N_1074);
and U3911 (N_3911,N_1329,N_283);
or U3912 (N_3912,N_1432,N_1644);
or U3913 (N_3913,N_983,N_136);
xnor U3914 (N_3914,N_1337,N_720);
nand U3915 (N_3915,N_861,N_108);
xor U3916 (N_3916,N_156,N_60);
nand U3917 (N_3917,N_238,N_53);
xor U3918 (N_3918,N_1503,N_426);
nand U3919 (N_3919,N_783,N_109);
nand U3920 (N_3920,N_806,N_959);
and U3921 (N_3921,N_1170,N_646);
xnor U3922 (N_3922,N_996,N_234);
xnor U3923 (N_3923,N_1243,N_192);
nand U3924 (N_3924,N_1238,N_1608);
and U3925 (N_3925,N_1045,N_631);
nand U3926 (N_3926,N_1803,N_961);
nand U3927 (N_3927,N_831,N_416);
nor U3928 (N_3928,N_1874,N_311);
and U3929 (N_3929,N_852,N_1502);
nor U3930 (N_3930,N_630,N_933);
nand U3931 (N_3931,N_1769,N_842);
xnor U3932 (N_3932,N_19,N_1093);
nor U3933 (N_3933,N_1771,N_1436);
nor U3934 (N_3934,N_253,N_368);
nor U3935 (N_3935,N_1477,N_1416);
or U3936 (N_3936,N_1756,N_245);
and U3937 (N_3937,N_1079,N_154);
nor U3938 (N_3938,N_1830,N_1036);
nand U3939 (N_3939,N_363,N_1678);
and U3940 (N_3940,N_506,N_1063);
or U3941 (N_3941,N_1420,N_1058);
xnor U3942 (N_3942,N_653,N_937);
nor U3943 (N_3943,N_1976,N_1040);
nor U3944 (N_3944,N_1448,N_1438);
or U3945 (N_3945,N_440,N_6);
nor U3946 (N_3946,N_1287,N_548);
xor U3947 (N_3947,N_1310,N_1202);
nor U3948 (N_3948,N_467,N_861);
nand U3949 (N_3949,N_1571,N_1694);
nor U3950 (N_3950,N_1755,N_808);
nor U3951 (N_3951,N_1101,N_124);
xnor U3952 (N_3952,N_488,N_1645);
nand U3953 (N_3953,N_1318,N_1753);
or U3954 (N_3954,N_693,N_474);
nor U3955 (N_3955,N_135,N_1319);
and U3956 (N_3956,N_757,N_335);
xnor U3957 (N_3957,N_581,N_124);
nand U3958 (N_3958,N_1116,N_9);
or U3959 (N_3959,N_1340,N_1344);
nand U3960 (N_3960,N_767,N_1190);
xor U3961 (N_3961,N_193,N_1295);
and U3962 (N_3962,N_722,N_1444);
xnor U3963 (N_3963,N_286,N_1844);
nand U3964 (N_3964,N_601,N_321);
or U3965 (N_3965,N_611,N_1912);
nor U3966 (N_3966,N_1289,N_1067);
nand U3967 (N_3967,N_1854,N_1117);
xnor U3968 (N_3968,N_25,N_47);
or U3969 (N_3969,N_1191,N_1897);
nor U3970 (N_3970,N_409,N_806);
and U3971 (N_3971,N_1294,N_1331);
xnor U3972 (N_3972,N_1832,N_824);
and U3973 (N_3973,N_120,N_1164);
and U3974 (N_3974,N_291,N_1072);
and U3975 (N_3975,N_1883,N_1222);
xor U3976 (N_3976,N_1117,N_817);
nor U3977 (N_3977,N_40,N_1441);
or U3978 (N_3978,N_1511,N_1436);
nand U3979 (N_3979,N_1970,N_68);
nand U3980 (N_3980,N_981,N_1147);
nor U3981 (N_3981,N_1291,N_1874);
or U3982 (N_3982,N_1548,N_1790);
or U3983 (N_3983,N_1668,N_1237);
xor U3984 (N_3984,N_749,N_70);
and U3985 (N_3985,N_1138,N_1818);
nand U3986 (N_3986,N_1985,N_703);
nor U3987 (N_3987,N_16,N_1680);
nor U3988 (N_3988,N_663,N_596);
and U3989 (N_3989,N_776,N_17);
and U3990 (N_3990,N_916,N_344);
xor U3991 (N_3991,N_1126,N_1839);
xnor U3992 (N_3992,N_1824,N_905);
xnor U3993 (N_3993,N_868,N_638);
or U3994 (N_3994,N_213,N_958);
and U3995 (N_3995,N_1131,N_564);
nor U3996 (N_3996,N_1966,N_1999);
xor U3997 (N_3997,N_1168,N_1359);
or U3998 (N_3998,N_1445,N_1549);
nand U3999 (N_3999,N_595,N_1031);
xor U4000 (N_4000,N_2670,N_3077);
or U4001 (N_4001,N_3816,N_2018);
or U4002 (N_4002,N_2465,N_2424);
or U4003 (N_4003,N_2351,N_2453);
and U4004 (N_4004,N_2743,N_3306);
xor U4005 (N_4005,N_3994,N_2655);
nor U4006 (N_4006,N_3741,N_2399);
or U4007 (N_4007,N_3424,N_3511);
nor U4008 (N_4008,N_2051,N_3045);
and U4009 (N_4009,N_3349,N_3315);
and U4010 (N_4010,N_2922,N_3549);
and U4011 (N_4011,N_3825,N_2024);
nand U4012 (N_4012,N_2067,N_2837);
nand U4013 (N_4013,N_2805,N_2813);
nor U4014 (N_4014,N_3481,N_3889);
xor U4015 (N_4015,N_3347,N_2840);
nor U4016 (N_4016,N_2419,N_2416);
nor U4017 (N_4017,N_3290,N_2050);
xor U4018 (N_4018,N_2558,N_2625);
nand U4019 (N_4019,N_3401,N_2337);
nor U4020 (N_4020,N_3057,N_3430);
nand U4021 (N_4021,N_2291,N_2197);
and U4022 (N_4022,N_2409,N_3689);
xor U4023 (N_4023,N_3409,N_2597);
nor U4024 (N_4024,N_2282,N_3348);
and U4025 (N_4025,N_3949,N_3415);
or U4026 (N_4026,N_3851,N_3947);
nand U4027 (N_4027,N_3420,N_2868);
and U4028 (N_4028,N_3343,N_2442);
xor U4029 (N_4029,N_2888,N_3761);
xor U4030 (N_4030,N_3721,N_2085);
and U4031 (N_4031,N_3973,N_2885);
xnor U4032 (N_4032,N_3356,N_3564);
and U4033 (N_4033,N_2973,N_3153);
and U4034 (N_4034,N_2091,N_3346);
xnor U4035 (N_4035,N_2231,N_2201);
and U4036 (N_4036,N_2943,N_3517);
and U4037 (N_4037,N_3119,N_3890);
nand U4038 (N_4038,N_2652,N_2967);
or U4039 (N_4039,N_3908,N_2335);
or U4040 (N_4040,N_2347,N_3768);
nand U4041 (N_4041,N_2503,N_3276);
and U4042 (N_4042,N_3699,N_3626);
xnor U4043 (N_4043,N_2115,N_3571);
nand U4044 (N_4044,N_3054,N_2154);
or U4045 (N_4045,N_2981,N_3282);
nor U4046 (N_4046,N_2947,N_2415);
and U4047 (N_4047,N_2788,N_2595);
and U4048 (N_4048,N_3053,N_2302);
nor U4049 (N_4049,N_2483,N_3203);
nand U4050 (N_4050,N_2948,N_2339);
nand U4051 (N_4051,N_3565,N_2002);
or U4052 (N_4052,N_2699,N_3774);
nand U4053 (N_4053,N_2375,N_3362);
xnor U4054 (N_4054,N_2066,N_2327);
nand U4055 (N_4055,N_2946,N_3064);
nand U4056 (N_4056,N_2603,N_3916);
nor U4057 (N_4057,N_3378,N_2792);
nand U4058 (N_4058,N_2763,N_3807);
nand U4059 (N_4059,N_3232,N_3185);
nand U4060 (N_4060,N_2544,N_2149);
and U4061 (N_4061,N_3940,N_3550);
nand U4062 (N_4062,N_3188,N_2945);
or U4063 (N_4063,N_3753,N_3164);
or U4064 (N_4064,N_3813,N_2410);
or U4065 (N_4065,N_2538,N_2906);
and U4066 (N_4066,N_2144,N_2646);
nand U4067 (N_4067,N_3441,N_2283);
and U4068 (N_4068,N_3151,N_3854);
nand U4069 (N_4069,N_3144,N_3285);
or U4070 (N_4070,N_2262,N_2555);
or U4071 (N_4071,N_2049,N_2128);
nor U4072 (N_4072,N_2610,N_2851);
nand U4073 (N_4073,N_2364,N_2371);
xnor U4074 (N_4074,N_3089,N_2999);
xnor U4075 (N_4075,N_3101,N_3927);
nand U4076 (N_4076,N_3193,N_3486);
nor U4077 (N_4077,N_3043,N_2669);
and U4078 (N_4078,N_3097,N_3291);
nor U4079 (N_4079,N_3403,N_2042);
nor U4080 (N_4080,N_3122,N_2346);
xnor U4081 (N_4081,N_3044,N_2377);
xor U4082 (N_4082,N_2532,N_3148);
xnor U4083 (N_4083,N_2378,N_2682);
xnor U4084 (N_4084,N_2621,N_2914);
or U4085 (N_4085,N_2804,N_3166);
and U4086 (N_4086,N_3312,N_2101);
nor U4087 (N_4087,N_2352,N_2268);
or U4088 (N_4088,N_3313,N_2498);
nor U4089 (N_4089,N_3658,N_3557);
nand U4090 (N_4090,N_3061,N_3995);
nor U4091 (N_4091,N_3039,N_2834);
xnor U4092 (N_4092,N_2462,N_2496);
xnor U4093 (N_4093,N_3546,N_3720);
and U4094 (N_4094,N_3515,N_2658);
or U4095 (N_4095,N_3673,N_2494);
nor U4096 (N_4096,N_2299,N_2866);
nand U4097 (N_4097,N_3011,N_3706);
and U4098 (N_4098,N_2517,N_3685);
nor U4099 (N_4099,N_2044,N_2394);
and U4100 (N_4100,N_2725,N_2168);
nand U4101 (N_4101,N_3765,N_2475);
or U4102 (N_4102,N_3860,N_3627);
xor U4103 (N_4103,N_3862,N_2978);
xnor U4104 (N_4104,N_3206,N_2854);
nor U4105 (N_4105,N_3398,N_2512);
and U4106 (N_4106,N_2566,N_3674);
nand U4107 (N_4107,N_3577,N_3771);
nand U4108 (N_4108,N_2100,N_3539);
nand U4109 (N_4109,N_3158,N_3671);
and U4110 (N_4110,N_2216,N_3233);
or U4111 (N_4111,N_3170,N_2272);
nand U4112 (N_4112,N_2321,N_3635);
and U4113 (N_4113,N_3609,N_2434);
nor U4114 (N_4114,N_2531,N_3829);
xnor U4115 (N_4115,N_2705,N_3462);
nand U4116 (N_4116,N_2092,N_3742);
and U4117 (N_4117,N_2842,N_3319);
and U4118 (N_4118,N_2037,N_2439);
xor U4119 (N_4119,N_2234,N_2872);
nand U4120 (N_4120,N_3163,N_2421);
and U4121 (N_4121,N_3922,N_2070);
and U4122 (N_4122,N_3836,N_2203);
and U4123 (N_4123,N_2784,N_3190);
or U4124 (N_4124,N_2015,N_2820);
xor U4125 (N_4125,N_2255,N_2361);
nor U4126 (N_4126,N_2464,N_2300);
nand U4127 (N_4127,N_3328,N_3501);
xnor U4128 (N_4128,N_2276,N_2677);
and U4129 (N_4129,N_3778,N_3124);
and U4130 (N_4130,N_2401,N_2642);
and U4131 (N_4131,N_2949,N_3650);
nand U4132 (N_4132,N_2153,N_2167);
xnor U4133 (N_4133,N_2936,N_3579);
nor U4134 (N_4134,N_3624,N_3220);
or U4135 (N_4135,N_2160,N_3437);
xnor U4136 (N_4136,N_3918,N_2976);
and U4137 (N_4137,N_3411,N_2501);
xor U4138 (N_4138,N_2379,N_3270);
nand U4139 (N_4139,N_3373,N_2040);
or U4140 (N_4140,N_3267,N_2608);
or U4141 (N_4141,N_3230,N_2703);
xnor U4142 (N_4142,N_3909,N_3805);
or U4143 (N_4143,N_3387,N_3562);
and U4144 (N_4144,N_2123,N_2278);
or U4145 (N_4145,N_3663,N_3581);
nand U4146 (N_4146,N_3811,N_3978);
nor U4147 (N_4147,N_3265,N_2955);
and U4148 (N_4148,N_3772,N_3243);
and U4149 (N_4149,N_3361,N_2106);
xor U4150 (N_4150,N_2515,N_2265);
nor U4151 (N_4151,N_2455,N_3570);
and U4152 (N_4152,N_2374,N_2087);
and U4153 (N_4153,N_3422,N_2176);
or U4154 (N_4154,N_2870,N_2098);
nor U4155 (N_4155,N_2251,N_2097);
or U4156 (N_4156,N_3902,N_3724);
and U4157 (N_4157,N_3035,N_3351);
xnor U4158 (N_4158,N_3913,N_2309);
nand U4159 (N_4159,N_2131,N_2794);
xnor U4160 (N_4160,N_3715,N_3677);
or U4161 (N_4161,N_3896,N_2175);
and U4162 (N_4162,N_3912,N_2565);
xnor U4163 (N_4163,N_3229,N_2103);
nand U4164 (N_4164,N_3817,N_3499);
or U4165 (N_4165,N_2769,N_2698);
nor U4166 (N_4166,N_3357,N_3228);
nor U4167 (N_4167,N_2504,N_2202);
nand U4168 (N_4168,N_2323,N_2264);
nand U4169 (N_4169,N_3618,N_3819);
and U4170 (N_4170,N_2457,N_3798);
nor U4171 (N_4171,N_2497,N_3344);
nand U4172 (N_4172,N_2893,N_3897);
nor U4173 (N_4173,N_2676,N_3558);
and U4174 (N_4174,N_2634,N_2916);
nand U4175 (N_4175,N_2900,N_3845);
and U4176 (N_4176,N_2675,N_3749);
or U4177 (N_4177,N_3885,N_3189);
or U4178 (N_4178,N_2289,N_3779);
xor U4179 (N_4179,N_2683,N_3784);
nor U4180 (N_4180,N_3429,N_2523);
or U4181 (N_4181,N_3264,N_2225);
nor U4182 (N_4182,N_2073,N_3612);
or U4183 (N_4183,N_2613,N_2545);
and U4184 (N_4184,N_2245,N_3605);
and U4185 (N_4185,N_3554,N_3544);
or U4186 (N_4186,N_3252,N_2127);
nand U4187 (N_4187,N_3591,N_3958);
xor U4188 (N_4188,N_2431,N_2065);
or U4189 (N_4189,N_3196,N_2172);
and U4190 (N_4190,N_2458,N_3414);
nand U4191 (N_4191,N_2965,N_2200);
or U4192 (N_4192,N_3510,N_3110);
nor U4193 (N_4193,N_3944,N_3421);
nand U4194 (N_4194,N_2749,N_3652);
and U4195 (N_4195,N_2731,N_2081);
and U4196 (N_4196,N_2724,N_3865);
xor U4197 (N_4197,N_3145,N_2240);
or U4198 (N_4198,N_3574,N_2719);
nor U4199 (N_4199,N_2112,N_2782);
and U4200 (N_4200,N_3251,N_2006);
nor U4201 (N_4201,N_2816,N_3714);
nor U4202 (N_4202,N_2461,N_3542);
or U4203 (N_4203,N_3079,N_2537);
or U4204 (N_4204,N_2672,N_2466);
nor U4205 (N_4205,N_2933,N_3425);
and U4206 (N_4206,N_2223,N_3777);
and U4207 (N_4207,N_3987,N_2806);
or U4208 (N_4208,N_3795,N_3732);
or U4209 (N_4209,N_2736,N_2329);
xor U4210 (N_4210,N_2564,N_2139);
xor U4211 (N_4211,N_3360,N_3575);
and U4212 (N_4212,N_2623,N_2078);
nand U4213 (N_4213,N_3876,N_2484);
xnor U4214 (N_4214,N_2579,N_2381);
nand U4215 (N_4215,N_3586,N_3314);
xnor U4216 (N_4216,N_3186,N_2875);
or U4217 (N_4217,N_2758,N_2190);
nor U4218 (N_4218,N_2985,N_2052);
xnor U4219 (N_4219,N_3849,N_3428);
or U4220 (N_4220,N_2954,N_3009);
nand U4221 (N_4221,N_2845,N_3100);
or U4222 (N_4222,N_2632,N_3582);
nand U4223 (N_4223,N_2372,N_2932);
and U4224 (N_4224,N_3369,N_3820);
or U4225 (N_4225,N_3456,N_3049);
nor U4226 (N_4226,N_3841,N_3921);
and U4227 (N_4227,N_2340,N_2395);
nand U4228 (N_4228,N_2576,N_2427);
or U4229 (N_4229,N_3967,N_3727);
or U4230 (N_4230,N_3178,N_2226);
xnor U4231 (N_4231,N_3480,N_2288);
nor U4232 (N_4232,N_2297,N_3971);
xor U4233 (N_4233,N_3096,N_2185);
nor U4234 (N_4234,N_2239,N_3996);
nand U4235 (N_4235,N_2867,N_3585);
xor U4236 (N_4236,N_2796,N_2312);
nand U4237 (N_4237,N_3269,N_3969);
or U4238 (N_4238,N_3638,N_3171);
nor U4239 (N_4239,N_3678,N_3262);
nor U4240 (N_4240,N_3036,N_2376);
nand U4241 (N_4241,N_3333,N_2486);
and U4242 (N_4242,N_2706,N_2310);
or U4243 (N_4243,N_2471,N_3878);
nand U4244 (N_4244,N_3823,N_2298);
nand U4245 (N_4245,N_2338,N_2666);
xor U4246 (N_4246,N_2193,N_2145);
nor U4247 (N_4247,N_2825,N_2133);
or U4248 (N_4248,N_3926,N_3274);
or U4249 (N_4249,N_3273,N_3263);
nand U4250 (N_4250,N_2490,N_3888);
nor U4251 (N_4251,N_2650,N_3078);
xor U4252 (N_4252,N_3466,N_2492);
xnor U4253 (N_4253,N_3358,N_2191);
or U4254 (N_4254,N_3129,N_3371);
xnor U4255 (N_4255,N_3234,N_3223);
or U4256 (N_4256,N_3479,N_2952);
and U4257 (N_4257,N_3716,N_3353);
and U4258 (N_4258,N_3470,N_2199);
or U4259 (N_4259,N_2445,N_3717);
and U4260 (N_4260,N_3729,N_2077);
and U4261 (N_4261,N_2207,N_2863);
and U4262 (N_4262,N_2068,N_3990);
xnor U4263 (N_4263,N_3152,N_3156);
or U4264 (N_4264,N_2311,N_3033);
and U4265 (N_4265,N_3906,N_2417);
and U4266 (N_4266,N_3394,N_2478);
and U4267 (N_4267,N_2720,N_2826);
nand U4268 (N_4268,N_2741,N_2083);
or U4269 (N_4269,N_3873,N_2522);
nand U4270 (N_4270,N_3527,N_2974);
or U4271 (N_4271,N_2930,N_2890);
or U4272 (N_4272,N_2815,N_2560);
xnor U4273 (N_4273,N_2228,N_3051);
nand U4274 (N_4274,N_2929,N_2937);
or U4275 (N_4275,N_3834,N_2041);
xnor U4276 (N_4276,N_3601,N_3307);
nor U4277 (N_4277,N_3238,N_3055);
xor U4278 (N_4278,N_3954,N_2204);
or U4279 (N_4279,N_3725,N_3381);
xnor U4280 (N_4280,N_3001,N_3676);
nand U4281 (N_4281,N_2832,N_2295);
xnor U4282 (N_4282,N_3628,N_2263);
nor U4283 (N_4283,N_2005,N_2111);
xor U4284 (N_4284,N_3694,N_2689);
xnor U4285 (N_4285,N_3484,N_2166);
xnor U4286 (N_4286,N_3696,N_3283);
or U4287 (N_4287,N_2437,N_2502);
and U4288 (N_4288,N_3194,N_3275);
nand U4289 (N_4289,N_2206,N_3372);
and U4290 (N_4290,N_2161,N_3058);
nand U4291 (N_4291,N_3580,N_3174);
xor U4292 (N_4292,N_3463,N_2607);
xor U4293 (N_4293,N_3117,N_2007);
nand U4294 (N_4294,N_3900,N_3250);
xnor U4295 (N_4295,N_2674,N_2817);
and U4296 (N_4296,N_3157,N_3123);
xnor U4297 (N_4297,N_2877,N_3211);
nand U4298 (N_4298,N_3801,N_2744);
or U4299 (N_4299,N_3733,N_3641);
nor U4300 (N_4300,N_3867,N_2107);
and U4301 (N_4301,N_2491,N_3329);
xnor U4302 (N_4302,N_2649,N_3740);
nand U4303 (N_4303,N_3653,N_3933);
xnor U4304 (N_4304,N_2902,N_3050);
nor U4305 (N_4305,N_2430,N_2156);
nand U4306 (N_4306,N_3320,N_2661);
xnor U4307 (N_4307,N_3533,N_2447);
and U4308 (N_4308,N_2671,N_2173);
nand U4309 (N_4309,N_3340,N_3367);
and U4310 (N_4310,N_3118,N_3986);
xor U4311 (N_4311,N_3620,N_3448);
or U4312 (N_4312,N_3983,N_3294);
nor U4313 (N_4313,N_2746,N_2992);
or U4314 (N_4314,N_3032,N_3938);
or U4315 (N_4315,N_2056,N_2126);
nor U4316 (N_4316,N_2961,N_3848);
nor U4317 (N_4317,N_3891,N_2186);
xor U4318 (N_4318,N_3828,N_3132);
nor U4319 (N_4319,N_3114,N_3611);
nand U4320 (N_4320,N_3402,N_2996);
xnor U4321 (N_4321,N_3426,N_2393);
or U4322 (N_4322,N_2177,N_2356);
and U4323 (N_4323,N_2257,N_2765);
nor U4324 (N_4324,N_3785,N_3710);
and U4325 (N_4325,N_2581,N_2861);
xor U4326 (N_4326,N_3091,N_2053);
xor U4327 (N_4327,N_2871,N_3702);
nand U4328 (N_4328,N_3094,N_3201);
or U4329 (N_4329,N_3826,N_3443);
nor U4330 (N_4330,N_2700,N_2909);
nor U4331 (N_4331,N_2624,N_3959);
xor U4332 (N_4332,N_2125,N_3111);
nor U4333 (N_4333,N_2857,N_3697);
and U4334 (N_4334,N_3690,N_2865);
or U4335 (N_4335,N_2891,N_3406);
nand U4336 (N_4336,N_2472,N_2102);
or U4337 (N_4337,N_3831,N_2386);
nor U4338 (N_4338,N_2275,N_3955);
or U4339 (N_4339,N_2680,N_3284);
xor U4340 (N_4340,N_2152,N_2456);
and U4341 (N_4341,N_3915,N_3300);
nor U4342 (N_4342,N_3842,N_2222);
xor U4343 (N_4343,N_2715,N_3520);
nor U4344 (N_4344,N_3334,N_3476);
or U4345 (N_4345,N_3625,N_3606);
nand U4346 (N_4346,N_2164,N_3984);
or U4347 (N_4347,N_2760,N_2058);
nand U4348 (N_4348,N_2489,N_3803);
nor U4349 (N_4349,N_2829,N_3667);
xor U4350 (N_4350,N_2991,N_2235);
xnor U4351 (N_4351,N_2679,N_2575);
nor U4352 (N_4352,N_2957,N_2198);
xnor U4353 (N_4353,N_2368,N_2232);
nand U4354 (N_4354,N_3532,N_3418);
nor U4355 (N_4355,N_3493,N_3404);
nand U4356 (N_4356,N_3634,N_3509);
nand U4357 (N_4357,N_3212,N_2830);
and U4358 (N_4358,N_2879,N_3668);
xnor U4359 (N_4359,N_2010,N_3098);
nand U4360 (N_4360,N_3109,N_2539);
nand U4361 (N_4361,N_3855,N_3442);
nor U4362 (N_4362,N_2884,N_3400);
and U4363 (N_4363,N_2525,N_2269);
nand U4364 (N_4364,N_2165,N_3695);
and U4365 (N_4365,N_2732,N_3128);
and U4366 (N_4366,N_3108,N_2433);
nand U4367 (N_4367,N_3713,N_2729);
nand U4368 (N_4368,N_3198,N_3245);
nor U4369 (N_4369,N_3258,N_3877);
or U4370 (N_4370,N_2350,N_2099);
and U4371 (N_4371,N_2307,N_3008);
or U4372 (N_4372,N_3863,N_2969);
or U4373 (N_4373,N_3370,N_3412);
or U4374 (N_4374,N_3134,N_2499);
nor U4375 (N_4375,N_2648,N_2249);
nor U4376 (N_4376,N_2305,N_2668);
and U4377 (N_4377,N_2205,N_3814);
or U4378 (N_4378,N_2398,N_2811);
xor U4379 (N_4379,N_3875,N_3964);
and U4380 (N_4380,N_3491,N_3524);
xnor U4381 (N_4381,N_2392,N_3553);
and U4382 (N_4382,N_2353,N_3543);
xnor U4383 (N_4383,N_2754,N_2904);
or U4384 (N_4384,N_2901,N_2827);
and U4385 (N_4385,N_2956,N_3461);
or U4386 (N_4386,N_2638,N_2448);
xnor U4387 (N_4387,N_2903,N_3281);
nand U4388 (N_4388,N_3576,N_2983);
or U4389 (N_4389,N_3155,N_2147);
or U4390 (N_4390,N_3376,N_2915);
or U4391 (N_4391,N_3856,N_3205);
or U4392 (N_4392,N_3730,N_3968);
xor U4393 (N_4393,N_2063,N_2046);
or U4394 (N_4394,N_2951,N_2285);
nor U4395 (N_4395,N_2778,N_2640);
and U4396 (N_4396,N_3278,N_3898);
xnor U4397 (N_4397,N_3536,N_2514);
nor U4398 (N_4398,N_3599,N_2331);
nor U4399 (N_4399,N_3683,N_2301);
xor U4400 (N_4400,N_2519,N_3594);
xor U4401 (N_4401,N_2941,N_3235);
or U4402 (N_4402,N_2384,N_2034);
xnor U4403 (N_4403,N_3997,N_3086);
and U4404 (N_4404,N_2839,N_2318);
nor U4405 (N_4405,N_3072,N_3615);
nand U4406 (N_4406,N_2690,N_3453);
or U4407 (N_4407,N_3088,N_3701);
or U4408 (N_4408,N_3385,N_3458);
nor U4409 (N_4409,N_2121,N_2209);
or U4410 (N_4410,N_3718,N_3604);
nand U4411 (N_4411,N_3503,N_3824);
xnor U4412 (N_4412,N_2020,N_2730);
nor U4413 (N_4413,N_3139,N_3081);
or U4414 (N_4414,N_2691,N_2117);
or U4415 (N_4415,N_3071,N_2896);
nand U4416 (N_4416,N_3127,N_2261);
xnor U4417 (N_4417,N_2477,N_2707);
or U4418 (N_4418,N_3872,N_3596);
or U4419 (N_4419,N_2776,N_3154);
xnor U4420 (N_4420,N_2214,N_3384);
xor U4421 (N_4421,N_2855,N_3248);
xnor U4422 (N_4422,N_2571,N_3953);
xnor U4423 (N_4423,N_3177,N_2391);
nand U4424 (N_4424,N_2143,N_2137);
nor U4425 (N_4425,N_2924,N_2894);
nor U4426 (N_4426,N_2075,N_3521);
and U4427 (N_4427,N_2345,N_2605);
nand U4428 (N_4428,N_3477,N_2609);
nor U4429 (N_4429,N_3861,N_3490);
nor U4430 (N_4430,N_3450,N_3810);
and U4431 (N_4431,N_3060,N_2182);
nor U4432 (N_4432,N_3998,N_2753);
nor U4433 (N_4433,N_3286,N_3893);
or U4434 (N_4434,N_2850,N_3600);
nor U4435 (N_4435,N_3126,N_2972);
nand U4436 (N_4436,N_2485,N_2270);
and U4437 (N_4437,N_3766,N_3946);
or U4438 (N_4438,N_3103,N_2614);
and U4439 (N_4439,N_3514,N_2230);
nand U4440 (N_4440,N_2667,N_3870);
nand U4441 (N_4441,N_2822,N_3272);
xor U4442 (N_4442,N_3950,N_3444);
nand U4443 (N_4443,N_2479,N_3037);
xnor U4444 (N_4444,N_2170,N_2516);
or U4445 (N_4445,N_2412,N_2030);
or U4446 (N_4446,N_2510,N_3452);
and U4447 (N_4447,N_3197,N_3208);
xnor U4448 (N_4448,N_2988,N_3240);
and U4449 (N_4449,N_3130,N_2777);
or U4450 (N_4450,N_3859,N_3762);
and U4451 (N_4451,N_3522,N_2195);
xor U4452 (N_4452,N_2071,N_2064);
and U4453 (N_4453,N_2836,N_2146);
nor U4454 (N_4454,N_2783,N_2124);
or U4455 (N_4455,N_2881,N_3743);
and U4456 (N_4456,N_2779,N_2799);
and U4457 (N_4457,N_3726,N_2158);
xor U4458 (N_4458,N_2362,N_2513);
xor U4459 (N_4459,N_3488,N_2968);
or U4460 (N_4460,N_2208,N_2509);
nand U4461 (N_4461,N_2174,N_2878);
or U4462 (N_4462,N_3722,N_2400);
nand U4463 (N_4463,N_2279,N_3843);
or U4464 (N_4464,N_3224,N_2267);
nor U4465 (N_4465,N_2027,N_3413);
or U4466 (N_4466,N_2495,N_3090);
nand U4467 (N_4467,N_3073,N_2292);
or U4468 (N_4468,N_2550,N_3654);
xor U4469 (N_4469,N_3665,N_2897);
xnor U4470 (N_4470,N_2459,N_3105);
or U4471 (N_4471,N_3095,N_3808);
nand U4472 (N_4472,N_2620,N_3982);
and U4473 (N_4473,N_2918,N_3815);
xor U4474 (N_4474,N_3309,N_2330);
or U4475 (N_4475,N_3711,N_2665);
nand U4476 (N_4476,N_3979,N_2762);
and U4477 (N_4477,N_3468,N_2118);
nor U4478 (N_4478,N_2481,N_2132);
xor U4479 (N_4479,N_3545,N_3438);
or U4480 (N_4480,N_3478,N_3603);
xnor U4481 (N_4481,N_2694,N_2599);
xnor U4482 (N_4482,N_3059,N_2684);
nor U4483 (N_4483,N_2835,N_2585);
and U4484 (N_4484,N_2563,N_2641);
or U4485 (N_4485,N_2761,N_3776);
xor U4486 (N_4486,N_3648,N_3709);
nand U4487 (N_4487,N_3253,N_3305);
and U4488 (N_4488,N_2358,N_3204);
nand U4489 (N_4489,N_3773,N_3631);
xor U4490 (N_4490,N_3492,N_2029);
xor U4491 (N_4491,N_2454,N_2786);
nor U4492 (N_4492,N_2217,N_2468);
nor U4493 (N_4493,N_3892,N_2443);
and U4494 (N_4494,N_2553,N_2882);
or U4495 (N_4495,N_2561,N_2592);
or U4496 (N_4496,N_3160,N_3882);
or U4497 (N_4497,N_3850,N_2953);
nand U4498 (N_4498,N_3167,N_2920);
or U4499 (N_4499,N_3822,N_3405);
nand U4500 (N_4500,N_3999,N_3303);
nor U4501 (N_4501,N_2413,N_3046);
nor U4502 (N_4502,N_2246,N_3181);
nor U4503 (N_4503,N_3786,N_2921);
and U4504 (N_4504,N_3146,N_3217);
and U4505 (N_4505,N_3473,N_3844);
or U4506 (N_4506,N_2506,N_2644);
or U4507 (N_4507,N_3316,N_3617);
or U4508 (N_4508,N_3952,N_2508);
nand U4509 (N_4509,N_2578,N_2582);
xor U4510 (N_4510,N_3149,N_3182);
or U4511 (N_4511,N_2254,N_2584);
and U4512 (N_4512,N_2714,N_2662);
xor U4513 (N_4513,N_3445,N_2540);
nor U4514 (N_4514,N_2348,N_3407);
and U4515 (N_4515,N_2460,N_3965);
and U4516 (N_4516,N_2480,N_3975);
or U4517 (N_4517,N_3084,N_2373);
and U4518 (N_4518,N_3988,N_3537);
or U4519 (N_4519,N_3295,N_3302);
nand U4520 (N_4520,N_3592,N_2045);
nand U4521 (N_4521,N_3395,N_2521);
xor U4522 (N_4522,N_3957,N_3669);
xor U4523 (N_4523,N_2322,N_3970);
nor U4524 (N_4524,N_2511,N_2527);
nand U4525 (N_4525,N_2643,N_2938);
xor U4526 (N_4526,N_3003,N_2993);
or U4527 (N_4527,N_2141,N_2033);
nor U4528 (N_4528,N_3708,N_3487);
nor U4529 (N_4529,N_3530,N_3780);
and U4530 (N_4530,N_3236,N_3002);
or U4531 (N_4531,N_3853,N_3221);
xor U4532 (N_4532,N_2789,N_3383);
and U4533 (N_4533,N_3389,N_2617);
or U4534 (N_4534,N_3956,N_3176);
nand U4535 (N_4535,N_3643,N_3924);
and U4536 (N_4536,N_3140,N_3244);
xor U4537 (N_4537,N_2096,N_2733);
nor U4538 (N_4538,N_2631,N_3962);
nand U4539 (N_4539,N_3213,N_2334);
nand U4540 (N_4540,N_2319,N_3021);
nand U4541 (N_4541,N_2023,N_2213);
nand U4542 (N_4542,N_3507,N_2151);
nor U4543 (N_4543,N_2728,N_2136);
and U4544 (N_4544,N_3857,N_2615);
and U4545 (N_4545,N_2917,N_2950);
nor U4546 (N_4546,N_3218,N_3607);
or U4547 (N_4547,N_2718,N_2241);
or U4548 (N_4548,N_2220,N_2600);
or U4549 (N_4549,N_2629,N_3419);
and U4550 (N_4550,N_3847,N_3439);
nand U4551 (N_4551,N_3573,N_2547);
or U4552 (N_4552,N_3354,N_2403);
nor U4553 (N_4553,N_3028,N_2543);
nand U4554 (N_4554,N_2179,N_3266);
and U4555 (N_4555,N_2341,N_3447);
nor U4556 (N_4556,N_2534,N_2975);
xor U4557 (N_4557,N_3756,N_3363);
or U4558 (N_4558,N_3764,N_2907);
nor U4559 (N_4559,N_3538,N_2536);
nor U4560 (N_4560,N_2113,N_3026);
nand U4561 (N_4561,N_3992,N_3326);
nor U4562 (N_4562,N_3548,N_2316);
and U4563 (N_4563,N_3184,N_3981);
nor U4564 (N_4564,N_3977,N_2734);
xnor U4565 (N_4565,N_2908,N_2619);
nor U4566 (N_4566,N_2739,N_3556);
xor U4567 (N_4567,N_2635,N_2385);
or U4568 (N_4568,N_3074,N_2692);
or U4569 (N_4569,N_2737,N_2047);
nor U4570 (N_4570,N_3647,N_2611);
or U4571 (N_4571,N_2678,N_2693);
xnor U4572 (N_4572,N_3723,N_3796);
nand U4573 (N_4573,N_2218,N_3904);
nor U4574 (N_4574,N_3559,N_3365);
nor U4575 (N_4575,N_2148,N_2653);
nand U4576 (N_4576,N_3006,N_2290);
xor U4577 (N_4577,N_3748,N_3399);
or U4578 (N_4578,N_3871,N_3219);
nor U4579 (N_4579,N_2864,N_2277);
or U4580 (N_4580,N_3242,N_2697);
xor U4581 (N_4581,N_3566,N_3014);
and U4582 (N_4582,N_3806,N_3868);
nor U4583 (N_4583,N_3679,N_3561);
nand U4584 (N_4584,N_2332,N_2838);
xnor U4585 (N_4585,N_3432,N_2601);
nor U4586 (N_4586,N_3593,N_3022);
or U4587 (N_4587,N_3525,N_3231);
or U4588 (N_4588,N_3299,N_2344);
and U4589 (N_4589,N_3738,N_3874);
nor U4590 (N_4590,N_2260,N_3731);
nand U4591 (N_4591,N_2435,N_3903);
nor U4592 (N_4592,N_2821,N_2911);
nor U4593 (N_4593,N_2696,N_3040);
nand U4594 (N_4594,N_3680,N_2554);
xnor U4595 (N_4595,N_3963,N_3980);
or U4596 (N_4596,N_2663,N_2673);
nand U4597 (N_4597,N_2627,N_2824);
or U4598 (N_4598,N_2004,N_3416);
and U4599 (N_4599,N_3832,N_3293);
nor U4600 (N_4600,N_3052,N_2647);
or U4601 (N_4601,N_3472,N_2966);
or U4602 (N_4602,N_2000,N_2236);
xnor U4603 (N_4603,N_3569,N_2304);
xor U4604 (N_4604,N_3589,N_3734);
nand U4605 (N_4605,N_3341,N_3168);
nor U4606 (N_4606,N_3567,N_2450);
and U4607 (N_4607,N_3065,N_3712);
xor U4608 (N_4608,N_2022,N_3688);
or U4609 (N_4609,N_3015,N_3636);
or U4610 (N_4610,N_3568,N_3787);
xnor U4611 (N_4611,N_3960,N_3112);
nor U4612 (N_4612,N_3737,N_2927);
and U4613 (N_4613,N_3031,N_3707);
and U4614 (N_4614,N_3700,N_2651);
and U4615 (N_4615,N_3173,N_2036);
xor U4616 (N_4616,N_3788,N_2695);
nor U4617 (N_4617,N_2129,N_2317);
nand U4618 (N_4618,N_3427,N_2998);
nor U4619 (N_4619,N_3930,N_2211);
nand U4620 (N_4620,N_2104,N_2895);
and U4621 (N_4621,N_2014,N_2899);
or U4622 (N_4622,N_3180,N_3120);
or U4623 (N_4623,N_3025,N_3649);
xnor U4624 (N_4624,N_2227,N_3018);
and U4625 (N_4625,N_2748,N_2090);
and U4626 (N_4626,N_3007,N_2809);
or U4627 (N_4627,N_3797,N_2685);
xnor U4628 (N_4628,N_2354,N_2408);
nor U4629 (N_4629,N_2574,N_3410);
and U4630 (N_4630,N_3297,N_2701);
nand U4631 (N_4631,N_2716,N_3526);
or U4632 (N_4632,N_2130,N_3719);
xnor U4633 (N_4633,N_2654,N_2404);
xor U4634 (N_4634,N_2664,N_2740);
xnor U4635 (N_4635,N_2287,N_2407);
or U4636 (N_4636,N_2557,N_3932);
nor U4637 (N_4637,N_2281,N_2402);
xor U4638 (N_4638,N_2819,N_3754);
or U4639 (N_4639,N_3255,N_3705);
xnor U4640 (N_4640,N_3063,N_2482);
nand U4641 (N_4641,N_3728,N_2583);
or U4642 (N_4642,N_2336,N_3321);
xnor U4643 (N_4643,N_3692,N_3989);
xnor U4644 (N_4644,N_2021,N_2926);
nand U4645 (N_4645,N_3608,N_2529);
nor U4646 (N_4646,N_3397,N_3417);
or U4647 (N_4647,N_3460,N_2723);
xnor U4648 (N_4648,N_2586,N_3209);
nor U4649 (N_4649,N_2883,N_2224);
or U4650 (N_4650,N_3789,N_2054);
or U4651 (N_4651,N_2406,N_2038);
xor U4652 (N_4652,N_2687,N_3451);
nand U4653 (N_4653,N_2791,N_3782);
and U4654 (N_4654,N_3662,N_3261);
or U4655 (N_4655,N_2823,N_3534);
or U4656 (N_4656,N_2055,N_3345);
nand U4657 (N_4657,N_3000,N_2181);
and U4658 (N_4658,N_3069,N_3366);
nor U4659 (N_4659,N_2810,N_2061);
xor U4660 (N_4660,N_2587,N_2438);
nand U4661 (N_4661,N_3335,N_2708);
nor U4662 (N_4662,N_3687,N_3379);
xor U4663 (N_4663,N_2048,N_3852);
nor U4664 (N_4664,N_2541,N_3894);
or U4665 (N_4665,N_2183,N_3241);
xor U4666 (N_4666,N_3763,N_3133);
nand U4667 (N_4667,N_2296,N_2852);
and U4668 (N_4668,N_2757,N_2488);
nor U4669 (N_4669,N_2849,N_3076);
nand U4670 (N_4670,N_3068,N_2742);
xnor U4671 (N_4671,N_2923,N_2962);
nor U4672 (N_4672,N_3436,N_3659);
nand U4673 (N_4673,N_3202,N_3976);
nor U4674 (N_4674,N_3482,N_3529);
nor U4675 (N_4675,N_2886,N_2383);
nand U4676 (N_4676,N_3016,N_2326);
and U4677 (N_4677,N_3489,N_2645);
nand U4678 (N_4678,N_2380,N_2781);
nand U4679 (N_4679,N_3656,N_2114);
or U4680 (N_4680,N_3675,N_2079);
and U4681 (N_4681,N_2844,N_3093);
or U4682 (N_4682,N_2271,N_2420);
nor U4683 (N_4683,N_2856,N_3939);
or U4684 (N_4684,N_2764,N_2846);
xnor U4685 (N_4685,N_3317,N_2140);
or U4686 (N_4686,N_2591,N_3388);
xor U4687 (N_4687,N_3210,N_2636);
nor U4688 (N_4688,N_3901,N_2382);
and U4689 (N_4689,N_3135,N_2470);
nand U4690 (N_4690,N_3616,N_3092);
and U4691 (N_4691,N_2569,N_2343);
and U4692 (N_4692,N_3866,N_2315);
nor U4693 (N_4693,N_2633,N_3840);
nor U4694 (N_4694,N_3833,N_2169);
nor U4695 (N_4695,N_2596,N_2589);
and U4696 (N_4696,N_3660,N_3937);
and U4697 (N_4697,N_2780,N_2418);
or U4698 (N_4698,N_2892,N_3513);
nor U4699 (N_4699,N_2082,N_3408);
nor U4700 (N_4700,N_2032,N_3881);
or U4701 (N_4701,N_3374,N_3147);
nor U4702 (N_4702,N_3619,N_3377);
or U4703 (N_4703,N_3614,N_3257);
or U4704 (N_4704,N_3972,N_2328);
and U4705 (N_4705,N_2568,N_3237);
xnor U4706 (N_4706,N_3138,N_3013);
and U4707 (N_4707,N_2688,N_3082);
nor U4708 (N_4708,N_2979,N_2812);
and U4709 (N_4709,N_2759,N_3745);
xor U4710 (N_4710,N_2717,N_3350);
nor U4711 (N_4711,N_3019,N_2449);
and U4712 (N_4712,N_3500,N_2057);
nor U4713 (N_4713,N_3433,N_2196);
nand U4714 (N_4714,N_2971,N_2474);
xor U4715 (N_4715,N_2785,N_3375);
nor U4716 (N_4716,N_2997,N_2750);
or U4717 (N_4717,N_3337,N_2752);
xor U4718 (N_4718,N_2549,N_2726);
xnor U4719 (N_4719,N_3042,N_3280);
xnor U4720 (N_4720,N_3698,N_3655);
xor U4721 (N_4721,N_2552,N_3633);
nand U4722 (N_4722,N_2889,N_2530);
xor U4723 (N_4723,N_3390,N_2986);
nor U4724 (N_4724,N_3943,N_2286);
xnor U4725 (N_4725,N_2294,N_3884);
nor U4726 (N_4726,N_3070,N_3535);
xnor U4727 (N_4727,N_3393,N_3195);
and U4728 (N_4728,N_3494,N_3116);
xnor U4729 (N_4729,N_2802,N_2159);
and U4730 (N_4730,N_3338,N_3464);
nor U4731 (N_4731,N_3598,N_2505);
nor U4732 (N_4732,N_3113,N_3651);
nor U4733 (N_4733,N_2243,N_3942);
nand U4734 (N_4734,N_3259,N_2588);
nand U4735 (N_4735,N_3640,N_2982);
xnor U4736 (N_4736,N_2093,N_3107);
nand U4737 (N_4737,N_3664,N_2274);
and U4738 (N_4738,N_3271,N_2977);
xnor U4739 (N_4739,N_3102,N_2026);
or U4740 (N_4740,N_2001,N_3308);
and U4741 (N_4741,N_2995,N_3519);
nand U4742 (N_4742,N_2808,N_2388);
nor U4743 (N_4743,N_3322,N_3632);
nor U4744 (N_4744,N_2841,N_2960);
and U4745 (N_4745,N_2942,N_3352);
nor U4746 (N_4746,N_3886,N_3691);
nor U4747 (N_4747,N_3516,N_2119);
xnor U4748 (N_4748,N_2134,N_3622);
nor U4749 (N_4749,N_2874,N_2306);
nand U4750 (N_4750,N_2266,N_2355);
xnor U4751 (N_4751,N_2367,N_2980);
xor U4752 (N_4752,N_3304,N_3023);
xor U4753 (N_4753,N_3225,N_3917);
or U4754 (N_4754,N_3216,N_2313);
nand U4755 (N_4755,N_3584,N_2848);
nor U4756 (N_4756,N_3684,N_3380);
or U4757 (N_4757,N_2019,N_2847);
nor U4758 (N_4758,N_2772,N_3793);
xnor U4759 (N_4759,N_3289,N_3595);
and U4760 (N_4760,N_2548,N_3504);
and U4761 (N_4761,N_2711,N_3948);
nor U4762 (N_4762,N_3791,N_2573);
and U4763 (N_4763,N_2365,N_2787);
nand U4764 (N_4764,N_2109,N_3910);
or U4765 (N_4765,N_3004,N_2189);
and U4766 (N_4766,N_3359,N_2440);
or U4767 (N_4767,N_3880,N_3336);
and U4768 (N_4768,N_3864,N_3794);
and U4769 (N_4769,N_2467,N_2735);
or U4770 (N_4770,N_2273,N_2713);
or U4771 (N_4771,N_2446,N_3911);
nor U4772 (N_4772,N_2898,N_3821);
nor U4773 (N_4773,N_3083,N_2756);
xnor U4774 (N_4774,N_2768,N_3301);
xor U4775 (N_4775,N_3704,N_2088);
nor U4776 (N_4776,N_2259,N_2925);
and U4777 (N_4777,N_2533,N_3750);
xor U4778 (N_4778,N_2814,N_2721);
and U4779 (N_4779,N_3547,N_2284);
nand U4780 (N_4780,N_2366,N_3639);
nor U4781 (N_4781,N_3459,N_3523);
and U4782 (N_4782,N_3657,N_2546);
or U4783 (N_4783,N_2622,N_3435);
or U4784 (N_4784,N_3246,N_2389);
nor U4785 (N_4785,N_2451,N_3034);
nand U4786 (N_4786,N_2238,N_2593);
nand U4787 (N_4787,N_3578,N_3125);
nor U4788 (N_4788,N_2233,N_2444);
xnor U4789 (N_4789,N_3518,N_3038);
and U4790 (N_4790,N_3087,N_3899);
or U4791 (N_4791,N_3672,N_2256);
or U4792 (N_4792,N_3630,N_2188);
nor U4793 (N_4793,N_2405,N_2308);
nand U4794 (N_4794,N_2559,N_3563);
or U4795 (N_4795,N_2500,N_2017);
and U4796 (N_4796,N_3686,N_2598);
and U4797 (N_4797,N_3809,N_2862);
xnor U4798 (N_4798,N_2526,N_3928);
xnor U4799 (N_4799,N_3931,N_3528);
or U4800 (N_4800,N_3508,N_2577);
xor U4801 (N_4801,N_3066,N_3311);
nor U4802 (N_4802,N_2219,N_2518);
nand U4803 (N_4803,N_2250,N_3030);
and U4804 (N_4804,N_3757,N_2606);
xor U4805 (N_4805,N_3279,N_3474);
and U4806 (N_4806,N_2069,N_3835);
xor U4807 (N_4807,N_3498,N_3214);
and U4808 (N_4808,N_3142,N_2244);
xor U4809 (N_4809,N_3682,N_2359);
and U4810 (N_4810,N_2441,N_3506);
xnor U4811 (N_4811,N_3175,N_3839);
nand U4812 (N_4812,N_2387,N_3318);
xnor U4813 (N_4813,N_2873,N_3846);
nor U4814 (N_4814,N_3895,N_2084);
and U4815 (N_4815,N_3541,N_3012);
nand U4816 (N_4816,N_3227,N_2637);
nor U4817 (N_4817,N_3277,N_3804);
xor U4818 (N_4818,N_3191,N_3324);
or U4819 (N_4819,N_3382,N_3239);
or U4820 (N_4820,N_3759,N_3935);
and U4821 (N_4821,N_2542,N_2828);
or U4822 (N_4822,N_3254,N_2076);
nor U4823 (N_4823,N_3830,N_2414);
nand U4824 (N_4824,N_3368,N_2162);
nor U4825 (N_4825,N_2989,N_3165);
nand U4826 (N_4826,N_2003,N_3512);
nand U4827 (N_4827,N_2628,N_3590);
xor U4828 (N_4828,N_2012,N_2108);
xnor U4829 (N_4829,N_2452,N_2016);
xnor U4830 (N_4830,N_3961,N_2436);
or U4831 (N_4831,N_2011,N_2712);
nand U4832 (N_4832,N_3799,N_2940);
xnor U4833 (N_4833,N_2360,N_3342);
nor U4834 (N_4834,N_3067,N_2876);
nor U4835 (N_4835,N_2639,N_3339);
and U4836 (N_4836,N_2105,N_2722);
xnor U4837 (N_4837,N_3483,N_2910);
nand U4838 (N_4838,N_3446,N_3179);
xor U4839 (N_4839,N_2887,N_3183);
nand U4840 (N_4840,N_3837,N_2035);
or U4841 (N_4841,N_2612,N_3131);
nor U4842 (N_4842,N_3905,N_2396);
xnor U4843 (N_4843,N_2163,N_3818);
nor U4844 (N_4844,N_3434,N_2656);
nand U4845 (N_4845,N_3887,N_3226);
nor U4846 (N_4846,N_3465,N_2178);
nor U4847 (N_4847,N_3364,N_3020);
nand U4848 (N_4848,N_2469,N_2994);
nor U4849 (N_4849,N_2429,N_3812);
and U4850 (N_4850,N_2931,N_3431);
or U4851 (N_4851,N_3923,N_2184);
nor U4852 (N_4852,N_3644,N_3945);
and U4853 (N_4853,N_3396,N_2192);
nand U4854 (N_4854,N_3739,N_3572);
and U4855 (N_4855,N_2325,N_2237);
nor U4856 (N_4856,N_2751,N_3161);
xnor U4857 (N_4857,N_2880,N_2423);
nor U4858 (N_4858,N_2710,N_2912);
nor U4859 (N_4859,N_2432,N_3215);
and U4860 (N_4860,N_3629,N_2681);
xnor U4861 (N_4861,N_2422,N_2142);
and U4862 (N_4862,N_2775,N_2747);
nor U4863 (N_4863,N_2293,N_2060);
or U4864 (N_4864,N_3222,N_3485);
xor U4865 (N_4865,N_3323,N_3587);
nor U4866 (N_4866,N_2630,N_3936);
xnor U4867 (N_4867,N_3467,N_3298);
or U4868 (N_4868,N_3914,N_3642);
nand U4869 (N_4869,N_3495,N_2320);
nor U4870 (N_4870,N_3661,N_2493);
nor U4871 (N_4871,N_2252,N_2426);
and U4872 (N_4872,N_3172,N_3137);
xnor U4873 (N_4873,N_3505,N_2934);
nand U4874 (N_4874,N_3693,N_3736);
nor U4875 (N_4875,N_2215,N_2411);
and U4876 (N_4876,N_2964,N_3471);
nand U4877 (N_4877,N_2798,N_3159);
or U4878 (N_4878,N_3802,N_3075);
xnor U4879 (N_4879,N_3056,N_2349);
or U4880 (N_4880,N_3330,N_2463);
xnor U4881 (N_4881,N_3838,N_3879);
or U4882 (N_4882,N_2524,N_3925);
and U4883 (N_4883,N_3790,N_3325);
nor U4884 (N_4884,N_2860,N_2970);
nor U4885 (N_4885,N_3747,N_2572);
and U4886 (N_4886,N_3310,N_3187);
and U4887 (N_4887,N_2935,N_3751);
nand U4888 (N_4888,N_2229,N_3010);
xor U4889 (N_4889,N_2766,N_3919);
and U4890 (N_4890,N_2807,N_2869);
and U4891 (N_4891,N_3991,N_3249);
and U4892 (N_4892,N_2556,N_3047);
and U4893 (N_4893,N_2280,N_3260);
nand U4894 (N_4894,N_3610,N_2818);
or U4895 (N_4895,N_2187,N_2210);
and U4896 (N_4896,N_2767,N_2773);
or U4897 (N_4897,N_3288,N_3941);
nor U4898 (N_4898,N_3744,N_3670);
xnor U4899 (N_4899,N_2905,N_2013);
xor U4900 (N_4900,N_2913,N_3993);
nor U4901 (N_4901,N_3602,N_2626);
xnor U4902 (N_4902,N_3755,N_2963);
xnor U4903 (N_4903,N_2797,N_2357);
and U4904 (N_4904,N_3985,N_3024);
or U4905 (N_4905,N_2194,N_3583);
or U4906 (N_4906,N_2770,N_2959);
and U4907 (N_4907,N_3502,N_3869);
or U4908 (N_4908,N_2487,N_3637);
xor U4909 (N_4909,N_3247,N_3735);
nand U4910 (N_4910,N_3005,N_2580);
and U4911 (N_4911,N_2984,N_2221);
nor U4912 (N_4912,N_3386,N_2138);
and U4913 (N_4913,N_3551,N_2657);
nand U4914 (N_4914,N_3666,N_3760);
and U4915 (N_4915,N_2535,N_2790);
nand U4916 (N_4916,N_3681,N_3085);
nand U4917 (N_4917,N_3457,N_3769);
nor U4918 (N_4918,N_2009,N_2771);
xor U4919 (N_4919,N_3783,N_3646);
nand U4920 (N_4920,N_2258,N_3162);
and U4921 (N_4921,N_3455,N_2155);
xnor U4922 (N_4922,N_2618,N_3440);
nor U4923 (N_4923,N_2801,N_3106);
xor U4924 (N_4924,N_3792,N_3752);
xor U4925 (N_4925,N_2008,N_3355);
and U4926 (N_4926,N_2476,N_3588);
or U4927 (N_4927,N_2507,N_2390);
nand U4928 (N_4928,N_3041,N_2616);
or U4929 (N_4929,N_2122,N_2089);
xor U4930 (N_4930,N_3104,N_2370);
nand U4931 (N_4931,N_2135,N_3613);
nand U4932 (N_4932,N_3497,N_2919);
nor U4933 (N_4933,N_2150,N_2602);
or U4934 (N_4934,N_2039,N_3974);
nor U4935 (N_4935,N_2604,N_3858);
and U4936 (N_4936,N_3331,N_3136);
nor U4937 (N_4937,N_2428,N_3966);
or U4938 (N_4938,N_2171,N_3531);
xnor U4939 (N_4939,N_3327,N_2116);
and U4940 (N_4940,N_2528,N_3296);
xnor U4941 (N_4941,N_2660,N_2793);
nor U4942 (N_4942,N_2939,N_3449);
nor U4943 (N_4943,N_3597,N_2028);
or U4944 (N_4944,N_3207,N_2369);
or U4945 (N_4945,N_2958,N_3199);
nor U4946 (N_4946,N_3029,N_2120);
nor U4947 (N_4947,N_2704,N_3540);
nor U4948 (N_4948,N_2248,N_2031);
and U4949 (N_4949,N_3560,N_3767);
and U4950 (N_4950,N_2059,N_3781);
and U4951 (N_4951,N_2072,N_2831);
nor U4952 (N_4952,N_2567,N_2738);
nand U4953 (N_4953,N_3496,N_2062);
and U4954 (N_4954,N_3555,N_3169);
nor U4955 (N_4955,N_2562,N_2110);
xor U4956 (N_4956,N_3621,N_2987);
or U4957 (N_4957,N_2180,N_3758);
xor U4958 (N_4958,N_3775,N_2324);
nand U4959 (N_4959,N_2800,N_2095);
or U4960 (N_4960,N_2990,N_2074);
xor U4961 (N_4961,N_3883,N_3770);
nor U4962 (N_4962,N_3048,N_3141);
or U4963 (N_4963,N_3929,N_3062);
and U4964 (N_4964,N_2025,N_3934);
and U4965 (N_4965,N_2803,N_3920);
or U4966 (N_4966,N_3746,N_2795);
xor U4967 (N_4967,N_2157,N_2944);
or U4968 (N_4968,N_3907,N_3150);
nor U4969 (N_4969,N_2727,N_2253);
and U4970 (N_4970,N_3292,N_3027);
and U4971 (N_4971,N_2363,N_2570);
or U4972 (N_4972,N_2303,N_3256);
nand U4973 (N_4973,N_2774,N_2590);
nand U4974 (N_4974,N_2520,N_2755);
nand U4975 (N_4975,N_3475,N_2342);
nor U4976 (N_4976,N_2080,N_2745);
nor U4977 (N_4977,N_2853,N_3287);
and U4978 (N_4978,N_2333,N_3645);
nor U4979 (N_4979,N_2425,N_2928);
nor U4980 (N_4980,N_3017,N_3200);
and U4981 (N_4981,N_2473,N_3268);
nand U4982 (N_4982,N_3454,N_3552);
nor U4983 (N_4983,N_3192,N_3423);
nand U4984 (N_4984,N_3827,N_3115);
and U4985 (N_4985,N_2659,N_2551);
or U4986 (N_4986,N_2397,N_3143);
and U4987 (N_4987,N_3800,N_3121);
nor U4988 (N_4988,N_3703,N_2843);
nor U4989 (N_4989,N_2858,N_2702);
and U4990 (N_4990,N_2247,N_2859);
or U4991 (N_4991,N_3469,N_2094);
nor U4992 (N_4992,N_2242,N_3391);
and U4993 (N_4993,N_3623,N_2212);
nor U4994 (N_4994,N_2594,N_2043);
and U4995 (N_4995,N_3951,N_2833);
nand U4996 (N_4996,N_3392,N_3332);
nand U4997 (N_4997,N_2314,N_3080);
xor U4998 (N_4998,N_2686,N_2086);
nor U4999 (N_4999,N_3099,N_2709);
and U5000 (N_5000,N_3126,N_3387);
xor U5001 (N_5001,N_3935,N_2244);
nor U5002 (N_5002,N_2263,N_3106);
or U5003 (N_5003,N_3841,N_3225);
or U5004 (N_5004,N_2564,N_3408);
nand U5005 (N_5005,N_3322,N_2367);
and U5006 (N_5006,N_2043,N_3544);
and U5007 (N_5007,N_2102,N_3517);
xor U5008 (N_5008,N_2936,N_3583);
or U5009 (N_5009,N_2254,N_2890);
or U5010 (N_5010,N_2649,N_2106);
xnor U5011 (N_5011,N_3639,N_2317);
or U5012 (N_5012,N_3133,N_2103);
xor U5013 (N_5013,N_3149,N_3646);
xnor U5014 (N_5014,N_3381,N_2710);
or U5015 (N_5015,N_2140,N_3274);
nand U5016 (N_5016,N_2933,N_2238);
nor U5017 (N_5017,N_3043,N_3227);
nor U5018 (N_5018,N_2967,N_3963);
and U5019 (N_5019,N_2408,N_3430);
and U5020 (N_5020,N_3627,N_3862);
nor U5021 (N_5021,N_2274,N_2612);
xnor U5022 (N_5022,N_3053,N_3276);
or U5023 (N_5023,N_3912,N_3668);
and U5024 (N_5024,N_2882,N_2895);
nor U5025 (N_5025,N_3147,N_2468);
nand U5026 (N_5026,N_3907,N_3323);
xnor U5027 (N_5027,N_2352,N_3430);
xor U5028 (N_5028,N_3202,N_2132);
and U5029 (N_5029,N_2252,N_3187);
nand U5030 (N_5030,N_2810,N_2897);
and U5031 (N_5031,N_3919,N_3094);
nor U5032 (N_5032,N_2190,N_3921);
xnor U5033 (N_5033,N_2063,N_3596);
nor U5034 (N_5034,N_2118,N_2408);
nor U5035 (N_5035,N_2432,N_3590);
nand U5036 (N_5036,N_3578,N_3923);
nand U5037 (N_5037,N_2324,N_3787);
xor U5038 (N_5038,N_3613,N_3064);
nand U5039 (N_5039,N_3088,N_2279);
nand U5040 (N_5040,N_3458,N_2990);
or U5041 (N_5041,N_3600,N_2050);
nand U5042 (N_5042,N_3748,N_2553);
nand U5043 (N_5043,N_2256,N_2255);
and U5044 (N_5044,N_2414,N_3963);
nand U5045 (N_5045,N_3424,N_2276);
and U5046 (N_5046,N_3458,N_3422);
or U5047 (N_5047,N_3148,N_3940);
xnor U5048 (N_5048,N_3025,N_3322);
or U5049 (N_5049,N_2892,N_2949);
and U5050 (N_5050,N_2806,N_2983);
nand U5051 (N_5051,N_2474,N_2453);
nand U5052 (N_5052,N_2277,N_2063);
nor U5053 (N_5053,N_3796,N_2847);
or U5054 (N_5054,N_3234,N_2150);
nand U5055 (N_5055,N_3030,N_2300);
xnor U5056 (N_5056,N_2309,N_2476);
and U5057 (N_5057,N_3136,N_2601);
xor U5058 (N_5058,N_2038,N_2374);
xor U5059 (N_5059,N_2390,N_2572);
or U5060 (N_5060,N_3940,N_3939);
and U5061 (N_5061,N_3767,N_2010);
or U5062 (N_5062,N_2362,N_3343);
or U5063 (N_5063,N_2566,N_3175);
and U5064 (N_5064,N_2737,N_3834);
or U5065 (N_5065,N_2962,N_3955);
nand U5066 (N_5066,N_2304,N_2365);
and U5067 (N_5067,N_2028,N_3212);
or U5068 (N_5068,N_3623,N_3174);
or U5069 (N_5069,N_2945,N_2076);
nand U5070 (N_5070,N_2919,N_2159);
nand U5071 (N_5071,N_2260,N_3593);
nor U5072 (N_5072,N_3648,N_3691);
nand U5073 (N_5073,N_3265,N_3649);
xor U5074 (N_5074,N_2010,N_2473);
or U5075 (N_5075,N_3059,N_3190);
and U5076 (N_5076,N_3679,N_3296);
nor U5077 (N_5077,N_2278,N_2616);
xnor U5078 (N_5078,N_2487,N_2053);
nand U5079 (N_5079,N_2277,N_2982);
nand U5080 (N_5080,N_3531,N_2559);
nand U5081 (N_5081,N_3725,N_3351);
nand U5082 (N_5082,N_3414,N_3841);
nor U5083 (N_5083,N_3101,N_2670);
nand U5084 (N_5084,N_3057,N_2564);
or U5085 (N_5085,N_3306,N_2242);
or U5086 (N_5086,N_2360,N_3236);
nand U5087 (N_5087,N_3686,N_3332);
nor U5088 (N_5088,N_2018,N_3779);
nand U5089 (N_5089,N_3539,N_3805);
or U5090 (N_5090,N_2758,N_2440);
xnor U5091 (N_5091,N_2871,N_3469);
nor U5092 (N_5092,N_2836,N_2053);
and U5093 (N_5093,N_3419,N_3431);
xor U5094 (N_5094,N_3808,N_2445);
nand U5095 (N_5095,N_2080,N_3843);
and U5096 (N_5096,N_2404,N_3705);
nand U5097 (N_5097,N_2743,N_3164);
xnor U5098 (N_5098,N_3996,N_2467);
xor U5099 (N_5099,N_3026,N_3504);
xor U5100 (N_5100,N_3067,N_3389);
nor U5101 (N_5101,N_3497,N_2672);
nand U5102 (N_5102,N_2185,N_2578);
or U5103 (N_5103,N_2174,N_2195);
and U5104 (N_5104,N_3796,N_2322);
nand U5105 (N_5105,N_2946,N_3087);
or U5106 (N_5106,N_2117,N_3250);
nor U5107 (N_5107,N_3577,N_2962);
and U5108 (N_5108,N_2600,N_2971);
nor U5109 (N_5109,N_2240,N_3162);
or U5110 (N_5110,N_3309,N_3991);
and U5111 (N_5111,N_3077,N_3573);
and U5112 (N_5112,N_2178,N_2097);
xnor U5113 (N_5113,N_3063,N_3026);
xor U5114 (N_5114,N_3716,N_3677);
nor U5115 (N_5115,N_2636,N_2392);
xor U5116 (N_5116,N_3031,N_3660);
nor U5117 (N_5117,N_3490,N_3208);
nor U5118 (N_5118,N_2718,N_3602);
xnor U5119 (N_5119,N_2441,N_3054);
nand U5120 (N_5120,N_2291,N_2506);
nor U5121 (N_5121,N_2262,N_2154);
xnor U5122 (N_5122,N_2001,N_2999);
xnor U5123 (N_5123,N_3436,N_2650);
nand U5124 (N_5124,N_3039,N_3937);
nor U5125 (N_5125,N_2931,N_3256);
nor U5126 (N_5126,N_2706,N_3739);
and U5127 (N_5127,N_2280,N_3607);
and U5128 (N_5128,N_3902,N_2429);
nor U5129 (N_5129,N_3421,N_3493);
nand U5130 (N_5130,N_2837,N_2155);
or U5131 (N_5131,N_2683,N_3835);
nand U5132 (N_5132,N_2463,N_3444);
and U5133 (N_5133,N_3409,N_2517);
nor U5134 (N_5134,N_3420,N_2961);
nand U5135 (N_5135,N_3811,N_2913);
and U5136 (N_5136,N_2429,N_2794);
and U5137 (N_5137,N_2350,N_2785);
nand U5138 (N_5138,N_2331,N_3495);
or U5139 (N_5139,N_3073,N_2572);
and U5140 (N_5140,N_3410,N_2617);
nand U5141 (N_5141,N_3413,N_2463);
and U5142 (N_5142,N_2706,N_2173);
xnor U5143 (N_5143,N_2608,N_3131);
and U5144 (N_5144,N_2151,N_2231);
xnor U5145 (N_5145,N_2318,N_3809);
or U5146 (N_5146,N_3187,N_3926);
nand U5147 (N_5147,N_2808,N_2850);
xor U5148 (N_5148,N_3146,N_3297);
nand U5149 (N_5149,N_3377,N_3616);
nand U5150 (N_5150,N_3708,N_3113);
and U5151 (N_5151,N_2948,N_2980);
or U5152 (N_5152,N_2498,N_3580);
and U5153 (N_5153,N_3321,N_2114);
or U5154 (N_5154,N_3820,N_3802);
nand U5155 (N_5155,N_3768,N_3408);
and U5156 (N_5156,N_3354,N_2784);
nand U5157 (N_5157,N_3259,N_2422);
nand U5158 (N_5158,N_3528,N_2830);
nor U5159 (N_5159,N_2882,N_2858);
and U5160 (N_5160,N_3315,N_3925);
and U5161 (N_5161,N_2121,N_2171);
nand U5162 (N_5162,N_3318,N_3134);
nand U5163 (N_5163,N_3280,N_3792);
xnor U5164 (N_5164,N_2342,N_3936);
and U5165 (N_5165,N_2073,N_3666);
or U5166 (N_5166,N_2156,N_3931);
nand U5167 (N_5167,N_2815,N_2429);
and U5168 (N_5168,N_2019,N_3715);
and U5169 (N_5169,N_2516,N_3736);
nand U5170 (N_5170,N_3748,N_3553);
nand U5171 (N_5171,N_3116,N_3711);
or U5172 (N_5172,N_2373,N_2510);
or U5173 (N_5173,N_2665,N_2349);
and U5174 (N_5174,N_3544,N_2117);
nor U5175 (N_5175,N_2339,N_2438);
nand U5176 (N_5176,N_2629,N_3180);
nor U5177 (N_5177,N_3429,N_2794);
nand U5178 (N_5178,N_3621,N_3639);
or U5179 (N_5179,N_3781,N_3919);
xnor U5180 (N_5180,N_3873,N_2991);
nand U5181 (N_5181,N_2591,N_3993);
nand U5182 (N_5182,N_3742,N_2272);
nand U5183 (N_5183,N_3539,N_3316);
or U5184 (N_5184,N_3543,N_3374);
nor U5185 (N_5185,N_2458,N_2992);
nand U5186 (N_5186,N_3346,N_2683);
nor U5187 (N_5187,N_3016,N_2095);
nor U5188 (N_5188,N_3593,N_2448);
nand U5189 (N_5189,N_3461,N_3135);
nor U5190 (N_5190,N_3801,N_2767);
xor U5191 (N_5191,N_2523,N_3796);
or U5192 (N_5192,N_3941,N_2068);
and U5193 (N_5193,N_3181,N_2708);
nand U5194 (N_5194,N_2373,N_3964);
nor U5195 (N_5195,N_2058,N_2148);
nor U5196 (N_5196,N_3566,N_3409);
nand U5197 (N_5197,N_2034,N_3829);
nand U5198 (N_5198,N_2698,N_3972);
and U5199 (N_5199,N_2013,N_3554);
xnor U5200 (N_5200,N_2603,N_3944);
nor U5201 (N_5201,N_2761,N_2206);
nand U5202 (N_5202,N_3586,N_2801);
nor U5203 (N_5203,N_2443,N_2763);
xor U5204 (N_5204,N_2945,N_2260);
nand U5205 (N_5205,N_3036,N_2068);
nand U5206 (N_5206,N_3586,N_2423);
nand U5207 (N_5207,N_2071,N_3726);
or U5208 (N_5208,N_2773,N_2264);
or U5209 (N_5209,N_2743,N_2672);
xnor U5210 (N_5210,N_2869,N_3269);
xnor U5211 (N_5211,N_3715,N_2001);
xor U5212 (N_5212,N_2962,N_3861);
nor U5213 (N_5213,N_3256,N_3478);
xnor U5214 (N_5214,N_2921,N_3109);
nor U5215 (N_5215,N_2499,N_2546);
nor U5216 (N_5216,N_3587,N_2777);
nand U5217 (N_5217,N_3929,N_3653);
or U5218 (N_5218,N_2624,N_2953);
nand U5219 (N_5219,N_2853,N_2014);
xnor U5220 (N_5220,N_2374,N_3368);
or U5221 (N_5221,N_2049,N_2693);
nand U5222 (N_5222,N_2247,N_3162);
nand U5223 (N_5223,N_2478,N_2408);
xnor U5224 (N_5224,N_3238,N_2719);
nand U5225 (N_5225,N_3830,N_3818);
and U5226 (N_5226,N_2334,N_2566);
xor U5227 (N_5227,N_3926,N_2196);
nor U5228 (N_5228,N_3635,N_2213);
nand U5229 (N_5229,N_3105,N_2410);
nand U5230 (N_5230,N_2506,N_3996);
and U5231 (N_5231,N_2086,N_2497);
and U5232 (N_5232,N_2977,N_3701);
xnor U5233 (N_5233,N_2896,N_2256);
nor U5234 (N_5234,N_2215,N_2617);
or U5235 (N_5235,N_3164,N_2109);
or U5236 (N_5236,N_3035,N_2392);
xor U5237 (N_5237,N_2024,N_3060);
or U5238 (N_5238,N_3073,N_3786);
xor U5239 (N_5239,N_2298,N_3565);
and U5240 (N_5240,N_3543,N_3354);
nand U5241 (N_5241,N_2848,N_2529);
and U5242 (N_5242,N_3268,N_3010);
nand U5243 (N_5243,N_3041,N_2575);
xnor U5244 (N_5244,N_3219,N_2565);
nand U5245 (N_5245,N_2947,N_3680);
nand U5246 (N_5246,N_3543,N_3413);
xnor U5247 (N_5247,N_2938,N_3970);
and U5248 (N_5248,N_2037,N_3212);
nand U5249 (N_5249,N_3011,N_2645);
or U5250 (N_5250,N_3661,N_3995);
xnor U5251 (N_5251,N_2636,N_2208);
xor U5252 (N_5252,N_3558,N_2903);
and U5253 (N_5253,N_3731,N_3657);
nand U5254 (N_5254,N_2905,N_2260);
or U5255 (N_5255,N_2213,N_2945);
nor U5256 (N_5256,N_2673,N_2833);
nand U5257 (N_5257,N_3814,N_2371);
nor U5258 (N_5258,N_3685,N_2498);
nand U5259 (N_5259,N_3515,N_2286);
xor U5260 (N_5260,N_3994,N_2425);
and U5261 (N_5261,N_3536,N_3250);
or U5262 (N_5262,N_3183,N_2077);
or U5263 (N_5263,N_3698,N_2526);
and U5264 (N_5264,N_2731,N_3495);
nand U5265 (N_5265,N_2927,N_3999);
nor U5266 (N_5266,N_3327,N_3703);
nor U5267 (N_5267,N_3024,N_2411);
nand U5268 (N_5268,N_2282,N_2882);
or U5269 (N_5269,N_3808,N_3427);
and U5270 (N_5270,N_2128,N_2270);
and U5271 (N_5271,N_3867,N_3641);
xnor U5272 (N_5272,N_2662,N_3699);
nand U5273 (N_5273,N_3404,N_2372);
or U5274 (N_5274,N_3803,N_2340);
nand U5275 (N_5275,N_2986,N_3426);
or U5276 (N_5276,N_3021,N_3444);
and U5277 (N_5277,N_2946,N_2187);
nor U5278 (N_5278,N_3344,N_3865);
or U5279 (N_5279,N_2187,N_3963);
and U5280 (N_5280,N_2956,N_2823);
nand U5281 (N_5281,N_3599,N_2400);
or U5282 (N_5282,N_3164,N_2182);
or U5283 (N_5283,N_2391,N_3866);
nand U5284 (N_5284,N_2788,N_2978);
nand U5285 (N_5285,N_3782,N_2792);
and U5286 (N_5286,N_3717,N_3191);
or U5287 (N_5287,N_3082,N_3092);
nand U5288 (N_5288,N_3047,N_3854);
or U5289 (N_5289,N_2251,N_3198);
xnor U5290 (N_5290,N_3534,N_2850);
or U5291 (N_5291,N_3542,N_2420);
and U5292 (N_5292,N_3264,N_3325);
nor U5293 (N_5293,N_3891,N_2629);
and U5294 (N_5294,N_3297,N_3922);
or U5295 (N_5295,N_2420,N_2249);
and U5296 (N_5296,N_2631,N_2336);
and U5297 (N_5297,N_2795,N_3449);
nand U5298 (N_5298,N_2174,N_3279);
nand U5299 (N_5299,N_3655,N_3541);
and U5300 (N_5300,N_2843,N_2050);
nand U5301 (N_5301,N_2158,N_2179);
or U5302 (N_5302,N_3846,N_3561);
or U5303 (N_5303,N_2416,N_2027);
xor U5304 (N_5304,N_3587,N_3485);
xnor U5305 (N_5305,N_2468,N_2552);
or U5306 (N_5306,N_3501,N_2696);
nor U5307 (N_5307,N_2945,N_2394);
nor U5308 (N_5308,N_3496,N_2481);
and U5309 (N_5309,N_2393,N_2326);
nor U5310 (N_5310,N_3923,N_2448);
and U5311 (N_5311,N_3025,N_3738);
xor U5312 (N_5312,N_2586,N_3926);
and U5313 (N_5313,N_2890,N_2998);
and U5314 (N_5314,N_3991,N_2233);
xnor U5315 (N_5315,N_3439,N_2048);
and U5316 (N_5316,N_3599,N_3799);
nand U5317 (N_5317,N_2022,N_2212);
nor U5318 (N_5318,N_2713,N_2080);
or U5319 (N_5319,N_2070,N_2377);
nand U5320 (N_5320,N_3437,N_2804);
and U5321 (N_5321,N_3779,N_3605);
or U5322 (N_5322,N_2807,N_3920);
and U5323 (N_5323,N_2642,N_2902);
or U5324 (N_5324,N_3337,N_3415);
nand U5325 (N_5325,N_2505,N_2270);
xnor U5326 (N_5326,N_3498,N_3018);
xor U5327 (N_5327,N_3896,N_2071);
or U5328 (N_5328,N_2178,N_3620);
nand U5329 (N_5329,N_3642,N_2575);
or U5330 (N_5330,N_3687,N_2304);
and U5331 (N_5331,N_2191,N_2285);
and U5332 (N_5332,N_3089,N_3410);
nand U5333 (N_5333,N_3040,N_3551);
nor U5334 (N_5334,N_3776,N_3471);
and U5335 (N_5335,N_3637,N_2556);
and U5336 (N_5336,N_2562,N_2792);
nor U5337 (N_5337,N_3441,N_3821);
xor U5338 (N_5338,N_2700,N_2970);
xor U5339 (N_5339,N_3213,N_3729);
or U5340 (N_5340,N_3574,N_2427);
or U5341 (N_5341,N_3515,N_3154);
or U5342 (N_5342,N_2817,N_2630);
nand U5343 (N_5343,N_2619,N_2987);
and U5344 (N_5344,N_2785,N_3351);
nand U5345 (N_5345,N_3823,N_2608);
nand U5346 (N_5346,N_3453,N_3333);
and U5347 (N_5347,N_2719,N_3491);
xnor U5348 (N_5348,N_2021,N_2150);
xnor U5349 (N_5349,N_3291,N_3007);
xnor U5350 (N_5350,N_3908,N_2397);
nor U5351 (N_5351,N_2113,N_3101);
or U5352 (N_5352,N_3006,N_3598);
nor U5353 (N_5353,N_2240,N_3281);
and U5354 (N_5354,N_2174,N_2746);
or U5355 (N_5355,N_2860,N_3711);
or U5356 (N_5356,N_3241,N_2626);
nand U5357 (N_5357,N_2310,N_3654);
nor U5358 (N_5358,N_3710,N_3786);
or U5359 (N_5359,N_3668,N_3151);
nor U5360 (N_5360,N_2526,N_3751);
nor U5361 (N_5361,N_3750,N_3987);
and U5362 (N_5362,N_2881,N_3102);
or U5363 (N_5363,N_3548,N_2464);
nand U5364 (N_5364,N_2956,N_2273);
and U5365 (N_5365,N_3384,N_2717);
nor U5366 (N_5366,N_3971,N_3611);
nor U5367 (N_5367,N_3301,N_3389);
or U5368 (N_5368,N_2730,N_2395);
nor U5369 (N_5369,N_2095,N_2470);
nor U5370 (N_5370,N_3371,N_3045);
xnor U5371 (N_5371,N_2222,N_3907);
xnor U5372 (N_5372,N_2193,N_3721);
nor U5373 (N_5373,N_2470,N_2913);
xnor U5374 (N_5374,N_2683,N_2086);
xor U5375 (N_5375,N_3663,N_2866);
nor U5376 (N_5376,N_3231,N_3954);
and U5377 (N_5377,N_3089,N_2151);
nor U5378 (N_5378,N_3865,N_3906);
and U5379 (N_5379,N_2464,N_3116);
xnor U5380 (N_5380,N_2489,N_2676);
nor U5381 (N_5381,N_2904,N_2422);
nand U5382 (N_5382,N_3792,N_2783);
xor U5383 (N_5383,N_2895,N_2218);
or U5384 (N_5384,N_3958,N_2045);
nand U5385 (N_5385,N_2844,N_3425);
or U5386 (N_5386,N_3509,N_2444);
and U5387 (N_5387,N_3212,N_3267);
xor U5388 (N_5388,N_2016,N_2675);
xor U5389 (N_5389,N_3787,N_3897);
and U5390 (N_5390,N_3718,N_3023);
xor U5391 (N_5391,N_3707,N_3927);
nor U5392 (N_5392,N_2431,N_3425);
or U5393 (N_5393,N_3759,N_3645);
xor U5394 (N_5394,N_3396,N_2161);
nor U5395 (N_5395,N_2330,N_3606);
or U5396 (N_5396,N_2713,N_2946);
nand U5397 (N_5397,N_2379,N_2228);
and U5398 (N_5398,N_3801,N_3166);
nor U5399 (N_5399,N_3025,N_3082);
xor U5400 (N_5400,N_2148,N_2678);
xnor U5401 (N_5401,N_2570,N_2668);
or U5402 (N_5402,N_2474,N_3573);
and U5403 (N_5403,N_3345,N_2155);
or U5404 (N_5404,N_2560,N_2545);
nor U5405 (N_5405,N_3215,N_3076);
xnor U5406 (N_5406,N_3983,N_3080);
or U5407 (N_5407,N_3343,N_2163);
nand U5408 (N_5408,N_3123,N_2219);
and U5409 (N_5409,N_2869,N_3937);
and U5410 (N_5410,N_3117,N_2735);
nor U5411 (N_5411,N_2602,N_2853);
or U5412 (N_5412,N_2015,N_2952);
xor U5413 (N_5413,N_3312,N_2059);
or U5414 (N_5414,N_2503,N_2990);
nand U5415 (N_5415,N_2684,N_3274);
xnor U5416 (N_5416,N_2676,N_2596);
xnor U5417 (N_5417,N_3725,N_2212);
or U5418 (N_5418,N_3050,N_2055);
and U5419 (N_5419,N_3354,N_3971);
nor U5420 (N_5420,N_3669,N_3996);
nand U5421 (N_5421,N_2304,N_3542);
or U5422 (N_5422,N_2350,N_2949);
nand U5423 (N_5423,N_2853,N_2659);
nor U5424 (N_5424,N_2254,N_3094);
nor U5425 (N_5425,N_3385,N_3172);
nor U5426 (N_5426,N_3642,N_3865);
nand U5427 (N_5427,N_2938,N_2934);
nor U5428 (N_5428,N_3357,N_3973);
or U5429 (N_5429,N_2113,N_2807);
or U5430 (N_5430,N_2486,N_3916);
nor U5431 (N_5431,N_3340,N_3819);
and U5432 (N_5432,N_3481,N_3432);
or U5433 (N_5433,N_3941,N_3169);
xor U5434 (N_5434,N_2156,N_3537);
xnor U5435 (N_5435,N_2917,N_2524);
nand U5436 (N_5436,N_3861,N_2277);
xnor U5437 (N_5437,N_2890,N_3839);
nor U5438 (N_5438,N_2733,N_2231);
nor U5439 (N_5439,N_3354,N_3463);
or U5440 (N_5440,N_3610,N_3557);
nor U5441 (N_5441,N_2208,N_2321);
or U5442 (N_5442,N_2634,N_3590);
nand U5443 (N_5443,N_3740,N_3613);
xor U5444 (N_5444,N_2304,N_2584);
or U5445 (N_5445,N_3447,N_2807);
xnor U5446 (N_5446,N_3544,N_3564);
nor U5447 (N_5447,N_2883,N_3241);
or U5448 (N_5448,N_2651,N_3284);
nand U5449 (N_5449,N_3478,N_3426);
nor U5450 (N_5450,N_3668,N_2713);
and U5451 (N_5451,N_3017,N_2816);
or U5452 (N_5452,N_3463,N_2399);
or U5453 (N_5453,N_3079,N_3902);
xor U5454 (N_5454,N_2003,N_3170);
nand U5455 (N_5455,N_3935,N_2303);
nand U5456 (N_5456,N_2500,N_2000);
and U5457 (N_5457,N_3247,N_2927);
nor U5458 (N_5458,N_2873,N_2915);
or U5459 (N_5459,N_3208,N_3544);
nor U5460 (N_5460,N_3908,N_3000);
or U5461 (N_5461,N_3066,N_3919);
or U5462 (N_5462,N_3936,N_2033);
nor U5463 (N_5463,N_2792,N_3744);
or U5464 (N_5464,N_3566,N_3810);
and U5465 (N_5465,N_2236,N_2462);
or U5466 (N_5466,N_2617,N_3653);
or U5467 (N_5467,N_2494,N_3802);
or U5468 (N_5468,N_2934,N_3909);
nand U5469 (N_5469,N_3510,N_2894);
nor U5470 (N_5470,N_2554,N_3702);
and U5471 (N_5471,N_2026,N_2341);
nor U5472 (N_5472,N_2465,N_2660);
nor U5473 (N_5473,N_2929,N_2411);
and U5474 (N_5474,N_3297,N_2146);
nor U5475 (N_5475,N_3403,N_3587);
nor U5476 (N_5476,N_2055,N_2511);
nor U5477 (N_5477,N_3231,N_3377);
nand U5478 (N_5478,N_3133,N_3959);
nor U5479 (N_5479,N_3160,N_3825);
and U5480 (N_5480,N_3041,N_3093);
or U5481 (N_5481,N_2841,N_2776);
nand U5482 (N_5482,N_3790,N_2218);
xor U5483 (N_5483,N_2478,N_2020);
xnor U5484 (N_5484,N_2934,N_2164);
xnor U5485 (N_5485,N_2157,N_2461);
xnor U5486 (N_5486,N_2925,N_3093);
nand U5487 (N_5487,N_2109,N_3610);
xnor U5488 (N_5488,N_2074,N_3500);
or U5489 (N_5489,N_3526,N_2687);
xnor U5490 (N_5490,N_2602,N_3955);
and U5491 (N_5491,N_3218,N_2639);
nand U5492 (N_5492,N_3482,N_3549);
xnor U5493 (N_5493,N_2139,N_3852);
or U5494 (N_5494,N_2076,N_3738);
and U5495 (N_5495,N_2197,N_2185);
or U5496 (N_5496,N_3855,N_2838);
xnor U5497 (N_5497,N_3303,N_2239);
or U5498 (N_5498,N_3248,N_2911);
nand U5499 (N_5499,N_3889,N_2309);
nor U5500 (N_5500,N_2255,N_3561);
or U5501 (N_5501,N_2510,N_3192);
nor U5502 (N_5502,N_3657,N_2663);
xnor U5503 (N_5503,N_2520,N_2556);
and U5504 (N_5504,N_3225,N_2895);
and U5505 (N_5505,N_3548,N_2149);
nor U5506 (N_5506,N_2528,N_2020);
nor U5507 (N_5507,N_2764,N_3144);
xor U5508 (N_5508,N_3705,N_3752);
nand U5509 (N_5509,N_2219,N_3312);
xor U5510 (N_5510,N_3954,N_2992);
xor U5511 (N_5511,N_3466,N_3266);
xor U5512 (N_5512,N_3618,N_2298);
xnor U5513 (N_5513,N_3822,N_2199);
nor U5514 (N_5514,N_3540,N_2791);
or U5515 (N_5515,N_2829,N_2593);
nor U5516 (N_5516,N_3943,N_3280);
nor U5517 (N_5517,N_3997,N_2708);
nor U5518 (N_5518,N_2310,N_2203);
or U5519 (N_5519,N_2600,N_3782);
or U5520 (N_5520,N_2074,N_2820);
xnor U5521 (N_5521,N_2450,N_2721);
and U5522 (N_5522,N_2163,N_2603);
and U5523 (N_5523,N_3286,N_2428);
or U5524 (N_5524,N_3747,N_2615);
or U5525 (N_5525,N_3950,N_2258);
xnor U5526 (N_5526,N_2742,N_2160);
or U5527 (N_5527,N_3974,N_2449);
nor U5528 (N_5528,N_3996,N_3726);
nor U5529 (N_5529,N_3940,N_3096);
xnor U5530 (N_5530,N_2096,N_3101);
and U5531 (N_5531,N_2041,N_3708);
nand U5532 (N_5532,N_3829,N_2821);
or U5533 (N_5533,N_3341,N_3905);
or U5534 (N_5534,N_2787,N_3281);
nor U5535 (N_5535,N_2945,N_3608);
nor U5536 (N_5536,N_3011,N_3563);
xor U5537 (N_5537,N_2860,N_3871);
and U5538 (N_5538,N_2213,N_3934);
and U5539 (N_5539,N_2686,N_3404);
xor U5540 (N_5540,N_3868,N_3462);
xnor U5541 (N_5541,N_3169,N_3869);
nor U5542 (N_5542,N_2150,N_3831);
xor U5543 (N_5543,N_2079,N_3125);
and U5544 (N_5544,N_2067,N_2079);
xnor U5545 (N_5545,N_3993,N_2833);
or U5546 (N_5546,N_3467,N_2865);
and U5547 (N_5547,N_3520,N_2635);
nand U5548 (N_5548,N_2180,N_2195);
and U5549 (N_5549,N_3618,N_2781);
nand U5550 (N_5550,N_2395,N_3492);
or U5551 (N_5551,N_2253,N_3628);
nor U5552 (N_5552,N_3304,N_3209);
xnor U5553 (N_5553,N_2345,N_2848);
or U5554 (N_5554,N_2380,N_2401);
or U5555 (N_5555,N_3728,N_2697);
and U5556 (N_5556,N_3771,N_2763);
xor U5557 (N_5557,N_3447,N_3322);
and U5558 (N_5558,N_2832,N_2861);
nand U5559 (N_5559,N_3611,N_2441);
and U5560 (N_5560,N_2608,N_3150);
and U5561 (N_5561,N_2702,N_3559);
xnor U5562 (N_5562,N_2425,N_3063);
or U5563 (N_5563,N_2128,N_2126);
nand U5564 (N_5564,N_2706,N_2410);
nand U5565 (N_5565,N_2101,N_3322);
nand U5566 (N_5566,N_3414,N_2596);
xor U5567 (N_5567,N_3086,N_3338);
or U5568 (N_5568,N_2284,N_3724);
and U5569 (N_5569,N_3135,N_2868);
or U5570 (N_5570,N_3798,N_2448);
nor U5571 (N_5571,N_3451,N_3973);
xor U5572 (N_5572,N_3724,N_2077);
xor U5573 (N_5573,N_2181,N_2152);
nand U5574 (N_5574,N_3395,N_3697);
xnor U5575 (N_5575,N_3142,N_2907);
nand U5576 (N_5576,N_2951,N_2735);
and U5577 (N_5577,N_2213,N_3412);
nand U5578 (N_5578,N_2123,N_2949);
or U5579 (N_5579,N_3097,N_2468);
nor U5580 (N_5580,N_2561,N_3198);
nand U5581 (N_5581,N_2993,N_3293);
nor U5582 (N_5582,N_3858,N_3795);
nand U5583 (N_5583,N_2364,N_2966);
or U5584 (N_5584,N_2651,N_3980);
or U5585 (N_5585,N_3936,N_2181);
and U5586 (N_5586,N_3105,N_2526);
and U5587 (N_5587,N_3442,N_3306);
and U5588 (N_5588,N_3111,N_2543);
nor U5589 (N_5589,N_2582,N_3654);
nor U5590 (N_5590,N_2719,N_2398);
and U5591 (N_5591,N_3788,N_2547);
nor U5592 (N_5592,N_2284,N_2055);
xor U5593 (N_5593,N_3513,N_3673);
nor U5594 (N_5594,N_2999,N_2469);
or U5595 (N_5595,N_2037,N_3954);
nand U5596 (N_5596,N_3158,N_3339);
or U5597 (N_5597,N_2583,N_2599);
nor U5598 (N_5598,N_3800,N_3458);
nand U5599 (N_5599,N_2798,N_3130);
nand U5600 (N_5600,N_2158,N_2487);
and U5601 (N_5601,N_3949,N_2068);
xor U5602 (N_5602,N_2014,N_3442);
xor U5603 (N_5603,N_2983,N_2586);
or U5604 (N_5604,N_3030,N_2485);
or U5605 (N_5605,N_2797,N_2354);
nand U5606 (N_5606,N_3294,N_3305);
or U5607 (N_5607,N_2456,N_3389);
xor U5608 (N_5608,N_2772,N_2878);
and U5609 (N_5609,N_3815,N_2669);
nand U5610 (N_5610,N_3822,N_2002);
or U5611 (N_5611,N_2363,N_3756);
and U5612 (N_5612,N_2364,N_2354);
xnor U5613 (N_5613,N_3708,N_2755);
or U5614 (N_5614,N_2966,N_2773);
or U5615 (N_5615,N_3323,N_2001);
xor U5616 (N_5616,N_3595,N_3388);
nor U5617 (N_5617,N_2410,N_3161);
xnor U5618 (N_5618,N_3486,N_2636);
or U5619 (N_5619,N_2422,N_2932);
nand U5620 (N_5620,N_2833,N_3717);
xnor U5621 (N_5621,N_2320,N_3488);
or U5622 (N_5622,N_3918,N_2859);
xnor U5623 (N_5623,N_3214,N_3456);
or U5624 (N_5624,N_2628,N_3311);
xnor U5625 (N_5625,N_2406,N_3693);
nand U5626 (N_5626,N_3051,N_3599);
xor U5627 (N_5627,N_3929,N_2316);
or U5628 (N_5628,N_2829,N_2419);
or U5629 (N_5629,N_3934,N_3730);
and U5630 (N_5630,N_2391,N_3545);
nand U5631 (N_5631,N_2440,N_2983);
and U5632 (N_5632,N_2184,N_3427);
and U5633 (N_5633,N_2606,N_3742);
xor U5634 (N_5634,N_3946,N_3384);
and U5635 (N_5635,N_2955,N_3443);
xnor U5636 (N_5636,N_2855,N_3149);
nand U5637 (N_5637,N_3073,N_3916);
and U5638 (N_5638,N_2614,N_3336);
or U5639 (N_5639,N_2342,N_2063);
or U5640 (N_5640,N_2027,N_2678);
nand U5641 (N_5641,N_3451,N_3135);
nand U5642 (N_5642,N_2396,N_2854);
xnor U5643 (N_5643,N_2757,N_2652);
or U5644 (N_5644,N_2731,N_2109);
and U5645 (N_5645,N_3363,N_2678);
nand U5646 (N_5646,N_2180,N_3856);
nor U5647 (N_5647,N_3637,N_2422);
xnor U5648 (N_5648,N_2294,N_3058);
or U5649 (N_5649,N_2608,N_3170);
xnor U5650 (N_5650,N_2164,N_3345);
xor U5651 (N_5651,N_2042,N_2625);
xor U5652 (N_5652,N_3491,N_3243);
nand U5653 (N_5653,N_2254,N_2899);
xor U5654 (N_5654,N_2467,N_3404);
nor U5655 (N_5655,N_3996,N_2693);
nor U5656 (N_5656,N_2103,N_2934);
nor U5657 (N_5657,N_3430,N_3202);
nand U5658 (N_5658,N_3058,N_3783);
or U5659 (N_5659,N_2671,N_2230);
nand U5660 (N_5660,N_2285,N_2124);
xor U5661 (N_5661,N_2454,N_2211);
nand U5662 (N_5662,N_3060,N_2311);
and U5663 (N_5663,N_3808,N_2924);
and U5664 (N_5664,N_2890,N_3408);
and U5665 (N_5665,N_3535,N_3964);
and U5666 (N_5666,N_3433,N_2012);
xor U5667 (N_5667,N_2843,N_3873);
nand U5668 (N_5668,N_2005,N_3920);
nand U5669 (N_5669,N_3467,N_2592);
nand U5670 (N_5670,N_3253,N_3667);
and U5671 (N_5671,N_3699,N_3998);
or U5672 (N_5672,N_2658,N_2869);
or U5673 (N_5673,N_2315,N_2411);
or U5674 (N_5674,N_2605,N_2421);
and U5675 (N_5675,N_3846,N_3165);
and U5676 (N_5676,N_3969,N_3609);
nor U5677 (N_5677,N_3591,N_3883);
xor U5678 (N_5678,N_3840,N_3176);
or U5679 (N_5679,N_2970,N_3139);
and U5680 (N_5680,N_2170,N_3953);
xor U5681 (N_5681,N_3999,N_2191);
and U5682 (N_5682,N_2785,N_3086);
and U5683 (N_5683,N_2282,N_3322);
nor U5684 (N_5684,N_3046,N_2157);
nand U5685 (N_5685,N_2022,N_3225);
xnor U5686 (N_5686,N_2144,N_3058);
and U5687 (N_5687,N_3395,N_3806);
xor U5688 (N_5688,N_2193,N_3780);
nor U5689 (N_5689,N_2347,N_2872);
or U5690 (N_5690,N_2160,N_3640);
xor U5691 (N_5691,N_3744,N_2593);
nand U5692 (N_5692,N_2925,N_3567);
or U5693 (N_5693,N_2043,N_3591);
and U5694 (N_5694,N_3674,N_3249);
or U5695 (N_5695,N_3811,N_3014);
nand U5696 (N_5696,N_2010,N_2437);
xnor U5697 (N_5697,N_2220,N_2576);
nor U5698 (N_5698,N_2689,N_3838);
xnor U5699 (N_5699,N_2686,N_3128);
or U5700 (N_5700,N_3346,N_2721);
nand U5701 (N_5701,N_2547,N_3885);
or U5702 (N_5702,N_2580,N_2493);
and U5703 (N_5703,N_2753,N_2163);
xor U5704 (N_5704,N_2633,N_3593);
xor U5705 (N_5705,N_2217,N_2270);
or U5706 (N_5706,N_3154,N_3903);
xor U5707 (N_5707,N_2749,N_3758);
nor U5708 (N_5708,N_2699,N_3803);
xnor U5709 (N_5709,N_2459,N_2466);
xnor U5710 (N_5710,N_3835,N_2637);
nand U5711 (N_5711,N_3743,N_3951);
and U5712 (N_5712,N_2715,N_2729);
or U5713 (N_5713,N_3010,N_2744);
nor U5714 (N_5714,N_2328,N_2828);
nor U5715 (N_5715,N_3249,N_3665);
or U5716 (N_5716,N_3016,N_3059);
xor U5717 (N_5717,N_2085,N_3494);
or U5718 (N_5718,N_3788,N_3869);
xor U5719 (N_5719,N_3552,N_2674);
nor U5720 (N_5720,N_3702,N_3727);
or U5721 (N_5721,N_2559,N_2077);
or U5722 (N_5722,N_3232,N_2147);
or U5723 (N_5723,N_2175,N_2043);
xor U5724 (N_5724,N_3032,N_3202);
nor U5725 (N_5725,N_3259,N_3307);
nand U5726 (N_5726,N_2079,N_2429);
or U5727 (N_5727,N_3252,N_3537);
nor U5728 (N_5728,N_3337,N_2306);
or U5729 (N_5729,N_3680,N_3739);
and U5730 (N_5730,N_2522,N_2711);
or U5731 (N_5731,N_2348,N_2356);
and U5732 (N_5732,N_2098,N_3276);
nor U5733 (N_5733,N_3394,N_3588);
xnor U5734 (N_5734,N_2647,N_2090);
nand U5735 (N_5735,N_3490,N_2705);
nand U5736 (N_5736,N_3991,N_2447);
nand U5737 (N_5737,N_3024,N_3968);
or U5738 (N_5738,N_3170,N_2230);
nor U5739 (N_5739,N_3378,N_3627);
nand U5740 (N_5740,N_2319,N_2437);
and U5741 (N_5741,N_2018,N_2776);
xor U5742 (N_5742,N_2096,N_2944);
nand U5743 (N_5743,N_3099,N_3318);
nand U5744 (N_5744,N_3174,N_3731);
xor U5745 (N_5745,N_2946,N_2597);
nor U5746 (N_5746,N_3149,N_2956);
or U5747 (N_5747,N_2839,N_2296);
nor U5748 (N_5748,N_3723,N_3942);
nand U5749 (N_5749,N_3858,N_3275);
nor U5750 (N_5750,N_3871,N_2417);
nor U5751 (N_5751,N_2194,N_3393);
nor U5752 (N_5752,N_2968,N_2154);
nand U5753 (N_5753,N_3767,N_3612);
xnor U5754 (N_5754,N_2268,N_2328);
nor U5755 (N_5755,N_3228,N_3571);
nor U5756 (N_5756,N_2295,N_3352);
xor U5757 (N_5757,N_3159,N_2707);
nand U5758 (N_5758,N_2592,N_2981);
nor U5759 (N_5759,N_3564,N_2556);
nand U5760 (N_5760,N_3690,N_3302);
xnor U5761 (N_5761,N_2311,N_3146);
or U5762 (N_5762,N_3570,N_3671);
nand U5763 (N_5763,N_3152,N_2974);
nor U5764 (N_5764,N_3998,N_3885);
xor U5765 (N_5765,N_3196,N_2843);
nand U5766 (N_5766,N_3776,N_2331);
or U5767 (N_5767,N_2915,N_2124);
and U5768 (N_5768,N_3869,N_2508);
xor U5769 (N_5769,N_2453,N_3666);
and U5770 (N_5770,N_2751,N_2833);
nor U5771 (N_5771,N_3297,N_3200);
nand U5772 (N_5772,N_2957,N_2223);
xor U5773 (N_5773,N_2836,N_2123);
nor U5774 (N_5774,N_3735,N_2164);
or U5775 (N_5775,N_2343,N_3330);
or U5776 (N_5776,N_3932,N_3490);
or U5777 (N_5777,N_3552,N_3615);
and U5778 (N_5778,N_2052,N_2893);
and U5779 (N_5779,N_2369,N_3600);
xnor U5780 (N_5780,N_3265,N_3689);
and U5781 (N_5781,N_3075,N_3314);
xnor U5782 (N_5782,N_2555,N_3350);
xnor U5783 (N_5783,N_2016,N_3307);
nand U5784 (N_5784,N_3184,N_2784);
nand U5785 (N_5785,N_2502,N_2130);
xnor U5786 (N_5786,N_3503,N_2725);
xnor U5787 (N_5787,N_2536,N_3590);
or U5788 (N_5788,N_3392,N_2915);
xnor U5789 (N_5789,N_2773,N_3727);
nor U5790 (N_5790,N_2553,N_3596);
or U5791 (N_5791,N_3451,N_3222);
and U5792 (N_5792,N_2365,N_3689);
nand U5793 (N_5793,N_2428,N_3125);
nand U5794 (N_5794,N_3485,N_3075);
nor U5795 (N_5795,N_3807,N_2479);
and U5796 (N_5796,N_2764,N_2826);
nor U5797 (N_5797,N_2250,N_2245);
or U5798 (N_5798,N_2365,N_3380);
nand U5799 (N_5799,N_3248,N_2633);
nor U5800 (N_5800,N_3962,N_2550);
and U5801 (N_5801,N_3951,N_2557);
nand U5802 (N_5802,N_2148,N_3286);
and U5803 (N_5803,N_3062,N_2616);
or U5804 (N_5804,N_2722,N_3862);
or U5805 (N_5805,N_2677,N_3555);
nor U5806 (N_5806,N_2888,N_3180);
or U5807 (N_5807,N_2917,N_3851);
or U5808 (N_5808,N_2649,N_2150);
nor U5809 (N_5809,N_3941,N_2694);
xnor U5810 (N_5810,N_3174,N_2077);
or U5811 (N_5811,N_3242,N_3354);
and U5812 (N_5812,N_2993,N_3722);
and U5813 (N_5813,N_2905,N_2327);
and U5814 (N_5814,N_2011,N_3135);
nor U5815 (N_5815,N_3514,N_2023);
nor U5816 (N_5816,N_3831,N_2106);
or U5817 (N_5817,N_3366,N_3655);
or U5818 (N_5818,N_2792,N_3000);
xnor U5819 (N_5819,N_3132,N_2327);
and U5820 (N_5820,N_3652,N_2177);
xnor U5821 (N_5821,N_3082,N_2967);
xor U5822 (N_5822,N_3418,N_3807);
nor U5823 (N_5823,N_2709,N_3750);
nand U5824 (N_5824,N_3779,N_3472);
and U5825 (N_5825,N_2180,N_3024);
xor U5826 (N_5826,N_3227,N_2769);
or U5827 (N_5827,N_2869,N_2273);
nor U5828 (N_5828,N_3274,N_2133);
and U5829 (N_5829,N_3142,N_2719);
nand U5830 (N_5830,N_3672,N_2921);
or U5831 (N_5831,N_3392,N_3201);
or U5832 (N_5832,N_3360,N_3822);
nor U5833 (N_5833,N_3243,N_3622);
and U5834 (N_5834,N_2772,N_3519);
or U5835 (N_5835,N_3018,N_3781);
nor U5836 (N_5836,N_3970,N_2960);
xor U5837 (N_5837,N_3270,N_2872);
nor U5838 (N_5838,N_3831,N_2638);
nand U5839 (N_5839,N_3346,N_2282);
nor U5840 (N_5840,N_2111,N_2701);
xor U5841 (N_5841,N_3348,N_3533);
or U5842 (N_5842,N_3561,N_2924);
nand U5843 (N_5843,N_3413,N_3908);
and U5844 (N_5844,N_3645,N_3590);
nand U5845 (N_5845,N_3452,N_2739);
or U5846 (N_5846,N_3345,N_2875);
or U5847 (N_5847,N_3756,N_2369);
xor U5848 (N_5848,N_2264,N_3707);
or U5849 (N_5849,N_2358,N_2880);
and U5850 (N_5850,N_2517,N_2695);
xnor U5851 (N_5851,N_3709,N_3376);
or U5852 (N_5852,N_3322,N_3712);
xnor U5853 (N_5853,N_3730,N_2810);
nand U5854 (N_5854,N_2929,N_3909);
xnor U5855 (N_5855,N_3678,N_3363);
and U5856 (N_5856,N_2666,N_2383);
nor U5857 (N_5857,N_2628,N_2041);
xor U5858 (N_5858,N_3526,N_3926);
nor U5859 (N_5859,N_2020,N_2367);
nor U5860 (N_5860,N_3945,N_2620);
nand U5861 (N_5861,N_3191,N_2044);
nor U5862 (N_5862,N_2416,N_3834);
or U5863 (N_5863,N_3324,N_3894);
or U5864 (N_5864,N_3532,N_2228);
or U5865 (N_5865,N_2739,N_3418);
or U5866 (N_5866,N_2780,N_3553);
and U5867 (N_5867,N_2360,N_2194);
nand U5868 (N_5868,N_3893,N_3832);
nand U5869 (N_5869,N_2518,N_2949);
and U5870 (N_5870,N_2231,N_2953);
and U5871 (N_5871,N_2342,N_2238);
and U5872 (N_5872,N_3968,N_2742);
xnor U5873 (N_5873,N_2116,N_2375);
nor U5874 (N_5874,N_3375,N_3003);
xor U5875 (N_5875,N_3613,N_2041);
and U5876 (N_5876,N_2390,N_2312);
xnor U5877 (N_5877,N_3456,N_2146);
nand U5878 (N_5878,N_2104,N_2467);
or U5879 (N_5879,N_2065,N_2869);
nand U5880 (N_5880,N_2355,N_3155);
xnor U5881 (N_5881,N_2568,N_3532);
nor U5882 (N_5882,N_2264,N_3498);
xnor U5883 (N_5883,N_3513,N_3707);
nand U5884 (N_5884,N_2907,N_3299);
nand U5885 (N_5885,N_3657,N_3859);
and U5886 (N_5886,N_3275,N_3503);
nand U5887 (N_5887,N_3019,N_2713);
and U5888 (N_5888,N_2722,N_3813);
nand U5889 (N_5889,N_2093,N_2907);
and U5890 (N_5890,N_2187,N_3981);
nand U5891 (N_5891,N_2304,N_3208);
and U5892 (N_5892,N_3294,N_2924);
nand U5893 (N_5893,N_3185,N_2682);
nor U5894 (N_5894,N_2690,N_2262);
nor U5895 (N_5895,N_2995,N_3881);
nor U5896 (N_5896,N_2713,N_3486);
nand U5897 (N_5897,N_3371,N_2029);
or U5898 (N_5898,N_2327,N_2540);
nand U5899 (N_5899,N_3115,N_3154);
or U5900 (N_5900,N_3230,N_3440);
or U5901 (N_5901,N_3556,N_3216);
xnor U5902 (N_5902,N_3438,N_3975);
and U5903 (N_5903,N_2119,N_2568);
and U5904 (N_5904,N_3640,N_3478);
nor U5905 (N_5905,N_3134,N_2300);
or U5906 (N_5906,N_2095,N_3345);
and U5907 (N_5907,N_3055,N_3178);
xor U5908 (N_5908,N_2119,N_3963);
nand U5909 (N_5909,N_3191,N_3890);
nor U5910 (N_5910,N_2599,N_3513);
nor U5911 (N_5911,N_3861,N_2512);
xnor U5912 (N_5912,N_3548,N_2998);
xor U5913 (N_5913,N_3220,N_2298);
and U5914 (N_5914,N_2186,N_2829);
xor U5915 (N_5915,N_2354,N_2352);
nor U5916 (N_5916,N_2884,N_2217);
nand U5917 (N_5917,N_2345,N_2709);
nand U5918 (N_5918,N_3490,N_2964);
nor U5919 (N_5919,N_2381,N_2720);
nand U5920 (N_5920,N_2076,N_2422);
and U5921 (N_5921,N_2275,N_3673);
or U5922 (N_5922,N_2810,N_3616);
or U5923 (N_5923,N_2325,N_3404);
nor U5924 (N_5924,N_3595,N_3544);
nand U5925 (N_5925,N_3389,N_3922);
nand U5926 (N_5926,N_3635,N_2414);
or U5927 (N_5927,N_3143,N_3890);
xor U5928 (N_5928,N_3304,N_3555);
or U5929 (N_5929,N_3142,N_3300);
xor U5930 (N_5930,N_3931,N_2669);
nand U5931 (N_5931,N_3336,N_3793);
and U5932 (N_5932,N_3385,N_3493);
or U5933 (N_5933,N_2973,N_3842);
and U5934 (N_5934,N_3415,N_3441);
nor U5935 (N_5935,N_2562,N_2069);
nand U5936 (N_5936,N_2179,N_2044);
nand U5937 (N_5937,N_3824,N_2438);
and U5938 (N_5938,N_2850,N_2349);
nand U5939 (N_5939,N_2372,N_3851);
xor U5940 (N_5940,N_2681,N_2708);
and U5941 (N_5941,N_2129,N_2400);
or U5942 (N_5942,N_2772,N_3710);
and U5943 (N_5943,N_3692,N_3331);
nand U5944 (N_5944,N_3631,N_2371);
nor U5945 (N_5945,N_3976,N_2784);
and U5946 (N_5946,N_3095,N_3416);
nor U5947 (N_5947,N_2539,N_2589);
and U5948 (N_5948,N_3354,N_3292);
nor U5949 (N_5949,N_2103,N_2633);
nand U5950 (N_5950,N_3530,N_2503);
or U5951 (N_5951,N_3589,N_3691);
nor U5952 (N_5952,N_2894,N_3383);
and U5953 (N_5953,N_3424,N_3189);
and U5954 (N_5954,N_3304,N_2045);
or U5955 (N_5955,N_3981,N_2759);
xnor U5956 (N_5956,N_3493,N_3378);
nor U5957 (N_5957,N_3757,N_3773);
and U5958 (N_5958,N_3080,N_3519);
xnor U5959 (N_5959,N_3820,N_2852);
nor U5960 (N_5960,N_3520,N_3947);
xor U5961 (N_5961,N_3436,N_2604);
xor U5962 (N_5962,N_2217,N_2798);
nand U5963 (N_5963,N_3023,N_2370);
or U5964 (N_5964,N_2012,N_3589);
or U5965 (N_5965,N_2912,N_3545);
nor U5966 (N_5966,N_2900,N_2250);
xor U5967 (N_5967,N_3222,N_2972);
or U5968 (N_5968,N_2103,N_2346);
nand U5969 (N_5969,N_3659,N_3236);
nor U5970 (N_5970,N_2939,N_3512);
and U5971 (N_5971,N_3106,N_3565);
xnor U5972 (N_5972,N_3365,N_2539);
nor U5973 (N_5973,N_2035,N_3196);
xnor U5974 (N_5974,N_3646,N_2840);
nor U5975 (N_5975,N_2462,N_3828);
nor U5976 (N_5976,N_2863,N_3216);
or U5977 (N_5977,N_2223,N_3032);
and U5978 (N_5978,N_2962,N_3926);
nor U5979 (N_5979,N_3266,N_3587);
xnor U5980 (N_5980,N_3139,N_3046);
nor U5981 (N_5981,N_2260,N_3428);
and U5982 (N_5982,N_2491,N_2016);
or U5983 (N_5983,N_2615,N_2058);
or U5984 (N_5984,N_3803,N_2215);
and U5985 (N_5985,N_3032,N_2840);
nor U5986 (N_5986,N_2836,N_3674);
and U5987 (N_5987,N_3220,N_2817);
nand U5988 (N_5988,N_2159,N_3146);
and U5989 (N_5989,N_2911,N_3067);
xor U5990 (N_5990,N_2174,N_2380);
and U5991 (N_5991,N_3481,N_3910);
nor U5992 (N_5992,N_2127,N_2417);
xnor U5993 (N_5993,N_2196,N_3663);
nor U5994 (N_5994,N_3434,N_3355);
or U5995 (N_5995,N_3727,N_2100);
or U5996 (N_5996,N_2725,N_3666);
nor U5997 (N_5997,N_2891,N_2987);
and U5998 (N_5998,N_3125,N_3844);
and U5999 (N_5999,N_3776,N_2559);
nor U6000 (N_6000,N_4457,N_5776);
nand U6001 (N_6001,N_4514,N_4219);
and U6002 (N_6002,N_4507,N_4986);
xor U6003 (N_6003,N_4797,N_4212);
or U6004 (N_6004,N_5948,N_4948);
xnor U6005 (N_6005,N_5018,N_5637);
or U6006 (N_6006,N_4819,N_5423);
and U6007 (N_6007,N_4754,N_4297);
xnor U6008 (N_6008,N_5288,N_5428);
nand U6009 (N_6009,N_5746,N_4666);
nand U6010 (N_6010,N_5082,N_4938);
nand U6011 (N_6011,N_5411,N_5897);
nor U6012 (N_6012,N_5756,N_4305);
nor U6013 (N_6013,N_5433,N_4114);
and U6014 (N_6014,N_4195,N_4939);
nor U6015 (N_6015,N_5346,N_5753);
nor U6016 (N_6016,N_5092,N_4815);
and U6017 (N_6017,N_4509,N_4975);
xor U6018 (N_6018,N_5914,N_4989);
and U6019 (N_6019,N_4907,N_5223);
nor U6020 (N_6020,N_5761,N_4474);
and U6021 (N_6021,N_5408,N_4607);
xor U6022 (N_6022,N_5364,N_5591);
or U6023 (N_6023,N_4537,N_5241);
or U6024 (N_6024,N_5685,N_4426);
xnor U6025 (N_6025,N_5075,N_4728);
xnor U6026 (N_6026,N_4866,N_4970);
xor U6027 (N_6027,N_4544,N_4676);
xnor U6028 (N_6028,N_4804,N_4940);
nand U6029 (N_6029,N_4742,N_5515);
or U6030 (N_6030,N_4477,N_4218);
xor U6031 (N_6031,N_4364,N_4057);
or U6032 (N_6032,N_4197,N_5283);
and U6033 (N_6033,N_5448,N_4181);
xor U6034 (N_6034,N_5904,N_5202);
nand U6035 (N_6035,N_4403,N_4769);
nor U6036 (N_6036,N_4420,N_5056);
or U6037 (N_6037,N_5226,N_5099);
and U6038 (N_6038,N_5021,N_4879);
and U6039 (N_6039,N_5994,N_5706);
and U6040 (N_6040,N_4997,N_4512);
or U6041 (N_6041,N_4822,N_5522);
nor U6042 (N_6042,N_4624,N_5959);
xor U6043 (N_6043,N_4148,N_5115);
or U6044 (N_6044,N_5945,N_4686);
nand U6045 (N_6045,N_5937,N_5874);
nor U6046 (N_6046,N_4731,N_5043);
nor U6047 (N_6047,N_5870,N_4838);
nor U6048 (N_6048,N_4153,N_4683);
xor U6049 (N_6049,N_4185,N_5440);
or U6050 (N_6050,N_5422,N_4448);
nor U6051 (N_6051,N_4752,N_5758);
nor U6052 (N_6052,N_4956,N_4347);
nor U6053 (N_6053,N_5209,N_5855);
nor U6054 (N_6054,N_4740,N_5326);
or U6055 (N_6055,N_4532,N_5881);
nand U6056 (N_6056,N_5104,N_4967);
or U6057 (N_6057,N_5555,N_4851);
nor U6058 (N_6058,N_5520,N_5337);
or U6059 (N_6059,N_4178,N_5619);
xor U6060 (N_6060,N_5536,N_4928);
or U6061 (N_6061,N_4471,N_5327);
or U6062 (N_6062,N_4620,N_5788);
nand U6063 (N_6063,N_5800,N_5750);
or U6064 (N_6064,N_4700,N_5880);
nand U6065 (N_6065,N_4430,N_5675);
nand U6066 (N_6066,N_4204,N_4213);
nor U6067 (N_6067,N_4722,N_4623);
and U6068 (N_6068,N_5741,N_4035);
and U6069 (N_6069,N_4521,N_5778);
xnor U6070 (N_6070,N_5234,N_5508);
or U6071 (N_6071,N_4706,N_4168);
nor U6072 (N_6072,N_5992,N_5033);
xnor U6073 (N_6073,N_5848,N_4422);
nand U6074 (N_6074,N_5186,N_4806);
and U6075 (N_6075,N_4753,N_4406);
nand U6076 (N_6076,N_4520,N_5794);
and U6077 (N_6077,N_5576,N_5453);
nor U6078 (N_6078,N_5495,N_5653);
and U6079 (N_6079,N_4570,N_4366);
nand U6080 (N_6080,N_4652,N_5529);
or U6081 (N_6081,N_5999,N_5939);
xnor U6082 (N_6082,N_5216,N_5986);
or U6083 (N_6083,N_5055,N_5771);
and U6084 (N_6084,N_4863,N_5641);
nor U6085 (N_6085,N_5500,N_4486);
nor U6086 (N_6086,N_5872,N_5291);
or U6087 (N_6087,N_4000,N_5916);
and U6088 (N_6088,N_4857,N_5340);
nor U6089 (N_6089,N_5414,N_5492);
or U6090 (N_6090,N_4875,N_5252);
nor U6091 (N_6091,N_5182,N_5251);
nor U6092 (N_6092,N_4777,N_4590);
nor U6093 (N_6093,N_5952,N_4318);
nand U6094 (N_6094,N_4429,N_4120);
or U6095 (N_6095,N_4376,N_4184);
nand U6096 (N_6096,N_4033,N_5654);
nand U6097 (N_6097,N_4449,N_4188);
and U6098 (N_6098,N_4559,N_4782);
nor U6099 (N_6099,N_4825,N_5569);
or U6100 (N_6100,N_4858,N_5073);
nand U6101 (N_6101,N_4309,N_5832);
and U6102 (N_6102,N_5566,N_5744);
or U6103 (N_6103,N_5635,N_4393);
and U6104 (N_6104,N_4664,N_4475);
nand U6105 (N_6105,N_5452,N_5137);
nor U6106 (N_6106,N_4447,N_4598);
nor U6107 (N_6107,N_4226,N_4924);
nor U6108 (N_6108,N_4021,N_4978);
nor U6109 (N_6109,N_5413,N_5665);
or U6110 (N_6110,N_5732,N_5793);
nand U6111 (N_6111,N_4355,N_4187);
or U6112 (N_6112,N_5834,N_5757);
nor U6113 (N_6113,N_5087,N_5048);
nand U6114 (N_6114,N_4174,N_5442);
xnor U6115 (N_6115,N_5564,N_4591);
nor U6116 (N_6116,N_5909,N_5212);
or U6117 (N_6117,N_4524,N_4844);
nand U6118 (N_6118,N_5678,N_5191);
xnor U6119 (N_6119,N_4059,N_5427);
xor U6120 (N_6120,N_5072,N_4555);
or U6121 (N_6121,N_5210,N_5541);
and U6122 (N_6122,N_5405,N_5815);
nand U6123 (N_6123,N_5893,N_4601);
and U6124 (N_6124,N_5640,N_5052);
nand U6125 (N_6125,N_5380,N_5378);
nor U6126 (N_6126,N_4301,N_4217);
or U6127 (N_6127,N_5604,N_5159);
xnor U6128 (N_6128,N_4070,N_4122);
and U6129 (N_6129,N_5165,N_5543);
xnor U6130 (N_6130,N_5098,N_4008);
and U6131 (N_6131,N_4054,N_5934);
nor U6132 (N_6132,N_4126,N_5585);
nand U6133 (N_6133,N_4250,N_4760);
xor U6134 (N_6134,N_4086,N_4412);
or U6135 (N_6135,N_5016,N_4194);
nand U6136 (N_6136,N_4464,N_4599);
and U6137 (N_6137,N_4667,N_5279);
nand U6138 (N_6138,N_5203,N_5702);
or U6139 (N_6139,N_4237,N_5459);
xor U6140 (N_6140,N_5501,N_4142);
xor U6141 (N_6141,N_5605,N_4698);
xnor U6142 (N_6142,N_4738,N_5140);
nor U6143 (N_6143,N_5973,N_4024);
or U6144 (N_6144,N_4182,N_5305);
nor U6145 (N_6145,N_4784,N_5740);
or U6146 (N_6146,N_5382,N_5280);
nand U6147 (N_6147,N_4893,N_4750);
nand U6148 (N_6148,N_4583,N_4717);
nand U6149 (N_6149,N_5766,N_5467);
nand U6150 (N_6150,N_5258,N_4402);
or U6151 (N_6151,N_5828,N_5620);
and U6152 (N_6152,N_5582,N_5592);
nand U6153 (N_6153,N_4762,N_4755);
or U6154 (N_6154,N_4594,N_4563);
or U6155 (N_6155,N_5730,N_4129);
or U6156 (N_6156,N_4418,N_4751);
or U6157 (N_6157,N_5147,N_4210);
nor U6158 (N_6158,N_5603,N_5805);
nor U6159 (N_6159,N_5972,N_5105);
nor U6160 (N_6160,N_5735,N_4534);
xnor U6161 (N_6161,N_5906,N_5601);
nand U6162 (N_6162,N_5636,N_4677);
nand U6163 (N_6163,N_5174,N_5630);
and U6164 (N_6164,N_5248,N_5008);
nand U6165 (N_6165,N_5519,N_4660);
xor U6166 (N_6166,N_4543,N_4873);
nand U6167 (N_6167,N_4074,N_5726);
nand U6168 (N_6168,N_4358,N_4159);
nand U6169 (N_6169,N_4209,N_5662);
or U6170 (N_6170,N_5957,N_5720);
or U6171 (N_6171,N_5797,N_4820);
nor U6172 (N_6172,N_4973,N_5511);
or U6173 (N_6173,N_4643,N_5849);
nand U6174 (N_6174,N_4650,N_4348);
and U6175 (N_6175,N_5229,N_4431);
and U6176 (N_6176,N_4006,N_4915);
nand U6177 (N_6177,N_5814,N_5377);
and U6178 (N_6178,N_5613,N_5692);
or U6179 (N_6179,N_5618,N_5712);
and U6180 (N_6180,N_5518,N_4561);
xnor U6181 (N_6181,N_5739,N_5928);
nor U6182 (N_6182,N_5704,N_5786);
nor U6183 (N_6183,N_5693,N_5953);
xnor U6184 (N_6184,N_5371,N_4971);
nor U6185 (N_6185,N_5141,N_5804);
or U6186 (N_6186,N_5527,N_5158);
nor U6187 (N_6187,N_4236,N_5397);
or U6188 (N_6188,N_5336,N_5782);
or U6189 (N_6189,N_4580,N_4719);
xor U6190 (N_6190,N_4143,N_5486);
or U6191 (N_6191,N_4007,N_5045);
nand U6192 (N_6192,N_4979,N_4200);
nand U6193 (N_6193,N_5911,N_5851);
xor U6194 (N_6194,N_5818,N_5319);
nor U6195 (N_6195,N_5193,N_4966);
nor U6196 (N_6196,N_4627,N_5850);
or U6197 (N_6197,N_4491,N_5164);
and U6198 (N_6198,N_5224,N_5717);
nand U6199 (N_6199,N_5360,N_4399);
and U6200 (N_6200,N_4028,N_5974);
nor U6201 (N_6201,N_5830,N_5854);
nor U6202 (N_6202,N_4397,N_4949);
nand U6203 (N_6203,N_5121,N_4988);
or U6204 (N_6204,N_4106,N_4465);
or U6205 (N_6205,N_5597,N_4541);
or U6206 (N_6206,N_4029,N_4339);
nor U6207 (N_6207,N_5131,N_5331);
nor U6208 (N_6208,N_5609,N_5009);
nand U6209 (N_6209,N_4014,N_5571);
nand U6210 (N_6210,N_5839,N_4302);
or U6211 (N_6211,N_4852,N_4190);
nor U6212 (N_6212,N_5051,N_5760);
nand U6213 (N_6213,N_4186,N_4617);
or U6214 (N_6214,N_4425,N_4155);
and U6215 (N_6215,N_5910,N_5544);
nand U6216 (N_6216,N_4082,N_4937);
nand U6217 (N_6217,N_4846,N_4703);
xor U6218 (N_6218,N_5296,N_4665);
and U6219 (N_6219,N_5088,N_5367);
xor U6220 (N_6220,N_5892,N_4482);
nand U6221 (N_6221,N_4638,N_5109);
or U6222 (N_6222,N_4952,N_5533);
and U6223 (N_6223,N_4729,N_5157);
or U6224 (N_6224,N_5769,N_5304);
or U6225 (N_6225,N_4062,N_5882);
nand U6226 (N_6226,N_5311,N_5456);
and U6227 (N_6227,N_4351,N_4454);
nand U6228 (N_6228,N_5049,N_4786);
and U6229 (N_6229,N_5328,N_5058);
and U6230 (N_6230,N_4523,N_5956);
or U6231 (N_6231,N_5431,N_4380);
nand U6232 (N_6232,N_5494,N_4201);
or U6233 (N_6233,N_4388,N_4001);
xnor U6234 (N_6234,N_4162,N_4642);
nor U6235 (N_6235,N_4778,N_4368);
nor U6236 (N_6236,N_4298,N_5531);
or U6237 (N_6237,N_4307,N_4352);
or U6238 (N_6238,N_4295,N_4055);
xor U6239 (N_6239,N_5035,N_5833);
and U6240 (N_6240,N_5310,N_4243);
and U6241 (N_6241,N_5868,N_4890);
and U6242 (N_6242,N_5517,N_4073);
xnor U6243 (N_6243,N_5153,N_4494);
nand U6244 (N_6244,N_4828,N_5196);
or U6245 (N_6245,N_5824,N_5388);
xnor U6246 (N_6246,N_5698,N_4342);
or U6247 (N_6247,N_4639,N_5689);
xor U6248 (N_6248,N_4827,N_4883);
xor U6249 (N_6249,N_5107,N_4690);
or U6250 (N_6250,N_5922,N_5984);
or U6251 (N_6251,N_5149,N_5138);
nor U6252 (N_6252,N_5097,N_5172);
xnor U6253 (N_6253,N_5211,N_4562);
xor U6254 (N_6254,N_4748,N_4249);
nand U6255 (N_6255,N_4096,N_4487);
nand U6256 (N_6256,N_5747,N_5436);
or U6257 (N_6257,N_4897,N_5374);
and U6258 (N_6258,N_4012,N_4221);
or U6259 (N_6259,N_4987,N_5985);
nand U6260 (N_6260,N_4771,N_5264);
or U6261 (N_6261,N_5743,N_5703);
xnor U6262 (N_6262,N_5837,N_4049);
nor U6263 (N_6263,N_5350,N_4904);
xor U6264 (N_6264,N_5709,N_5711);
nor U6265 (N_6265,N_4177,N_4668);
nor U6266 (N_6266,N_5923,N_5053);
nor U6267 (N_6267,N_5345,N_4687);
xnor U6268 (N_6268,N_5425,N_5568);
or U6269 (N_6269,N_5315,N_4409);
nand U6270 (N_6270,N_4341,N_5444);
or U6271 (N_6271,N_4203,N_5130);
nand U6272 (N_6272,N_4892,N_5989);
nor U6273 (N_6273,N_4957,N_4790);
and U6274 (N_6274,N_4291,N_5488);
nand U6275 (N_6275,N_5490,N_4060);
xor U6276 (N_6276,N_4821,N_4392);
nand U6277 (N_6277,N_4536,N_5602);
xnor U6278 (N_6278,N_4444,N_5590);
nand U6279 (N_6279,N_4548,N_4985);
nor U6280 (N_6280,N_5243,N_5451);
or U6281 (N_6281,N_5086,N_5156);
or U6282 (N_6282,N_4041,N_5574);
nor U6283 (N_6283,N_5316,N_5421);
nor U6284 (N_6284,N_4003,N_5335);
and U6285 (N_6285,N_5827,N_4993);
nand U6286 (N_6286,N_4066,N_4228);
xor U6287 (N_6287,N_5809,N_5022);
xnor U6288 (N_6288,N_5161,N_4972);
xnor U6289 (N_6289,N_5466,N_5545);
or U6290 (N_6290,N_5046,N_4075);
xor U6291 (N_6291,N_5355,N_5188);
nor U6292 (N_6292,N_4635,N_5250);
and U6293 (N_6293,N_4472,N_4888);
or U6294 (N_6294,N_4708,N_5132);
xnor U6295 (N_6295,N_5729,N_4776);
nor U6296 (N_6296,N_4357,N_4493);
nand U6297 (N_6297,N_4315,N_4092);
nand U6298 (N_6298,N_5863,N_4572);
nor U6299 (N_6299,N_5721,N_5417);
or U6300 (N_6300,N_4269,N_4390);
or U6301 (N_6301,N_5287,N_4108);
and U6302 (N_6302,N_5190,N_5951);
or U6303 (N_6303,N_4552,N_4905);
or U6304 (N_6304,N_4946,N_5622);
nor U6305 (N_6305,N_5866,N_5903);
nand U6306 (N_6306,N_4871,N_5458);
nand U6307 (N_6307,N_4467,N_4490);
xnor U6308 (N_6308,N_5633,N_5476);
nor U6309 (N_6309,N_4522,N_5700);
and U6310 (N_6310,N_4775,N_5943);
nand U6311 (N_6311,N_5399,N_4485);
or U6312 (N_6312,N_4914,N_5240);
nor U6313 (N_6313,N_4688,N_5347);
or U6314 (N_6314,N_5068,N_5742);
nand U6315 (N_6315,N_5817,N_5171);
xor U6316 (N_6316,N_5370,N_5435);
and U6317 (N_6317,N_4146,N_4027);
nand U6318 (N_6318,N_4878,N_5179);
or U6319 (N_6319,N_4774,N_4816);
xor U6320 (N_6320,N_4763,N_4785);
nor U6321 (N_6321,N_5710,N_5323);
nor U6322 (N_6322,N_4919,N_5713);
and U6323 (N_6323,N_5524,N_5840);
nand U6324 (N_6324,N_5219,N_4943);
nor U6325 (N_6325,N_4255,N_5067);
xnor U6326 (N_6326,N_4304,N_4078);
nor U6327 (N_6327,N_5135,N_4282);
nand U6328 (N_6328,N_4176,N_5811);
and U6329 (N_6329,N_5737,N_5256);
nor U6330 (N_6330,N_5783,N_4196);
nand U6331 (N_6331,N_5807,N_4648);
or U6332 (N_6332,N_4408,N_5332);
or U6333 (N_6333,N_5607,N_4363);
nor U6334 (N_6334,N_5204,N_4272);
or U6335 (N_6335,N_4280,N_4980);
nand U6336 (N_6336,N_4216,N_4932);
and U6337 (N_6337,N_5168,N_5542);
nand U6338 (N_6338,N_4983,N_4245);
xor U6339 (N_6339,N_5375,N_5728);
or U6340 (N_6340,N_4047,N_4225);
and U6341 (N_6341,N_4959,N_4423);
nor U6342 (N_6342,N_5557,N_4323);
nand U6343 (N_6343,N_5192,N_4343);
nor U6344 (N_6344,N_4587,N_4415);
nand U6345 (N_6345,N_5719,N_5480);
or U6346 (N_6346,N_4894,N_5026);
or U6347 (N_6347,N_5499,N_5962);
and U6348 (N_6348,N_5349,N_5651);
and U6349 (N_6349,N_4606,N_4414);
or U6350 (N_6350,N_4991,N_5813);
nand U6351 (N_6351,N_5773,N_4720);
nor U6352 (N_6352,N_4571,N_4670);
or U6353 (N_6353,N_4505,N_4835);
and U6354 (N_6354,N_5077,N_4626);
nand U6355 (N_6355,N_5669,N_5074);
xor U6356 (N_6356,N_4749,N_4726);
and U6357 (N_6357,N_5981,N_4446);
nand U6358 (N_6358,N_4103,N_5979);
nand U6359 (N_6359,N_5676,N_5586);
or U6360 (N_6360,N_5487,N_4084);
xor U6361 (N_6361,N_5100,N_5460);
and U6362 (N_6362,N_4829,N_5801);
and U6363 (N_6363,N_5019,N_4040);
and U6364 (N_6364,N_4499,N_4123);
and U6365 (N_6365,N_5069,N_5852);
nand U6366 (N_6366,N_4920,N_5667);
or U6367 (N_6367,N_4109,N_4325);
nand U6368 (N_6368,N_4547,N_5129);
or U6369 (N_6369,N_4313,N_4818);
and U6370 (N_6370,N_4709,N_5372);
nor U6371 (N_6371,N_5781,N_5514);
nand U6372 (N_6372,N_4300,N_5942);
xnor U6373 (N_6373,N_4276,N_5695);
xor U6374 (N_6374,N_4018,N_5434);
and U6375 (N_6375,N_5247,N_5078);
nand U6376 (N_6376,N_4337,N_4419);
xor U6377 (N_6377,N_4134,N_4546);
nor U6378 (N_6378,N_4179,N_4533);
nor U6379 (N_6379,N_5755,N_4005);
or U6380 (N_6380,N_4634,N_4922);
nand U6381 (N_6381,N_4809,N_4525);
nand U6382 (N_6382,N_5201,N_5464);
nand U6383 (N_6383,N_5356,N_5023);
xor U6384 (N_6384,N_5883,N_5173);
xnor U6385 (N_6385,N_4372,N_4649);
or U6386 (N_6386,N_5905,N_4947);
nor U6387 (N_6387,N_5816,N_4288);
nor U6388 (N_6388,N_5477,N_5503);
and U6389 (N_6389,N_4359,N_5206);
nor U6390 (N_6390,N_4768,N_4923);
or U6391 (N_6391,N_4868,N_4538);
nand U6392 (N_6392,N_4068,N_4274);
xnor U6393 (N_6393,N_4792,N_4141);
nand U6394 (N_6394,N_5232,N_5856);
or U6395 (N_6395,N_5111,N_5961);
and U6396 (N_6396,N_4805,N_4721);
nor U6397 (N_6397,N_4759,N_5510);
and U6398 (N_6398,N_5385,N_4810);
nor U6399 (N_6399,N_5090,N_5220);
xor U6400 (N_6400,N_5825,N_5627);
nand U6401 (N_6401,N_4091,N_5913);
xor U6402 (N_6402,N_4680,N_4167);
xnor U6403 (N_6403,N_4646,N_4421);
nor U6404 (N_6404,N_5277,N_4540);
xor U6405 (N_6405,N_5221,N_5102);
nor U6406 (N_6406,N_4707,N_5632);
or U6407 (N_6407,N_5313,N_5964);
and U6408 (N_6408,N_4672,N_5617);
xor U6409 (N_6409,N_5736,N_5420);
xor U6410 (N_6410,N_5393,N_5474);
nor U6411 (N_6411,N_5123,N_5955);
nand U6412 (N_6412,N_5154,N_4745);
and U6413 (N_6413,N_4737,N_5738);
xnor U6414 (N_6414,N_5977,N_4331);
or U6415 (N_6415,N_5844,N_4231);
nand U6416 (N_6416,N_5643,N_4856);
xor U6417 (N_6417,N_4568,N_4299);
and U6418 (N_6418,N_5039,N_4861);
nor U6419 (N_6419,N_5608,N_4906);
xor U6420 (N_6420,N_5249,N_5772);
and U6421 (N_6421,N_5389,N_4279);
nand U6422 (N_6422,N_4385,N_4371);
nand U6423 (N_6423,N_4974,N_4597);
nor U6424 (N_6424,N_5938,N_5845);
xnor U6425 (N_6425,N_4595,N_4503);
or U6426 (N_6426,N_5924,N_4391);
and U6427 (N_6427,N_4814,N_4038);
nand U6428 (N_6428,N_5255,N_4773);
xnor U6429 (N_6429,N_4602,N_4675);
nand U6430 (N_6430,N_5160,N_5506);
and U6431 (N_6431,N_5341,N_5344);
xnor U6432 (N_6432,N_4618,N_5185);
xor U6433 (N_6433,N_5749,N_5321);
and U6434 (N_6434,N_5236,N_4310);
xor U6435 (N_6435,N_4381,N_4992);
or U6436 (N_6436,N_5847,N_4247);
nor U6437 (N_6437,N_5152,N_4389);
or U6438 (N_6438,N_5473,N_5925);
nand U6439 (N_6439,N_5301,N_5081);
or U6440 (N_6440,N_5644,N_5183);
nand U6441 (N_6441,N_5180,N_4910);
nand U6442 (N_6442,N_5200,N_4767);
nor U6443 (N_6443,N_4616,N_5638);
nor U6444 (N_6444,N_4895,N_4193);
and U6445 (N_6445,N_4138,N_5290);
nor U6446 (N_6446,N_4410,N_5207);
and U6447 (N_6447,N_5812,N_5461);
nand U6448 (N_6448,N_4631,N_5767);
or U6449 (N_6449,N_4977,N_4679);
or U6450 (N_6450,N_4515,N_5418);
or U6451 (N_6451,N_5261,N_5862);
or U6452 (N_6452,N_5365,N_4294);
nand U6453 (N_6453,N_4461,N_4743);
nand U6454 (N_6454,N_4211,N_4206);
or U6455 (N_6455,N_4744,N_4424);
or U6456 (N_6456,N_4527,N_5861);
xor U6457 (N_6457,N_4115,N_4799);
and U6458 (N_6458,N_5752,N_4896);
xor U6459 (N_6459,N_4135,N_4741);
and U6460 (N_6460,N_5199,N_5819);
or U6461 (N_6461,N_5274,N_5929);
and U6462 (N_6462,N_5314,N_5696);
and U6463 (N_6463,N_5976,N_4151);
xor U6464 (N_6464,N_5386,N_5062);
nor U6465 (N_6465,N_4518,N_5113);
nand U6466 (N_6466,N_5886,N_5106);
xor U6467 (N_6467,N_4127,N_5409);
and U6468 (N_6468,N_4052,N_4281);
or U6469 (N_6469,N_4320,N_5539);
nand U6470 (N_6470,N_4612,N_4953);
xnor U6471 (N_6471,N_4880,N_5468);
or U6472 (N_6472,N_4043,N_5538);
and U6473 (N_6473,N_4781,N_5795);
and U6474 (N_6474,N_4031,N_5502);
nand U6475 (N_6475,N_5128,N_4470);
nand U6476 (N_6476,N_5975,N_4887);
nand U6477 (N_6477,N_5231,N_5358);
xnor U6478 (N_6478,N_5670,N_5649);
xnor U6479 (N_6479,N_4849,N_4042);
xnor U6480 (N_6480,N_4229,N_4899);
and U6481 (N_6481,N_5765,N_4715);
nor U6482 (N_6482,N_4723,N_5610);
or U6483 (N_6483,N_4629,N_5491);
nor U6484 (N_6484,N_4519,N_5338);
and U6485 (N_6485,N_4145,N_5921);
nor U6486 (N_6486,N_5278,N_5228);
xnor U6487 (N_6487,N_4198,N_4479);
nand U6488 (N_6488,N_5083,N_5554);
nor U6489 (N_6489,N_4160,N_4098);
nand U6490 (N_6490,N_4224,N_4968);
and U6491 (N_6491,N_5927,N_4716);
nor U6492 (N_6492,N_4289,N_4625);
and U6493 (N_6493,N_5133,N_4508);
xnor U6494 (N_6494,N_4417,N_4692);
xor U6495 (N_6495,N_5257,N_4874);
and U6496 (N_6496,N_5064,N_5679);
and U6497 (N_6497,N_5213,N_4584);
nand U6498 (N_6498,N_4466,N_4076);
or U6499 (N_6499,N_5139,N_4063);
xor U6500 (N_6500,N_4659,N_5426);
and U6501 (N_6501,N_5446,N_4296);
nor U6502 (N_6502,N_4733,N_5112);
and U6503 (N_6503,N_4656,N_4316);
xnor U6504 (N_6504,N_4758,N_4962);
and U6505 (N_6505,N_5733,N_5563);
or U6506 (N_6506,N_4175,N_5798);
xnor U6507 (N_6507,N_4094,N_5791);
nor U6508 (N_6508,N_5122,N_4710);
or U6509 (N_6509,N_4131,N_5065);
and U6510 (N_6510,N_4222,N_5189);
xor U6511 (N_6511,N_5918,N_4292);
nor U6512 (N_6512,N_4684,N_5917);
xnor U6513 (N_6513,N_4002,N_5658);
nor U6514 (N_6514,N_4253,N_4862);
xor U6515 (N_6515,N_4287,N_5803);
or U6516 (N_6516,N_5616,N_4085);
and U6517 (N_6517,N_5307,N_5003);
nand U6518 (N_6518,N_5070,N_5898);
and U6519 (N_6519,N_5400,N_5671);
or U6520 (N_6520,N_4689,N_5177);
nor U6521 (N_6521,N_5483,N_5908);
or U6522 (N_6522,N_4439,N_5659);
and U6523 (N_6523,N_5691,N_5263);
and U6524 (N_6524,N_5664,N_4395);
or U6525 (N_6525,N_5672,N_4800);
nand U6526 (N_6526,N_4982,N_5978);
nor U6527 (N_6527,N_5784,N_5876);
and U6528 (N_6528,N_4484,N_4925);
xnor U6529 (N_6529,N_5329,N_4845);
and U6530 (N_6530,N_4192,N_4020);
nor U6531 (N_6531,N_4916,N_4233);
nor U6532 (N_6532,N_4855,N_4370);
nor U6533 (N_6533,N_4104,N_4277);
or U6534 (N_6534,N_4244,N_5657);
nor U6535 (N_6535,N_5325,N_4811);
xnor U6536 (N_6536,N_5621,N_4263);
nand U6537 (N_6537,N_5899,N_4564);
nand U6538 (N_6538,N_4165,N_4576);
nor U6539 (N_6539,N_4791,N_5724);
nor U6540 (N_6540,N_5050,N_5036);
nor U6541 (N_6541,N_5103,N_4902);
xnor U6542 (N_6542,N_5686,N_5965);
and U6543 (N_6543,N_4869,N_4132);
nor U6544 (N_6544,N_4889,N_4711);
and U6545 (N_6545,N_4739,N_4876);
nor U6546 (N_6546,N_5373,N_5178);
nand U6547 (N_6547,N_4171,N_5958);
nand U6548 (N_6548,N_4645,N_4614);
or U6549 (N_6549,N_4958,N_4251);
xor U6550 (N_6550,N_5683,N_4156);
and U6551 (N_6551,N_4839,N_4090);
or U6552 (N_6552,N_5233,N_5652);
and U6553 (N_6553,N_4268,N_5663);
nand U6554 (N_6554,N_5674,N_4099);
nand U6555 (N_6555,N_4927,N_5991);
nor U6556 (N_6556,N_5155,N_5528);
xor U6557 (N_6557,N_4859,N_5395);
or U6558 (N_6558,N_5725,N_4398);
xor U6559 (N_6559,N_5935,N_4051);
nand U6560 (N_6560,N_5504,N_5915);
nand U6561 (N_6561,N_4332,N_5877);
nor U6562 (N_6562,N_4262,N_4511);
nand U6563 (N_6563,N_4585,N_4111);
nand U6564 (N_6564,N_4833,N_5013);
and U6565 (N_6565,N_4516,N_4933);
and U6566 (N_6566,N_4473,N_5521);
nand U6567 (N_6567,N_5887,N_5846);
and U6568 (N_6568,N_5581,N_4560);
nor U6569 (N_6569,N_4384,N_5628);
xor U6570 (N_6570,N_5919,N_4207);
nand U6571 (N_6571,N_5996,N_4275);
nand U6572 (N_6572,N_4764,N_5754);
or U6573 (N_6573,N_5465,N_5034);
nor U6574 (N_6574,N_5842,N_4694);
nor U6575 (N_6575,N_4630,N_4961);
nand U6576 (N_6576,N_5276,N_4954);
or U6577 (N_6577,N_5281,N_5303);
or U6578 (N_6578,N_4912,N_4865);
xor U6579 (N_6579,N_4427,N_5163);
and U6580 (N_6580,N_4458,N_4841);
nor U6581 (N_6581,N_5745,N_5215);
or U6582 (N_6582,N_5768,N_4998);
nand U6583 (N_6583,N_5297,N_4565);
xnor U6584 (N_6584,N_5478,N_4658);
or U6585 (N_6585,N_4019,N_5029);
xnor U6586 (N_6586,N_4330,N_5246);
and U6587 (N_6587,N_5785,N_5869);
nand U6588 (N_6588,N_4673,N_4346);
xnor U6589 (N_6589,N_4586,N_5673);
or U6590 (N_6590,N_5432,N_5507);
xnor U6591 (N_6591,N_4045,N_5963);
or U6592 (N_6592,N_4152,N_5450);
nand U6593 (N_6593,N_5025,N_5266);
nor U6594 (N_6594,N_4695,N_5513);
and U6595 (N_6595,N_4401,N_5967);
and U6596 (N_6596,N_5823,N_5789);
nand U6597 (N_6597,N_4433,N_5573);
or U6598 (N_6598,N_4747,N_5988);
and U6599 (N_6599,N_4260,N_5454);
and U6600 (N_6600,N_5612,N_4154);
xnor U6601 (N_6601,N_4671,N_4377);
nor U6602 (N_6602,N_5968,N_4539);
and U6603 (N_6603,N_4238,N_5512);
nand U6604 (N_6604,N_5888,N_5265);
or U6605 (N_6605,N_5143,N_5998);
and U6606 (N_6606,N_5273,N_5006);
nand U6607 (N_6607,N_5176,N_4095);
nand U6608 (N_6608,N_5108,N_4202);
or U6609 (N_6609,N_5150,N_4022);
xnor U6610 (N_6610,N_5879,N_5751);
nand U6611 (N_6611,N_5799,N_4647);
nor U6612 (N_6612,N_5089,N_5391);
xor U6613 (N_6613,N_5596,N_5639);
xnor U6614 (N_6614,N_5714,N_4886);
and U6615 (N_6615,N_4173,N_4550);
xor U6616 (N_6616,N_4557,N_4794);
nand U6617 (N_6617,N_4469,N_5493);
or U6618 (N_6618,N_5394,N_4901);
nand U6619 (N_6619,N_4405,N_5871);
or U6620 (N_6620,N_4633,N_5320);
nand U6621 (N_6621,N_4267,N_4622);
or U6622 (N_6622,N_4964,N_5552);
and U6623 (N_6623,N_5194,N_4817);
or U6624 (N_6624,N_5534,N_4502);
or U6625 (N_6625,N_4191,N_5699);
and U6626 (N_6626,N_5390,N_5770);
nor U6627 (N_6627,N_4831,N_5116);
nor U6628 (N_6628,N_5443,N_4394);
or U6629 (N_6629,N_4340,N_5227);
or U6630 (N_6630,N_4009,N_5010);
nor U6631 (N_6631,N_5293,N_5600);
nand U6632 (N_6632,N_4452,N_4459);
nor U6633 (N_6633,N_5169,N_4746);
nand U6634 (N_6634,N_4592,N_4147);
xor U6635 (N_6635,N_5646,N_5060);
nand U6636 (N_6636,N_5629,N_4283);
and U6637 (N_6637,N_4034,N_4365);
xnor U6638 (N_6638,N_4678,N_4918);
nand U6639 (N_6639,N_4528,N_4725);
or U6640 (N_6640,N_5983,N_4199);
xnor U6641 (N_6641,N_4116,N_4801);
xnor U6642 (N_6642,N_5101,N_5110);
xor U6643 (N_6643,N_4312,N_5406);
and U6644 (N_6644,N_5148,N_4504);
nand U6645 (N_6645,N_4079,N_5271);
nor U6646 (N_6646,N_5595,N_5032);
nor U6647 (N_6647,N_4483,N_5860);
nand U6648 (N_6648,N_5864,N_5439);
nor U6649 (N_6649,N_4780,N_4712);
nor U6650 (N_6650,N_4387,N_5343);
nor U6651 (N_6651,N_5599,N_4701);
xor U6652 (N_6652,N_4266,N_4496);
xnor U6653 (N_6653,N_4354,N_4900);
nand U6654 (N_6654,N_5498,N_4566);
and U6655 (N_6655,N_4662,N_5170);
or U6656 (N_6656,N_5063,N_5526);
xor U6657 (N_6657,N_4558,N_5810);
nand U6658 (N_6658,N_4220,N_4913);
nor U6659 (N_6659,N_4327,N_4898);
or U6660 (N_6660,N_5059,N_5626);
nor U6661 (N_6661,N_5634,N_4969);
nand U6662 (N_6662,N_4010,N_4999);
or U6663 (N_6663,N_5885,N_5334);
xnor U6664 (N_6664,N_4303,N_5763);
nor U6665 (N_6665,N_4015,N_4061);
and U6666 (N_6666,N_5895,N_4329);
and U6667 (N_6667,N_4468,N_5438);
or U6668 (N_6668,N_5368,N_4577);
xor U6669 (N_6669,N_5836,N_4832);
xnor U6670 (N_6670,N_4161,N_5469);
nand U6671 (N_6671,N_4089,N_5875);
xor U6672 (N_6672,N_4117,N_5701);
and U6673 (N_6673,N_4926,N_4437);
nand U6674 (N_6674,N_5270,N_5214);
and U6675 (N_6675,N_5884,N_5858);
or U6676 (N_6676,N_5615,N_5677);
nand U6677 (N_6677,N_4338,N_4336);
nand U6678 (N_6678,N_4489,N_4230);
and U6679 (N_6679,N_4549,N_4942);
nor U6680 (N_6680,N_5031,N_5080);
and U6681 (N_6681,N_5530,N_4013);
nor U6682 (N_6682,N_5449,N_4872);
and U6683 (N_6683,N_5748,N_4789);
or U6684 (N_6684,N_4450,N_4367);
nand U6685 (N_6685,N_4124,N_4356);
and U6686 (N_6686,N_5462,N_4362);
or U6687 (N_6687,N_4691,N_4088);
and U6688 (N_6688,N_5235,N_5404);
or U6689 (N_6689,N_4110,N_5120);
and U6690 (N_6690,N_4682,N_4651);
or U6691 (N_6691,N_4453,N_5625);
xnor U6692 (N_6692,N_4609,N_4882);
nand U6693 (N_6693,N_5392,N_4573);
xnor U6694 (N_6694,N_5057,N_4802);
nor U6695 (N_6695,N_5339,N_4628);
and U6696 (N_6696,N_4637,N_4037);
xor U6697 (N_6697,N_5230,N_4102);
or U6698 (N_6698,N_4319,N_5481);
xnor U6699 (N_6699,N_4257,N_5218);
xor U6700 (N_6700,N_4840,N_4588);
and U6701 (N_6701,N_5949,N_4101);
and U6702 (N_6702,N_4107,N_5285);
nor U6703 (N_6703,N_5777,N_5482);
and U6704 (N_6704,N_5873,N_4083);
nor U6705 (N_6705,N_4663,N_5412);
and U6706 (N_6706,N_5642,N_5516);
nand U6707 (N_6707,N_5987,N_5550);
nor U6708 (N_6708,N_5071,N_4644);
or U6709 (N_6709,N_5167,N_4077);
or U6710 (N_6710,N_5484,N_5125);
and U6711 (N_6711,N_4344,N_5902);
nand U6712 (N_6712,N_4478,N_4166);
nand U6713 (N_6713,N_5145,N_5594);
nand U6714 (N_6714,N_5966,N_4158);
xnor U6715 (N_6715,N_4046,N_5037);
and U6716 (N_6716,N_5041,N_4039);
xnor U6717 (N_6717,N_5993,N_5079);
xor U6718 (N_6718,N_4130,N_5429);
and U6719 (N_6719,N_4259,N_5437);
nor U6720 (N_6720,N_5085,N_5997);
xnor U6721 (N_6721,N_4480,N_5790);
or U6722 (N_6722,N_4067,N_5723);
or U6723 (N_6723,N_5308,N_4333);
nor U6724 (N_6724,N_5020,N_5680);
and U6725 (N_6725,N_4596,N_4456);
and U6726 (N_6726,N_4308,N_4205);
nand U6727 (N_6727,N_5244,N_4843);
nand U6728 (N_6728,N_5859,N_4349);
or U6729 (N_6729,N_4125,N_4657);
or U6730 (N_6730,N_4556,N_5472);
nand U6731 (N_6731,N_5831,N_5727);
xor U6732 (N_6732,N_5187,N_4965);
xnor U6733 (N_6733,N_4891,N_5294);
and U6734 (N_6734,N_4379,N_4854);
xor U6735 (N_6735,N_5969,N_4944);
nor U6736 (N_6736,N_4242,N_4383);
xnor U6737 (N_6737,N_5166,N_4517);
xnor U6738 (N_6738,N_5286,N_4984);
nor U6739 (N_6739,N_5118,N_5584);
and U6740 (N_6740,N_4326,N_4133);
nand U6741 (N_6741,N_5901,N_4837);
nor U6742 (N_6742,N_4870,N_5558);
nand U6743 (N_6743,N_4779,N_5471);
and U6744 (N_6744,N_5260,N_4234);
and U6745 (N_6745,N_4261,N_5697);
and U6746 (N_6746,N_4172,N_5061);
nor U6747 (N_6747,N_4121,N_5284);
nor U6748 (N_6748,N_4069,N_5361);
xor U6749 (N_6749,N_4438,N_5357);
and U6750 (N_6750,N_4736,N_4436);
nor U6751 (N_6751,N_5546,N_4795);
and U6752 (N_6752,N_5445,N_5990);
nor U6753 (N_6753,N_5559,N_4441);
nand U6754 (N_6754,N_4498,N_4462);
and U6755 (N_6755,N_5694,N_4921);
or U6756 (N_6756,N_5455,N_5759);
or U6757 (N_6757,N_4432,N_5195);
nand U6758 (N_6758,N_5366,N_5655);
and U6759 (N_6759,N_4834,N_4693);
xnor U6760 (N_6760,N_5403,N_4796);
or U6761 (N_6761,N_5030,N_5017);
nand U6762 (N_6762,N_4705,N_4286);
and U6763 (N_6763,N_4072,N_5878);
nand U6764 (N_6764,N_4065,N_4285);
nand U6765 (N_6765,N_5066,N_4492);
nand U6766 (N_6766,N_5575,N_5716);
nor U6767 (N_6767,N_4730,N_4793);
nor U6768 (N_6768,N_4334,N_4306);
xnor U6769 (N_6769,N_5774,N_5525);
nand U6770 (N_6770,N_5684,N_4945);
nand U6771 (N_6771,N_4252,N_4271);
xnor U6772 (N_6772,N_4050,N_4375);
nand U6773 (N_6773,N_4575,N_5117);
nand U6774 (N_6774,N_5096,N_5567);
nand U6775 (N_6775,N_5463,N_5342);
nand U6776 (N_6776,N_5982,N_4113);
nor U6777 (N_6777,N_5136,N_5532);
and U6778 (N_6778,N_4278,N_4488);
nor U6779 (N_6779,N_5926,N_4345);
xnor U6780 (N_6780,N_5907,N_5764);
nand U6781 (N_6781,N_5457,N_5920);
xnor U6782 (N_6782,N_4569,N_5647);
or U6783 (N_6783,N_4995,N_4321);
or U6784 (N_6784,N_4080,N_4081);
or U6785 (N_6785,N_5004,N_4885);
or U6786 (N_6786,N_4322,N_4128);
nor U6787 (N_6787,N_4600,N_5940);
and U6788 (N_6788,N_5094,N_5205);
nor U6789 (N_6789,N_4284,N_4163);
and U6790 (N_6790,N_4807,N_4144);
and U6791 (N_6791,N_4150,N_5047);
xnor U6792 (N_6792,N_5587,N_4981);
xnor U6793 (N_6793,N_4823,N_5282);
or U6794 (N_6794,N_4661,N_5668);
nor U6795 (N_6795,N_5623,N_5262);
nand U6796 (N_6796,N_5042,N_4017);
and U6797 (N_6797,N_4254,N_5707);
nor U6798 (N_6798,N_4976,N_4118);
nor U6799 (N_6799,N_5867,N_5401);
or U6800 (N_6800,N_4311,N_5820);
nand U6801 (N_6801,N_5889,N_5645);
and U6802 (N_6802,N_4501,N_5424);
xnor U6803 (N_6803,N_4579,N_4772);
nand U6804 (N_6804,N_5447,N_5275);
nand U6805 (N_6805,N_4783,N_5000);
nor U6806 (N_6806,N_5298,N_4613);
and U6807 (N_6807,N_4654,N_4481);
xnor U6808 (N_6808,N_4451,N_4058);
and U6809 (N_6809,N_5091,N_4463);
and U6810 (N_6810,N_4044,N_5217);
xnor U6811 (N_6811,N_4223,N_5324);
or U6812 (N_6812,N_5577,N_4542);
xnor U6813 (N_6813,N_5843,N_5731);
nor U6814 (N_6814,N_4936,N_4328);
xnor U6815 (N_6815,N_4030,N_4697);
nand U6816 (N_6816,N_5802,N_5624);
or U6817 (N_6817,N_5208,N_5479);
nand U6818 (N_6818,N_4713,N_5475);
nand U6819 (N_6819,N_4770,N_5690);
nand U6820 (N_6820,N_5396,N_4554);
and U6821 (N_6821,N_4093,N_5441);
nand U6822 (N_6822,N_5722,N_5162);
or U6823 (N_6823,N_4813,N_4189);
nor U6824 (N_6824,N_4026,N_4004);
xnor U6825 (N_6825,N_4836,N_4324);
or U6826 (N_6826,N_4445,N_5238);
or U6827 (N_6827,N_4374,N_4714);
xor U6828 (N_6828,N_5362,N_5496);
or U6829 (N_6829,N_5775,N_4407);
nor U6830 (N_6830,N_5001,N_4903);
nor U6831 (N_6831,N_5095,N_5359);
or U6832 (N_6832,N_4053,N_4112);
and U6833 (N_6833,N_4669,N_4350);
xnor U6834 (N_6834,N_5762,N_5853);
nor U6835 (N_6835,N_5470,N_5292);
and U6836 (N_6836,N_5225,N_5354);
nand U6837 (N_6837,N_4265,N_4137);
or U6838 (N_6838,N_5708,N_4619);
nand U6839 (N_6839,N_5896,N_5588);
xor U6840 (N_6840,N_4064,N_4963);
and U6841 (N_6841,N_5718,N_5317);
nor U6842 (N_6842,N_5259,N_5253);
nand U6843 (N_6843,N_5578,N_5309);
nor U6844 (N_6844,N_5779,N_5835);
nand U6845 (N_6845,N_5027,N_4950);
nand U6846 (N_6846,N_4413,N_5239);
or U6847 (N_6847,N_5146,N_5272);
or U6848 (N_6848,N_5254,N_4674);
and U6849 (N_6849,N_5681,N_4574);
or U6850 (N_6850,N_5944,N_4757);
and U6851 (N_6851,N_4908,N_4732);
nor U6852 (N_6852,N_4023,N_4442);
xnor U6853 (N_6853,N_4960,N_5363);
nand U6854 (N_6854,N_4353,N_5330);
nor U6855 (N_6855,N_5144,N_4955);
nor U6856 (N_6856,N_5549,N_5142);
and U6857 (N_6857,N_4551,N_5666);
xnor U6858 (N_6858,N_4361,N_5093);
and U6859 (N_6859,N_4139,N_5302);
nor U6860 (N_6860,N_5489,N_5631);
or U6861 (N_6861,N_5351,N_4610);
and U6862 (N_6862,N_4756,N_5841);
and U6863 (N_6863,N_4848,N_4264);
nand U6864 (N_6864,N_5570,N_4632);
nand U6865 (N_6865,N_5682,N_5995);
or U6866 (N_6866,N_5379,N_4812);
xor U6867 (N_6867,N_4808,N_5044);
and U6868 (N_6868,N_5237,N_4164);
nand U6869 (N_6869,N_5197,N_4860);
nor U6870 (N_6870,N_4235,N_5941);
or U6871 (N_6871,N_5787,N_4830);
nor U6872 (N_6872,N_4495,N_4685);
and U6873 (N_6873,N_5583,N_5054);
and U6874 (N_6874,N_4611,N_4699);
and U6875 (N_6875,N_5005,N_5119);
or U6876 (N_6876,N_4105,N_4884);
nand U6877 (N_6877,N_5971,N_4246);
nor U6878 (N_6878,N_5333,N_5548);
nor U6879 (N_6879,N_5381,N_5611);
nor U6880 (N_6880,N_4929,N_5808);
nand U6881 (N_6881,N_5579,N_4718);
xor U6882 (N_6882,N_5383,N_4149);
and U6883 (N_6883,N_5430,N_5269);
nor U6884 (N_6884,N_4593,N_5306);
or U6885 (N_6885,N_4608,N_4119);
xor U6886 (N_6886,N_5865,N_4136);
nand U6887 (N_6887,N_4476,N_5410);
xor U6888 (N_6888,N_5407,N_4214);
or U6889 (N_6889,N_4787,N_4881);
and U6890 (N_6890,N_5648,N_4317);
and U6891 (N_6891,N_5792,N_4208);
nand U6892 (N_6892,N_5181,N_4788);
and U6893 (N_6893,N_5384,N_4853);
xnor U6894 (N_6894,N_5560,N_5126);
nor U6895 (N_6895,N_5402,N_5299);
nand U6896 (N_6896,N_4455,N_4911);
xor U6897 (N_6897,N_5012,N_4850);
nand U6898 (N_6898,N_4724,N_4909);
nand U6899 (N_6899,N_5589,N_5821);
nor U6900 (N_6900,N_5606,N_4605);
nand U6901 (N_6901,N_4513,N_4867);
and U6902 (N_6902,N_4655,N_4056);
nand U6903 (N_6903,N_4727,N_5289);
and U6904 (N_6904,N_5954,N_4766);
nor U6905 (N_6905,N_5040,N_4256);
nor U6906 (N_6906,N_4378,N_5705);
nor U6907 (N_6907,N_5134,N_4404);
and U6908 (N_6908,N_4290,N_4140);
nand U6909 (N_6909,N_5024,N_5348);
and U6910 (N_6910,N_5505,N_4553);
nor U6911 (N_6911,N_5890,N_4183);
xnor U6912 (N_6912,N_5715,N_5485);
nand U6913 (N_6913,N_4702,N_5980);
nand U6914 (N_6914,N_4097,N_5387);
xor U6915 (N_6915,N_5198,N_5509);
nor U6916 (N_6916,N_5734,N_4510);
nor U6917 (N_6917,N_4400,N_5572);
nand U6918 (N_6918,N_4545,N_4036);
xnor U6919 (N_6919,N_5523,N_5780);
nand U6920 (N_6920,N_5838,N_4396);
nand U6921 (N_6921,N_5561,N_4435);
or U6922 (N_6922,N_5084,N_4798);
nor U6923 (N_6923,N_5826,N_4931);
and U6924 (N_6924,N_4087,N_5222);
and U6925 (N_6925,N_4877,N_5946);
nand U6926 (N_6926,N_5556,N_4994);
xnor U6927 (N_6927,N_5540,N_4239);
or U6928 (N_6928,N_5950,N_4460);
nor U6929 (N_6929,N_4258,N_4360);
or U6930 (N_6930,N_5933,N_4636);
xor U6931 (N_6931,N_4864,N_4293);
xor U6932 (N_6932,N_5661,N_5295);
nor U6933 (N_6933,N_5076,N_5398);
xor U6934 (N_6934,N_5127,N_5614);
or U6935 (N_6935,N_5598,N_4603);
nand U6936 (N_6936,N_4416,N_4011);
nor U6937 (N_6937,N_5415,N_4842);
and U6938 (N_6938,N_4930,N_4373);
or U6939 (N_6939,N_5322,N_4640);
and U6940 (N_6940,N_4578,N_5932);
or U6941 (N_6941,N_4100,N_5245);
xnor U6942 (N_6942,N_5376,N_4232);
nor U6943 (N_6943,N_5822,N_4335);
or U6944 (N_6944,N_4434,N_4615);
xor U6945 (N_6945,N_4696,N_4428);
xnor U6946 (N_6946,N_5151,N_5416);
and U6947 (N_6947,N_4529,N_5537);
nand U6948 (N_6948,N_4734,N_4535);
and U6949 (N_6949,N_4025,N_4589);
nand U6950 (N_6950,N_4273,N_4016);
nor U6951 (N_6951,N_4996,N_5947);
nand U6952 (N_6952,N_4582,N_4526);
xnor U6953 (N_6953,N_5930,N_4531);
nor U6954 (N_6954,N_4735,N_5497);
nand U6955 (N_6955,N_5267,N_4382);
nand U6956 (N_6956,N_5353,N_5551);
xnor U6957 (N_6957,N_5806,N_5931);
or U6958 (N_6958,N_4847,N_5007);
or U6959 (N_6959,N_4641,N_5015);
xor U6960 (N_6960,N_4826,N_4621);
or U6961 (N_6961,N_4314,N_4951);
xor U6962 (N_6962,N_5565,N_5660);
nand U6963 (N_6963,N_5936,N_4248);
and U6964 (N_6964,N_4215,N_5894);
nor U6965 (N_6965,N_5891,N_4934);
xor U6966 (N_6966,N_5562,N_5796);
nand U6967 (N_6967,N_4803,N_5547);
and U6968 (N_6968,N_5312,N_4581);
nor U6969 (N_6969,N_4048,N_5900);
xor U6970 (N_6970,N_5650,N_4990);
nor U6971 (N_6971,N_4157,N_4824);
nor U6972 (N_6972,N_5184,N_5268);
and U6973 (N_6973,N_5175,N_4180);
xor U6974 (N_6974,N_4506,N_5242);
xnor U6975 (N_6975,N_5960,N_5656);
or U6976 (N_6976,N_4241,N_5002);
nand U6977 (N_6977,N_5419,N_4604);
nor U6978 (N_6978,N_4169,N_4032);
or U6979 (N_6979,N_5028,N_4071);
nand U6980 (N_6980,N_5011,N_4500);
and U6981 (N_6981,N_4227,N_5369);
nand U6982 (N_6982,N_4704,N_5687);
nand U6983 (N_6983,N_5857,N_4765);
nand U6984 (N_6984,N_4653,N_4270);
nor U6985 (N_6985,N_4567,N_4369);
nand U6986 (N_6986,N_5300,N_4170);
nor U6987 (N_6987,N_4411,N_4530);
xnor U6988 (N_6988,N_5970,N_4497);
and U6989 (N_6989,N_5038,N_4917);
xnor U6990 (N_6990,N_4681,N_5580);
xor U6991 (N_6991,N_5352,N_5912);
and U6992 (N_6992,N_5114,N_4443);
nand U6993 (N_6993,N_4935,N_5124);
or U6994 (N_6994,N_5688,N_4240);
and U6995 (N_6995,N_5318,N_5553);
nand U6996 (N_6996,N_5829,N_4941);
or U6997 (N_6997,N_4761,N_5593);
or U6998 (N_6998,N_4386,N_5535);
nand U6999 (N_6999,N_4440,N_5014);
and U7000 (N_7000,N_4376,N_4907);
xor U7001 (N_7001,N_5105,N_5755);
or U7002 (N_7002,N_5950,N_4337);
nor U7003 (N_7003,N_5141,N_5196);
nor U7004 (N_7004,N_5326,N_5707);
and U7005 (N_7005,N_5477,N_4172);
xnor U7006 (N_7006,N_4690,N_4144);
xnor U7007 (N_7007,N_5050,N_4855);
and U7008 (N_7008,N_5407,N_4308);
nor U7009 (N_7009,N_5484,N_5375);
and U7010 (N_7010,N_4077,N_4487);
and U7011 (N_7011,N_5584,N_5974);
nor U7012 (N_7012,N_5087,N_5098);
nor U7013 (N_7013,N_5815,N_5385);
xor U7014 (N_7014,N_5285,N_4473);
nor U7015 (N_7015,N_5933,N_4234);
nor U7016 (N_7016,N_4221,N_4333);
or U7017 (N_7017,N_5823,N_5965);
and U7018 (N_7018,N_5600,N_5758);
xnor U7019 (N_7019,N_4609,N_4860);
and U7020 (N_7020,N_4162,N_5981);
or U7021 (N_7021,N_4494,N_5691);
nand U7022 (N_7022,N_4108,N_5555);
nand U7023 (N_7023,N_5083,N_5609);
nand U7024 (N_7024,N_5639,N_4725);
or U7025 (N_7025,N_4692,N_4217);
nand U7026 (N_7026,N_5778,N_5576);
and U7027 (N_7027,N_5614,N_4519);
nand U7028 (N_7028,N_4460,N_5549);
or U7029 (N_7029,N_4337,N_4040);
and U7030 (N_7030,N_4028,N_4119);
xor U7031 (N_7031,N_4138,N_4810);
nor U7032 (N_7032,N_4379,N_5148);
xor U7033 (N_7033,N_4379,N_5835);
xnor U7034 (N_7034,N_5940,N_5641);
and U7035 (N_7035,N_5840,N_4164);
nor U7036 (N_7036,N_4827,N_4308);
xnor U7037 (N_7037,N_4822,N_4092);
or U7038 (N_7038,N_5928,N_5506);
xor U7039 (N_7039,N_5319,N_4738);
or U7040 (N_7040,N_4430,N_5040);
and U7041 (N_7041,N_4334,N_5205);
xor U7042 (N_7042,N_4887,N_5133);
nand U7043 (N_7043,N_4817,N_4712);
or U7044 (N_7044,N_5947,N_5034);
nand U7045 (N_7045,N_4820,N_5221);
nor U7046 (N_7046,N_5723,N_5034);
and U7047 (N_7047,N_5633,N_5630);
and U7048 (N_7048,N_5258,N_4717);
or U7049 (N_7049,N_4064,N_4351);
and U7050 (N_7050,N_5504,N_5569);
nor U7051 (N_7051,N_5307,N_4122);
nor U7052 (N_7052,N_4228,N_4036);
xnor U7053 (N_7053,N_4690,N_4937);
nor U7054 (N_7054,N_5789,N_4560);
xnor U7055 (N_7055,N_4555,N_4900);
nand U7056 (N_7056,N_5296,N_5790);
xnor U7057 (N_7057,N_5923,N_5302);
nand U7058 (N_7058,N_4056,N_4895);
nand U7059 (N_7059,N_4850,N_5727);
nor U7060 (N_7060,N_4673,N_4504);
or U7061 (N_7061,N_5372,N_5550);
and U7062 (N_7062,N_4254,N_4001);
nand U7063 (N_7063,N_5948,N_4196);
and U7064 (N_7064,N_4707,N_4034);
xnor U7065 (N_7065,N_5394,N_5785);
or U7066 (N_7066,N_4682,N_5413);
nor U7067 (N_7067,N_4690,N_5650);
or U7068 (N_7068,N_5222,N_5845);
xnor U7069 (N_7069,N_5831,N_4958);
xor U7070 (N_7070,N_4853,N_5217);
nand U7071 (N_7071,N_5097,N_5183);
xor U7072 (N_7072,N_5120,N_4641);
or U7073 (N_7073,N_5092,N_4764);
and U7074 (N_7074,N_5097,N_5710);
nor U7075 (N_7075,N_5096,N_5358);
nor U7076 (N_7076,N_5142,N_4011);
nor U7077 (N_7077,N_4927,N_4691);
xnor U7078 (N_7078,N_5798,N_4505);
or U7079 (N_7079,N_5902,N_5286);
or U7080 (N_7080,N_5646,N_5626);
xor U7081 (N_7081,N_4234,N_5992);
xnor U7082 (N_7082,N_4474,N_5148);
and U7083 (N_7083,N_4722,N_4993);
or U7084 (N_7084,N_4086,N_4671);
and U7085 (N_7085,N_5513,N_5742);
nor U7086 (N_7086,N_5282,N_5487);
or U7087 (N_7087,N_4175,N_5871);
nor U7088 (N_7088,N_5092,N_4156);
nor U7089 (N_7089,N_5325,N_5920);
or U7090 (N_7090,N_5288,N_5113);
nor U7091 (N_7091,N_4309,N_4134);
xnor U7092 (N_7092,N_5034,N_4821);
nand U7093 (N_7093,N_5463,N_4445);
or U7094 (N_7094,N_4668,N_4980);
nor U7095 (N_7095,N_5770,N_4868);
nor U7096 (N_7096,N_5730,N_5233);
or U7097 (N_7097,N_5856,N_4430);
nand U7098 (N_7098,N_4601,N_5364);
and U7099 (N_7099,N_4066,N_4216);
xnor U7100 (N_7100,N_4923,N_4396);
nand U7101 (N_7101,N_4823,N_4266);
or U7102 (N_7102,N_5207,N_4003);
and U7103 (N_7103,N_4197,N_4074);
and U7104 (N_7104,N_5341,N_5502);
nor U7105 (N_7105,N_5594,N_5999);
or U7106 (N_7106,N_5440,N_5421);
and U7107 (N_7107,N_5397,N_4232);
and U7108 (N_7108,N_5906,N_5199);
xnor U7109 (N_7109,N_5848,N_4458);
and U7110 (N_7110,N_5403,N_5326);
or U7111 (N_7111,N_5850,N_4108);
or U7112 (N_7112,N_4784,N_4901);
xnor U7113 (N_7113,N_5841,N_5024);
nand U7114 (N_7114,N_5272,N_4636);
nand U7115 (N_7115,N_4997,N_5940);
nand U7116 (N_7116,N_4964,N_4492);
xor U7117 (N_7117,N_4461,N_5399);
and U7118 (N_7118,N_5563,N_4094);
nand U7119 (N_7119,N_5184,N_4529);
xor U7120 (N_7120,N_4055,N_5679);
xnor U7121 (N_7121,N_5638,N_5443);
nor U7122 (N_7122,N_5213,N_4992);
nor U7123 (N_7123,N_4593,N_5126);
and U7124 (N_7124,N_4403,N_5948);
xor U7125 (N_7125,N_4417,N_4523);
and U7126 (N_7126,N_5608,N_5381);
or U7127 (N_7127,N_5470,N_4050);
nor U7128 (N_7128,N_5220,N_4342);
and U7129 (N_7129,N_5769,N_4283);
and U7130 (N_7130,N_4150,N_5471);
or U7131 (N_7131,N_5586,N_4563);
nand U7132 (N_7132,N_4877,N_4390);
or U7133 (N_7133,N_4474,N_5540);
or U7134 (N_7134,N_4457,N_4007);
nand U7135 (N_7135,N_4244,N_5880);
nand U7136 (N_7136,N_4592,N_4009);
and U7137 (N_7137,N_5014,N_4076);
and U7138 (N_7138,N_5173,N_4426);
and U7139 (N_7139,N_4942,N_5376);
nor U7140 (N_7140,N_5799,N_4033);
or U7141 (N_7141,N_4879,N_4195);
nor U7142 (N_7142,N_4706,N_4165);
nor U7143 (N_7143,N_5261,N_5212);
xnor U7144 (N_7144,N_5437,N_5765);
or U7145 (N_7145,N_4737,N_4003);
or U7146 (N_7146,N_5057,N_4124);
xor U7147 (N_7147,N_4301,N_5736);
xor U7148 (N_7148,N_4156,N_5489);
nand U7149 (N_7149,N_5625,N_5959);
or U7150 (N_7150,N_5126,N_5158);
or U7151 (N_7151,N_4164,N_5093);
nor U7152 (N_7152,N_4443,N_4063);
and U7153 (N_7153,N_4650,N_4927);
or U7154 (N_7154,N_4127,N_5429);
or U7155 (N_7155,N_5257,N_5141);
xnor U7156 (N_7156,N_5392,N_5914);
or U7157 (N_7157,N_5452,N_4713);
nand U7158 (N_7158,N_5031,N_4839);
and U7159 (N_7159,N_5602,N_5725);
or U7160 (N_7160,N_4525,N_5345);
and U7161 (N_7161,N_4249,N_5213);
nand U7162 (N_7162,N_5992,N_5252);
xnor U7163 (N_7163,N_5879,N_4233);
nor U7164 (N_7164,N_4381,N_5469);
xnor U7165 (N_7165,N_4983,N_4641);
nor U7166 (N_7166,N_4716,N_5734);
xor U7167 (N_7167,N_5620,N_4901);
xor U7168 (N_7168,N_5349,N_4026);
xor U7169 (N_7169,N_4692,N_5887);
or U7170 (N_7170,N_4905,N_4559);
nand U7171 (N_7171,N_5609,N_5826);
nand U7172 (N_7172,N_5037,N_5503);
or U7173 (N_7173,N_4603,N_5822);
or U7174 (N_7174,N_4054,N_4331);
and U7175 (N_7175,N_4015,N_4428);
and U7176 (N_7176,N_4876,N_5679);
xor U7177 (N_7177,N_5614,N_4388);
and U7178 (N_7178,N_5084,N_5049);
nor U7179 (N_7179,N_5716,N_4429);
nand U7180 (N_7180,N_5832,N_4373);
and U7181 (N_7181,N_5837,N_4933);
or U7182 (N_7182,N_5960,N_5669);
xor U7183 (N_7183,N_4102,N_4478);
and U7184 (N_7184,N_5206,N_5550);
nand U7185 (N_7185,N_5445,N_4050);
and U7186 (N_7186,N_4030,N_4382);
or U7187 (N_7187,N_5159,N_5271);
xor U7188 (N_7188,N_5048,N_5076);
xnor U7189 (N_7189,N_5944,N_4112);
nor U7190 (N_7190,N_5840,N_4026);
and U7191 (N_7191,N_5879,N_5439);
nand U7192 (N_7192,N_5283,N_5394);
xnor U7193 (N_7193,N_5804,N_4125);
or U7194 (N_7194,N_4161,N_4168);
nand U7195 (N_7195,N_4626,N_4949);
nor U7196 (N_7196,N_4537,N_5617);
nor U7197 (N_7197,N_4113,N_4766);
and U7198 (N_7198,N_5714,N_4442);
nand U7199 (N_7199,N_5582,N_4812);
xnor U7200 (N_7200,N_4165,N_4128);
nand U7201 (N_7201,N_4412,N_5430);
nor U7202 (N_7202,N_5480,N_5696);
xnor U7203 (N_7203,N_5740,N_5056);
or U7204 (N_7204,N_5182,N_5136);
nand U7205 (N_7205,N_5340,N_5898);
nor U7206 (N_7206,N_4407,N_4883);
nor U7207 (N_7207,N_5217,N_5911);
xor U7208 (N_7208,N_5436,N_5859);
or U7209 (N_7209,N_4436,N_5077);
nor U7210 (N_7210,N_4443,N_4320);
nor U7211 (N_7211,N_4269,N_5405);
xnor U7212 (N_7212,N_5104,N_4495);
nand U7213 (N_7213,N_4226,N_4662);
nand U7214 (N_7214,N_5128,N_4177);
and U7215 (N_7215,N_5864,N_4713);
and U7216 (N_7216,N_5959,N_5285);
or U7217 (N_7217,N_5657,N_5740);
and U7218 (N_7218,N_4815,N_5982);
or U7219 (N_7219,N_5586,N_4243);
nor U7220 (N_7220,N_5734,N_4852);
nor U7221 (N_7221,N_4249,N_5251);
xnor U7222 (N_7222,N_5660,N_4015);
nor U7223 (N_7223,N_5317,N_5710);
nand U7224 (N_7224,N_4423,N_4911);
and U7225 (N_7225,N_4235,N_5815);
xnor U7226 (N_7226,N_4650,N_4716);
or U7227 (N_7227,N_4424,N_4560);
or U7228 (N_7228,N_5883,N_5659);
nor U7229 (N_7229,N_5315,N_5181);
and U7230 (N_7230,N_5138,N_5323);
or U7231 (N_7231,N_5235,N_4390);
nor U7232 (N_7232,N_4886,N_5914);
and U7233 (N_7233,N_5747,N_4218);
xnor U7234 (N_7234,N_4619,N_5389);
nor U7235 (N_7235,N_5571,N_5130);
and U7236 (N_7236,N_5660,N_5960);
xor U7237 (N_7237,N_5101,N_5901);
nor U7238 (N_7238,N_5098,N_4690);
or U7239 (N_7239,N_5698,N_4668);
and U7240 (N_7240,N_4831,N_4904);
and U7241 (N_7241,N_4239,N_5568);
nand U7242 (N_7242,N_4499,N_4965);
nor U7243 (N_7243,N_5049,N_4172);
xnor U7244 (N_7244,N_5985,N_4762);
and U7245 (N_7245,N_5247,N_4207);
and U7246 (N_7246,N_4379,N_5217);
or U7247 (N_7247,N_5226,N_5807);
and U7248 (N_7248,N_4383,N_5685);
nand U7249 (N_7249,N_4349,N_5023);
xor U7250 (N_7250,N_5420,N_5621);
nand U7251 (N_7251,N_4910,N_5985);
nor U7252 (N_7252,N_4532,N_4987);
and U7253 (N_7253,N_4628,N_5214);
nor U7254 (N_7254,N_4278,N_5245);
xnor U7255 (N_7255,N_5129,N_5362);
xor U7256 (N_7256,N_4089,N_5386);
or U7257 (N_7257,N_4198,N_5398);
nor U7258 (N_7258,N_4002,N_5196);
nand U7259 (N_7259,N_4113,N_4081);
nand U7260 (N_7260,N_4244,N_5396);
nor U7261 (N_7261,N_4445,N_4305);
nand U7262 (N_7262,N_5069,N_5697);
xnor U7263 (N_7263,N_4654,N_5108);
nand U7264 (N_7264,N_5498,N_4479);
nor U7265 (N_7265,N_4547,N_4653);
nand U7266 (N_7266,N_5375,N_5547);
nand U7267 (N_7267,N_5428,N_5821);
or U7268 (N_7268,N_4493,N_5289);
and U7269 (N_7269,N_4790,N_4494);
or U7270 (N_7270,N_5054,N_4432);
and U7271 (N_7271,N_4552,N_4358);
or U7272 (N_7272,N_4227,N_4433);
and U7273 (N_7273,N_5950,N_5956);
and U7274 (N_7274,N_5436,N_5271);
nor U7275 (N_7275,N_5878,N_4902);
nor U7276 (N_7276,N_5256,N_5802);
or U7277 (N_7277,N_5065,N_4783);
nor U7278 (N_7278,N_5534,N_5650);
or U7279 (N_7279,N_5003,N_4247);
and U7280 (N_7280,N_5023,N_4919);
or U7281 (N_7281,N_5265,N_4596);
and U7282 (N_7282,N_4369,N_5819);
or U7283 (N_7283,N_5757,N_5084);
or U7284 (N_7284,N_4144,N_4531);
nor U7285 (N_7285,N_4147,N_4451);
and U7286 (N_7286,N_5652,N_4048);
xor U7287 (N_7287,N_5518,N_4979);
xor U7288 (N_7288,N_5261,N_4410);
nor U7289 (N_7289,N_4862,N_5169);
and U7290 (N_7290,N_5417,N_4247);
xor U7291 (N_7291,N_4025,N_5526);
nand U7292 (N_7292,N_4449,N_5177);
or U7293 (N_7293,N_5935,N_5459);
xor U7294 (N_7294,N_4036,N_5432);
nor U7295 (N_7295,N_4582,N_4297);
nand U7296 (N_7296,N_4872,N_5188);
xor U7297 (N_7297,N_5281,N_5144);
xnor U7298 (N_7298,N_5904,N_4262);
or U7299 (N_7299,N_5063,N_4991);
or U7300 (N_7300,N_4623,N_5751);
xor U7301 (N_7301,N_4194,N_4270);
nand U7302 (N_7302,N_5242,N_5656);
xor U7303 (N_7303,N_5546,N_5691);
nor U7304 (N_7304,N_5627,N_5775);
xor U7305 (N_7305,N_4854,N_5257);
nor U7306 (N_7306,N_5558,N_4154);
xnor U7307 (N_7307,N_4973,N_5325);
nor U7308 (N_7308,N_5968,N_5451);
xnor U7309 (N_7309,N_4233,N_4991);
and U7310 (N_7310,N_4453,N_5250);
or U7311 (N_7311,N_4774,N_5201);
nor U7312 (N_7312,N_5312,N_4593);
nand U7313 (N_7313,N_5583,N_4005);
nand U7314 (N_7314,N_4006,N_5498);
or U7315 (N_7315,N_4715,N_5413);
xor U7316 (N_7316,N_5657,N_4776);
or U7317 (N_7317,N_4820,N_4348);
and U7318 (N_7318,N_4332,N_4607);
or U7319 (N_7319,N_5356,N_5449);
nor U7320 (N_7320,N_5743,N_4338);
nand U7321 (N_7321,N_4614,N_4062);
nand U7322 (N_7322,N_5029,N_4468);
nand U7323 (N_7323,N_5114,N_5896);
nor U7324 (N_7324,N_4309,N_5619);
and U7325 (N_7325,N_5240,N_5300);
and U7326 (N_7326,N_5781,N_4445);
xnor U7327 (N_7327,N_5870,N_4543);
nor U7328 (N_7328,N_4201,N_4680);
nor U7329 (N_7329,N_5915,N_5152);
xnor U7330 (N_7330,N_4961,N_4071);
and U7331 (N_7331,N_4145,N_5390);
or U7332 (N_7332,N_5930,N_4512);
or U7333 (N_7333,N_4218,N_5551);
xor U7334 (N_7334,N_4744,N_4500);
and U7335 (N_7335,N_4707,N_5424);
nor U7336 (N_7336,N_4259,N_5353);
or U7337 (N_7337,N_5199,N_4309);
nand U7338 (N_7338,N_5152,N_5144);
nor U7339 (N_7339,N_4224,N_4676);
nor U7340 (N_7340,N_4600,N_4816);
xor U7341 (N_7341,N_5940,N_4389);
nand U7342 (N_7342,N_5837,N_4262);
nand U7343 (N_7343,N_4051,N_5911);
or U7344 (N_7344,N_4850,N_5304);
xnor U7345 (N_7345,N_5629,N_5897);
nand U7346 (N_7346,N_4674,N_5696);
and U7347 (N_7347,N_5891,N_5155);
or U7348 (N_7348,N_5102,N_5617);
xnor U7349 (N_7349,N_4065,N_4024);
or U7350 (N_7350,N_4195,N_5866);
nand U7351 (N_7351,N_5477,N_4275);
or U7352 (N_7352,N_4685,N_5970);
or U7353 (N_7353,N_5854,N_5766);
or U7354 (N_7354,N_5564,N_5370);
and U7355 (N_7355,N_5747,N_4638);
nor U7356 (N_7356,N_5657,N_5963);
xnor U7357 (N_7357,N_5122,N_5134);
nand U7358 (N_7358,N_4571,N_5272);
nor U7359 (N_7359,N_5220,N_4572);
nand U7360 (N_7360,N_5589,N_4825);
nand U7361 (N_7361,N_4975,N_5352);
xnor U7362 (N_7362,N_4062,N_4377);
and U7363 (N_7363,N_5540,N_5818);
nor U7364 (N_7364,N_4131,N_4698);
or U7365 (N_7365,N_5980,N_5489);
nand U7366 (N_7366,N_4167,N_5429);
and U7367 (N_7367,N_4694,N_4323);
nand U7368 (N_7368,N_4473,N_5238);
and U7369 (N_7369,N_4649,N_5556);
nor U7370 (N_7370,N_5166,N_4914);
xnor U7371 (N_7371,N_5760,N_4442);
nor U7372 (N_7372,N_4713,N_4638);
xnor U7373 (N_7373,N_5541,N_5164);
nor U7374 (N_7374,N_5829,N_5954);
nand U7375 (N_7375,N_5752,N_4134);
xnor U7376 (N_7376,N_4929,N_5674);
nor U7377 (N_7377,N_5969,N_5753);
or U7378 (N_7378,N_4420,N_5092);
and U7379 (N_7379,N_4326,N_5320);
and U7380 (N_7380,N_4476,N_4400);
nor U7381 (N_7381,N_4672,N_5999);
nand U7382 (N_7382,N_5026,N_5414);
nor U7383 (N_7383,N_5060,N_4693);
xnor U7384 (N_7384,N_5054,N_5765);
nor U7385 (N_7385,N_4341,N_5347);
or U7386 (N_7386,N_5923,N_5598);
nand U7387 (N_7387,N_4660,N_4304);
nor U7388 (N_7388,N_4061,N_4608);
or U7389 (N_7389,N_5001,N_4357);
nand U7390 (N_7390,N_4428,N_4876);
nor U7391 (N_7391,N_4640,N_4819);
xnor U7392 (N_7392,N_5057,N_5512);
nor U7393 (N_7393,N_4228,N_5385);
and U7394 (N_7394,N_5557,N_4943);
nor U7395 (N_7395,N_4927,N_4131);
or U7396 (N_7396,N_4608,N_5051);
nor U7397 (N_7397,N_5619,N_4187);
and U7398 (N_7398,N_5472,N_4831);
and U7399 (N_7399,N_5237,N_5061);
xnor U7400 (N_7400,N_4292,N_5129);
nor U7401 (N_7401,N_5499,N_4137);
xnor U7402 (N_7402,N_4336,N_5123);
and U7403 (N_7403,N_5032,N_4632);
and U7404 (N_7404,N_4852,N_5543);
nand U7405 (N_7405,N_4140,N_4812);
xnor U7406 (N_7406,N_4770,N_4915);
xor U7407 (N_7407,N_5932,N_5533);
nor U7408 (N_7408,N_4378,N_5497);
and U7409 (N_7409,N_5302,N_5637);
nor U7410 (N_7410,N_5839,N_5203);
or U7411 (N_7411,N_4640,N_4509);
nor U7412 (N_7412,N_4068,N_5178);
xnor U7413 (N_7413,N_4907,N_5558);
xnor U7414 (N_7414,N_4312,N_5641);
or U7415 (N_7415,N_4143,N_4705);
nand U7416 (N_7416,N_5532,N_4961);
nor U7417 (N_7417,N_4757,N_4958);
xnor U7418 (N_7418,N_5440,N_4170);
nor U7419 (N_7419,N_4261,N_4678);
nand U7420 (N_7420,N_4665,N_4007);
and U7421 (N_7421,N_4848,N_5991);
nor U7422 (N_7422,N_5813,N_5458);
or U7423 (N_7423,N_4111,N_4422);
and U7424 (N_7424,N_5119,N_4285);
xnor U7425 (N_7425,N_4054,N_5066);
nand U7426 (N_7426,N_5393,N_4167);
nand U7427 (N_7427,N_5219,N_4550);
nand U7428 (N_7428,N_5828,N_4215);
or U7429 (N_7429,N_5920,N_5333);
or U7430 (N_7430,N_4053,N_5155);
or U7431 (N_7431,N_4625,N_4784);
nor U7432 (N_7432,N_5615,N_5704);
or U7433 (N_7433,N_5841,N_4453);
nand U7434 (N_7434,N_5654,N_5479);
nor U7435 (N_7435,N_4018,N_4302);
nand U7436 (N_7436,N_4671,N_4055);
nor U7437 (N_7437,N_4306,N_5610);
nand U7438 (N_7438,N_4496,N_4592);
and U7439 (N_7439,N_4574,N_5220);
nor U7440 (N_7440,N_4155,N_5999);
or U7441 (N_7441,N_4927,N_4536);
and U7442 (N_7442,N_4877,N_5278);
or U7443 (N_7443,N_5707,N_4048);
nand U7444 (N_7444,N_4636,N_4590);
and U7445 (N_7445,N_5556,N_5314);
or U7446 (N_7446,N_4937,N_4344);
xor U7447 (N_7447,N_4159,N_4292);
or U7448 (N_7448,N_5842,N_4002);
and U7449 (N_7449,N_4676,N_5986);
or U7450 (N_7450,N_5464,N_4957);
nor U7451 (N_7451,N_4882,N_5924);
nand U7452 (N_7452,N_4410,N_4400);
xnor U7453 (N_7453,N_4840,N_5522);
nand U7454 (N_7454,N_5230,N_5518);
or U7455 (N_7455,N_4970,N_5229);
or U7456 (N_7456,N_4913,N_4943);
nand U7457 (N_7457,N_4572,N_4676);
or U7458 (N_7458,N_5681,N_4555);
nor U7459 (N_7459,N_5630,N_5364);
nor U7460 (N_7460,N_4757,N_4858);
and U7461 (N_7461,N_4732,N_5440);
or U7462 (N_7462,N_5226,N_4863);
or U7463 (N_7463,N_4397,N_5918);
nand U7464 (N_7464,N_5386,N_5465);
and U7465 (N_7465,N_5056,N_4326);
nand U7466 (N_7466,N_4474,N_5221);
nor U7467 (N_7467,N_4368,N_4619);
and U7468 (N_7468,N_5019,N_5183);
and U7469 (N_7469,N_5307,N_5576);
nand U7470 (N_7470,N_5151,N_4753);
xnor U7471 (N_7471,N_4674,N_4678);
nor U7472 (N_7472,N_4908,N_5165);
xor U7473 (N_7473,N_4703,N_5129);
xor U7474 (N_7474,N_5237,N_4739);
nand U7475 (N_7475,N_5412,N_4856);
nor U7476 (N_7476,N_4131,N_4472);
and U7477 (N_7477,N_5420,N_5903);
and U7478 (N_7478,N_4573,N_5677);
xor U7479 (N_7479,N_5978,N_5274);
nor U7480 (N_7480,N_5983,N_5676);
nand U7481 (N_7481,N_4531,N_4281);
nand U7482 (N_7482,N_5434,N_5964);
nor U7483 (N_7483,N_5160,N_5144);
nand U7484 (N_7484,N_4696,N_4895);
nor U7485 (N_7485,N_4474,N_5056);
nand U7486 (N_7486,N_5200,N_5039);
and U7487 (N_7487,N_4010,N_5513);
nor U7488 (N_7488,N_4526,N_5009);
xor U7489 (N_7489,N_5886,N_4819);
nand U7490 (N_7490,N_5830,N_4252);
and U7491 (N_7491,N_5292,N_4412);
nor U7492 (N_7492,N_5113,N_4043);
or U7493 (N_7493,N_4392,N_5151);
nor U7494 (N_7494,N_4313,N_4728);
or U7495 (N_7495,N_4879,N_4578);
xnor U7496 (N_7496,N_4347,N_4112);
nor U7497 (N_7497,N_5383,N_5732);
xnor U7498 (N_7498,N_4668,N_5416);
nor U7499 (N_7499,N_5117,N_4527);
or U7500 (N_7500,N_5303,N_5635);
nand U7501 (N_7501,N_5534,N_5230);
nor U7502 (N_7502,N_5990,N_5953);
nor U7503 (N_7503,N_4894,N_5090);
nand U7504 (N_7504,N_5004,N_4556);
xnor U7505 (N_7505,N_5502,N_4244);
nand U7506 (N_7506,N_4276,N_4173);
nor U7507 (N_7507,N_4210,N_4734);
nor U7508 (N_7508,N_4936,N_5130);
nor U7509 (N_7509,N_4099,N_4806);
and U7510 (N_7510,N_5117,N_5728);
nand U7511 (N_7511,N_5181,N_5509);
xor U7512 (N_7512,N_5322,N_5822);
and U7513 (N_7513,N_4299,N_5885);
xor U7514 (N_7514,N_4984,N_4048);
and U7515 (N_7515,N_5073,N_4311);
nor U7516 (N_7516,N_5405,N_5493);
nor U7517 (N_7517,N_4938,N_4074);
and U7518 (N_7518,N_5363,N_4913);
nand U7519 (N_7519,N_5300,N_5734);
and U7520 (N_7520,N_4001,N_5726);
nor U7521 (N_7521,N_4060,N_5595);
and U7522 (N_7522,N_5433,N_4377);
xnor U7523 (N_7523,N_5677,N_5617);
nand U7524 (N_7524,N_4631,N_4655);
nor U7525 (N_7525,N_5070,N_4658);
nand U7526 (N_7526,N_4354,N_4390);
xor U7527 (N_7527,N_4637,N_5471);
nor U7528 (N_7528,N_5207,N_4306);
nand U7529 (N_7529,N_4665,N_4447);
or U7530 (N_7530,N_4560,N_5688);
xnor U7531 (N_7531,N_5898,N_5270);
xnor U7532 (N_7532,N_5843,N_5143);
and U7533 (N_7533,N_4001,N_5198);
nor U7534 (N_7534,N_4025,N_5841);
or U7535 (N_7535,N_5804,N_4326);
nor U7536 (N_7536,N_5068,N_5181);
and U7537 (N_7537,N_4174,N_4510);
nand U7538 (N_7538,N_5864,N_4565);
nor U7539 (N_7539,N_5447,N_4584);
or U7540 (N_7540,N_5467,N_5403);
nand U7541 (N_7541,N_5327,N_5814);
nand U7542 (N_7542,N_5732,N_4519);
and U7543 (N_7543,N_5707,N_4229);
nor U7544 (N_7544,N_4652,N_5336);
or U7545 (N_7545,N_5621,N_4157);
nor U7546 (N_7546,N_4024,N_4697);
or U7547 (N_7547,N_4296,N_4422);
nor U7548 (N_7548,N_4488,N_4583);
and U7549 (N_7549,N_5898,N_4508);
or U7550 (N_7550,N_4514,N_5389);
or U7551 (N_7551,N_5656,N_4440);
and U7552 (N_7552,N_4227,N_5141);
and U7553 (N_7553,N_4642,N_5305);
or U7554 (N_7554,N_5521,N_4169);
or U7555 (N_7555,N_4744,N_4170);
or U7556 (N_7556,N_5783,N_4154);
nand U7557 (N_7557,N_4672,N_4400);
xor U7558 (N_7558,N_5548,N_4280);
and U7559 (N_7559,N_5290,N_5072);
or U7560 (N_7560,N_4141,N_5654);
and U7561 (N_7561,N_4285,N_5637);
or U7562 (N_7562,N_5894,N_4943);
and U7563 (N_7563,N_4440,N_5430);
and U7564 (N_7564,N_5308,N_5749);
nor U7565 (N_7565,N_4723,N_5205);
nand U7566 (N_7566,N_4292,N_4109);
or U7567 (N_7567,N_5362,N_5444);
xor U7568 (N_7568,N_5552,N_5860);
nor U7569 (N_7569,N_5362,N_5870);
nand U7570 (N_7570,N_4326,N_5315);
nor U7571 (N_7571,N_5069,N_5571);
and U7572 (N_7572,N_5039,N_4545);
xnor U7573 (N_7573,N_4086,N_4622);
nor U7574 (N_7574,N_5659,N_4600);
nor U7575 (N_7575,N_4123,N_4049);
or U7576 (N_7576,N_5622,N_4041);
nor U7577 (N_7577,N_4160,N_5951);
xnor U7578 (N_7578,N_5569,N_5841);
xor U7579 (N_7579,N_4218,N_4942);
nand U7580 (N_7580,N_4960,N_4097);
nor U7581 (N_7581,N_4340,N_5783);
nor U7582 (N_7582,N_4493,N_4934);
xnor U7583 (N_7583,N_5632,N_5755);
and U7584 (N_7584,N_5267,N_4978);
nand U7585 (N_7585,N_4522,N_5321);
and U7586 (N_7586,N_4079,N_4264);
nand U7587 (N_7587,N_5361,N_5953);
nor U7588 (N_7588,N_4938,N_4706);
nand U7589 (N_7589,N_5472,N_4920);
nor U7590 (N_7590,N_4865,N_4617);
nand U7591 (N_7591,N_4207,N_4672);
and U7592 (N_7592,N_4995,N_4566);
nand U7593 (N_7593,N_4105,N_5627);
nand U7594 (N_7594,N_5481,N_4820);
nor U7595 (N_7595,N_4185,N_4538);
nand U7596 (N_7596,N_5981,N_5619);
nor U7597 (N_7597,N_5264,N_5494);
nand U7598 (N_7598,N_4101,N_4587);
nand U7599 (N_7599,N_4348,N_5082);
nand U7600 (N_7600,N_5675,N_4512);
nand U7601 (N_7601,N_5138,N_5552);
nor U7602 (N_7602,N_5386,N_5999);
or U7603 (N_7603,N_4428,N_4316);
and U7604 (N_7604,N_4151,N_5003);
nor U7605 (N_7605,N_4656,N_5837);
nor U7606 (N_7606,N_4716,N_4615);
nand U7607 (N_7607,N_5880,N_4279);
nor U7608 (N_7608,N_5059,N_5946);
nand U7609 (N_7609,N_4056,N_4834);
or U7610 (N_7610,N_4756,N_4236);
nand U7611 (N_7611,N_5182,N_4031);
or U7612 (N_7612,N_4349,N_4616);
xnor U7613 (N_7613,N_4379,N_5081);
and U7614 (N_7614,N_4447,N_5365);
nor U7615 (N_7615,N_4295,N_5760);
or U7616 (N_7616,N_5224,N_5278);
nor U7617 (N_7617,N_5368,N_5766);
nand U7618 (N_7618,N_4973,N_5667);
nand U7619 (N_7619,N_4548,N_5168);
or U7620 (N_7620,N_5160,N_5653);
nor U7621 (N_7621,N_5200,N_5536);
xor U7622 (N_7622,N_4701,N_4345);
nand U7623 (N_7623,N_5653,N_5665);
nor U7624 (N_7624,N_4238,N_5273);
nor U7625 (N_7625,N_4916,N_5200);
nor U7626 (N_7626,N_5751,N_4959);
xor U7627 (N_7627,N_4541,N_4893);
nand U7628 (N_7628,N_5755,N_4518);
xnor U7629 (N_7629,N_4469,N_5334);
nor U7630 (N_7630,N_4414,N_4656);
and U7631 (N_7631,N_4025,N_4729);
and U7632 (N_7632,N_5119,N_5219);
and U7633 (N_7633,N_5421,N_5007);
or U7634 (N_7634,N_5029,N_5328);
and U7635 (N_7635,N_4275,N_4510);
nand U7636 (N_7636,N_4624,N_5942);
or U7637 (N_7637,N_4670,N_5918);
or U7638 (N_7638,N_4405,N_4451);
and U7639 (N_7639,N_4303,N_5890);
nand U7640 (N_7640,N_5885,N_5125);
nor U7641 (N_7641,N_5797,N_4002);
nand U7642 (N_7642,N_5020,N_4435);
or U7643 (N_7643,N_5176,N_5535);
nor U7644 (N_7644,N_5430,N_4736);
and U7645 (N_7645,N_4720,N_5572);
or U7646 (N_7646,N_4732,N_5593);
nand U7647 (N_7647,N_4634,N_5889);
nor U7648 (N_7648,N_4477,N_5368);
nand U7649 (N_7649,N_5604,N_4265);
xnor U7650 (N_7650,N_5432,N_5883);
nand U7651 (N_7651,N_5630,N_4464);
and U7652 (N_7652,N_4316,N_5755);
and U7653 (N_7653,N_4706,N_5514);
nand U7654 (N_7654,N_4420,N_5892);
xor U7655 (N_7655,N_5622,N_4979);
nand U7656 (N_7656,N_4224,N_4732);
xnor U7657 (N_7657,N_4172,N_5279);
nor U7658 (N_7658,N_5704,N_5805);
or U7659 (N_7659,N_5836,N_4625);
and U7660 (N_7660,N_5153,N_5793);
and U7661 (N_7661,N_4758,N_4970);
nor U7662 (N_7662,N_5736,N_5701);
and U7663 (N_7663,N_4481,N_5604);
nor U7664 (N_7664,N_5131,N_5156);
nor U7665 (N_7665,N_5209,N_4446);
xnor U7666 (N_7666,N_5098,N_4053);
nor U7667 (N_7667,N_5262,N_5592);
nand U7668 (N_7668,N_4151,N_4782);
and U7669 (N_7669,N_4720,N_4668);
nor U7670 (N_7670,N_5546,N_5969);
xor U7671 (N_7671,N_4012,N_4996);
nand U7672 (N_7672,N_5156,N_4892);
nor U7673 (N_7673,N_5415,N_5344);
xor U7674 (N_7674,N_5252,N_4431);
and U7675 (N_7675,N_4825,N_5684);
and U7676 (N_7676,N_4526,N_5264);
nand U7677 (N_7677,N_4859,N_4151);
xnor U7678 (N_7678,N_5500,N_4638);
and U7679 (N_7679,N_4591,N_4809);
nand U7680 (N_7680,N_5492,N_4095);
nor U7681 (N_7681,N_4255,N_4095);
nand U7682 (N_7682,N_4792,N_4833);
xor U7683 (N_7683,N_5161,N_5366);
and U7684 (N_7684,N_5930,N_4231);
xor U7685 (N_7685,N_4779,N_5106);
or U7686 (N_7686,N_5423,N_4092);
xnor U7687 (N_7687,N_5424,N_5716);
and U7688 (N_7688,N_5269,N_4436);
nand U7689 (N_7689,N_5341,N_4941);
nor U7690 (N_7690,N_5241,N_4285);
or U7691 (N_7691,N_4736,N_5961);
nand U7692 (N_7692,N_5004,N_5873);
or U7693 (N_7693,N_4251,N_5767);
or U7694 (N_7694,N_5231,N_5196);
nor U7695 (N_7695,N_4302,N_4800);
nor U7696 (N_7696,N_5311,N_4175);
and U7697 (N_7697,N_4032,N_5445);
xnor U7698 (N_7698,N_4529,N_4284);
xnor U7699 (N_7699,N_4704,N_5479);
and U7700 (N_7700,N_5305,N_5116);
or U7701 (N_7701,N_5461,N_5452);
and U7702 (N_7702,N_4596,N_5951);
nand U7703 (N_7703,N_5263,N_4909);
nor U7704 (N_7704,N_5922,N_4963);
and U7705 (N_7705,N_4190,N_4649);
nor U7706 (N_7706,N_4720,N_4900);
and U7707 (N_7707,N_5656,N_5016);
and U7708 (N_7708,N_4347,N_5577);
or U7709 (N_7709,N_4778,N_4515);
nor U7710 (N_7710,N_4807,N_5448);
xnor U7711 (N_7711,N_5151,N_5216);
and U7712 (N_7712,N_4779,N_4463);
nand U7713 (N_7713,N_4840,N_4618);
xor U7714 (N_7714,N_5245,N_5279);
or U7715 (N_7715,N_5262,N_5572);
and U7716 (N_7716,N_5992,N_4036);
nor U7717 (N_7717,N_4413,N_5790);
and U7718 (N_7718,N_4877,N_4038);
or U7719 (N_7719,N_5601,N_5743);
and U7720 (N_7720,N_4961,N_5072);
and U7721 (N_7721,N_4002,N_5317);
nand U7722 (N_7722,N_5842,N_5793);
nand U7723 (N_7723,N_4816,N_4979);
xor U7724 (N_7724,N_4743,N_4527);
nand U7725 (N_7725,N_5613,N_5709);
and U7726 (N_7726,N_4198,N_4450);
nand U7727 (N_7727,N_5009,N_5739);
nor U7728 (N_7728,N_4533,N_4792);
nor U7729 (N_7729,N_5350,N_4073);
xor U7730 (N_7730,N_5239,N_4719);
xor U7731 (N_7731,N_5034,N_5206);
xnor U7732 (N_7732,N_5107,N_4904);
nor U7733 (N_7733,N_4290,N_4166);
nand U7734 (N_7734,N_4343,N_5464);
and U7735 (N_7735,N_5006,N_5612);
and U7736 (N_7736,N_4311,N_5463);
and U7737 (N_7737,N_5620,N_5286);
or U7738 (N_7738,N_4987,N_5552);
nor U7739 (N_7739,N_4585,N_4676);
xnor U7740 (N_7740,N_5794,N_4843);
nor U7741 (N_7741,N_5780,N_4167);
nand U7742 (N_7742,N_4760,N_4328);
nor U7743 (N_7743,N_5361,N_4806);
nor U7744 (N_7744,N_4286,N_4168);
nor U7745 (N_7745,N_5298,N_4152);
and U7746 (N_7746,N_4981,N_5179);
xor U7747 (N_7747,N_4910,N_5040);
xnor U7748 (N_7748,N_5509,N_4532);
nor U7749 (N_7749,N_4024,N_4672);
or U7750 (N_7750,N_4635,N_4045);
and U7751 (N_7751,N_4549,N_5058);
xor U7752 (N_7752,N_5574,N_5383);
nor U7753 (N_7753,N_5330,N_4173);
nand U7754 (N_7754,N_4475,N_4874);
and U7755 (N_7755,N_4856,N_5728);
xor U7756 (N_7756,N_5612,N_4897);
nand U7757 (N_7757,N_5801,N_5239);
and U7758 (N_7758,N_5429,N_5393);
xor U7759 (N_7759,N_4620,N_5659);
or U7760 (N_7760,N_5037,N_4775);
nor U7761 (N_7761,N_5065,N_5786);
xnor U7762 (N_7762,N_4933,N_5716);
xnor U7763 (N_7763,N_5307,N_5066);
and U7764 (N_7764,N_4573,N_4668);
and U7765 (N_7765,N_5724,N_4806);
nand U7766 (N_7766,N_4298,N_4638);
xnor U7767 (N_7767,N_5162,N_5663);
or U7768 (N_7768,N_4317,N_5061);
xnor U7769 (N_7769,N_4594,N_5612);
nor U7770 (N_7770,N_4806,N_5205);
nor U7771 (N_7771,N_4030,N_5628);
or U7772 (N_7772,N_4613,N_4018);
xnor U7773 (N_7773,N_5541,N_4546);
and U7774 (N_7774,N_4434,N_4910);
and U7775 (N_7775,N_5021,N_5742);
xnor U7776 (N_7776,N_4547,N_4823);
nand U7777 (N_7777,N_5760,N_4315);
or U7778 (N_7778,N_5399,N_5340);
xnor U7779 (N_7779,N_5681,N_5513);
xnor U7780 (N_7780,N_5622,N_4423);
nor U7781 (N_7781,N_4539,N_5159);
nand U7782 (N_7782,N_4122,N_4580);
and U7783 (N_7783,N_5633,N_5093);
xor U7784 (N_7784,N_5170,N_5106);
nor U7785 (N_7785,N_5795,N_4264);
xor U7786 (N_7786,N_5423,N_4705);
xor U7787 (N_7787,N_5883,N_4035);
xor U7788 (N_7788,N_5584,N_4976);
and U7789 (N_7789,N_4931,N_5028);
or U7790 (N_7790,N_5969,N_5831);
nand U7791 (N_7791,N_4902,N_5555);
xnor U7792 (N_7792,N_4912,N_5581);
xnor U7793 (N_7793,N_5926,N_5500);
nand U7794 (N_7794,N_4971,N_4553);
xor U7795 (N_7795,N_4732,N_4346);
xor U7796 (N_7796,N_4593,N_4679);
nand U7797 (N_7797,N_4242,N_4735);
nor U7798 (N_7798,N_4102,N_5246);
or U7799 (N_7799,N_5861,N_5697);
xnor U7800 (N_7800,N_5416,N_5920);
nor U7801 (N_7801,N_5806,N_5425);
nand U7802 (N_7802,N_4931,N_5176);
nand U7803 (N_7803,N_4948,N_5409);
xor U7804 (N_7804,N_5670,N_5800);
and U7805 (N_7805,N_5427,N_5714);
and U7806 (N_7806,N_4314,N_4851);
and U7807 (N_7807,N_4139,N_4881);
nor U7808 (N_7808,N_4345,N_5944);
nor U7809 (N_7809,N_5477,N_5087);
or U7810 (N_7810,N_4031,N_5563);
xor U7811 (N_7811,N_4222,N_4554);
or U7812 (N_7812,N_5272,N_4256);
nor U7813 (N_7813,N_4459,N_4023);
or U7814 (N_7814,N_4857,N_5695);
and U7815 (N_7815,N_4018,N_5566);
xnor U7816 (N_7816,N_4978,N_5731);
nand U7817 (N_7817,N_4998,N_4488);
nor U7818 (N_7818,N_5363,N_4497);
and U7819 (N_7819,N_5105,N_5341);
nor U7820 (N_7820,N_4302,N_5240);
or U7821 (N_7821,N_4411,N_4667);
nand U7822 (N_7822,N_4130,N_5024);
or U7823 (N_7823,N_5862,N_4664);
and U7824 (N_7824,N_4030,N_5480);
and U7825 (N_7825,N_4639,N_4085);
nor U7826 (N_7826,N_4270,N_4960);
or U7827 (N_7827,N_4214,N_4029);
nand U7828 (N_7828,N_5691,N_4384);
nor U7829 (N_7829,N_4867,N_4802);
or U7830 (N_7830,N_5641,N_4413);
xnor U7831 (N_7831,N_5628,N_5637);
and U7832 (N_7832,N_5226,N_5502);
or U7833 (N_7833,N_5208,N_4554);
nand U7834 (N_7834,N_5451,N_5824);
nor U7835 (N_7835,N_4771,N_4266);
nor U7836 (N_7836,N_5680,N_5395);
xor U7837 (N_7837,N_5018,N_4579);
nor U7838 (N_7838,N_4541,N_4086);
xnor U7839 (N_7839,N_4397,N_5920);
and U7840 (N_7840,N_5452,N_4504);
nor U7841 (N_7841,N_5660,N_4837);
nand U7842 (N_7842,N_5967,N_5750);
or U7843 (N_7843,N_4881,N_5633);
xor U7844 (N_7844,N_5564,N_4198);
nor U7845 (N_7845,N_5440,N_4213);
nor U7846 (N_7846,N_5178,N_5089);
and U7847 (N_7847,N_5231,N_4754);
nor U7848 (N_7848,N_4886,N_5138);
xor U7849 (N_7849,N_4164,N_5005);
and U7850 (N_7850,N_4403,N_5491);
or U7851 (N_7851,N_4782,N_4585);
and U7852 (N_7852,N_4960,N_5166);
nor U7853 (N_7853,N_4615,N_5261);
xor U7854 (N_7854,N_5535,N_4439);
or U7855 (N_7855,N_4529,N_4918);
nand U7856 (N_7856,N_4441,N_4682);
nor U7857 (N_7857,N_4957,N_5829);
nand U7858 (N_7858,N_5537,N_4905);
and U7859 (N_7859,N_5216,N_5780);
and U7860 (N_7860,N_4503,N_4311);
nor U7861 (N_7861,N_4503,N_5782);
xor U7862 (N_7862,N_5361,N_4789);
and U7863 (N_7863,N_4083,N_4366);
nor U7864 (N_7864,N_5475,N_4202);
nor U7865 (N_7865,N_5314,N_4806);
nor U7866 (N_7866,N_4919,N_4659);
xor U7867 (N_7867,N_5939,N_4416);
or U7868 (N_7868,N_5511,N_4219);
and U7869 (N_7869,N_4460,N_5379);
nand U7870 (N_7870,N_4383,N_4690);
nand U7871 (N_7871,N_5922,N_5361);
or U7872 (N_7872,N_4860,N_4282);
nand U7873 (N_7873,N_4008,N_4804);
nor U7874 (N_7874,N_5307,N_5040);
nor U7875 (N_7875,N_5430,N_5182);
and U7876 (N_7876,N_4562,N_4041);
nor U7877 (N_7877,N_4403,N_5364);
and U7878 (N_7878,N_4445,N_4996);
nand U7879 (N_7879,N_5238,N_5232);
nand U7880 (N_7880,N_4836,N_4950);
and U7881 (N_7881,N_4654,N_4577);
or U7882 (N_7882,N_5200,N_5045);
nand U7883 (N_7883,N_5855,N_5219);
nor U7884 (N_7884,N_4309,N_5241);
or U7885 (N_7885,N_4375,N_5914);
or U7886 (N_7886,N_5693,N_4788);
and U7887 (N_7887,N_4798,N_4230);
xnor U7888 (N_7888,N_5928,N_4569);
xnor U7889 (N_7889,N_4968,N_5237);
and U7890 (N_7890,N_5631,N_4103);
xor U7891 (N_7891,N_5087,N_5119);
or U7892 (N_7892,N_5078,N_5766);
nand U7893 (N_7893,N_4007,N_5419);
or U7894 (N_7894,N_4078,N_4150);
or U7895 (N_7895,N_4112,N_4095);
nor U7896 (N_7896,N_5894,N_4570);
nor U7897 (N_7897,N_4036,N_5572);
and U7898 (N_7898,N_5540,N_5544);
nor U7899 (N_7899,N_4776,N_4819);
nor U7900 (N_7900,N_5209,N_5531);
or U7901 (N_7901,N_5968,N_5035);
nand U7902 (N_7902,N_5002,N_4254);
nand U7903 (N_7903,N_5637,N_4820);
nand U7904 (N_7904,N_4222,N_5261);
nor U7905 (N_7905,N_5901,N_4985);
nor U7906 (N_7906,N_4356,N_5820);
nor U7907 (N_7907,N_5715,N_4526);
nand U7908 (N_7908,N_5735,N_4525);
nor U7909 (N_7909,N_5896,N_5096);
nand U7910 (N_7910,N_4836,N_4368);
and U7911 (N_7911,N_5579,N_5886);
xnor U7912 (N_7912,N_4268,N_4512);
xnor U7913 (N_7913,N_5993,N_5849);
or U7914 (N_7914,N_4153,N_4468);
and U7915 (N_7915,N_4175,N_5116);
nand U7916 (N_7916,N_4617,N_4201);
nor U7917 (N_7917,N_4522,N_4200);
nor U7918 (N_7918,N_4133,N_4437);
or U7919 (N_7919,N_4287,N_4586);
nand U7920 (N_7920,N_4387,N_5515);
xor U7921 (N_7921,N_4879,N_4553);
and U7922 (N_7922,N_5237,N_4524);
or U7923 (N_7923,N_5425,N_5327);
or U7924 (N_7924,N_5300,N_4191);
and U7925 (N_7925,N_5208,N_5727);
or U7926 (N_7926,N_5855,N_4120);
nor U7927 (N_7927,N_5133,N_5991);
and U7928 (N_7928,N_5839,N_5662);
and U7929 (N_7929,N_5029,N_4978);
nor U7930 (N_7930,N_5430,N_4902);
xnor U7931 (N_7931,N_5728,N_5077);
nor U7932 (N_7932,N_5272,N_5406);
and U7933 (N_7933,N_5677,N_5743);
nand U7934 (N_7934,N_4122,N_4161);
and U7935 (N_7935,N_5634,N_4664);
nand U7936 (N_7936,N_4818,N_4144);
xor U7937 (N_7937,N_4431,N_4911);
nor U7938 (N_7938,N_4965,N_5261);
nand U7939 (N_7939,N_4519,N_4384);
and U7940 (N_7940,N_4703,N_5058);
nand U7941 (N_7941,N_4835,N_4893);
xnor U7942 (N_7942,N_5355,N_4299);
nor U7943 (N_7943,N_4972,N_5843);
and U7944 (N_7944,N_5300,N_5397);
xnor U7945 (N_7945,N_5503,N_5732);
or U7946 (N_7946,N_5413,N_4823);
or U7947 (N_7947,N_5274,N_5613);
and U7948 (N_7948,N_5657,N_5545);
nand U7949 (N_7949,N_5574,N_4099);
nor U7950 (N_7950,N_5119,N_4045);
nor U7951 (N_7951,N_4957,N_5573);
nand U7952 (N_7952,N_5610,N_4262);
nor U7953 (N_7953,N_4576,N_5745);
nand U7954 (N_7954,N_4697,N_4838);
xor U7955 (N_7955,N_4097,N_4493);
xnor U7956 (N_7956,N_4974,N_4785);
nor U7957 (N_7957,N_4752,N_5230);
or U7958 (N_7958,N_4903,N_4038);
and U7959 (N_7959,N_4880,N_4548);
and U7960 (N_7960,N_5537,N_4255);
xor U7961 (N_7961,N_4317,N_5195);
nor U7962 (N_7962,N_5577,N_5151);
xnor U7963 (N_7963,N_5655,N_4889);
or U7964 (N_7964,N_4288,N_4154);
xnor U7965 (N_7965,N_4833,N_4483);
xor U7966 (N_7966,N_4239,N_4824);
xnor U7967 (N_7967,N_5653,N_4427);
or U7968 (N_7968,N_4270,N_5180);
or U7969 (N_7969,N_4709,N_5986);
and U7970 (N_7970,N_5537,N_4664);
xor U7971 (N_7971,N_5778,N_5837);
and U7972 (N_7972,N_5309,N_5668);
and U7973 (N_7973,N_5170,N_5185);
and U7974 (N_7974,N_4063,N_4706);
xor U7975 (N_7975,N_4073,N_5484);
nand U7976 (N_7976,N_4460,N_4542);
xor U7977 (N_7977,N_5601,N_4759);
and U7978 (N_7978,N_5710,N_5520);
or U7979 (N_7979,N_4464,N_5104);
xnor U7980 (N_7980,N_4862,N_5227);
nand U7981 (N_7981,N_4000,N_5748);
nand U7982 (N_7982,N_4362,N_4011);
xor U7983 (N_7983,N_4015,N_4129);
and U7984 (N_7984,N_4369,N_5888);
nand U7985 (N_7985,N_5344,N_4919);
or U7986 (N_7986,N_5184,N_5793);
nand U7987 (N_7987,N_5844,N_4644);
xnor U7988 (N_7988,N_4796,N_4465);
xor U7989 (N_7989,N_4635,N_4055);
nand U7990 (N_7990,N_5262,N_5879);
xor U7991 (N_7991,N_4812,N_4267);
xnor U7992 (N_7992,N_5530,N_4794);
xnor U7993 (N_7993,N_5139,N_4049);
nand U7994 (N_7994,N_5178,N_4066);
nor U7995 (N_7995,N_5155,N_4023);
xnor U7996 (N_7996,N_5912,N_5518);
xnor U7997 (N_7997,N_4510,N_4836);
nand U7998 (N_7998,N_4527,N_5411);
and U7999 (N_7999,N_5330,N_4274);
xor U8000 (N_8000,N_7378,N_7765);
xnor U8001 (N_8001,N_6644,N_7586);
or U8002 (N_8002,N_6845,N_6656);
nor U8003 (N_8003,N_6496,N_6968);
xnor U8004 (N_8004,N_7697,N_7166);
or U8005 (N_8005,N_6293,N_6985);
and U8006 (N_8006,N_6577,N_6659);
and U8007 (N_8007,N_6389,N_7076);
xnor U8008 (N_8008,N_7556,N_6828);
nand U8009 (N_8009,N_6226,N_6144);
or U8010 (N_8010,N_7183,N_6383);
nand U8011 (N_8011,N_7093,N_7473);
or U8012 (N_8012,N_7426,N_7600);
or U8013 (N_8013,N_6454,N_7597);
nand U8014 (N_8014,N_6660,N_6098);
nand U8015 (N_8015,N_7333,N_6569);
or U8016 (N_8016,N_6614,N_6765);
and U8017 (N_8017,N_6083,N_6865);
nor U8018 (N_8018,N_7495,N_7810);
nor U8019 (N_8019,N_6195,N_7956);
and U8020 (N_8020,N_6394,N_7288);
nor U8021 (N_8021,N_7014,N_6155);
nor U8022 (N_8022,N_6088,N_7063);
and U8023 (N_8023,N_6814,N_6740);
nor U8024 (N_8024,N_7943,N_6450);
nor U8025 (N_8025,N_6837,N_6709);
nand U8026 (N_8026,N_7270,N_6286);
nor U8027 (N_8027,N_6125,N_6752);
nor U8028 (N_8028,N_6579,N_7368);
and U8029 (N_8029,N_6060,N_7976);
nand U8030 (N_8030,N_7030,N_6846);
or U8031 (N_8031,N_7027,N_6217);
or U8032 (N_8032,N_7787,N_7138);
nor U8033 (N_8033,N_7879,N_6610);
or U8034 (N_8034,N_7646,N_7411);
or U8035 (N_8035,N_6482,N_6469);
nand U8036 (N_8036,N_6710,N_6984);
and U8037 (N_8037,N_6992,N_7724);
xnor U8038 (N_8038,N_7779,N_6794);
xor U8039 (N_8039,N_6576,N_7256);
xnor U8040 (N_8040,N_7221,N_6595);
and U8041 (N_8041,N_7583,N_7730);
and U8042 (N_8042,N_7712,N_6178);
nor U8043 (N_8043,N_7169,N_7066);
xor U8044 (N_8044,N_6434,N_6929);
xor U8045 (N_8045,N_6042,N_6866);
or U8046 (N_8046,N_6906,N_6091);
and U8047 (N_8047,N_6957,N_6547);
and U8048 (N_8048,N_6014,N_6243);
or U8049 (N_8049,N_6292,N_6111);
nand U8050 (N_8050,N_6067,N_7994);
nor U8051 (N_8051,N_6002,N_6522);
nor U8052 (N_8052,N_6463,N_7132);
or U8053 (N_8053,N_7992,N_7963);
xnor U8054 (N_8054,N_6649,N_7734);
nand U8055 (N_8055,N_6089,N_7342);
or U8056 (N_8056,N_6065,N_6702);
nand U8057 (N_8057,N_7369,N_7893);
nor U8058 (N_8058,N_6035,N_6953);
nor U8059 (N_8059,N_7627,N_6824);
and U8060 (N_8060,N_6330,N_6673);
and U8061 (N_8061,N_7782,N_7385);
or U8062 (N_8062,N_7991,N_7885);
or U8063 (N_8063,N_6544,N_6749);
nand U8064 (N_8064,N_6820,N_6112);
nor U8065 (N_8065,N_7259,N_7029);
xor U8066 (N_8066,N_7868,N_7798);
and U8067 (N_8067,N_6113,N_7609);
nand U8068 (N_8068,N_6848,N_6907);
and U8069 (N_8069,N_7479,N_6304);
xnor U8070 (N_8070,N_7317,N_6689);
and U8071 (N_8071,N_6215,N_6407);
nor U8072 (N_8072,N_6607,N_7691);
nor U8073 (N_8073,N_7575,N_7968);
xor U8074 (N_8074,N_7837,N_7630);
or U8075 (N_8075,N_6104,N_7995);
or U8076 (N_8076,N_6225,N_6591);
and U8077 (N_8077,N_7075,N_7817);
nor U8078 (N_8078,N_6315,N_7933);
nor U8079 (N_8079,N_7960,N_6952);
and U8080 (N_8080,N_7329,N_6753);
nor U8081 (N_8081,N_6885,N_6543);
and U8082 (N_8082,N_7710,N_6021);
nor U8083 (N_8083,N_6402,N_6258);
nor U8084 (N_8084,N_7663,N_6766);
nand U8085 (N_8085,N_6365,N_6223);
and U8086 (N_8086,N_7927,N_7682);
nor U8087 (N_8087,N_6371,N_6031);
nand U8088 (N_8088,N_7072,N_6274);
xnor U8089 (N_8089,N_7695,N_6367);
and U8090 (N_8090,N_7122,N_6821);
xnor U8091 (N_8091,N_7967,N_7334);
or U8092 (N_8092,N_7178,N_6829);
or U8093 (N_8093,N_6206,N_6108);
nor U8094 (N_8094,N_6197,N_6196);
and U8095 (N_8095,N_6880,N_7338);
or U8096 (N_8096,N_6151,N_7536);
xor U8097 (N_8097,N_7618,N_7962);
nor U8098 (N_8098,N_6140,N_6433);
and U8099 (N_8099,N_7105,N_7661);
nor U8100 (N_8100,N_7624,N_6387);
nor U8101 (N_8101,N_6411,N_7899);
or U8102 (N_8102,N_6686,N_7409);
xnor U8103 (N_8103,N_7892,N_7750);
or U8104 (N_8104,N_7263,N_6359);
nand U8105 (N_8105,N_6316,N_6982);
and U8106 (N_8106,N_7584,N_6988);
nor U8107 (N_8107,N_6935,N_6527);
and U8108 (N_8108,N_6375,N_6882);
or U8109 (N_8109,N_6976,N_7662);
xnor U8110 (N_8110,N_6210,N_7325);
and U8111 (N_8111,N_6449,N_7469);
and U8112 (N_8112,N_6627,N_7635);
or U8113 (N_8113,N_7234,N_6729);
and U8114 (N_8114,N_7891,N_6425);
nand U8115 (N_8115,N_7861,N_7977);
xnor U8116 (N_8116,N_6755,N_6194);
and U8117 (N_8117,N_6926,N_6071);
xnor U8118 (N_8118,N_7327,N_7870);
xnor U8119 (N_8119,N_6468,N_7195);
nor U8120 (N_8120,N_6064,N_6989);
nor U8121 (N_8121,N_6580,N_6983);
or U8122 (N_8122,N_6924,N_7971);
or U8123 (N_8123,N_6581,N_7621);
nand U8124 (N_8124,N_7500,N_7135);
and U8125 (N_8125,N_7362,N_7973);
and U8126 (N_8126,N_7110,N_6492);
nor U8127 (N_8127,N_7652,N_6305);
xor U8128 (N_8128,N_7504,N_6199);
or U8129 (N_8129,N_6693,N_6205);
and U8130 (N_8130,N_7328,N_6096);
and U8131 (N_8131,N_7518,N_7370);
and U8132 (N_8132,N_6027,N_7211);
xnor U8133 (N_8133,N_6115,N_6373);
nor U8134 (N_8134,N_7755,N_7843);
and U8135 (N_8135,N_7688,N_7533);
nor U8136 (N_8136,N_7241,N_6235);
nand U8137 (N_8137,N_6748,N_6903);
nand U8138 (N_8138,N_7477,N_7754);
xnor U8139 (N_8139,N_7738,N_7881);
nor U8140 (N_8140,N_7488,N_7939);
xnor U8141 (N_8141,N_6323,N_7796);
nand U8142 (N_8142,N_6704,N_7209);
xnor U8143 (N_8143,N_7161,N_7539);
or U8144 (N_8144,N_6545,N_6203);
xnor U8145 (N_8145,N_7783,N_6222);
xor U8146 (N_8146,N_6176,N_7000);
and U8147 (N_8147,N_7445,N_7350);
nor U8148 (N_8148,N_7985,N_7527);
nor U8149 (N_8149,N_6959,N_6084);
nand U8150 (N_8150,N_6028,N_7756);
or U8151 (N_8151,N_7714,N_6272);
nand U8152 (N_8152,N_7393,N_7483);
and U8153 (N_8153,N_7410,N_6921);
nand U8154 (N_8154,N_6675,N_7223);
nor U8155 (N_8155,N_7875,N_6987);
nor U8156 (N_8156,N_6583,N_6836);
or U8157 (N_8157,N_7711,N_7692);
nand U8158 (N_8158,N_6590,N_7282);
nor U8159 (N_8159,N_6619,N_7450);
xor U8160 (N_8160,N_6052,N_6440);
and U8161 (N_8161,N_6932,N_7098);
and U8162 (N_8162,N_7626,N_7744);
nand U8163 (N_8163,N_7677,N_6066);
nor U8164 (N_8164,N_6979,N_7103);
xnor U8165 (N_8165,N_6737,N_6174);
nor U8166 (N_8166,N_7847,N_7401);
and U8167 (N_8167,N_7202,N_7516);
nand U8168 (N_8168,N_7153,N_7954);
nand U8169 (N_8169,N_6382,N_6401);
nor U8170 (N_8170,N_6894,N_6445);
nor U8171 (N_8171,N_6722,N_7038);
and U8172 (N_8172,N_7036,N_7471);
and U8173 (N_8173,N_7789,N_6940);
or U8174 (N_8174,N_6967,N_6117);
and U8175 (N_8175,N_7743,N_6193);
and U8176 (N_8176,N_7139,N_7366);
nor U8177 (N_8177,N_7900,N_6757);
nand U8178 (N_8178,N_7945,N_7811);
nor U8179 (N_8179,N_6951,N_7045);
or U8180 (N_8180,N_6708,N_6105);
nor U8181 (N_8181,N_6731,N_7874);
nand U8182 (N_8182,N_6900,N_6531);
nor U8183 (N_8183,N_7502,N_6484);
or U8184 (N_8184,N_6805,N_6779);
nand U8185 (N_8185,N_7084,N_7622);
nand U8186 (N_8186,N_7467,N_6654);
nor U8187 (N_8187,N_6519,N_6661);
xor U8188 (N_8188,N_6655,N_6038);
or U8189 (N_8189,N_7951,N_7305);
nand U8190 (N_8190,N_7242,N_6310);
nor U8191 (N_8191,N_7880,N_7696);
and U8192 (N_8192,N_6221,N_7763);
or U8193 (N_8193,N_7753,N_6851);
and U8194 (N_8194,N_6504,N_6278);
nor U8195 (N_8195,N_6284,N_6134);
nor U8196 (N_8196,N_7433,N_6819);
xor U8197 (N_8197,N_7484,N_7895);
nand U8198 (N_8198,N_7905,N_7854);
xor U8199 (N_8199,N_7372,N_6170);
nand U8200 (N_8200,N_6996,N_6141);
xor U8201 (N_8201,N_6691,N_7942);
nand U8202 (N_8202,N_6931,N_6279);
and U8203 (N_8203,N_6335,N_6896);
and U8204 (N_8204,N_7509,N_7689);
or U8205 (N_8205,N_7448,N_7913);
xnor U8206 (N_8206,N_7348,N_7210);
and U8207 (N_8207,N_6281,N_6299);
or U8208 (N_8208,N_7394,N_7812);
or U8209 (N_8209,N_6349,N_7131);
nor U8210 (N_8210,N_7482,N_6036);
xor U8211 (N_8211,N_6441,N_7284);
nor U8212 (N_8212,N_7363,N_7059);
and U8213 (N_8213,N_6131,N_7489);
or U8214 (N_8214,N_6506,N_7940);
nand U8215 (N_8215,N_6574,N_7774);
or U8216 (N_8216,N_6501,N_7540);
nand U8217 (N_8217,N_6791,N_6540);
and U8218 (N_8218,N_6497,N_7508);
or U8219 (N_8219,N_7670,N_7416);
xnor U8220 (N_8220,N_6128,N_6844);
xor U8221 (N_8221,N_7659,N_6937);
nor U8222 (N_8222,N_7449,N_6741);
nand U8223 (N_8223,N_6876,N_7883);
or U8224 (N_8224,N_6670,N_6818);
nand U8225 (N_8225,N_7587,N_6054);
and U8226 (N_8226,N_6780,N_6346);
nor U8227 (N_8227,N_7447,N_7571);
xnor U8228 (N_8228,N_7308,N_6229);
nor U8229 (N_8229,N_6838,N_7949);
and U8230 (N_8230,N_7232,N_6725);
xnor U8231 (N_8231,N_7761,N_7970);
nor U8232 (N_8232,N_7155,N_7716);
and U8233 (N_8233,N_7759,N_7343);
xor U8234 (N_8234,N_7717,N_6928);
and U8235 (N_8235,N_6474,N_6253);
nand U8236 (N_8236,N_7154,N_6114);
or U8237 (N_8237,N_7156,N_6008);
or U8238 (N_8238,N_6460,N_6516);
xnor U8239 (N_8239,N_6006,N_6622);
and U8240 (N_8240,N_6062,N_6201);
or U8241 (N_8241,N_6313,N_6628);
xor U8242 (N_8242,N_6216,N_6700);
nand U8243 (N_8243,N_6009,N_6404);
nand U8244 (N_8244,N_6625,N_7307);
xnor U8245 (N_8245,N_6130,N_7543);
nand U8246 (N_8246,N_6910,N_7123);
nor U8247 (N_8247,N_6398,N_6776);
or U8248 (N_8248,N_7046,N_6396);
nor U8249 (N_8249,N_6297,N_6030);
nor U8250 (N_8250,N_7922,N_6695);
or U8251 (N_8251,N_6589,N_7632);
or U8252 (N_8252,N_6245,N_7251);
or U8253 (N_8253,N_7846,N_7920);
nand U8254 (N_8254,N_6645,N_6895);
and U8255 (N_8255,N_7236,N_7560);
xor U8256 (N_8256,N_6934,N_7345);
xnor U8257 (N_8257,N_7576,N_7687);
and U8258 (N_8258,N_6942,N_6904);
nor U8259 (N_8259,N_6397,N_7313);
nor U8260 (N_8260,N_6267,N_7672);
or U8261 (N_8261,N_7912,N_6439);
and U8262 (N_8262,N_6961,N_7102);
or U8263 (N_8263,N_7948,N_6386);
or U8264 (N_8264,N_7375,N_7315);
and U8265 (N_8265,N_6056,N_6047);
xnor U8266 (N_8266,N_7914,N_7193);
nand U8267 (N_8267,N_6796,N_6448);
nor U8268 (N_8268,N_7092,N_7054);
nand U8269 (N_8269,N_7396,N_7071);
and U8270 (N_8270,N_7398,N_7603);
nor U8271 (N_8271,N_6594,N_6321);
or U8272 (N_8272,N_6202,N_7849);
and U8273 (N_8273,N_6019,N_6826);
nand U8274 (N_8274,N_6956,N_7785);
or U8275 (N_8275,N_7009,N_6073);
nor U8276 (N_8276,N_6852,N_6751);
or U8277 (N_8277,N_6798,N_6687);
or U8278 (N_8278,N_6472,N_6771);
nor U8279 (N_8279,N_6809,N_6560);
and U8280 (N_8280,N_6939,N_6033);
nor U8281 (N_8281,N_6761,N_7941);
or U8282 (N_8282,N_7051,N_6945);
nand U8283 (N_8283,N_7816,N_7146);
xnor U8284 (N_8284,N_6786,N_6638);
and U8285 (N_8285,N_6116,N_6643);
xor U8286 (N_8286,N_7124,N_6273);
nor U8287 (N_8287,N_7786,N_6790);
and U8288 (N_8288,N_7598,N_6338);
xor U8289 (N_8289,N_6582,N_6877);
and U8290 (N_8290,N_7095,N_7454);
or U8291 (N_8291,N_7637,N_6133);
nand U8292 (N_8292,N_7808,N_7220);
nor U8293 (N_8293,N_6572,N_6763);
xnor U8294 (N_8294,N_6403,N_6517);
nand U8295 (N_8295,N_6802,N_7192);
or U8296 (N_8296,N_6287,N_6525);
or U8297 (N_8297,N_6494,N_6584);
nand U8298 (N_8298,N_7311,N_6620);
nor U8299 (N_8299,N_7058,N_6181);
nand U8300 (N_8300,N_6657,N_7612);
xnor U8301 (N_8301,N_6259,N_6552);
or U8302 (N_8302,N_7041,N_7017);
and U8303 (N_8303,N_7392,N_7830);
xnor U8304 (N_8304,N_6830,N_7474);
nor U8305 (N_8305,N_7184,N_6684);
xor U8306 (N_8306,N_6483,N_6750);
nor U8307 (N_8307,N_6973,N_7048);
nand U8308 (N_8308,N_6612,N_6171);
nand U8309 (N_8309,N_7128,N_6300);
or U8310 (N_8310,N_7676,N_6135);
or U8311 (N_8311,N_6018,N_7455);
and U8312 (N_8312,N_6094,N_7821);
and U8313 (N_8313,N_6129,N_7856);
or U8314 (N_8314,N_6465,N_7395);
nor U8315 (N_8315,N_7053,N_6041);
and U8316 (N_8316,N_7399,N_6853);
and U8317 (N_8317,N_7421,N_6892);
xnor U8318 (N_8318,N_6077,N_7459);
xnor U8319 (N_8319,N_6797,N_6343);
and U8320 (N_8320,N_6424,N_7807);
nand U8321 (N_8321,N_6345,N_6344);
and U8322 (N_8322,N_6807,N_6639);
xnor U8323 (N_8323,N_6562,N_6784);
nand U8324 (N_8324,N_7780,N_6082);
and U8325 (N_8325,N_6319,N_7625);
nand U8326 (N_8326,N_7228,N_6280);
xor U8327 (N_8327,N_7446,N_6723);
and U8328 (N_8328,N_6162,N_6488);
nor U8329 (N_8329,N_7314,N_7056);
or U8330 (N_8330,N_7390,N_7475);
xor U8331 (N_8331,N_6551,N_6804);
xor U8332 (N_8332,N_6012,N_7965);
nor U8333 (N_8333,N_7173,N_7641);
nand U8334 (N_8334,N_7257,N_7294);
nor U8335 (N_8335,N_6553,N_7835);
or U8336 (N_8336,N_7726,N_6524);
xor U8337 (N_8337,N_7279,N_7277);
and U8338 (N_8338,N_6409,N_6156);
xor U8339 (N_8339,N_7408,N_6461);
xor U8340 (N_8340,N_6586,N_7091);
nor U8341 (N_8341,N_7096,N_6936);
and U8342 (N_8342,N_7911,N_7638);
nor U8343 (N_8343,N_7840,N_7073);
xnor U8344 (N_8344,N_7403,N_6159);
and U8345 (N_8345,N_7736,N_6611);
and U8346 (N_8346,N_7297,N_7081);
nor U8347 (N_8347,N_6682,N_7094);
and U8348 (N_8348,N_7797,N_6822);
xnor U8349 (N_8349,N_6587,N_7778);
nor U8350 (N_8350,N_7909,N_7718);
and U8351 (N_8351,N_6575,N_7722);
and U8352 (N_8352,N_6414,N_7099);
nand U8353 (N_8353,N_7330,N_6847);
nor U8354 (N_8354,N_7212,N_6833);
nor U8355 (N_8355,N_6107,N_7916);
and U8356 (N_8356,N_7032,N_7562);
xor U8357 (N_8357,N_7214,N_7651);
nor U8358 (N_8358,N_6099,N_7993);
or U8359 (N_8359,N_6801,N_6095);
nor U8360 (N_8360,N_6864,N_7510);
xor U8361 (N_8361,N_6558,N_6863);
nor U8362 (N_8362,N_7768,N_6873);
nand U8363 (N_8363,N_6971,N_6240);
and U8364 (N_8364,N_6331,N_6473);
or U8365 (N_8365,N_6435,N_7354);
nor U8366 (N_8366,N_7042,N_6658);
xor U8367 (N_8367,N_6430,N_7112);
or U8368 (N_8368,N_6055,N_7983);
nor U8369 (N_8369,N_7608,N_7190);
xor U8370 (N_8370,N_7665,N_6870);
nand U8371 (N_8371,N_7741,N_7319);
xnor U8372 (N_8372,N_7133,N_7715);
nor U8373 (N_8373,N_6362,N_6220);
or U8374 (N_8374,N_7181,N_7271);
or U8375 (N_8375,N_6475,N_7964);
or U8376 (N_8376,N_6485,N_7530);
and U8377 (N_8377,N_7501,N_7737);
xor U8378 (N_8378,N_6775,N_6462);
xnor U8379 (N_8379,N_7140,N_6566);
xor U8380 (N_8380,N_7125,N_6518);
nor U8381 (N_8381,N_7152,N_6182);
nor U8382 (N_8382,N_6913,N_6856);
xnor U8383 (N_8383,N_6539,N_6044);
and U8384 (N_8384,N_7578,N_6231);
xor U8385 (N_8385,N_6571,N_6326);
nand U8386 (N_8386,N_6511,N_7443);
nor U8387 (N_8387,N_6227,N_6767);
nand U8388 (N_8388,N_7005,N_6537);
nand U8389 (N_8389,N_7436,N_6263);
and U8390 (N_8390,N_6466,N_7148);
nand U8391 (N_8391,N_7269,N_7425);
xor U8392 (N_8392,N_6613,N_6093);
xor U8393 (N_8393,N_6538,N_7230);
or U8394 (N_8394,N_7115,N_6302);
and U8395 (N_8395,N_7287,N_6123);
xnor U8396 (N_8396,N_7019,N_7438);
xnor U8397 (N_8397,N_6680,N_7727);
xnor U8398 (N_8398,N_6831,N_6179);
xnor U8399 (N_8399,N_7777,N_7799);
nor U8400 (N_8400,N_7801,N_7052);
xnor U8401 (N_8401,N_7851,N_6384);
nand U8402 (N_8402,N_7130,N_7767);
nand U8403 (N_8403,N_7616,N_6421);
xor U8404 (N_8404,N_6512,N_6887);
nor U8405 (N_8405,N_7100,N_7011);
or U8406 (N_8406,N_6908,N_6758);
nand U8407 (N_8407,N_6533,N_7357);
and U8408 (N_8408,N_7231,N_7003);
and U8409 (N_8409,N_7008,N_6604);
xnor U8410 (N_8410,N_7580,N_6455);
nand U8411 (N_8411,N_7302,N_7289);
or U8412 (N_8412,N_6438,N_6555);
nor U8413 (N_8413,N_6214,N_6585);
or U8414 (N_8414,N_7189,N_6624);
nand U8415 (N_8415,N_6621,N_7884);
xnor U8416 (N_8416,N_6510,N_6211);
and U8417 (N_8417,N_7966,N_6148);
nor U8418 (N_8418,N_7928,N_7491);
and U8419 (N_8419,N_7567,N_7273);
and U8420 (N_8420,N_6209,N_7953);
or U8421 (N_8421,N_6916,N_6161);
xor U8422 (N_8422,N_7684,N_7719);
xnor U8423 (N_8423,N_6672,N_7740);
xor U8424 (N_8424,N_6557,N_7018);
xor U8425 (N_8425,N_7222,N_6489);
xor U8426 (N_8426,N_7175,N_6958);
nand U8427 (N_8427,N_7998,N_7171);
and U8428 (N_8428,N_6001,N_7020);
or U8429 (N_8429,N_7944,N_6158);
nand U8430 (N_8430,N_6121,N_7291);
or U8431 (N_8431,N_6683,N_7623);
or U8432 (N_8432,N_6549,N_7721);
nand U8433 (N_8433,N_7177,N_6964);
and U8434 (N_8434,N_6868,N_6696);
nand U8435 (N_8435,N_6126,N_6678);
xnor U8436 (N_8436,N_6422,N_7605);
nor U8437 (N_8437,N_7134,N_6641);
or U8438 (N_8438,N_6888,N_7592);
or U8439 (N_8439,N_7957,N_6219);
or U8440 (N_8440,N_7034,N_7423);
nand U8441 (N_8441,N_6799,N_7364);
and U8442 (N_8442,N_7602,N_6406);
and U8443 (N_8443,N_6734,N_7946);
nor U8444 (N_8444,N_6254,N_6860);
xnor U8445 (N_8445,N_7186,N_6596);
xor U8446 (N_8446,N_6013,N_6879);
xnor U8447 (N_8447,N_6334,N_7633);
xor U8448 (N_8448,N_6238,N_7182);
nand U8449 (N_8449,N_6354,N_6630);
xor U8450 (N_8450,N_7028,N_7648);
nand U8451 (N_8451,N_7904,N_6995);
nor U8452 (N_8452,N_6050,N_7188);
xor U8453 (N_8453,N_6187,N_7206);
or U8454 (N_8454,N_7557,N_7143);
and U8455 (N_8455,N_6842,N_6999);
or U8456 (N_8456,N_6667,N_7582);
and U8457 (N_8457,N_7855,N_7006);
nand U8458 (N_8458,N_7686,N_7295);
xor U8459 (N_8459,N_7323,N_7620);
xnor U8460 (N_8460,N_6541,N_7035);
xnor U8461 (N_8461,N_6993,N_6043);
or U8462 (N_8462,N_6481,N_6634);
or U8463 (N_8463,N_7158,N_7187);
or U8464 (N_8464,N_7336,N_7321);
or U8465 (N_8465,N_7857,N_7551);
and U8466 (N_8466,N_6642,N_7478);
nor U8467 (N_8467,N_6663,N_6291);
xor U8468 (N_8468,N_6391,N_7611);
and U8469 (N_8469,N_6234,N_7453);
and U8470 (N_8470,N_6754,N_7800);
nand U8471 (N_8471,N_7419,N_6721);
and U8472 (N_8472,N_6320,N_6173);
nor U8473 (N_8473,N_6283,N_7658);
or U8474 (N_8474,N_6762,N_7590);
xnor U8475 (N_8475,N_7699,N_6556);
and U8476 (N_8476,N_7528,N_6003);
nor U8477 (N_8477,N_7109,N_7978);
nand U8478 (N_8478,N_7457,N_7068);
xnor U8479 (N_8479,N_6699,N_7040);
nand U8480 (N_8480,N_7404,N_6016);
nand U8481 (N_8481,N_6314,N_7280);
nor U8482 (N_8482,N_7629,N_6498);
xor U8483 (N_8483,N_6565,N_7397);
nor U8484 (N_8484,N_7299,N_7713);
nand U8485 (N_8485,N_6294,N_6608);
or U8486 (N_8486,N_7465,N_6318);
nor U8487 (N_8487,N_6972,N_7456);
xor U8488 (N_8488,N_6228,N_7561);
xor U8489 (N_8489,N_7380,N_6416);
nand U8490 (N_8490,N_7371,N_6676);
nand U8491 (N_8491,N_6078,N_6163);
nand U8492 (N_8492,N_7274,N_7167);
and U8493 (N_8493,N_7031,N_7701);
or U8494 (N_8494,N_7923,N_7349);
and U8495 (N_8495,N_7064,N_7827);
xor U8496 (N_8496,N_6881,N_6266);
nand U8497 (N_8497,N_6370,N_6812);
or U8498 (N_8498,N_6532,N_7150);
or U8499 (N_8499,N_6208,N_7538);
nor U8500 (N_8500,N_7987,N_7639);
and U8501 (N_8501,N_7203,N_6295);
or U8502 (N_8502,N_7168,N_6233);
or U8503 (N_8503,N_7432,N_6479);
xnor U8504 (N_8504,N_6901,N_6875);
nand U8505 (N_8505,N_6379,N_7434);
or U8506 (N_8506,N_6898,N_6204);
and U8507 (N_8507,N_6177,N_7116);
xor U8508 (N_8508,N_6692,N_7534);
and U8509 (N_8509,N_7548,N_7706);
nand U8510 (N_8510,N_7037,N_7969);
xnor U8511 (N_8511,N_6180,N_6534);
nor U8512 (N_8512,N_6919,N_7959);
nor U8513 (N_8513,N_6415,N_7858);
nand U8514 (N_8514,N_7374,N_7239);
or U8515 (N_8515,N_6769,N_6905);
and U8516 (N_8516,N_7907,N_7930);
nor U8517 (N_8517,N_7283,N_6495);
nor U8518 (N_8518,N_6787,N_6015);
and U8519 (N_8519,N_7332,N_6470);
and U8520 (N_8520,N_6535,N_7669);
nor U8521 (N_8521,N_7194,N_6167);
or U8522 (N_8522,N_6962,N_7926);
or U8523 (N_8523,N_7873,N_7979);
or U8524 (N_8524,N_6954,N_7877);
nand U8525 (N_8525,N_7346,N_6070);
nand U8526 (N_8526,N_6122,N_6669);
and U8527 (N_8527,N_6736,N_6647);
xor U8528 (N_8528,N_7468,N_6248);
or U8529 (N_8529,N_7872,N_7831);
or U8530 (N_8530,N_6559,N_6867);
nand U8531 (N_8531,N_6085,N_7981);
nand U8532 (N_8532,N_7896,N_6189);
and U8533 (N_8533,N_6332,N_6328);
and U8534 (N_8534,N_7268,N_7248);
nor U8535 (N_8535,N_7890,N_7876);
or U8536 (N_8536,N_7065,N_7205);
or U8537 (N_8537,N_6000,N_7818);
xor U8538 (N_8538,N_7244,N_6927);
or U8539 (N_8539,N_7640,N_7272);
or U8540 (N_8540,N_7929,N_7180);
nand U8541 (N_8541,N_7568,N_7420);
and U8542 (N_8542,N_7300,N_7472);
or U8543 (N_8543,N_6453,N_6137);
nor U8544 (N_8544,N_6022,N_7062);
nor U8545 (N_8545,N_6688,N_7650);
and U8546 (N_8546,N_6004,N_6718);
and U8547 (N_8547,N_7645,N_7990);
xnor U8548 (N_8548,N_6528,N_7674);
or U8549 (N_8549,N_7141,N_7381);
xnor U8550 (N_8550,N_7865,N_7255);
nor U8551 (N_8551,N_6268,N_7809);
or U8552 (N_8552,N_6811,N_6045);
nand U8553 (N_8553,N_7225,N_7373);
xor U8554 (N_8554,N_7137,N_7524);
xnor U8555 (N_8555,N_7039,N_6862);
and U8556 (N_8556,N_6413,N_7958);
nor U8557 (N_8557,N_7085,N_6324);
or U8558 (N_8558,N_6074,N_7417);
nand U8559 (N_8559,N_6388,N_6327);
xnor U8560 (N_8560,N_7026,N_7772);
nor U8561 (N_8561,N_7550,N_7376);
nor U8562 (N_8562,N_6783,N_7089);
nor U8563 (N_8563,N_7451,N_7022);
xor U8564 (N_8564,N_7573,N_6190);
and U8565 (N_8565,N_6650,N_6719);
and U8566 (N_8566,N_6183,N_7704);
or U8567 (N_8567,N_7480,N_7841);
xnor U8568 (N_8568,N_6270,N_7898);
or U8569 (N_8569,N_7379,N_6859);
xnor U8570 (N_8570,N_6247,N_7720);
xor U8571 (N_8571,N_6735,N_6759);
nor U8572 (N_8572,N_6858,N_7747);
nor U8573 (N_8573,N_6428,N_6990);
nand U8574 (N_8574,N_7149,N_7588);
or U8575 (N_8575,N_6289,N_6941);
nor U8576 (N_8576,N_6322,N_6977);
and U8577 (N_8577,N_6476,N_7795);
nor U8578 (N_8578,N_6154,N_7878);
nand U8579 (N_8579,N_6184,N_6017);
and U8580 (N_8580,N_7703,N_7108);
or U8581 (N_8581,N_6947,N_7791);
nand U8582 (N_8582,N_6909,N_7207);
nand U8583 (N_8583,N_7725,N_6897);
xor U8584 (N_8584,N_7229,N_6843);
nor U8585 (N_8585,N_7326,N_7521);
xor U8586 (N_8586,N_6733,N_7276);
or U8587 (N_8587,N_6306,N_7523);
nand U8588 (N_8588,N_6742,N_6770);
nand U8589 (N_8589,N_7581,N_7679);
or U8590 (N_8590,N_6350,N_7264);
or U8591 (N_8591,N_7698,N_7015);
nand U8592 (N_8592,N_7544,N_6800);
nand U8593 (N_8593,N_6994,N_7243);
nand U8594 (N_8594,N_7466,N_7402);
nand U8595 (N_8595,N_7844,N_7262);
nand U8596 (N_8596,N_7729,N_6269);
and U8597 (N_8597,N_6412,N_7216);
nand U8598 (N_8598,N_7077,N_6458);
and U8599 (N_8599,N_6339,N_7126);
xor U8600 (N_8600,N_7897,N_6264);
nor U8601 (N_8601,N_6106,N_6697);
nand U8602 (N_8602,N_6542,N_6025);
xnor U8603 (N_8603,N_6026,N_6353);
xnor U8604 (N_8604,N_7921,N_6720);
nand U8605 (N_8605,N_6813,N_6726);
nor U8606 (N_8606,N_6514,N_7546);
or U8607 (N_8607,N_7164,N_6296);
nor U8608 (N_8608,N_7080,N_6186);
and U8609 (N_8609,N_6857,N_6823);
or U8610 (N_8610,N_7606,N_7903);
and U8611 (N_8611,N_6573,N_6119);
nor U8612 (N_8612,N_6616,N_6617);
xnor U8613 (N_8613,N_6609,N_6503);
xor U8614 (N_8614,N_6832,N_6480);
and U8615 (N_8615,N_7850,N_6405);
xnor U8616 (N_8616,N_6285,N_7882);
xor U8617 (N_8617,N_6188,N_6290);
nand U8618 (N_8618,N_7867,N_6615);
nor U8619 (N_8619,N_6023,N_6920);
nand U8620 (N_8620,N_6633,N_7430);
nand U8621 (N_8621,N_6275,N_7529);
nor U8622 (N_8622,N_6793,N_6564);
nand U8623 (N_8623,N_7004,N_6457);
and U8624 (N_8624,N_6974,N_7862);
nor U8625 (N_8625,N_7604,N_6076);
and U8626 (N_8626,N_7010,N_6745);
nor U8627 (N_8627,N_6578,N_7781);
and U8628 (N_8628,N_6378,N_7353);
and U8629 (N_8629,N_7925,N_7224);
or U8630 (N_8630,N_6526,N_6712);
nor U8631 (N_8631,N_6175,N_7825);
or U8632 (N_8632,N_7770,N_7515);
nand U8633 (N_8633,N_6252,N_6966);
and U8634 (N_8634,N_6103,N_7938);
and U8635 (N_8635,N_6143,N_6390);
nor U8636 (N_8636,N_6239,N_7083);
or U8637 (N_8637,N_6922,N_6102);
or U8638 (N_8638,N_7814,N_6301);
or U8639 (N_8639,N_6677,N_6768);
xnor U8640 (N_8640,N_6850,N_6459);
nor U8641 (N_8641,N_6385,N_7599);
nand U8642 (N_8642,N_7179,N_6124);
nand U8643 (N_8643,N_7113,N_7162);
and U8644 (N_8644,N_6991,N_6410);
nand U8645 (N_8645,N_6399,N_6444);
xnor U8646 (N_8646,N_6288,N_6058);
nand U8647 (N_8647,N_6629,N_6963);
and U8648 (N_8648,N_6948,N_7117);
or U8649 (N_8649,N_6808,N_7120);
and U8650 (N_8650,N_7834,N_6086);
nand U8651 (N_8651,N_6810,N_6442);
xor U8652 (N_8652,N_7050,N_6943);
xnor U8653 (N_8653,N_7919,N_7200);
nor U8654 (N_8654,N_6059,N_6303);
nand U8655 (N_8655,N_7823,N_7090);
xnor U8656 (N_8656,N_7352,N_7499);
nand U8657 (N_8657,N_6400,N_7127);
or U8658 (N_8658,N_6855,N_6849);
or U8659 (N_8659,N_6981,N_6536);
nand U8660 (N_8660,N_6081,N_7306);
nand U8661 (N_8661,N_7424,N_6165);
nand U8662 (N_8662,N_7918,N_6717);
nand U8663 (N_8663,N_7078,N_6363);
or U8664 (N_8664,N_6153,N_7441);
nand U8665 (N_8665,N_6311,N_7191);
nor U8666 (N_8666,N_7174,N_7245);
or U8667 (N_8667,N_6308,N_7428);
and U8668 (N_8668,N_6032,N_7413);
nand U8669 (N_8669,N_7683,N_6393);
and U8670 (N_8670,N_7776,N_6491);
xnor U8671 (N_8671,N_7748,N_7237);
or U8672 (N_8672,N_6886,N_7752);
xor U8673 (N_8673,N_6090,N_6020);
nor U8674 (N_8674,N_7871,N_7732);
xnor U8675 (N_8675,N_7261,N_7247);
or U8676 (N_8676,N_7542,N_7384);
or U8677 (N_8677,N_7057,N_6431);
nand U8678 (N_8678,N_7647,N_6730);
nor U8679 (N_8679,N_6902,N_6640);
or U8680 (N_8680,N_6727,N_7498);
or U8681 (N_8681,N_6241,N_6172);
or U8682 (N_8682,N_7129,N_7044);
nand U8683 (N_8683,N_6487,N_7001);
and U8684 (N_8684,N_7845,N_7119);
or U8685 (N_8685,N_7462,N_7655);
xor U8686 (N_8686,N_6637,N_6356);
or U8687 (N_8687,N_6145,N_7577);
or U8688 (N_8688,N_6773,N_6772);
and U8689 (N_8689,N_7060,N_6010);
nand U8690 (N_8690,N_7889,N_7114);
or U8691 (N_8691,N_7702,N_6871);
nor U8692 (N_8692,N_6490,N_7318);
or U8693 (N_8693,N_7997,N_7757);
or U8694 (N_8694,N_6738,N_7163);
nand U8695 (N_8695,N_7769,N_6706);
or U8696 (N_8696,N_7439,N_7490);
or U8697 (N_8697,N_6282,N_7226);
nand U8698 (N_8698,N_7157,N_6230);
or U8699 (N_8699,N_6703,N_6732);
nor U8700 (N_8700,N_6869,N_6606);
xor U8701 (N_8701,N_6011,N_6452);
nand U8702 (N_8702,N_6164,N_7301);
or U8703 (N_8703,N_6515,N_6361);
and U8704 (N_8704,N_7335,N_6040);
xor U8705 (N_8705,N_7429,N_6563);
or U8706 (N_8706,N_6185,N_7233);
and U8707 (N_8707,N_7803,N_6369);
xnor U8708 (N_8708,N_6599,N_7771);
nand U8709 (N_8709,N_7145,N_6705);
nor U8710 (N_8710,N_6778,N_7464);
or U8711 (N_8711,N_6408,N_7503);
nor U8712 (N_8712,N_6419,N_7347);
xnor U8713 (N_8713,N_6307,N_7074);
nor U8714 (N_8714,N_6664,N_7418);
xnor U8715 (N_8715,N_7506,N_6046);
nand U8716 (N_8716,N_7554,N_6456);
nand U8717 (N_8717,N_7107,N_7525);
and U8718 (N_8718,N_6337,N_6110);
xnor U8719 (N_8719,N_7848,N_6890);
or U8720 (N_8720,N_7246,N_7290);
nor U8721 (N_8721,N_7520,N_7198);
nor U8722 (N_8722,N_7838,N_6260);
and U8723 (N_8723,N_6933,N_7170);
or U8724 (N_8724,N_6236,N_6834);
nand U8725 (N_8725,N_7915,N_6598);
or U8726 (N_8726,N_7160,N_6447);
xor U8727 (N_8727,N_6965,N_7709);
nor U8728 (N_8728,N_6340,N_6146);
and U8729 (N_8729,N_6618,N_6652);
nand U8730 (N_8730,N_6502,N_6998);
or U8731 (N_8731,N_7613,N_7852);
or U8732 (N_8732,N_6500,N_7906);
nand U8733 (N_8733,N_7541,N_6716);
and U8734 (N_8734,N_7975,N_7794);
nand U8735 (N_8735,N_6372,N_6884);
xnor U8736 (N_8736,N_7388,N_7427);
nor U8737 (N_8737,N_7458,N_7298);
nand U8738 (N_8738,N_6374,N_6980);
nor U8739 (N_8739,N_7526,N_7894);
and U8740 (N_8740,N_6191,N_6142);
nand U8741 (N_8741,N_7917,N_6883);
nand U8742 (N_8742,N_6333,N_7278);
or U8743 (N_8743,N_6530,N_6080);
nand U8744 (N_8744,N_6246,N_7104);
xnor U8745 (N_8745,N_7470,N_7185);
and U8746 (N_8746,N_6944,N_6147);
nand U8747 (N_8747,N_7351,N_6632);
and U8748 (N_8748,N_6341,N_6878);
nand U8749 (N_8749,N_6923,N_6237);
or U8750 (N_8750,N_6464,N_7517);
or U8751 (N_8751,N_6561,N_6915);
nand U8752 (N_8752,N_6646,N_7549);
or U8753 (N_8753,N_7007,N_7805);
nand U8754 (N_8754,N_6166,N_6568);
nor U8755 (N_8755,N_7383,N_7386);
and U8756 (N_8756,N_7266,N_7654);
nor U8757 (N_8757,N_7505,N_6739);
xor U8758 (N_8758,N_6978,N_6366);
or U8759 (N_8759,N_6891,N_7931);
and U8760 (N_8760,N_7493,N_7545);
or U8761 (N_8761,N_6803,N_6911);
nor U8762 (N_8762,N_7910,N_7492);
xor U8763 (N_8763,N_6781,N_7766);
and U8764 (N_8764,N_7365,N_6651);
nand U8765 (N_8765,N_6168,N_6101);
xor U8766 (N_8766,N_7121,N_6679);
or U8767 (N_8767,N_7218,N_6546);
or U8768 (N_8768,N_6242,N_6747);
nor U8769 (N_8769,N_7547,N_6312);
nor U8770 (N_8770,N_7461,N_6665);
or U8771 (N_8771,N_7341,N_6946);
or U8772 (N_8772,N_7219,N_6605);
and U8773 (N_8773,N_7728,N_6623);
nor U8774 (N_8774,N_7111,N_6261);
or U8775 (N_8775,N_7790,N_6249);
nand U8776 (N_8776,N_6034,N_7643);
nor U8777 (N_8777,N_6764,N_6380);
or U8778 (N_8778,N_7615,N_6499);
xor U8779 (N_8779,N_6674,N_7355);
nand U8780 (N_8780,N_6950,N_7486);
and U8781 (N_8781,N_7215,N_6816);
and U8782 (N_8782,N_6097,N_7553);
xnor U8783 (N_8783,N_7815,N_7869);
xor U8784 (N_8784,N_6777,N_7485);
or U8785 (N_8785,N_7511,N_6429);
xnor U8786 (N_8786,N_7367,N_7552);
nor U8787 (N_8787,N_7569,N_6376);
nor U8788 (N_8788,N_7440,N_6120);
or U8789 (N_8789,N_7859,N_6600);
or U8790 (N_8790,N_6899,N_6997);
and U8791 (N_8791,N_7745,N_7565);
nand U8792 (N_8792,N_6061,N_6662);
and U8793 (N_8793,N_6841,N_6690);
nand U8794 (N_8794,N_6256,N_6960);
xnor U8795 (N_8795,N_7764,N_6602);
and U8796 (N_8796,N_6364,N_7888);
and U8797 (N_8797,N_6149,N_6198);
or U8798 (N_8798,N_6521,N_7055);
xnor U8799 (N_8799,N_7988,N_6785);
or U8800 (N_8800,N_7452,N_6118);
and U8801 (N_8801,N_7079,N_7937);
xnor U8802 (N_8802,N_7176,N_7025);
or U8803 (N_8803,N_7537,N_6358);
nor U8804 (N_8804,N_7924,N_7494);
xor U8805 (N_8805,N_7316,N_6486);
xor U8806 (N_8806,N_6970,N_6724);
nand U8807 (N_8807,N_7197,N_7819);
and U8808 (N_8808,N_6707,N_6825);
or U8809 (N_8809,N_6276,N_7566);
xnor U8810 (N_8810,N_7002,N_7558);
xor U8811 (N_8811,N_7980,N_7784);
and U8812 (N_8812,N_6192,N_7512);
or U8813 (N_8813,N_7309,N_7033);
or U8814 (N_8814,N_7559,N_7656);
and U8815 (N_8815,N_7829,N_7668);
xnor U8816 (N_8816,N_6597,N_7513);
xnor U8817 (N_8817,N_7594,N_7358);
and U8818 (N_8818,N_7360,N_6918);
nand U8819 (N_8819,N_6782,N_7773);
or U8820 (N_8820,N_7680,N_6523);
nand U8821 (N_8821,N_7644,N_7240);
xor U8822 (N_8822,N_7675,N_6636);
xnor U8823 (N_8823,N_6477,N_6774);
and U8824 (N_8824,N_6788,N_7460);
xnor U8825 (N_8825,N_6914,N_7864);
xnor U8826 (N_8826,N_6681,N_7972);
or U8827 (N_8827,N_7607,N_7833);
and U8828 (N_8828,N_6792,N_6427);
xor U8829 (N_8829,N_7406,N_7101);
and U8830 (N_8830,N_7961,N_7296);
and U8831 (N_8831,N_7555,N_7708);
xnor U8832 (N_8832,N_6872,N_7731);
nand U8833 (N_8833,N_6508,N_7227);
or U8834 (N_8834,N_6109,N_6554);
and U8835 (N_8835,N_6037,N_6938);
xnor U8836 (N_8836,N_7595,N_7023);
nor U8837 (N_8837,N_7749,N_6806);
nor U8838 (N_8838,N_7442,N_6024);
xnor U8839 (N_8839,N_6063,N_7252);
nand U8840 (N_8840,N_6049,N_7681);
nor U8841 (N_8841,N_6232,N_7739);
nand U8842 (N_8842,N_6746,N_7070);
and U8843 (N_8843,N_7106,N_6251);
nand U8844 (N_8844,N_6213,N_7619);
or U8845 (N_8845,N_7901,N_7793);
xnor U8846 (N_8846,N_7320,N_6271);
nor U8847 (N_8847,N_6671,N_6840);
nand U8848 (N_8848,N_7069,N_6436);
or U8849 (N_8849,N_6309,N_7596);
nand U8850 (N_8850,N_6360,N_6152);
xor U8851 (N_8851,N_7217,N_7281);
xor U8852 (N_8852,N_6685,N_7853);
nor U8853 (N_8853,N_6053,N_7707);
xnor U8854 (N_8854,N_7151,N_7047);
or U8855 (N_8855,N_6467,N_7824);
nand U8856 (N_8856,N_7118,N_6478);
xnor U8857 (N_8857,N_6352,N_6930);
xor U8858 (N_8858,N_7519,N_6244);
or U8859 (N_8859,N_7086,N_6626);
xnor U8860 (N_8860,N_6005,N_6426);
nor U8861 (N_8861,N_7685,N_6420);
xor U8862 (N_8862,N_6548,N_7996);
nor U8863 (N_8863,N_7673,N_6986);
nor U8864 (N_8864,N_6854,N_7660);
nor U8865 (N_8865,N_7826,N_7657);
nand U8866 (N_8866,N_7642,N_7043);
nand U8867 (N_8867,N_6347,N_6160);
or U8868 (N_8868,N_7013,N_6418);
xor U8869 (N_8869,N_7340,N_6635);
or U8870 (N_8870,N_7213,N_7312);
nand U8871 (N_8871,N_6357,N_6505);
nand U8872 (N_8872,N_7391,N_7628);
and U8873 (N_8873,N_6048,N_7267);
nand U8874 (N_8874,N_7235,N_6451);
and U8875 (N_8875,N_6912,N_6257);
nand U8876 (N_8876,N_7792,N_7208);
nand U8877 (N_8877,N_6417,N_7693);
and U8878 (N_8878,N_7405,N_6567);
nand U8879 (N_8879,N_7012,N_7407);
xor U8880 (N_8880,N_6075,N_6355);
nor U8881 (N_8881,N_6835,N_7999);
nand U8882 (N_8882,N_7589,N_7649);
xnor U8883 (N_8883,N_7437,N_7762);
nand U8884 (N_8884,N_7258,N_7690);
xnor U8885 (N_8885,N_7286,N_7361);
and U8886 (N_8886,N_6975,N_7344);
nand U8887 (N_8887,N_7671,N_7863);
nand U8888 (N_8888,N_7842,N_7260);
nor U8889 (N_8889,N_7310,N_7984);
nand U8890 (N_8890,N_7813,N_7507);
or U8891 (N_8891,N_6493,N_6817);
or U8892 (N_8892,N_7678,N_6051);
nand U8893 (N_8893,N_7563,N_7275);
and U8894 (N_8894,N_7088,N_6069);
or U8895 (N_8895,N_6423,N_7989);
and U8896 (N_8896,N_6955,N_6150);
and U8897 (N_8897,N_7955,N_6603);
nor U8898 (N_8898,N_6348,N_7382);
nor U8899 (N_8899,N_7285,N_6756);
and U8900 (N_8900,N_7775,N_7412);
nor U8901 (N_8901,N_6949,N_6368);
and U8902 (N_8902,N_7199,N_7067);
nand U8903 (N_8903,N_7804,N_7936);
and U8904 (N_8904,N_7497,N_6513);
nand U8905 (N_8905,N_7463,N_7723);
nand U8906 (N_8906,N_7172,N_7860);
and U8907 (N_8907,N_7735,N_7634);
nor U8908 (N_8908,N_7304,N_6446);
and U8909 (N_8909,N_7947,N_6529);
nor U8910 (N_8910,N_7481,N_6443);
xor U8911 (N_8911,N_6157,N_6298);
and U8912 (N_8912,N_7820,N_6507);
nand U8913 (N_8913,N_6588,N_7389);
and U8914 (N_8914,N_6136,N_7886);
and U8915 (N_8915,N_7974,N_7908);
nor U8916 (N_8916,N_6007,N_7496);
and U8917 (N_8917,N_7952,N_6169);
nand U8918 (N_8918,N_6057,N_7265);
or U8919 (N_8919,N_6711,N_6795);
or U8920 (N_8920,N_7097,N_7532);
nand U8921 (N_8921,N_6277,N_7359);
or U8922 (N_8922,N_6653,N_6648);
nand U8923 (N_8923,N_6701,N_7636);
nand U8924 (N_8924,N_6789,N_7249);
xor U8925 (N_8925,N_7666,N_7254);
and U8926 (N_8926,N_6039,N_7839);
nand U8927 (N_8927,N_6925,N_7303);
nor U8928 (N_8928,N_6336,N_7144);
nor U8929 (N_8929,N_7836,N_7293);
nor U8930 (N_8930,N_7387,N_7806);
nor U8931 (N_8931,N_7934,N_7866);
and U8932 (N_8932,N_6550,N_6092);
or U8933 (N_8933,N_7514,N_6342);
and U8934 (N_8934,N_6744,N_6127);
nor U8935 (N_8935,N_7204,N_7802);
nor U8936 (N_8936,N_7564,N_7337);
xnor U8937 (N_8937,N_6743,N_7356);
nor U8938 (N_8938,N_7832,N_6839);
xnor U8939 (N_8939,N_7610,N_6668);
or U8940 (N_8940,N_7165,N_6395);
and U8941 (N_8941,N_7570,N_7617);
nand U8942 (N_8942,N_7667,N_7292);
xnor U8943 (N_8943,N_7572,N_7196);
or U8944 (N_8944,N_7986,N_7574);
xor U8945 (N_8945,N_6520,N_6760);
nor U8946 (N_8946,N_7535,N_6570);
xor U8947 (N_8947,N_7331,N_6200);
xnor U8948 (N_8948,N_6874,N_6351);
xor U8949 (N_8949,N_7147,N_6728);
and U8950 (N_8950,N_7694,N_6969);
nand U8951 (N_8951,N_6666,N_7082);
xor U8952 (N_8952,N_7339,N_7061);
nor U8953 (N_8953,N_6079,N_6325);
or U8954 (N_8954,N_7742,N_7705);
and U8955 (N_8955,N_6329,N_7322);
xnor U8956 (N_8956,N_6100,N_6509);
or U8957 (N_8957,N_6255,N_7760);
nor U8958 (N_8958,N_7887,N_6377);
or U8959 (N_8959,N_6207,N_7950);
and U8960 (N_8960,N_6072,N_7400);
or U8961 (N_8961,N_6714,N_7758);
or U8962 (N_8962,N_6593,N_7982);
nor U8963 (N_8963,N_6815,N_7751);
and U8964 (N_8964,N_6250,N_6917);
and U8965 (N_8965,N_7935,N_7016);
nor U8966 (N_8966,N_7664,N_7531);
nor U8967 (N_8967,N_7746,N_7136);
or U8968 (N_8968,N_6029,N_7142);
or U8969 (N_8969,N_7902,N_7653);
nand U8970 (N_8970,N_7087,N_6471);
or U8971 (N_8971,N_6893,N_6715);
or U8972 (N_8972,N_7631,N_6713);
or U8973 (N_8973,N_6087,N_7049);
or U8974 (N_8974,N_7614,N_6262);
nand U8975 (N_8975,N_7487,N_6218);
and U8976 (N_8976,N_7201,N_6139);
nand U8977 (N_8977,N_6437,N_7601);
xor U8978 (N_8978,N_6212,N_6592);
xor U8979 (N_8979,N_6889,N_7788);
nor U8980 (N_8980,N_7435,N_6138);
nor U8981 (N_8981,N_6392,N_7476);
or U8982 (N_8982,N_7444,N_7414);
xor U8983 (N_8983,N_7828,N_7822);
and U8984 (N_8984,N_6698,N_7324);
nand U8985 (N_8985,N_6631,N_6827);
nand U8986 (N_8986,N_6381,N_7700);
nand U8987 (N_8987,N_6317,N_6601);
xor U8988 (N_8988,N_7585,N_6068);
xor U8989 (N_8989,N_6861,N_7238);
or U8990 (N_8990,N_6132,N_6694);
or U8991 (N_8991,N_6432,N_7579);
nand U8992 (N_8992,N_7250,N_7024);
nor U8993 (N_8993,N_7159,N_7522);
or U8994 (N_8994,N_6224,N_7431);
or U8995 (N_8995,N_7733,N_7253);
xnor U8996 (N_8996,N_7422,N_6265);
nand U8997 (N_8997,N_7591,N_7415);
nor U8998 (N_8998,N_7593,N_7932);
nor U8999 (N_8999,N_7021,N_7377);
or U9000 (N_9000,N_6273,N_6132);
nor U9001 (N_9001,N_6243,N_6585);
xnor U9002 (N_9002,N_7333,N_7955);
nor U9003 (N_9003,N_6586,N_6711);
nand U9004 (N_9004,N_7637,N_7773);
nor U9005 (N_9005,N_6781,N_6693);
nor U9006 (N_9006,N_7722,N_7475);
xnor U9007 (N_9007,N_6578,N_7432);
or U9008 (N_9008,N_6802,N_6127);
or U9009 (N_9009,N_7802,N_7035);
nand U9010 (N_9010,N_7810,N_6539);
or U9011 (N_9011,N_7705,N_6177);
or U9012 (N_9012,N_7667,N_7029);
nand U9013 (N_9013,N_6393,N_6957);
and U9014 (N_9014,N_7077,N_6812);
or U9015 (N_9015,N_6748,N_7392);
nor U9016 (N_9016,N_6526,N_7406);
nand U9017 (N_9017,N_6972,N_7475);
or U9018 (N_9018,N_6453,N_7129);
and U9019 (N_9019,N_6303,N_6554);
nor U9020 (N_9020,N_7981,N_6342);
nand U9021 (N_9021,N_6081,N_7234);
or U9022 (N_9022,N_7723,N_7365);
nor U9023 (N_9023,N_6136,N_7672);
xor U9024 (N_9024,N_6115,N_6849);
xnor U9025 (N_9025,N_7630,N_6280);
nand U9026 (N_9026,N_6527,N_7188);
nand U9027 (N_9027,N_6034,N_6423);
or U9028 (N_9028,N_7444,N_7714);
or U9029 (N_9029,N_7439,N_7038);
and U9030 (N_9030,N_6990,N_7971);
and U9031 (N_9031,N_6935,N_7910);
nand U9032 (N_9032,N_7741,N_6896);
or U9033 (N_9033,N_6912,N_6989);
nor U9034 (N_9034,N_7821,N_6722);
nor U9035 (N_9035,N_7913,N_6883);
xnor U9036 (N_9036,N_7821,N_6355);
nand U9037 (N_9037,N_7834,N_7643);
nor U9038 (N_9038,N_6445,N_6298);
xnor U9039 (N_9039,N_6244,N_6781);
xor U9040 (N_9040,N_7359,N_6256);
and U9041 (N_9041,N_7849,N_6003);
and U9042 (N_9042,N_6972,N_6838);
xor U9043 (N_9043,N_7150,N_7196);
nand U9044 (N_9044,N_7996,N_6150);
nand U9045 (N_9045,N_7688,N_6035);
xnor U9046 (N_9046,N_7711,N_7027);
nor U9047 (N_9047,N_6670,N_7529);
or U9048 (N_9048,N_6109,N_7999);
nand U9049 (N_9049,N_6409,N_6912);
and U9050 (N_9050,N_7803,N_7077);
xor U9051 (N_9051,N_6333,N_7793);
nor U9052 (N_9052,N_6241,N_7255);
or U9053 (N_9053,N_6270,N_7247);
xnor U9054 (N_9054,N_6445,N_7121);
nand U9055 (N_9055,N_7973,N_7169);
nor U9056 (N_9056,N_7100,N_6792);
nand U9057 (N_9057,N_6326,N_6903);
or U9058 (N_9058,N_6713,N_7052);
nor U9059 (N_9059,N_7211,N_6061);
and U9060 (N_9060,N_7566,N_7693);
nor U9061 (N_9061,N_6357,N_7076);
or U9062 (N_9062,N_7430,N_6599);
or U9063 (N_9063,N_6184,N_6165);
nor U9064 (N_9064,N_6295,N_6016);
and U9065 (N_9065,N_7276,N_7360);
or U9066 (N_9066,N_6594,N_7180);
nor U9067 (N_9067,N_7181,N_6335);
nand U9068 (N_9068,N_6387,N_6357);
xor U9069 (N_9069,N_7914,N_6767);
and U9070 (N_9070,N_7549,N_6880);
and U9071 (N_9071,N_6917,N_7530);
and U9072 (N_9072,N_7263,N_6687);
and U9073 (N_9073,N_6190,N_7461);
nand U9074 (N_9074,N_7336,N_7242);
and U9075 (N_9075,N_6979,N_6227);
xor U9076 (N_9076,N_7312,N_7470);
nand U9077 (N_9077,N_6216,N_7927);
xor U9078 (N_9078,N_7718,N_7963);
and U9079 (N_9079,N_6750,N_6776);
and U9080 (N_9080,N_7677,N_6050);
xnor U9081 (N_9081,N_6643,N_6896);
or U9082 (N_9082,N_7056,N_6894);
and U9083 (N_9083,N_6692,N_7846);
xor U9084 (N_9084,N_6035,N_7843);
xnor U9085 (N_9085,N_7332,N_6421);
or U9086 (N_9086,N_7764,N_7771);
and U9087 (N_9087,N_7025,N_7161);
or U9088 (N_9088,N_6819,N_6297);
nand U9089 (N_9089,N_6531,N_7441);
or U9090 (N_9090,N_7688,N_6127);
nand U9091 (N_9091,N_6032,N_6228);
or U9092 (N_9092,N_7716,N_6606);
nand U9093 (N_9093,N_7412,N_6278);
nand U9094 (N_9094,N_7639,N_6255);
xor U9095 (N_9095,N_7616,N_6184);
nand U9096 (N_9096,N_6033,N_7663);
nor U9097 (N_9097,N_7025,N_6313);
nor U9098 (N_9098,N_7720,N_6129);
xnor U9099 (N_9099,N_6664,N_7867);
xnor U9100 (N_9100,N_7962,N_7558);
or U9101 (N_9101,N_7234,N_7777);
nor U9102 (N_9102,N_7474,N_7825);
or U9103 (N_9103,N_7291,N_6685);
xor U9104 (N_9104,N_7765,N_6220);
nor U9105 (N_9105,N_7672,N_6414);
and U9106 (N_9106,N_7168,N_7972);
and U9107 (N_9107,N_6059,N_6080);
or U9108 (N_9108,N_7806,N_7602);
or U9109 (N_9109,N_6816,N_6744);
nor U9110 (N_9110,N_7981,N_6287);
nor U9111 (N_9111,N_6179,N_7038);
nand U9112 (N_9112,N_7324,N_7654);
nand U9113 (N_9113,N_6359,N_6631);
nand U9114 (N_9114,N_7994,N_6649);
or U9115 (N_9115,N_7551,N_7071);
and U9116 (N_9116,N_6749,N_6720);
nor U9117 (N_9117,N_7584,N_7296);
or U9118 (N_9118,N_7337,N_6885);
nand U9119 (N_9119,N_6823,N_6168);
xor U9120 (N_9120,N_6323,N_7842);
nand U9121 (N_9121,N_6044,N_7891);
nand U9122 (N_9122,N_6788,N_7528);
and U9123 (N_9123,N_6159,N_7475);
or U9124 (N_9124,N_6200,N_7450);
or U9125 (N_9125,N_7678,N_6648);
or U9126 (N_9126,N_6966,N_7130);
nand U9127 (N_9127,N_7644,N_7721);
nor U9128 (N_9128,N_7432,N_6096);
and U9129 (N_9129,N_7884,N_7113);
xnor U9130 (N_9130,N_7542,N_7075);
nand U9131 (N_9131,N_6598,N_6578);
and U9132 (N_9132,N_7867,N_7740);
nor U9133 (N_9133,N_7446,N_7367);
xor U9134 (N_9134,N_6051,N_6033);
nand U9135 (N_9135,N_6197,N_7475);
and U9136 (N_9136,N_7493,N_6642);
and U9137 (N_9137,N_6588,N_6417);
and U9138 (N_9138,N_6161,N_6706);
nor U9139 (N_9139,N_6900,N_6817);
or U9140 (N_9140,N_6379,N_6229);
nand U9141 (N_9141,N_6073,N_6933);
nand U9142 (N_9142,N_6179,N_6671);
nor U9143 (N_9143,N_7275,N_6208);
or U9144 (N_9144,N_7963,N_6194);
or U9145 (N_9145,N_6121,N_6624);
and U9146 (N_9146,N_7093,N_6697);
nor U9147 (N_9147,N_6462,N_6152);
xnor U9148 (N_9148,N_6760,N_6338);
xor U9149 (N_9149,N_6194,N_7738);
or U9150 (N_9150,N_6698,N_6588);
nor U9151 (N_9151,N_6287,N_7550);
and U9152 (N_9152,N_7521,N_6199);
or U9153 (N_9153,N_7390,N_6148);
nor U9154 (N_9154,N_6374,N_7405);
and U9155 (N_9155,N_7640,N_6497);
nor U9156 (N_9156,N_6341,N_6972);
or U9157 (N_9157,N_7064,N_6283);
nor U9158 (N_9158,N_6601,N_6409);
nor U9159 (N_9159,N_7494,N_7700);
and U9160 (N_9160,N_6427,N_7280);
xnor U9161 (N_9161,N_7427,N_7007);
nor U9162 (N_9162,N_7029,N_6469);
nand U9163 (N_9163,N_7639,N_7516);
or U9164 (N_9164,N_7664,N_6510);
nand U9165 (N_9165,N_6953,N_6431);
nor U9166 (N_9166,N_6155,N_7167);
xnor U9167 (N_9167,N_6235,N_7794);
and U9168 (N_9168,N_7926,N_6030);
xor U9169 (N_9169,N_6485,N_7882);
nand U9170 (N_9170,N_6409,N_6139);
or U9171 (N_9171,N_7447,N_7660);
nor U9172 (N_9172,N_6403,N_7712);
and U9173 (N_9173,N_7820,N_6273);
or U9174 (N_9174,N_6768,N_6710);
nor U9175 (N_9175,N_7916,N_7531);
nor U9176 (N_9176,N_7749,N_6557);
nor U9177 (N_9177,N_6799,N_6824);
xnor U9178 (N_9178,N_6295,N_6670);
nor U9179 (N_9179,N_6718,N_6772);
nand U9180 (N_9180,N_7408,N_6816);
xnor U9181 (N_9181,N_6613,N_7537);
nand U9182 (N_9182,N_6236,N_6250);
and U9183 (N_9183,N_6080,N_7050);
nor U9184 (N_9184,N_7344,N_7887);
or U9185 (N_9185,N_6152,N_6070);
or U9186 (N_9186,N_6217,N_7039);
and U9187 (N_9187,N_6804,N_6204);
and U9188 (N_9188,N_7211,N_7636);
nand U9189 (N_9189,N_7566,N_7694);
or U9190 (N_9190,N_7624,N_7496);
or U9191 (N_9191,N_6095,N_6292);
nor U9192 (N_9192,N_7244,N_7828);
and U9193 (N_9193,N_6592,N_7440);
xnor U9194 (N_9194,N_6842,N_6837);
nor U9195 (N_9195,N_7929,N_7291);
xnor U9196 (N_9196,N_6064,N_7569);
nor U9197 (N_9197,N_7747,N_6293);
nor U9198 (N_9198,N_7930,N_6095);
and U9199 (N_9199,N_6055,N_6352);
xnor U9200 (N_9200,N_6989,N_7819);
and U9201 (N_9201,N_7687,N_7222);
and U9202 (N_9202,N_7005,N_7576);
or U9203 (N_9203,N_6887,N_7303);
xnor U9204 (N_9204,N_6351,N_7913);
or U9205 (N_9205,N_6194,N_7951);
or U9206 (N_9206,N_7720,N_6222);
nor U9207 (N_9207,N_7424,N_7369);
nand U9208 (N_9208,N_6724,N_7822);
xor U9209 (N_9209,N_6641,N_6190);
and U9210 (N_9210,N_6062,N_7851);
nor U9211 (N_9211,N_7732,N_6694);
and U9212 (N_9212,N_7146,N_6431);
and U9213 (N_9213,N_6437,N_7918);
nor U9214 (N_9214,N_6146,N_6586);
nand U9215 (N_9215,N_6499,N_6875);
or U9216 (N_9216,N_6190,N_6239);
and U9217 (N_9217,N_6554,N_6313);
nand U9218 (N_9218,N_7058,N_7570);
xnor U9219 (N_9219,N_6563,N_7461);
nor U9220 (N_9220,N_6042,N_6269);
xor U9221 (N_9221,N_6316,N_7803);
and U9222 (N_9222,N_7883,N_7543);
nor U9223 (N_9223,N_7775,N_7648);
nor U9224 (N_9224,N_7353,N_7040);
nor U9225 (N_9225,N_6686,N_7250);
nor U9226 (N_9226,N_6575,N_6361);
and U9227 (N_9227,N_6440,N_6293);
or U9228 (N_9228,N_6191,N_6766);
nand U9229 (N_9229,N_7462,N_6689);
nor U9230 (N_9230,N_7461,N_7471);
nor U9231 (N_9231,N_6704,N_7872);
nand U9232 (N_9232,N_7169,N_6609);
nor U9233 (N_9233,N_6773,N_6151);
nor U9234 (N_9234,N_6321,N_7971);
and U9235 (N_9235,N_6369,N_7698);
or U9236 (N_9236,N_6948,N_7174);
xnor U9237 (N_9237,N_7795,N_6683);
nor U9238 (N_9238,N_7331,N_6606);
and U9239 (N_9239,N_7921,N_6658);
xnor U9240 (N_9240,N_7030,N_7689);
xor U9241 (N_9241,N_7442,N_6404);
or U9242 (N_9242,N_6023,N_7061);
and U9243 (N_9243,N_7317,N_6846);
and U9244 (N_9244,N_7903,N_7483);
and U9245 (N_9245,N_6619,N_6809);
nand U9246 (N_9246,N_6291,N_6054);
and U9247 (N_9247,N_7188,N_7725);
or U9248 (N_9248,N_7727,N_6905);
nand U9249 (N_9249,N_7974,N_6450);
or U9250 (N_9250,N_6593,N_7302);
and U9251 (N_9251,N_6652,N_7506);
or U9252 (N_9252,N_6188,N_7950);
and U9253 (N_9253,N_6427,N_7993);
nand U9254 (N_9254,N_6781,N_6997);
xor U9255 (N_9255,N_7722,N_7845);
nor U9256 (N_9256,N_6691,N_7615);
nor U9257 (N_9257,N_7189,N_7605);
or U9258 (N_9258,N_7401,N_7426);
and U9259 (N_9259,N_7517,N_7866);
nand U9260 (N_9260,N_7025,N_6733);
xor U9261 (N_9261,N_7691,N_6980);
nor U9262 (N_9262,N_6299,N_6412);
nor U9263 (N_9263,N_6104,N_6283);
nand U9264 (N_9264,N_7021,N_7126);
and U9265 (N_9265,N_7224,N_6111);
nand U9266 (N_9266,N_6016,N_6893);
nor U9267 (N_9267,N_7092,N_7608);
nand U9268 (N_9268,N_7065,N_7972);
and U9269 (N_9269,N_7193,N_7520);
nor U9270 (N_9270,N_6438,N_6942);
nor U9271 (N_9271,N_6138,N_6783);
and U9272 (N_9272,N_6430,N_6956);
or U9273 (N_9273,N_7405,N_7600);
nand U9274 (N_9274,N_7431,N_6774);
nor U9275 (N_9275,N_6440,N_6671);
and U9276 (N_9276,N_7591,N_7700);
and U9277 (N_9277,N_6627,N_6696);
or U9278 (N_9278,N_7289,N_6595);
nand U9279 (N_9279,N_7656,N_7920);
nand U9280 (N_9280,N_7355,N_6597);
xor U9281 (N_9281,N_6792,N_6400);
nor U9282 (N_9282,N_6993,N_7289);
or U9283 (N_9283,N_6540,N_7016);
nand U9284 (N_9284,N_6496,N_6492);
nand U9285 (N_9285,N_6873,N_7956);
and U9286 (N_9286,N_6619,N_6707);
nand U9287 (N_9287,N_7656,N_7383);
xor U9288 (N_9288,N_7403,N_7144);
or U9289 (N_9289,N_7660,N_6157);
xnor U9290 (N_9290,N_6348,N_7989);
and U9291 (N_9291,N_6808,N_7368);
or U9292 (N_9292,N_7215,N_6050);
and U9293 (N_9293,N_6154,N_6847);
nand U9294 (N_9294,N_6278,N_7532);
nor U9295 (N_9295,N_6403,N_7655);
xnor U9296 (N_9296,N_7640,N_7157);
nand U9297 (N_9297,N_7239,N_7703);
or U9298 (N_9298,N_7419,N_6319);
xnor U9299 (N_9299,N_7003,N_6156);
nand U9300 (N_9300,N_7764,N_6727);
xor U9301 (N_9301,N_7399,N_7689);
xnor U9302 (N_9302,N_6933,N_6186);
and U9303 (N_9303,N_6923,N_7354);
or U9304 (N_9304,N_6109,N_6293);
or U9305 (N_9305,N_7322,N_7423);
nor U9306 (N_9306,N_6662,N_7900);
xor U9307 (N_9307,N_7323,N_7386);
nand U9308 (N_9308,N_7999,N_7462);
or U9309 (N_9309,N_7023,N_6207);
or U9310 (N_9310,N_6513,N_6603);
nor U9311 (N_9311,N_7908,N_7534);
and U9312 (N_9312,N_6143,N_6670);
nor U9313 (N_9313,N_6861,N_6823);
or U9314 (N_9314,N_7102,N_6510);
nand U9315 (N_9315,N_6151,N_7563);
xor U9316 (N_9316,N_7065,N_6603);
xor U9317 (N_9317,N_6308,N_6720);
nand U9318 (N_9318,N_7798,N_7018);
nor U9319 (N_9319,N_7360,N_6051);
nor U9320 (N_9320,N_6831,N_7475);
nor U9321 (N_9321,N_6387,N_6167);
or U9322 (N_9322,N_6086,N_6656);
and U9323 (N_9323,N_7605,N_6690);
nor U9324 (N_9324,N_7006,N_7696);
or U9325 (N_9325,N_7033,N_7552);
and U9326 (N_9326,N_6246,N_7042);
and U9327 (N_9327,N_6723,N_6557);
xnor U9328 (N_9328,N_7423,N_6733);
and U9329 (N_9329,N_6000,N_7736);
nor U9330 (N_9330,N_7750,N_7456);
or U9331 (N_9331,N_7842,N_6876);
xor U9332 (N_9332,N_6949,N_7174);
nor U9333 (N_9333,N_7979,N_7226);
nor U9334 (N_9334,N_7209,N_7791);
xor U9335 (N_9335,N_6045,N_6837);
xor U9336 (N_9336,N_6864,N_6943);
xor U9337 (N_9337,N_6554,N_6065);
or U9338 (N_9338,N_6108,N_7996);
nor U9339 (N_9339,N_6467,N_7129);
xnor U9340 (N_9340,N_7094,N_7670);
and U9341 (N_9341,N_7796,N_7686);
or U9342 (N_9342,N_6192,N_6150);
nor U9343 (N_9343,N_6308,N_6233);
nand U9344 (N_9344,N_7815,N_7451);
xnor U9345 (N_9345,N_7974,N_6010);
nor U9346 (N_9346,N_6890,N_7571);
and U9347 (N_9347,N_6715,N_6945);
and U9348 (N_9348,N_7653,N_7950);
nand U9349 (N_9349,N_6844,N_6913);
nor U9350 (N_9350,N_7045,N_6861);
nor U9351 (N_9351,N_6016,N_6933);
and U9352 (N_9352,N_7721,N_7192);
nand U9353 (N_9353,N_6994,N_7692);
or U9354 (N_9354,N_6016,N_6101);
nor U9355 (N_9355,N_6469,N_7042);
and U9356 (N_9356,N_6535,N_7406);
or U9357 (N_9357,N_7586,N_7188);
xor U9358 (N_9358,N_6128,N_7747);
xor U9359 (N_9359,N_7486,N_6995);
and U9360 (N_9360,N_7551,N_7520);
and U9361 (N_9361,N_7822,N_6834);
and U9362 (N_9362,N_6794,N_7785);
nor U9363 (N_9363,N_7460,N_7663);
and U9364 (N_9364,N_7322,N_6740);
nand U9365 (N_9365,N_7951,N_6066);
xor U9366 (N_9366,N_6186,N_7101);
or U9367 (N_9367,N_6753,N_6702);
nand U9368 (N_9368,N_7690,N_7315);
and U9369 (N_9369,N_6733,N_6218);
nor U9370 (N_9370,N_7532,N_6422);
nand U9371 (N_9371,N_7013,N_6944);
and U9372 (N_9372,N_6272,N_6512);
or U9373 (N_9373,N_6238,N_7108);
nor U9374 (N_9374,N_6555,N_7743);
and U9375 (N_9375,N_6745,N_7091);
and U9376 (N_9376,N_7005,N_6283);
or U9377 (N_9377,N_6850,N_7448);
xor U9378 (N_9378,N_7629,N_6845);
and U9379 (N_9379,N_7295,N_7460);
and U9380 (N_9380,N_6704,N_6428);
nor U9381 (N_9381,N_7147,N_6278);
nor U9382 (N_9382,N_6062,N_6589);
nand U9383 (N_9383,N_7377,N_6864);
or U9384 (N_9384,N_7872,N_7145);
or U9385 (N_9385,N_6960,N_6280);
or U9386 (N_9386,N_6166,N_7043);
and U9387 (N_9387,N_6937,N_6468);
nor U9388 (N_9388,N_6477,N_6273);
or U9389 (N_9389,N_6778,N_7410);
nand U9390 (N_9390,N_7318,N_6809);
nor U9391 (N_9391,N_6578,N_6892);
and U9392 (N_9392,N_6479,N_6871);
xnor U9393 (N_9393,N_7405,N_6223);
or U9394 (N_9394,N_7548,N_7168);
nor U9395 (N_9395,N_7623,N_6265);
nor U9396 (N_9396,N_6550,N_7954);
xor U9397 (N_9397,N_7443,N_6488);
nor U9398 (N_9398,N_6603,N_7449);
or U9399 (N_9399,N_6807,N_7539);
nor U9400 (N_9400,N_7789,N_6018);
xor U9401 (N_9401,N_7367,N_7161);
and U9402 (N_9402,N_7101,N_7359);
xnor U9403 (N_9403,N_7098,N_6219);
xor U9404 (N_9404,N_6309,N_7988);
nor U9405 (N_9405,N_6356,N_6676);
or U9406 (N_9406,N_6302,N_7301);
nor U9407 (N_9407,N_7596,N_7886);
and U9408 (N_9408,N_6394,N_7857);
nor U9409 (N_9409,N_6678,N_7173);
nor U9410 (N_9410,N_7512,N_7921);
or U9411 (N_9411,N_6325,N_7496);
xor U9412 (N_9412,N_6424,N_7012);
nor U9413 (N_9413,N_6250,N_6933);
nand U9414 (N_9414,N_7125,N_7941);
or U9415 (N_9415,N_6888,N_7877);
xor U9416 (N_9416,N_7874,N_7270);
and U9417 (N_9417,N_6628,N_7995);
nor U9418 (N_9418,N_6944,N_7830);
and U9419 (N_9419,N_7870,N_7707);
xor U9420 (N_9420,N_6911,N_6746);
xnor U9421 (N_9421,N_7702,N_6193);
and U9422 (N_9422,N_6936,N_6807);
nor U9423 (N_9423,N_6909,N_7824);
xor U9424 (N_9424,N_7786,N_7805);
nor U9425 (N_9425,N_7792,N_6874);
xor U9426 (N_9426,N_6335,N_6624);
and U9427 (N_9427,N_7943,N_6488);
or U9428 (N_9428,N_7345,N_6560);
or U9429 (N_9429,N_6747,N_7886);
nor U9430 (N_9430,N_6573,N_6394);
nor U9431 (N_9431,N_7090,N_7388);
xnor U9432 (N_9432,N_6480,N_7537);
nor U9433 (N_9433,N_6561,N_7911);
and U9434 (N_9434,N_6938,N_7521);
nand U9435 (N_9435,N_7521,N_6584);
or U9436 (N_9436,N_6321,N_7118);
nor U9437 (N_9437,N_7330,N_6364);
xor U9438 (N_9438,N_7892,N_7815);
nor U9439 (N_9439,N_7482,N_7085);
and U9440 (N_9440,N_6318,N_7956);
xor U9441 (N_9441,N_6926,N_7545);
and U9442 (N_9442,N_7157,N_6728);
xnor U9443 (N_9443,N_7656,N_6393);
and U9444 (N_9444,N_7362,N_6893);
nand U9445 (N_9445,N_6754,N_7994);
and U9446 (N_9446,N_6167,N_6925);
and U9447 (N_9447,N_7143,N_6805);
nand U9448 (N_9448,N_6477,N_7444);
nand U9449 (N_9449,N_7638,N_6004);
nor U9450 (N_9450,N_7457,N_6415);
nor U9451 (N_9451,N_6976,N_7009);
nand U9452 (N_9452,N_6099,N_6475);
nor U9453 (N_9453,N_6032,N_6659);
nand U9454 (N_9454,N_7342,N_7398);
nor U9455 (N_9455,N_7952,N_6243);
nor U9456 (N_9456,N_7691,N_6297);
and U9457 (N_9457,N_6218,N_6781);
nor U9458 (N_9458,N_6032,N_6175);
and U9459 (N_9459,N_6362,N_7776);
and U9460 (N_9460,N_7816,N_6619);
or U9461 (N_9461,N_7956,N_6990);
nand U9462 (N_9462,N_6096,N_6448);
nor U9463 (N_9463,N_6095,N_7594);
nor U9464 (N_9464,N_7673,N_7616);
xor U9465 (N_9465,N_6418,N_7346);
nand U9466 (N_9466,N_7470,N_7092);
and U9467 (N_9467,N_6960,N_6908);
and U9468 (N_9468,N_6325,N_7474);
or U9469 (N_9469,N_6123,N_6891);
and U9470 (N_9470,N_7800,N_7735);
xnor U9471 (N_9471,N_7143,N_6774);
or U9472 (N_9472,N_7579,N_7067);
nand U9473 (N_9473,N_6147,N_7859);
xor U9474 (N_9474,N_7859,N_6438);
xor U9475 (N_9475,N_7924,N_7137);
xor U9476 (N_9476,N_7934,N_6380);
and U9477 (N_9477,N_7821,N_7993);
nor U9478 (N_9478,N_7538,N_6423);
and U9479 (N_9479,N_7211,N_7489);
and U9480 (N_9480,N_6633,N_6921);
or U9481 (N_9481,N_6434,N_6730);
or U9482 (N_9482,N_7952,N_6395);
or U9483 (N_9483,N_6056,N_6166);
or U9484 (N_9484,N_6659,N_6460);
or U9485 (N_9485,N_6696,N_6044);
and U9486 (N_9486,N_7761,N_6069);
xor U9487 (N_9487,N_7727,N_7838);
xnor U9488 (N_9488,N_6954,N_6677);
and U9489 (N_9489,N_7191,N_6167);
nand U9490 (N_9490,N_7676,N_6746);
or U9491 (N_9491,N_7346,N_6431);
nand U9492 (N_9492,N_6449,N_6901);
xnor U9493 (N_9493,N_7779,N_6981);
nor U9494 (N_9494,N_6389,N_6947);
and U9495 (N_9495,N_7356,N_6110);
nand U9496 (N_9496,N_6603,N_6009);
and U9497 (N_9497,N_7663,N_6864);
or U9498 (N_9498,N_6922,N_7890);
or U9499 (N_9499,N_6834,N_6056);
xor U9500 (N_9500,N_6136,N_6040);
or U9501 (N_9501,N_6102,N_6970);
nand U9502 (N_9502,N_6937,N_6447);
and U9503 (N_9503,N_7539,N_7318);
and U9504 (N_9504,N_7283,N_6960);
and U9505 (N_9505,N_6340,N_6227);
nand U9506 (N_9506,N_6498,N_7274);
xor U9507 (N_9507,N_6121,N_6435);
nand U9508 (N_9508,N_6814,N_7946);
xnor U9509 (N_9509,N_6911,N_6796);
or U9510 (N_9510,N_7155,N_7256);
or U9511 (N_9511,N_6094,N_7949);
nor U9512 (N_9512,N_6092,N_6171);
xor U9513 (N_9513,N_6064,N_6781);
and U9514 (N_9514,N_7675,N_7172);
xnor U9515 (N_9515,N_7985,N_6105);
and U9516 (N_9516,N_6411,N_6884);
xnor U9517 (N_9517,N_7163,N_6829);
or U9518 (N_9518,N_7542,N_6687);
xnor U9519 (N_9519,N_6560,N_7159);
nand U9520 (N_9520,N_6140,N_6560);
nand U9521 (N_9521,N_6026,N_7074);
and U9522 (N_9522,N_6777,N_7983);
nor U9523 (N_9523,N_6045,N_6752);
or U9524 (N_9524,N_7721,N_7478);
and U9525 (N_9525,N_7060,N_7446);
nand U9526 (N_9526,N_7720,N_6221);
nor U9527 (N_9527,N_7385,N_7791);
and U9528 (N_9528,N_6742,N_7611);
and U9529 (N_9529,N_7618,N_7931);
or U9530 (N_9530,N_7222,N_6477);
nand U9531 (N_9531,N_6922,N_7924);
or U9532 (N_9532,N_6418,N_6954);
xor U9533 (N_9533,N_6652,N_7019);
xnor U9534 (N_9534,N_7743,N_7961);
nor U9535 (N_9535,N_6269,N_6319);
and U9536 (N_9536,N_7285,N_6230);
xor U9537 (N_9537,N_6161,N_6819);
nor U9538 (N_9538,N_7801,N_6920);
xnor U9539 (N_9539,N_6149,N_7609);
xnor U9540 (N_9540,N_6333,N_7504);
and U9541 (N_9541,N_7376,N_6004);
nor U9542 (N_9542,N_7849,N_7060);
nand U9543 (N_9543,N_6387,N_7217);
or U9544 (N_9544,N_6053,N_7865);
or U9545 (N_9545,N_7333,N_7225);
nor U9546 (N_9546,N_6124,N_7705);
xnor U9547 (N_9547,N_7475,N_6393);
xor U9548 (N_9548,N_7003,N_6522);
or U9549 (N_9549,N_7845,N_7231);
and U9550 (N_9550,N_7528,N_6994);
and U9551 (N_9551,N_7295,N_7794);
nand U9552 (N_9552,N_6773,N_7993);
nand U9553 (N_9553,N_7584,N_6265);
nor U9554 (N_9554,N_7205,N_6063);
or U9555 (N_9555,N_6388,N_7330);
nand U9556 (N_9556,N_7676,N_7705);
nand U9557 (N_9557,N_6225,N_7860);
xnor U9558 (N_9558,N_6126,N_6898);
nor U9559 (N_9559,N_6732,N_7730);
nor U9560 (N_9560,N_6208,N_6677);
nand U9561 (N_9561,N_6919,N_7978);
xnor U9562 (N_9562,N_7105,N_6643);
xnor U9563 (N_9563,N_6701,N_6429);
and U9564 (N_9564,N_6238,N_6110);
nand U9565 (N_9565,N_7319,N_7776);
nor U9566 (N_9566,N_6178,N_6867);
and U9567 (N_9567,N_7969,N_7190);
nand U9568 (N_9568,N_7413,N_7785);
xnor U9569 (N_9569,N_7831,N_7119);
nand U9570 (N_9570,N_6865,N_6068);
and U9571 (N_9571,N_6688,N_6814);
nor U9572 (N_9572,N_6378,N_6661);
nand U9573 (N_9573,N_7937,N_7199);
nand U9574 (N_9574,N_6494,N_7200);
and U9575 (N_9575,N_6246,N_6549);
or U9576 (N_9576,N_7562,N_7732);
or U9577 (N_9577,N_7494,N_6870);
xor U9578 (N_9578,N_6724,N_7540);
or U9579 (N_9579,N_7519,N_6546);
or U9580 (N_9580,N_7933,N_6445);
nand U9581 (N_9581,N_7161,N_7958);
xnor U9582 (N_9582,N_7821,N_7939);
nand U9583 (N_9583,N_7093,N_6766);
or U9584 (N_9584,N_6776,N_7131);
nand U9585 (N_9585,N_7663,N_6496);
xor U9586 (N_9586,N_7148,N_7417);
nor U9587 (N_9587,N_7654,N_6840);
nand U9588 (N_9588,N_6782,N_7014);
and U9589 (N_9589,N_6957,N_7847);
or U9590 (N_9590,N_7462,N_6939);
nor U9591 (N_9591,N_6871,N_6848);
and U9592 (N_9592,N_6724,N_6270);
or U9593 (N_9593,N_6021,N_6892);
xor U9594 (N_9594,N_6126,N_6625);
xnor U9595 (N_9595,N_7888,N_6761);
nor U9596 (N_9596,N_7009,N_7429);
and U9597 (N_9597,N_6580,N_7871);
nand U9598 (N_9598,N_7025,N_7181);
nor U9599 (N_9599,N_6426,N_7681);
nand U9600 (N_9600,N_7344,N_6839);
nand U9601 (N_9601,N_6812,N_6215);
nand U9602 (N_9602,N_6713,N_6524);
nor U9603 (N_9603,N_6697,N_7262);
or U9604 (N_9604,N_6144,N_6758);
and U9605 (N_9605,N_6716,N_7148);
nor U9606 (N_9606,N_7148,N_7903);
nand U9607 (N_9607,N_7207,N_7361);
nor U9608 (N_9608,N_7493,N_6993);
or U9609 (N_9609,N_7728,N_6599);
and U9610 (N_9610,N_7985,N_7815);
or U9611 (N_9611,N_7359,N_7013);
nor U9612 (N_9612,N_7731,N_7944);
and U9613 (N_9613,N_6151,N_7535);
or U9614 (N_9614,N_7729,N_7061);
and U9615 (N_9615,N_6165,N_6577);
nand U9616 (N_9616,N_6066,N_6344);
nand U9617 (N_9617,N_6384,N_7043);
or U9618 (N_9618,N_6142,N_7440);
or U9619 (N_9619,N_6818,N_6243);
nand U9620 (N_9620,N_7086,N_7737);
nand U9621 (N_9621,N_7384,N_6415);
xnor U9622 (N_9622,N_6947,N_7747);
or U9623 (N_9623,N_7426,N_7666);
and U9624 (N_9624,N_7592,N_6070);
nor U9625 (N_9625,N_6313,N_6672);
nand U9626 (N_9626,N_7672,N_7099);
or U9627 (N_9627,N_6202,N_6287);
nand U9628 (N_9628,N_7019,N_7260);
nand U9629 (N_9629,N_6583,N_7076);
nand U9630 (N_9630,N_7382,N_7028);
or U9631 (N_9631,N_7285,N_7866);
nand U9632 (N_9632,N_7860,N_6043);
nand U9633 (N_9633,N_7233,N_7750);
xnor U9634 (N_9634,N_6209,N_6782);
nor U9635 (N_9635,N_6902,N_7308);
xor U9636 (N_9636,N_7348,N_6166);
nand U9637 (N_9637,N_7299,N_7770);
nor U9638 (N_9638,N_7895,N_7400);
or U9639 (N_9639,N_7617,N_7755);
or U9640 (N_9640,N_7681,N_7972);
and U9641 (N_9641,N_7755,N_7356);
and U9642 (N_9642,N_6584,N_7505);
or U9643 (N_9643,N_6368,N_7157);
xnor U9644 (N_9644,N_7238,N_7486);
or U9645 (N_9645,N_7352,N_6650);
nor U9646 (N_9646,N_6984,N_7251);
xor U9647 (N_9647,N_7237,N_7397);
or U9648 (N_9648,N_7008,N_7366);
or U9649 (N_9649,N_6541,N_6754);
xor U9650 (N_9650,N_6454,N_7265);
or U9651 (N_9651,N_6230,N_7712);
and U9652 (N_9652,N_6815,N_6564);
nor U9653 (N_9653,N_7793,N_7851);
or U9654 (N_9654,N_7098,N_6702);
xor U9655 (N_9655,N_7152,N_7269);
nor U9656 (N_9656,N_6229,N_7059);
or U9657 (N_9657,N_7623,N_6714);
xnor U9658 (N_9658,N_7182,N_7919);
or U9659 (N_9659,N_6232,N_7171);
nand U9660 (N_9660,N_7689,N_6535);
nand U9661 (N_9661,N_7227,N_7632);
nand U9662 (N_9662,N_6701,N_7470);
or U9663 (N_9663,N_7269,N_6496);
nand U9664 (N_9664,N_6216,N_6105);
nand U9665 (N_9665,N_6956,N_7011);
nor U9666 (N_9666,N_7687,N_6999);
nand U9667 (N_9667,N_7197,N_7323);
and U9668 (N_9668,N_6384,N_7503);
and U9669 (N_9669,N_6905,N_7070);
or U9670 (N_9670,N_6861,N_6022);
nand U9671 (N_9671,N_7378,N_6866);
nor U9672 (N_9672,N_7551,N_7439);
nand U9673 (N_9673,N_7682,N_6143);
xor U9674 (N_9674,N_7049,N_7851);
nor U9675 (N_9675,N_7234,N_6152);
or U9676 (N_9676,N_7650,N_7383);
xor U9677 (N_9677,N_7214,N_6135);
nor U9678 (N_9678,N_6784,N_7867);
and U9679 (N_9679,N_6155,N_6408);
nor U9680 (N_9680,N_6429,N_7819);
and U9681 (N_9681,N_6217,N_7360);
and U9682 (N_9682,N_6137,N_6698);
nor U9683 (N_9683,N_7516,N_6831);
nand U9684 (N_9684,N_7032,N_6488);
nand U9685 (N_9685,N_7704,N_6823);
nor U9686 (N_9686,N_7612,N_7689);
nand U9687 (N_9687,N_7032,N_6757);
or U9688 (N_9688,N_6321,N_7401);
nor U9689 (N_9689,N_7854,N_7307);
nor U9690 (N_9690,N_6715,N_7259);
xnor U9691 (N_9691,N_7983,N_6872);
or U9692 (N_9692,N_6531,N_6812);
xor U9693 (N_9693,N_7062,N_6528);
and U9694 (N_9694,N_6058,N_6287);
nor U9695 (N_9695,N_6318,N_7147);
xor U9696 (N_9696,N_7149,N_7682);
nand U9697 (N_9697,N_7662,N_7483);
or U9698 (N_9698,N_7192,N_6575);
xnor U9699 (N_9699,N_7350,N_6629);
nand U9700 (N_9700,N_6124,N_7886);
or U9701 (N_9701,N_7855,N_6030);
xnor U9702 (N_9702,N_7327,N_7278);
or U9703 (N_9703,N_7204,N_7165);
nor U9704 (N_9704,N_6752,N_6924);
xor U9705 (N_9705,N_6596,N_7559);
and U9706 (N_9706,N_7161,N_6825);
nor U9707 (N_9707,N_6585,N_7756);
nand U9708 (N_9708,N_7735,N_7657);
nor U9709 (N_9709,N_7626,N_6279);
or U9710 (N_9710,N_6589,N_7758);
nor U9711 (N_9711,N_6011,N_6930);
or U9712 (N_9712,N_6345,N_7174);
and U9713 (N_9713,N_7179,N_7957);
nor U9714 (N_9714,N_7208,N_6813);
nand U9715 (N_9715,N_6016,N_6119);
nor U9716 (N_9716,N_6842,N_6239);
xor U9717 (N_9717,N_6229,N_6582);
nor U9718 (N_9718,N_7812,N_7802);
nor U9719 (N_9719,N_6959,N_7692);
nand U9720 (N_9720,N_7929,N_6238);
nand U9721 (N_9721,N_6512,N_6404);
nand U9722 (N_9722,N_6535,N_7465);
or U9723 (N_9723,N_6479,N_7973);
nor U9724 (N_9724,N_7201,N_7103);
nor U9725 (N_9725,N_6006,N_7767);
xnor U9726 (N_9726,N_7224,N_7661);
nand U9727 (N_9727,N_6252,N_7472);
xnor U9728 (N_9728,N_7437,N_6754);
or U9729 (N_9729,N_7978,N_6683);
and U9730 (N_9730,N_6128,N_7729);
or U9731 (N_9731,N_6987,N_7006);
or U9732 (N_9732,N_6929,N_6164);
or U9733 (N_9733,N_7893,N_7624);
or U9734 (N_9734,N_7321,N_7525);
and U9735 (N_9735,N_7295,N_6820);
xor U9736 (N_9736,N_6112,N_6589);
nand U9737 (N_9737,N_7591,N_6876);
xnor U9738 (N_9738,N_6629,N_7670);
nand U9739 (N_9739,N_7664,N_6182);
nor U9740 (N_9740,N_7757,N_6523);
or U9741 (N_9741,N_7591,N_7518);
nand U9742 (N_9742,N_6397,N_7693);
nor U9743 (N_9743,N_6884,N_7956);
nand U9744 (N_9744,N_6547,N_7802);
and U9745 (N_9745,N_6623,N_7051);
and U9746 (N_9746,N_6983,N_6056);
and U9747 (N_9747,N_6346,N_6302);
xnor U9748 (N_9748,N_6246,N_6726);
xor U9749 (N_9749,N_7653,N_6244);
and U9750 (N_9750,N_6410,N_6916);
nor U9751 (N_9751,N_6690,N_6149);
nand U9752 (N_9752,N_6743,N_6491);
and U9753 (N_9753,N_7337,N_6842);
nor U9754 (N_9754,N_7223,N_7196);
and U9755 (N_9755,N_7451,N_6754);
and U9756 (N_9756,N_6949,N_7493);
nor U9757 (N_9757,N_6737,N_7381);
nor U9758 (N_9758,N_7625,N_7019);
xor U9759 (N_9759,N_7432,N_6277);
or U9760 (N_9760,N_7090,N_7841);
xor U9761 (N_9761,N_7357,N_6712);
or U9762 (N_9762,N_6205,N_6288);
nor U9763 (N_9763,N_6185,N_6021);
xor U9764 (N_9764,N_7474,N_7450);
nor U9765 (N_9765,N_6211,N_7381);
xor U9766 (N_9766,N_7955,N_7958);
or U9767 (N_9767,N_6806,N_7808);
nand U9768 (N_9768,N_6993,N_7726);
xor U9769 (N_9769,N_7612,N_7577);
and U9770 (N_9770,N_7940,N_7026);
or U9771 (N_9771,N_6038,N_7853);
or U9772 (N_9772,N_6160,N_7888);
nor U9773 (N_9773,N_6254,N_7745);
nand U9774 (N_9774,N_6044,N_6380);
or U9775 (N_9775,N_7033,N_7607);
nand U9776 (N_9776,N_7185,N_7419);
nor U9777 (N_9777,N_6169,N_6252);
and U9778 (N_9778,N_7854,N_6206);
xnor U9779 (N_9779,N_7778,N_6585);
nand U9780 (N_9780,N_7473,N_7542);
nor U9781 (N_9781,N_7191,N_7649);
xnor U9782 (N_9782,N_7714,N_7979);
xnor U9783 (N_9783,N_6706,N_6176);
nor U9784 (N_9784,N_6262,N_7663);
and U9785 (N_9785,N_6704,N_7814);
or U9786 (N_9786,N_7093,N_6620);
nor U9787 (N_9787,N_7851,N_6766);
and U9788 (N_9788,N_7599,N_6265);
and U9789 (N_9789,N_7386,N_7548);
nand U9790 (N_9790,N_6688,N_6857);
and U9791 (N_9791,N_6332,N_7828);
or U9792 (N_9792,N_7064,N_7858);
xor U9793 (N_9793,N_6791,N_7084);
nand U9794 (N_9794,N_7768,N_6496);
and U9795 (N_9795,N_6176,N_6062);
and U9796 (N_9796,N_7800,N_7021);
xor U9797 (N_9797,N_6936,N_6089);
or U9798 (N_9798,N_6884,N_6463);
and U9799 (N_9799,N_6871,N_7175);
nand U9800 (N_9800,N_7923,N_6601);
xor U9801 (N_9801,N_6446,N_6943);
or U9802 (N_9802,N_6366,N_6250);
xnor U9803 (N_9803,N_7436,N_7210);
nor U9804 (N_9804,N_7092,N_6144);
nor U9805 (N_9805,N_7139,N_7293);
xnor U9806 (N_9806,N_7806,N_6529);
or U9807 (N_9807,N_6895,N_6344);
xor U9808 (N_9808,N_7988,N_6742);
or U9809 (N_9809,N_6572,N_7648);
xnor U9810 (N_9810,N_7452,N_6807);
and U9811 (N_9811,N_7986,N_7493);
nor U9812 (N_9812,N_7102,N_7925);
or U9813 (N_9813,N_6650,N_6741);
xnor U9814 (N_9814,N_7908,N_6487);
nor U9815 (N_9815,N_7972,N_6094);
or U9816 (N_9816,N_7156,N_7160);
xnor U9817 (N_9817,N_7397,N_7123);
xor U9818 (N_9818,N_6546,N_6087);
and U9819 (N_9819,N_7774,N_6402);
xnor U9820 (N_9820,N_7399,N_6392);
nand U9821 (N_9821,N_7441,N_6221);
xnor U9822 (N_9822,N_6617,N_7484);
or U9823 (N_9823,N_7649,N_7871);
or U9824 (N_9824,N_6657,N_7625);
nor U9825 (N_9825,N_7612,N_6777);
and U9826 (N_9826,N_7525,N_6135);
or U9827 (N_9827,N_7828,N_7266);
and U9828 (N_9828,N_7183,N_6363);
nand U9829 (N_9829,N_6444,N_7206);
and U9830 (N_9830,N_6187,N_7839);
nand U9831 (N_9831,N_7283,N_7900);
xor U9832 (N_9832,N_7831,N_6935);
nand U9833 (N_9833,N_7323,N_6898);
nor U9834 (N_9834,N_7684,N_7473);
and U9835 (N_9835,N_7229,N_6136);
xnor U9836 (N_9836,N_7896,N_6567);
nor U9837 (N_9837,N_6026,N_6662);
or U9838 (N_9838,N_7217,N_7037);
xnor U9839 (N_9839,N_6622,N_7527);
nand U9840 (N_9840,N_7109,N_6778);
xnor U9841 (N_9841,N_6699,N_6259);
nor U9842 (N_9842,N_6679,N_6265);
nand U9843 (N_9843,N_7237,N_7544);
or U9844 (N_9844,N_7930,N_6585);
and U9845 (N_9845,N_6018,N_6089);
xor U9846 (N_9846,N_6514,N_7804);
nand U9847 (N_9847,N_6209,N_7725);
nand U9848 (N_9848,N_6907,N_7132);
and U9849 (N_9849,N_6061,N_6069);
or U9850 (N_9850,N_6509,N_7250);
nor U9851 (N_9851,N_7263,N_6174);
nor U9852 (N_9852,N_7422,N_7282);
nand U9853 (N_9853,N_6074,N_6798);
nor U9854 (N_9854,N_7434,N_7043);
or U9855 (N_9855,N_7565,N_7445);
xnor U9856 (N_9856,N_6879,N_6026);
nand U9857 (N_9857,N_7667,N_7030);
nand U9858 (N_9858,N_7369,N_6361);
nand U9859 (N_9859,N_7836,N_6570);
or U9860 (N_9860,N_6765,N_7409);
nand U9861 (N_9861,N_7827,N_6054);
and U9862 (N_9862,N_7380,N_7597);
nand U9863 (N_9863,N_6586,N_7866);
xor U9864 (N_9864,N_6298,N_7137);
and U9865 (N_9865,N_6453,N_7609);
and U9866 (N_9866,N_6802,N_6266);
nor U9867 (N_9867,N_7386,N_6680);
and U9868 (N_9868,N_7060,N_6069);
xor U9869 (N_9869,N_6825,N_6392);
xor U9870 (N_9870,N_7082,N_7097);
and U9871 (N_9871,N_6682,N_7830);
xor U9872 (N_9872,N_7241,N_7794);
nor U9873 (N_9873,N_7007,N_7665);
nand U9874 (N_9874,N_6758,N_7393);
and U9875 (N_9875,N_6362,N_6997);
nor U9876 (N_9876,N_7651,N_6823);
or U9877 (N_9877,N_6404,N_6381);
nand U9878 (N_9878,N_7097,N_6313);
and U9879 (N_9879,N_7564,N_7442);
and U9880 (N_9880,N_6577,N_6830);
nor U9881 (N_9881,N_6264,N_6928);
nor U9882 (N_9882,N_7508,N_7024);
xnor U9883 (N_9883,N_6177,N_6758);
and U9884 (N_9884,N_7083,N_6146);
xnor U9885 (N_9885,N_7984,N_6491);
or U9886 (N_9886,N_6438,N_6199);
nor U9887 (N_9887,N_7758,N_7683);
or U9888 (N_9888,N_6397,N_7375);
xor U9889 (N_9889,N_7746,N_6583);
xor U9890 (N_9890,N_7205,N_6929);
nor U9891 (N_9891,N_6983,N_7289);
nand U9892 (N_9892,N_6862,N_6129);
nor U9893 (N_9893,N_6013,N_6692);
and U9894 (N_9894,N_6826,N_7864);
nor U9895 (N_9895,N_7581,N_6219);
nand U9896 (N_9896,N_7853,N_6598);
or U9897 (N_9897,N_7242,N_7254);
or U9898 (N_9898,N_6825,N_7820);
nand U9899 (N_9899,N_7735,N_6085);
or U9900 (N_9900,N_6288,N_7675);
or U9901 (N_9901,N_6216,N_6288);
xnor U9902 (N_9902,N_7956,N_7703);
or U9903 (N_9903,N_7615,N_7093);
and U9904 (N_9904,N_7798,N_6761);
xor U9905 (N_9905,N_7684,N_7668);
nor U9906 (N_9906,N_7613,N_7383);
nand U9907 (N_9907,N_6451,N_7724);
nor U9908 (N_9908,N_7204,N_7592);
nand U9909 (N_9909,N_6607,N_7655);
nand U9910 (N_9910,N_6976,N_6722);
and U9911 (N_9911,N_6379,N_6804);
and U9912 (N_9912,N_6045,N_7103);
and U9913 (N_9913,N_6591,N_7622);
and U9914 (N_9914,N_6907,N_7857);
nand U9915 (N_9915,N_7373,N_6197);
or U9916 (N_9916,N_6422,N_6673);
or U9917 (N_9917,N_6060,N_6035);
nor U9918 (N_9918,N_7451,N_6609);
or U9919 (N_9919,N_7224,N_6056);
xor U9920 (N_9920,N_7624,N_6081);
or U9921 (N_9921,N_7710,N_7337);
and U9922 (N_9922,N_6610,N_7669);
nand U9923 (N_9923,N_7615,N_6864);
nor U9924 (N_9924,N_7722,N_6117);
and U9925 (N_9925,N_7833,N_6390);
and U9926 (N_9926,N_7227,N_7540);
nand U9927 (N_9927,N_7778,N_6739);
nor U9928 (N_9928,N_7702,N_6766);
nand U9929 (N_9929,N_7427,N_6569);
and U9930 (N_9930,N_7351,N_7006);
and U9931 (N_9931,N_6844,N_7067);
nor U9932 (N_9932,N_6584,N_7370);
nand U9933 (N_9933,N_7297,N_7169);
nand U9934 (N_9934,N_7694,N_7644);
or U9935 (N_9935,N_7105,N_6926);
nor U9936 (N_9936,N_7513,N_6164);
nand U9937 (N_9937,N_7416,N_7328);
and U9938 (N_9938,N_7627,N_7923);
xor U9939 (N_9939,N_7890,N_6998);
and U9940 (N_9940,N_7289,N_7314);
nand U9941 (N_9941,N_6283,N_6999);
nor U9942 (N_9942,N_6942,N_6593);
xnor U9943 (N_9943,N_6684,N_6666);
nand U9944 (N_9944,N_6910,N_6901);
nand U9945 (N_9945,N_6473,N_7950);
and U9946 (N_9946,N_7548,N_7287);
or U9947 (N_9947,N_6957,N_7492);
or U9948 (N_9948,N_6202,N_7597);
nor U9949 (N_9949,N_7062,N_6114);
nor U9950 (N_9950,N_7344,N_6059);
nor U9951 (N_9951,N_7896,N_7031);
and U9952 (N_9952,N_7192,N_6303);
and U9953 (N_9953,N_6897,N_6361);
nor U9954 (N_9954,N_6780,N_7198);
xor U9955 (N_9955,N_7114,N_6478);
or U9956 (N_9956,N_7473,N_7376);
nor U9957 (N_9957,N_6726,N_7024);
nor U9958 (N_9958,N_7581,N_6023);
and U9959 (N_9959,N_7241,N_6676);
nor U9960 (N_9960,N_7772,N_7115);
xnor U9961 (N_9961,N_6316,N_7238);
nor U9962 (N_9962,N_7290,N_7335);
and U9963 (N_9963,N_6168,N_6980);
nand U9964 (N_9964,N_6636,N_7472);
and U9965 (N_9965,N_6255,N_7968);
nand U9966 (N_9966,N_6338,N_7556);
nand U9967 (N_9967,N_7151,N_6150);
xor U9968 (N_9968,N_6599,N_7205);
and U9969 (N_9969,N_7922,N_6431);
nor U9970 (N_9970,N_6333,N_7984);
nor U9971 (N_9971,N_7733,N_6192);
or U9972 (N_9972,N_6893,N_7749);
nor U9973 (N_9973,N_6981,N_7836);
and U9974 (N_9974,N_7047,N_6429);
xor U9975 (N_9975,N_7278,N_6745);
nand U9976 (N_9976,N_7819,N_6963);
nand U9977 (N_9977,N_7454,N_7339);
nand U9978 (N_9978,N_7865,N_7742);
xnor U9979 (N_9979,N_7792,N_7610);
xnor U9980 (N_9980,N_6737,N_6356);
nor U9981 (N_9981,N_7806,N_6918);
nor U9982 (N_9982,N_6993,N_7658);
xor U9983 (N_9983,N_7328,N_6614);
nor U9984 (N_9984,N_7668,N_7117);
and U9985 (N_9985,N_6560,N_7703);
nand U9986 (N_9986,N_6354,N_6921);
nor U9987 (N_9987,N_7072,N_7964);
nor U9988 (N_9988,N_7431,N_6871);
nand U9989 (N_9989,N_6985,N_7769);
nor U9990 (N_9990,N_7098,N_6691);
and U9991 (N_9991,N_6290,N_7940);
nand U9992 (N_9992,N_6226,N_7046);
nor U9993 (N_9993,N_7189,N_7212);
and U9994 (N_9994,N_7191,N_6203);
xor U9995 (N_9995,N_6178,N_6585);
xnor U9996 (N_9996,N_6739,N_7770);
nor U9997 (N_9997,N_7115,N_6189);
nor U9998 (N_9998,N_6201,N_6714);
or U9999 (N_9999,N_6228,N_7711);
nand U10000 (N_10000,N_9367,N_9207);
or U10001 (N_10001,N_8333,N_9497);
nand U10002 (N_10002,N_8827,N_8036);
and U10003 (N_10003,N_9603,N_8566);
and U10004 (N_10004,N_9307,N_8221);
or U10005 (N_10005,N_8606,N_9788);
nor U10006 (N_10006,N_9801,N_8964);
and U10007 (N_10007,N_8884,N_8934);
xor U10008 (N_10008,N_9827,N_9547);
nor U10009 (N_10009,N_8336,N_9115);
nor U10010 (N_10010,N_9310,N_9672);
or U10011 (N_10011,N_9750,N_8233);
and U10012 (N_10012,N_9107,N_8503);
and U10013 (N_10013,N_8726,N_9121);
xnor U10014 (N_10014,N_8498,N_8058);
nand U10015 (N_10015,N_9783,N_8139);
or U10016 (N_10016,N_8168,N_8829);
nand U10017 (N_10017,N_9102,N_8390);
and U10018 (N_10018,N_8300,N_8688);
xnor U10019 (N_10019,N_8536,N_9594);
or U10020 (N_10020,N_8105,N_8895);
nand U10021 (N_10021,N_8999,N_8419);
or U10022 (N_10022,N_8148,N_9640);
nand U10023 (N_10023,N_8949,N_9432);
nor U10024 (N_10024,N_8764,N_9063);
and U10025 (N_10025,N_8893,N_9909);
nand U10026 (N_10026,N_8299,N_8159);
nor U10027 (N_10027,N_8821,N_9775);
nand U10028 (N_10028,N_8152,N_8238);
and U10029 (N_10029,N_8444,N_9957);
xnor U10030 (N_10030,N_8945,N_8201);
nand U10031 (N_10031,N_8661,N_8578);
or U10032 (N_10032,N_8741,N_8252);
nand U10033 (N_10033,N_8158,N_8106);
or U10034 (N_10034,N_9571,N_9154);
xnor U10035 (N_10035,N_8396,N_9913);
or U10036 (N_10036,N_9297,N_9092);
nor U10037 (N_10037,N_9634,N_9922);
or U10038 (N_10038,N_9091,N_8856);
nand U10039 (N_10039,N_9064,N_8501);
xor U10040 (N_10040,N_8351,N_9689);
nand U10041 (N_10041,N_9335,N_9744);
xnor U10042 (N_10042,N_8530,N_8488);
nand U10043 (N_10043,N_9030,N_9430);
and U10044 (N_10044,N_9058,N_8611);
xnor U10045 (N_10045,N_9879,N_9460);
or U10046 (N_10046,N_8743,N_9401);
nor U10047 (N_10047,N_9683,N_9149);
and U10048 (N_10048,N_9085,N_8185);
and U10049 (N_10049,N_8648,N_8593);
or U10050 (N_10050,N_8886,N_9165);
xnor U10051 (N_10051,N_8507,N_9754);
and U10052 (N_10052,N_8795,N_9444);
and U10053 (N_10053,N_8868,N_9026);
or U10054 (N_10054,N_8265,N_8627);
nand U10055 (N_10055,N_9374,N_9388);
nand U10056 (N_10056,N_9656,N_8974);
xnor U10057 (N_10057,N_8967,N_9824);
or U10058 (N_10058,N_8124,N_8410);
nor U10059 (N_10059,N_9000,N_8815);
nor U10060 (N_10060,N_8184,N_8830);
nor U10061 (N_10061,N_9190,N_8307);
xnor U10062 (N_10062,N_9771,N_8164);
and U10063 (N_10063,N_8162,N_9988);
nor U10064 (N_10064,N_8271,N_9059);
nor U10065 (N_10065,N_8891,N_8885);
nor U10066 (N_10066,N_9562,N_9025);
nor U10067 (N_10067,N_8630,N_8855);
nor U10068 (N_10068,N_8644,N_9070);
and U10069 (N_10069,N_8604,N_8624);
nor U10070 (N_10070,N_9651,N_9461);
xor U10071 (N_10071,N_8607,N_9816);
nor U10072 (N_10072,N_8052,N_8636);
or U10073 (N_10073,N_8582,N_9280);
nor U10074 (N_10074,N_9291,N_8090);
xnor U10075 (N_10075,N_9693,N_9441);
or U10076 (N_10076,N_8181,N_9790);
and U10077 (N_10077,N_9109,N_9383);
nor U10078 (N_10078,N_8719,N_9930);
or U10079 (N_10079,N_9950,N_8235);
xnor U10080 (N_10080,N_9815,N_9035);
nor U10081 (N_10081,N_8260,N_9474);
nor U10082 (N_10082,N_9238,N_9519);
and U10083 (N_10083,N_8588,N_8357);
nand U10084 (N_10084,N_9223,N_8877);
nand U10085 (N_10085,N_8943,N_9597);
and U10086 (N_10086,N_8971,N_8857);
and U10087 (N_10087,N_9073,N_9283);
xnor U10088 (N_10088,N_8454,N_8635);
and U10089 (N_10089,N_9966,N_8851);
or U10090 (N_10090,N_9061,N_8189);
or U10091 (N_10091,N_8672,N_8383);
xor U10092 (N_10092,N_8215,N_8027);
or U10093 (N_10093,N_8755,N_9228);
xnor U10094 (N_10094,N_8273,N_8988);
nor U10095 (N_10095,N_8477,N_9567);
and U10096 (N_10096,N_8136,N_9210);
nor U10097 (N_10097,N_8114,N_8178);
xnor U10098 (N_10098,N_9943,N_8825);
and U10099 (N_10099,N_9602,N_8640);
nor U10100 (N_10100,N_9890,N_9434);
xor U10101 (N_10101,N_8750,N_8873);
xnor U10102 (N_10102,N_9256,N_9493);
nor U10103 (N_10103,N_8129,N_8978);
or U10104 (N_10104,N_8199,N_8362);
and U10105 (N_10105,N_9364,N_9264);
nor U10106 (N_10106,N_9160,N_9792);
nand U10107 (N_10107,N_9752,N_8668);
and U10108 (N_10108,N_9103,N_8086);
and U10109 (N_10109,N_8375,N_8935);
nand U10110 (N_10110,N_8789,N_8660);
nand U10111 (N_10111,N_8474,N_9494);
nor U10112 (N_10112,N_9686,N_9868);
xnor U10113 (N_10113,N_9227,N_9077);
and U10114 (N_10114,N_9196,N_8278);
xor U10115 (N_10115,N_9005,N_8443);
or U10116 (N_10116,N_9611,N_9558);
and U10117 (N_10117,N_8460,N_8259);
and U10118 (N_10118,N_8870,N_8203);
xnor U10119 (N_10119,N_9517,N_9167);
nand U10120 (N_10120,N_9089,N_8339);
nor U10121 (N_10121,N_8956,N_9038);
nor U10122 (N_10122,N_9373,N_9701);
nor U10123 (N_10123,N_8338,N_8962);
nand U10124 (N_10124,N_8898,N_9525);
nor U10125 (N_10125,N_8172,N_9831);
nor U10126 (N_10126,N_8930,N_8631);
xnor U10127 (N_10127,N_9886,N_9755);
xor U10128 (N_10128,N_9576,N_8732);
or U10129 (N_10129,N_9719,N_9990);
xnor U10130 (N_10130,N_9372,N_8369);
and U10131 (N_10131,N_9963,N_8428);
xnor U10132 (N_10132,N_8526,N_8775);
and U10133 (N_10133,N_8133,N_9054);
and U10134 (N_10134,N_9318,N_8716);
nor U10135 (N_10135,N_9599,N_8564);
xnor U10136 (N_10136,N_9095,N_9222);
nand U10137 (N_10137,N_8277,N_9407);
and U10138 (N_10138,N_8093,N_9176);
nor U10139 (N_10139,N_8850,N_9637);
nor U10140 (N_10140,N_9437,N_8788);
xnor U10141 (N_10141,N_9426,N_8349);
xor U10142 (N_10142,N_8984,N_8459);
and U10143 (N_10143,N_8950,N_9969);
xnor U10144 (N_10144,N_8697,N_8391);
or U10145 (N_10145,N_9546,N_9045);
and U10146 (N_10146,N_9342,N_9803);
xor U10147 (N_10147,N_8149,N_9111);
and U10148 (N_10148,N_9654,N_8513);
nand U10149 (N_10149,N_9496,N_8031);
nor U10150 (N_10150,N_9086,N_8236);
xnor U10151 (N_10151,N_8476,N_8427);
and U10152 (N_10152,N_8774,N_9202);
xor U10153 (N_10153,N_9609,N_8026);
nand U10154 (N_10154,N_9200,N_8916);
nor U10155 (N_10155,N_8959,N_9022);
xnor U10156 (N_10156,N_9266,N_8389);
or U10157 (N_10157,N_8785,N_8304);
nor U10158 (N_10158,N_8563,N_8506);
xor U10159 (N_10159,N_8596,N_8126);
xnor U10160 (N_10160,N_8077,N_9216);
nand U10161 (N_10161,N_9302,N_8312);
or U10162 (N_10162,N_8276,N_9076);
nand U10163 (N_10163,N_8509,N_9564);
nor U10164 (N_10164,N_9958,N_9606);
nor U10165 (N_10165,N_8899,N_9764);
and U10166 (N_10166,N_9860,N_8284);
or U10167 (N_10167,N_8489,N_9666);
nand U10168 (N_10168,N_9285,N_8973);
and U10169 (N_10169,N_9119,N_9117);
or U10170 (N_10170,N_9315,N_9986);
nor U10171 (N_10171,N_9728,N_8534);
xor U10172 (N_10172,N_9415,N_8352);
nor U10173 (N_10173,N_9970,N_8330);
and U10174 (N_10174,N_8034,N_9604);
nor U10175 (N_10175,N_8681,N_8257);
or U10176 (N_10176,N_8388,N_9774);
nor U10177 (N_10177,N_9233,N_8229);
xor U10178 (N_10178,N_8294,N_9902);
nor U10179 (N_10179,N_9057,N_9447);
nand U10180 (N_10180,N_8659,N_9428);
xor U10181 (N_10181,N_9470,N_9747);
nor U10182 (N_10182,N_9685,N_9305);
nand U10183 (N_10183,N_9742,N_8015);
and U10184 (N_10184,N_9811,N_8571);
and U10185 (N_10185,N_8552,N_9463);
xor U10186 (N_10186,N_8261,N_8160);
xnor U10187 (N_10187,N_9659,N_8426);
or U10188 (N_10188,N_8332,N_8224);
xnor U10189 (N_10189,N_9559,N_8429);
or U10190 (N_10190,N_8628,N_9144);
nand U10191 (N_10191,N_8790,N_8544);
and U10192 (N_10192,N_9158,N_8134);
xor U10193 (N_10193,N_9633,N_8197);
nand U10194 (N_10194,N_8061,N_9492);
and U10195 (N_10195,N_9273,N_9338);
xor U10196 (N_10196,N_9612,N_8449);
nor U10197 (N_10197,N_8654,N_9740);
nand U10198 (N_10198,N_8110,N_9096);
or U10199 (N_10199,N_8594,N_9584);
and U10200 (N_10200,N_9487,N_9588);
or U10201 (N_10201,N_9613,N_9593);
xor U10202 (N_10202,N_9143,N_8655);
or U10203 (N_10203,N_8558,N_9263);
and U10204 (N_10204,N_8980,N_9359);
xor U10205 (N_10205,N_8359,N_8046);
nand U10206 (N_10206,N_9776,N_9015);
nor U10207 (N_10207,N_8639,N_8206);
nor U10208 (N_10208,N_8976,N_8067);
nand U10209 (N_10209,N_9646,N_9229);
and U10210 (N_10210,N_9334,N_9994);
or U10211 (N_10211,N_9218,N_9258);
nand U10212 (N_10212,N_8752,N_9292);
nor U10213 (N_10213,N_9810,N_8609);
nand U10214 (N_10214,N_9748,N_8524);
and U10215 (N_10215,N_9753,N_9473);
xnor U10216 (N_10216,N_9381,N_8314);
nor U10217 (N_10217,N_9676,N_8065);
nor U10218 (N_10218,N_8037,N_8615);
and U10219 (N_10219,N_8953,N_9137);
nor U10220 (N_10220,N_9684,N_8985);
xor U10221 (N_10221,N_8580,N_8423);
or U10222 (N_10222,N_8363,N_8869);
xnor U10223 (N_10223,N_9433,N_9142);
nand U10224 (N_10224,N_8192,N_9320);
nand U10225 (N_10225,N_9959,N_8220);
and U10226 (N_10226,N_8119,N_9663);
xor U10227 (N_10227,N_8658,N_8603);
and U10228 (N_10228,N_9365,N_9925);
or U10229 (N_10229,N_9888,N_8335);
xor U10230 (N_10230,N_8499,N_8007);
and U10231 (N_10231,N_9467,N_9056);
xor U10232 (N_10232,N_9452,N_9583);
xor U10233 (N_10233,N_9246,N_8882);
xnor U10234 (N_10234,N_9626,N_8667);
nand U10235 (N_10235,N_9175,N_9449);
nand U10236 (N_10236,N_9671,N_8135);
and U10237 (N_10237,N_8466,N_8584);
or U10238 (N_10238,N_9491,N_8103);
nor U10239 (N_10239,N_9270,N_9234);
nor U10240 (N_10240,N_8434,N_9806);
nor U10241 (N_10241,N_8720,N_8242);
or U10242 (N_10242,N_8770,N_8263);
nand U10243 (N_10243,N_9841,N_8432);
or U10244 (N_10244,N_9608,N_8515);
or U10245 (N_10245,N_9768,N_8979);
or U10246 (N_10246,N_8002,N_8791);
and U10247 (N_10247,N_9239,N_8048);
or U10248 (N_10248,N_9509,N_8938);
xor U10249 (N_10249,N_9729,N_8468);
xnor U10250 (N_10250,N_8568,N_8188);
xor U10251 (N_10251,N_8812,N_9206);
and U10252 (N_10252,N_8853,N_9314);
or U10253 (N_10253,N_9923,N_9514);
and U10254 (N_10254,N_8703,N_8068);
nand U10255 (N_10255,N_8900,N_9380);
nand U10256 (N_10256,N_9842,N_8486);
nor U10257 (N_10257,N_8292,N_9850);
nor U10258 (N_10258,N_8217,N_8577);
or U10259 (N_10259,N_9653,N_8792);
nand U10260 (N_10260,N_9741,N_9173);
xnor U10261 (N_10261,N_9697,N_9155);
xnor U10262 (N_10262,N_9882,N_8347);
nor U10263 (N_10263,N_9442,N_8707);
and U10264 (N_10264,N_8940,N_8019);
nand U10265 (N_10265,N_8711,N_9766);
xnor U10266 (N_10266,N_8632,N_9551);
or U10267 (N_10267,N_9087,N_8927);
nor U10268 (N_10268,N_8418,N_9717);
or U10269 (N_10269,N_9533,N_9066);
nand U10270 (N_10270,N_9260,N_9140);
nand U10271 (N_10271,N_9733,N_8968);
nor U10272 (N_10272,N_8574,N_9642);
xnor U10273 (N_10273,N_8128,N_9503);
or U10274 (N_10274,N_8537,N_8166);
or U10275 (N_10275,N_9550,N_8921);
nor U10276 (N_10276,N_8431,N_8480);
xor U10277 (N_10277,N_9907,N_9631);
nor U10278 (N_10278,N_9080,N_9431);
nor U10279 (N_10279,N_9702,N_8003);
nor U10280 (N_10280,N_8186,N_9134);
nor U10281 (N_10281,N_9561,N_9548);
and U10282 (N_10282,N_8863,N_8520);
or U10283 (N_10283,N_9100,N_9139);
and U10284 (N_10284,N_9802,N_8319);
or U10285 (N_10285,N_9664,N_8137);
and U10286 (N_10286,N_9472,N_9483);
or U10287 (N_10287,N_8424,N_8478);
nand U10288 (N_10288,N_8266,N_9813);
xnor U10289 (N_10289,N_9756,N_8992);
nor U10290 (N_10290,N_8806,N_8514);
xnor U10291 (N_10291,N_9214,N_8457);
and U10292 (N_10292,N_8017,N_9869);
xor U10293 (N_10293,N_8044,N_9569);
nor U10294 (N_10294,N_8972,N_8049);
or U10295 (N_10295,N_9481,N_8694);
and U10296 (N_10296,N_9624,N_9168);
xor U10297 (N_10297,N_9031,N_9510);
or U10298 (N_10298,N_8268,N_8724);
nor U10299 (N_10299,N_9647,N_9159);
nor U10300 (N_10300,N_9895,N_8715);
and U10301 (N_10301,N_9166,N_9241);
nor U10302 (N_10302,N_9678,N_8011);
xor U10303 (N_10303,N_8780,N_8174);
nor U10304 (N_10304,N_8547,N_9982);
or U10305 (N_10305,N_9275,N_8808);
xnor U10306 (N_10306,N_9615,N_8045);
nor U10307 (N_10307,N_9319,N_8226);
xor U10308 (N_10308,N_8686,N_9469);
nor U10309 (N_10309,N_9462,N_9544);
nor U10310 (N_10310,N_9712,N_9713);
nand U10311 (N_10311,N_9985,N_8932);
and U10312 (N_10312,N_9916,N_9249);
nand U10313 (N_10313,N_9820,N_9013);
nand U10314 (N_10314,N_8028,N_8532);
xor U10315 (N_10315,N_9526,N_9759);
nand U10316 (N_10316,N_9295,N_8545);
and U10317 (N_10317,N_9761,N_9377);
nand U10318 (N_10318,N_9681,N_9967);
xor U10319 (N_10319,N_9975,N_8907);
nand U10320 (N_10320,N_9037,N_8308);
nand U10321 (N_10321,N_8413,N_8961);
or U10322 (N_10322,N_9069,N_8010);
and U10323 (N_10323,N_9534,N_8098);
nor U10324 (N_10324,N_9688,N_8915);
nor U10325 (N_10325,N_8747,N_8843);
and U10326 (N_10326,N_8749,N_9255);
or U10327 (N_10327,N_9090,N_8144);
nand U10328 (N_10328,N_9271,N_8100);
xor U10329 (N_10329,N_9772,N_9456);
xnor U10330 (N_10330,N_9901,N_9696);
or U10331 (N_10331,N_9789,N_8182);
or U10332 (N_10332,N_8387,N_9502);
nand U10333 (N_10333,N_9840,N_9252);
nand U10334 (N_10334,N_8784,N_9829);
xor U10335 (N_10335,N_8190,N_9240);
or U10336 (N_10336,N_9511,N_8511);
xor U10337 (N_10337,N_8009,N_9834);
and U10338 (N_10338,N_8324,N_8112);
nand U10339 (N_10339,N_8161,N_8380);
or U10340 (N_10340,N_9455,N_8062);
nand U10341 (N_10341,N_9627,N_8113);
nor U10342 (N_10342,N_8165,N_8701);
or U10343 (N_10343,N_9410,N_8523);
or U10344 (N_10344,N_9505,N_9589);
xor U10345 (N_10345,N_9288,N_8376);
and U10346 (N_10346,N_8721,N_9849);
nand U10347 (N_10347,N_8327,N_8814);
xnor U10348 (N_10348,N_9284,N_8579);
nand U10349 (N_10349,N_8072,N_9644);
xnor U10350 (N_10350,N_8625,N_9971);
xor U10351 (N_10351,N_8794,N_8782);
and U10352 (N_10352,N_8573,N_9325);
and U10353 (N_10353,N_9354,N_8231);
or U10354 (N_10354,N_9230,N_9204);
xor U10355 (N_10355,N_9443,N_9478);
xnor U10356 (N_10356,N_8592,N_8177);
nand U10357 (N_10357,N_8772,N_9313);
and U10358 (N_10358,N_8321,N_8282);
and U10359 (N_10359,N_9565,N_9244);
and U10360 (N_10360,N_8766,N_9545);
or U10361 (N_10361,N_9440,N_9339);
or U10362 (N_10362,N_9570,N_9859);
nand U10363 (N_10363,N_9251,N_9427);
and U10364 (N_10364,N_8228,N_9261);
xnor U10365 (N_10365,N_8797,N_8078);
xor U10366 (N_10366,N_9865,N_8102);
xnor U10367 (N_10367,N_9527,N_8286);
nor U10368 (N_10368,N_8483,N_9413);
nand U10369 (N_10369,N_8080,N_8251);
nand U10370 (N_10370,N_8920,N_8637);
nor U10371 (N_10371,N_9189,N_8709);
nor U10372 (N_10372,N_8723,N_8810);
nor U10373 (N_10373,N_8942,N_9516);
and U10374 (N_10374,N_9199,N_9224);
nand U10375 (N_10375,N_8073,N_8533);
or U10376 (N_10376,N_9992,N_9253);
xor U10377 (N_10377,N_9557,N_9304);
or U10378 (N_10378,N_8929,N_8529);
nor U10379 (N_10379,N_9675,N_8140);
xnor U10380 (N_10380,N_9453,N_9591);
nor U10381 (N_10381,N_8946,N_9484);
nand U10382 (N_10382,N_9983,N_8704);
nor U10383 (N_10383,N_9580,N_9282);
or U10384 (N_10384,N_9918,N_8663);
or U10385 (N_10385,N_9408,N_8575);
xnor U10386 (N_10386,N_8816,N_9108);
or U10387 (N_10387,N_9632,N_9984);
and U10388 (N_10388,N_9823,N_9924);
xor U10389 (N_10389,N_8131,N_8315);
nor U10390 (N_10390,N_9822,N_9454);
xnor U10391 (N_10391,N_9543,N_8599);
nor U10392 (N_10392,N_8370,N_8902);
or U10393 (N_10393,N_8130,N_9861);
nand U10394 (N_10394,N_9358,N_8281);
and U10395 (N_10395,N_9785,N_8598);
or U10396 (N_10396,N_8991,N_9677);
nor U10397 (N_10397,N_8095,N_8758);
nor U10398 (N_10398,N_9231,N_9274);
and U10399 (N_10399,N_9172,N_9851);
nand U10400 (N_10400,N_9660,N_9395);
nor U10401 (N_10401,N_8469,N_9931);
and U10402 (N_10402,N_9787,N_9948);
or U10403 (N_10403,N_9555,N_8381);
or U10404 (N_10404,N_8504,N_8951);
and U10405 (N_10405,N_9769,N_8092);
nand U10406 (N_10406,N_9217,N_8082);
nor U10407 (N_10407,N_9997,N_8289);
and U10408 (N_10408,N_8997,N_9120);
or U10409 (N_10409,N_9186,N_8183);
and U10410 (N_10410,N_8502,N_8412);
or U10411 (N_10411,N_8646,N_9665);
and U10412 (N_10412,N_8919,N_9060);
and U10413 (N_10413,N_8645,N_9021);
nand U10414 (N_10414,N_8737,N_8617);
xor U10415 (N_10415,N_8691,N_9670);
nand U10416 (N_10416,N_9479,N_9575);
nand U10417 (N_10417,N_9418,N_9490);
nand U10418 (N_10418,N_8302,N_8897);
nand U10419 (N_10419,N_9438,N_9873);
nand U10420 (N_10420,N_8731,N_8892);
nor U10421 (N_10421,N_9385,N_8053);
nor U10422 (N_10422,N_9743,N_8804);
or U10423 (N_10423,N_9906,N_9760);
nand U10424 (N_10424,N_9489,N_9695);
nor U10425 (N_10425,N_8342,N_9301);
nor U10426 (N_10426,N_9537,N_8417);
nor U10427 (N_10427,N_9679,N_8416);
nor U10428 (N_10428,N_8211,N_9682);
and U10429 (N_10429,N_9530,N_9250);
xnor U10430 (N_10430,N_9641,N_8683);
xnor U10431 (N_10431,N_8084,N_8005);
or U10432 (N_10432,N_9912,N_9457);
nand U10433 (N_10433,N_9303,N_9587);
xnor U10434 (N_10434,N_8690,N_8727);
nand U10435 (N_10435,N_8982,N_8702);
or U10436 (N_10436,N_8759,N_9830);
or U10437 (N_10437,N_8908,N_9786);
and U10438 (N_10438,N_8518,N_8372);
or U10439 (N_10439,N_9836,N_8297);
nand U10440 (N_10440,N_8029,N_8056);
or U10441 (N_10441,N_8783,N_9933);
or U10442 (N_10442,N_8569,N_9177);
nand U10443 (N_10443,N_8484,N_9541);
nand U10444 (N_10444,N_8762,N_9855);
nand U10445 (N_10445,N_9480,N_8662);
and U10446 (N_10446,N_8722,N_8024);
nand U10447 (N_10447,N_9193,N_9075);
nor U10448 (N_10448,N_9600,N_9347);
or U10449 (N_10449,N_9884,N_8831);
xor U10450 (N_10450,N_9420,N_9122);
xnor U10451 (N_10451,N_9521,N_9795);
xor U10452 (N_10452,N_9732,N_9114);
or U10453 (N_10453,N_8364,N_9356);
nor U10454 (N_10454,N_9046,N_8666);
nor U10455 (N_10455,N_9093,N_8121);
nand U10456 (N_10456,N_9390,N_8448);
nor U10457 (N_10457,N_9917,N_9024);
xor U10458 (N_10458,N_9581,N_8917);
or U10459 (N_10459,N_9536,N_8393);
nor U10460 (N_10460,N_8904,N_8420);
and U10461 (N_10461,N_8554,N_8652);
nand U10462 (N_10462,N_8032,N_8865);
or U10463 (N_10463,N_8163,N_8777);
nor U10464 (N_10464,N_8763,N_9343);
or U10465 (N_10465,N_8358,N_8958);
or U10466 (N_10466,N_8329,N_9235);
xor U10467 (N_10467,N_9048,N_9928);
nor U10468 (N_10468,N_8400,N_8993);
nor U10469 (N_10469,N_9911,N_8151);
nor U10470 (N_10470,N_9028,N_8482);
nand U10471 (N_10471,N_8353,N_8481);
or U10472 (N_10472,N_9208,N_8705);
and U10473 (N_10473,N_9616,N_8600);
xnor U10474 (N_10474,N_9946,N_9691);
nand U10475 (N_10475,N_9017,N_9745);
nor U10476 (N_10476,N_9082,N_9498);
or U10477 (N_10477,N_8006,N_8208);
nand U10478 (N_10478,N_8793,N_8279);
or U10479 (N_10479,N_9553,N_9586);
nand U10480 (N_10480,N_8415,N_8022);
xor U10481 (N_10481,N_9138,N_9248);
nor U10482 (N_10482,N_8998,N_9673);
nand U10483 (N_10483,N_9905,N_8728);
nand U10484 (N_10484,N_9953,N_9996);
or U10485 (N_10485,N_9826,N_8097);
xor U10486 (N_10486,N_8733,N_8800);
nand U10487 (N_10487,N_8685,N_9221);
and U10488 (N_10488,N_8761,N_9891);
and U10489 (N_10489,N_8861,N_8633);
or U10490 (N_10490,N_9191,N_8004);
or U10491 (N_10491,N_9819,N_9780);
and U10492 (N_10492,N_8512,N_9052);
nand U10493 (N_10493,N_9669,N_9779);
nor U10494 (N_10494,N_8404,N_9724);
and U10495 (N_10495,N_9044,N_8854);
nand U10496 (N_10496,N_9018,N_9378);
or U10497 (N_10497,N_8495,N_8414);
nor U10498 (N_10498,N_8205,N_9722);
xnor U10499 (N_10499,N_9770,N_8778);
xor U10500 (N_10500,N_8346,N_9084);
nor U10501 (N_10501,N_9704,N_8977);
and U10502 (N_10502,N_9105,N_9366);
nand U10503 (N_10503,N_9707,N_8247);
and U10504 (N_10504,N_8179,N_9466);
nor U10505 (N_10505,N_8207,N_8440);
nor U10506 (N_10506,N_9535,N_9500);
or U10507 (N_10507,N_9808,N_8933);
nor U10508 (N_10508,N_8223,N_9773);
or U10509 (N_10509,N_9579,N_9952);
nand U10510 (N_10510,N_8910,N_9327);
and U10511 (N_10511,N_9552,N_8280);
nor U10512 (N_10512,N_9399,N_8407);
xnor U10513 (N_10513,N_8613,N_8670);
nand U10514 (N_10514,N_8008,N_8167);
xor U10515 (N_10515,N_9636,N_8669);
and U10516 (N_10516,N_9311,N_9972);
xor U10517 (N_10517,N_8653,N_8210);
nand U10518 (N_10518,N_8757,N_9951);
nor U10519 (N_10519,N_8647,N_8708);
xnor U10520 (N_10520,N_8664,N_8612);
or U10521 (N_10521,N_9614,N_9978);
or U10522 (N_10522,N_9286,N_9904);
and U10523 (N_10523,N_8425,N_9881);
or U10524 (N_10524,N_9147,N_8948);
xnor U10525 (N_10525,N_8535,N_8249);
and U10526 (N_10526,N_9170,N_9574);
or U10527 (N_10527,N_8127,N_8805);
nor U10528 (N_10528,N_8883,N_9345);
nor U10529 (N_10529,N_8714,N_9932);
or U10530 (N_10530,N_9039,N_9556);
nor U10531 (N_10531,N_8881,N_9053);
or U10532 (N_10532,N_9324,N_9099);
and U10533 (N_10533,N_9947,N_8014);
or U10534 (N_10534,N_9939,N_8587);
or U10535 (N_10535,N_8813,N_8066);
nand U10536 (N_10536,N_8879,N_9718);
xor U10537 (N_10537,N_8202,N_8059);
xor U10538 (N_10538,N_8698,N_8699);
or U10539 (N_10539,N_8994,N_8505);
nand U10540 (N_10540,N_8385,N_8889);
nor U10541 (N_10541,N_8963,N_9921);
and U10542 (N_10542,N_8435,N_9871);
xnor U10543 (N_10543,N_9384,N_9723);
and U10544 (N_10544,N_9033,N_9910);
nor U10545 (N_10545,N_9645,N_9885);
nand U10546 (N_10546,N_9781,N_8754);
xnor U10547 (N_10547,N_9237,N_8550);
nor U10548 (N_10548,N_9362,N_8142);
xor U10549 (N_10549,N_8384,N_9839);
nand U10550 (N_10550,N_9965,N_8291);
nor U10551 (N_10551,N_8510,N_9330);
xnor U10552 (N_10552,N_8786,N_9499);
nor U10553 (N_10553,N_8490,N_9908);
or U10554 (N_10554,N_8340,N_8913);
or U10555 (N_10555,N_8194,N_9268);
xor U10556 (N_10556,N_9735,N_9486);
xor U10557 (N_10557,N_9226,N_8000);
or U10558 (N_10558,N_9605,N_8925);
and U10559 (N_10559,N_9876,N_9520);
and U10560 (N_10560,N_8043,N_9353);
or U10561 (N_10561,N_9817,N_8155);
xor U10562 (N_10562,N_9949,N_9414);
xnor U10563 (N_10563,N_9412,N_8693);
nand U10564 (N_10564,N_8912,N_9488);
nor U10565 (N_10565,N_8840,N_9185);
or U10566 (N_10566,N_9051,N_9955);
nand U10567 (N_10567,N_8906,N_8088);
nor U10568 (N_10568,N_9094,N_8562);
nand U10569 (N_10569,N_8303,N_9267);
or U10570 (N_10570,N_9777,N_9716);
or U10571 (N_10571,N_9515,N_9123);
or U10572 (N_10572,N_9162,N_8542);
xnor U10573 (N_10573,N_8802,N_8862);
xnor U10574 (N_10574,N_8473,N_8819);
xnor U10575 (N_10575,N_9814,N_8262);
nor U10576 (N_10576,N_9153,N_8331);
nor U10577 (N_10577,N_8436,N_9308);
xnor U10578 (N_10578,N_8341,N_9898);
or U10579 (N_10579,N_8888,N_9538);
and U10580 (N_10580,N_9648,N_9577);
and U10581 (N_10581,N_9393,N_8348);
and U10582 (N_10582,N_8608,N_8253);
xnor U10583 (N_10583,N_9845,N_9629);
or U10584 (N_10584,N_9734,N_9794);
nand U10585 (N_10585,N_8494,N_8641);
and U10586 (N_10586,N_9419,N_8595);
xnor U10587 (N_10587,N_9477,N_8619);
nor U10588 (N_10588,N_8695,N_8894);
xnor U10589 (N_10589,N_8651,N_9623);
xor U10590 (N_10590,N_8366,N_8572);
and U10591 (N_10591,N_9409,N_8960);
and U10592 (N_10592,N_9899,N_9767);
or U10593 (N_10593,N_9265,N_8560);
xnor U10594 (N_10594,N_9620,N_8649);
nor U10595 (N_10595,N_9299,N_9857);
and U10596 (N_10596,N_9655,N_9513);
or U10597 (N_10597,N_9067,N_9833);
and U10598 (N_10598,N_8195,N_9336);
or U10599 (N_10599,N_9661,N_9179);
and U10600 (N_10600,N_9294,N_8479);
and U10601 (N_10601,N_8154,N_9807);
or U10602 (N_10602,N_8467,N_9690);
and U10603 (N_10603,N_8125,N_8849);
or U10604 (N_10604,N_8403,N_9880);
and U10605 (N_10605,N_8779,N_8887);
or U10606 (N_10606,N_8108,N_8272);
and U10607 (N_10607,N_8634,N_8039);
nand U10608 (N_10608,N_8230,N_8665);
or U10609 (N_10609,N_9711,N_8241);
nor U10610 (N_10610,N_8471,N_9009);
nand U10611 (N_10611,N_9391,N_8845);
and U10612 (N_10612,N_9706,N_8621);
xor U10613 (N_10613,N_8620,N_9436);
nor U10614 (N_10614,N_9406,N_9317);
and U10615 (N_10615,N_8063,N_9269);
nor U10616 (N_10616,N_9981,N_8169);
nand U10617 (N_10617,N_8903,N_9793);
nand U10618 (N_10618,N_9194,N_9348);
nor U10619 (N_10619,N_8016,N_8947);
nand U10620 (N_10620,N_9800,N_8150);
nand U10621 (N_10621,N_9281,N_9145);
or U10622 (N_10622,N_8955,N_8911);
nor U10623 (N_10623,N_9797,N_9116);
nor U10624 (N_10624,N_8213,N_8767);
and U10625 (N_10625,N_8876,N_9867);
xor U10626 (N_10626,N_8225,N_9146);
xor U10627 (N_10627,N_8567,N_9279);
and U10628 (N_10628,N_8739,N_8328);
nand U10629 (N_10629,N_8710,N_8406);
or U10630 (N_10630,N_8836,N_9687);
or U10631 (N_10631,N_8064,N_9680);
nand U10632 (N_10632,N_8405,N_9872);
and U10633 (N_10633,N_9607,N_9023);
nand U10634 (N_10634,N_8408,N_8047);
nand U10635 (N_10635,N_8138,N_8656);
xor U10636 (N_10636,N_8275,N_9425);
or U10637 (N_10637,N_8966,N_9163);
or U10638 (N_10638,N_8222,N_8549);
or U10639 (N_10639,N_9088,N_9980);
nand U10640 (N_10640,N_8847,N_8838);
or U10641 (N_10641,N_9812,N_9529);
xnor U10642 (N_10642,N_8890,N_8288);
nor U10643 (N_10643,N_8023,N_9277);
or U10644 (N_10644,N_8191,N_8954);
nor U10645 (N_10645,N_9954,N_8018);
nor U10646 (N_10646,N_9847,N_8117);
and U10647 (N_10647,N_9055,N_8101);
or U10648 (N_10648,N_8451,N_9370);
nand U10649 (N_10649,N_8492,N_8751);
nand U10650 (N_10650,N_9298,N_8132);
nand U10651 (N_10651,N_8475,N_8555);
xnor U10652 (N_10652,N_9394,N_9012);
or U10653 (N_10653,N_8543,N_8123);
nor U10654 (N_10654,N_9762,N_8522);
and U10655 (N_10655,N_8712,N_9131);
xnor U10656 (N_10656,N_9936,N_9598);
xor U10657 (N_10657,N_9278,N_8025);
xnor U10658 (N_10658,N_8232,N_8089);
nor U10659 (N_10659,N_9763,N_9007);
xnor U10660 (N_10660,N_9411,N_9259);
nand U10661 (N_10661,N_9848,N_9350);
or U10662 (N_10662,N_9508,N_8957);
nand U10663 (N_10663,N_8834,N_9796);
or U10664 (N_10664,N_8343,N_9262);
xnor U10665 (N_10665,N_8107,N_8219);
nand U10666 (N_10666,N_8674,N_9977);
nor U10667 (N_10667,N_9662,N_9862);
and U10668 (N_10668,N_8776,N_8682);
nor U10669 (N_10669,N_9464,N_8528);
or U10670 (N_10670,N_9549,N_8030);
nand U10671 (N_10671,N_8296,N_8246);
or U10672 (N_10672,N_9074,N_8638);
nor U10673 (N_10673,N_9874,N_8866);
nor U10674 (N_10674,N_8736,N_8872);
nand U10675 (N_10675,N_8643,N_8931);
xor U10676 (N_10676,N_8500,N_9821);
nand U10677 (N_10677,N_8941,N_8760);
nand U10678 (N_10678,N_9198,N_9184);
or U10679 (N_10679,N_9476,N_9065);
xor U10680 (N_10680,N_8824,N_9495);
nand U10681 (N_10681,N_8801,N_8990);
nand U10682 (N_10682,N_8622,N_8684);
and U10683 (N_10683,N_9991,N_9531);
xnor U10684 (N_10684,N_9858,N_8673);
and U10685 (N_10685,N_8392,N_8875);
nor U10686 (N_10686,N_9316,N_8051);
and U10687 (N_10687,N_9344,N_8896);
or U10688 (N_10688,N_9081,N_9136);
nand U10689 (N_10689,N_9746,N_8074);
xnor U10690 (N_10690,N_8811,N_8020);
or U10691 (N_10691,N_8965,N_9195);
nand U10692 (N_10692,N_9150,N_9995);
and U10693 (N_10693,N_9694,N_9903);
or U10694 (N_10694,N_9507,N_9225);
nor U10695 (N_10695,N_8243,N_9504);
nand U10696 (N_10696,N_8334,N_9751);
nand U10697 (N_10697,N_9894,N_8924);
or U10698 (N_10698,N_8987,N_8995);
nor U10699 (N_10699,N_9778,N_9458);
nor U10700 (N_10700,N_8939,N_8399);
and U10701 (N_10701,N_9188,N_9323);
nand U10702 (N_10702,N_8521,N_8290);
and U10703 (N_10703,N_8936,N_9127);
and U10704 (N_10704,N_8700,N_9601);
or U10705 (N_10705,N_9877,N_9448);
nor U10706 (N_10706,N_9582,N_9595);
nand U10707 (N_10707,N_8525,N_9652);
or U10708 (N_10708,N_8311,N_9328);
or U10709 (N_10709,N_9445,N_8070);
xnor U10710 (N_10710,N_8325,N_9113);
nor U10711 (N_10711,N_9171,N_8013);
xor U10712 (N_10712,N_8493,N_8799);
and U10713 (N_10713,N_8298,N_9585);
or U10714 (N_10714,N_8270,N_8527);
and U10715 (N_10715,N_9287,N_8147);
nand U10716 (N_10716,N_9201,N_8832);
nand U10717 (N_10717,N_9212,N_8379);
or U10718 (N_10718,N_9398,N_9112);
or U10719 (N_10719,N_8255,N_8461);
nand U10720 (N_10720,N_8878,N_9043);
xnor U10721 (N_10721,N_8844,N_8085);
xor U10722 (N_10722,N_9156,N_9889);
nor U10723 (N_10723,N_9019,N_9828);
nor U10724 (N_10724,N_9878,N_9765);
and U10725 (N_10725,N_9126,N_8446);
and U10726 (N_10726,N_9182,N_9405);
nand U10727 (N_10727,N_9209,N_9110);
and U10728 (N_10728,N_8310,N_8175);
xor U10729 (N_10729,N_8245,N_8170);
nor U10730 (N_10730,N_9396,N_8871);
or U10731 (N_10731,N_8326,N_8283);
nand U10732 (N_10732,N_9290,N_9563);
nor U10733 (N_10733,N_9832,N_9197);
nand U10734 (N_10734,N_9387,N_9124);
xor U10735 (N_10735,N_8218,N_9423);
nand U10736 (N_10736,N_9389,N_9938);
and U10737 (N_10737,N_8354,N_8553);
or U10738 (N_10738,N_8610,N_9245);
nor U10739 (N_10739,N_9183,N_9866);
and U10740 (N_10740,N_8038,N_9731);
or U10741 (N_10741,N_8173,N_9475);
xnor U10742 (N_10742,N_9625,N_9720);
nand U10743 (N_10743,N_8001,N_8905);
nor U10744 (N_10744,N_9485,N_9083);
nand U10745 (N_10745,N_9326,N_9976);
or U10746 (N_10746,N_9192,N_9942);
or U10747 (N_10747,N_8874,N_8438);
nand U10748 (N_10748,N_8519,N_8371);
xor U10749 (N_10749,N_9072,N_9178);
and U10750 (N_10750,N_8538,N_8350);
and U10751 (N_10751,N_9993,N_8305);
nor U10752 (N_10752,N_8143,N_8671);
nor U10753 (N_10753,N_9130,N_9528);
nor U10754 (N_10754,N_9446,N_9386);
or U10755 (N_10755,N_8601,N_8970);
or U10756 (N_10756,N_9900,N_9376);
xnor U10757 (N_10757,N_8605,N_9011);
xnor U10758 (N_10758,N_9312,N_9337);
and U10759 (N_10759,N_9161,N_8198);
nor U10760 (N_10760,N_9883,N_8557);
and U10761 (N_10761,N_9349,N_8926);
nor U10762 (N_10762,N_9003,N_8180);
nor U10763 (N_10763,N_8293,N_8626);
nand U10764 (N_10764,N_8781,N_9825);
and U10765 (N_10765,N_9439,N_8590);
and U10766 (N_10766,N_9243,N_8422);
nor U10767 (N_10767,N_8923,N_9101);
nand U10768 (N_10768,N_8196,N_9726);
nor U10769 (N_10769,N_8463,N_9118);
nor U10770 (N_10770,N_8952,N_9960);
or U10771 (N_10771,N_9592,N_9272);
nor U10772 (N_10772,N_9036,N_8453);
or U10773 (N_10773,N_9417,N_9935);
and U10774 (N_10774,N_9758,N_8678);
nand U10775 (N_10775,N_9791,N_8200);
nand U10776 (N_10776,N_8337,N_9920);
nand U10777 (N_10777,N_8616,N_8583);
xor U10778 (N_10778,N_8050,N_8817);
and U10779 (N_10779,N_8042,N_9148);
or U10780 (N_10780,N_8642,N_8746);
or U10781 (N_10781,N_8983,N_9875);
and U10782 (N_10782,N_8937,N_8914);
nand U10783 (N_10783,N_8969,N_9020);
nand U10784 (N_10784,N_8239,N_8864);
nor U10785 (N_10785,N_9482,N_9838);
or U10786 (N_10786,N_8909,N_9749);
nor U10787 (N_10787,N_8581,N_9940);
and U10788 (N_10788,N_8576,N_9340);
and U10789 (N_10789,N_8398,N_8287);
and U10790 (N_10790,N_8922,N_8367);
or U10791 (N_10791,N_9341,N_8356);
and U10792 (N_10792,N_8551,N_8437);
xnor U10793 (N_10793,N_8409,N_9518);
nand U10794 (N_10794,N_8753,N_9635);
nand U10795 (N_10795,N_9512,N_8629);
nand U10796 (N_10796,N_9008,N_8837);
nand U10797 (N_10797,N_8718,N_9962);
or U10798 (N_10798,N_9071,N_9351);
nor U10799 (N_10799,N_9180,N_8441);
nor U10800 (N_10800,N_8585,N_8768);
or U10801 (N_10801,N_9042,N_8445);
xnor U10802 (N_10802,N_8378,N_8848);
and U10803 (N_10803,N_8254,N_8455);
nand U10804 (N_10804,N_8111,N_8040);
xnor U10805 (N_10805,N_9361,N_8104);
or U10806 (N_10806,N_9979,N_8989);
xnor U10807 (N_10807,N_8057,N_8301);
or U10808 (N_10808,N_8204,N_8559);
nand U10809 (N_10809,N_8081,N_8244);
and U10810 (N_10810,N_9181,N_8320);
or U10811 (N_10811,N_9657,N_8306);
or U10812 (N_10812,N_8828,N_8809);
nor U10813 (N_10813,N_9782,N_9232);
nand U10814 (N_10814,N_9404,N_9674);
xnor U10815 (N_10815,N_9034,N_8462);
and U10816 (N_10816,N_9375,N_9435);
nor U10817 (N_10817,N_9360,N_8738);
nor U10818 (N_10818,N_9961,N_8382);
and U10819 (N_10819,N_9289,N_8250);
xor U10820 (N_10820,N_8918,N_9539);
nor U10821 (N_10821,N_9738,N_8730);
nor U10822 (N_10822,N_9560,N_9628);
or U10823 (N_10823,N_8264,N_8614);
nor U10824 (N_10824,N_9554,N_9737);
xor U10825 (N_10825,N_9157,N_8773);
or U10826 (N_10826,N_9956,N_9332);
and U10827 (N_10827,N_9424,N_8565);
xnor U10828 (N_10828,N_8803,N_9610);
and U10829 (N_10829,N_9125,N_9129);
or U10830 (N_10830,N_9835,N_8833);
nand U10831 (N_10831,N_9852,N_9974);
and U10832 (N_10832,N_9798,N_9805);
nand U10833 (N_10833,N_9566,N_8060);
or U10834 (N_10834,N_8680,N_9730);
nand U10835 (N_10835,N_8706,N_9128);
or U10836 (N_10836,N_9300,N_8623);
nand U10837 (N_10837,N_8546,N_8485);
and U10838 (N_10838,N_9915,N_8087);
xnor U10839 (N_10839,N_8240,N_8470);
nor U10840 (N_10840,N_8589,N_8541);
xor U10841 (N_10841,N_8374,N_9914);
or U10842 (N_10842,N_9220,N_8115);
and U10843 (N_10843,N_9215,N_8021);
nand U10844 (N_10844,N_9944,N_8237);
nand U10845 (N_10845,N_8570,N_8452);
or U10846 (N_10846,N_9211,N_9524);
nand U10847 (N_10847,N_8083,N_9700);
nand U10848 (N_10848,N_9169,N_8713);
nor U10849 (N_10849,N_9369,N_8487);
xnor U10850 (N_10850,N_8361,N_9422);
nor U10851 (N_10851,N_9929,N_8735);
or U10852 (N_10852,N_9047,N_9715);
nor U10853 (N_10853,N_8787,N_8091);
nand U10854 (N_10854,N_9941,N_8450);
xnor U10855 (N_10855,N_8901,N_8540);
and U10856 (N_10856,N_8256,N_9896);
or U10857 (N_10857,N_9667,N_9864);
xor U10858 (N_10858,N_9618,N_8548);
xor U10859 (N_10859,N_8012,N_8496);
xor U10860 (N_10860,N_8096,N_9973);
and U10861 (N_10861,N_8397,N_8071);
nor U10862 (N_10862,N_9247,N_8216);
or U10863 (N_10863,N_8075,N_8839);
and U10864 (N_10864,N_9471,N_9346);
and U10865 (N_10865,N_8234,N_9870);
and U10866 (N_10866,N_8986,N_9709);
nand U10867 (N_10867,N_9998,N_8464);
and U10868 (N_10868,N_8439,N_8394);
nor U10869 (N_10869,N_9368,N_8055);
or U10870 (N_10870,N_8798,N_8248);
or U10871 (N_10871,N_9151,N_8586);
xor U10872 (N_10872,N_8725,N_9402);
nand U10873 (N_10873,N_9465,N_9721);
or U10874 (N_10874,N_9621,N_8316);
xor U10875 (N_10875,N_8472,N_9331);
nor U10876 (N_10876,N_9133,N_9152);
nor U10877 (N_10877,N_8675,N_8365);
and U10878 (N_10878,N_8122,N_9293);
nor U10879 (N_10879,N_9727,N_9987);
nor U10880 (N_10880,N_8373,N_8345);
or U10881 (N_10881,N_8187,N_9506);
or U10882 (N_10882,N_8852,N_9863);
nand U10883 (N_10883,N_9050,N_8650);
or U10884 (N_10884,N_9329,N_9242);
nand U10885 (N_10885,N_9989,N_8212);
nand U10886 (N_10886,N_8402,N_9135);
nor U10887 (N_10887,N_8386,N_8740);
nor U10888 (N_10888,N_9400,N_8076);
and U10889 (N_10889,N_9236,N_9078);
nand U10890 (N_10890,N_9968,N_9416);
nor U10891 (N_10891,N_8313,N_9106);
nand U10892 (N_10892,N_9843,N_8771);
nand U10893 (N_10893,N_9403,N_8069);
nor U10894 (N_10894,N_9049,N_8355);
nor U10895 (N_10895,N_9010,N_9379);
or U10896 (N_10896,N_9104,N_8285);
nor U10897 (N_10897,N_8561,N_8344);
nand U10898 (N_10898,N_9698,N_8274);
and U10899 (N_10899,N_8323,N_9818);
xnor U10900 (N_10900,N_8602,N_8322);
and U10901 (N_10901,N_9964,N_9897);
or U10902 (N_10902,N_9837,N_9450);
or U10903 (N_10903,N_8846,N_8657);
or U10904 (N_10904,N_8928,N_8258);
and U10905 (N_10905,N_9649,N_9041);
or U10906 (N_10906,N_8267,N_8465);
xor U10907 (N_10907,N_9357,N_8597);
nand U10908 (N_10908,N_9322,N_9999);
nor U10909 (N_10909,N_8377,N_9532);
and U10910 (N_10910,N_9522,N_8171);
xor U10911 (N_10911,N_9296,N_8176);
or U10912 (N_10912,N_9934,N_8822);
nor U10913 (N_10913,N_9333,N_9027);
and U10914 (N_10914,N_8156,N_8295);
or U10915 (N_10915,N_8035,N_8689);
and U10916 (N_10916,N_8497,N_9309);
or U10917 (N_10917,N_8099,N_8858);
or U10918 (N_10918,N_8430,N_9132);
nand U10919 (N_10919,N_8227,N_9757);
nor U10920 (N_10920,N_9630,N_8796);
xor U10921 (N_10921,N_9382,N_8679);
nor U10922 (N_10922,N_9799,N_9703);
nor U10923 (N_10923,N_8823,N_8765);
nor U10924 (N_10924,N_8835,N_8859);
nor U10925 (N_10925,N_9219,N_8269);
nor U10926 (N_10926,N_8517,N_8309);
or U10927 (N_10927,N_9352,N_8880);
and U10928 (N_10928,N_8692,N_9945);
or U10929 (N_10929,N_8756,N_9014);
or U10930 (N_10930,N_8491,N_9174);
or U10931 (N_10931,N_9306,N_8826);
or U10932 (N_10932,N_8841,N_9068);
or U10933 (N_10933,N_9540,N_9736);
and U10934 (N_10934,N_8860,N_9501);
nor U10935 (N_10935,N_8867,N_8748);
xnor U10936 (N_10936,N_9926,N_9187);
and U10937 (N_10937,N_9429,N_9459);
nor U10938 (N_10938,N_9893,N_9451);
xor U10939 (N_10939,N_9638,N_9578);
xnor U10940 (N_10940,N_9213,N_9804);
xnor U10941 (N_10941,N_9468,N_9542);
nor U10942 (N_10942,N_9205,N_8842);
nand U10943 (N_10943,N_8676,N_8508);
nand U10944 (N_10944,N_8146,N_8442);
xnor U10945 (N_10945,N_9650,N_8214);
nor U10946 (N_10946,N_9892,N_9854);
nand U10947 (N_10947,N_9853,N_9040);
nand U10948 (N_10948,N_8317,N_9937);
nor U10949 (N_10949,N_9739,N_8116);
nand U10950 (N_10950,N_8094,N_8395);
xor U10951 (N_10951,N_8041,N_8458);
and U10952 (N_10952,N_8447,N_9619);
nor U10953 (N_10953,N_8996,N_9708);
and U10954 (N_10954,N_9321,N_8769);
or U10955 (N_10955,N_8033,N_9705);
or U10956 (N_10956,N_8981,N_9523);
and U10957 (N_10957,N_8687,N_8145);
xor U10958 (N_10958,N_9809,N_8591);
or U10959 (N_10959,N_9006,N_8745);
nand U10960 (N_10960,N_9927,N_8411);
and U10961 (N_10961,N_8729,N_9164);
or U10962 (N_10962,N_9097,N_9714);
nand U10963 (N_10963,N_9371,N_9001);
xnor U10964 (N_10964,N_9098,N_8944);
or U10965 (N_10965,N_9856,N_8209);
and U10966 (N_10966,N_8807,N_9725);
and U10967 (N_10967,N_8556,N_8153);
nor U10968 (N_10968,N_8120,N_9355);
xnor U10969 (N_10969,N_8079,N_9254);
nand U10970 (N_10970,N_9004,N_9692);
xor U10971 (N_10971,N_9572,N_8531);
nor U10972 (N_10972,N_9257,N_8742);
or U10973 (N_10973,N_8360,N_9029);
or U10974 (N_10974,N_8818,N_8118);
nor U10975 (N_10975,N_9919,N_9421);
nor U10976 (N_10976,N_8539,N_8368);
and U10977 (N_10977,N_9846,N_8717);
xor U10978 (N_10978,N_9276,N_8734);
nand U10979 (N_10979,N_9639,N_8677);
and U10980 (N_10980,N_8109,N_8820);
xnor U10981 (N_10981,N_9032,N_9568);
or U10982 (N_10982,N_8744,N_9062);
or U10983 (N_10983,N_9203,N_9397);
and U10984 (N_10984,N_9710,N_9784);
nor U10985 (N_10985,N_9002,N_8318);
and U10986 (N_10986,N_9643,N_9617);
or U10987 (N_10987,N_8975,N_9699);
nand U10988 (N_10988,N_8054,N_8421);
or U10989 (N_10989,N_9079,N_8157);
nor U10990 (N_10990,N_9622,N_8401);
and U10991 (N_10991,N_8618,N_9596);
and U10992 (N_10992,N_8141,N_8516);
nor U10993 (N_10993,N_8696,N_8456);
xor U10994 (N_10994,N_9887,N_9590);
nand U10995 (N_10995,N_9668,N_8193);
and U10996 (N_10996,N_9141,N_9658);
xor U10997 (N_10997,N_9392,N_9844);
xor U10998 (N_10998,N_9363,N_9016);
nor U10999 (N_10999,N_8433,N_9573);
xnor U11000 (N_11000,N_8442,N_9784);
nand U11001 (N_11001,N_8416,N_8449);
and U11002 (N_11002,N_8696,N_8822);
nor U11003 (N_11003,N_8576,N_8930);
or U11004 (N_11004,N_8880,N_8851);
or U11005 (N_11005,N_8061,N_9878);
nor U11006 (N_11006,N_9967,N_9966);
and U11007 (N_11007,N_8798,N_9779);
nand U11008 (N_11008,N_9462,N_8207);
or U11009 (N_11009,N_8693,N_8651);
or U11010 (N_11010,N_8559,N_8067);
xor U11011 (N_11011,N_9378,N_9764);
or U11012 (N_11012,N_8031,N_8990);
nand U11013 (N_11013,N_9918,N_8126);
nor U11014 (N_11014,N_8534,N_9686);
nor U11015 (N_11015,N_9865,N_9851);
and U11016 (N_11016,N_9135,N_9532);
or U11017 (N_11017,N_8646,N_9743);
or U11018 (N_11018,N_8415,N_9976);
nor U11019 (N_11019,N_8062,N_8750);
and U11020 (N_11020,N_9223,N_9989);
and U11021 (N_11021,N_8575,N_8247);
or U11022 (N_11022,N_8328,N_9857);
nand U11023 (N_11023,N_9372,N_9503);
xnor U11024 (N_11024,N_9873,N_8669);
nand U11025 (N_11025,N_9523,N_8480);
nor U11026 (N_11026,N_8660,N_9670);
xnor U11027 (N_11027,N_9951,N_9818);
xnor U11028 (N_11028,N_8557,N_8369);
or U11029 (N_11029,N_9699,N_9441);
nor U11030 (N_11030,N_9928,N_8639);
and U11031 (N_11031,N_8546,N_8541);
nand U11032 (N_11032,N_9898,N_8077);
nand U11033 (N_11033,N_9400,N_8265);
xor U11034 (N_11034,N_9167,N_8680);
and U11035 (N_11035,N_9657,N_9972);
nor U11036 (N_11036,N_8973,N_8091);
nor U11037 (N_11037,N_9096,N_8901);
or U11038 (N_11038,N_8201,N_9298);
or U11039 (N_11039,N_9654,N_8889);
nand U11040 (N_11040,N_9029,N_8480);
or U11041 (N_11041,N_8051,N_9760);
nor U11042 (N_11042,N_9845,N_9272);
nand U11043 (N_11043,N_9041,N_8000);
nor U11044 (N_11044,N_9815,N_8202);
nor U11045 (N_11045,N_8780,N_8966);
or U11046 (N_11046,N_8233,N_9813);
xor U11047 (N_11047,N_9841,N_9155);
xnor U11048 (N_11048,N_8886,N_8182);
nand U11049 (N_11049,N_9996,N_8703);
or U11050 (N_11050,N_9871,N_9752);
or U11051 (N_11051,N_9529,N_8365);
or U11052 (N_11052,N_8812,N_9315);
and U11053 (N_11053,N_9200,N_8043);
or U11054 (N_11054,N_8384,N_9212);
xor U11055 (N_11055,N_9795,N_8197);
nand U11056 (N_11056,N_9957,N_9888);
xnor U11057 (N_11057,N_9893,N_8139);
or U11058 (N_11058,N_8795,N_9815);
or U11059 (N_11059,N_8825,N_8834);
and U11060 (N_11060,N_9438,N_9028);
nand U11061 (N_11061,N_8893,N_8978);
nor U11062 (N_11062,N_8350,N_9909);
or U11063 (N_11063,N_8825,N_9766);
xnor U11064 (N_11064,N_9168,N_8770);
nor U11065 (N_11065,N_9294,N_9700);
nor U11066 (N_11066,N_9284,N_9365);
xnor U11067 (N_11067,N_8822,N_8037);
nand U11068 (N_11068,N_9977,N_8259);
nand U11069 (N_11069,N_9931,N_8333);
nor U11070 (N_11070,N_9590,N_9603);
or U11071 (N_11071,N_9806,N_8370);
nor U11072 (N_11072,N_9241,N_8516);
nand U11073 (N_11073,N_8067,N_8534);
or U11074 (N_11074,N_8274,N_9441);
nand U11075 (N_11075,N_8399,N_8050);
nand U11076 (N_11076,N_8020,N_8310);
nand U11077 (N_11077,N_9480,N_8944);
or U11078 (N_11078,N_9920,N_8833);
nor U11079 (N_11079,N_8739,N_8407);
or U11080 (N_11080,N_8755,N_8342);
xor U11081 (N_11081,N_8591,N_9882);
nor U11082 (N_11082,N_9595,N_9600);
nor U11083 (N_11083,N_9653,N_8529);
nand U11084 (N_11084,N_9681,N_9656);
nor U11085 (N_11085,N_8181,N_9381);
and U11086 (N_11086,N_8227,N_9687);
xor U11087 (N_11087,N_8283,N_9277);
nor U11088 (N_11088,N_9679,N_9990);
or U11089 (N_11089,N_8322,N_8567);
nor U11090 (N_11090,N_9597,N_9063);
nor U11091 (N_11091,N_9473,N_9543);
or U11092 (N_11092,N_8347,N_9260);
or U11093 (N_11093,N_9850,N_8960);
nand U11094 (N_11094,N_9673,N_9656);
and U11095 (N_11095,N_9103,N_9636);
nand U11096 (N_11096,N_9423,N_9384);
or U11097 (N_11097,N_9914,N_9582);
and U11098 (N_11098,N_8142,N_9351);
and U11099 (N_11099,N_9186,N_8275);
nand U11100 (N_11100,N_8499,N_9919);
nand U11101 (N_11101,N_8701,N_8635);
nand U11102 (N_11102,N_9175,N_9195);
xor U11103 (N_11103,N_9151,N_9580);
nand U11104 (N_11104,N_9727,N_9566);
xor U11105 (N_11105,N_8824,N_9013);
or U11106 (N_11106,N_8796,N_9660);
xor U11107 (N_11107,N_9666,N_9121);
nand U11108 (N_11108,N_8561,N_8894);
xor U11109 (N_11109,N_8397,N_8218);
or U11110 (N_11110,N_8685,N_9557);
nand U11111 (N_11111,N_9445,N_9901);
nand U11112 (N_11112,N_9595,N_9365);
and U11113 (N_11113,N_8477,N_8866);
or U11114 (N_11114,N_9375,N_8718);
and U11115 (N_11115,N_9581,N_8918);
xor U11116 (N_11116,N_8527,N_9142);
and U11117 (N_11117,N_9754,N_9013);
nor U11118 (N_11118,N_9574,N_9699);
nor U11119 (N_11119,N_8463,N_8906);
and U11120 (N_11120,N_8240,N_8867);
nand U11121 (N_11121,N_8916,N_9485);
and U11122 (N_11122,N_8763,N_9307);
nor U11123 (N_11123,N_8799,N_9374);
nand U11124 (N_11124,N_8421,N_9874);
or U11125 (N_11125,N_9854,N_9427);
nor U11126 (N_11126,N_8177,N_9715);
and U11127 (N_11127,N_9619,N_9512);
xor U11128 (N_11128,N_9085,N_9494);
xor U11129 (N_11129,N_8536,N_8274);
nor U11130 (N_11130,N_8896,N_9026);
or U11131 (N_11131,N_8424,N_9951);
xnor U11132 (N_11132,N_9722,N_9305);
nor U11133 (N_11133,N_8959,N_9695);
xor U11134 (N_11134,N_9447,N_8897);
and U11135 (N_11135,N_9274,N_9121);
and U11136 (N_11136,N_9282,N_8399);
nor U11137 (N_11137,N_8779,N_9092);
nand U11138 (N_11138,N_9712,N_8055);
nand U11139 (N_11139,N_9265,N_8926);
nor U11140 (N_11140,N_9019,N_8159);
xor U11141 (N_11141,N_8776,N_9843);
and U11142 (N_11142,N_8032,N_8645);
xor U11143 (N_11143,N_9720,N_9144);
xor U11144 (N_11144,N_9338,N_9989);
xnor U11145 (N_11145,N_8831,N_8640);
xor U11146 (N_11146,N_9938,N_8459);
nor U11147 (N_11147,N_9290,N_8714);
xnor U11148 (N_11148,N_8958,N_9723);
nand U11149 (N_11149,N_9727,N_8565);
or U11150 (N_11150,N_9064,N_9508);
nor U11151 (N_11151,N_8821,N_8878);
nor U11152 (N_11152,N_9061,N_9999);
xnor U11153 (N_11153,N_9654,N_8292);
or U11154 (N_11154,N_8262,N_9977);
xnor U11155 (N_11155,N_9997,N_8934);
xor U11156 (N_11156,N_9488,N_8971);
nor U11157 (N_11157,N_9357,N_9338);
or U11158 (N_11158,N_9416,N_9630);
nand U11159 (N_11159,N_9422,N_9559);
nand U11160 (N_11160,N_9961,N_9661);
or U11161 (N_11161,N_8836,N_9123);
nand U11162 (N_11162,N_9133,N_8876);
xor U11163 (N_11163,N_8684,N_8090);
xor U11164 (N_11164,N_9154,N_8237);
and U11165 (N_11165,N_9582,N_9540);
and U11166 (N_11166,N_8906,N_8031);
nand U11167 (N_11167,N_9509,N_9364);
nor U11168 (N_11168,N_9309,N_9793);
nand U11169 (N_11169,N_9011,N_9791);
and U11170 (N_11170,N_9517,N_8676);
or U11171 (N_11171,N_9930,N_9266);
or U11172 (N_11172,N_9757,N_8349);
xor U11173 (N_11173,N_9281,N_9410);
nand U11174 (N_11174,N_8312,N_8475);
nor U11175 (N_11175,N_9796,N_8055);
or U11176 (N_11176,N_9736,N_8755);
xor U11177 (N_11177,N_9778,N_8767);
and U11178 (N_11178,N_8555,N_9337);
nor U11179 (N_11179,N_8785,N_9203);
xor U11180 (N_11180,N_8314,N_9711);
nand U11181 (N_11181,N_8006,N_8524);
xnor U11182 (N_11182,N_9189,N_9081);
nor U11183 (N_11183,N_8459,N_9791);
and U11184 (N_11184,N_9109,N_8280);
and U11185 (N_11185,N_8988,N_9698);
xnor U11186 (N_11186,N_9647,N_9825);
and U11187 (N_11187,N_8667,N_8630);
nand U11188 (N_11188,N_8766,N_8852);
xnor U11189 (N_11189,N_8476,N_8190);
xor U11190 (N_11190,N_9335,N_8603);
nor U11191 (N_11191,N_9472,N_9565);
or U11192 (N_11192,N_8294,N_8224);
nand U11193 (N_11193,N_8311,N_9527);
and U11194 (N_11194,N_8098,N_8293);
xor U11195 (N_11195,N_8700,N_8379);
xor U11196 (N_11196,N_8587,N_9619);
xor U11197 (N_11197,N_8004,N_8838);
xnor U11198 (N_11198,N_8668,N_8326);
nor U11199 (N_11199,N_9091,N_8989);
or U11200 (N_11200,N_9193,N_9386);
nand U11201 (N_11201,N_8855,N_8697);
or U11202 (N_11202,N_9063,N_9704);
and U11203 (N_11203,N_9367,N_8030);
or U11204 (N_11204,N_8665,N_8937);
nand U11205 (N_11205,N_9018,N_9361);
nor U11206 (N_11206,N_8948,N_9191);
xor U11207 (N_11207,N_8746,N_9557);
and U11208 (N_11208,N_9464,N_8501);
nor U11209 (N_11209,N_8269,N_8364);
xor U11210 (N_11210,N_9797,N_9602);
or U11211 (N_11211,N_8896,N_9944);
or U11212 (N_11212,N_8247,N_9681);
nand U11213 (N_11213,N_8736,N_8692);
nand U11214 (N_11214,N_9703,N_8268);
xnor U11215 (N_11215,N_8115,N_9040);
nand U11216 (N_11216,N_8000,N_9240);
xor U11217 (N_11217,N_8912,N_9343);
nand U11218 (N_11218,N_9903,N_9369);
or U11219 (N_11219,N_9906,N_8451);
or U11220 (N_11220,N_9498,N_9639);
xor U11221 (N_11221,N_9887,N_8857);
nand U11222 (N_11222,N_8710,N_8096);
and U11223 (N_11223,N_9357,N_9810);
xnor U11224 (N_11224,N_8116,N_8708);
xnor U11225 (N_11225,N_8011,N_8029);
xnor U11226 (N_11226,N_9233,N_9804);
xor U11227 (N_11227,N_9454,N_9286);
or U11228 (N_11228,N_9071,N_9834);
and U11229 (N_11229,N_8304,N_8964);
nor U11230 (N_11230,N_9671,N_9474);
nand U11231 (N_11231,N_8437,N_9080);
nand U11232 (N_11232,N_9899,N_9441);
nand U11233 (N_11233,N_9186,N_9152);
and U11234 (N_11234,N_8698,N_9965);
xor U11235 (N_11235,N_8504,N_8196);
and U11236 (N_11236,N_9228,N_9689);
and U11237 (N_11237,N_9339,N_9247);
nor U11238 (N_11238,N_9655,N_9858);
or U11239 (N_11239,N_8115,N_9699);
nand U11240 (N_11240,N_9457,N_8158);
or U11241 (N_11241,N_9881,N_8514);
or U11242 (N_11242,N_9643,N_8053);
and U11243 (N_11243,N_9444,N_9516);
xor U11244 (N_11244,N_9709,N_8233);
and U11245 (N_11245,N_8929,N_9111);
or U11246 (N_11246,N_8626,N_8884);
and U11247 (N_11247,N_9934,N_9169);
and U11248 (N_11248,N_8500,N_8511);
nand U11249 (N_11249,N_8964,N_9538);
nor U11250 (N_11250,N_8134,N_9546);
nand U11251 (N_11251,N_9204,N_8609);
nor U11252 (N_11252,N_8779,N_8218);
xnor U11253 (N_11253,N_8137,N_9010);
nand U11254 (N_11254,N_9195,N_8375);
nand U11255 (N_11255,N_8479,N_8822);
nand U11256 (N_11256,N_8464,N_9765);
nor U11257 (N_11257,N_8193,N_9140);
and U11258 (N_11258,N_8500,N_8802);
nor U11259 (N_11259,N_9851,N_8541);
nand U11260 (N_11260,N_8440,N_9753);
nand U11261 (N_11261,N_9733,N_8553);
nand U11262 (N_11262,N_9049,N_9186);
or U11263 (N_11263,N_9767,N_8172);
nand U11264 (N_11264,N_9076,N_9242);
nor U11265 (N_11265,N_8419,N_9117);
or U11266 (N_11266,N_9718,N_9096);
nor U11267 (N_11267,N_9648,N_8857);
and U11268 (N_11268,N_8144,N_8710);
or U11269 (N_11269,N_9501,N_8133);
nor U11270 (N_11270,N_9600,N_8078);
and U11271 (N_11271,N_8470,N_9549);
nand U11272 (N_11272,N_9995,N_9154);
and U11273 (N_11273,N_9943,N_8954);
nand U11274 (N_11274,N_9309,N_9508);
nand U11275 (N_11275,N_8529,N_9905);
and U11276 (N_11276,N_9951,N_9222);
and U11277 (N_11277,N_8223,N_9714);
nor U11278 (N_11278,N_9674,N_8820);
nor U11279 (N_11279,N_9212,N_9038);
and U11280 (N_11280,N_8202,N_9936);
or U11281 (N_11281,N_9859,N_9546);
nor U11282 (N_11282,N_8618,N_8318);
or U11283 (N_11283,N_9478,N_9647);
xor U11284 (N_11284,N_8137,N_9816);
and U11285 (N_11285,N_9002,N_8860);
and U11286 (N_11286,N_8834,N_9267);
nand U11287 (N_11287,N_8063,N_9451);
nand U11288 (N_11288,N_8568,N_8645);
nand U11289 (N_11289,N_9827,N_8724);
and U11290 (N_11290,N_9745,N_9466);
nand U11291 (N_11291,N_9204,N_8607);
nand U11292 (N_11292,N_9141,N_9307);
and U11293 (N_11293,N_9344,N_9340);
nand U11294 (N_11294,N_9884,N_8692);
and U11295 (N_11295,N_8055,N_9106);
nand U11296 (N_11296,N_9956,N_8963);
and U11297 (N_11297,N_8950,N_9857);
xor U11298 (N_11298,N_8670,N_9820);
xor U11299 (N_11299,N_9457,N_9950);
and U11300 (N_11300,N_8207,N_8340);
and U11301 (N_11301,N_9352,N_9723);
xor U11302 (N_11302,N_8010,N_8506);
nand U11303 (N_11303,N_8677,N_8012);
xor U11304 (N_11304,N_8559,N_8786);
xor U11305 (N_11305,N_8856,N_8297);
or U11306 (N_11306,N_9961,N_9276);
xor U11307 (N_11307,N_8484,N_9524);
nor U11308 (N_11308,N_8192,N_9052);
or U11309 (N_11309,N_8834,N_9091);
nand U11310 (N_11310,N_9404,N_9282);
and U11311 (N_11311,N_8901,N_9974);
nor U11312 (N_11312,N_9521,N_9007);
xnor U11313 (N_11313,N_8519,N_8745);
nor U11314 (N_11314,N_9894,N_8474);
or U11315 (N_11315,N_8694,N_9671);
nand U11316 (N_11316,N_9250,N_8069);
xnor U11317 (N_11317,N_9567,N_8555);
and U11318 (N_11318,N_8744,N_8479);
or U11319 (N_11319,N_9543,N_8497);
nor U11320 (N_11320,N_9397,N_8396);
xnor U11321 (N_11321,N_9569,N_8309);
or U11322 (N_11322,N_9101,N_9670);
nor U11323 (N_11323,N_8984,N_8176);
nor U11324 (N_11324,N_9017,N_9241);
nor U11325 (N_11325,N_8979,N_8216);
or U11326 (N_11326,N_9488,N_9710);
xor U11327 (N_11327,N_9517,N_9795);
xor U11328 (N_11328,N_9176,N_8297);
and U11329 (N_11329,N_8202,N_9510);
nand U11330 (N_11330,N_8723,N_8518);
or U11331 (N_11331,N_9990,N_9282);
nor U11332 (N_11332,N_8136,N_9342);
and U11333 (N_11333,N_8605,N_9973);
nand U11334 (N_11334,N_8334,N_9552);
xnor U11335 (N_11335,N_8744,N_8049);
nor U11336 (N_11336,N_9894,N_9889);
nor U11337 (N_11337,N_9365,N_9148);
nor U11338 (N_11338,N_9151,N_9376);
nor U11339 (N_11339,N_8781,N_8626);
nor U11340 (N_11340,N_9271,N_8585);
nand U11341 (N_11341,N_9473,N_9076);
nand U11342 (N_11342,N_8345,N_9704);
or U11343 (N_11343,N_8872,N_8645);
nand U11344 (N_11344,N_9714,N_8848);
and U11345 (N_11345,N_8691,N_9837);
nor U11346 (N_11346,N_8937,N_9551);
and U11347 (N_11347,N_8332,N_8251);
or U11348 (N_11348,N_8125,N_8313);
and U11349 (N_11349,N_8882,N_8887);
nor U11350 (N_11350,N_8099,N_8669);
or U11351 (N_11351,N_8819,N_9899);
or U11352 (N_11352,N_9727,N_9461);
xor U11353 (N_11353,N_8961,N_9116);
nor U11354 (N_11354,N_9591,N_8189);
nand U11355 (N_11355,N_9185,N_8615);
nand U11356 (N_11356,N_9506,N_9675);
nand U11357 (N_11357,N_9359,N_9968);
xnor U11358 (N_11358,N_9587,N_8110);
or U11359 (N_11359,N_8199,N_9668);
or U11360 (N_11360,N_9748,N_9579);
nand U11361 (N_11361,N_8290,N_8887);
or U11362 (N_11362,N_9232,N_9408);
and U11363 (N_11363,N_8718,N_8110);
xor U11364 (N_11364,N_9141,N_9065);
nand U11365 (N_11365,N_8023,N_8248);
xor U11366 (N_11366,N_8269,N_9522);
xor U11367 (N_11367,N_9511,N_8303);
or U11368 (N_11368,N_9262,N_9827);
or U11369 (N_11369,N_8257,N_9723);
nand U11370 (N_11370,N_8723,N_9325);
nor U11371 (N_11371,N_8000,N_8033);
nor U11372 (N_11372,N_8588,N_9086);
or U11373 (N_11373,N_9839,N_8931);
xnor U11374 (N_11374,N_9238,N_9681);
nand U11375 (N_11375,N_9368,N_8555);
and U11376 (N_11376,N_9145,N_9833);
nor U11377 (N_11377,N_9659,N_8817);
nand U11378 (N_11378,N_9187,N_9534);
nor U11379 (N_11379,N_8513,N_8241);
and U11380 (N_11380,N_9735,N_9395);
nand U11381 (N_11381,N_9991,N_9725);
xor U11382 (N_11382,N_9264,N_8969);
and U11383 (N_11383,N_9436,N_8403);
and U11384 (N_11384,N_8351,N_8035);
nand U11385 (N_11385,N_8176,N_8680);
nor U11386 (N_11386,N_9916,N_8084);
nor U11387 (N_11387,N_9034,N_9144);
nand U11388 (N_11388,N_9044,N_8119);
nand U11389 (N_11389,N_8419,N_8947);
xor U11390 (N_11390,N_9461,N_8153);
and U11391 (N_11391,N_9645,N_9803);
and U11392 (N_11392,N_8191,N_8609);
nor U11393 (N_11393,N_8967,N_9962);
or U11394 (N_11394,N_9936,N_9540);
nand U11395 (N_11395,N_8725,N_9079);
nand U11396 (N_11396,N_8785,N_9811);
nor U11397 (N_11397,N_9475,N_8653);
xor U11398 (N_11398,N_8188,N_9090);
nand U11399 (N_11399,N_9761,N_9814);
and U11400 (N_11400,N_9370,N_9984);
xnor U11401 (N_11401,N_9370,N_8999);
or U11402 (N_11402,N_9950,N_8610);
nor U11403 (N_11403,N_9064,N_9167);
nand U11404 (N_11404,N_9180,N_8988);
nand U11405 (N_11405,N_9162,N_9726);
nor U11406 (N_11406,N_9783,N_9852);
nand U11407 (N_11407,N_8524,N_9818);
nand U11408 (N_11408,N_8224,N_8223);
or U11409 (N_11409,N_8592,N_8923);
xnor U11410 (N_11410,N_8481,N_9730);
or U11411 (N_11411,N_9134,N_9932);
or U11412 (N_11412,N_8790,N_9138);
or U11413 (N_11413,N_9270,N_8050);
nor U11414 (N_11414,N_9264,N_8357);
nand U11415 (N_11415,N_9326,N_9855);
xnor U11416 (N_11416,N_8063,N_8020);
xnor U11417 (N_11417,N_9103,N_8452);
xor U11418 (N_11418,N_8201,N_8408);
nor U11419 (N_11419,N_9929,N_8880);
xnor U11420 (N_11420,N_8671,N_9770);
or U11421 (N_11421,N_9105,N_9589);
xor U11422 (N_11422,N_9675,N_9046);
or U11423 (N_11423,N_8620,N_9754);
xor U11424 (N_11424,N_9443,N_8135);
xor U11425 (N_11425,N_9912,N_8073);
nor U11426 (N_11426,N_8557,N_9976);
and U11427 (N_11427,N_8111,N_9061);
nor U11428 (N_11428,N_8128,N_9882);
nor U11429 (N_11429,N_9398,N_9114);
xnor U11430 (N_11430,N_9713,N_8147);
nor U11431 (N_11431,N_8123,N_9166);
nand U11432 (N_11432,N_8215,N_9336);
nor U11433 (N_11433,N_8131,N_9076);
nand U11434 (N_11434,N_9878,N_9710);
or U11435 (N_11435,N_8869,N_9677);
and U11436 (N_11436,N_8708,N_8256);
xnor U11437 (N_11437,N_8237,N_9041);
xnor U11438 (N_11438,N_9679,N_9868);
or U11439 (N_11439,N_9510,N_9770);
and U11440 (N_11440,N_8628,N_9847);
and U11441 (N_11441,N_9755,N_9058);
and U11442 (N_11442,N_8989,N_9246);
nor U11443 (N_11443,N_9245,N_9426);
and U11444 (N_11444,N_8893,N_9581);
nand U11445 (N_11445,N_9749,N_9487);
and U11446 (N_11446,N_8312,N_8710);
xnor U11447 (N_11447,N_8358,N_8350);
nand U11448 (N_11448,N_9589,N_9358);
or U11449 (N_11449,N_8999,N_8424);
xnor U11450 (N_11450,N_9836,N_9198);
nor U11451 (N_11451,N_8385,N_8529);
or U11452 (N_11452,N_8576,N_9129);
xor U11453 (N_11453,N_8003,N_9985);
xnor U11454 (N_11454,N_9858,N_9835);
and U11455 (N_11455,N_8735,N_9579);
nand U11456 (N_11456,N_8944,N_9173);
nor U11457 (N_11457,N_9166,N_8740);
nand U11458 (N_11458,N_8108,N_9748);
and U11459 (N_11459,N_9229,N_8750);
and U11460 (N_11460,N_9938,N_9998);
nand U11461 (N_11461,N_9760,N_9989);
or U11462 (N_11462,N_8737,N_8075);
nand U11463 (N_11463,N_8908,N_9593);
xnor U11464 (N_11464,N_9291,N_8731);
and U11465 (N_11465,N_9735,N_8246);
nand U11466 (N_11466,N_9912,N_8036);
nand U11467 (N_11467,N_9072,N_9185);
nand U11468 (N_11468,N_8575,N_8310);
and U11469 (N_11469,N_9058,N_8741);
xor U11470 (N_11470,N_9909,N_8490);
nor U11471 (N_11471,N_9602,N_9869);
and U11472 (N_11472,N_9772,N_8901);
or U11473 (N_11473,N_8615,N_8825);
nand U11474 (N_11474,N_9072,N_9611);
or U11475 (N_11475,N_8044,N_9748);
xnor U11476 (N_11476,N_9102,N_8088);
and U11477 (N_11477,N_9383,N_9358);
nand U11478 (N_11478,N_8105,N_8461);
and U11479 (N_11479,N_9684,N_8190);
nor U11480 (N_11480,N_8472,N_9993);
nand U11481 (N_11481,N_9321,N_9930);
nand U11482 (N_11482,N_9998,N_8455);
and U11483 (N_11483,N_8058,N_8076);
and U11484 (N_11484,N_9463,N_8760);
or U11485 (N_11485,N_9573,N_8816);
and U11486 (N_11486,N_9305,N_9974);
or U11487 (N_11487,N_9469,N_8245);
or U11488 (N_11488,N_8125,N_9539);
and U11489 (N_11489,N_8741,N_9297);
xor U11490 (N_11490,N_8306,N_8879);
and U11491 (N_11491,N_9482,N_8846);
nand U11492 (N_11492,N_9097,N_8933);
xor U11493 (N_11493,N_9350,N_9275);
xnor U11494 (N_11494,N_8239,N_9894);
xor U11495 (N_11495,N_8594,N_9541);
and U11496 (N_11496,N_8530,N_9591);
and U11497 (N_11497,N_9579,N_8211);
and U11498 (N_11498,N_9220,N_8683);
and U11499 (N_11499,N_8643,N_9201);
and U11500 (N_11500,N_8643,N_9287);
and U11501 (N_11501,N_8042,N_8812);
or U11502 (N_11502,N_8368,N_9490);
xnor U11503 (N_11503,N_9629,N_9331);
or U11504 (N_11504,N_8171,N_8580);
nand U11505 (N_11505,N_8497,N_8880);
xor U11506 (N_11506,N_8339,N_9759);
or U11507 (N_11507,N_9952,N_8143);
nor U11508 (N_11508,N_8519,N_8268);
nand U11509 (N_11509,N_8583,N_8736);
nand U11510 (N_11510,N_8548,N_9833);
nand U11511 (N_11511,N_8108,N_8717);
or U11512 (N_11512,N_9281,N_8037);
nor U11513 (N_11513,N_8513,N_9302);
and U11514 (N_11514,N_8756,N_8848);
and U11515 (N_11515,N_8491,N_8634);
nand U11516 (N_11516,N_9135,N_8475);
xnor U11517 (N_11517,N_9334,N_9747);
or U11518 (N_11518,N_9107,N_9328);
xnor U11519 (N_11519,N_8390,N_9556);
nor U11520 (N_11520,N_8112,N_8454);
xnor U11521 (N_11521,N_9730,N_9935);
and U11522 (N_11522,N_8008,N_9197);
nor U11523 (N_11523,N_9975,N_8219);
and U11524 (N_11524,N_8482,N_9258);
or U11525 (N_11525,N_8396,N_9920);
nand U11526 (N_11526,N_8251,N_9991);
or U11527 (N_11527,N_8421,N_9571);
and U11528 (N_11528,N_8183,N_8439);
or U11529 (N_11529,N_8872,N_9425);
or U11530 (N_11530,N_9086,N_9124);
nand U11531 (N_11531,N_9004,N_9295);
and U11532 (N_11532,N_9511,N_9734);
xor U11533 (N_11533,N_8096,N_9953);
nor U11534 (N_11534,N_9367,N_9007);
and U11535 (N_11535,N_8412,N_9708);
xnor U11536 (N_11536,N_9455,N_8374);
or U11537 (N_11537,N_8793,N_8423);
nor U11538 (N_11538,N_9946,N_9532);
or U11539 (N_11539,N_9043,N_9870);
xor U11540 (N_11540,N_9471,N_8579);
nor U11541 (N_11541,N_8748,N_8029);
nor U11542 (N_11542,N_8340,N_9752);
xnor U11543 (N_11543,N_9022,N_9716);
nand U11544 (N_11544,N_8134,N_9579);
xor U11545 (N_11545,N_9410,N_9077);
or U11546 (N_11546,N_8693,N_8331);
xnor U11547 (N_11547,N_9141,N_8620);
or U11548 (N_11548,N_8209,N_9683);
or U11549 (N_11549,N_9923,N_9021);
nand U11550 (N_11550,N_8808,N_9596);
or U11551 (N_11551,N_8159,N_9272);
nor U11552 (N_11552,N_8386,N_9712);
or U11553 (N_11553,N_9682,N_9615);
xor U11554 (N_11554,N_8326,N_9786);
xnor U11555 (N_11555,N_9452,N_8509);
nand U11556 (N_11556,N_9844,N_8258);
nor U11557 (N_11557,N_8379,N_9896);
and U11558 (N_11558,N_8191,N_9310);
nor U11559 (N_11559,N_9039,N_8015);
nand U11560 (N_11560,N_8260,N_8173);
or U11561 (N_11561,N_9496,N_8663);
or U11562 (N_11562,N_8368,N_9159);
nand U11563 (N_11563,N_9958,N_9562);
nand U11564 (N_11564,N_9125,N_8704);
xnor U11565 (N_11565,N_8215,N_9554);
xor U11566 (N_11566,N_8927,N_8512);
nor U11567 (N_11567,N_9687,N_9350);
nand U11568 (N_11568,N_9297,N_8894);
nand U11569 (N_11569,N_8866,N_8442);
or U11570 (N_11570,N_8463,N_9190);
nor U11571 (N_11571,N_9115,N_8549);
and U11572 (N_11572,N_8107,N_9176);
xnor U11573 (N_11573,N_9004,N_8513);
nor U11574 (N_11574,N_8992,N_9623);
nor U11575 (N_11575,N_8950,N_9936);
nor U11576 (N_11576,N_8363,N_8612);
nor U11577 (N_11577,N_9015,N_9734);
nand U11578 (N_11578,N_9794,N_8827);
and U11579 (N_11579,N_8241,N_9398);
nor U11580 (N_11580,N_9848,N_8926);
xor U11581 (N_11581,N_8787,N_8493);
or U11582 (N_11582,N_9092,N_9237);
and U11583 (N_11583,N_8965,N_9387);
nand U11584 (N_11584,N_8214,N_9894);
and U11585 (N_11585,N_9019,N_9687);
nand U11586 (N_11586,N_9783,N_9263);
xor U11587 (N_11587,N_8404,N_8751);
nand U11588 (N_11588,N_8455,N_8578);
xnor U11589 (N_11589,N_8199,N_9122);
nor U11590 (N_11590,N_9011,N_8198);
xnor U11591 (N_11591,N_9629,N_9113);
nor U11592 (N_11592,N_8231,N_8877);
xor U11593 (N_11593,N_8100,N_9240);
nor U11594 (N_11594,N_9663,N_8445);
nor U11595 (N_11595,N_9160,N_9584);
nand U11596 (N_11596,N_8885,N_9822);
and U11597 (N_11597,N_9760,N_8681);
xor U11598 (N_11598,N_8567,N_8949);
nand U11599 (N_11599,N_9588,N_8856);
nand U11600 (N_11600,N_9380,N_8130);
or U11601 (N_11601,N_9573,N_9179);
and U11602 (N_11602,N_8623,N_9350);
or U11603 (N_11603,N_9060,N_8048);
nor U11604 (N_11604,N_8050,N_8012);
nand U11605 (N_11605,N_9234,N_8676);
nor U11606 (N_11606,N_8277,N_9083);
xor U11607 (N_11607,N_8198,N_9099);
nor U11608 (N_11608,N_9477,N_9854);
xnor U11609 (N_11609,N_8423,N_9505);
nand U11610 (N_11610,N_8121,N_9436);
nor U11611 (N_11611,N_8526,N_8756);
nor U11612 (N_11612,N_8383,N_8532);
nor U11613 (N_11613,N_9971,N_8820);
and U11614 (N_11614,N_9556,N_9479);
or U11615 (N_11615,N_9628,N_8287);
nand U11616 (N_11616,N_8890,N_9160);
nand U11617 (N_11617,N_9765,N_8760);
and U11618 (N_11618,N_8015,N_9243);
and U11619 (N_11619,N_9733,N_9601);
and U11620 (N_11620,N_9238,N_8459);
nor U11621 (N_11621,N_9310,N_9968);
nand U11622 (N_11622,N_8052,N_9205);
and U11623 (N_11623,N_9546,N_9048);
nor U11624 (N_11624,N_9603,N_9605);
nor U11625 (N_11625,N_8095,N_8775);
or U11626 (N_11626,N_8189,N_9065);
and U11627 (N_11627,N_9264,N_9017);
xnor U11628 (N_11628,N_8622,N_9534);
xnor U11629 (N_11629,N_9008,N_9189);
nand U11630 (N_11630,N_8635,N_8939);
nor U11631 (N_11631,N_8480,N_8889);
or U11632 (N_11632,N_9668,N_9039);
and U11633 (N_11633,N_9879,N_9871);
xnor U11634 (N_11634,N_8766,N_9229);
nand U11635 (N_11635,N_9296,N_8381);
nor U11636 (N_11636,N_8723,N_9681);
and U11637 (N_11637,N_9950,N_8549);
and U11638 (N_11638,N_9167,N_8218);
and U11639 (N_11639,N_8019,N_8033);
and U11640 (N_11640,N_8454,N_9938);
and U11641 (N_11641,N_9492,N_9305);
xor U11642 (N_11642,N_9152,N_9405);
xnor U11643 (N_11643,N_9942,N_9980);
nand U11644 (N_11644,N_9505,N_8416);
and U11645 (N_11645,N_8025,N_9548);
xor U11646 (N_11646,N_9528,N_8771);
xnor U11647 (N_11647,N_8419,N_8690);
nor U11648 (N_11648,N_8495,N_9628);
xnor U11649 (N_11649,N_8747,N_9570);
or U11650 (N_11650,N_9708,N_9435);
nand U11651 (N_11651,N_9018,N_9290);
and U11652 (N_11652,N_9428,N_9350);
nand U11653 (N_11653,N_9959,N_9137);
or U11654 (N_11654,N_8703,N_9206);
or U11655 (N_11655,N_8304,N_8708);
nand U11656 (N_11656,N_8996,N_9445);
nand U11657 (N_11657,N_9897,N_8942);
nor U11658 (N_11658,N_8781,N_8127);
xor U11659 (N_11659,N_9030,N_9332);
or U11660 (N_11660,N_9941,N_9831);
and U11661 (N_11661,N_9888,N_8183);
nor U11662 (N_11662,N_9067,N_8926);
nor U11663 (N_11663,N_9793,N_9301);
nand U11664 (N_11664,N_8151,N_9483);
or U11665 (N_11665,N_9180,N_9887);
and U11666 (N_11666,N_9081,N_8350);
nor U11667 (N_11667,N_9186,N_8632);
nor U11668 (N_11668,N_9121,N_9155);
and U11669 (N_11669,N_9627,N_9334);
xnor U11670 (N_11670,N_8717,N_9808);
nor U11671 (N_11671,N_8527,N_8328);
nand U11672 (N_11672,N_9511,N_9311);
or U11673 (N_11673,N_8380,N_9370);
xor U11674 (N_11674,N_8248,N_8898);
or U11675 (N_11675,N_8443,N_8318);
nor U11676 (N_11676,N_9213,N_8322);
nor U11677 (N_11677,N_9092,N_8924);
and U11678 (N_11678,N_9489,N_9615);
xor U11679 (N_11679,N_8377,N_8026);
nand U11680 (N_11680,N_8988,N_9007);
nor U11681 (N_11681,N_8714,N_9719);
or U11682 (N_11682,N_8726,N_9916);
and U11683 (N_11683,N_9410,N_8997);
nand U11684 (N_11684,N_8740,N_9120);
nand U11685 (N_11685,N_9250,N_8795);
nor U11686 (N_11686,N_9245,N_8521);
and U11687 (N_11687,N_9761,N_9974);
nor U11688 (N_11688,N_8943,N_9267);
nand U11689 (N_11689,N_8514,N_9271);
xor U11690 (N_11690,N_9320,N_8969);
nor U11691 (N_11691,N_9019,N_9583);
xor U11692 (N_11692,N_8919,N_9721);
xor U11693 (N_11693,N_8159,N_9963);
or U11694 (N_11694,N_9722,N_8191);
xor U11695 (N_11695,N_8292,N_9799);
xnor U11696 (N_11696,N_9549,N_8406);
xnor U11697 (N_11697,N_9999,N_8484);
or U11698 (N_11698,N_9406,N_8961);
nand U11699 (N_11699,N_9229,N_9686);
nor U11700 (N_11700,N_8520,N_9406);
xnor U11701 (N_11701,N_8675,N_8384);
and U11702 (N_11702,N_8106,N_9494);
xor U11703 (N_11703,N_9768,N_9907);
or U11704 (N_11704,N_9376,N_9668);
nand U11705 (N_11705,N_8217,N_9573);
and U11706 (N_11706,N_9471,N_8958);
xor U11707 (N_11707,N_9976,N_8754);
nor U11708 (N_11708,N_8956,N_8574);
xnor U11709 (N_11709,N_8267,N_9348);
xor U11710 (N_11710,N_8320,N_8228);
xnor U11711 (N_11711,N_9312,N_9887);
nor U11712 (N_11712,N_9019,N_9295);
xor U11713 (N_11713,N_9081,N_9717);
xnor U11714 (N_11714,N_8443,N_9310);
xor U11715 (N_11715,N_9729,N_8441);
or U11716 (N_11716,N_9670,N_8832);
xnor U11717 (N_11717,N_9123,N_8019);
xnor U11718 (N_11718,N_8755,N_9623);
nand U11719 (N_11719,N_8160,N_8427);
nor U11720 (N_11720,N_9280,N_8391);
nor U11721 (N_11721,N_9439,N_9608);
and U11722 (N_11722,N_8682,N_8606);
or U11723 (N_11723,N_8750,N_9881);
xor U11724 (N_11724,N_8241,N_9293);
and U11725 (N_11725,N_8974,N_8833);
nand U11726 (N_11726,N_8255,N_8328);
nor U11727 (N_11727,N_9369,N_9010);
nor U11728 (N_11728,N_9536,N_9100);
or U11729 (N_11729,N_8601,N_9236);
nor U11730 (N_11730,N_8608,N_9927);
and U11731 (N_11731,N_8109,N_9507);
nor U11732 (N_11732,N_9836,N_9660);
nor U11733 (N_11733,N_9050,N_8938);
nand U11734 (N_11734,N_9065,N_8484);
or U11735 (N_11735,N_8535,N_8341);
xor U11736 (N_11736,N_9423,N_9600);
xnor U11737 (N_11737,N_8746,N_9837);
nand U11738 (N_11738,N_8953,N_8529);
nor U11739 (N_11739,N_9615,N_8378);
or U11740 (N_11740,N_9182,N_8626);
and U11741 (N_11741,N_9462,N_9146);
nor U11742 (N_11742,N_8092,N_8015);
nand U11743 (N_11743,N_9045,N_8835);
and U11744 (N_11744,N_8211,N_9842);
nor U11745 (N_11745,N_9023,N_9721);
nand U11746 (N_11746,N_8510,N_9674);
xnor U11747 (N_11747,N_9746,N_8121);
xnor U11748 (N_11748,N_8992,N_8605);
nand U11749 (N_11749,N_8154,N_9045);
xnor U11750 (N_11750,N_9092,N_8859);
xnor U11751 (N_11751,N_8519,N_9452);
xnor U11752 (N_11752,N_8569,N_8807);
nand U11753 (N_11753,N_8176,N_8872);
and U11754 (N_11754,N_9788,N_8990);
xnor U11755 (N_11755,N_8402,N_9221);
nand U11756 (N_11756,N_8892,N_9508);
nand U11757 (N_11757,N_8429,N_9572);
nand U11758 (N_11758,N_8619,N_8124);
xnor U11759 (N_11759,N_8454,N_8110);
and U11760 (N_11760,N_9621,N_8109);
and U11761 (N_11761,N_8640,N_8325);
or U11762 (N_11762,N_8030,N_9204);
or U11763 (N_11763,N_8341,N_8874);
nand U11764 (N_11764,N_8266,N_9817);
xnor U11765 (N_11765,N_8340,N_8357);
or U11766 (N_11766,N_9243,N_8410);
nand U11767 (N_11767,N_8099,N_9321);
and U11768 (N_11768,N_8973,N_8172);
or U11769 (N_11769,N_8368,N_8059);
and U11770 (N_11770,N_8362,N_8289);
nand U11771 (N_11771,N_9281,N_9665);
and U11772 (N_11772,N_9239,N_9195);
and U11773 (N_11773,N_9182,N_9834);
xor U11774 (N_11774,N_9748,N_9515);
nand U11775 (N_11775,N_9723,N_9557);
and U11776 (N_11776,N_8172,N_8785);
nand U11777 (N_11777,N_9988,N_8805);
nand U11778 (N_11778,N_9505,N_9143);
xnor U11779 (N_11779,N_9353,N_9297);
xor U11780 (N_11780,N_9874,N_8635);
or U11781 (N_11781,N_9576,N_8813);
nand U11782 (N_11782,N_9513,N_9571);
or U11783 (N_11783,N_8130,N_9383);
or U11784 (N_11784,N_9722,N_9757);
and U11785 (N_11785,N_9184,N_9371);
xor U11786 (N_11786,N_9277,N_8554);
nand U11787 (N_11787,N_9756,N_9245);
or U11788 (N_11788,N_8372,N_9949);
xnor U11789 (N_11789,N_9008,N_8356);
xnor U11790 (N_11790,N_8341,N_9831);
nor U11791 (N_11791,N_9089,N_9344);
or U11792 (N_11792,N_9094,N_8095);
or U11793 (N_11793,N_8235,N_8532);
or U11794 (N_11794,N_9126,N_9818);
and U11795 (N_11795,N_8121,N_9302);
xor U11796 (N_11796,N_8640,N_8476);
nand U11797 (N_11797,N_8475,N_8334);
nor U11798 (N_11798,N_9970,N_8482);
nand U11799 (N_11799,N_9377,N_8111);
or U11800 (N_11800,N_8984,N_8014);
nor U11801 (N_11801,N_8467,N_9271);
xnor U11802 (N_11802,N_8982,N_9854);
or U11803 (N_11803,N_9680,N_8820);
or U11804 (N_11804,N_9588,N_9158);
nand U11805 (N_11805,N_8366,N_9745);
and U11806 (N_11806,N_9803,N_9935);
or U11807 (N_11807,N_9491,N_9931);
or U11808 (N_11808,N_9507,N_8149);
xnor U11809 (N_11809,N_9728,N_8986);
and U11810 (N_11810,N_9163,N_9652);
xor U11811 (N_11811,N_8237,N_9004);
or U11812 (N_11812,N_8800,N_9982);
xnor U11813 (N_11813,N_8716,N_8465);
or U11814 (N_11814,N_9574,N_9263);
xor U11815 (N_11815,N_9571,N_8032);
nand U11816 (N_11816,N_8605,N_8157);
or U11817 (N_11817,N_9445,N_8498);
and U11818 (N_11818,N_9037,N_9433);
nor U11819 (N_11819,N_9465,N_8547);
and U11820 (N_11820,N_9286,N_8005);
xor U11821 (N_11821,N_8743,N_9793);
xnor U11822 (N_11822,N_8902,N_9828);
and U11823 (N_11823,N_8993,N_8361);
and U11824 (N_11824,N_8965,N_9955);
nor U11825 (N_11825,N_8097,N_8302);
nor U11826 (N_11826,N_8372,N_8395);
and U11827 (N_11827,N_9916,N_9788);
nor U11828 (N_11828,N_9243,N_8088);
xnor U11829 (N_11829,N_8262,N_9273);
or U11830 (N_11830,N_9755,N_9243);
nor U11831 (N_11831,N_8035,N_9895);
and U11832 (N_11832,N_8095,N_9748);
nand U11833 (N_11833,N_9700,N_9530);
and U11834 (N_11834,N_8094,N_8305);
nor U11835 (N_11835,N_9727,N_8451);
nand U11836 (N_11836,N_9550,N_8264);
or U11837 (N_11837,N_8187,N_9194);
nand U11838 (N_11838,N_9820,N_8665);
and U11839 (N_11839,N_9179,N_8507);
nand U11840 (N_11840,N_9831,N_8069);
xnor U11841 (N_11841,N_8803,N_9985);
xnor U11842 (N_11842,N_8593,N_9421);
xor U11843 (N_11843,N_9497,N_9981);
or U11844 (N_11844,N_9841,N_8846);
or U11845 (N_11845,N_9590,N_9672);
nor U11846 (N_11846,N_8915,N_8666);
xnor U11847 (N_11847,N_8657,N_8251);
or U11848 (N_11848,N_8444,N_8578);
nand U11849 (N_11849,N_8673,N_8486);
nand U11850 (N_11850,N_8128,N_9094);
nor U11851 (N_11851,N_8009,N_9325);
or U11852 (N_11852,N_9040,N_8278);
or U11853 (N_11853,N_8617,N_9419);
and U11854 (N_11854,N_8211,N_8088);
nor U11855 (N_11855,N_9416,N_8462);
xnor U11856 (N_11856,N_9696,N_8062);
nor U11857 (N_11857,N_8977,N_9963);
or U11858 (N_11858,N_9019,N_8526);
and U11859 (N_11859,N_8188,N_8533);
nand U11860 (N_11860,N_8194,N_9978);
nand U11861 (N_11861,N_9178,N_9186);
xnor U11862 (N_11862,N_9133,N_9371);
or U11863 (N_11863,N_8341,N_9083);
xnor U11864 (N_11864,N_9392,N_8498);
xor U11865 (N_11865,N_9336,N_8112);
xnor U11866 (N_11866,N_8424,N_8893);
nor U11867 (N_11867,N_8952,N_8323);
xnor U11868 (N_11868,N_8010,N_8041);
xnor U11869 (N_11869,N_9162,N_8443);
and U11870 (N_11870,N_9014,N_8458);
nor U11871 (N_11871,N_8749,N_8473);
nor U11872 (N_11872,N_8071,N_9927);
or U11873 (N_11873,N_9890,N_9374);
xor U11874 (N_11874,N_9327,N_9328);
or U11875 (N_11875,N_8145,N_8748);
and U11876 (N_11876,N_9088,N_8956);
nor U11877 (N_11877,N_9415,N_8252);
or U11878 (N_11878,N_9273,N_9470);
or U11879 (N_11879,N_9418,N_8278);
nor U11880 (N_11880,N_9721,N_9082);
nand U11881 (N_11881,N_8797,N_8068);
xnor U11882 (N_11882,N_8443,N_9582);
nor U11883 (N_11883,N_9969,N_9081);
or U11884 (N_11884,N_8487,N_8146);
or U11885 (N_11885,N_8136,N_8773);
nand U11886 (N_11886,N_9222,N_9576);
nand U11887 (N_11887,N_9682,N_9916);
nand U11888 (N_11888,N_8492,N_8221);
or U11889 (N_11889,N_8050,N_9910);
xor U11890 (N_11890,N_9440,N_9303);
nand U11891 (N_11891,N_9587,N_9262);
and U11892 (N_11892,N_8858,N_8544);
nand U11893 (N_11893,N_8938,N_8817);
xnor U11894 (N_11894,N_8150,N_8526);
and U11895 (N_11895,N_9691,N_9683);
nor U11896 (N_11896,N_8598,N_8007);
nor U11897 (N_11897,N_9013,N_8680);
xnor U11898 (N_11898,N_9616,N_9138);
xor U11899 (N_11899,N_9147,N_8142);
and U11900 (N_11900,N_8186,N_9070);
nor U11901 (N_11901,N_8801,N_8099);
xnor U11902 (N_11902,N_8867,N_8901);
nor U11903 (N_11903,N_8889,N_9003);
or U11904 (N_11904,N_9337,N_9422);
nand U11905 (N_11905,N_9810,N_8516);
or U11906 (N_11906,N_8185,N_8619);
and U11907 (N_11907,N_8569,N_9573);
and U11908 (N_11908,N_9465,N_8338);
and U11909 (N_11909,N_8681,N_9993);
and U11910 (N_11910,N_8869,N_9115);
or U11911 (N_11911,N_9881,N_9690);
xor U11912 (N_11912,N_8543,N_9591);
nor U11913 (N_11913,N_8373,N_8934);
and U11914 (N_11914,N_9522,N_8312);
and U11915 (N_11915,N_9952,N_8718);
nor U11916 (N_11916,N_9251,N_8170);
and U11917 (N_11917,N_9409,N_8975);
and U11918 (N_11918,N_9573,N_8421);
xor U11919 (N_11919,N_9546,N_9377);
or U11920 (N_11920,N_9284,N_9854);
and U11921 (N_11921,N_9036,N_9320);
nor U11922 (N_11922,N_9504,N_9458);
or U11923 (N_11923,N_8615,N_8395);
and U11924 (N_11924,N_8325,N_8411);
nor U11925 (N_11925,N_8972,N_9735);
nand U11926 (N_11926,N_9937,N_9384);
nor U11927 (N_11927,N_9726,N_9969);
or U11928 (N_11928,N_8518,N_8279);
xnor U11929 (N_11929,N_8947,N_9082);
or U11930 (N_11930,N_9394,N_8882);
xor U11931 (N_11931,N_8824,N_9127);
nor U11932 (N_11932,N_9969,N_8497);
and U11933 (N_11933,N_9483,N_9959);
nor U11934 (N_11934,N_9421,N_8014);
or U11935 (N_11935,N_8334,N_9760);
nand U11936 (N_11936,N_8220,N_9526);
or U11937 (N_11937,N_9090,N_8063);
nor U11938 (N_11938,N_9567,N_8337);
nor U11939 (N_11939,N_9809,N_9622);
and U11940 (N_11940,N_9984,N_9922);
xor U11941 (N_11941,N_8311,N_9459);
and U11942 (N_11942,N_9578,N_9170);
xnor U11943 (N_11943,N_8624,N_9701);
and U11944 (N_11944,N_9545,N_9209);
nor U11945 (N_11945,N_8181,N_8678);
or U11946 (N_11946,N_9088,N_9808);
and U11947 (N_11947,N_8493,N_8267);
nand U11948 (N_11948,N_9581,N_8495);
and U11949 (N_11949,N_9366,N_9512);
nand U11950 (N_11950,N_8988,N_9720);
nand U11951 (N_11951,N_9902,N_8213);
or U11952 (N_11952,N_8254,N_8812);
nor U11953 (N_11953,N_8182,N_9134);
or U11954 (N_11954,N_9436,N_9341);
nand U11955 (N_11955,N_9199,N_9693);
nand U11956 (N_11956,N_9148,N_8597);
nand U11957 (N_11957,N_8187,N_9099);
xor U11958 (N_11958,N_9100,N_8601);
nor U11959 (N_11959,N_9110,N_9989);
nor U11960 (N_11960,N_9668,N_8813);
xor U11961 (N_11961,N_8780,N_9353);
nor U11962 (N_11962,N_8060,N_8845);
xnor U11963 (N_11963,N_8207,N_9216);
xnor U11964 (N_11964,N_9339,N_9306);
nor U11965 (N_11965,N_9848,N_8912);
nand U11966 (N_11966,N_8093,N_9895);
or U11967 (N_11967,N_9353,N_9691);
xor U11968 (N_11968,N_9293,N_8847);
nand U11969 (N_11969,N_9600,N_9704);
and U11970 (N_11970,N_9947,N_9244);
and U11971 (N_11971,N_8772,N_9161);
and U11972 (N_11972,N_9685,N_8143);
nand U11973 (N_11973,N_9080,N_9918);
nor U11974 (N_11974,N_9248,N_9199);
nand U11975 (N_11975,N_9718,N_9058);
and U11976 (N_11976,N_9082,N_9381);
nand U11977 (N_11977,N_8132,N_8889);
or U11978 (N_11978,N_9187,N_8952);
or U11979 (N_11979,N_9784,N_8908);
xnor U11980 (N_11980,N_9606,N_8212);
or U11981 (N_11981,N_8838,N_8324);
nand U11982 (N_11982,N_9489,N_9814);
and U11983 (N_11983,N_9674,N_8905);
nand U11984 (N_11984,N_9767,N_8844);
xor U11985 (N_11985,N_9835,N_9405);
nand U11986 (N_11986,N_9664,N_9865);
or U11987 (N_11987,N_9589,N_8965);
nand U11988 (N_11988,N_9620,N_9127);
nor U11989 (N_11989,N_9770,N_8530);
and U11990 (N_11990,N_8755,N_8698);
nor U11991 (N_11991,N_9662,N_9821);
xnor U11992 (N_11992,N_8449,N_8321);
nand U11993 (N_11993,N_8908,N_9290);
nand U11994 (N_11994,N_8133,N_9358);
nand U11995 (N_11995,N_8928,N_8146);
and U11996 (N_11996,N_8550,N_9650);
nor U11997 (N_11997,N_8462,N_9735);
and U11998 (N_11998,N_9324,N_9529);
nor U11999 (N_11999,N_9268,N_8350);
nand U12000 (N_12000,N_10858,N_11433);
nand U12001 (N_12001,N_10430,N_10410);
or U12002 (N_12002,N_11247,N_11168);
nor U12003 (N_12003,N_10747,N_11937);
or U12004 (N_12004,N_10202,N_10805);
xor U12005 (N_12005,N_10975,N_11870);
and U12006 (N_12006,N_11879,N_10273);
or U12007 (N_12007,N_11628,N_10487);
nor U12008 (N_12008,N_10740,N_11051);
nor U12009 (N_12009,N_10292,N_10844);
nor U12010 (N_12010,N_11416,N_10614);
nor U12011 (N_12011,N_10655,N_11243);
nor U12012 (N_12012,N_11312,N_11999);
nand U12013 (N_12013,N_10117,N_10812);
nand U12014 (N_12014,N_11471,N_11455);
nand U12015 (N_12015,N_10676,N_10257);
or U12016 (N_12016,N_11677,N_10768);
xor U12017 (N_12017,N_11876,N_10016);
nand U12018 (N_12018,N_11304,N_10985);
and U12019 (N_12019,N_10871,N_10228);
nor U12020 (N_12020,N_10640,N_10759);
or U12021 (N_12021,N_11743,N_10903);
and U12022 (N_12022,N_11667,N_11380);
and U12023 (N_12023,N_11162,N_10279);
and U12024 (N_12024,N_11156,N_10637);
or U12025 (N_12025,N_11078,N_11596);
nand U12026 (N_12026,N_10245,N_11354);
and U12027 (N_12027,N_11980,N_10824);
xnor U12028 (N_12028,N_10666,N_11270);
and U12029 (N_12029,N_10719,N_11214);
or U12030 (N_12030,N_10504,N_11967);
nor U12031 (N_12031,N_11314,N_10745);
nand U12032 (N_12032,N_10814,N_11127);
xor U12033 (N_12033,N_11176,N_10393);
or U12034 (N_12034,N_11113,N_11619);
xnor U12035 (N_12035,N_10026,N_10645);
and U12036 (N_12036,N_11276,N_10936);
or U12037 (N_12037,N_10823,N_11396);
nand U12038 (N_12038,N_10594,N_10052);
or U12039 (N_12039,N_11068,N_10071);
nand U12040 (N_12040,N_11442,N_10875);
or U12041 (N_12041,N_10479,N_10746);
and U12042 (N_12042,N_11607,N_10529);
or U12043 (N_12043,N_10998,N_11942);
nor U12044 (N_12044,N_11634,N_11561);
nand U12045 (N_12045,N_11456,N_10475);
and U12046 (N_12046,N_11252,N_10857);
and U12047 (N_12047,N_10851,N_10883);
or U12048 (N_12048,N_11853,N_11324);
nor U12049 (N_12049,N_11576,N_10786);
or U12050 (N_12050,N_11079,N_10471);
or U12051 (N_12051,N_10456,N_11180);
and U12052 (N_12052,N_10911,N_10895);
or U12053 (N_12053,N_10653,N_10012);
and U12054 (N_12054,N_10760,N_10271);
nand U12055 (N_12055,N_11459,N_11152);
xor U12056 (N_12056,N_10879,N_10684);
nand U12057 (N_12057,N_10313,N_10801);
and U12058 (N_12058,N_11842,N_11787);
nand U12059 (N_12059,N_11222,N_10061);
nand U12060 (N_12060,N_10981,N_10606);
xor U12061 (N_12061,N_11328,N_11602);
and U12062 (N_12062,N_11150,N_11680);
or U12063 (N_12063,N_10333,N_11423);
or U12064 (N_12064,N_11378,N_11479);
nor U12065 (N_12065,N_10582,N_11262);
nand U12066 (N_12066,N_11996,N_11740);
nor U12067 (N_12067,N_11548,N_11827);
xor U12068 (N_12068,N_10596,N_10371);
and U12069 (N_12069,N_10652,N_10821);
nor U12070 (N_12070,N_11851,N_10656);
and U12071 (N_12071,N_10997,N_11541);
nand U12072 (N_12072,N_11374,N_10528);
nand U12073 (N_12073,N_11509,N_10396);
and U12074 (N_12074,N_11806,N_10015);
nor U12075 (N_12075,N_10426,N_10962);
nor U12076 (N_12076,N_10832,N_11462);
nor U12077 (N_12077,N_11552,N_11178);
and U12078 (N_12078,N_11791,N_10314);
xor U12079 (N_12079,N_10892,N_10711);
and U12080 (N_12080,N_10847,N_10086);
xor U12081 (N_12081,N_10534,N_11390);
or U12082 (N_12082,N_11935,N_11441);
or U12083 (N_12083,N_10349,N_11460);
xor U12084 (N_12084,N_11155,N_11898);
and U12085 (N_12085,N_10518,N_11090);
or U12086 (N_12086,N_11540,N_11712);
and U12087 (N_12087,N_11124,N_10638);
nand U12088 (N_12088,N_10930,N_10323);
nor U12089 (N_12089,N_10498,N_11517);
nor U12090 (N_12090,N_10695,N_10605);
nor U12091 (N_12091,N_10242,N_10113);
nor U12092 (N_12092,N_10904,N_11687);
or U12093 (N_12093,N_11313,N_11165);
and U12094 (N_12094,N_10566,N_11151);
nor U12095 (N_12095,N_10486,N_11543);
or U12096 (N_12096,N_10727,N_11398);
nor U12097 (N_12097,N_11055,N_11788);
nand U12098 (N_12098,N_10960,N_11816);
nor U12099 (N_12099,N_10675,N_10384);
nand U12100 (N_12100,N_10576,N_11504);
nor U12101 (N_12101,N_11902,N_11131);
or U12102 (N_12102,N_11502,N_11235);
and U12103 (N_12103,N_11148,N_10046);
nor U12104 (N_12104,N_10833,N_10574);
and U12105 (N_12105,N_11877,N_11708);
nand U12106 (N_12106,N_11317,N_10598);
nand U12107 (N_12107,N_10156,N_11869);
nor U12108 (N_12108,N_10386,N_11803);
and U12109 (N_12109,N_10929,N_11862);
xor U12110 (N_12110,N_10581,N_10575);
nor U12111 (N_12111,N_11301,N_10469);
nor U12112 (N_12112,N_10957,N_10146);
and U12113 (N_12113,N_11044,N_10216);
nand U12114 (N_12114,N_11624,N_10180);
xnor U12115 (N_12115,N_11498,N_11578);
or U12116 (N_12116,N_10618,N_11611);
nand U12117 (N_12117,N_10415,N_10934);
and U12118 (N_12118,N_10561,N_11261);
nor U12119 (N_12119,N_11691,N_10771);
nor U12120 (N_12120,N_11794,N_10447);
and U12121 (N_12121,N_11701,N_11973);
or U12122 (N_12122,N_11491,N_11207);
xnor U12123 (N_12123,N_11355,N_10753);
nand U12124 (N_12124,N_10213,N_10686);
nor U12125 (N_12125,N_11950,N_10478);
and U12126 (N_12126,N_11205,N_10733);
and U12127 (N_12127,N_11971,N_11177);
and U12128 (N_12128,N_11265,N_11626);
and U12129 (N_12129,N_10165,N_10115);
xnor U12130 (N_12130,N_10112,N_11285);
xor U12131 (N_12131,N_10119,N_11143);
or U12132 (N_12132,N_10214,N_11409);
xor U12133 (N_12133,N_11651,N_11434);
and U12134 (N_12134,N_10910,N_11329);
nor U12135 (N_12135,N_10099,N_11315);
xor U12136 (N_12136,N_11221,N_11437);
nand U12137 (N_12137,N_11196,N_10129);
or U12138 (N_12138,N_10822,N_10861);
nand U12139 (N_12139,N_10670,N_11883);
xnor U12140 (N_12140,N_10784,N_11192);
nand U12141 (N_12141,N_10192,N_11861);
or U12142 (N_12142,N_11856,N_10922);
nand U12143 (N_12143,N_10993,N_10405);
xnor U12144 (N_12144,N_11500,N_11960);
nor U12145 (N_12145,N_11213,N_10674);
xnor U12146 (N_12146,N_11257,N_11894);
xor U12147 (N_12147,N_11726,N_10246);
nor U12148 (N_12148,N_11103,N_11901);
or U12149 (N_12149,N_10159,N_10346);
and U12150 (N_12150,N_10231,N_11910);
nand U12151 (N_12151,N_10158,N_11246);
nor U12152 (N_12152,N_10151,N_11513);
or U12153 (N_12153,N_10427,N_10943);
and U12154 (N_12154,N_11287,N_10308);
nor U12155 (N_12155,N_11319,N_11425);
and U12156 (N_12156,N_10878,N_10380);
or U12157 (N_12157,N_11264,N_11949);
or U12158 (N_12158,N_11122,N_11318);
nor U12159 (N_12159,N_11091,N_10491);
xor U12160 (N_12160,N_10403,N_10586);
xor U12161 (N_12161,N_10890,N_10210);
and U12162 (N_12162,N_10541,N_11332);
nor U12163 (N_12163,N_10521,N_11917);
nor U12164 (N_12164,N_10697,N_11427);
nor U12165 (N_12165,N_11022,N_11195);
and U12166 (N_12166,N_11534,N_11941);
or U12167 (N_12167,N_11197,N_11719);
and U12168 (N_12168,N_10971,N_10177);
xnor U12169 (N_12169,N_10924,N_11623);
nor U12170 (N_12170,N_10630,N_10408);
and U12171 (N_12171,N_10704,N_11133);
nand U12172 (N_12172,N_10651,N_11249);
nor U12173 (N_12173,N_10796,N_10305);
nor U12174 (N_12174,N_10164,N_10340);
or U12175 (N_12175,N_10463,N_10546);
and U12176 (N_12176,N_11403,N_11684);
xnor U12177 (N_12177,N_10923,N_10064);
nand U12178 (N_12178,N_11410,N_10197);
and U12179 (N_12179,N_11829,N_11516);
or U12180 (N_12180,N_10963,N_11704);
or U12181 (N_12181,N_10617,N_11228);
nand U12182 (N_12182,N_10307,N_11369);
or U12183 (N_12183,N_11136,N_10100);
xor U12184 (N_12184,N_11105,N_11888);
or U12185 (N_12185,N_11116,N_10110);
nand U12186 (N_12186,N_10783,N_10735);
xor U12187 (N_12187,N_11190,N_11343);
and U12188 (N_12188,N_11050,N_11797);
or U12189 (N_12189,N_11102,N_11974);
xnor U12190 (N_12190,N_11957,N_11464);
nand U12191 (N_12191,N_10927,N_11563);
or U12192 (N_12192,N_10668,N_11478);
xor U12193 (N_12193,N_11027,N_10458);
or U12194 (N_12194,N_10664,N_11485);
and U12195 (N_12195,N_11017,N_10425);
or U12196 (N_12196,N_11739,N_10190);
nand U12197 (N_12197,N_11826,N_10820);
nand U12198 (N_12198,N_11036,N_11873);
xor U12199 (N_12199,N_11913,N_11008);
xor U12200 (N_12200,N_10979,N_11020);
nor U12201 (N_12201,N_10788,N_10438);
nor U12202 (N_12202,N_10986,N_11363);
and U12203 (N_12203,N_10310,N_11492);
xor U12204 (N_12204,N_10327,N_10633);
or U12205 (N_12205,N_11655,N_10530);
xnor U12206 (N_12206,N_11145,N_10264);
nor U12207 (N_12207,N_11832,N_11072);
xnor U12208 (N_12208,N_11801,N_10700);
nand U12209 (N_12209,N_11401,N_11557);
nor U12210 (N_12210,N_11411,N_10660);
nand U12211 (N_12211,N_11346,N_11848);
and U12212 (N_12212,N_11585,N_10692);
or U12213 (N_12213,N_11834,N_11203);
nor U12214 (N_12214,N_10553,N_10022);
or U12215 (N_12215,N_11223,N_10418);
nand U12216 (N_12216,N_10194,N_10090);
xor U12217 (N_12217,N_10466,N_11554);
xor U12218 (N_12218,N_11309,N_10807);
nand U12219 (N_12219,N_10073,N_11605);
nor U12220 (N_12220,N_10365,N_10034);
xnor U12221 (N_12221,N_10829,N_11533);
xor U12222 (N_12222,N_10564,N_10716);
and U12223 (N_12223,N_10688,N_10818);
and U12224 (N_12224,N_10137,N_11639);
nand U12225 (N_12225,N_10791,N_11250);
or U12226 (N_12226,N_11780,N_10226);
nand U12227 (N_12227,N_10414,N_10636);
or U12228 (N_12228,N_10173,N_11362);
nand U12229 (N_12229,N_10669,N_11279);
nor U12230 (N_12230,N_11393,N_10603);
and U12231 (N_12231,N_10162,N_11187);
or U12232 (N_12232,N_11277,N_10862);
nand U12233 (N_12233,N_11924,N_10799);
nor U12234 (N_12234,N_10992,N_10894);
or U12235 (N_12235,N_11449,N_11310);
nor U12236 (N_12236,N_10632,N_11544);
xnor U12237 (N_12237,N_11037,N_11920);
nor U12238 (N_12238,N_11060,N_11745);
nor U12239 (N_12239,N_10348,N_11340);
nand U12240 (N_12240,N_11388,N_11256);
xnor U12241 (N_12241,N_10610,N_10251);
xor U12242 (N_12242,N_10170,N_11397);
and U12243 (N_12243,N_10008,N_10255);
nor U12244 (N_12244,N_11087,N_10265);
xnor U12245 (N_12245,N_10131,N_11865);
nor U12246 (N_12246,N_11737,N_10145);
nor U12247 (N_12247,N_11731,N_11843);
xnor U12248 (N_12248,N_11267,N_10286);
and U12249 (N_12249,N_11721,N_10256);
nand U12250 (N_12250,N_11104,N_10247);
nand U12251 (N_12251,N_11665,N_10352);
and U12252 (N_12252,N_11515,N_10876);
and U12253 (N_12253,N_10881,N_11217);
or U12254 (N_12254,N_11367,N_10813);
nor U12255 (N_12255,N_10370,N_10258);
and U12256 (N_12256,N_11927,N_10542);
nand U12257 (N_12257,N_11146,N_10087);
nand U12258 (N_12258,N_11736,N_11850);
nor U12259 (N_12259,N_10056,N_10600);
nand U12260 (N_12260,N_10001,N_10284);
nand U12261 (N_12261,N_11061,N_11041);
and U12262 (N_12262,N_11738,N_10693);
nor U12263 (N_12263,N_11164,N_10472);
nand U12264 (N_12264,N_11053,N_11139);
nand U12265 (N_12265,N_10423,N_10299);
nor U12266 (N_12266,N_11450,N_10902);
xor U12267 (N_12267,N_11402,N_11753);
nor U12268 (N_12268,N_10744,N_11286);
and U12269 (N_12269,N_11336,N_11604);
nor U12270 (N_12270,N_10678,N_10317);
and U12271 (N_12271,N_10969,N_10767);
and U12272 (N_12272,N_10077,N_10958);
xnor U12273 (N_12273,N_10130,N_11849);
nand U12274 (N_12274,N_10374,N_10268);
xnor U12275 (N_12275,N_10267,N_10092);
nor U12276 (N_12276,N_11621,N_11505);
xnor U12277 (N_12277,N_11781,N_10175);
xnor U12278 (N_12278,N_11972,N_11184);
nand U12279 (N_12279,N_10188,N_11356);
nor U12280 (N_12280,N_10035,N_10182);
nand U12281 (N_12281,N_10762,N_11507);
nor U12282 (N_12282,N_11963,N_10391);
nand U12283 (N_12283,N_11887,N_11720);
nand U12284 (N_12284,N_11654,N_10815);
nor U12285 (N_12285,N_10913,N_10721);
xnor U12286 (N_12286,N_10587,N_11206);
or U12287 (N_12287,N_11334,N_10204);
nand U12288 (N_12288,N_10045,N_10431);
nor U12289 (N_12289,N_10094,N_11115);
and U12290 (N_12290,N_10989,N_10672);
nor U12291 (N_12291,N_10053,N_10178);
xnor U12292 (N_12292,N_10454,N_11609);
xor U12293 (N_12293,N_10749,N_11527);
nand U12294 (N_12294,N_10446,N_11703);
nand U12295 (N_12295,N_11348,N_10342);
or U12296 (N_12296,N_11063,N_10005);
xnor U12297 (N_12297,N_10863,N_10355);
or U12298 (N_12298,N_11379,N_11013);
nor U12299 (N_12299,N_11417,N_11762);
or U12300 (N_12300,N_11512,N_10161);
and U12301 (N_12301,N_11292,N_10114);
xnor U12302 (N_12302,N_10850,N_10207);
nand U12303 (N_12303,N_11149,N_10263);
or U12304 (N_12304,N_10461,N_11930);
or U12305 (N_12305,N_11606,N_11368);
xor U12306 (N_12306,N_11289,N_11137);
nor U12307 (N_12307,N_10961,N_11891);
nor U12308 (N_12308,N_10452,N_10383);
and U12309 (N_12309,N_11682,N_11538);
xor U12310 (N_12310,N_10450,N_11043);
nor U12311 (N_12311,N_10517,N_10144);
nor U12312 (N_12312,N_10545,N_11531);
xor U12313 (N_12313,N_10489,N_11792);
nand U12314 (N_12314,N_10728,N_11198);
or U12315 (N_12315,N_11990,N_10625);
nand U12316 (N_12316,N_11487,N_10168);
and U12317 (N_12317,N_10877,N_10773);
nand U12318 (N_12318,N_11448,N_11351);
or U12319 (N_12319,N_11350,N_10124);
nand U12320 (N_12320,N_10048,N_10017);
nor U12321 (N_12321,N_11650,N_11618);
and U12322 (N_12322,N_11057,N_11352);
nor U12323 (N_12323,N_11627,N_10027);
and U12324 (N_12324,N_11412,N_10031);
or U12325 (N_12325,N_10041,N_10069);
nand U12326 (N_12326,N_11486,N_11947);
nand U12327 (N_12327,N_10134,N_10933);
and U12328 (N_12328,N_11640,N_10343);
or U12329 (N_12329,N_10044,N_11391);
nand U12330 (N_12330,N_11642,N_11964);
and U12331 (N_12331,N_10908,N_10531);
xnor U12332 (N_12332,N_11290,N_11868);
nor U12333 (N_12333,N_10250,N_10217);
xor U12334 (N_12334,N_10921,N_11128);
xor U12335 (N_12335,N_11934,N_10649);
nor U12336 (N_12336,N_11896,N_11673);
xor U12337 (N_12337,N_11705,N_11847);
or U12338 (N_12338,N_11241,N_11763);
or U12339 (N_12339,N_10855,N_11988);
or U12340 (N_12340,N_10341,N_11259);
xnor U12341 (N_12341,N_11039,N_11546);
and U12342 (N_12342,N_11494,N_11188);
nand U12343 (N_12343,N_11166,N_11857);
nand U12344 (N_12344,N_10419,N_10220);
nor U12345 (N_12345,N_11777,N_11524);
nor U12346 (N_12346,N_10457,N_11383);
xor U12347 (N_12347,N_11770,N_11657);
xor U12348 (N_12348,N_11696,N_11229);
nor U12349 (N_12349,N_10339,N_10269);
or U12350 (N_12350,N_10780,N_11831);
xnor U12351 (N_12351,N_10208,N_10368);
xor U12352 (N_12352,N_10646,N_11824);
and U12353 (N_12353,N_11610,N_11638);
nand U12354 (N_12354,N_10639,N_10382);
nand U12355 (N_12355,N_10287,N_10750);
and U12356 (N_12356,N_11732,N_10535);
nand U12357 (N_12357,N_10502,N_11019);
and U12358 (N_12358,N_11723,N_10387);
or U12359 (N_12359,N_10853,N_11539);
and U12360 (N_12360,N_10560,N_11194);
nor U12361 (N_12361,N_10854,N_10098);
nor U12362 (N_12362,N_10155,N_10680);
nand U12363 (N_12363,N_10573,N_10211);
nand U12364 (N_12364,N_10532,N_10499);
or U12365 (N_12365,N_10888,N_11233);
or U12366 (N_12366,N_11923,N_11906);
nor U12367 (N_12367,N_10289,N_10239);
nand U12368 (N_12368,N_11929,N_10009);
nand U12369 (N_12369,N_11260,N_10301);
or U12370 (N_12370,N_10449,N_10353);
and U12371 (N_12371,N_10578,N_10991);
xnor U12372 (N_12372,N_11316,N_10905);
xnor U12373 (N_12373,N_11365,N_10623);
nor U12374 (N_12374,N_11339,N_11706);
nand U12375 (N_12375,N_11697,N_10650);
xnor U12376 (N_12376,N_10331,N_10174);
nor U12377 (N_12377,N_11987,N_11566);
nor U12378 (N_12378,N_11132,N_10729);
and U12379 (N_12379,N_10501,N_10334);
or U12380 (N_12380,N_10906,N_11303);
xor U12381 (N_12381,N_10482,N_11702);
and U12382 (N_12382,N_11945,N_10435);
and U12383 (N_12383,N_11900,N_10572);
or U12384 (N_12384,N_11083,N_10032);
xor U12385 (N_12385,N_11958,N_10831);
or U12386 (N_12386,N_11893,N_10337);
nor U12387 (N_12387,N_11892,N_11004);
xor U12388 (N_12388,N_10109,N_10551);
nand U12389 (N_12389,N_10677,N_11174);
or U12390 (N_12390,N_11200,N_10335);
nand U12391 (N_12391,N_10555,N_11911);
or U12392 (N_12392,N_11422,N_11191);
xor U12393 (N_12393,N_11889,N_11445);
xnor U12394 (N_12394,N_10152,N_11615);
and U12395 (N_12395,N_10051,N_10058);
and U12396 (N_12396,N_11179,N_10898);
nand U12397 (N_12397,N_10437,N_11820);
nand U12398 (N_12398,N_11981,N_11588);
xnor U12399 (N_12399,N_11674,N_11614);
nor U12400 (N_12400,N_10412,N_11522);
nand U12401 (N_12401,N_11147,N_10140);
or U12402 (N_12402,N_10607,N_11798);
xor U12403 (N_12403,N_10293,N_10148);
xor U12404 (N_12404,N_10141,N_10970);
nor U12405 (N_12405,N_10084,N_11685);
or U12406 (N_12406,N_11293,N_10955);
xor U12407 (N_12407,N_10054,N_11031);
or U12408 (N_12408,N_10602,N_10076);
nand U12409 (N_12409,N_11713,N_11404);
nor U12410 (N_12410,N_11899,N_11288);
nor U12411 (N_12411,N_11863,N_11240);
xnor U12412 (N_12412,N_11109,N_11111);
nand U12413 (N_12413,N_10253,N_10734);
or U12414 (N_12414,N_11431,N_10848);
and U12415 (N_12415,N_10329,N_11825);
nor U12416 (N_12416,N_10798,N_11234);
xnor U12417 (N_12417,N_10741,N_10549);
nand U12418 (N_12418,N_11038,N_10770);
xor U12419 (N_12419,N_11660,N_10235);
nor U12420 (N_12420,N_11699,N_11581);
xor U12421 (N_12421,N_10916,N_10667);
nor U12422 (N_12422,N_10224,N_11991);
nand U12423 (N_12423,N_10232,N_11098);
and U12424 (N_12424,N_10185,N_10731);
or U12425 (N_12425,N_11989,N_11366);
xnor U12426 (N_12426,N_10332,N_11428);
xor U12427 (N_12427,N_11926,N_11129);
or U12428 (N_12428,N_11421,N_10123);
and U12429 (N_12429,N_11590,N_10659);
nor U12430 (N_12430,N_11734,N_11466);
nand U12431 (N_12431,N_11413,N_10941);
nand U12432 (N_12432,N_10448,N_11962);
or U12433 (N_12433,N_10794,N_10626);
and U12434 (N_12434,N_10417,N_10066);
or U12435 (N_12435,N_10947,N_11473);
and U12436 (N_12436,N_11571,N_10931);
xor U12437 (N_12437,N_10023,N_11230);
nor U12438 (N_12438,N_11062,N_11707);
xor U12439 (N_12439,N_10774,N_10516);
or U12440 (N_12440,N_10462,N_10390);
xnor U12441 (N_12441,N_10157,N_10070);
xor U12442 (N_12442,N_11864,N_10205);
or U12443 (N_12443,N_11786,N_11694);
nand U12444 (N_12444,N_10868,N_10357);
nand U12445 (N_12445,N_10358,N_10184);
xnor U12446 (N_12446,N_11570,N_11599);
nor U12447 (N_12447,N_10834,N_11406);
or U12448 (N_12448,N_11114,N_11360);
nor U12449 (N_12449,N_10690,N_10689);
nand U12450 (N_12450,N_10477,N_11364);
nor U12451 (N_12451,N_11529,N_10647);
xnor U12452 (N_12452,N_11501,N_11756);
nand U12453 (N_12453,N_10938,N_10480);
xnor U12454 (N_12454,N_11955,N_10093);
or U12455 (N_12455,N_11922,N_11595);
xor U12456 (N_12456,N_11978,N_10275);
nand U12457 (N_12457,N_11302,N_10866);
or U12458 (N_12458,N_11817,N_10852);
or U12459 (N_12459,N_10554,N_11813);
nor U12460 (N_12460,N_10682,N_10738);
or U12461 (N_12461,N_10270,N_10359);
nor U12462 (N_12462,N_11014,N_11600);
xnor U12463 (N_12463,N_11679,N_11330);
nor U12464 (N_12464,N_11046,N_10191);
and U12465 (N_12465,N_10559,N_11714);
nor U12466 (N_12466,N_11603,N_11943);
and U12467 (N_12467,N_11633,N_10360);
or U12468 (N_12468,N_11451,N_10047);
or U12469 (N_12469,N_11749,N_10203);
or U12470 (N_12470,N_10000,N_11577);
xor U12471 (N_12471,N_10956,N_11185);
and U12472 (N_12472,N_10127,N_11536);
nor U12473 (N_12473,N_10918,N_11419);
and U12474 (N_12474,N_10136,N_11802);
nand U12475 (N_12475,N_10932,N_11371);
nand U12476 (N_12476,N_11426,N_11630);
and U12477 (N_12477,N_11054,N_11637);
nor U12478 (N_12478,N_10153,N_11938);
nor U12479 (N_12479,N_11347,N_11866);
nor U12480 (N_12480,N_11569,N_10404);
or U12481 (N_12481,N_10298,N_10379);
xnor U12482 (N_12482,N_11931,N_10886);
and U12483 (N_12483,N_10186,N_11231);
or U12484 (N_12484,N_10336,N_10976);
and U12485 (N_12485,N_10849,N_10588);
xnor U12486 (N_12486,N_10303,N_10550);
or U12487 (N_12487,N_11664,N_11649);
nor U12488 (N_12488,N_10830,N_10392);
and U12489 (N_12489,N_10608,N_10002);
and U12490 (N_12490,N_10252,N_10920);
and U12491 (N_12491,N_11181,N_11112);
or U12492 (N_12492,N_10460,N_10385);
nor U12493 (N_12493,N_10589,N_11333);
nand U12494 (N_12494,N_11032,N_11689);
or U12495 (N_12495,N_11890,N_11273);
nor U12496 (N_12496,N_10797,N_10497);
xor U12497 (N_12497,N_11154,N_10954);
nor U12498 (N_12498,N_11495,N_10965);
xor U12499 (N_12499,N_11503,N_11094);
nand U12500 (N_12500,N_11306,N_11698);
xor U12501 (N_12501,N_11307,N_11204);
or U12502 (N_12502,N_10864,N_10778);
or U12503 (N_12503,N_11182,N_11123);
nor U12504 (N_12504,N_11381,N_10030);
nand U12505 (N_12505,N_10615,N_10266);
or U12506 (N_12506,N_10540,N_10538);
nor U12507 (N_12507,N_11724,N_10199);
xnor U12508 (N_12508,N_11158,N_10154);
xnor U12509 (N_12509,N_11954,N_11555);
and U12510 (N_12510,N_10720,N_10973);
xor U12511 (N_12511,N_10227,N_10563);
nand U12512 (N_12512,N_11345,N_10928);
nor U12513 (N_12513,N_10484,N_11026);
nor U12514 (N_12514,N_11754,N_10003);
nor U12515 (N_12515,N_10409,N_11553);
and U12516 (N_12516,N_10398,N_11747);
and U12517 (N_12517,N_11729,N_10837);
xnor U12518 (N_12518,N_11526,N_10221);
xor U12519 (N_12519,N_10262,N_10974);
or U12520 (N_12520,N_11477,N_11484);
and U12521 (N_12521,N_10240,N_10867);
nand U12522 (N_12522,N_10732,N_10513);
and U12523 (N_12523,N_10751,N_11525);
nor U12524 (N_12524,N_10413,N_10241);
or U12525 (N_12525,N_10590,N_11499);
or U12526 (N_12526,N_11582,N_11771);
or U12527 (N_12527,N_10095,N_11659);
nor U12528 (N_12528,N_11173,N_11925);
nand U12529 (N_12529,N_11916,N_10362);
or U12530 (N_12530,N_11767,N_11171);
nor U12531 (N_12531,N_11676,N_11769);
xnor U12532 (N_12532,N_10291,N_11983);
or U12533 (N_12533,N_10951,N_11728);
and U12534 (N_12534,N_10490,N_10089);
xnor U12535 (N_12535,N_11744,N_11764);
or U12536 (N_12536,N_11444,N_10421);
or U12537 (N_12537,N_11224,N_11430);
xor U12538 (N_12538,N_10593,N_11021);
or U12539 (N_12539,N_10388,N_11092);
xor U12540 (N_12540,N_10597,N_10726);
nor U12541 (N_12541,N_11438,N_11097);
xnor U12542 (N_12542,N_11757,N_11066);
xnor U12543 (N_12543,N_10189,N_11040);
or U12544 (N_12544,N_11647,N_11349);
and U12545 (N_12545,N_10366,N_11994);
xor U12546 (N_12546,N_10067,N_10118);
or U12547 (N_12547,N_10433,N_11635);
or U12548 (N_12548,N_10533,N_11153);
nand U12549 (N_12549,N_10811,N_10354);
nor U12550 (N_12550,N_10967,N_11594);
or U12551 (N_12551,N_11034,N_10982);
nor U12552 (N_12552,N_10420,N_10539);
or U12553 (N_12553,N_10787,N_10785);
xnor U12554 (N_12554,N_11966,N_11237);
or U12555 (N_12555,N_11752,N_11928);
nand U12556 (N_12556,N_10887,N_11497);
and U12557 (N_12557,N_11049,N_11956);
xor U12558 (N_12558,N_11997,N_11625);
and U12559 (N_12559,N_11772,N_11119);
or U12560 (N_12560,N_10043,N_10116);
or U12561 (N_12561,N_10663,N_10743);
or U12562 (N_12562,N_10776,N_10520);
xor U12563 (N_12563,N_11608,N_11521);
xor U12564 (N_12564,N_11056,N_10580);
xor U12565 (N_12565,N_10707,N_10781);
nand U12566 (N_12566,N_10063,N_10036);
or U12567 (N_12567,N_10212,N_10133);
and U12568 (N_12568,N_10193,N_11810);
and U12569 (N_12569,N_11483,N_10244);
nor U12570 (N_12570,N_11007,N_10968);
xnor U12571 (N_12571,N_11574,N_10166);
xor U12572 (N_12572,N_10020,N_11523);
and U12573 (N_12573,N_11932,N_11912);
nor U12574 (N_12574,N_10160,N_10397);
nor U12575 (N_12575,N_11481,N_11386);
nor U12576 (N_12576,N_11436,N_11556);
nor U12577 (N_12577,N_10278,N_10453);
xor U12578 (N_12578,N_10024,N_11750);
or U12579 (N_12579,N_11337,N_11117);
and U12580 (N_12580,N_10592,N_10896);
nand U12581 (N_12581,N_11085,N_11361);
xnor U12582 (N_12582,N_10167,N_11511);
and U12583 (N_12583,N_10758,N_11075);
and U12584 (N_12584,N_11778,N_10147);
and U12585 (N_12585,N_11331,N_11035);
nand U12586 (N_12586,N_10978,N_11266);
nor U12587 (N_12587,N_11447,N_10309);
nand U12588 (N_12588,N_11535,N_11975);
nor U12589 (N_12589,N_10406,N_11760);
xor U12590 (N_12590,N_11807,N_11562);
nand U12591 (N_12591,N_10013,N_11789);
nor U12592 (N_12592,N_11245,N_11822);
xor U12593 (N_12593,N_11933,N_10500);
and U12594 (N_12594,N_10150,N_10233);
or U12595 (N_12595,N_11993,N_10643);
nand U12596 (N_12596,N_10795,N_11661);
nor U12597 (N_12597,N_11952,N_10565);
nand U12598 (N_12598,N_11951,N_11836);
and U12599 (N_12599,N_10282,N_11220);
and U12600 (N_12600,N_10584,N_11446);
nor U12601 (N_12601,N_11641,N_10940);
nor U12602 (N_12602,N_10401,N_10075);
or U12603 (N_12603,N_11226,N_10229);
nor U12604 (N_12604,N_11296,N_10378);
nor U12605 (N_12605,N_11755,N_11089);
nand U12606 (N_12606,N_11170,N_10874);
nor U12607 (N_12607,N_10543,N_11215);
xor U12608 (N_12608,N_11108,N_11846);
nor U12609 (N_12609,N_11692,N_10694);
xor U12610 (N_12610,N_10736,N_11016);
and U12611 (N_12611,N_10737,N_10761);
xor U12612 (N_12612,N_11457,N_10914);
or U12613 (N_12613,N_10277,N_10488);
nor U12614 (N_12614,N_10330,N_11811);
nand U12615 (N_12615,N_11939,N_10121);
nor U12616 (N_12616,N_10828,N_11844);
xnor U12617 (N_12617,N_10869,N_10619);
xor U12618 (N_12618,N_11283,N_10570);
nand U12619 (N_12619,N_11631,N_11295);
xor U12620 (N_12620,N_10826,N_11718);
xor U12621 (N_12621,N_11453,N_11167);
xnor U12622 (N_12622,N_11668,N_10808);
nand U12623 (N_12623,N_10884,N_11159);
and U12624 (N_12624,N_11389,N_11959);
nor U12625 (N_12625,N_10964,N_10966);
nor U12626 (N_12626,N_11311,N_10126);
xnor U12627 (N_12627,N_11297,N_10455);
nor U12628 (N_12628,N_10839,N_11686);
or U12629 (N_12629,N_10351,N_11979);
and U12630 (N_12630,N_11323,N_10018);
xor U12631 (N_12631,N_10757,N_10705);
or U12632 (N_12632,N_11727,N_11251);
nor U12633 (N_12633,N_11579,N_11835);
and U12634 (N_12634,N_10514,N_10754);
xnor U12635 (N_12635,N_10369,N_11622);
and U12636 (N_12636,N_10345,N_11418);
or U12637 (N_12637,N_11208,N_11800);
xor U12638 (N_12638,N_10096,N_11216);
nor U12639 (N_12639,N_11045,N_11096);
xnor U12640 (N_12640,N_10451,N_11884);
and U12641 (N_12641,N_10080,N_10508);
xor U12642 (N_12642,N_11305,N_11908);
xor U12643 (N_12643,N_10708,N_11711);
xnor U12644 (N_12644,N_11073,N_10503);
nor U12645 (N_12645,N_10583,N_10143);
or U12646 (N_12646,N_10492,N_10809);
nand U12647 (N_12647,N_10394,N_10524);
nand U12648 (N_12648,N_11169,N_11586);
or U12649 (N_12649,N_11520,N_11394);
nand U12650 (N_12650,N_11838,N_11768);
nor U12651 (N_12651,N_11775,N_10915);
or U12652 (N_12652,N_10326,N_10297);
nor U12653 (N_12653,N_10724,N_10860);
and U12654 (N_12654,N_10465,N_11465);
xnor U12655 (N_12655,N_11130,N_11201);
or U12656 (N_12656,N_10183,N_10710);
nor U12657 (N_12657,N_11280,N_10440);
xor U12658 (N_12658,N_10347,N_11766);
xor U12659 (N_12659,N_11918,N_11710);
nand U12660 (N_12660,N_11818,N_11023);
nand U12661 (N_12661,N_11812,N_11878);
and U12662 (N_12662,N_10055,N_11424);
nor U12663 (N_12663,N_11867,N_11144);
nand U12664 (N_12664,N_10613,N_11189);
nor U12665 (N_12665,N_10558,N_11909);
nand U12666 (N_12666,N_10389,N_10105);
nand U12667 (N_12667,N_11488,N_11833);
or U12668 (N_12668,N_10880,N_11670);
or U12669 (N_12669,N_10436,N_10079);
or U12670 (N_12670,N_11110,N_10375);
nand U12671 (N_12671,N_11904,N_10443);
nand U12672 (N_12672,N_11429,N_10980);
or U12673 (N_12673,N_10789,N_11468);
nor U12674 (N_12674,N_11968,N_10004);
xor U12675 (N_12675,N_10128,N_11489);
xnor U12676 (N_12676,N_10082,N_10222);
xor U12677 (N_12677,N_11341,N_10621);
nand U12678 (N_12678,N_10703,N_11746);
nand U12679 (N_12679,N_10782,N_10912);
or U12680 (N_12680,N_10698,N_11321);
nand U12681 (N_12681,N_11617,N_11258);
xor U12682 (N_12682,N_10644,N_10999);
nor U12683 (N_12683,N_10039,N_10944);
or U12684 (N_12684,N_11735,N_11254);
xnor U12685 (N_12685,N_10765,N_10428);
or U12686 (N_12686,N_11439,N_11395);
xnor U12687 (N_12687,N_11528,N_11976);
and U12688 (N_12688,N_10132,N_11461);
and U12689 (N_12689,N_10515,N_10952);
and U12690 (N_12690,N_10028,N_10085);
xor U12691 (N_12691,N_10562,N_10439);
or U12692 (N_12692,N_10803,N_10445);
nor U12693 (N_12693,N_11255,N_10671);
or U12694 (N_12694,N_10604,N_11058);
xnor U12695 (N_12695,N_11809,N_11567);
nor U12696 (N_12696,N_11669,N_11903);
and U12697 (N_12697,N_10648,N_10376);
or U12698 (N_12698,N_10654,N_11067);
and U12699 (N_12699,N_11944,N_10769);
nor U12700 (N_12700,N_11469,N_11052);
or U12701 (N_12701,N_11474,N_10470);
or U12702 (N_12702,N_11069,N_11443);
nor U12703 (N_12703,N_10476,N_10990);
or U12704 (N_12704,N_10779,N_10842);
nor U12705 (N_12705,N_10817,N_10350);
and U12706 (N_12706,N_11140,N_10907);
xor U12707 (N_12707,N_11064,N_10571);
xor U12708 (N_12708,N_10236,N_11193);
and U12709 (N_12709,N_11248,N_10622);
or U12710 (N_12710,N_11783,N_10935);
nor U12711 (N_12711,N_10523,N_10714);
and U12712 (N_12712,N_10328,N_10101);
or U12713 (N_12713,N_11385,N_11584);
xnor U12714 (N_12714,N_11210,N_10557);
nand U12715 (N_12715,N_10010,N_10025);
nor U12716 (N_12716,N_11860,N_11518);
and U12717 (N_12717,N_10033,N_10103);
nand U12718 (N_12718,N_11033,N_10198);
xnor U12719 (N_12719,N_11161,N_11612);
xnor U12720 (N_12720,N_10288,N_11070);
nand U12721 (N_12721,N_11080,N_10373);
and U12722 (N_12722,N_10631,N_11134);
and U12723 (N_12723,N_11709,N_11881);
or U12724 (N_12724,N_10062,N_11001);
nor U12725 (N_12725,N_11028,N_11163);
nand U12726 (N_12726,N_10172,N_11308);
nand U12727 (N_12727,N_11088,N_10984);
or U12728 (N_12728,N_10081,N_11010);
nand U12729 (N_12729,N_10169,N_11871);
nand U12730 (N_12730,N_11852,N_11560);
or U12731 (N_12731,N_11435,N_10699);
nand U12732 (N_12732,N_11805,N_10804);
xor U12733 (N_12733,N_10163,N_11244);
nor U12734 (N_12734,N_10909,N_10901);
and U12735 (N_12735,N_11326,N_11678);
xor U12736 (N_12736,N_10249,N_11629);
and U12737 (N_12737,N_10040,N_10616);
and U12738 (N_12738,N_10142,N_10544);
nand U12739 (N_12739,N_10712,N_10701);
and U12740 (N_12740,N_11452,N_11683);
nor U12741 (N_12741,N_10792,N_10122);
or U12742 (N_12742,N_10983,N_10261);
and U12743 (N_12743,N_11322,N_11202);
or U12744 (N_12744,N_11758,N_10318);
xnor U12745 (N_12745,N_10942,N_10548);
or U12746 (N_12746,N_10296,N_11885);
xnor U12747 (N_12747,N_11272,N_11344);
nand U12748 (N_12748,N_10206,N_10917);
xnor U12749 (N_12749,N_11828,N_10802);
xor U12750 (N_12750,N_11716,N_11093);
nor U12751 (N_12751,N_10237,N_10870);
and U12752 (N_12752,N_11965,N_10841);
nor U12753 (N_12753,N_11796,N_10635);
or U12754 (N_12754,N_11616,N_11225);
and U12755 (N_12755,N_10097,N_11558);
nand U12756 (N_12756,N_11157,N_10037);
nand U12757 (N_12757,N_11537,N_10179);
xor U12758 (N_12758,N_11765,N_11232);
nand U12759 (N_12759,N_10819,N_10091);
xor U12760 (N_12760,N_10074,N_10525);
and U12761 (N_12761,N_10280,N_11717);
nor U12762 (N_12762,N_11907,N_10657);
nand U12763 (N_12763,N_11646,N_10628);
nor U12764 (N_12764,N_11282,N_11940);
nand U12765 (N_12765,N_11011,N_11730);
nor U12766 (N_12766,N_11029,N_10407);
nand U12767 (N_12767,N_10764,N_11886);
nand U12768 (N_12768,N_10338,N_11681);
or U12769 (N_12769,N_11141,N_11227);
nand U12770 (N_12770,N_10953,N_11840);
xnor U12771 (N_12771,N_10464,N_10139);
and U12772 (N_12772,N_11593,N_11175);
and U12773 (N_12773,N_10507,N_11476);
xor U12774 (N_12774,N_10715,N_10537);
nand U12775 (N_12775,N_11977,N_11773);
xnor U12776 (N_12776,N_10579,N_10777);
and U12777 (N_12777,N_11126,N_11373);
xor U12778 (N_12778,N_11024,N_11821);
or U12779 (N_12779,N_11905,N_10364);
xnor U12780 (N_12780,N_10843,N_10591);
or U12781 (N_12781,N_11632,N_11874);
nor U12782 (N_12782,N_11510,N_11759);
and U12783 (N_12783,N_10441,N_11793);
and U12784 (N_12784,N_10474,N_10624);
and U12785 (N_12785,N_11671,N_11015);
nor U12786 (N_12786,N_11142,N_11815);
or U12787 (N_12787,N_10840,N_11002);
nor U12788 (N_12788,N_11785,N_10691);
nor U12789 (N_12789,N_11921,N_10416);
nand U12790 (N_12790,N_10363,N_10872);
or U12791 (N_12791,N_10395,N_11841);
xnor U12792 (N_12792,N_11086,N_11294);
or U12793 (N_12793,N_10315,N_10473);
and U12794 (N_12794,N_10512,N_11795);
nor U12795 (N_12795,N_10283,N_10215);
nand U12796 (N_12796,N_10810,N_10243);
or U12797 (N_12797,N_11653,N_11172);
nor U12798 (N_12798,N_10505,N_10059);
xor U12799 (N_12799,N_10138,N_11636);
and U12800 (N_12800,N_10948,N_11666);
and U12801 (N_12801,N_11325,N_10687);
xnor U12802 (N_12802,N_11101,N_11376);
and U12803 (N_12803,N_10014,N_11725);
or U12804 (N_12804,N_10367,N_11408);
xnor U12805 (N_12805,N_10065,N_10083);
and U12806 (N_12806,N_10344,N_10629);
nor U12807 (N_12807,N_11077,N_11100);
xnor U12808 (N_12808,N_11672,N_10107);
or U12809 (N_12809,N_10411,N_10361);
nor U12810 (N_12810,N_10994,N_10722);
and U12811 (N_12811,N_11338,N_11663);
or U12812 (N_12812,N_11018,N_10434);
and U12813 (N_12813,N_11644,N_10467);
or U12814 (N_12814,N_11998,N_10945);
xor U12815 (N_12815,N_11858,N_10899);
or U12816 (N_12816,N_10422,N_10891);
or U12817 (N_12817,N_11872,N_10424);
or U12818 (N_12818,N_11375,N_10937);
nand U12819 (N_12819,N_11839,N_10495);
nand U12820 (N_12820,N_10181,N_11662);
and U12821 (N_12821,N_10552,N_11219);
nor U12822 (N_12822,N_10510,N_11387);
nor U12823 (N_12823,N_11327,N_11915);
xnor U12824 (N_12824,N_10432,N_10281);
nor U12825 (N_12825,N_11583,N_10569);
or U12826 (N_12826,N_10919,N_11186);
or U12827 (N_12827,N_10007,N_11218);
xnor U12828 (N_12828,N_11414,N_11580);
nor U12829 (N_12829,N_10285,N_11587);
and U12830 (N_12830,N_11358,N_11969);
xnor U12831 (N_12831,N_11992,N_11377);
or U12832 (N_12832,N_10609,N_11009);
and U12833 (N_12833,N_11742,N_10889);
or U12834 (N_12834,N_10290,N_11542);
nand U12835 (N_12835,N_10634,N_10276);
and U12836 (N_12836,N_11550,N_10681);
nor U12837 (N_12837,N_11138,N_10611);
nor U12838 (N_12838,N_10149,N_11774);
and U12839 (N_12839,N_11565,N_10709);
and U12840 (N_12840,N_10859,N_10248);
nand U12841 (N_12841,N_11690,N_11382);
xnor U12842 (N_12842,N_11482,N_10356);
nand U12843 (N_12843,N_10377,N_10752);
or U12844 (N_12844,N_11480,N_10793);
nand U12845 (N_12845,N_10196,N_11278);
nor U12846 (N_12846,N_10950,N_11875);
and U12847 (N_12847,N_10620,N_11199);
or U12848 (N_12848,N_10325,N_11514);
xor U12849 (N_12849,N_10209,N_11790);
and U12850 (N_12850,N_10120,N_10519);
nand U12851 (N_12851,N_11291,N_11591);
nor U12852 (N_12852,N_11658,N_10259);
and U12853 (N_12853,N_11081,N_10585);
nor U12854 (N_12854,N_10577,N_10527);
xnor U12855 (N_12855,N_10068,N_11985);
or U12856 (N_12856,N_10302,N_11645);
nand U12857 (N_12857,N_10234,N_10755);
or U12858 (N_12858,N_10790,N_11372);
nand U12859 (N_12859,N_11601,N_10225);
nand U12860 (N_12860,N_10702,N_11568);
and U12861 (N_12861,N_11082,N_11135);
or U12862 (N_12862,N_10885,N_11532);
nand U12863 (N_12863,N_11946,N_10536);
or U12864 (N_12864,N_10468,N_11047);
or U12865 (N_12865,N_10713,N_11970);
nor U12866 (N_12866,N_10050,N_10972);
nor U12867 (N_12867,N_11025,N_11242);
nor U12868 (N_12868,N_11508,N_11722);
xnor U12869 (N_12869,N_10320,N_11120);
nand U12870 (N_12870,N_10522,N_11779);
and U12871 (N_12871,N_11420,N_10511);
nand U12872 (N_12872,N_11005,N_10200);
nand U12873 (N_12873,N_11961,N_10900);
and U12874 (N_12874,N_10195,N_11107);
nand U12875 (N_12875,N_11353,N_11733);
and U12876 (N_12876,N_11776,N_11106);
or U12877 (N_12877,N_11936,N_11823);
or U12878 (N_12878,N_10021,N_11239);
nor U12879 (N_12879,N_10845,N_10111);
xnor U12880 (N_12880,N_11125,N_10319);
xor U12881 (N_12881,N_10742,N_10219);
xor U12882 (N_12882,N_11253,N_10176);
nor U12883 (N_12883,N_10104,N_11059);
nor U12884 (N_12884,N_10772,N_10627);
nor U12885 (N_12885,N_11000,N_10612);
or U12886 (N_12886,N_10595,N_10493);
and U12887 (N_12887,N_11549,N_10661);
or U12888 (N_12888,N_11099,N_11012);
xor U12889 (N_12889,N_10042,N_11300);
xnor U12890 (N_12890,N_10836,N_11342);
xor U12891 (N_12891,N_11357,N_10506);
nand U12892 (N_12892,N_11880,N_11564);
nor U12893 (N_12893,N_11006,N_10816);
nor U12894 (N_12894,N_11095,N_10483);
xnor U12895 (N_12895,N_10106,N_11656);
xor U12896 (N_12896,N_10925,N_10223);
or U12897 (N_12897,N_11804,N_11209);
and U12898 (N_12898,N_11493,N_10088);
and U12899 (N_12899,N_11895,N_11048);
nor U12900 (N_12900,N_10775,N_10723);
or U12901 (N_12901,N_11652,N_11643);
nor U12902 (N_12902,N_11613,N_11897);
and U12903 (N_12903,N_10825,N_11271);
nand U12904 (N_12904,N_10171,N_10946);
xor U12905 (N_12905,N_10995,N_10254);
nand U12906 (N_12906,N_10057,N_11597);
or U12907 (N_12907,N_10856,N_11320);
and U12908 (N_12908,N_11814,N_11384);
nand U12909 (N_12909,N_10949,N_11986);
or U12910 (N_12910,N_11782,N_10274);
and U12911 (N_12911,N_10311,N_10187);
nand U12912 (N_12912,N_11715,N_10987);
xnor U12913 (N_12913,N_11238,N_10049);
nand U12914 (N_12914,N_11845,N_11405);
nand U12915 (N_12915,N_11953,N_11761);
nor U12916 (N_12916,N_11212,N_10429);
or U12917 (N_12917,N_11859,N_10547);
nand U12918 (N_12918,N_11071,N_10599);
nand U12919 (N_12919,N_10567,N_11160);
nand U12920 (N_12920,N_11432,N_10218);
and U12921 (N_12921,N_11003,N_10135);
xnor U12922 (N_12922,N_11030,N_11592);
nor U12923 (N_12923,N_10683,N_10102);
and U12924 (N_12924,N_11589,N_10019);
nor U12925 (N_12925,N_11598,N_10662);
and U12926 (N_12926,N_11370,N_11458);
and U12927 (N_12927,N_11984,N_11392);
or U12928 (N_12928,N_10316,N_10442);
nor U12929 (N_12929,N_11274,N_10496);
nor U12930 (N_12930,N_10996,N_10730);
and U12931 (N_12931,N_10642,N_11519);
nand U12932 (N_12932,N_10873,N_11074);
nand U12933 (N_12933,N_10272,N_11919);
xnor U12934 (N_12934,N_11236,N_11799);
or U12935 (N_12935,N_11855,N_11688);
or U12936 (N_12936,N_11675,N_10679);
or U12937 (N_12937,N_10230,N_10006);
nor U12938 (N_12938,N_11084,N_10568);
nor U12939 (N_12939,N_11530,N_10939);
nand U12940 (N_12940,N_11547,N_11837);
nor U12941 (N_12941,N_11400,N_10897);
xnor U12942 (N_12942,N_10763,N_11472);
nand U12943 (N_12943,N_11275,N_11042);
or U12944 (N_12944,N_10658,N_11808);
nor U12945 (N_12945,N_11545,N_11819);
xnor U12946 (N_12946,N_10806,N_11948);
xor U12947 (N_12947,N_10260,N_11121);
nand U12948 (N_12948,N_11299,N_10526);
and U12949 (N_12949,N_10717,N_11572);
nor U12950 (N_12950,N_10835,N_10402);
or U12951 (N_12951,N_10029,N_11407);
and U12952 (N_12952,N_10494,N_10988);
nand U12953 (N_12953,N_11335,N_11882);
nand U12954 (N_12954,N_11693,N_11475);
nand U12955 (N_12955,N_11748,N_11830);
nor U12956 (N_12956,N_10381,N_10846);
nand U12957 (N_12957,N_10011,N_10706);
and U12958 (N_12958,N_10959,N_11415);
nand U12959 (N_12959,N_10324,N_11700);
or U12960 (N_12960,N_10696,N_11470);
nand U12961 (N_12961,N_10673,N_11914);
and U12962 (N_12962,N_11751,N_10800);
nor U12963 (N_12963,N_11281,N_11463);
xnor U12964 (N_12964,N_10306,N_10865);
nor U12965 (N_12965,N_11211,N_11467);
nor U12966 (N_12966,N_10748,N_10312);
or U12967 (N_12967,N_10685,N_10485);
xor U12968 (N_12968,N_11573,N_11506);
or U12969 (N_12969,N_11399,N_10078);
nand U12970 (N_12970,N_11854,N_10300);
or U12971 (N_12971,N_11359,N_10295);
nor U12972 (N_12972,N_10641,N_10322);
or U12973 (N_12973,N_10481,N_10372);
nor U12974 (N_12974,N_11065,N_11559);
nand U12975 (N_12975,N_10400,N_10556);
nor U12976 (N_12976,N_10838,N_10766);
or U12977 (N_12977,N_11298,N_11263);
nor U12978 (N_12978,N_11454,N_11183);
or U12979 (N_12979,N_11118,N_10321);
nor U12980 (N_12980,N_11620,N_11551);
nor U12981 (N_12981,N_10060,N_10201);
nor U12982 (N_12982,N_10926,N_11076);
nand U12983 (N_12983,N_11741,N_10238);
and U12984 (N_12984,N_10601,N_10038);
nor U12985 (N_12985,N_10108,N_11648);
or U12986 (N_12986,N_10893,N_11284);
xor U12987 (N_12987,N_10725,N_10739);
and U12988 (N_12988,N_11982,N_11440);
nor U12989 (N_12989,N_10509,N_10444);
and U12990 (N_12990,N_10072,N_10827);
xor U12991 (N_12991,N_10294,N_11784);
nand U12992 (N_12992,N_11269,N_11695);
nand U12993 (N_12993,N_10882,N_10718);
nor U12994 (N_12994,N_11268,N_10459);
nor U12995 (N_12995,N_10399,N_10304);
nor U12996 (N_12996,N_11496,N_11995);
nand U12997 (N_12997,N_10125,N_11490);
nor U12998 (N_12998,N_10977,N_10756);
nor U12999 (N_12999,N_11575,N_10665);
or U13000 (N_13000,N_11270,N_11098);
xor U13001 (N_13001,N_10071,N_10908);
nand U13002 (N_13002,N_10913,N_11598);
nand U13003 (N_13003,N_11654,N_11405);
or U13004 (N_13004,N_10019,N_11421);
nand U13005 (N_13005,N_11137,N_10062);
nor U13006 (N_13006,N_11512,N_11288);
nor U13007 (N_13007,N_11736,N_11386);
nor U13008 (N_13008,N_11956,N_10013);
nor U13009 (N_13009,N_11757,N_11532);
nor U13010 (N_13010,N_10678,N_10982);
and U13011 (N_13011,N_10275,N_10729);
or U13012 (N_13012,N_10847,N_10057);
nor U13013 (N_13013,N_11646,N_11375);
and U13014 (N_13014,N_11399,N_11412);
xor U13015 (N_13015,N_10438,N_11753);
xor U13016 (N_13016,N_10745,N_11822);
xnor U13017 (N_13017,N_10359,N_11263);
and U13018 (N_13018,N_11327,N_10085);
and U13019 (N_13019,N_11672,N_10337);
nand U13020 (N_13020,N_10509,N_10500);
xnor U13021 (N_13021,N_11727,N_11692);
nor U13022 (N_13022,N_10872,N_10023);
nor U13023 (N_13023,N_11744,N_11356);
or U13024 (N_13024,N_11802,N_10971);
and U13025 (N_13025,N_10712,N_10792);
xnor U13026 (N_13026,N_10061,N_10581);
or U13027 (N_13027,N_10750,N_11410);
and U13028 (N_13028,N_10094,N_10270);
nor U13029 (N_13029,N_10461,N_11721);
xnor U13030 (N_13030,N_10617,N_10614);
and U13031 (N_13031,N_10222,N_11101);
or U13032 (N_13032,N_11158,N_11777);
nor U13033 (N_13033,N_11143,N_11403);
nor U13034 (N_13034,N_11551,N_11542);
xor U13035 (N_13035,N_10397,N_10108);
xor U13036 (N_13036,N_10979,N_11604);
nand U13037 (N_13037,N_10811,N_10019);
and U13038 (N_13038,N_11557,N_11217);
nand U13039 (N_13039,N_10713,N_10291);
and U13040 (N_13040,N_11196,N_10908);
nor U13041 (N_13041,N_11820,N_10996);
nand U13042 (N_13042,N_11844,N_11121);
xnor U13043 (N_13043,N_11962,N_11108);
xnor U13044 (N_13044,N_11494,N_11714);
nor U13045 (N_13045,N_10345,N_11211);
and U13046 (N_13046,N_10407,N_11314);
nand U13047 (N_13047,N_11321,N_11254);
xor U13048 (N_13048,N_11953,N_11178);
nand U13049 (N_13049,N_11000,N_11930);
nand U13050 (N_13050,N_11657,N_11627);
xor U13051 (N_13051,N_11959,N_10480);
xor U13052 (N_13052,N_10316,N_10419);
or U13053 (N_13053,N_10514,N_11645);
nor U13054 (N_13054,N_10941,N_10475);
xnor U13055 (N_13055,N_10313,N_10077);
and U13056 (N_13056,N_10861,N_11047);
nor U13057 (N_13057,N_11428,N_11791);
nand U13058 (N_13058,N_10305,N_10201);
xor U13059 (N_13059,N_10040,N_11622);
or U13060 (N_13060,N_10265,N_10924);
and U13061 (N_13061,N_11346,N_11743);
nor U13062 (N_13062,N_11261,N_10318);
or U13063 (N_13063,N_10612,N_11372);
and U13064 (N_13064,N_10212,N_11041);
xor U13065 (N_13065,N_11487,N_11723);
xnor U13066 (N_13066,N_11050,N_11809);
nor U13067 (N_13067,N_11676,N_11062);
xor U13068 (N_13068,N_10413,N_11348);
xor U13069 (N_13069,N_10457,N_10522);
or U13070 (N_13070,N_10775,N_10391);
nor U13071 (N_13071,N_11261,N_11119);
and U13072 (N_13072,N_10673,N_10714);
and U13073 (N_13073,N_11479,N_11213);
nor U13074 (N_13074,N_11071,N_10349);
nand U13075 (N_13075,N_10750,N_10974);
or U13076 (N_13076,N_11310,N_11001);
nor U13077 (N_13077,N_11823,N_10290);
nand U13078 (N_13078,N_10663,N_11621);
nand U13079 (N_13079,N_11609,N_11635);
nor U13080 (N_13080,N_11350,N_10828);
and U13081 (N_13081,N_10026,N_11622);
nand U13082 (N_13082,N_11023,N_11888);
xnor U13083 (N_13083,N_10138,N_10556);
and U13084 (N_13084,N_10237,N_11386);
xor U13085 (N_13085,N_10377,N_10595);
or U13086 (N_13086,N_10222,N_11351);
nor U13087 (N_13087,N_10942,N_10360);
and U13088 (N_13088,N_11873,N_11655);
xor U13089 (N_13089,N_10259,N_11359);
xnor U13090 (N_13090,N_10327,N_11681);
nand U13091 (N_13091,N_11267,N_10551);
and U13092 (N_13092,N_11048,N_10696);
and U13093 (N_13093,N_10579,N_10318);
nand U13094 (N_13094,N_10314,N_10886);
or U13095 (N_13095,N_10239,N_11896);
and U13096 (N_13096,N_10244,N_11930);
nor U13097 (N_13097,N_11120,N_10455);
nand U13098 (N_13098,N_11913,N_11602);
and U13099 (N_13099,N_10598,N_11804);
or U13100 (N_13100,N_11641,N_10938);
nand U13101 (N_13101,N_10892,N_11977);
xnor U13102 (N_13102,N_11035,N_11334);
xor U13103 (N_13103,N_10120,N_11230);
and U13104 (N_13104,N_11141,N_11566);
xor U13105 (N_13105,N_10756,N_11863);
or U13106 (N_13106,N_11345,N_10747);
and U13107 (N_13107,N_10302,N_11601);
and U13108 (N_13108,N_11553,N_10170);
nor U13109 (N_13109,N_11040,N_10226);
nand U13110 (N_13110,N_11366,N_10193);
or U13111 (N_13111,N_11740,N_10684);
and U13112 (N_13112,N_11809,N_11575);
nand U13113 (N_13113,N_11752,N_11306);
nor U13114 (N_13114,N_11736,N_11973);
nor U13115 (N_13115,N_10754,N_10454);
or U13116 (N_13116,N_10970,N_10674);
and U13117 (N_13117,N_10347,N_11770);
nand U13118 (N_13118,N_11725,N_10090);
and U13119 (N_13119,N_11635,N_10377);
nand U13120 (N_13120,N_11254,N_10958);
or U13121 (N_13121,N_10088,N_10947);
or U13122 (N_13122,N_10695,N_10748);
xnor U13123 (N_13123,N_10307,N_11469);
or U13124 (N_13124,N_11008,N_10607);
nor U13125 (N_13125,N_11350,N_11846);
nand U13126 (N_13126,N_10491,N_10521);
and U13127 (N_13127,N_10919,N_10832);
nor U13128 (N_13128,N_11360,N_10223);
xor U13129 (N_13129,N_11021,N_10948);
or U13130 (N_13130,N_10934,N_11576);
nor U13131 (N_13131,N_10161,N_11319);
nand U13132 (N_13132,N_10727,N_11745);
and U13133 (N_13133,N_11490,N_10474);
or U13134 (N_13134,N_11323,N_11681);
and U13135 (N_13135,N_10434,N_11260);
nand U13136 (N_13136,N_11481,N_10853);
and U13137 (N_13137,N_11231,N_10014);
or U13138 (N_13138,N_10580,N_10533);
nor U13139 (N_13139,N_11433,N_11656);
or U13140 (N_13140,N_10913,N_10544);
xnor U13141 (N_13141,N_10162,N_10887);
or U13142 (N_13142,N_10228,N_10544);
and U13143 (N_13143,N_11226,N_10596);
and U13144 (N_13144,N_11722,N_11140);
xnor U13145 (N_13145,N_10173,N_11221);
or U13146 (N_13146,N_10202,N_11900);
and U13147 (N_13147,N_11080,N_11790);
and U13148 (N_13148,N_10184,N_11970);
nor U13149 (N_13149,N_10198,N_11403);
and U13150 (N_13150,N_11031,N_10096);
xor U13151 (N_13151,N_11879,N_10213);
or U13152 (N_13152,N_11948,N_11940);
xor U13153 (N_13153,N_10946,N_10446);
and U13154 (N_13154,N_11778,N_10945);
or U13155 (N_13155,N_11099,N_10598);
or U13156 (N_13156,N_11121,N_10264);
nand U13157 (N_13157,N_11315,N_10993);
nor U13158 (N_13158,N_11431,N_10940);
and U13159 (N_13159,N_10233,N_11014);
xnor U13160 (N_13160,N_11829,N_11709);
nor U13161 (N_13161,N_10132,N_11222);
and U13162 (N_13162,N_10952,N_11369);
xnor U13163 (N_13163,N_10800,N_10301);
xnor U13164 (N_13164,N_10305,N_10661);
or U13165 (N_13165,N_10636,N_10537);
and U13166 (N_13166,N_10753,N_10252);
nor U13167 (N_13167,N_11654,N_10282);
and U13168 (N_13168,N_10086,N_11461);
and U13169 (N_13169,N_10109,N_10167);
nor U13170 (N_13170,N_10365,N_10572);
or U13171 (N_13171,N_10073,N_10006);
xor U13172 (N_13172,N_11608,N_10380);
nand U13173 (N_13173,N_10040,N_10763);
and U13174 (N_13174,N_10626,N_10128);
or U13175 (N_13175,N_11141,N_10366);
nor U13176 (N_13176,N_10662,N_11072);
nor U13177 (N_13177,N_10366,N_11367);
nand U13178 (N_13178,N_10369,N_10348);
and U13179 (N_13179,N_10524,N_11998);
nor U13180 (N_13180,N_11685,N_10607);
nand U13181 (N_13181,N_10724,N_10816);
or U13182 (N_13182,N_11278,N_11638);
xnor U13183 (N_13183,N_10175,N_10826);
nor U13184 (N_13184,N_10262,N_11086);
or U13185 (N_13185,N_11293,N_10521);
and U13186 (N_13186,N_11885,N_10692);
nor U13187 (N_13187,N_11314,N_11669);
or U13188 (N_13188,N_11910,N_10825);
and U13189 (N_13189,N_10033,N_10946);
and U13190 (N_13190,N_11558,N_10369);
or U13191 (N_13191,N_10972,N_11553);
nor U13192 (N_13192,N_10884,N_11981);
nand U13193 (N_13193,N_11115,N_11288);
and U13194 (N_13194,N_10574,N_10944);
nand U13195 (N_13195,N_10663,N_11034);
nor U13196 (N_13196,N_10840,N_10622);
or U13197 (N_13197,N_10341,N_11246);
or U13198 (N_13198,N_11312,N_10534);
and U13199 (N_13199,N_10677,N_11695);
nor U13200 (N_13200,N_10182,N_11957);
and U13201 (N_13201,N_11859,N_10938);
or U13202 (N_13202,N_11957,N_10675);
and U13203 (N_13203,N_11027,N_11194);
or U13204 (N_13204,N_11854,N_11416);
or U13205 (N_13205,N_11351,N_11639);
or U13206 (N_13206,N_11327,N_10137);
nand U13207 (N_13207,N_11622,N_11521);
or U13208 (N_13208,N_11497,N_11643);
nand U13209 (N_13209,N_10239,N_11508);
and U13210 (N_13210,N_10855,N_10069);
nor U13211 (N_13211,N_10999,N_10756);
nand U13212 (N_13212,N_10003,N_10515);
xor U13213 (N_13213,N_11365,N_10769);
nor U13214 (N_13214,N_11898,N_10300);
nand U13215 (N_13215,N_10292,N_11234);
nor U13216 (N_13216,N_11248,N_11311);
or U13217 (N_13217,N_10004,N_10418);
xor U13218 (N_13218,N_11179,N_11028);
nor U13219 (N_13219,N_10654,N_10879);
and U13220 (N_13220,N_10189,N_11375);
nor U13221 (N_13221,N_10521,N_10368);
xnor U13222 (N_13222,N_10167,N_10860);
xnor U13223 (N_13223,N_11014,N_11811);
nand U13224 (N_13224,N_11551,N_11197);
and U13225 (N_13225,N_10229,N_11513);
and U13226 (N_13226,N_10083,N_11378);
or U13227 (N_13227,N_10913,N_10794);
nor U13228 (N_13228,N_11323,N_10641);
nand U13229 (N_13229,N_10466,N_11026);
or U13230 (N_13230,N_11538,N_10554);
nand U13231 (N_13231,N_10966,N_10088);
or U13232 (N_13232,N_11012,N_10504);
nand U13233 (N_13233,N_10185,N_10713);
nor U13234 (N_13234,N_11751,N_11755);
nor U13235 (N_13235,N_11979,N_11213);
nor U13236 (N_13236,N_11151,N_10060);
xnor U13237 (N_13237,N_10489,N_10415);
and U13238 (N_13238,N_10166,N_11478);
xor U13239 (N_13239,N_10677,N_10886);
xor U13240 (N_13240,N_10846,N_10567);
or U13241 (N_13241,N_10316,N_11323);
or U13242 (N_13242,N_10173,N_11523);
xor U13243 (N_13243,N_11140,N_11600);
nand U13244 (N_13244,N_10922,N_11703);
or U13245 (N_13245,N_10240,N_10850);
nand U13246 (N_13246,N_11117,N_11633);
xor U13247 (N_13247,N_10506,N_11409);
xor U13248 (N_13248,N_11096,N_10568);
nand U13249 (N_13249,N_11524,N_11228);
and U13250 (N_13250,N_11621,N_10838);
and U13251 (N_13251,N_11032,N_10113);
and U13252 (N_13252,N_10248,N_10756);
and U13253 (N_13253,N_11742,N_11666);
xor U13254 (N_13254,N_11470,N_11041);
and U13255 (N_13255,N_10799,N_10095);
nor U13256 (N_13256,N_11747,N_11666);
nand U13257 (N_13257,N_10339,N_10228);
or U13258 (N_13258,N_10469,N_11953);
xor U13259 (N_13259,N_10422,N_11142);
and U13260 (N_13260,N_11838,N_11627);
or U13261 (N_13261,N_11342,N_11928);
xnor U13262 (N_13262,N_10299,N_10923);
and U13263 (N_13263,N_10340,N_10144);
and U13264 (N_13264,N_11761,N_10027);
or U13265 (N_13265,N_10613,N_10458);
nor U13266 (N_13266,N_11915,N_11189);
nor U13267 (N_13267,N_10288,N_11623);
xnor U13268 (N_13268,N_10144,N_10830);
xor U13269 (N_13269,N_10207,N_11527);
and U13270 (N_13270,N_11386,N_11087);
xor U13271 (N_13271,N_10254,N_11029);
xor U13272 (N_13272,N_10881,N_11826);
or U13273 (N_13273,N_11515,N_10929);
and U13274 (N_13274,N_10335,N_10895);
or U13275 (N_13275,N_11909,N_10851);
or U13276 (N_13276,N_10854,N_11702);
and U13277 (N_13277,N_10029,N_11175);
and U13278 (N_13278,N_10773,N_11111);
xor U13279 (N_13279,N_11960,N_10716);
and U13280 (N_13280,N_10932,N_11352);
and U13281 (N_13281,N_11218,N_11960);
and U13282 (N_13282,N_11342,N_10551);
nor U13283 (N_13283,N_10615,N_10538);
xor U13284 (N_13284,N_11834,N_10995);
nor U13285 (N_13285,N_11440,N_10210);
xor U13286 (N_13286,N_11760,N_11330);
nand U13287 (N_13287,N_11187,N_11810);
xor U13288 (N_13288,N_11699,N_10928);
or U13289 (N_13289,N_11744,N_11076);
or U13290 (N_13290,N_11615,N_10448);
nand U13291 (N_13291,N_11038,N_11078);
nand U13292 (N_13292,N_10868,N_11405);
and U13293 (N_13293,N_11500,N_10968);
nor U13294 (N_13294,N_10329,N_11211);
and U13295 (N_13295,N_11810,N_11985);
nor U13296 (N_13296,N_10523,N_11128);
and U13297 (N_13297,N_10591,N_11604);
xnor U13298 (N_13298,N_10339,N_11601);
nor U13299 (N_13299,N_10481,N_11735);
nor U13300 (N_13300,N_10283,N_10572);
nand U13301 (N_13301,N_10928,N_11672);
and U13302 (N_13302,N_11807,N_10807);
nor U13303 (N_13303,N_10658,N_11054);
nor U13304 (N_13304,N_10052,N_10838);
nand U13305 (N_13305,N_11734,N_10723);
nor U13306 (N_13306,N_10368,N_10922);
nor U13307 (N_13307,N_10929,N_10235);
xnor U13308 (N_13308,N_11367,N_11464);
and U13309 (N_13309,N_11925,N_11333);
or U13310 (N_13310,N_10605,N_10860);
nand U13311 (N_13311,N_11630,N_10844);
and U13312 (N_13312,N_11873,N_11323);
nand U13313 (N_13313,N_11531,N_10647);
xnor U13314 (N_13314,N_10356,N_10634);
or U13315 (N_13315,N_11212,N_10345);
xnor U13316 (N_13316,N_11253,N_10398);
nor U13317 (N_13317,N_10566,N_10348);
nor U13318 (N_13318,N_10812,N_11050);
or U13319 (N_13319,N_11460,N_11301);
or U13320 (N_13320,N_10049,N_10474);
and U13321 (N_13321,N_10989,N_11940);
xnor U13322 (N_13322,N_10960,N_10971);
nor U13323 (N_13323,N_11231,N_10864);
and U13324 (N_13324,N_11869,N_10107);
and U13325 (N_13325,N_10493,N_10815);
or U13326 (N_13326,N_11594,N_11950);
and U13327 (N_13327,N_11050,N_10088);
and U13328 (N_13328,N_11836,N_11623);
and U13329 (N_13329,N_10607,N_10146);
nand U13330 (N_13330,N_11392,N_10514);
or U13331 (N_13331,N_10506,N_11197);
or U13332 (N_13332,N_10197,N_10498);
nand U13333 (N_13333,N_10559,N_10823);
xor U13334 (N_13334,N_10594,N_11185);
nor U13335 (N_13335,N_11697,N_10356);
nand U13336 (N_13336,N_11587,N_11586);
xnor U13337 (N_13337,N_10611,N_10313);
xnor U13338 (N_13338,N_11882,N_10789);
nor U13339 (N_13339,N_11622,N_10055);
xnor U13340 (N_13340,N_11635,N_11457);
xor U13341 (N_13341,N_11580,N_10105);
or U13342 (N_13342,N_10167,N_10342);
nor U13343 (N_13343,N_10969,N_10413);
xnor U13344 (N_13344,N_11838,N_10405);
and U13345 (N_13345,N_11748,N_11044);
nand U13346 (N_13346,N_10684,N_11403);
and U13347 (N_13347,N_10249,N_11628);
xor U13348 (N_13348,N_10128,N_11657);
nor U13349 (N_13349,N_11083,N_11539);
nand U13350 (N_13350,N_11937,N_10063);
or U13351 (N_13351,N_10811,N_11395);
or U13352 (N_13352,N_10109,N_10057);
nand U13353 (N_13353,N_10649,N_10662);
nor U13354 (N_13354,N_11068,N_11006);
nor U13355 (N_13355,N_11637,N_10963);
or U13356 (N_13356,N_11990,N_10839);
nand U13357 (N_13357,N_11375,N_11323);
and U13358 (N_13358,N_10726,N_10903);
and U13359 (N_13359,N_11307,N_10453);
nor U13360 (N_13360,N_11316,N_11453);
nor U13361 (N_13361,N_11919,N_11890);
xnor U13362 (N_13362,N_10433,N_10655);
or U13363 (N_13363,N_10957,N_11680);
nand U13364 (N_13364,N_11722,N_11283);
xnor U13365 (N_13365,N_10401,N_11406);
nand U13366 (N_13366,N_10717,N_10751);
nor U13367 (N_13367,N_11787,N_11129);
xnor U13368 (N_13368,N_10375,N_11637);
and U13369 (N_13369,N_11337,N_11870);
and U13370 (N_13370,N_11516,N_10051);
xnor U13371 (N_13371,N_10058,N_11769);
nand U13372 (N_13372,N_10926,N_10540);
or U13373 (N_13373,N_11585,N_10551);
xnor U13374 (N_13374,N_11180,N_11600);
nand U13375 (N_13375,N_10685,N_11398);
or U13376 (N_13376,N_10130,N_11506);
nand U13377 (N_13377,N_11606,N_11695);
nor U13378 (N_13378,N_10950,N_11656);
nor U13379 (N_13379,N_11041,N_10943);
or U13380 (N_13380,N_10654,N_10512);
or U13381 (N_13381,N_11919,N_10671);
nor U13382 (N_13382,N_11739,N_11751);
and U13383 (N_13383,N_11211,N_10597);
nor U13384 (N_13384,N_10940,N_10454);
nor U13385 (N_13385,N_11434,N_11849);
nand U13386 (N_13386,N_10963,N_10776);
xor U13387 (N_13387,N_11863,N_10859);
nand U13388 (N_13388,N_11722,N_10066);
nor U13389 (N_13389,N_10011,N_10816);
nand U13390 (N_13390,N_11438,N_10619);
nand U13391 (N_13391,N_11464,N_11223);
xnor U13392 (N_13392,N_10353,N_10589);
nand U13393 (N_13393,N_11108,N_11864);
nand U13394 (N_13394,N_10393,N_10409);
or U13395 (N_13395,N_10518,N_11040);
nand U13396 (N_13396,N_10407,N_11685);
or U13397 (N_13397,N_11726,N_11277);
nor U13398 (N_13398,N_11432,N_11853);
nor U13399 (N_13399,N_11447,N_10916);
xor U13400 (N_13400,N_10880,N_11293);
xor U13401 (N_13401,N_11269,N_11674);
or U13402 (N_13402,N_10107,N_11428);
xor U13403 (N_13403,N_11233,N_11726);
or U13404 (N_13404,N_11221,N_10124);
xnor U13405 (N_13405,N_10166,N_11540);
nor U13406 (N_13406,N_11832,N_11569);
and U13407 (N_13407,N_10253,N_11360);
and U13408 (N_13408,N_10048,N_10262);
xnor U13409 (N_13409,N_10851,N_10029);
nor U13410 (N_13410,N_11057,N_10219);
and U13411 (N_13411,N_11379,N_10927);
or U13412 (N_13412,N_11797,N_10888);
or U13413 (N_13413,N_10444,N_11555);
nor U13414 (N_13414,N_11647,N_11174);
nor U13415 (N_13415,N_10474,N_10517);
nand U13416 (N_13416,N_10438,N_11393);
and U13417 (N_13417,N_10674,N_11080);
and U13418 (N_13418,N_11749,N_10849);
and U13419 (N_13419,N_11246,N_11085);
nand U13420 (N_13420,N_10948,N_11297);
nand U13421 (N_13421,N_10868,N_10964);
nor U13422 (N_13422,N_11629,N_11926);
or U13423 (N_13423,N_11436,N_10725);
nor U13424 (N_13424,N_11633,N_11608);
nand U13425 (N_13425,N_10970,N_10181);
nand U13426 (N_13426,N_10358,N_10464);
xnor U13427 (N_13427,N_10825,N_10837);
nand U13428 (N_13428,N_10062,N_10450);
and U13429 (N_13429,N_10736,N_11761);
nor U13430 (N_13430,N_10439,N_11647);
nor U13431 (N_13431,N_11446,N_10997);
nand U13432 (N_13432,N_11922,N_11857);
xnor U13433 (N_13433,N_11930,N_10448);
and U13434 (N_13434,N_10359,N_10876);
nand U13435 (N_13435,N_10270,N_11833);
nor U13436 (N_13436,N_11076,N_10215);
and U13437 (N_13437,N_10963,N_11968);
and U13438 (N_13438,N_10026,N_10804);
xor U13439 (N_13439,N_10405,N_10041);
xnor U13440 (N_13440,N_10053,N_10953);
xor U13441 (N_13441,N_11693,N_11374);
nand U13442 (N_13442,N_10324,N_10083);
and U13443 (N_13443,N_11531,N_11416);
xnor U13444 (N_13444,N_10584,N_11453);
nand U13445 (N_13445,N_11419,N_10342);
xor U13446 (N_13446,N_11141,N_11172);
nor U13447 (N_13447,N_11041,N_11263);
and U13448 (N_13448,N_10272,N_10528);
and U13449 (N_13449,N_11864,N_10526);
nor U13450 (N_13450,N_11545,N_11382);
or U13451 (N_13451,N_10120,N_11587);
nand U13452 (N_13452,N_10246,N_10725);
nand U13453 (N_13453,N_10451,N_10880);
and U13454 (N_13454,N_10616,N_11650);
xnor U13455 (N_13455,N_11605,N_11343);
xnor U13456 (N_13456,N_11959,N_10960);
xnor U13457 (N_13457,N_11501,N_11239);
and U13458 (N_13458,N_11860,N_11530);
xor U13459 (N_13459,N_10082,N_11065);
nor U13460 (N_13460,N_10238,N_10712);
nand U13461 (N_13461,N_11533,N_11749);
and U13462 (N_13462,N_10173,N_10742);
nor U13463 (N_13463,N_11429,N_10070);
xnor U13464 (N_13464,N_11023,N_11397);
nand U13465 (N_13465,N_11439,N_11366);
nand U13466 (N_13466,N_10803,N_11424);
or U13467 (N_13467,N_10127,N_11474);
nand U13468 (N_13468,N_10437,N_10636);
nand U13469 (N_13469,N_10540,N_10419);
nand U13470 (N_13470,N_11011,N_11595);
or U13471 (N_13471,N_11551,N_10385);
or U13472 (N_13472,N_11798,N_10624);
nand U13473 (N_13473,N_10551,N_11496);
nor U13474 (N_13474,N_10255,N_10740);
nor U13475 (N_13475,N_11647,N_11281);
nor U13476 (N_13476,N_10539,N_11840);
and U13477 (N_13477,N_11438,N_11200);
or U13478 (N_13478,N_10607,N_10833);
and U13479 (N_13479,N_10890,N_10903);
nor U13480 (N_13480,N_11409,N_11767);
or U13481 (N_13481,N_11361,N_10254);
xnor U13482 (N_13482,N_10180,N_11311);
nand U13483 (N_13483,N_10117,N_11864);
xor U13484 (N_13484,N_10082,N_11944);
nor U13485 (N_13485,N_11313,N_11233);
xor U13486 (N_13486,N_11494,N_11862);
and U13487 (N_13487,N_10056,N_10404);
or U13488 (N_13488,N_10711,N_10173);
nor U13489 (N_13489,N_10838,N_11581);
nand U13490 (N_13490,N_11764,N_11057);
nand U13491 (N_13491,N_10120,N_11734);
and U13492 (N_13492,N_11320,N_11082);
xnor U13493 (N_13493,N_10385,N_11474);
xnor U13494 (N_13494,N_10682,N_11323);
xnor U13495 (N_13495,N_10524,N_11426);
xor U13496 (N_13496,N_10900,N_11665);
or U13497 (N_13497,N_10982,N_11817);
nand U13498 (N_13498,N_10276,N_10053);
or U13499 (N_13499,N_11142,N_11808);
nor U13500 (N_13500,N_10159,N_11250);
or U13501 (N_13501,N_10584,N_10000);
xor U13502 (N_13502,N_10829,N_11322);
and U13503 (N_13503,N_10275,N_10894);
nor U13504 (N_13504,N_10673,N_11915);
nand U13505 (N_13505,N_11267,N_10111);
nor U13506 (N_13506,N_11127,N_11526);
nor U13507 (N_13507,N_10767,N_10292);
nor U13508 (N_13508,N_10669,N_10108);
xnor U13509 (N_13509,N_10674,N_10825);
and U13510 (N_13510,N_10338,N_11759);
xnor U13511 (N_13511,N_11487,N_10862);
or U13512 (N_13512,N_10301,N_11716);
nor U13513 (N_13513,N_11109,N_11633);
xor U13514 (N_13514,N_11114,N_11860);
xnor U13515 (N_13515,N_10455,N_11917);
nand U13516 (N_13516,N_11554,N_10177);
nor U13517 (N_13517,N_10223,N_10582);
nor U13518 (N_13518,N_11440,N_10376);
and U13519 (N_13519,N_11631,N_10258);
and U13520 (N_13520,N_10051,N_10285);
xor U13521 (N_13521,N_11263,N_10025);
nor U13522 (N_13522,N_11817,N_11883);
and U13523 (N_13523,N_10718,N_11417);
and U13524 (N_13524,N_10217,N_10391);
or U13525 (N_13525,N_10728,N_11652);
nor U13526 (N_13526,N_11898,N_10407);
and U13527 (N_13527,N_11350,N_10117);
and U13528 (N_13528,N_11191,N_10912);
nand U13529 (N_13529,N_10212,N_11846);
and U13530 (N_13530,N_11811,N_11977);
nand U13531 (N_13531,N_11402,N_10826);
xor U13532 (N_13532,N_11284,N_11604);
xor U13533 (N_13533,N_10410,N_11234);
nor U13534 (N_13534,N_10704,N_10255);
or U13535 (N_13535,N_11955,N_11004);
xnor U13536 (N_13536,N_11423,N_11562);
and U13537 (N_13537,N_10893,N_11276);
nor U13538 (N_13538,N_11010,N_11457);
and U13539 (N_13539,N_11898,N_10051);
or U13540 (N_13540,N_10573,N_11846);
nor U13541 (N_13541,N_10835,N_11183);
xor U13542 (N_13542,N_10892,N_11242);
or U13543 (N_13543,N_11622,N_10177);
nor U13544 (N_13544,N_10104,N_10834);
xor U13545 (N_13545,N_10880,N_10125);
xnor U13546 (N_13546,N_10148,N_11127);
and U13547 (N_13547,N_11381,N_10507);
nand U13548 (N_13548,N_10077,N_10835);
xor U13549 (N_13549,N_11138,N_10974);
nand U13550 (N_13550,N_11160,N_10409);
xor U13551 (N_13551,N_10052,N_10263);
or U13552 (N_13552,N_10919,N_10654);
nand U13553 (N_13553,N_10585,N_10102);
or U13554 (N_13554,N_10836,N_11686);
or U13555 (N_13555,N_11203,N_11555);
or U13556 (N_13556,N_10170,N_10762);
or U13557 (N_13557,N_11732,N_10720);
xnor U13558 (N_13558,N_10834,N_11459);
nor U13559 (N_13559,N_11501,N_11443);
and U13560 (N_13560,N_10638,N_10713);
and U13561 (N_13561,N_10094,N_10596);
nand U13562 (N_13562,N_11664,N_10815);
nor U13563 (N_13563,N_10861,N_10918);
xor U13564 (N_13564,N_11171,N_11879);
or U13565 (N_13565,N_11509,N_10932);
nand U13566 (N_13566,N_11040,N_10424);
and U13567 (N_13567,N_11187,N_11909);
and U13568 (N_13568,N_11080,N_10463);
nor U13569 (N_13569,N_11742,N_10399);
and U13570 (N_13570,N_10480,N_11418);
nand U13571 (N_13571,N_11888,N_10273);
or U13572 (N_13572,N_10337,N_11425);
and U13573 (N_13573,N_10965,N_10513);
and U13574 (N_13574,N_11846,N_11388);
and U13575 (N_13575,N_11003,N_10246);
nand U13576 (N_13576,N_10549,N_11398);
or U13577 (N_13577,N_10818,N_11281);
nand U13578 (N_13578,N_11273,N_10007);
nor U13579 (N_13579,N_11070,N_11369);
nand U13580 (N_13580,N_11253,N_11729);
or U13581 (N_13581,N_11711,N_10872);
nand U13582 (N_13582,N_10367,N_11153);
and U13583 (N_13583,N_11568,N_10657);
or U13584 (N_13584,N_10170,N_11761);
and U13585 (N_13585,N_11942,N_11855);
and U13586 (N_13586,N_10326,N_10989);
and U13587 (N_13587,N_11948,N_10200);
and U13588 (N_13588,N_10163,N_10603);
nand U13589 (N_13589,N_10648,N_10714);
nand U13590 (N_13590,N_11775,N_11248);
nor U13591 (N_13591,N_10103,N_11004);
nor U13592 (N_13592,N_11037,N_10511);
and U13593 (N_13593,N_11185,N_11159);
or U13594 (N_13594,N_11673,N_11798);
nor U13595 (N_13595,N_11413,N_11481);
or U13596 (N_13596,N_10723,N_10741);
or U13597 (N_13597,N_10871,N_11928);
or U13598 (N_13598,N_10245,N_10702);
and U13599 (N_13599,N_11726,N_10181);
nor U13600 (N_13600,N_11309,N_10694);
nor U13601 (N_13601,N_11448,N_10599);
or U13602 (N_13602,N_10310,N_11342);
nand U13603 (N_13603,N_11946,N_11844);
xnor U13604 (N_13604,N_11703,N_11600);
or U13605 (N_13605,N_11286,N_10833);
nor U13606 (N_13606,N_10599,N_10992);
nand U13607 (N_13607,N_11492,N_10812);
or U13608 (N_13608,N_10321,N_11285);
nand U13609 (N_13609,N_10829,N_11282);
and U13610 (N_13610,N_11584,N_10075);
nand U13611 (N_13611,N_11898,N_10050);
or U13612 (N_13612,N_10456,N_11743);
xor U13613 (N_13613,N_11100,N_10336);
or U13614 (N_13614,N_10335,N_10689);
or U13615 (N_13615,N_11603,N_11414);
or U13616 (N_13616,N_10646,N_11026);
and U13617 (N_13617,N_11701,N_11155);
nand U13618 (N_13618,N_10722,N_11695);
or U13619 (N_13619,N_10052,N_11116);
and U13620 (N_13620,N_10615,N_11591);
xor U13621 (N_13621,N_10253,N_11349);
or U13622 (N_13622,N_10672,N_11207);
nand U13623 (N_13623,N_10748,N_11355);
nand U13624 (N_13624,N_10551,N_10448);
and U13625 (N_13625,N_10727,N_11416);
nor U13626 (N_13626,N_11667,N_10062);
nand U13627 (N_13627,N_11539,N_10281);
and U13628 (N_13628,N_11608,N_10179);
nor U13629 (N_13629,N_11778,N_10262);
nor U13630 (N_13630,N_10440,N_10898);
xor U13631 (N_13631,N_11984,N_11916);
xnor U13632 (N_13632,N_10119,N_11791);
xor U13633 (N_13633,N_11376,N_10129);
nand U13634 (N_13634,N_11299,N_10680);
nand U13635 (N_13635,N_11019,N_10933);
and U13636 (N_13636,N_11418,N_11110);
xnor U13637 (N_13637,N_10431,N_11064);
and U13638 (N_13638,N_11847,N_10738);
nor U13639 (N_13639,N_11455,N_11037);
xnor U13640 (N_13640,N_11421,N_11069);
nor U13641 (N_13641,N_10777,N_10372);
nor U13642 (N_13642,N_11590,N_10653);
or U13643 (N_13643,N_11641,N_11161);
and U13644 (N_13644,N_11635,N_11374);
xnor U13645 (N_13645,N_11666,N_10803);
and U13646 (N_13646,N_10967,N_11621);
or U13647 (N_13647,N_11191,N_11686);
and U13648 (N_13648,N_11823,N_10504);
nand U13649 (N_13649,N_10852,N_10106);
and U13650 (N_13650,N_11889,N_10732);
or U13651 (N_13651,N_10439,N_11964);
nor U13652 (N_13652,N_10750,N_10404);
or U13653 (N_13653,N_11716,N_10736);
nand U13654 (N_13654,N_11096,N_10440);
nor U13655 (N_13655,N_11354,N_11375);
nor U13656 (N_13656,N_10977,N_10495);
nand U13657 (N_13657,N_11865,N_10354);
or U13658 (N_13658,N_10522,N_10136);
nand U13659 (N_13659,N_10173,N_10098);
and U13660 (N_13660,N_11450,N_11389);
and U13661 (N_13661,N_10615,N_11183);
nand U13662 (N_13662,N_11463,N_10917);
nand U13663 (N_13663,N_11724,N_10812);
nand U13664 (N_13664,N_11378,N_11929);
xnor U13665 (N_13665,N_10095,N_11790);
and U13666 (N_13666,N_11284,N_11111);
and U13667 (N_13667,N_10553,N_11907);
or U13668 (N_13668,N_11910,N_10014);
nor U13669 (N_13669,N_10307,N_11703);
and U13670 (N_13670,N_11462,N_11209);
xor U13671 (N_13671,N_11997,N_11802);
xor U13672 (N_13672,N_11047,N_10940);
xnor U13673 (N_13673,N_10712,N_10207);
or U13674 (N_13674,N_10112,N_11512);
nand U13675 (N_13675,N_10068,N_11374);
or U13676 (N_13676,N_11709,N_10943);
and U13677 (N_13677,N_10321,N_10607);
nand U13678 (N_13678,N_11082,N_11824);
nand U13679 (N_13679,N_10516,N_10220);
nor U13680 (N_13680,N_10610,N_10642);
and U13681 (N_13681,N_11035,N_11104);
and U13682 (N_13682,N_11483,N_10518);
xor U13683 (N_13683,N_10881,N_10236);
xnor U13684 (N_13684,N_11444,N_11330);
nor U13685 (N_13685,N_10688,N_10044);
nand U13686 (N_13686,N_10162,N_10630);
xor U13687 (N_13687,N_11736,N_11310);
nand U13688 (N_13688,N_10474,N_10747);
nand U13689 (N_13689,N_10622,N_11426);
or U13690 (N_13690,N_10351,N_11966);
nor U13691 (N_13691,N_10252,N_11683);
nand U13692 (N_13692,N_11354,N_10779);
and U13693 (N_13693,N_11481,N_11737);
xnor U13694 (N_13694,N_10855,N_10869);
or U13695 (N_13695,N_11322,N_10801);
nor U13696 (N_13696,N_10650,N_11797);
or U13697 (N_13697,N_10679,N_10957);
nand U13698 (N_13698,N_11235,N_10900);
xnor U13699 (N_13699,N_10914,N_10487);
or U13700 (N_13700,N_11065,N_10628);
and U13701 (N_13701,N_10600,N_10567);
or U13702 (N_13702,N_11779,N_10772);
and U13703 (N_13703,N_11590,N_10867);
nor U13704 (N_13704,N_11834,N_11901);
nor U13705 (N_13705,N_11168,N_10467);
and U13706 (N_13706,N_10469,N_10367);
or U13707 (N_13707,N_11525,N_10259);
nor U13708 (N_13708,N_10362,N_10831);
nor U13709 (N_13709,N_11991,N_11156);
or U13710 (N_13710,N_11837,N_10755);
xnor U13711 (N_13711,N_11258,N_11914);
and U13712 (N_13712,N_11217,N_10166);
nor U13713 (N_13713,N_11298,N_10666);
or U13714 (N_13714,N_11588,N_10174);
nor U13715 (N_13715,N_10541,N_11589);
or U13716 (N_13716,N_10161,N_10824);
or U13717 (N_13717,N_11491,N_10597);
xor U13718 (N_13718,N_11070,N_10024);
xor U13719 (N_13719,N_11281,N_10813);
nand U13720 (N_13720,N_11610,N_10660);
nor U13721 (N_13721,N_11165,N_10443);
nand U13722 (N_13722,N_11521,N_10906);
nand U13723 (N_13723,N_10910,N_11043);
xor U13724 (N_13724,N_11303,N_10052);
nor U13725 (N_13725,N_10968,N_11033);
and U13726 (N_13726,N_10964,N_11617);
or U13727 (N_13727,N_10632,N_10055);
xor U13728 (N_13728,N_11527,N_10436);
xor U13729 (N_13729,N_10312,N_10109);
and U13730 (N_13730,N_11213,N_10901);
xor U13731 (N_13731,N_10308,N_10099);
nor U13732 (N_13732,N_10867,N_11157);
nor U13733 (N_13733,N_10569,N_11672);
nand U13734 (N_13734,N_10822,N_11680);
or U13735 (N_13735,N_10601,N_11146);
nand U13736 (N_13736,N_10329,N_11393);
xor U13737 (N_13737,N_11366,N_10968);
nor U13738 (N_13738,N_10376,N_11173);
or U13739 (N_13739,N_11584,N_10231);
or U13740 (N_13740,N_11190,N_10288);
xnor U13741 (N_13741,N_11128,N_10971);
nand U13742 (N_13742,N_11328,N_11390);
and U13743 (N_13743,N_10751,N_11055);
nor U13744 (N_13744,N_10332,N_10053);
nor U13745 (N_13745,N_10702,N_10180);
nor U13746 (N_13746,N_11172,N_11749);
xnor U13747 (N_13747,N_10467,N_10690);
xnor U13748 (N_13748,N_10093,N_11111);
and U13749 (N_13749,N_10810,N_10340);
or U13750 (N_13750,N_11232,N_10949);
or U13751 (N_13751,N_11427,N_11835);
nor U13752 (N_13752,N_11209,N_11808);
xnor U13753 (N_13753,N_11183,N_11330);
and U13754 (N_13754,N_11957,N_10245);
xor U13755 (N_13755,N_11850,N_10277);
and U13756 (N_13756,N_11184,N_11019);
nor U13757 (N_13757,N_10885,N_10859);
xnor U13758 (N_13758,N_10031,N_11484);
nand U13759 (N_13759,N_10801,N_10289);
or U13760 (N_13760,N_10920,N_11240);
nand U13761 (N_13761,N_10664,N_10026);
and U13762 (N_13762,N_11469,N_10002);
nor U13763 (N_13763,N_10399,N_10929);
or U13764 (N_13764,N_11877,N_10740);
and U13765 (N_13765,N_10671,N_11239);
nand U13766 (N_13766,N_10718,N_10317);
xor U13767 (N_13767,N_10417,N_11317);
nor U13768 (N_13768,N_10654,N_10870);
or U13769 (N_13769,N_11890,N_10765);
or U13770 (N_13770,N_10209,N_10054);
or U13771 (N_13771,N_10866,N_11985);
or U13772 (N_13772,N_11560,N_10074);
or U13773 (N_13773,N_11281,N_10530);
nand U13774 (N_13774,N_11174,N_11889);
nor U13775 (N_13775,N_11233,N_10519);
and U13776 (N_13776,N_11937,N_11744);
and U13777 (N_13777,N_11768,N_10636);
nand U13778 (N_13778,N_11495,N_10692);
xor U13779 (N_13779,N_10336,N_11828);
nand U13780 (N_13780,N_10910,N_10552);
and U13781 (N_13781,N_11132,N_11199);
nor U13782 (N_13782,N_11908,N_10234);
or U13783 (N_13783,N_11646,N_11505);
xnor U13784 (N_13784,N_10647,N_10098);
or U13785 (N_13785,N_11110,N_10848);
and U13786 (N_13786,N_10112,N_10102);
xnor U13787 (N_13787,N_10110,N_10472);
or U13788 (N_13788,N_10599,N_11989);
and U13789 (N_13789,N_11994,N_10435);
or U13790 (N_13790,N_11588,N_11426);
xor U13791 (N_13791,N_10648,N_11363);
nor U13792 (N_13792,N_11066,N_11159);
nor U13793 (N_13793,N_10755,N_11522);
xor U13794 (N_13794,N_10758,N_11931);
or U13795 (N_13795,N_10640,N_11420);
xnor U13796 (N_13796,N_10025,N_10338);
nand U13797 (N_13797,N_11640,N_10053);
nand U13798 (N_13798,N_11418,N_11254);
and U13799 (N_13799,N_10785,N_10957);
and U13800 (N_13800,N_10349,N_10724);
xor U13801 (N_13801,N_11813,N_11716);
and U13802 (N_13802,N_11299,N_10200);
nand U13803 (N_13803,N_11888,N_10849);
nor U13804 (N_13804,N_10737,N_11356);
nor U13805 (N_13805,N_11842,N_11831);
and U13806 (N_13806,N_11777,N_11210);
xnor U13807 (N_13807,N_11956,N_11700);
xnor U13808 (N_13808,N_11498,N_11142);
nor U13809 (N_13809,N_11075,N_11529);
nor U13810 (N_13810,N_10863,N_11986);
or U13811 (N_13811,N_11685,N_11052);
nand U13812 (N_13812,N_11818,N_10496);
and U13813 (N_13813,N_11715,N_10781);
or U13814 (N_13814,N_10870,N_10484);
or U13815 (N_13815,N_11376,N_11677);
nor U13816 (N_13816,N_10174,N_11411);
and U13817 (N_13817,N_11506,N_11851);
and U13818 (N_13818,N_10576,N_11380);
nand U13819 (N_13819,N_11162,N_10239);
and U13820 (N_13820,N_11528,N_10217);
nor U13821 (N_13821,N_10211,N_10845);
nand U13822 (N_13822,N_11854,N_10625);
xor U13823 (N_13823,N_11788,N_10450);
nor U13824 (N_13824,N_11146,N_11537);
nor U13825 (N_13825,N_11766,N_10446);
nor U13826 (N_13826,N_10055,N_11893);
and U13827 (N_13827,N_10240,N_10647);
nor U13828 (N_13828,N_10698,N_11533);
nor U13829 (N_13829,N_11754,N_11978);
nor U13830 (N_13830,N_10713,N_11715);
or U13831 (N_13831,N_10989,N_11248);
and U13832 (N_13832,N_11012,N_11715);
and U13833 (N_13833,N_11562,N_11636);
nor U13834 (N_13834,N_10145,N_10019);
and U13835 (N_13835,N_11199,N_10803);
and U13836 (N_13836,N_10937,N_10315);
nor U13837 (N_13837,N_10465,N_10110);
or U13838 (N_13838,N_10343,N_10189);
and U13839 (N_13839,N_10184,N_11867);
or U13840 (N_13840,N_11473,N_10238);
and U13841 (N_13841,N_10548,N_11316);
or U13842 (N_13842,N_11858,N_10420);
xnor U13843 (N_13843,N_11911,N_10464);
or U13844 (N_13844,N_10041,N_11696);
and U13845 (N_13845,N_11479,N_11630);
and U13846 (N_13846,N_11373,N_11038);
nor U13847 (N_13847,N_11634,N_11615);
xnor U13848 (N_13848,N_10217,N_11794);
nand U13849 (N_13849,N_11668,N_10304);
and U13850 (N_13850,N_10070,N_10348);
or U13851 (N_13851,N_11606,N_10797);
nand U13852 (N_13852,N_11916,N_10563);
xor U13853 (N_13853,N_11050,N_10054);
nor U13854 (N_13854,N_10062,N_11969);
and U13855 (N_13855,N_10917,N_11051);
nand U13856 (N_13856,N_11876,N_10991);
and U13857 (N_13857,N_11582,N_10552);
nand U13858 (N_13858,N_11313,N_11102);
xor U13859 (N_13859,N_10818,N_10559);
nand U13860 (N_13860,N_11888,N_11192);
and U13861 (N_13861,N_10679,N_11026);
and U13862 (N_13862,N_11981,N_11192);
nand U13863 (N_13863,N_10064,N_10718);
xnor U13864 (N_13864,N_11872,N_10905);
or U13865 (N_13865,N_10738,N_11335);
nor U13866 (N_13866,N_11320,N_11139);
and U13867 (N_13867,N_10201,N_10164);
nor U13868 (N_13868,N_11027,N_10820);
nor U13869 (N_13869,N_11762,N_10256);
xnor U13870 (N_13870,N_10774,N_10737);
xor U13871 (N_13871,N_11860,N_11775);
xor U13872 (N_13872,N_11099,N_10272);
and U13873 (N_13873,N_10904,N_11604);
nand U13874 (N_13874,N_11143,N_10193);
xor U13875 (N_13875,N_11578,N_10816);
nor U13876 (N_13876,N_11294,N_10318);
xor U13877 (N_13877,N_10878,N_11847);
xnor U13878 (N_13878,N_10038,N_11585);
and U13879 (N_13879,N_11721,N_10786);
xnor U13880 (N_13880,N_11124,N_10330);
nor U13881 (N_13881,N_10394,N_11752);
and U13882 (N_13882,N_11922,N_11689);
nor U13883 (N_13883,N_10040,N_10800);
nor U13884 (N_13884,N_11660,N_11041);
nand U13885 (N_13885,N_11482,N_11307);
or U13886 (N_13886,N_11002,N_11260);
xnor U13887 (N_13887,N_10323,N_11427);
and U13888 (N_13888,N_11782,N_11212);
xnor U13889 (N_13889,N_10989,N_11180);
and U13890 (N_13890,N_11642,N_11734);
nor U13891 (N_13891,N_11241,N_10692);
nand U13892 (N_13892,N_11437,N_11421);
xnor U13893 (N_13893,N_11259,N_11864);
and U13894 (N_13894,N_11241,N_11369);
and U13895 (N_13895,N_10724,N_11378);
nand U13896 (N_13896,N_10641,N_11373);
xnor U13897 (N_13897,N_11213,N_10368);
nor U13898 (N_13898,N_11631,N_10959);
or U13899 (N_13899,N_10890,N_10119);
nor U13900 (N_13900,N_11523,N_10599);
and U13901 (N_13901,N_10348,N_10260);
xor U13902 (N_13902,N_11899,N_10714);
or U13903 (N_13903,N_10371,N_10912);
and U13904 (N_13904,N_11148,N_11131);
or U13905 (N_13905,N_10163,N_11365);
xor U13906 (N_13906,N_10756,N_10127);
nand U13907 (N_13907,N_11126,N_10772);
and U13908 (N_13908,N_10098,N_10902);
or U13909 (N_13909,N_10238,N_11734);
xnor U13910 (N_13910,N_10839,N_11126);
xnor U13911 (N_13911,N_10430,N_11455);
and U13912 (N_13912,N_10297,N_11282);
nor U13913 (N_13913,N_10646,N_11476);
and U13914 (N_13914,N_11080,N_11294);
or U13915 (N_13915,N_10852,N_11263);
nor U13916 (N_13916,N_11108,N_10115);
and U13917 (N_13917,N_11431,N_10065);
or U13918 (N_13918,N_10243,N_11698);
nor U13919 (N_13919,N_10222,N_11138);
nor U13920 (N_13920,N_10668,N_11708);
and U13921 (N_13921,N_11347,N_11075);
nand U13922 (N_13922,N_11956,N_10529);
and U13923 (N_13923,N_11020,N_10717);
nand U13924 (N_13924,N_10431,N_10553);
or U13925 (N_13925,N_11191,N_11967);
xor U13926 (N_13926,N_11784,N_11228);
and U13927 (N_13927,N_10344,N_11294);
and U13928 (N_13928,N_10396,N_10585);
nor U13929 (N_13929,N_10200,N_10316);
and U13930 (N_13930,N_11033,N_11161);
nand U13931 (N_13931,N_11271,N_11596);
and U13932 (N_13932,N_10862,N_11627);
or U13933 (N_13933,N_11789,N_10383);
or U13934 (N_13934,N_10565,N_11905);
xnor U13935 (N_13935,N_10839,N_11572);
nor U13936 (N_13936,N_11003,N_10358);
and U13937 (N_13937,N_10660,N_11346);
or U13938 (N_13938,N_11089,N_10831);
nand U13939 (N_13939,N_11130,N_11215);
or U13940 (N_13940,N_11001,N_10423);
nor U13941 (N_13941,N_10864,N_11598);
or U13942 (N_13942,N_11818,N_10952);
and U13943 (N_13943,N_10474,N_11589);
nor U13944 (N_13944,N_10616,N_11639);
nor U13945 (N_13945,N_11076,N_10789);
xor U13946 (N_13946,N_10846,N_11384);
and U13947 (N_13947,N_10839,N_10959);
or U13948 (N_13948,N_11010,N_10518);
and U13949 (N_13949,N_10042,N_11443);
nand U13950 (N_13950,N_11948,N_10514);
nor U13951 (N_13951,N_10599,N_10506);
and U13952 (N_13952,N_11161,N_11740);
or U13953 (N_13953,N_10666,N_10047);
xnor U13954 (N_13954,N_11447,N_11876);
nand U13955 (N_13955,N_11375,N_11680);
nor U13956 (N_13956,N_10834,N_10452);
and U13957 (N_13957,N_11946,N_10983);
nor U13958 (N_13958,N_11008,N_11621);
nor U13959 (N_13959,N_11530,N_10084);
nand U13960 (N_13960,N_11886,N_11857);
nand U13961 (N_13961,N_11345,N_10842);
nand U13962 (N_13962,N_11656,N_11467);
xor U13963 (N_13963,N_11449,N_10331);
nand U13964 (N_13964,N_11693,N_10205);
xor U13965 (N_13965,N_11147,N_11467);
xor U13966 (N_13966,N_10382,N_10873);
or U13967 (N_13967,N_10225,N_11490);
and U13968 (N_13968,N_11065,N_11373);
xor U13969 (N_13969,N_10193,N_10447);
or U13970 (N_13970,N_10904,N_11620);
or U13971 (N_13971,N_10396,N_11009);
nor U13972 (N_13972,N_10995,N_10828);
and U13973 (N_13973,N_10338,N_11308);
nor U13974 (N_13974,N_10304,N_11083);
xnor U13975 (N_13975,N_11850,N_10328);
xor U13976 (N_13976,N_10503,N_11737);
or U13977 (N_13977,N_11183,N_11982);
xor U13978 (N_13978,N_10962,N_11814);
or U13979 (N_13979,N_11316,N_11540);
xnor U13980 (N_13980,N_10218,N_11797);
xnor U13981 (N_13981,N_10252,N_10274);
or U13982 (N_13982,N_10266,N_10993);
xnor U13983 (N_13983,N_10801,N_11952);
nor U13984 (N_13984,N_11031,N_11380);
nor U13985 (N_13985,N_11739,N_10473);
and U13986 (N_13986,N_10235,N_10472);
xor U13987 (N_13987,N_11826,N_11885);
or U13988 (N_13988,N_10207,N_10506);
or U13989 (N_13989,N_10363,N_11243);
xor U13990 (N_13990,N_10130,N_11829);
and U13991 (N_13991,N_10381,N_10514);
nand U13992 (N_13992,N_11893,N_11366);
and U13993 (N_13993,N_11188,N_11194);
or U13994 (N_13994,N_11265,N_11179);
and U13995 (N_13995,N_11854,N_11399);
or U13996 (N_13996,N_10862,N_11727);
or U13997 (N_13997,N_11484,N_10347);
nand U13998 (N_13998,N_10396,N_10752);
and U13999 (N_13999,N_11078,N_10132);
xor U14000 (N_14000,N_13978,N_12134);
and U14001 (N_14001,N_13801,N_12319);
or U14002 (N_14002,N_12784,N_12282);
nor U14003 (N_14003,N_12076,N_12079);
or U14004 (N_14004,N_12305,N_12202);
or U14005 (N_14005,N_12201,N_12107);
or U14006 (N_14006,N_12336,N_13662);
xnor U14007 (N_14007,N_12140,N_13555);
and U14008 (N_14008,N_13982,N_13397);
and U14009 (N_14009,N_12346,N_12944);
nor U14010 (N_14010,N_12804,N_12169);
nand U14011 (N_14011,N_12837,N_13847);
or U14012 (N_14012,N_13696,N_13528);
nor U14013 (N_14013,N_13332,N_13558);
nand U14014 (N_14014,N_13326,N_13583);
nand U14015 (N_14015,N_13330,N_12936);
nand U14016 (N_14016,N_13607,N_13349);
and U14017 (N_14017,N_13041,N_12329);
nand U14018 (N_14018,N_12602,N_13989);
nand U14019 (N_14019,N_12137,N_12953);
nand U14020 (N_14020,N_13814,N_12779);
or U14021 (N_14021,N_13757,N_12309);
xnor U14022 (N_14022,N_12586,N_12067);
nand U14023 (N_14023,N_12218,N_13712);
and U14024 (N_14024,N_13535,N_12177);
and U14025 (N_14025,N_12019,N_12776);
xnor U14026 (N_14026,N_13548,N_13911);
or U14027 (N_14027,N_13632,N_12046);
nand U14028 (N_14028,N_13896,N_13722);
xnor U14029 (N_14029,N_13087,N_12184);
nand U14030 (N_14030,N_12334,N_12517);
and U14031 (N_14031,N_13432,N_13043);
nand U14032 (N_14032,N_13078,N_12012);
nand U14033 (N_14033,N_13142,N_12082);
or U14034 (N_14034,N_13199,N_13498);
nor U14035 (N_14035,N_13366,N_12750);
and U14036 (N_14036,N_13539,N_12498);
nor U14037 (N_14037,N_12916,N_12131);
or U14038 (N_14038,N_13953,N_12527);
nor U14039 (N_14039,N_12114,N_13151);
xnor U14040 (N_14040,N_13540,N_13772);
xor U14041 (N_14041,N_13530,N_13994);
nand U14042 (N_14042,N_12490,N_12760);
nor U14043 (N_14043,N_13392,N_12627);
nand U14044 (N_14044,N_12644,N_13123);
and U14045 (N_14045,N_13531,N_12382);
xnor U14046 (N_14046,N_13179,N_13709);
nor U14047 (N_14047,N_13054,N_12203);
and U14048 (N_14048,N_13538,N_13117);
xnor U14049 (N_14049,N_13973,N_12731);
nor U14050 (N_14050,N_12905,N_12587);
or U14051 (N_14051,N_12959,N_13479);
nand U14052 (N_14052,N_13158,N_12600);
and U14053 (N_14053,N_12249,N_12962);
or U14054 (N_14054,N_12590,N_12833);
and U14055 (N_14055,N_12207,N_12118);
nand U14056 (N_14056,N_13003,N_12073);
nor U14057 (N_14057,N_12027,N_13287);
nand U14058 (N_14058,N_13312,N_12482);
nand U14059 (N_14059,N_13371,N_12084);
nor U14060 (N_14060,N_13324,N_12990);
nor U14061 (N_14061,N_12420,N_12443);
or U14062 (N_14062,N_13972,N_12045);
or U14063 (N_14063,N_13520,N_13616);
xor U14064 (N_14064,N_12754,N_13372);
and U14065 (N_14065,N_12033,N_12466);
xor U14066 (N_14066,N_12967,N_13603);
nand U14067 (N_14067,N_12630,N_12465);
xnor U14068 (N_14068,N_12263,N_13950);
or U14069 (N_14069,N_13033,N_13170);
nor U14070 (N_14070,N_12922,N_13282);
or U14071 (N_14071,N_12846,N_13215);
nand U14072 (N_14072,N_13737,N_12687);
nor U14073 (N_14073,N_13610,N_12771);
xnor U14074 (N_14074,N_13387,N_12455);
nor U14075 (N_14075,N_12402,N_13898);
nor U14076 (N_14076,N_13309,N_12987);
xnor U14077 (N_14077,N_13321,N_12564);
xnor U14078 (N_14078,N_12255,N_13850);
nand U14079 (N_14079,N_12597,N_13466);
xnor U14080 (N_14080,N_12742,N_13651);
xnor U14081 (N_14081,N_13820,N_12688);
nor U14082 (N_14082,N_12505,N_13723);
or U14083 (N_14083,N_13979,N_12631);
and U14084 (N_14084,N_13486,N_13654);
xor U14085 (N_14085,N_13985,N_12938);
or U14086 (N_14086,N_13034,N_12599);
xor U14087 (N_14087,N_13475,N_12237);
nand U14088 (N_14088,N_12499,N_12277);
nand U14089 (N_14089,N_12749,N_12926);
or U14090 (N_14090,N_13005,N_12244);
nand U14091 (N_14091,N_13529,N_12328);
and U14092 (N_14092,N_12349,N_13146);
or U14093 (N_14093,N_13104,N_13881);
and U14094 (N_14094,N_12040,N_12311);
nor U14095 (N_14095,N_13909,N_12875);
or U14096 (N_14096,N_13629,N_13788);
nand U14097 (N_14097,N_12350,N_12735);
nand U14098 (N_14098,N_13537,N_12380);
or U14099 (N_14099,N_13357,N_13437);
xor U14100 (N_14100,N_12185,N_13344);
nand U14101 (N_14101,N_13490,N_12512);
nand U14102 (N_14102,N_12072,N_12155);
or U14103 (N_14103,N_12874,N_13243);
xor U14104 (N_14104,N_13298,N_12321);
nor U14105 (N_14105,N_12999,N_12819);
or U14106 (N_14106,N_12813,N_12643);
nor U14107 (N_14107,N_13731,N_12619);
nor U14108 (N_14108,N_12325,N_12717);
xor U14109 (N_14109,N_13351,N_13506);
and U14110 (N_14110,N_13557,N_13415);
nand U14111 (N_14111,N_13811,N_12224);
nor U14112 (N_14112,N_12622,N_12909);
or U14113 (N_14113,N_12852,N_13461);
xor U14114 (N_14114,N_12370,N_13252);
and U14115 (N_14115,N_12421,N_12092);
nor U14116 (N_14116,N_13792,N_12091);
xor U14117 (N_14117,N_13345,N_13889);
xor U14118 (N_14118,N_13083,N_13921);
nand U14119 (N_14119,N_12149,N_12032);
nand U14120 (N_14120,N_13864,N_13517);
and U14121 (N_14121,N_12411,N_12474);
and U14122 (N_14122,N_12727,N_13133);
nand U14123 (N_14123,N_12009,N_12522);
xnor U14124 (N_14124,N_12920,N_13956);
or U14125 (N_14125,N_13325,N_12154);
and U14126 (N_14126,N_13114,N_12457);
xor U14127 (N_14127,N_13752,N_13334);
and U14128 (N_14128,N_13231,N_12947);
and U14129 (N_14129,N_13477,N_12553);
nor U14130 (N_14130,N_13768,N_12887);
or U14131 (N_14131,N_12121,N_13706);
nand U14132 (N_14132,N_12354,N_12550);
nand U14133 (N_14133,N_12842,N_13892);
xor U14134 (N_14134,N_13927,N_13077);
and U14135 (N_14135,N_13789,N_13617);
nor U14136 (N_14136,N_13627,N_12798);
and U14137 (N_14137,N_12811,N_12437);
nor U14138 (N_14138,N_12188,N_13521);
xnor U14139 (N_14139,N_13804,N_13882);
and U14140 (N_14140,N_12528,N_12348);
and U14141 (N_14141,N_12608,N_13377);
nand U14142 (N_14142,N_13389,N_12398);
nand U14143 (N_14143,N_12623,N_13150);
and U14144 (N_14144,N_12005,N_13713);
and U14145 (N_14145,N_13840,N_13379);
or U14146 (N_14146,N_13758,N_13181);
nor U14147 (N_14147,N_12106,N_12954);
and U14148 (N_14148,N_13667,N_12678);
nand U14149 (N_14149,N_12693,N_13605);
or U14150 (N_14150,N_13522,N_12200);
xor U14151 (N_14151,N_13888,N_13944);
nand U14152 (N_14152,N_13541,N_12649);
nand U14153 (N_14153,N_13549,N_12486);
and U14154 (N_14154,N_12089,N_12790);
nor U14155 (N_14155,N_12476,N_13575);
xor U14156 (N_14156,N_13405,N_13593);
nor U14157 (N_14157,N_12662,N_12931);
or U14158 (N_14158,N_13813,N_13621);
nor U14159 (N_14159,N_12043,N_12062);
and U14160 (N_14160,N_12880,N_12379);
or U14161 (N_14161,N_13842,N_12980);
or U14162 (N_14162,N_12573,N_12217);
nand U14163 (N_14163,N_13070,N_12275);
nor U14164 (N_14164,N_13701,N_12971);
and U14165 (N_14165,N_12316,N_13863);
nor U14166 (N_14166,N_12123,N_13987);
nand U14167 (N_14167,N_12740,N_12101);
and U14168 (N_14168,N_12044,N_12481);
or U14169 (N_14169,N_12889,N_12775);
or U14170 (N_14170,N_13428,N_13496);
or U14171 (N_14171,N_12552,N_12291);
or U14172 (N_14172,N_13843,N_13218);
and U14173 (N_14173,N_12708,N_13419);
or U14174 (N_14174,N_13767,N_12637);
xnor U14175 (N_14175,N_12502,N_13481);
and U14176 (N_14176,N_12042,N_12489);
and U14177 (N_14177,N_12758,N_13986);
nand U14178 (N_14178,N_13472,N_13659);
xnor U14179 (N_14179,N_13431,N_13128);
nor U14180 (N_14180,N_13578,N_13217);
or U14181 (N_14181,N_13093,N_13519);
xor U14182 (N_14182,N_12356,N_12341);
nor U14183 (N_14183,N_13550,N_13364);
or U14184 (N_14184,N_13076,N_12215);
xor U14185 (N_14185,N_13444,N_13849);
and U14186 (N_14186,N_13665,N_13905);
nand U14187 (N_14187,N_13410,N_13203);
nand U14188 (N_14188,N_13229,N_12707);
nor U14189 (N_14189,N_13119,N_13178);
and U14190 (N_14190,N_12709,N_12054);
or U14191 (N_14191,N_13715,N_12585);
and U14192 (N_14192,N_12322,N_13977);
xor U14193 (N_14193,N_12095,N_13173);
or U14194 (N_14194,N_13141,N_13676);
or U14195 (N_14195,N_12229,N_13042);
xnor U14196 (N_14196,N_13048,N_12447);
nor U14197 (N_14197,N_13658,N_12533);
nor U14198 (N_14198,N_13590,N_12178);
nand U14199 (N_14199,N_13725,N_12763);
or U14200 (N_14200,N_12911,N_13716);
xnor U14201 (N_14201,N_12087,N_12407);
or U14202 (N_14202,N_13805,N_13851);
xor U14203 (N_14203,N_12960,N_13500);
nand U14204 (N_14204,N_13401,N_13859);
nand U14205 (N_14205,N_13099,N_13028);
nor U14206 (N_14206,N_13436,N_13495);
or U14207 (N_14207,N_12615,N_13525);
xnor U14208 (N_14208,N_13560,N_13124);
nand U14209 (N_14209,N_12344,N_13105);
nor U14210 (N_14210,N_13259,N_12259);
xor U14211 (N_14211,N_13571,N_12061);
nor U14212 (N_14212,N_13641,N_13081);
nand U14213 (N_14213,N_13206,N_13049);
and U14214 (N_14214,N_12471,N_13245);
or U14215 (N_14215,N_13013,N_12239);
nand U14216 (N_14216,N_13682,N_13680);
or U14217 (N_14217,N_12272,N_12598);
and U14218 (N_14218,N_13228,N_12901);
nor U14219 (N_14219,N_12351,N_13524);
and U14220 (N_14220,N_13726,N_12741);
nand U14221 (N_14221,N_12878,N_12940);
nand U14222 (N_14222,N_12186,N_13802);
nor U14223 (N_14223,N_13899,N_13009);
and U14224 (N_14224,N_13289,N_13579);
xor U14225 (N_14225,N_12633,N_12994);
and U14226 (N_14226,N_12016,N_13413);
or U14227 (N_14227,N_13239,N_12614);
xnor U14228 (N_14228,N_12289,N_12732);
nor U14229 (N_14229,N_12983,N_13272);
nand U14230 (N_14230,N_13305,N_13692);
nand U14231 (N_14231,N_12985,N_12231);
or U14232 (N_14232,N_13942,N_12514);
nand U14233 (N_14233,N_13396,N_13702);
nor U14234 (N_14234,N_12803,N_13266);
and U14235 (N_14235,N_12260,N_13363);
nand U14236 (N_14236,N_12523,N_13748);
xnor U14237 (N_14237,N_13169,N_12559);
xnor U14238 (N_14238,N_12392,N_12904);
nand U14239 (N_14239,N_13816,N_13232);
nand U14240 (N_14240,N_12831,N_12330);
xnor U14241 (N_14241,N_12252,N_12782);
and U14242 (N_14242,N_13144,N_12570);
xor U14243 (N_14243,N_13573,N_13874);
nand U14244 (N_14244,N_12069,N_12176);
or U14245 (N_14245,N_13137,N_13168);
and U14246 (N_14246,N_13580,N_13202);
nand U14247 (N_14247,N_12870,N_13071);
or U14248 (N_14248,N_13824,N_13399);
and U14249 (N_14249,N_13800,N_13102);
nor U14250 (N_14250,N_12098,N_13753);
xnor U14251 (N_14251,N_12978,N_13817);
nor U14252 (N_14252,N_12766,N_12205);
nor U14253 (N_14253,N_12925,N_12433);
nor U14254 (N_14254,N_12400,N_13876);
xor U14255 (N_14255,N_13335,N_12128);
xnor U14256 (N_14256,N_13165,N_13314);
or U14257 (N_14257,N_12795,N_12171);
nand U14258 (N_14258,N_13039,N_13599);
xnor U14259 (N_14259,N_13000,N_13318);
and U14260 (N_14260,N_13462,N_13831);
and U14261 (N_14261,N_13201,N_13191);
and U14262 (N_14262,N_13965,N_13559);
or U14263 (N_14263,N_13582,N_12737);
nand U14264 (N_14264,N_13255,N_13683);
or U14265 (N_14265,N_12562,N_12891);
xor U14266 (N_14266,N_13294,N_12666);
and U14267 (N_14267,N_12770,N_13106);
xnor U14268 (N_14268,N_12966,N_13148);
or U14269 (N_14269,N_13354,N_12792);
or U14270 (N_14270,N_12669,N_12712);
nand U14271 (N_14271,N_12315,N_13090);
nand U14272 (N_14272,N_13836,N_13235);
xor U14273 (N_14273,N_13194,N_12247);
nor U14274 (N_14274,N_13685,N_13670);
and U14275 (N_14275,N_12996,N_13742);
or U14276 (N_14276,N_12450,N_13027);
nor U14277 (N_14277,N_13422,N_13210);
xor U14278 (N_14278,N_13200,N_12357);
xor U14279 (N_14279,N_13552,N_13058);
nand U14280 (N_14280,N_13834,N_13380);
nor U14281 (N_14281,N_13618,N_13101);
and U14282 (N_14282,N_13736,N_13935);
or U14283 (N_14283,N_12789,N_12163);
nand U14284 (N_14284,N_13474,N_12416);
nand U14285 (N_14285,N_13333,N_13853);
nor U14286 (N_14286,N_12968,N_13807);
xor U14287 (N_14287,N_13516,N_12204);
or U14288 (N_14288,N_12725,N_12338);
xnor U14289 (N_14289,N_13400,N_13771);
or U14290 (N_14290,N_13435,N_13016);
xor U14291 (N_14291,N_13342,N_12172);
nand U14292 (N_14292,N_12537,N_12057);
nor U14293 (N_14293,N_13417,N_12817);
xor U14294 (N_14294,N_13187,N_12526);
nand U14295 (N_14295,N_12501,N_13446);
or U14296 (N_14296,N_12897,N_13916);
nand U14297 (N_14297,N_12521,N_13854);
or U14298 (N_14298,N_13460,N_12663);
xor U14299 (N_14299,N_13769,N_13830);
nor U14300 (N_14300,N_12679,N_12461);
nand U14301 (N_14301,N_13955,N_12406);
xor U14302 (N_14302,N_12074,N_12093);
nor U14303 (N_14303,N_12028,N_12273);
or U14304 (N_14304,N_12892,N_13910);
xor U14305 (N_14305,N_12838,N_13361);
xor U14306 (N_14306,N_12504,N_12757);
nor U14307 (N_14307,N_13328,N_12661);
or U14308 (N_14308,N_12561,N_13125);
xor U14309 (N_14309,N_13553,N_13221);
or U14310 (N_14310,N_12697,N_12367);
nor U14311 (N_14311,N_12848,N_12135);
nand U14312 (N_14312,N_12815,N_12997);
xnor U14313 (N_14313,N_13852,N_13393);
nor U14314 (N_14314,N_13595,N_13732);
xnor U14315 (N_14315,N_13046,N_13728);
or U14316 (N_14316,N_13508,N_13694);
and U14317 (N_14317,N_13832,N_13609);
nor U14318 (N_14318,N_13086,N_12657);
nor U14319 (N_14319,N_13798,N_12377);
xor U14320 (N_14320,N_13420,N_12306);
or U14321 (N_14321,N_12146,N_13269);
nor U14322 (N_14322,N_12167,N_12964);
xnor U14323 (N_14323,N_13409,N_13080);
and U14324 (N_14324,N_12744,N_12442);
nor U14325 (N_14325,N_13708,N_13063);
or U14326 (N_14326,N_12584,N_12048);
and U14327 (N_14327,N_12013,N_12793);
or U14328 (N_14328,N_13275,N_13035);
xor U14329 (N_14329,N_12518,N_13988);
nor U14330 (N_14330,N_13633,N_12935);
nand U14331 (N_14331,N_13711,N_12108);
or U14332 (N_14332,N_13004,N_13310);
nand U14333 (N_14333,N_12112,N_12122);
and U14334 (N_14334,N_12414,N_12410);
xor U14335 (N_14335,N_12100,N_12762);
nand U14336 (N_14336,N_12068,N_12371);
nor U14337 (N_14337,N_13126,N_13710);
or U14338 (N_14338,N_13299,N_13597);
or U14339 (N_14339,N_13780,N_12826);
or U14340 (N_14340,N_12243,N_12460);
nor U14341 (N_14341,N_12799,N_12908);
and U14342 (N_14342,N_12153,N_13390);
or U14343 (N_14343,N_12132,N_13554);
nor U14344 (N_14344,N_12448,N_13879);
or U14345 (N_14345,N_13964,N_12064);
or U14346 (N_14346,N_13268,N_12543);
nor U14347 (N_14347,N_13626,N_12943);
and U14348 (N_14348,N_12660,N_13643);
and U14349 (N_14349,N_13196,N_13439);
nor U14350 (N_14350,N_13515,N_12434);
nand U14351 (N_14351,N_12475,N_12182);
or U14352 (N_14352,N_12384,N_12147);
and U14353 (N_14353,N_13503,N_12110);
xnor U14354 (N_14354,N_13285,N_13613);
nand U14355 (N_14355,N_13073,N_12656);
xor U14356 (N_14356,N_12360,N_13329);
xnor U14357 (N_14357,N_12119,N_13880);
nor U14358 (N_14358,N_13796,N_13047);
or U14359 (N_14359,N_13295,N_13040);
nand U14360 (N_14360,N_13205,N_12796);
or U14361 (N_14361,N_12729,N_12293);
and U14362 (N_14362,N_12839,N_12393);
or U14363 (N_14363,N_13457,N_13327);
or U14364 (N_14364,N_13652,N_13981);
xnor U14365 (N_14365,N_12668,N_13250);
xor U14366 (N_14366,N_12814,N_13190);
nand U14367 (N_14367,N_12748,N_13029);
or U14368 (N_14368,N_13374,N_13384);
xor U14369 (N_14369,N_12756,N_12834);
or U14370 (N_14370,N_13724,N_13068);
and U14371 (N_14371,N_12853,N_13739);
nor U14372 (N_14372,N_12212,N_12444);
nor U14373 (N_14373,N_12365,N_13877);
nor U14374 (N_14374,N_12432,N_13219);
and U14375 (N_14375,N_12036,N_13302);
nand U14376 (N_14376,N_13214,N_13693);
xor U14377 (N_14377,N_13958,N_12594);
xor U14378 (N_14378,N_12209,N_12609);
nor U14379 (N_14379,N_13208,N_13565);
nor U14380 (N_14380,N_13793,N_12075);
nand U14381 (N_14381,N_12047,N_12423);
or U14382 (N_14382,N_13216,N_12720);
or U14383 (N_14383,N_12820,N_13720);
nor U14384 (N_14384,N_13037,N_13307);
or U14385 (N_14385,N_13969,N_12919);
nand U14386 (N_14386,N_13904,N_12066);
xor U14387 (N_14387,N_12428,N_13476);
nand U14388 (N_14388,N_13425,N_13167);
xor U14389 (N_14389,N_13222,N_13097);
nor U14390 (N_14390,N_12917,N_13154);
or U14391 (N_14391,N_13267,N_12713);
xnor U14392 (N_14392,N_13404,N_12109);
or U14393 (N_14393,N_12438,N_12928);
nand U14394 (N_14394,N_12618,N_13300);
xor U14395 (N_14395,N_13060,N_13441);
or U14396 (N_14396,N_13795,N_13963);
and U14397 (N_14397,N_12366,N_12507);
or U14398 (N_14398,N_12519,N_13913);
xnor U14399 (N_14399,N_13402,N_13092);
xnor U14400 (N_14400,N_12056,N_13934);
nand U14401 (N_14401,N_13572,N_12722);
or U14402 (N_14402,N_13499,N_12183);
or U14403 (N_14403,N_13587,N_12358);
nand U14404 (N_14404,N_13543,N_12752);
nand U14405 (N_14405,N_12284,N_13601);
and U14406 (N_14406,N_12548,N_12927);
or U14407 (N_14407,N_13943,N_13829);
nor U14408 (N_14408,N_13427,N_13248);
and U14409 (N_14409,N_12648,N_13929);
or U14410 (N_14410,N_12187,N_12989);
nor U14411 (N_14411,N_12477,N_12099);
nor U14412 (N_14412,N_13338,N_12642);
nand U14413 (N_14413,N_12018,N_12710);
nor U14414 (N_14414,N_12234,N_13075);
and U14415 (N_14415,N_12164,N_12781);
and U14416 (N_14416,N_13017,N_13118);
or U14417 (N_14417,N_12680,N_13906);
nor U14418 (N_14418,N_13765,N_13823);
nand U14419 (N_14419,N_12422,N_13395);
nand U14420 (N_14420,N_12923,N_13962);
or U14421 (N_14421,N_13391,N_13251);
nand U14422 (N_14422,N_13264,N_13738);
or U14423 (N_14423,N_12847,N_13429);
nor U14424 (N_14424,N_13244,N_12213);
xnor U14425 (N_14425,N_13131,N_12190);
or U14426 (N_14426,N_12385,N_13501);
and U14427 (N_14427,N_13866,N_13747);
nand U14428 (N_14428,N_13976,N_13233);
nor U14429 (N_14429,N_12791,N_12454);
nor U14430 (N_14430,N_12483,N_12439);
and U14431 (N_14431,N_13157,N_13564);
xor U14432 (N_14432,N_13908,N_12478);
xnor U14433 (N_14433,N_12413,N_13642);
and U14434 (N_14434,N_12802,N_13514);
and U14435 (N_14435,N_13954,N_13727);
xor U14436 (N_14436,N_13611,N_12280);
and U14437 (N_14437,N_12885,N_12684);
and U14438 (N_14438,N_13172,N_12105);
nor U14439 (N_14439,N_12686,N_13821);
and U14440 (N_14440,N_12773,N_13630);
nor U14441 (N_14441,N_12716,N_12787);
and U14442 (N_14442,N_13261,N_13375);
xnor U14443 (N_14443,N_13975,N_13108);
xor U14444 (N_14444,N_12011,N_12287);
nor U14445 (N_14445,N_13782,N_13007);
xnor U14446 (N_14446,N_12138,N_13115);
nand U14447 (N_14447,N_13766,N_12806);
or U14448 (N_14448,N_13220,N_12397);
nand U14449 (N_14449,N_13143,N_13209);
xor U14450 (N_14450,N_12298,N_12863);
xnor U14451 (N_14451,N_12728,N_12557);
and U14452 (N_14452,N_13822,N_13127);
xnor U14453 (N_14453,N_13370,N_12540);
xnor U14454 (N_14454,N_12854,N_13337);
and U14455 (N_14455,N_13797,N_13835);
or U14456 (N_14456,N_13140,N_13411);
nand U14457 (N_14457,N_13511,N_13421);
nand U14458 (N_14458,N_13922,N_12524);
xor U14459 (N_14459,N_12331,N_13171);
nand U14460 (N_14460,N_12596,N_12362);
nand U14461 (N_14461,N_12788,N_12085);
xor U14462 (N_14462,N_13991,N_12473);
and U14463 (N_14463,N_12672,N_13585);
xor U14464 (N_14464,N_12628,N_12025);
or U14465 (N_14465,N_12823,N_12934);
nand U14466 (N_14466,N_12391,N_13914);
and U14467 (N_14467,N_12015,N_12228);
nand U14468 (N_14468,N_12801,N_12952);
and U14469 (N_14469,N_12638,N_12440);
or U14470 (N_14470,N_13438,N_12001);
and U14471 (N_14471,N_12060,N_12671);
and U14472 (N_14472,N_12950,N_12038);
xnor U14473 (N_14473,N_13576,N_12577);
or U14474 (N_14474,N_12867,N_12446);
and U14475 (N_14475,N_12877,N_13038);
or U14476 (N_14476,N_12453,N_12431);
xnor U14477 (N_14477,N_12975,N_13050);
xor U14478 (N_14478,N_13939,N_12408);
nor U14479 (N_14479,N_13414,N_13920);
nor U14480 (N_14480,N_12857,N_13980);
nand U14481 (N_14481,N_13925,N_13542);
nand U14482 (N_14482,N_13584,N_13699);
xor U14483 (N_14483,N_13669,N_13290);
xor U14484 (N_14484,N_13620,N_13177);
nor U14485 (N_14485,N_13504,N_13674);
xnor U14486 (N_14486,N_13453,N_13488);
and U14487 (N_14487,N_13403,N_13907);
or U14488 (N_14488,N_12462,N_13074);
nor U14489 (N_14489,N_12583,N_12858);
xor U14490 (N_14490,N_13089,N_13900);
and U14491 (N_14491,N_13808,N_13998);
and U14492 (N_14492,N_13452,N_12246);
and U14493 (N_14493,N_12719,N_13455);
xnor U14494 (N_14494,N_13188,N_12267);
or U14495 (N_14495,N_12565,N_13717);
or U14496 (N_14496,N_12851,N_13871);
nand U14497 (N_14497,N_13577,N_12957);
nand U14498 (N_14498,N_12174,N_13803);
xnor U14499 (N_14499,N_12900,N_13376);
or U14500 (N_14500,N_12250,N_12222);
xor U14501 (N_14501,N_13163,N_12353);
and U14502 (N_14502,N_12472,N_13442);
nor U14503 (N_14503,N_13084,N_12401);
nor U14504 (N_14504,N_13263,N_12278);
nor U14505 (N_14505,N_13303,N_13993);
nor U14506 (N_14506,N_13271,N_12743);
xnor U14507 (N_14507,N_12861,N_13164);
or U14508 (N_14508,N_12601,N_13113);
and U14509 (N_14509,N_13598,N_12828);
and U14510 (N_14510,N_12242,N_13509);
xnor U14511 (N_14511,N_13489,N_12097);
xnor U14512 (N_14512,N_13968,N_13751);
nor U14513 (N_14513,N_12865,N_12469);
xor U14514 (N_14514,N_12078,N_12302);
and U14515 (N_14515,N_13828,N_13469);
and U14516 (N_14516,N_13687,N_13861);
nand U14517 (N_14517,N_12970,N_13502);
and U14518 (N_14518,N_13348,N_12734);
or U14519 (N_14519,N_12612,N_12368);
nor U14520 (N_14520,N_13482,N_12253);
nand U14521 (N_14521,N_12361,N_13663);
nor U14522 (N_14522,N_13024,N_12288);
and U14523 (N_14523,N_13688,N_13735);
or U14524 (N_14524,N_12318,N_12317);
nor U14525 (N_14525,N_13897,N_12591);
nand U14526 (N_14526,N_12254,N_12511);
xor U14527 (N_14527,N_12175,N_12199);
nand U14528 (N_14528,N_12409,N_13176);
and U14529 (N_14529,N_12574,N_12195);
nor U14530 (N_14530,N_12604,N_12510);
nand U14531 (N_14531,N_13533,N_12780);
xor U14532 (N_14532,N_13666,N_12767);
and U14533 (N_14533,N_12080,N_12616);
xor U14534 (N_14534,N_12197,N_13534);
or U14535 (N_14535,N_12206,N_12037);
nor U14536 (N_14536,N_13147,N_13574);
xor U14537 (N_14537,N_13650,N_13448);
xnor U14538 (N_14538,N_13946,N_13783);
nand U14539 (N_14539,N_12159,N_13385);
nand U14540 (N_14540,N_13407,N_12855);
and U14541 (N_14541,N_12494,N_12969);
and U14542 (N_14542,N_13262,N_13635);
nand U14543 (N_14543,N_13484,N_13031);
xnor U14544 (N_14544,N_12211,N_12738);
nand U14545 (N_14545,N_12558,N_13394);
nand U14546 (N_14546,N_13570,N_12166);
or U14547 (N_14547,N_12491,N_12323);
xnor U14548 (N_14548,N_12860,N_12810);
nand U14549 (N_14549,N_12946,N_12539);
nand U14550 (N_14550,N_12389,N_13249);
or U14551 (N_14551,N_13957,N_13454);
nand U14552 (N_14552,N_13776,N_12226);
nand U14553 (N_14553,N_12000,N_13066);
nor U14554 (N_14554,N_13690,N_12977);
or U14555 (N_14555,N_13812,N_12715);
xnor U14556 (N_14556,N_12721,N_12290);
xnor U14557 (N_14557,N_13426,N_13020);
or U14558 (N_14558,N_12300,N_12896);
xnor U14559 (N_14559,N_13278,N_12951);
nand U14560 (N_14560,N_12148,N_13246);
and U14561 (N_14561,N_12310,N_12699);
or U14562 (N_14562,N_12065,N_12133);
xnor U14563 (N_14563,N_13608,N_12157);
and U14564 (N_14564,N_13240,N_12768);
nor U14565 (N_14565,N_12181,N_12233);
or U14566 (N_14566,N_12024,N_12198);
nor U14567 (N_14567,N_12626,N_13719);
nand U14568 (N_14568,N_12636,N_13779);
nand U14569 (N_14569,N_12850,N_12059);
and U14570 (N_14570,N_13107,N_13799);
or U14571 (N_14571,N_13507,N_13478);
and U14572 (N_14572,N_12827,N_13381);
nor U14573 (N_14573,N_13291,N_12546);
or U14574 (N_14574,N_13195,N_13062);
nand U14575 (N_14575,N_13936,N_13156);
nor U14576 (N_14576,N_12051,N_13161);
nor U14577 (N_14577,N_13948,N_13591);
nor U14578 (N_14578,N_13661,N_13624);
and U14579 (N_14579,N_13527,N_13924);
or U14580 (N_14580,N_12755,N_12324);
or U14581 (N_14581,N_12595,N_12151);
or U14582 (N_14582,N_12274,N_12375);
and U14583 (N_14583,N_13491,N_12470);
or U14584 (N_14584,N_12216,N_13226);
xor U14585 (N_14585,N_13211,N_12006);
nor U14586 (N_14586,N_12988,N_13778);
nor U14587 (N_14587,N_13433,N_13770);
xor U14588 (N_14588,N_12825,N_13649);
or U14589 (N_14589,N_13388,N_13860);
or U14590 (N_14590,N_13513,N_13971);
nor U14591 (N_14591,N_13926,N_12783);
nor U14592 (N_14592,N_12653,N_12426);
and U14593 (N_14593,N_12264,N_12193);
nor U14594 (N_14594,N_13518,N_13346);
nand U14595 (N_14595,N_13365,N_13698);
and U14596 (N_14596,N_13369,N_13858);
and U14597 (N_14597,N_12120,N_12299);
nor U14598 (N_14598,N_13999,N_13762);
or U14599 (N_14599,N_12071,N_12915);
nand U14600 (N_14600,N_13149,N_13445);
or U14601 (N_14601,N_12941,N_12261);
or U14602 (N_14602,N_12189,N_12841);
and U14603 (N_14603,N_12545,N_13129);
or U14604 (N_14604,N_12683,N_12677);
and U14605 (N_14605,N_13313,N_12876);
nand U14606 (N_14606,N_13185,N_12022);
nand U14607 (N_14607,N_13061,N_12063);
xnor U14608 (N_14608,N_12580,N_13378);
xnor U14609 (N_14609,N_12281,N_12429);
or U14610 (N_14610,N_13931,N_13023);
nand U14611 (N_14611,N_12031,N_13002);
xnor U14612 (N_14612,N_12949,N_12778);
nor U14613 (N_14613,N_12441,N_12493);
nor U14614 (N_14614,N_13510,N_12320);
nand U14615 (N_14615,N_12808,N_13886);
and U14616 (N_14616,N_13594,N_12238);
or U14617 (N_14617,N_12150,N_12670);
xor U14618 (N_14618,N_12158,N_12830);
and U14619 (N_14619,N_13120,N_13734);
nand U14620 (N_14620,N_12530,N_12010);
nand U14621 (N_14621,N_13276,N_13465);
nand U14622 (N_14622,N_13749,N_12563);
nand U14623 (N_14623,N_13707,N_12531);
nand U14624 (N_14624,N_12049,N_12307);
nand U14625 (N_14625,N_13664,N_13997);
nor U14626 (N_14626,N_12294,N_12308);
and U14627 (N_14627,N_13464,N_13257);
xnor U14628 (N_14628,N_12924,N_12534);
or U14629 (N_14629,N_12265,N_12270);
and U14630 (N_14630,N_13657,N_13006);
and U14631 (N_14631,N_12961,N_13912);
nand U14632 (N_14632,N_12751,N_13044);
and U14633 (N_14633,N_12142,N_12445);
nand U14634 (N_14634,N_13602,N_12077);
xnor U14635 (N_14635,N_12963,N_13116);
xnor U14636 (N_14636,N_13760,N_13794);
and U14637 (N_14637,N_13951,N_13634);
xor U14638 (N_14638,N_12279,N_13301);
nor U14639 (N_14639,N_13468,N_13625);
and U14640 (N_14640,N_12883,N_12673);
nand U14641 (N_14641,N_12807,N_13703);
nand U14642 (N_14642,N_13152,N_12094);
and U14643 (N_14643,N_12283,N_12945);
and U14644 (N_14644,N_12753,N_12948);
or U14645 (N_14645,N_13743,N_13940);
and U14646 (N_14646,N_13110,N_13112);
or U14647 (N_14647,N_12117,N_13343);
xnor U14648 (N_14648,N_13756,N_13204);
nand U14649 (N_14649,N_13283,N_13012);
or U14650 (N_14650,N_13901,N_13505);
nor U14651 (N_14651,N_12718,N_13051);
nand U14652 (N_14652,N_12225,N_13868);
and U14653 (N_14653,N_13056,N_13026);
xor U14654 (N_14654,N_12332,N_13754);
nand U14655 (N_14655,N_12337,N_12034);
nor U14656 (N_14656,N_12906,N_12399);
nand U14657 (N_14657,N_12747,N_13064);
nor U14658 (N_14658,N_12606,N_12021);
xnor U14659 (N_14659,N_12497,N_12029);
or U14660 (N_14660,N_13011,N_12425);
nand U14661 (N_14661,N_12496,N_12388);
nor U14662 (N_14662,N_13207,N_12488);
xor U14663 (N_14663,N_12879,N_13260);
and U14664 (N_14664,N_12345,N_13341);
nand U14665 (N_14665,N_12369,N_13192);
nand U14666 (N_14666,N_12232,N_13848);
and U14667 (N_14667,N_12333,N_13600);
or U14668 (N_14668,N_12464,N_13362);
nand U14669 (N_14669,N_13648,N_13919);
xor U14670 (N_14670,N_13636,N_12376);
nor U14671 (N_14671,N_12544,N_13984);
nor U14672 (N_14672,N_12984,N_13759);
xnor U14673 (N_14673,N_12339,N_13689);
xnor U14674 (N_14674,N_12821,N_13589);
nand U14675 (N_14675,N_13656,N_12381);
nand U14676 (N_14676,N_12822,N_12314);
nand U14677 (N_14677,N_12386,N_13561);
xnor U14678 (N_14678,N_13470,N_13718);
and U14679 (N_14679,N_13974,N_12664);
nand U14680 (N_14680,N_13008,N_12886);
nor U14681 (N_14681,N_12862,N_13839);
and U14682 (N_14682,N_13225,N_13937);
and U14683 (N_14683,N_12116,N_13952);
and U14684 (N_14684,N_12956,N_13355);
and U14685 (N_14685,N_12127,N_13885);
and U14686 (N_14686,N_12844,N_12219);
and U14687 (N_14687,N_12881,N_13155);
xor U14688 (N_14688,N_13160,N_13639);
nor U14689 (N_14689,N_13055,N_13671);
and U14690 (N_14690,N_13838,N_12292);
or U14691 (N_14691,N_13787,N_12918);
nor U14692 (N_14692,N_12611,N_13227);
nor U14693 (N_14693,N_13644,N_12864);
or U14694 (N_14694,N_13894,N_12418);
nand U14695 (N_14695,N_13022,N_13945);
and U14696 (N_14696,N_12667,N_13615);
or U14697 (N_14697,N_13856,N_12170);
and U14698 (N_14698,N_12610,N_13449);
xor U14699 (N_14699,N_13563,N_12039);
nand U14700 (N_14700,N_13619,N_12374);
and U14701 (N_14701,N_13130,N_12703);
nor U14702 (N_14702,N_12266,N_13406);
xor U14703 (N_14703,N_12589,N_12739);
or U14704 (N_14704,N_12355,N_13032);
xnor U14705 (N_14705,N_12173,N_13494);
and U14706 (N_14706,N_12532,N_13837);
nand U14707 (N_14707,N_12220,N_13668);
nand U14708 (N_14708,N_13750,N_13098);
xnor U14709 (N_14709,N_13774,N_13546);
nor U14710 (N_14710,N_13010,N_12003);
xnor U14711 (N_14711,N_13189,N_12685);
nor U14712 (N_14712,N_12130,N_12403);
nand U14713 (N_14713,N_13569,N_12578);
or U14714 (N_14714,N_12342,N_12295);
nand U14715 (N_14715,N_13996,N_12002);
or U14716 (N_14716,N_13640,N_13741);
or U14717 (N_14717,N_12335,N_13675);
and U14718 (N_14718,N_13467,N_13001);
nor U14719 (N_14719,N_12452,N_12786);
and U14720 (N_14720,N_13132,N_12480);
xnor U14721 (N_14721,N_13562,N_12986);
or U14722 (N_14722,N_13057,N_13279);
nand U14723 (N_14723,N_13785,N_13434);
nor U14724 (N_14724,N_12824,N_13878);
nor U14725 (N_14725,N_13492,N_12023);
nor U14726 (N_14726,N_13704,N_12592);
nand U14727 (N_14727,N_12998,N_13288);
or U14728 (N_14728,N_13875,N_13180);
and U14729 (N_14729,N_12343,N_12458);
nor U14730 (N_14730,N_12468,N_13292);
nand U14731 (N_14731,N_12965,N_12241);
or U14732 (N_14732,N_12235,N_13319);
xor U14733 (N_14733,N_13637,N_12152);
nor U14734 (N_14734,N_13270,N_12690);
and U14735 (N_14735,N_12888,N_13067);
or U14736 (N_14736,N_12733,N_13862);
nor U14737 (N_14737,N_12124,N_12240);
or U14738 (N_14738,N_12191,N_13806);
nand U14739 (N_14739,N_12903,N_13424);
or U14740 (N_14740,N_12646,N_12866);
nand U14741 (N_14741,N_13052,N_12868);
nor U14742 (N_14742,N_12890,N_12921);
or U14743 (N_14743,N_12625,N_12579);
nand U14744 (N_14744,N_13966,N_13018);
or U14745 (N_14745,N_13777,N_13311);
xor U14746 (N_14746,N_12593,N_12041);
or U14747 (N_14747,N_13695,N_13628);
nand U14748 (N_14748,N_12509,N_12296);
nand U14749 (N_14749,N_13359,N_13162);
or U14750 (N_14750,N_13079,N_13197);
or U14751 (N_14751,N_12696,N_12898);
xor U14752 (N_14752,N_12372,N_13322);
xor U14753 (N_14753,N_12104,N_12939);
nand U14754 (N_14754,N_12088,N_13923);
and U14755 (N_14755,N_13103,N_13781);
or U14756 (N_14756,N_13673,N_13684);
nand U14757 (N_14757,N_12859,N_13891);
nand U14758 (N_14758,N_13247,N_12007);
xor U14759 (N_14759,N_12102,N_13159);
xor U14760 (N_14760,N_12894,N_12008);
xor U14761 (N_14761,N_13320,N_13512);
xor U14762 (N_14762,N_12659,N_12214);
nor U14763 (N_14763,N_13581,N_12829);
or U14764 (N_14764,N_12378,N_12582);
and U14765 (N_14765,N_13526,N_13493);
and U14766 (N_14766,N_12058,N_12620);
and U14767 (N_14767,N_12603,N_12340);
nand U14768 (N_14768,N_12081,N_12227);
xor U14769 (N_14769,N_13566,N_13733);
nor U14770 (N_14770,N_13021,N_13186);
nand U14771 (N_14771,N_13122,N_13631);
xnor U14772 (N_14772,N_12014,N_12125);
or U14773 (N_14773,N_12895,N_13135);
or U14774 (N_14774,N_12702,N_12508);
nand U14775 (N_14775,N_12665,N_13825);
nand U14776 (N_14776,N_12451,N_12581);
xnor U14777 (N_14777,N_13786,N_12258);
xor U14778 (N_14778,N_12326,N_12568);
nand U14779 (N_14779,N_12566,N_12103);
and U14780 (N_14780,N_12647,N_13645);
nor U14781 (N_14781,N_12785,N_13638);
nand U14782 (N_14782,N_13352,N_13691);
nand U14783 (N_14783,N_12800,N_13224);
xnor U14784 (N_14784,N_13418,N_13819);
nor U14785 (N_14785,N_12845,N_12650);
xor U14786 (N_14786,N_12700,N_13845);
nor U14787 (N_14787,N_12724,N_13895);
nand U14788 (N_14788,N_12529,N_13970);
or U14789 (N_14789,N_12230,N_13223);
and U14790 (N_14790,N_12843,N_12774);
nor U14791 (N_14791,N_12641,N_13212);
nor U14792 (N_14792,N_12050,N_12812);
nor U14793 (N_14793,N_13855,N_12495);
and U14794 (N_14794,N_13681,N_13903);
xor U14795 (N_14795,N_12761,N_13761);
nand U14796 (N_14796,N_12869,N_12705);
or U14797 (N_14797,N_13015,N_13463);
or U14798 (N_14798,N_13930,N_12542);
or U14799 (N_14799,N_13293,N_13556);
xnor U14800 (N_14800,N_12674,N_12053);
and U14801 (N_14801,N_12588,N_12955);
xor U14802 (N_14802,N_13995,N_12479);
and U14803 (N_14803,N_13763,N_13567);
and U14804 (N_14804,N_12210,N_13672);
and U14805 (N_14805,N_13323,N_12872);
xor U14806 (N_14806,N_12736,N_12485);
and U14807 (N_14807,N_13382,N_13316);
or U14808 (N_14808,N_12096,N_12373);
nand U14809 (N_14809,N_13865,N_13088);
xor U14810 (N_14810,N_12363,N_12745);
nand U14811 (N_14811,N_12139,N_13740);
nor U14812 (N_14812,N_13136,N_12435);
xnor U14813 (N_14813,N_13714,N_12764);
nor U14814 (N_14814,N_13095,N_12145);
nor U14815 (N_14815,N_13746,N_12536);
and U14816 (N_14816,N_13383,N_12576);
or U14817 (N_14817,N_12675,N_13459);
nand U14818 (N_14818,N_13791,N_13347);
xnor U14819 (N_14819,N_13340,N_13588);
and U14820 (N_14820,N_12516,N_13990);
nor U14821 (N_14821,N_13241,N_12136);
nor U14822 (N_14822,N_12506,N_12262);
and U14823 (N_14823,N_13893,N_12160);
nor U14824 (N_14824,N_13065,N_12208);
or U14825 (N_14825,N_13536,N_12179);
and U14826 (N_14826,N_13398,N_12629);
xnor U14827 (N_14827,N_13606,N_12083);
and U14828 (N_14828,N_13523,N_12560);
nor U14829 (N_14829,N_13237,N_12704);
nand U14830 (N_14830,N_13072,N_12285);
xnor U14831 (N_14831,N_12698,N_12541);
and U14832 (N_14832,N_12301,N_13592);
and U14833 (N_14833,N_13872,N_12463);
xor U14834 (N_14834,N_12304,N_13254);
nand U14835 (N_14835,N_12982,N_12676);
and U14836 (N_14836,N_13841,N_12569);
nor U14837 (N_14837,N_13890,N_13480);
xor U14838 (N_14838,N_12958,N_12849);
nor U14839 (N_14839,N_13622,N_12515);
and U14840 (N_14840,N_13532,N_13373);
xor U14841 (N_14841,N_13408,N_13121);
nand U14842 (N_14842,N_12652,N_13679);
xnor U14843 (N_14843,N_12929,N_13810);
nor U14844 (N_14844,N_12899,N_12605);
nor U14845 (N_14845,N_12567,N_12635);
nor U14846 (N_14846,N_12257,N_13308);
and U14847 (N_14847,N_12692,N_12017);
nor U14848 (N_14848,N_12236,N_12395);
nand U14849 (N_14849,N_12549,N_12893);
or U14850 (N_14850,N_13145,N_13336);
or U14851 (N_14851,N_13818,N_12639);
nand U14852 (N_14852,N_13918,N_12196);
and U14853 (N_14853,N_13932,N_12313);
nand U14854 (N_14854,N_12256,N_12525);
or U14855 (N_14855,N_12777,N_12995);
nor U14856 (N_14856,N_13568,N_12932);
nand U14857 (N_14857,N_13274,N_13545);
nand U14858 (N_14858,N_13697,N_13604);
nand U14859 (N_14859,N_12459,N_12052);
or U14860 (N_14860,N_12910,N_13745);
nor U14861 (N_14861,N_13045,N_12976);
nor U14862 (N_14862,N_13306,N_12914);
or U14863 (N_14863,N_13961,N_13139);
nand U14864 (N_14864,N_12882,N_13253);
and U14865 (N_14865,N_12503,N_12640);
nor U14866 (N_14866,N_12359,N_12902);
xnor U14867 (N_14867,N_13096,N_13623);
nor U14868 (N_14868,N_13721,N_13094);
nand U14869 (N_14869,N_13473,N_12913);
nor U14870 (N_14870,N_12513,N_12695);
or U14871 (N_14871,N_12245,N_13451);
xnor U14872 (N_14872,N_12871,N_13273);
and U14873 (N_14873,N_13947,N_13827);
nand U14874 (N_14874,N_13138,N_13331);
xor U14875 (N_14875,N_12551,N_13019);
xor U14876 (N_14876,N_12269,N_12417);
nand U14877 (N_14877,N_12055,N_12624);
xor U14878 (N_14878,N_13416,N_13483);
and U14879 (N_14879,N_12126,N_12759);
or U14880 (N_14880,N_13933,N_13339);
and U14881 (N_14881,N_12192,N_13655);
nor U14882 (N_14882,N_13153,N_13456);
nand U14883 (N_14883,N_13755,N_13025);
nand U14884 (N_14884,N_12682,N_13487);
and U14885 (N_14885,N_12538,N_12658);
nand U14886 (N_14886,N_13551,N_13109);
or U14887 (N_14887,N_13960,N_12271);
and U14888 (N_14888,N_12427,N_13902);
nor U14889 (N_14889,N_13809,N_12930);
nand U14890 (N_14890,N_13317,N_13846);
nor U14891 (N_14891,N_12547,N_12312);
nor U14892 (N_14892,N_12818,N_12701);
or U14893 (N_14893,N_12090,N_13238);
xor U14894 (N_14894,N_13297,N_13386);
xor U14895 (N_14895,N_13887,N_13353);
nand U14896 (N_14896,N_12645,N_13586);
and U14897 (N_14897,N_12973,N_12556);
xnor U14898 (N_14898,N_13350,N_13174);
nor U14899 (N_14899,N_12168,N_12364);
or U14900 (N_14900,N_13983,N_13884);
xor U14901 (N_14901,N_12467,N_12706);
and U14902 (N_14902,N_13443,N_12730);
xor U14903 (N_14903,N_13280,N_13915);
or U14904 (N_14904,N_12419,N_12387);
or U14905 (N_14905,N_12492,N_13367);
or U14906 (N_14906,N_12180,N_12805);
xor U14907 (N_14907,N_13236,N_12165);
nand U14908 (N_14908,N_13647,N_13368);
nor U14909 (N_14909,N_13992,N_12691);
xor U14910 (N_14910,N_13193,N_12424);
nand U14911 (N_14911,N_13730,N_12694);
or U14912 (N_14912,N_12297,N_13356);
and U14913 (N_14913,N_12726,N_13256);
xor U14914 (N_14914,N_12832,N_13242);
nand U14915 (N_14915,N_13184,N_12070);
or U14916 (N_14916,N_12026,N_13358);
nand U14917 (N_14917,N_13447,N_12681);
nor U14918 (N_14918,N_13082,N_12161);
nor U14919 (N_14919,N_12404,N_13967);
and U14920 (N_14920,N_12993,N_13686);
xor U14921 (N_14921,N_12436,N_13873);
nand U14922 (N_14922,N_12746,N_12711);
nand U14923 (N_14923,N_12613,N_12268);
nor U14924 (N_14924,N_13234,N_12129);
nor U14925 (N_14925,N_12816,N_13458);
or U14926 (N_14926,N_12020,N_13059);
xnor U14927 (N_14927,N_13286,N_13612);
xor U14928 (N_14928,N_13069,N_12689);
and U14929 (N_14929,N_13646,N_12555);
and U14930 (N_14930,N_12634,N_12723);
and U14931 (N_14931,N_13182,N_12194);
nor U14932 (N_14932,N_12617,N_13412);
and U14933 (N_14933,N_13660,N_13036);
and U14934 (N_14934,N_13014,N_13134);
or U14935 (N_14935,N_12143,N_12907);
nand U14936 (N_14936,N_13949,N_13596);
and U14937 (N_14937,N_13826,N_12449);
nand U14938 (N_14938,N_12772,N_12856);
or U14939 (N_14939,N_13284,N_12654);
nand U14940 (N_14940,N_13440,N_13844);
nor U14941 (N_14941,N_12113,N_13497);
and U14942 (N_14942,N_12992,N_13705);
nand U14943 (N_14943,N_13175,N_12035);
and U14944 (N_14944,N_13166,N_12430);
or U14945 (N_14945,N_13941,N_13277);
xor U14946 (N_14946,N_12840,N_13360);
nor U14947 (N_14947,N_13729,N_12912);
xnor U14948 (N_14948,N_13869,N_12030);
or U14949 (N_14949,N_12415,N_13883);
nand U14950 (N_14950,N_12394,N_12991);
or U14951 (N_14951,N_12937,N_13471);
xor U14952 (N_14952,N_13867,N_12144);
and U14953 (N_14953,N_13775,N_12972);
or U14954 (N_14954,N_13544,N_12347);
nand U14955 (N_14955,N_13030,N_13744);
nand U14956 (N_14956,N_13485,N_13111);
nand U14957 (N_14957,N_12396,N_12554);
and U14958 (N_14958,N_13678,N_12156);
or U14959 (N_14959,N_12111,N_13653);
nor U14960 (N_14960,N_12390,N_13938);
or U14961 (N_14961,N_12327,N_12405);
nor U14962 (N_14962,N_12412,N_13183);
and U14963 (N_14963,N_12484,N_12004);
nand U14964 (N_14964,N_13959,N_12276);
nand U14965 (N_14965,N_13815,N_12714);
or U14966 (N_14966,N_12248,N_13764);
or U14967 (N_14967,N_12520,N_12141);
xnor U14968 (N_14968,N_12500,N_12383);
or U14969 (N_14969,N_12571,N_12535);
or U14970 (N_14970,N_13213,N_12835);
and U14971 (N_14971,N_12086,N_13614);
nand U14972 (N_14972,N_13265,N_13677);
xnor U14973 (N_14973,N_12873,N_12223);
xor U14974 (N_14974,N_12942,N_12632);
xnor U14975 (N_14975,N_12115,N_13423);
nor U14976 (N_14976,N_12352,N_12979);
xnor U14977 (N_14977,N_12809,N_13928);
or U14978 (N_14978,N_13315,N_12981);
nor U14979 (N_14979,N_12974,N_13784);
and U14980 (N_14980,N_13296,N_13304);
nand U14981 (N_14981,N_13790,N_13917);
or U14982 (N_14982,N_12884,N_13870);
and U14983 (N_14983,N_12286,N_12765);
and U14984 (N_14984,N_13700,N_13230);
or U14985 (N_14985,N_13773,N_13281);
nand U14986 (N_14986,N_13450,N_12251);
nand U14987 (N_14987,N_12933,N_13198);
nor U14988 (N_14988,N_12797,N_12303);
and U14989 (N_14989,N_12794,N_13430);
and U14990 (N_14990,N_12572,N_12836);
nand U14991 (N_14991,N_13833,N_12162);
nor U14992 (N_14992,N_12769,N_13085);
nand U14993 (N_14993,N_12487,N_12651);
nand U14994 (N_14994,N_12575,N_13857);
and U14995 (N_14995,N_13053,N_12655);
xor U14996 (N_14996,N_13258,N_13547);
nor U14997 (N_14997,N_13100,N_12221);
xnor U14998 (N_14998,N_13091,N_12607);
xnor U14999 (N_14999,N_12456,N_12621);
nand U15000 (N_15000,N_12833,N_12734);
and U15001 (N_15001,N_13444,N_13040);
nand U15002 (N_15002,N_13491,N_13423);
nor U15003 (N_15003,N_12312,N_12640);
xor U15004 (N_15004,N_13421,N_12710);
xnor U15005 (N_15005,N_13391,N_12902);
nand U15006 (N_15006,N_13329,N_12290);
nand U15007 (N_15007,N_12592,N_12015);
xnor U15008 (N_15008,N_13642,N_12346);
or U15009 (N_15009,N_12284,N_12291);
nor U15010 (N_15010,N_12961,N_12013);
xor U15011 (N_15011,N_13698,N_13471);
nand U15012 (N_15012,N_12995,N_12081);
or U15013 (N_15013,N_13003,N_12369);
or U15014 (N_15014,N_13998,N_13056);
nor U15015 (N_15015,N_12956,N_13477);
and U15016 (N_15016,N_13589,N_12774);
and U15017 (N_15017,N_13808,N_12406);
xor U15018 (N_15018,N_13058,N_12473);
xor U15019 (N_15019,N_12390,N_12816);
xor U15020 (N_15020,N_12595,N_12439);
xor U15021 (N_15021,N_13267,N_12327);
nand U15022 (N_15022,N_13204,N_12646);
nor U15023 (N_15023,N_12879,N_12529);
xnor U15024 (N_15024,N_12778,N_13439);
or U15025 (N_15025,N_13614,N_12678);
nor U15026 (N_15026,N_13468,N_12521);
nor U15027 (N_15027,N_12828,N_13434);
xnor U15028 (N_15028,N_12054,N_12556);
nand U15029 (N_15029,N_13989,N_13229);
xnor U15030 (N_15030,N_13219,N_12366);
or U15031 (N_15031,N_13726,N_12754);
nor U15032 (N_15032,N_13849,N_13643);
xor U15033 (N_15033,N_13927,N_13800);
or U15034 (N_15034,N_12818,N_12744);
nor U15035 (N_15035,N_12725,N_13137);
nand U15036 (N_15036,N_12060,N_13609);
nor U15037 (N_15037,N_12997,N_13176);
and U15038 (N_15038,N_12135,N_12828);
xnor U15039 (N_15039,N_12663,N_12794);
and U15040 (N_15040,N_12796,N_13716);
nand U15041 (N_15041,N_13731,N_13204);
or U15042 (N_15042,N_12533,N_13737);
or U15043 (N_15043,N_12009,N_12892);
nor U15044 (N_15044,N_12031,N_12130);
xnor U15045 (N_15045,N_13257,N_12831);
nor U15046 (N_15046,N_12345,N_12004);
xor U15047 (N_15047,N_12632,N_12800);
or U15048 (N_15048,N_12439,N_13428);
and U15049 (N_15049,N_13698,N_13720);
nor U15050 (N_15050,N_12226,N_13778);
and U15051 (N_15051,N_13441,N_13472);
or U15052 (N_15052,N_12805,N_12278);
nor U15053 (N_15053,N_13019,N_12197);
nand U15054 (N_15054,N_13164,N_12182);
or U15055 (N_15055,N_13057,N_12695);
and U15056 (N_15056,N_12549,N_12154);
xor U15057 (N_15057,N_12636,N_12986);
nor U15058 (N_15058,N_13518,N_12414);
nor U15059 (N_15059,N_12399,N_13049);
nand U15060 (N_15060,N_13439,N_13493);
and U15061 (N_15061,N_13227,N_13205);
and U15062 (N_15062,N_12335,N_12726);
or U15063 (N_15063,N_12280,N_13939);
nand U15064 (N_15064,N_12760,N_12020);
or U15065 (N_15065,N_12260,N_12294);
or U15066 (N_15066,N_12412,N_12330);
nand U15067 (N_15067,N_13221,N_13857);
nor U15068 (N_15068,N_13204,N_13506);
nor U15069 (N_15069,N_13571,N_13254);
and U15070 (N_15070,N_13498,N_12169);
xor U15071 (N_15071,N_12680,N_12356);
and U15072 (N_15072,N_12793,N_12581);
nor U15073 (N_15073,N_13332,N_12616);
or U15074 (N_15074,N_12963,N_13411);
nor U15075 (N_15075,N_13121,N_12530);
and U15076 (N_15076,N_12537,N_13619);
or U15077 (N_15077,N_12576,N_13931);
nor U15078 (N_15078,N_12728,N_12794);
nor U15079 (N_15079,N_13580,N_12291);
or U15080 (N_15080,N_13108,N_13337);
xor U15081 (N_15081,N_12312,N_13181);
or U15082 (N_15082,N_12313,N_13918);
or U15083 (N_15083,N_13448,N_12367);
or U15084 (N_15084,N_12074,N_13195);
nand U15085 (N_15085,N_13611,N_12049);
xnor U15086 (N_15086,N_12856,N_12092);
nand U15087 (N_15087,N_12216,N_13451);
and U15088 (N_15088,N_13312,N_12458);
nand U15089 (N_15089,N_13817,N_12231);
nor U15090 (N_15090,N_13686,N_12885);
and U15091 (N_15091,N_13293,N_12855);
nand U15092 (N_15092,N_12466,N_12251);
nor U15093 (N_15093,N_12504,N_13174);
nand U15094 (N_15094,N_12484,N_12754);
and U15095 (N_15095,N_13484,N_13860);
nand U15096 (N_15096,N_13614,N_12397);
or U15097 (N_15097,N_12359,N_13543);
xor U15098 (N_15098,N_12261,N_12784);
xor U15099 (N_15099,N_12338,N_13781);
nand U15100 (N_15100,N_13157,N_12908);
nor U15101 (N_15101,N_13238,N_13075);
or U15102 (N_15102,N_13446,N_12683);
and U15103 (N_15103,N_13689,N_13910);
nor U15104 (N_15104,N_12272,N_12388);
nand U15105 (N_15105,N_13165,N_12218);
nor U15106 (N_15106,N_13896,N_13437);
nand U15107 (N_15107,N_13559,N_12923);
nor U15108 (N_15108,N_13057,N_12566);
nor U15109 (N_15109,N_12608,N_12144);
nand U15110 (N_15110,N_13914,N_12334);
and U15111 (N_15111,N_12256,N_13945);
and U15112 (N_15112,N_13134,N_13184);
or U15113 (N_15113,N_12681,N_12247);
xor U15114 (N_15114,N_13478,N_13163);
xnor U15115 (N_15115,N_13575,N_13827);
or U15116 (N_15116,N_13559,N_13170);
nor U15117 (N_15117,N_13768,N_12449);
and U15118 (N_15118,N_13751,N_12814);
xor U15119 (N_15119,N_12497,N_12106);
or U15120 (N_15120,N_13804,N_12971);
xnor U15121 (N_15121,N_13080,N_13245);
nor U15122 (N_15122,N_13650,N_12756);
nor U15123 (N_15123,N_13803,N_13757);
or U15124 (N_15124,N_12092,N_12774);
or U15125 (N_15125,N_13565,N_12945);
xor U15126 (N_15126,N_13960,N_13665);
or U15127 (N_15127,N_12021,N_12822);
xor U15128 (N_15128,N_13306,N_13530);
nor U15129 (N_15129,N_13583,N_12045);
xnor U15130 (N_15130,N_13787,N_12901);
xor U15131 (N_15131,N_13543,N_12926);
nor U15132 (N_15132,N_12996,N_12384);
nor U15133 (N_15133,N_13355,N_13098);
xor U15134 (N_15134,N_12961,N_13868);
or U15135 (N_15135,N_12615,N_12510);
xnor U15136 (N_15136,N_12528,N_13786);
or U15137 (N_15137,N_12510,N_13052);
nor U15138 (N_15138,N_12719,N_13678);
nor U15139 (N_15139,N_12801,N_13314);
nor U15140 (N_15140,N_13735,N_12332);
and U15141 (N_15141,N_12153,N_13611);
xnor U15142 (N_15142,N_13677,N_12769);
or U15143 (N_15143,N_13782,N_13423);
xor U15144 (N_15144,N_12792,N_13057);
or U15145 (N_15145,N_13185,N_13681);
and U15146 (N_15146,N_13724,N_13924);
or U15147 (N_15147,N_12655,N_12204);
nor U15148 (N_15148,N_13181,N_12315);
and U15149 (N_15149,N_13448,N_12203);
nor U15150 (N_15150,N_12040,N_13612);
and U15151 (N_15151,N_12033,N_13839);
nand U15152 (N_15152,N_13547,N_12672);
nor U15153 (N_15153,N_12094,N_13616);
or U15154 (N_15154,N_13623,N_12113);
xor U15155 (N_15155,N_13221,N_13951);
and U15156 (N_15156,N_13429,N_12983);
or U15157 (N_15157,N_13659,N_12852);
or U15158 (N_15158,N_13179,N_12603);
or U15159 (N_15159,N_13924,N_13461);
and U15160 (N_15160,N_12065,N_12992);
nor U15161 (N_15161,N_13352,N_12651);
nand U15162 (N_15162,N_12199,N_13910);
nor U15163 (N_15163,N_13928,N_12606);
or U15164 (N_15164,N_12547,N_12420);
xor U15165 (N_15165,N_12386,N_13493);
or U15166 (N_15166,N_12670,N_12464);
nor U15167 (N_15167,N_13085,N_12628);
nand U15168 (N_15168,N_13322,N_13095);
and U15169 (N_15169,N_12651,N_13882);
nand U15170 (N_15170,N_12679,N_13187);
xnor U15171 (N_15171,N_12322,N_12460);
xnor U15172 (N_15172,N_12187,N_12782);
or U15173 (N_15173,N_13818,N_12960);
or U15174 (N_15174,N_12282,N_13175);
nand U15175 (N_15175,N_12063,N_13318);
nand U15176 (N_15176,N_12729,N_13298);
nor U15177 (N_15177,N_13265,N_12054);
and U15178 (N_15178,N_13802,N_13992);
xor U15179 (N_15179,N_13915,N_12435);
nor U15180 (N_15180,N_12966,N_12060);
nor U15181 (N_15181,N_12017,N_12757);
nor U15182 (N_15182,N_13721,N_12479);
xor U15183 (N_15183,N_12516,N_12049);
nor U15184 (N_15184,N_13892,N_12514);
nand U15185 (N_15185,N_13781,N_12566);
or U15186 (N_15186,N_13943,N_13588);
and U15187 (N_15187,N_13037,N_13775);
xnor U15188 (N_15188,N_13333,N_13328);
nor U15189 (N_15189,N_12812,N_13703);
or U15190 (N_15190,N_12598,N_12606);
and U15191 (N_15191,N_12944,N_13992);
nor U15192 (N_15192,N_13650,N_12058);
and U15193 (N_15193,N_13086,N_13972);
nand U15194 (N_15194,N_12672,N_12071);
and U15195 (N_15195,N_13338,N_12511);
nand U15196 (N_15196,N_12650,N_13622);
xnor U15197 (N_15197,N_13281,N_12141);
nor U15198 (N_15198,N_12156,N_13601);
and U15199 (N_15199,N_12866,N_13538);
and U15200 (N_15200,N_12565,N_12072);
nor U15201 (N_15201,N_13465,N_13370);
xnor U15202 (N_15202,N_12215,N_13662);
nor U15203 (N_15203,N_13475,N_13084);
and U15204 (N_15204,N_13734,N_13067);
nand U15205 (N_15205,N_12734,N_13535);
or U15206 (N_15206,N_12538,N_12777);
or U15207 (N_15207,N_12103,N_13055);
nand U15208 (N_15208,N_13062,N_13434);
or U15209 (N_15209,N_12134,N_13558);
xnor U15210 (N_15210,N_13897,N_12723);
nand U15211 (N_15211,N_13110,N_12957);
xor U15212 (N_15212,N_12747,N_12565);
and U15213 (N_15213,N_13963,N_13057);
nand U15214 (N_15214,N_13030,N_13906);
or U15215 (N_15215,N_12391,N_12291);
or U15216 (N_15216,N_13115,N_13676);
or U15217 (N_15217,N_12831,N_13148);
and U15218 (N_15218,N_13997,N_12779);
nor U15219 (N_15219,N_12683,N_12133);
nor U15220 (N_15220,N_13955,N_13953);
and U15221 (N_15221,N_13009,N_12541);
or U15222 (N_15222,N_12372,N_13130);
nor U15223 (N_15223,N_13474,N_12301);
nand U15224 (N_15224,N_12946,N_12838);
nand U15225 (N_15225,N_13027,N_13070);
nand U15226 (N_15226,N_13315,N_13254);
or U15227 (N_15227,N_13648,N_12336);
xor U15228 (N_15228,N_13728,N_12980);
or U15229 (N_15229,N_13142,N_12085);
xor U15230 (N_15230,N_13648,N_13266);
and U15231 (N_15231,N_13747,N_12208);
or U15232 (N_15232,N_12019,N_12466);
xnor U15233 (N_15233,N_13000,N_13707);
or U15234 (N_15234,N_12964,N_13066);
or U15235 (N_15235,N_13313,N_13047);
nor U15236 (N_15236,N_13122,N_12894);
nand U15237 (N_15237,N_13931,N_13378);
nand U15238 (N_15238,N_13605,N_13864);
and U15239 (N_15239,N_12582,N_13028);
and U15240 (N_15240,N_13606,N_13790);
or U15241 (N_15241,N_12806,N_13104);
or U15242 (N_15242,N_12245,N_13652);
nand U15243 (N_15243,N_12375,N_12857);
and U15244 (N_15244,N_13717,N_13017);
nor U15245 (N_15245,N_12247,N_12094);
nand U15246 (N_15246,N_12044,N_12663);
and U15247 (N_15247,N_12618,N_13129);
xnor U15248 (N_15248,N_13808,N_12975);
or U15249 (N_15249,N_13899,N_12958);
nor U15250 (N_15250,N_13128,N_13033);
or U15251 (N_15251,N_12121,N_12425);
and U15252 (N_15252,N_13487,N_12950);
nor U15253 (N_15253,N_13105,N_13623);
or U15254 (N_15254,N_13649,N_13716);
or U15255 (N_15255,N_13303,N_13414);
nor U15256 (N_15256,N_12206,N_13536);
or U15257 (N_15257,N_13484,N_13041);
nand U15258 (N_15258,N_12157,N_13980);
or U15259 (N_15259,N_12980,N_12520);
and U15260 (N_15260,N_13877,N_12401);
nor U15261 (N_15261,N_12337,N_12371);
nor U15262 (N_15262,N_13037,N_12958);
or U15263 (N_15263,N_13561,N_13712);
and U15264 (N_15264,N_12985,N_12719);
xor U15265 (N_15265,N_13162,N_12575);
nor U15266 (N_15266,N_12346,N_13522);
nor U15267 (N_15267,N_13710,N_12223);
nor U15268 (N_15268,N_12049,N_12930);
nand U15269 (N_15269,N_13504,N_13129);
or U15270 (N_15270,N_12413,N_13692);
or U15271 (N_15271,N_12851,N_12896);
xor U15272 (N_15272,N_12138,N_12567);
nor U15273 (N_15273,N_12566,N_13283);
xnor U15274 (N_15274,N_13528,N_12303);
nand U15275 (N_15275,N_12974,N_12567);
nor U15276 (N_15276,N_12230,N_13228);
and U15277 (N_15277,N_13872,N_13783);
nor U15278 (N_15278,N_13829,N_13527);
xor U15279 (N_15279,N_12380,N_12605);
and U15280 (N_15280,N_13045,N_12755);
nand U15281 (N_15281,N_13462,N_12202);
nor U15282 (N_15282,N_12235,N_12606);
nor U15283 (N_15283,N_13622,N_12192);
and U15284 (N_15284,N_13123,N_12347);
or U15285 (N_15285,N_12182,N_13001);
nand U15286 (N_15286,N_13166,N_12812);
nand U15287 (N_15287,N_13051,N_13467);
and U15288 (N_15288,N_12916,N_12201);
nand U15289 (N_15289,N_12466,N_13364);
xnor U15290 (N_15290,N_12308,N_12745);
xnor U15291 (N_15291,N_13670,N_12764);
and U15292 (N_15292,N_13207,N_12281);
xnor U15293 (N_15293,N_12002,N_13409);
or U15294 (N_15294,N_12320,N_13842);
and U15295 (N_15295,N_13485,N_13172);
and U15296 (N_15296,N_13827,N_12225);
nand U15297 (N_15297,N_12951,N_13830);
nor U15298 (N_15298,N_12366,N_12285);
or U15299 (N_15299,N_12806,N_13863);
nor U15300 (N_15300,N_13518,N_13797);
or U15301 (N_15301,N_13825,N_12794);
xor U15302 (N_15302,N_12497,N_12223);
nor U15303 (N_15303,N_13926,N_12348);
nor U15304 (N_15304,N_12779,N_13292);
or U15305 (N_15305,N_12534,N_12507);
nor U15306 (N_15306,N_13013,N_12766);
nor U15307 (N_15307,N_12678,N_12724);
nand U15308 (N_15308,N_13560,N_13818);
xnor U15309 (N_15309,N_12738,N_13792);
nand U15310 (N_15310,N_13163,N_13944);
nor U15311 (N_15311,N_12288,N_12549);
xor U15312 (N_15312,N_13022,N_12611);
or U15313 (N_15313,N_13309,N_12264);
or U15314 (N_15314,N_13121,N_12468);
xnor U15315 (N_15315,N_13386,N_13016);
nand U15316 (N_15316,N_13639,N_13468);
nand U15317 (N_15317,N_12794,N_12761);
nand U15318 (N_15318,N_12017,N_13631);
nor U15319 (N_15319,N_12206,N_13935);
and U15320 (N_15320,N_13758,N_13589);
nand U15321 (N_15321,N_13616,N_12575);
nand U15322 (N_15322,N_12567,N_12277);
nor U15323 (N_15323,N_13520,N_13507);
or U15324 (N_15324,N_13771,N_12721);
nand U15325 (N_15325,N_13178,N_13082);
or U15326 (N_15326,N_13284,N_12880);
nand U15327 (N_15327,N_12451,N_13373);
and U15328 (N_15328,N_12484,N_13296);
or U15329 (N_15329,N_13415,N_12977);
nand U15330 (N_15330,N_12282,N_12870);
xnor U15331 (N_15331,N_13768,N_13787);
nand U15332 (N_15332,N_13808,N_12215);
and U15333 (N_15333,N_12030,N_13831);
nand U15334 (N_15334,N_13708,N_13840);
or U15335 (N_15335,N_12319,N_13364);
or U15336 (N_15336,N_13547,N_13494);
and U15337 (N_15337,N_12815,N_13456);
nand U15338 (N_15338,N_12900,N_12237);
nor U15339 (N_15339,N_12887,N_12360);
xnor U15340 (N_15340,N_13583,N_13225);
or U15341 (N_15341,N_12633,N_12882);
and U15342 (N_15342,N_12785,N_12300);
xor U15343 (N_15343,N_13560,N_12233);
nor U15344 (N_15344,N_12889,N_12990);
nor U15345 (N_15345,N_12004,N_12793);
and U15346 (N_15346,N_13188,N_13633);
nor U15347 (N_15347,N_12979,N_12534);
or U15348 (N_15348,N_13885,N_13491);
xnor U15349 (N_15349,N_12299,N_13266);
nand U15350 (N_15350,N_13509,N_12448);
xor U15351 (N_15351,N_12163,N_12501);
and U15352 (N_15352,N_13758,N_13150);
and U15353 (N_15353,N_13321,N_12800);
or U15354 (N_15354,N_12330,N_12080);
and U15355 (N_15355,N_13450,N_13770);
or U15356 (N_15356,N_13260,N_12193);
xor U15357 (N_15357,N_12351,N_12890);
nor U15358 (N_15358,N_12442,N_12682);
and U15359 (N_15359,N_12947,N_13814);
and U15360 (N_15360,N_12233,N_13946);
nor U15361 (N_15361,N_13043,N_13846);
or U15362 (N_15362,N_12017,N_12651);
nand U15363 (N_15363,N_12224,N_13909);
or U15364 (N_15364,N_12135,N_13807);
and U15365 (N_15365,N_13463,N_13972);
nand U15366 (N_15366,N_12999,N_13501);
nor U15367 (N_15367,N_13422,N_13078);
or U15368 (N_15368,N_13461,N_12804);
or U15369 (N_15369,N_13801,N_12046);
nand U15370 (N_15370,N_12978,N_13057);
xnor U15371 (N_15371,N_12034,N_12360);
and U15372 (N_15372,N_12458,N_12000);
or U15373 (N_15373,N_13336,N_12423);
or U15374 (N_15374,N_12143,N_12359);
or U15375 (N_15375,N_13032,N_13073);
and U15376 (N_15376,N_13657,N_13071);
xnor U15377 (N_15377,N_12098,N_13973);
and U15378 (N_15378,N_12433,N_12111);
and U15379 (N_15379,N_13884,N_12539);
or U15380 (N_15380,N_12888,N_12325);
nor U15381 (N_15381,N_12468,N_12815);
nor U15382 (N_15382,N_12889,N_12712);
and U15383 (N_15383,N_12522,N_12231);
and U15384 (N_15384,N_12553,N_12304);
nor U15385 (N_15385,N_13306,N_13023);
or U15386 (N_15386,N_12636,N_13227);
nor U15387 (N_15387,N_13757,N_12272);
or U15388 (N_15388,N_12649,N_13037);
xor U15389 (N_15389,N_13261,N_12648);
nor U15390 (N_15390,N_12126,N_12940);
nor U15391 (N_15391,N_12890,N_13438);
and U15392 (N_15392,N_12273,N_13841);
xnor U15393 (N_15393,N_13102,N_13404);
nand U15394 (N_15394,N_13579,N_12127);
and U15395 (N_15395,N_13755,N_12824);
xor U15396 (N_15396,N_13722,N_13171);
xnor U15397 (N_15397,N_13399,N_12309);
and U15398 (N_15398,N_12464,N_13251);
and U15399 (N_15399,N_12472,N_12078);
and U15400 (N_15400,N_12631,N_12219);
nor U15401 (N_15401,N_12342,N_13831);
and U15402 (N_15402,N_12850,N_12079);
or U15403 (N_15403,N_12952,N_12926);
or U15404 (N_15404,N_13725,N_12295);
and U15405 (N_15405,N_12157,N_12071);
or U15406 (N_15406,N_13498,N_12429);
xor U15407 (N_15407,N_12958,N_12597);
or U15408 (N_15408,N_12636,N_12424);
or U15409 (N_15409,N_13289,N_12188);
nand U15410 (N_15410,N_13812,N_13715);
nand U15411 (N_15411,N_13885,N_12874);
xor U15412 (N_15412,N_12395,N_13818);
nor U15413 (N_15413,N_13337,N_12538);
xor U15414 (N_15414,N_13052,N_13919);
nand U15415 (N_15415,N_12002,N_12651);
nand U15416 (N_15416,N_13479,N_12736);
and U15417 (N_15417,N_12181,N_13609);
nor U15418 (N_15418,N_12635,N_12063);
or U15419 (N_15419,N_12426,N_12222);
or U15420 (N_15420,N_13657,N_13301);
nand U15421 (N_15421,N_12768,N_12602);
and U15422 (N_15422,N_12520,N_13190);
nor U15423 (N_15423,N_12236,N_12747);
xnor U15424 (N_15424,N_13016,N_12764);
and U15425 (N_15425,N_13215,N_12313);
xor U15426 (N_15426,N_13477,N_13619);
xor U15427 (N_15427,N_12074,N_13691);
and U15428 (N_15428,N_12333,N_13472);
nand U15429 (N_15429,N_13667,N_13167);
and U15430 (N_15430,N_13138,N_13272);
xor U15431 (N_15431,N_12913,N_12830);
xor U15432 (N_15432,N_12692,N_12199);
xor U15433 (N_15433,N_12362,N_12570);
nand U15434 (N_15434,N_12620,N_12515);
nand U15435 (N_15435,N_13360,N_13692);
nor U15436 (N_15436,N_12790,N_13920);
nand U15437 (N_15437,N_13522,N_13832);
nand U15438 (N_15438,N_12378,N_13752);
or U15439 (N_15439,N_13592,N_12348);
nor U15440 (N_15440,N_12202,N_13089);
xor U15441 (N_15441,N_13211,N_13765);
nor U15442 (N_15442,N_13267,N_12115);
or U15443 (N_15443,N_12663,N_12010);
nand U15444 (N_15444,N_13819,N_13981);
xor U15445 (N_15445,N_12968,N_12735);
nand U15446 (N_15446,N_13114,N_12670);
nor U15447 (N_15447,N_12312,N_12028);
or U15448 (N_15448,N_12804,N_12135);
nand U15449 (N_15449,N_13128,N_12417);
or U15450 (N_15450,N_12018,N_12914);
nand U15451 (N_15451,N_13094,N_13437);
xor U15452 (N_15452,N_13829,N_13277);
xor U15453 (N_15453,N_12894,N_13601);
xor U15454 (N_15454,N_13906,N_12200);
xnor U15455 (N_15455,N_12141,N_13993);
and U15456 (N_15456,N_13351,N_12611);
xor U15457 (N_15457,N_12327,N_13717);
nand U15458 (N_15458,N_12555,N_13137);
or U15459 (N_15459,N_12574,N_12073);
nand U15460 (N_15460,N_13363,N_12832);
nand U15461 (N_15461,N_13307,N_13202);
and U15462 (N_15462,N_12608,N_13658);
nand U15463 (N_15463,N_13557,N_13954);
nor U15464 (N_15464,N_13936,N_12068);
and U15465 (N_15465,N_12999,N_13774);
nor U15466 (N_15466,N_13412,N_13457);
xor U15467 (N_15467,N_13555,N_13501);
or U15468 (N_15468,N_12357,N_12637);
xnor U15469 (N_15469,N_13131,N_13790);
and U15470 (N_15470,N_12023,N_13725);
or U15471 (N_15471,N_12673,N_12983);
xnor U15472 (N_15472,N_13077,N_12109);
or U15473 (N_15473,N_13743,N_13058);
and U15474 (N_15474,N_13921,N_12162);
xor U15475 (N_15475,N_13300,N_12622);
or U15476 (N_15476,N_13928,N_13600);
and U15477 (N_15477,N_12145,N_12148);
nand U15478 (N_15478,N_13497,N_13926);
and U15479 (N_15479,N_12915,N_13353);
and U15480 (N_15480,N_13966,N_13856);
xor U15481 (N_15481,N_13268,N_12792);
nor U15482 (N_15482,N_13453,N_12078);
nand U15483 (N_15483,N_12795,N_12281);
and U15484 (N_15484,N_13693,N_12415);
xnor U15485 (N_15485,N_12585,N_12829);
and U15486 (N_15486,N_13634,N_12299);
nor U15487 (N_15487,N_13899,N_13871);
nand U15488 (N_15488,N_13668,N_13502);
nand U15489 (N_15489,N_13463,N_13723);
nand U15490 (N_15490,N_13955,N_12838);
and U15491 (N_15491,N_13897,N_12480);
nand U15492 (N_15492,N_12666,N_13372);
nor U15493 (N_15493,N_12138,N_12780);
and U15494 (N_15494,N_13734,N_13752);
nor U15495 (N_15495,N_12817,N_12134);
or U15496 (N_15496,N_12788,N_13526);
or U15497 (N_15497,N_13194,N_12878);
and U15498 (N_15498,N_13164,N_12771);
or U15499 (N_15499,N_13211,N_12243);
xnor U15500 (N_15500,N_12397,N_13090);
or U15501 (N_15501,N_12194,N_12067);
or U15502 (N_15502,N_13031,N_13939);
nand U15503 (N_15503,N_12984,N_12510);
nor U15504 (N_15504,N_12628,N_13003);
nor U15505 (N_15505,N_13414,N_12236);
or U15506 (N_15506,N_13205,N_13512);
nor U15507 (N_15507,N_13209,N_12501);
and U15508 (N_15508,N_12852,N_12778);
xnor U15509 (N_15509,N_13392,N_12471);
nor U15510 (N_15510,N_13000,N_12603);
or U15511 (N_15511,N_13995,N_13143);
nor U15512 (N_15512,N_13086,N_12108);
or U15513 (N_15513,N_13896,N_13026);
or U15514 (N_15514,N_12049,N_12914);
nand U15515 (N_15515,N_13248,N_13202);
or U15516 (N_15516,N_12565,N_12433);
xnor U15517 (N_15517,N_12544,N_12894);
and U15518 (N_15518,N_13278,N_13431);
and U15519 (N_15519,N_12886,N_12697);
xnor U15520 (N_15520,N_13418,N_13376);
and U15521 (N_15521,N_13321,N_13062);
xnor U15522 (N_15522,N_12839,N_13734);
nor U15523 (N_15523,N_13735,N_13285);
nor U15524 (N_15524,N_13154,N_12307);
nand U15525 (N_15525,N_13871,N_13033);
nor U15526 (N_15526,N_12057,N_12615);
and U15527 (N_15527,N_12305,N_12116);
nand U15528 (N_15528,N_13164,N_12441);
nand U15529 (N_15529,N_12162,N_12953);
nor U15530 (N_15530,N_13264,N_13016);
and U15531 (N_15531,N_12172,N_13212);
nor U15532 (N_15532,N_13472,N_12646);
nor U15533 (N_15533,N_13797,N_13682);
nor U15534 (N_15534,N_13537,N_13371);
nor U15535 (N_15535,N_13691,N_12597);
and U15536 (N_15536,N_13488,N_13661);
nor U15537 (N_15537,N_13597,N_12937);
nor U15538 (N_15538,N_12099,N_12443);
or U15539 (N_15539,N_13626,N_13453);
nand U15540 (N_15540,N_12142,N_13977);
and U15541 (N_15541,N_13386,N_13348);
xnor U15542 (N_15542,N_12742,N_13356);
xnor U15543 (N_15543,N_13458,N_13968);
xnor U15544 (N_15544,N_12246,N_12530);
nor U15545 (N_15545,N_13785,N_13563);
and U15546 (N_15546,N_12834,N_12517);
and U15547 (N_15547,N_13976,N_13741);
and U15548 (N_15548,N_13937,N_12559);
nor U15549 (N_15549,N_12500,N_13659);
or U15550 (N_15550,N_12545,N_13112);
nor U15551 (N_15551,N_13265,N_12033);
nand U15552 (N_15552,N_13087,N_12190);
nor U15553 (N_15553,N_13234,N_12101);
xor U15554 (N_15554,N_13389,N_12761);
and U15555 (N_15555,N_12006,N_13037);
and U15556 (N_15556,N_13736,N_13162);
or U15557 (N_15557,N_13333,N_13582);
and U15558 (N_15558,N_12216,N_13237);
and U15559 (N_15559,N_12758,N_12554);
nand U15560 (N_15560,N_13426,N_12501);
nand U15561 (N_15561,N_13475,N_12815);
xnor U15562 (N_15562,N_13535,N_13704);
or U15563 (N_15563,N_12008,N_13641);
or U15564 (N_15564,N_12861,N_13136);
or U15565 (N_15565,N_13978,N_12943);
or U15566 (N_15566,N_12135,N_13929);
nor U15567 (N_15567,N_13363,N_13917);
and U15568 (N_15568,N_13627,N_12191);
nand U15569 (N_15569,N_13591,N_12763);
nand U15570 (N_15570,N_12719,N_12510);
xor U15571 (N_15571,N_13704,N_12239);
nor U15572 (N_15572,N_13929,N_13687);
or U15573 (N_15573,N_12402,N_12501);
xor U15574 (N_15574,N_13175,N_13273);
and U15575 (N_15575,N_13679,N_12856);
nand U15576 (N_15576,N_12349,N_12106);
nor U15577 (N_15577,N_13845,N_13932);
nand U15578 (N_15578,N_12565,N_13150);
or U15579 (N_15579,N_12858,N_13374);
nor U15580 (N_15580,N_12820,N_13743);
nor U15581 (N_15581,N_13444,N_12412);
nand U15582 (N_15582,N_12362,N_13242);
nand U15583 (N_15583,N_13886,N_12182);
xnor U15584 (N_15584,N_12005,N_12599);
nor U15585 (N_15585,N_12381,N_13368);
xnor U15586 (N_15586,N_13568,N_12724);
nand U15587 (N_15587,N_13553,N_13861);
or U15588 (N_15588,N_13123,N_12157);
nor U15589 (N_15589,N_12438,N_13952);
nor U15590 (N_15590,N_12989,N_13235);
or U15591 (N_15591,N_13520,N_13807);
xnor U15592 (N_15592,N_12760,N_12892);
and U15593 (N_15593,N_13597,N_13986);
nand U15594 (N_15594,N_13735,N_12491);
and U15595 (N_15595,N_12152,N_12040);
xnor U15596 (N_15596,N_13423,N_13178);
nor U15597 (N_15597,N_12336,N_12325);
nor U15598 (N_15598,N_12108,N_12594);
nor U15599 (N_15599,N_12738,N_13969);
nor U15600 (N_15600,N_12451,N_13186);
xor U15601 (N_15601,N_13590,N_13752);
nand U15602 (N_15602,N_13359,N_13676);
xnor U15603 (N_15603,N_12361,N_13528);
xnor U15604 (N_15604,N_12141,N_13720);
or U15605 (N_15605,N_12638,N_12878);
nand U15606 (N_15606,N_12578,N_13396);
nand U15607 (N_15607,N_12958,N_13569);
or U15608 (N_15608,N_13868,N_13053);
nand U15609 (N_15609,N_13448,N_13479);
and U15610 (N_15610,N_12458,N_13555);
and U15611 (N_15611,N_13436,N_12830);
nor U15612 (N_15612,N_13128,N_13013);
or U15613 (N_15613,N_12485,N_12743);
or U15614 (N_15614,N_12426,N_12208);
and U15615 (N_15615,N_12708,N_12520);
nand U15616 (N_15616,N_13421,N_12645);
and U15617 (N_15617,N_13450,N_12469);
or U15618 (N_15618,N_13973,N_12379);
nand U15619 (N_15619,N_13752,N_12994);
nor U15620 (N_15620,N_13204,N_13990);
or U15621 (N_15621,N_12409,N_13335);
and U15622 (N_15622,N_13267,N_12689);
nor U15623 (N_15623,N_13505,N_12686);
nand U15624 (N_15624,N_12934,N_12008);
or U15625 (N_15625,N_12879,N_13498);
nand U15626 (N_15626,N_12331,N_13151);
xor U15627 (N_15627,N_12789,N_13641);
nand U15628 (N_15628,N_12816,N_13138);
or U15629 (N_15629,N_12463,N_13230);
xor U15630 (N_15630,N_13739,N_12347);
nand U15631 (N_15631,N_13321,N_13733);
nand U15632 (N_15632,N_12316,N_13993);
and U15633 (N_15633,N_13621,N_13464);
and U15634 (N_15634,N_12626,N_12639);
nand U15635 (N_15635,N_13319,N_12513);
nand U15636 (N_15636,N_13663,N_13358);
xor U15637 (N_15637,N_12809,N_12874);
xor U15638 (N_15638,N_12843,N_13221);
or U15639 (N_15639,N_13117,N_12512);
or U15640 (N_15640,N_12829,N_12519);
xnor U15641 (N_15641,N_13634,N_12173);
nor U15642 (N_15642,N_12891,N_12659);
and U15643 (N_15643,N_13729,N_13403);
and U15644 (N_15644,N_12458,N_12553);
or U15645 (N_15645,N_12512,N_12101);
xnor U15646 (N_15646,N_13973,N_13498);
and U15647 (N_15647,N_12363,N_12907);
xor U15648 (N_15648,N_12852,N_13928);
and U15649 (N_15649,N_13663,N_12273);
and U15650 (N_15650,N_13975,N_13448);
nor U15651 (N_15651,N_12034,N_12032);
xnor U15652 (N_15652,N_13769,N_13638);
xnor U15653 (N_15653,N_13542,N_13757);
and U15654 (N_15654,N_12814,N_12823);
and U15655 (N_15655,N_12660,N_13812);
nor U15656 (N_15656,N_12566,N_13497);
xnor U15657 (N_15657,N_13039,N_13310);
nand U15658 (N_15658,N_12598,N_13982);
or U15659 (N_15659,N_13267,N_12917);
and U15660 (N_15660,N_12018,N_12485);
or U15661 (N_15661,N_12238,N_13200);
xor U15662 (N_15662,N_12267,N_13622);
or U15663 (N_15663,N_13835,N_12877);
or U15664 (N_15664,N_12767,N_12125);
nand U15665 (N_15665,N_13096,N_12544);
xor U15666 (N_15666,N_12409,N_12526);
xnor U15667 (N_15667,N_13524,N_13169);
nor U15668 (N_15668,N_12091,N_12785);
or U15669 (N_15669,N_12984,N_13292);
xor U15670 (N_15670,N_12180,N_13303);
nor U15671 (N_15671,N_12434,N_13997);
nand U15672 (N_15672,N_13573,N_13311);
and U15673 (N_15673,N_12601,N_13789);
xnor U15674 (N_15674,N_13083,N_12923);
nand U15675 (N_15675,N_12127,N_13593);
and U15676 (N_15676,N_13889,N_13017);
or U15677 (N_15677,N_13876,N_12585);
and U15678 (N_15678,N_13914,N_12375);
and U15679 (N_15679,N_12056,N_13677);
nand U15680 (N_15680,N_12539,N_13356);
and U15681 (N_15681,N_13963,N_12403);
nor U15682 (N_15682,N_12832,N_13816);
and U15683 (N_15683,N_13364,N_12390);
and U15684 (N_15684,N_12192,N_13719);
and U15685 (N_15685,N_13444,N_12579);
and U15686 (N_15686,N_13751,N_13865);
and U15687 (N_15687,N_13871,N_13745);
or U15688 (N_15688,N_12079,N_13905);
xor U15689 (N_15689,N_12265,N_12695);
nor U15690 (N_15690,N_12219,N_12676);
xnor U15691 (N_15691,N_13592,N_13820);
xor U15692 (N_15692,N_12768,N_13575);
and U15693 (N_15693,N_12052,N_12712);
xnor U15694 (N_15694,N_13428,N_12266);
nand U15695 (N_15695,N_13858,N_12993);
and U15696 (N_15696,N_13446,N_12016);
xnor U15697 (N_15697,N_13835,N_12739);
nand U15698 (N_15698,N_12200,N_12583);
nand U15699 (N_15699,N_12826,N_13552);
or U15700 (N_15700,N_12984,N_13689);
xnor U15701 (N_15701,N_13438,N_13449);
xor U15702 (N_15702,N_12568,N_13781);
or U15703 (N_15703,N_13301,N_13044);
or U15704 (N_15704,N_12827,N_13523);
nor U15705 (N_15705,N_13231,N_12369);
or U15706 (N_15706,N_12705,N_13002);
xor U15707 (N_15707,N_12288,N_12902);
nand U15708 (N_15708,N_12817,N_12246);
nor U15709 (N_15709,N_13290,N_12912);
and U15710 (N_15710,N_13954,N_13357);
and U15711 (N_15711,N_12720,N_13957);
or U15712 (N_15712,N_12423,N_13086);
or U15713 (N_15713,N_12159,N_12405);
and U15714 (N_15714,N_12507,N_12640);
and U15715 (N_15715,N_12223,N_12665);
and U15716 (N_15716,N_12593,N_12809);
nor U15717 (N_15717,N_13072,N_13398);
or U15718 (N_15718,N_13300,N_13183);
nor U15719 (N_15719,N_13309,N_13265);
nor U15720 (N_15720,N_12449,N_12107);
xnor U15721 (N_15721,N_13077,N_12444);
nand U15722 (N_15722,N_12623,N_13233);
xor U15723 (N_15723,N_13155,N_12834);
or U15724 (N_15724,N_13686,N_13261);
nor U15725 (N_15725,N_12959,N_12068);
xor U15726 (N_15726,N_13939,N_12767);
nand U15727 (N_15727,N_12770,N_13799);
nor U15728 (N_15728,N_13951,N_13106);
nand U15729 (N_15729,N_12769,N_12487);
nand U15730 (N_15730,N_12776,N_12633);
nor U15731 (N_15731,N_13038,N_13609);
nand U15732 (N_15732,N_13651,N_13682);
nor U15733 (N_15733,N_12369,N_13527);
and U15734 (N_15734,N_12537,N_13735);
or U15735 (N_15735,N_12119,N_12676);
or U15736 (N_15736,N_13596,N_12770);
and U15737 (N_15737,N_12035,N_12008);
and U15738 (N_15738,N_12625,N_13144);
or U15739 (N_15739,N_13509,N_13016);
nor U15740 (N_15740,N_13635,N_12828);
or U15741 (N_15741,N_12769,N_12471);
xnor U15742 (N_15742,N_12539,N_13549);
nor U15743 (N_15743,N_12030,N_13116);
nor U15744 (N_15744,N_13455,N_13458);
and U15745 (N_15745,N_13457,N_13711);
nor U15746 (N_15746,N_13285,N_13817);
nor U15747 (N_15747,N_12295,N_12587);
or U15748 (N_15748,N_12169,N_13000);
or U15749 (N_15749,N_13498,N_13028);
nand U15750 (N_15750,N_12372,N_12480);
or U15751 (N_15751,N_13893,N_13186);
or U15752 (N_15752,N_12945,N_13939);
nor U15753 (N_15753,N_12510,N_12384);
or U15754 (N_15754,N_12253,N_12470);
xor U15755 (N_15755,N_12177,N_13877);
or U15756 (N_15756,N_13466,N_12803);
or U15757 (N_15757,N_13043,N_12898);
nor U15758 (N_15758,N_12687,N_13868);
or U15759 (N_15759,N_12720,N_12800);
nor U15760 (N_15760,N_12484,N_12070);
nor U15761 (N_15761,N_13279,N_12270);
and U15762 (N_15762,N_13725,N_12078);
or U15763 (N_15763,N_13842,N_13567);
or U15764 (N_15764,N_12773,N_12840);
nor U15765 (N_15765,N_12660,N_12463);
nand U15766 (N_15766,N_13359,N_12376);
nand U15767 (N_15767,N_12727,N_12722);
and U15768 (N_15768,N_12426,N_13955);
nor U15769 (N_15769,N_12663,N_12239);
or U15770 (N_15770,N_12885,N_13756);
nor U15771 (N_15771,N_12982,N_13484);
or U15772 (N_15772,N_13367,N_13455);
or U15773 (N_15773,N_12268,N_13638);
and U15774 (N_15774,N_12879,N_12008);
or U15775 (N_15775,N_12187,N_12741);
nor U15776 (N_15776,N_13228,N_13615);
or U15777 (N_15777,N_13240,N_13709);
nand U15778 (N_15778,N_13678,N_13977);
xnor U15779 (N_15779,N_13079,N_12277);
or U15780 (N_15780,N_12903,N_13395);
xor U15781 (N_15781,N_13094,N_12851);
and U15782 (N_15782,N_12455,N_13529);
xnor U15783 (N_15783,N_12193,N_13825);
nand U15784 (N_15784,N_12815,N_13481);
and U15785 (N_15785,N_13165,N_12375);
nor U15786 (N_15786,N_13011,N_13202);
xnor U15787 (N_15787,N_13023,N_13341);
and U15788 (N_15788,N_13366,N_12057);
nand U15789 (N_15789,N_12853,N_12287);
nor U15790 (N_15790,N_12796,N_12880);
and U15791 (N_15791,N_13053,N_13435);
xor U15792 (N_15792,N_12417,N_13157);
and U15793 (N_15793,N_13616,N_13660);
nor U15794 (N_15794,N_12888,N_12992);
nand U15795 (N_15795,N_12359,N_12332);
or U15796 (N_15796,N_13044,N_12172);
nor U15797 (N_15797,N_13357,N_12505);
nor U15798 (N_15798,N_13396,N_13104);
and U15799 (N_15799,N_12326,N_13033);
nand U15800 (N_15800,N_12636,N_13941);
and U15801 (N_15801,N_12526,N_13776);
nand U15802 (N_15802,N_12275,N_13720);
or U15803 (N_15803,N_12918,N_13323);
or U15804 (N_15804,N_13117,N_12000);
nand U15805 (N_15805,N_13936,N_13772);
nand U15806 (N_15806,N_12777,N_12903);
nand U15807 (N_15807,N_12533,N_13756);
nor U15808 (N_15808,N_13413,N_12636);
nor U15809 (N_15809,N_13671,N_13856);
nor U15810 (N_15810,N_13539,N_13569);
nor U15811 (N_15811,N_12993,N_13993);
and U15812 (N_15812,N_12508,N_13276);
and U15813 (N_15813,N_13148,N_13618);
nand U15814 (N_15814,N_12899,N_12529);
nor U15815 (N_15815,N_12815,N_12647);
nor U15816 (N_15816,N_12708,N_12338);
nor U15817 (N_15817,N_12032,N_13145);
or U15818 (N_15818,N_12102,N_13511);
xor U15819 (N_15819,N_13129,N_13117);
nand U15820 (N_15820,N_12398,N_13224);
nor U15821 (N_15821,N_12851,N_13381);
or U15822 (N_15822,N_12570,N_12337);
and U15823 (N_15823,N_12703,N_12314);
xnor U15824 (N_15824,N_13313,N_13817);
xnor U15825 (N_15825,N_13171,N_13198);
or U15826 (N_15826,N_12377,N_13026);
nor U15827 (N_15827,N_13260,N_12099);
xor U15828 (N_15828,N_12208,N_12560);
xor U15829 (N_15829,N_12622,N_13593);
nand U15830 (N_15830,N_12556,N_13925);
and U15831 (N_15831,N_13111,N_12995);
nor U15832 (N_15832,N_12334,N_13672);
nand U15833 (N_15833,N_12038,N_12433);
nand U15834 (N_15834,N_13206,N_12618);
and U15835 (N_15835,N_12882,N_13746);
xnor U15836 (N_15836,N_13307,N_12314);
and U15837 (N_15837,N_12720,N_12272);
nand U15838 (N_15838,N_13525,N_13529);
xor U15839 (N_15839,N_12473,N_13985);
and U15840 (N_15840,N_13068,N_13562);
xnor U15841 (N_15841,N_13912,N_12080);
and U15842 (N_15842,N_13187,N_12823);
nor U15843 (N_15843,N_12899,N_12338);
or U15844 (N_15844,N_13472,N_13516);
xnor U15845 (N_15845,N_12330,N_13938);
and U15846 (N_15846,N_13386,N_12478);
nor U15847 (N_15847,N_13786,N_12591);
and U15848 (N_15848,N_12973,N_12560);
or U15849 (N_15849,N_13274,N_13369);
xnor U15850 (N_15850,N_12330,N_13011);
and U15851 (N_15851,N_13565,N_12125);
nand U15852 (N_15852,N_13917,N_12816);
or U15853 (N_15853,N_12265,N_13861);
nor U15854 (N_15854,N_13831,N_12545);
nand U15855 (N_15855,N_12946,N_13671);
nor U15856 (N_15856,N_13418,N_12259);
nand U15857 (N_15857,N_12425,N_12081);
xnor U15858 (N_15858,N_13278,N_13378);
nand U15859 (N_15859,N_12802,N_12351);
nor U15860 (N_15860,N_13675,N_12975);
nor U15861 (N_15861,N_12066,N_12104);
nand U15862 (N_15862,N_13690,N_12561);
xnor U15863 (N_15863,N_13138,N_12725);
nor U15864 (N_15864,N_12469,N_13318);
xor U15865 (N_15865,N_13734,N_13499);
nand U15866 (N_15866,N_12307,N_13684);
nand U15867 (N_15867,N_13249,N_13245);
or U15868 (N_15868,N_12235,N_13416);
or U15869 (N_15869,N_12674,N_12625);
nand U15870 (N_15870,N_13493,N_13889);
or U15871 (N_15871,N_13090,N_13300);
nor U15872 (N_15872,N_12141,N_12968);
or U15873 (N_15873,N_13479,N_13054);
and U15874 (N_15874,N_13523,N_12406);
and U15875 (N_15875,N_12609,N_12692);
and U15876 (N_15876,N_13342,N_13726);
nor U15877 (N_15877,N_12238,N_12988);
and U15878 (N_15878,N_13665,N_13901);
xnor U15879 (N_15879,N_13063,N_13973);
or U15880 (N_15880,N_12536,N_13740);
nand U15881 (N_15881,N_13402,N_12608);
nand U15882 (N_15882,N_12814,N_12169);
and U15883 (N_15883,N_13471,N_12558);
and U15884 (N_15884,N_13774,N_12686);
nand U15885 (N_15885,N_13186,N_12285);
and U15886 (N_15886,N_12905,N_12957);
nor U15887 (N_15887,N_13154,N_13929);
nor U15888 (N_15888,N_13551,N_12554);
nor U15889 (N_15889,N_12273,N_13478);
xor U15890 (N_15890,N_12532,N_13097);
nor U15891 (N_15891,N_12410,N_12557);
nand U15892 (N_15892,N_12449,N_13478);
nor U15893 (N_15893,N_12820,N_13990);
nor U15894 (N_15894,N_12882,N_12039);
nand U15895 (N_15895,N_13081,N_12378);
xor U15896 (N_15896,N_12189,N_12568);
xnor U15897 (N_15897,N_13220,N_13151);
nand U15898 (N_15898,N_13157,N_13237);
and U15899 (N_15899,N_12295,N_12416);
or U15900 (N_15900,N_13826,N_12848);
xor U15901 (N_15901,N_13317,N_13310);
and U15902 (N_15902,N_13633,N_13228);
and U15903 (N_15903,N_13630,N_12105);
nand U15904 (N_15904,N_13464,N_12502);
or U15905 (N_15905,N_12148,N_13168);
or U15906 (N_15906,N_12923,N_13284);
and U15907 (N_15907,N_13477,N_12532);
or U15908 (N_15908,N_13862,N_13008);
and U15909 (N_15909,N_12371,N_13201);
nor U15910 (N_15910,N_12923,N_13606);
and U15911 (N_15911,N_12594,N_12805);
nand U15912 (N_15912,N_12671,N_13431);
and U15913 (N_15913,N_12654,N_13846);
nand U15914 (N_15914,N_12891,N_12691);
nand U15915 (N_15915,N_12373,N_13454);
nand U15916 (N_15916,N_13528,N_13498);
xnor U15917 (N_15917,N_13951,N_12682);
or U15918 (N_15918,N_13762,N_12833);
or U15919 (N_15919,N_12541,N_12412);
xor U15920 (N_15920,N_13037,N_12233);
xnor U15921 (N_15921,N_13331,N_13934);
nor U15922 (N_15922,N_13375,N_13859);
or U15923 (N_15923,N_13103,N_12952);
or U15924 (N_15924,N_12957,N_12665);
nand U15925 (N_15925,N_13587,N_12544);
or U15926 (N_15926,N_13124,N_12754);
or U15927 (N_15927,N_12737,N_13812);
nor U15928 (N_15928,N_12761,N_13550);
nand U15929 (N_15929,N_12204,N_13358);
xor U15930 (N_15930,N_12913,N_12641);
nor U15931 (N_15931,N_12916,N_12239);
and U15932 (N_15932,N_13017,N_13311);
nand U15933 (N_15933,N_13599,N_13687);
nand U15934 (N_15934,N_13202,N_12320);
and U15935 (N_15935,N_12746,N_13185);
nor U15936 (N_15936,N_12696,N_13578);
xor U15937 (N_15937,N_13006,N_13508);
nand U15938 (N_15938,N_12484,N_13421);
xor U15939 (N_15939,N_12301,N_13897);
nand U15940 (N_15940,N_12562,N_13597);
xor U15941 (N_15941,N_13010,N_12669);
nand U15942 (N_15942,N_13943,N_13548);
nor U15943 (N_15943,N_12368,N_12725);
nor U15944 (N_15944,N_13658,N_13628);
or U15945 (N_15945,N_12226,N_12999);
nor U15946 (N_15946,N_13655,N_12740);
xor U15947 (N_15947,N_12902,N_13816);
nand U15948 (N_15948,N_12159,N_12250);
nand U15949 (N_15949,N_13669,N_12914);
nand U15950 (N_15950,N_12222,N_13408);
nand U15951 (N_15951,N_13212,N_12733);
and U15952 (N_15952,N_12883,N_12650);
or U15953 (N_15953,N_13115,N_12889);
or U15954 (N_15954,N_13048,N_12552);
nand U15955 (N_15955,N_12020,N_12190);
nor U15956 (N_15956,N_13974,N_12085);
and U15957 (N_15957,N_13353,N_12835);
and U15958 (N_15958,N_13391,N_12589);
or U15959 (N_15959,N_12856,N_13747);
xnor U15960 (N_15960,N_12250,N_13700);
nor U15961 (N_15961,N_13850,N_12245);
nand U15962 (N_15962,N_12431,N_12781);
and U15963 (N_15963,N_12027,N_12072);
and U15964 (N_15964,N_12223,N_13984);
and U15965 (N_15965,N_12812,N_12352);
nor U15966 (N_15966,N_12431,N_12021);
nand U15967 (N_15967,N_13664,N_12852);
nand U15968 (N_15968,N_12119,N_12968);
and U15969 (N_15969,N_12673,N_12704);
or U15970 (N_15970,N_13693,N_13555);
or U15971 (N_15971,N_13014,N_13889);
nor U15972 (N_15972,N_12618,N_13430);
nand U15973 (N_15973,N_13696,N_12133);
nor U15974 (N_15974,N_13047,N_13067);
nor U15975 (N_15975,N_13896,N_12602);
nand U15976 (N_15976,N_13092,N_12618);
and U15977 (N_15977,N_12779,N_13074);
and U15978 (N_15978,N_13335,N_12181);
xnor U15979 (N_15979,N_13837,N_12907);
nand U15980 (N_15980,N_13004,N_12515);
and U15981 (N_15981,N_12916,N_12893);
or U15982 (N_15982,N_13742,N_13527);
xnor U15983 (N_15983,N_12440,N_13729);
nor U15984 (N_15984,N_12670,N_13065);
and U15985 (N_15985,N_12679,N_13752);
xnor U15986 (N_15986,N_13313,N_13157);
nand U15987 (N_15987,N_13984,N_12624);
nand U15988 (N_15988,N_12181,N_13152);
xnor U15989 (N_15989,N_12320,N_12688);
or U15990 (N_15990,N_12660,N_13667);
nor U15991 (N_15991,N_13469,N_12841);
nand U15992 (N_15992,N_12559,N_13472);
nor U15993 (N_15993,N_12916,N_12156);
nor U15994 (N_15994,N_12499,N_13570);
and U15995 (N_15995,N_13222,N_13077);
xor U15996 (N_15996,N_13719,N_12207);
nor U15997 (N_15997,N_12889,N_13722);
nand U15998 (N_15998,N_12038,N_12949);
nand U15999 (N_15999,N_12490,N_12252);
nor U16000 (N_16000,N_14319,N_14074);
nor U16001 (N_16001,N_14532,N_15482);
nor U16002 (N_16002,N_15571,N_15661);
nor U16003 (N_16003,N_15142,N_15486);
and U16004 (N_16004,N_14215,N_14525);
and U16005 (N_16005,N_15930,N_15502);
and U16006 (N_16006,N_15783,N_15311);
nand U16007 (N_16007,N_15401,N_14576);
xor U16008 (N_16008,N_14632,N_15043);
nor U16009 (N_16009,N_15594,N_14137);
xnor U16010 (N_16010,N_15505,N_15052);
and U16011 (N_16011,N_14340,N_14879);
and U16012 (N_16012,N_15682,N_15325);
and U16013 (N_16013,N_14551,N_15229);
and U16014 (N_16014,N_15789,N_15061);
nand U16015 (N_16015,N_15515,N_14564);
or U16016 (N_16016,N_15357,N_15485);
or U16017 (N_16017,N_14891,N_15901);
or U16018 (N_16018,N_14989,N_14219);
nor U16019 (N_16019,N_14958,N_15341);
and U16020 (N_16020,N_15655,N_14981);
nor U16021 (N_16021,N_14560,N_15751);
xnor U16022 (N_16022,N_14755,N_14933);
xor U16023 (N_16023,N_14617,N_14987);
xor U16024 (N_16024,N_15266,N_14880);
and U16025 (N_16025,N_14589,N_15034);
and U16026 (N_16026,N_14101,N_15340);
xor U16027 (N_16027,N_15808,N_15512);
or U16028 (N_16028,N_14012,N_14918);
nand U16029 (N_16029,N_15533,N_14250);
nor U16030 (N_16030,N_14552,N_15336);
and U16031 (N_16031,N_15902,N_15723);
or U16032 (N_16032,N_14407,N_15439);
nand U16033 (N_16033,N_15246,N_15601);
or U16034 (N_16034,N_14019,N_14457);
nor U16035 (N_16035,N_14896,N_15781);
nand U16036 (N_16036,N_15016,N_15890);
or U16037 (N_16037,N_15350,N_15648);
and U16038 (N_16038,N_14713,N_14009);
or U16039 (N_16039,N_14226,N_15787);
or U16040 (N_16040,N_14050,N_15529);
xor U16041 (N_16041,N_15245,N_14418);
or U16042 (N_16042,N_14485,N_15826);
nand U16043 (N_16043,N_14768,N_15907);
xnor U16044 (N_16044,N_14416,N_15123);
xnor U16045 (N_16045,N_14124,N_15164);
and U16046 (N_16046,N_15839,N_15276);
nand U16047 (N_16047,N_14373,N_15875);
xor U16048 (N_16048,N_15520,N_15656);
or U16049 (N_16049,N_14115,N_14053);
xnor U16050 (N_16050,N_14893,N_15924);
or U16051 (N_16051,N_14079,N_15690);
xor U16052 (N_16052,N_15898,N_14410);
nand U16053 (N_16053,N_14682,N_15095);
nand U16054 (N_16054,N_14433,N_15260);
xnor U16055 (N_16055,N_15014,N_15630);
or U16056 (N_16056,N_14609,N_15064);
and U16057 (N_16057,N_14696,N_14213);
or U16058 (N_16058,N_14583,N_15605);
or U16059 (N_16059,N_14098,N_14363);
nand U16060 (N_16060,N_14235,N_14973);
xor U16061 (N_16061,N_15835,N_15651);
nor U16062 (N_16062,N_14670,N_14310);
nor U16063 (N_16063,N_15855,N_14200);
and U16064 (N_16064,N_15730,N_15674);
nor U16065 (N_16065,N_15171,N_15582);
and U16066 (N_16066,N_14593,N_14761);
nand U16067 (N_16067,N_14287,N_14204);
xor U16068 (N_16068,N_14198,N_15560);
and U16069 (N_16069,N_15085,N_15137);
nor U16070 (N_16070,N_15188,N_15242);
xor U16071 (N_16071,N_14435,N_14106);
or U16072 (N_16072,N_15249,N_15030);
nand U16073 (N_16073,N_15870,N_14645);
nor U16074 (N_16074,N_14292,N_14983);
nand U16075 (N_16075,N_14470,N_15076);
nand U16076 (N_16076,N_15152,N_15319);
xnor U16077 (N_16077,N_14392,N_14205);
nor U16078 (N_16078,N_15672,N_14874);
nor U16079 (N_16079,N_14206,N_14188);
nand U16080 (N_16080,N_14661,N_15935);
nor U16081 (N_16081,N_14417,N_14312);
nor U16082 (N_16082,N_15255,N_14791);
or U16083 (N_16083,N_14174,N_14790);
xor U16084 (N_16084,N_15250,N_15253);
and U16085 (N_16085,N_15563,N_14045);
nand U16086 (N_16086,N_14163,N_14917);
and U16087 (N_16087,N_15827,N_15926);
or U16088 (N_16088,N_14212,N_15063);
or U16089 (N_16089,N_15905,N_14329);
xnor U16090 (N_16090,N_14674,N_15465);
xnor U16091 (N_16091,N_14280,N_15277);
nand U16092 (N_16092,N_15768,N_15252);
nor U16093 (N_16093,N_14068,N_15694);
and U16094 (N_16094,N_14949,N_14788);
nor U16095 (N_16095,N_15192,N_14863);
or U16096 (N_16096,N_14595,N_15603);
nor U16097 (N_16097,N_14716,N_14786);
nor U16098 (N_16098,N_14102,N_15284);
nor U16099 (N_16099,N_15353,N_14400);
and U16100 (N_16100,N_14151,N_14704);
nor U16101 (N_16101,N_14956,N_15286);
and U16102 (N_16102,N_14831,N_14377);
nand U16103 (N_16103,N_15722,N_14071);
xnor U16104 (N_16104,N_14652,N_14351);
or U16105 (N_16105,N_14527,N_14342);
nor U16106 (N_16106,N_14764,N_15693);
and U16107 (N_16107,N_14912,N_15203);
or U16108 (N_16108,N_15208,N_15066);
and U16109 (N_16109,N_14428,N_15844);
and U16110 (N_16110,N_14862,N_14272);
nand U16111 (N_16111,N_14133,N_15766);
and U16112 (N_16112,N_15770,N_14534);
xnor U16113 (N_16113,N_14544,N_15370);
nor U16114 (N_16114,N_15062,N_15200);
and U16115 (N_16115,N_14962,N_15632);
nand U16116 (N_16116,N_14675,N_15876);
or U16117 (N_16117,N_14636,N_14061);
nor U16118 (N_16118,N_14175,N_15814);
nor U16119 (N_16119,N_14107,N_15356);
or U16120 (N_16120,N_14922,N_15753);
nor U16121 (N_16121,N_14358,N_14669);
nor U16122 (N_16122,N_15071,N_15606);
or U16123 (N_16123,N_15704,N_14224);
or U16124 (N_16124,N_15960,N_14082);
nor U16125 (N_16125,N_15358,N_14461);
and U16126 (N_16126,N_14864,N_14847);
or U16127 (N_16127,N_15013,N_15925);
nand U16128 (N_16128,N_14253,N_15848);
xnor U16129 (N_16129,N_15927,N_15184);
nor U16130 (N_16130,N_14739,N_14815);
nor U16131 (N_16131,N_14998,N_15310);
or U16132 (N_16132,N_15005,N_14972);
nand U16133 (N_16133,N_14612,N_14376);
and U16134 (N_16134,N_15892,N_15148);
and U16135 (N_16135,N_14970,N_15000);
xor U16136 (N_16136,N_15012,N_14961);
nor U16137 (N_16137,N_15743,N_14699);
nor U16138 (N_16138,N_15989,N_14383);
xor U16139 (N_16139,N_14227,N_15338);
nand U16140 (N_16140,N_15039,N_14240);
nand U16141 (N_16141,N_15681,N_15920);
and U16142 (N_16142,N_15343,N_14315);
or U16143 (N_16143,N_14969,N_14619);
xnor U16144 (N_16144,N_15720,N_15718);
xnor U16145 (N_16145,N_14056,N_14828);
nor U16146 (N_16146,N_15498,N_15161);
xor U16147 (N_16147,N_15351,N_15469);
and U16148 (N_16148,N_15579,N_15049);
nor U16149 (N_16149,N_14776,N_14112);
nand U16150 (N_16150,N_14839,N_14386);
nor U16151 (N_16151,N_15938,N_14299);
nand U16152 (N_16152,N_15506,N_14694);
nor U16153 (N_16153,N_15423,N_15421);
and U16154 (N_16154,N_14466,N_15524);
nand U16155 (N_16155,N_15549,N_15492);
and U16156 (N_16156,N_14538,N_15050);
xor U16157 (N_16157,N_15238,N_14086);
and U16158 (N_16158,N_14714,N_15600);
xnor U16159 (N_16159,N_15257,N_14982);
xor U16160 (N_16160,N_15991,N_14024);
xnor U16161 (N_16161,N_14763,N_14710);
or U16162 (N_16162,N_14859,N_14677);
or U16163 (N_16163,N_14026,N_14231);
and U16164 (N_16164,N_14167,N_14925);
and U16165 (N_16165,N_15241,N_15265);
and U16166 (N_16166,N_14994,N_14873);
or U16167 (N_16167,N_15895,N_14297);
nand U16168 (N_16168,N_14084,N_14440);
xnor U16169 (N_16169,N_14246,N_14008);
xor U16170 (N_16170,N_14731,N_15141);
nand U16171 (N_16171,N_15510,N_15130);
nand U16172 (N_16172,N_15068,N_14742);
and U16173 (N_16173,N_14749,N_15503);
and U16174 (N_16174,N_15966,N_14812);
nor U16175 (N_16175,N_14622,N_15214);
nand U16176 (N_16176,N_15735,N_14031);
and U16177 (N_16177,N_14931,N_14401);
or U16178 (N_16178,N_15795,N_15422);
or U16179 (N_16179,N_14001,N_14087);
and U16180 (N_16180,N_15160,N_14996);
xnor U16181 (N_16181,N_15654,N_15324);
xor U16182 (N_16182,N_14181,N_15554);
xnor U16183 (N_16183,N_15390,N_14493);
xor U16184 (N_16184,N_14429,N_14268);
xnor U16185 (N_16185,N_15734,N_14035);
or U16186 (N_16186,N_15696,N_14284);
or U16187 (N_16187,N_14540,N_15596);
xnor U16188 (N_16188,N_14797,N_15897);
or U16189 (N_16189,N_14190,N_14968);
nor U16190 (N_16190,N_15174,N_14260);
or U16191 (N_16191,N_14692,N_15680);
nor U16192 (N_16192,N_15584,N_15282);
or U16193 (N_16193,N_14316,N_15083);
nor U16194 (N_16194,N_15060,N_15289);
nand U16195 (N_16195,N_14464,N_15536);
and U16196 (N_16196,N_15443,N_14676);
xnor U16197 (N_16197,N_15086,N_15132);
nor U16198 (N_16198,N_14060,N_15231);
nor U16199 (N_16199,N_15023,N_14562);
or U16200 (N_16200,N_14817,N_15225);
nor U16201 (N_16201,N_15806,N_14614);
nand U16202 (N_16202,N_15322,N_15263);
and U16203 (N_16203,N_15391,N_15084);
or U16204 (N_16204,N_15937,N_15106);
and U16205 (N_16205,N_15836,N_14225);
xor U16206 (N_16206,N_15215,N_14449);
nor U16207 (N_16207,N_15635,N_15593);
nand U16208 (N_16208,N_15793,N_14221);
nand U16209 (N_16209,N_14591,N_15149);
nand U16210 (N_16210,N_14179,N_15580);
nor U16211 (N_16211,N_15275,N_14502);
nor U16212 (N_16212,N_15928,N_15233);
or U16213 (N_16213,N_15569,N_15099);
and U16214 (N_16214,N_14057,N_14793);
or U16215 (N_16215,N_15900,N_14478);
nor U16216 (N_16216,N_15687,N_14085);
xor U16217 (N_16217,N_14604,N_15198);
nand U16218 (N_16218,N_14189,N_14594);
nor U16219 (N_16219,N_14556,N_14630);
and U16220 (N_16220,N_15824,N_14499);
nand U16221 (N_16221,N_14887,N_14536);
or U16222 (N_16222,N_15178,N_14999);
nor U16223 (N_16223,N_14802,N_15228);
and U16224 (N_16224,N_15355,N_14520);
or U16225 (N_16225,N_15139,N_14055);
and U16226 (N_16226,N_15756,N_14575);
xnor U16227 (N_16227,N_14930,N_14733);
and U16228 (N_16228,N_14463,N_15058);
xnor U16229 (N_16229,N_15135,N_14033);
xnor U16230 (N_16230,N_15678,N_15940);
and U16231 (N_16231,N_14004,N_15981);
nand U16232 (N_16232,N_15535,N_15755);
nand U16233 (N_16233,N_15679,N_15670);
xnor U16234 (N_16234,N_14805,N_15811);
nor U16235 (N_16235,N_14201,N_14770);
xor U16236 (N_16236,N_14446,N_15332);
nor U16237 (N_16237,N_14671,N_15543);
and U16238 (N_16238,N_14685,N_15491);
nor U16239 (N_16239,N_15978,N_15595);
nand U16240 (N_16240,N_15035,N_14191);
nor U16241 (N_16241,N_15096,N_15757);
xor U16242 (N_16242,N_15361,N_15407);
or U16243 (N_16243,N_15404,N_14715);
nor U16244 (N_16244,N_15020,N_15706);
and U16245 (N_16245,N_15763,N_15180);
or U16246 (N_16246,N_15446,N_15107);
or U16247 (N_16247,N_15965,N_15169);
xnor U16248 (N_16248,N_14217,N_15864);
xnor U16249 (N_16249,N_14244,N_14518);
or U16250 (N_16250,N_14803,N_14172);
xor U16251 (N_16251,N_15101,N_15080);
or U16252 (N_16252,N_15202,N_14984);
nor U16253 (N_16253,N_15954,N_14153);
nand U16254 (N_16254,N_15797,N_14585);
or U16255 (N_16255,N_14557,N_15758);
xor U16256 (N_16256,N_15660,N_14993);
or U16257 (N_16257,N_15312,N_14897);
nand U16258 (N_16258,N_15197,N_14991);
nand U16259 (N_16259,N_15326,N_14489);
xor U16260 (N_16260,N_15015,N_14357);
xor U16261 (N_16261,N_14195,N_15731);
and U16262 (N_16262,N_15963,N_14480);
and U16263 (N_16263,N_14236,N_15205);
or U16264 (N_16264,N_15344,N_14391);
and U16265 (N_16265,N_15158,N_14018);
nand U16266 (N_16266,N_15075,N_15652);
nand U16267 (N_16267,N_15568,N_15841);
nand U16268 (N_16268,N_14475,N_14458);
or U16269 (N_16269,N_14798,N_15140);
nand U16270 (N_16270,N_15955,N_15359);
nand U16271 (N_16271,N_15643,N_15074);
or U16272 (N_16272,N_14472,N_14159);
or U16273 (N_16273,N_14020,N_14114);
nand U16274 (N_16274,N_15967,N_15645);
xor U16275 (N_16275,N_14368,N_14281);
and U16276 (N_16276,N_14097,N_14597);
xor U16277 (N_16277,N_15663,N_14605);
nand U16278 (N_16278,N_14496,N_14131);
or U16279 (N_16279,N_15933,N_15547);
xnor U16280 (N_16280,N_15894,N_14963);
nor U16281 (N_16281,N_15379,N_15859);
or U16282 (N_16282,N_14596,N_14385);
nor U16283 (N_16283,N_15784,N_14384);
or U16284 (N_16284,N_15367,N_14599);
nor U16285 (N_16285,N_15377,N_15558);
xnor U16286 (N_16286,N_15832,N_15261);
or U16287 (N_16287,N_14929,N_14216);
xnor U16288 (N_16288,N_15126,N_14712);
xor U16289 (N_16289,N_14016,N_15114);
nand U16290 (N_16290,N_15460,N_14571);
nor U16291 (N_16291,N_14431,N_14992);
nand U16292 (N_16292,N_15154,N_15010);
nand U16293 (N_16293,N_15182,N_15226);
and U16294 (N_16294,N_15318,N_15669);
nand U16295 (N_16295,N_15749,N_14199);
xnor U16296 (N_16296,N_15611,N_15112);
nor U16297 (N_16297,N_15614,N_14708);
nand U16298 (N_16298,N_15285,N_14054);
nand U16299 (N_16299,N_14809,N_15659);
nand U16300 (N_16300,N_14078,N_14040);
and U16301 (N_16301,N_14794,N_14354);
and U16302 (N_16302,N_15153,N_14590);
nor U16303 (N_16303,N_15903,N_15666);
nor U16304 (N_16304,N_14081,N_14876);
or U16305 (N_16305,N_14834,N_15204);
nor U16306 (N_16306,N_14130,N_15576);
and U16307 (N_16307,N_15992,N_14323);
nor U16308 (N_16308,N_14664,N_14408);
xor U16309 (N_16309,N_15065,N_15179);
nand U16310 (N_16310,N_14214,N_14419);
and U16311 (N_16311,N_14286,N_15771);
xnor U16312 (N_16312,N_14207,N_14814);
nand U16313 (N_16313,N_14005,N_14379);
nand U16314 (N_16314,N_15544,N_14838);
or U16315 (N_16315,N_15251,N_15037);
xor U16316 (N_16316,N_15974,N_15767);
or U16317 (N_16317,N_15733,N_14883);
nor U16318 (N_16318,N_15562,N_15385);
nor U16319 (N_16319,N_14125,N_14077);
nor U16320 (N_16320,N_15009,N_14616);
nand U16321 (N_16321,N_14627,N_14550);
nand U16322 (N_16322,N_14023,N_14158);
or U16323 (N_16323,N_14454,N_15452);
and U16324 (N_16324,N_14187,N_14986);
nand U16325 (N_16325,N_14155,N_15473);
and U16326 (N_16326,N_15125,N_14491);
xnor U16327 (N_16327,N_14483,N_14600);
or U16328 (N_16328,N_14570,N_14196);
nor U16329 (N_16329,N_15923,N_14801);
nand U16330 (N_16330,N_15786,N_15438);
nor U16331 (N_16331,N_15742,N_14890);
or U16332 (N_16332,N_15858,N_14735);
xor U16333 (N_16333,N_15274,N_14683);
nor U16334 (N_16334,N_14402,N_15267);
or U16335 (N_16335,N_15412,N_15513);
xor U16336 (N_16336,N_14964,N_14277);
nand U16337 (N_16337,N_15293,N_14471);
xor U16338 (N_16338,N_14736,N_14412);
nand U16339 (N_16339,N_14309,N_14313);
xnor U16340 (N_16340,N_14854,N_15082);
xor U16341 (N_16341,N_15525,N_15383);
nand U16342 (N_16342,N_14398,N_15931);
nand U16343 (N_16343,N_15829,N_15805);
nor U16344 (N_16344,N_15024,N_14453);
and U16345 (N_16345,N_14903,N_14924);
and U16346 (N_16346,N_14635,N_15240);
nand U16347 (N_16347,N_15586,N_14043);
xnor U16348 (N_16348,N_14719,N_15166);
or U16349 (N_16349,N_14047,N_15780);
nor U16350 (N_16350,N_14651,N_14288);
nor U16351 (N_16351,N_15769,N_15468);
xor U16352 (N_16352,N_15921,N_14051);
xnor U16353 (N_16353,N_14729,N_15975);
nor U16354 (N_16354,N_14840,N_15511);
nor U16355 (N_16355,N_14065,N_15219);
and U16356 (N_16356,N_14751,N_14946);
xor U16357 (N_16357,N_15583,N_14516);
and U16358 (N_16358,N_15480,N_14180);
or U16359 (N_16359,N_15910,N_14041);
xnor U16360 (N_16360,N_15941,N_15857);
or U16361 (N_16361,N_15364,N_15707);
nor U16362 (N_16362,N_14509,N_14448);
or U16363 (N_16363,N_14680,N_14484);
and U16364 (N_16364,N_14775,N_15919);
and U16365 (N_16365,N_14531,N_14730);
or U16366 (N_16366,N_15629,N_14422);
xnor U16367 (N_16367,N_14586,N_15761);
and U16368 (N_16368,N_14545,N_15887);
xor U16369 (N_16369,N_14278,N_15235);
nand U16370 (N_16370,N_15778,N_15541);
or U16371 (N_16371,N_14951,N_14711);
and U16372 (N_16372,N_15737,N_14662);
nor U16373 (N_16373,N_14271,N_14378);
nor U16374 (N_16374,N_15397,N_14262);
xor U16375 (N_16375,N_14149,N_14177);
nand U16376 (N_16376,N_14362,N_14083);
nor U16377 (N_16377,N_14765,N_15962);
and U16378 (N_16378,N_14420,N_14306);
nor U16379 (N_16379,N_14783,N_14346);
nor U16380 (N_16380,N_14942,N_15913);
nor U16381 (N_16381,N_14663,N_14767);
nand U16382 (N_16382,N_15155,N_14166);
or U16383 (N_16383,N_14257,N_14366);
xnor U16384 (N_16384,N_14760,N_14811);
and U16385 (N_16385,N_15048,N_14853);
xor U16386 (N_16386,N_14073,N_15741);
or U16387 (N_16387,N_14935,N_15157);
or U16388 (N_16388,N_15922,N_15990);
nor U16389 (N_16389,N_14526,N_15297);
or U16390 (N_16390,N_15320,N_14923);
xnor U16391 (N_16391,N_14787,N_14587);
nor U16392 (N_16392,N_15295,N_14553);
or U16393 (N_16393,N_15456,N_14360);
and U16394 (N_16394,N_14965,N_15042);
or U16395 (N_16395,N_15948,N_15879);
or U16396 (N_16396,N_14267,N_14608);
nor U16397 (N_16397,N_15360,N_15163);
nand U16398 (N_16398,N_14171,N_14176);
nor U16399 (N_16399,N_14256,N_15059);
nand U16400 (N_16400,N_14707,N_14744);
and U16401 (N_16401,N_15017,N_15958);
nand U16402 (N_16402,N_14184,N_15462);
nand U16403 (N_16403,N_14654,N_15791);
xnor U16404 (N_16404,N_15402,N_15574);
or U16405 (N_16405,N_15070,N_14845);
nor U16406 (N_16406,N_14655,N_14255);
nand U16407 (N_16407,N_14233,N_14826);
or U16408 (N_16408,N_14906,N_14795);
xor U16409 (N_16409,N_15287,N_14328);
xor U16410 (N_16410,N_15712,N_15956);
and U16411 (N_16411,N_14613,N_14944);
xnor U16412 (N_16412,N_14285,N_14487);
xor U16413 (N_16413,N_14036,N_14537);
and U16414 (N_16414,N_15715,N_15838);
xor U16415 (N_16415,N_15862,N_14959);
nor U16416 (N_16416,N_15463,N_14533);
and U16417 (N_16417,N_14170,N_15500);
xor U16418 (N_16418,N_14741,N_14111);
nor U16419 (N_16419,N_15381,N_15038);
and U16420 (N_16420,N_14169,N_14558);
nor U16421 (N_16421,N_14481,N_15077);
and U16422 (N_16422,N_14905,N_15572);
and U16423 (N_16423,N_15342,N_15081);
and U16424 (N_16424,N_15530,N_15514);
nand U16425 (N_16425,N_15256,N_14067);
and U16426 (N_16426,N_14252,N_14220);
nor U16427 (N_16427,N_14620,N_14870);
nand U16428 (N_16428,N_14581,N_14872);
or U16429 (N_16429,N_15888,N_15110);
and U16430 (N_16430,N_14218,N_15980);
or U16431 (N_16431,N_15054,N_14772);
nor U16432 (N_16432,N_15258,N_15776);
nor U16433 (N_16433,N_15994,N_15244);
nor U16434 (N_16434,N_14697,N_15453);
nand U16435 (N_16435,N_15833,N_15847);
nand U16436 (N_16436,N_15615,N_15705);
or U16437 (N_16437,N_14091,N_15591);
or U16438 (N_16438,N_14985,N_14274);
or U16439 (N_16439,N_15053,N_14681);
or U16440 (N_16440,N_15429,N_14724);
nand U16441 (N_16441,N_14535,N_14606);
nor U16442 (N_16442,N_15531,N_14460);
nand U16443 (N_16443,N_14465,N_15882);
and U16444 (N_16444,N_15909,N_14726);
xor U16445 (N_16445,N_14211,N_14348);
nor U16446 (N_16446,N_14186,N_15458);
and U16447 (N_16447,N_14479,N_14565);
xnor U16448 (N_16448,N_15891,N_14781);
or U16449 (N_16449,N_14350,N_15072);
nor U16450 (N_16450,N_15395,N_15116);
or U16451 (N_16451,N_14232,N_14030);
xor U16452 (N_16452,N_15764,N_15585);
nand U16453 (N_16453,N_14455,N_15658);
and U16454 (N_16454,N_15291,N_14601);
nand U16455 (N_16455,N_14249,N_15995);
xnor U16456 (N_16456,N_15747,N_15883);
and U16457 (N_16457,N_14147,N_15548);
and U16458 (N_16458,N_15561,N_14995);
nor U16459 (N_16459,N_14103,N_14549);
xor U16460 (N_16460,N_14421,N_14720);
nor U16461 (N_16461,N_15527,N_14052);
and U16462 (N_16462,N_15392,N_14754);
and U16463 (N_16463,N_14325,N_15186);
xor U16464 (N_16464,N_14443,N_14424);
xnor U16465 (N_16465,N_14395,N_14150);
or U16466 (N_16466,N_15803,N_15633);
or U16467 (N_16467,N_14672,N_14359);
nor U16468 (N_16468,N_15959,N_14894);
nor U16469 (N_16469,N_15363,N_15851);
nand U16470 (N_16470,N_15650,N_15002);
nor U16471 (N_16471,N_15842,N_15637);
nor U16472 (N_16472,N_14279,N_15380);
or U16473 (N_16473,N_15971,N_14966);
or U16474 (N_16474,N_15435,N_15430);
xnor U16475 (N_16475,N_14469,N_14957);
nand U16476 (N_16476,N_14841,N_14554);
nor U16477 (N_16477,N_15415,N_14975);
nand U16478 (N_16478,N_15794,N_14135);
nand U16479 (N_16479,N_14173,N_14732);
or U16480 (N_16480,N_15268,N_14911);
xnor U16481 (N_16481,N_14762,N_15352);
nor U16482 (N_16482,N_14241,N_15952);
and U16483 (N_16483,N_14641,N_14851);
nand U16484 (N_16484,N_15713,N_15055);
nand U16485 (N_16485,N_14437,N_14820);
and U16486 (N_16486,N_15775,N_14633);
xor U16487 (N_16487,N_15211,N_15728);
xor U16488 (N_16488,N_15212,N_14816);
xnor U16489 (N_16489,N_14152,N_14514);
nor U16490 (N_16490,N_14611,N_14588);
xor U16491 (N_16491,N_15045,N_14746);
or U16492 (N_16492,N_14546,N_15998);
or U16493 (N_16493,N_14178,N_14517);
nor U16494 (N_16494,N_15945,N_15812);
or U16495 (N_16495,N_15011,N_15863);
xor U16496 (N_16496,N_15934,N_14773);
nor U16497 (N_16497,N_15671,N_14568);
and U16498 (N_16498,N_14182,N_15523);
or U16499 (N_16499,N_15738,N_15201);
xor U16500 (N_16500,N_14117,N_14938);
or U16501 (N_16501,N_14778,N_14881);
nor U16502 (N_16502,N_15032,N_14850);
nand U16503 (N_16503,N_14647,N_14860);
nand U16504 (N_16504,N_14066,N_15714);
or U16505 (N_16505,N_14193,N_14021);
xnor U16506 (N_16506,N_15427,N_14940);
and U16507 (N_16507,N_14361,N_15478);
nand U16508 (N_16508,N_14245,N_15471);
nor U16509 (N_16509,N_14784,N_14042);
and U16510 (N_16510,N_15914,N_15224);
nor U16511 (N_16511,N_14058,N_15779);
nand U16512 (N_16512,N_15969,N_15001);
nand U16513 (N_16513,N_14307,N_15540);
or U16514 (N_16514,N_15484,N_15816);
nand U16515 (N_16515,N_14495,N_14028);
xnor U16516 (N_16516,N_14476,N_14119);
or U16517 (N_16517,N_15475,N_15399);
and U16518 (N_16518,N_14118,N_15156);
or U16519 (N_16519,N_15942,N_14341);
or U16520 (N_16520,N_15589,N_15944);
or U16521 (N_16521,N_14702,N_14251);
and U16522 (N_16522,N_14559,N_15303);
and U16523 (N_16523,N_14618,N_14497);
nor U16524 (N_16524,N_14919,N_14806);
nand U16525 (N_16525,N_15398,N_15296);
xor U16526 (N_16526,N_15098,N_15018);
nand U16527 (N_16527,N_14819,N_15067);
and U16528 (N_16528,N_15634,N_15624);
nor U16529 (N_16529,N_14679,N_14785);
and U16530 (N_16530,N_15599,N_15418);
nor U16531 (N_16531,N_14411,N_15474);
nand U16532 (N_16532,N_14301,N_14441);
xor U16533 (N_16533,N_15581,N_14907);
nand U16534 (N_16534,N_14771,N_15159);
xor U16535 (N_16535,N_14322,N_14978);
and U16536 (N_16536,N_15004,N_15993);
nand U16537 (N_16537,N_14748,N_14920);
and U16538 (N_16538,N_15092,N_14844);
nor U16539 (N_16539,N_15866,N_15748);
xnor U16540 (N_16540,N_14639,N_15647);
nand U16541 (N_16541,N_14910,N_14039);
nand U16542 (N_16542,N_15698,N_15578);
and U16543 (N_16543,N_15167,N_14709);
xnor U16544 (N_16544,N_15248,N_15646);
nand U16545 (N_16545,N_14242,N_14503);
nand U16546 (N_16546,N_14011,N_15454);
and U16547 (N_16547,N_15968,N_14542);
and U16548 (N_16548,N_14988,N_15987);
or U16549 (N_16549,N_15825,N_14034);
nand U16550 (N_16550,N_14157,N_15437);
nand U16551 (N_16551,N_15221,N_15517);
nor U16552 (N_16552,N_15729,N_14238);
or U16553 (N_16553,N_14302,N_15988);
nor U16554 (N_16554,N_14291,N_15622);
and U16555 (N_16555,N_15041,N_15191);
or U16556 (N_16556,N_15301,N_15328);
and U16557 (N_16557,N_14515,N_14311);
xnor U16558 (N_16558,N_14168,N_14387);
and U16559 (N_16559,N_14892,N_15555);
xnor U16560 (N_16560,N_15684,N_15104);
and U16561 (N_16561,N_15709,N_14276);
nand U16562 (N_16562,N_15288,N_15732);
and U16563 (N_16563,N_15716,N_14474);
nand U16564 (N_16564,N_15300,N_14752);
or U16565 (N_16565,N_15830,N_15809);
xnor U16566 (N_16566,N_15368,N_15686);
and U16567 (N_16567,N_14868,N_14504);
nor U16568 (N_16568,N_14566,N_15602);
nand U16569 (N_16569,N_15818,N_15801);
or U16570 (N_16570,N_15745,N_14136);
xor U16571 (N_16571,N_14528,N_15317);
and U16572 (N_16572,N_14865,N_14473);
and U16573 (N_16573,N_15853,N_14108);
nor U16574 (N_16574,N_14740,N_14955);
nand U16575 (N_16575,N_15871,N_15997);
xor U16576 (N_16576,N_14294,N_15662);
and U16577 (N_16577,N_15929,N_15269);
or U16578 (N_16578,N_14976,N_14547);
nand U16579 (N_16579,N_14070,N_14888);
or U16580 (N_16580,N_15347,N_15610);
nand U16581 (N_16581,N_14832,N_14822);
nand U16582 (N_16582,N_14727,N_14336);
xor U16583 (N_16583,N_14367,N_14582);
nand U16584 (N_16584,N_14861,N_14634);
xor U16585 (N_16585,N_15136,N_14837);
and U16586 (N_16586,N_15828,N_15823);
or U16587 (N_16587,N_14657,N_14427);
and U16588 (N_16588,N_15393,N_14967);
and U16589 (N_16589,N_14725,N_14110);
nand U16590 (N_16590,N_15947,N_14327);
xor U16591 (N_16591,N_15436,N_15145);
xnor U16592 (N_16592,N_14388,N_14782);
xnor U16593 (N_16593,N_14263,N_15575);
nor U16594 (N_16594,N_14369,N_15683);
and U16595 (N_16595,N_14849,N_14698);
xnor U16596 (N_16596,N_14197,N_15754);
nand U16597 (N_16597,N_15330,N_14825);
nand U16598 (N_16598,N_14842,N_15939);
and U16599 (N_16599,N_15612,N_15649);
nor U16600 (N_16600,N_14898,N_14637);
or U16601 (N_16601,N_14304,N_15725);
or U16602 (N_16602,N_15127,N_14403);
nor U16603 (N_16603,N_14908,N_15115);
xor U16604 (N_16604,N_15964,N_15493);
and U16605 (N_16605,N_14414,N_15384);
nand U16606 (N_16606,N_15532,N_15321);
xor U16607 (N_16607,N_14722,N_14062);
or U16608 (N_16608,N_14653,N_15079);
nand U16609 (N_16609,N_14140,N_15607);
nand U16610 (N_16610,N_14703,N_15762);
or U16611 (N_16611,N_15522,N_14977);
xnor U16612 (N_16612,N_15736,N_14122);
nand U16613 (N_16613,N_15566,N_15457);
nand U16614 (N_16614,N_14393,N_14813);
nor U16615 (N_16615,N_14413,N_15129);
xor U16616 (N_16616,N_14574,N_15676);
nand U16617 (N_16617,N_15983,N_15122);
xor U16618 (N_16618,N_14756,N_14258);
nor U16619 (N_16619,N_15817,N_14759);
xor U16620 (N_16620,N_15376,N_15592);
nor U16621 (N_16621,N_14185,N_14567);
or U16622 (N_16622,N_15711,N_15984);
or U16623 (N_16623,N_15867,N_14505);
and U16624 (N_16624,N_15752,N_15893);
or U16625 (N_16625,N_15102,N_15621);
xor U16626 (N_16626,N_14138,N_14332);
or U16627 (N_16627,N_15886,N_14769);
and U16628 (N_16628,N_15477,N_14728);
or U16629 (N_16629,N_14230,N_14548);
nor U16630 (N_16630,N_15528,N_15590);
or U16631 (N_16631,N_15986,N_15047);
nand U16632 (N_16632,N_14830,N_15917);
and U16633 (N_16633,N_15144,N_14640);
nor U16634 (N_16634,N_15588,N_15073);
nor U16635 (N_16635,N_15627,N_14953);
xnor U16636 (N_16636,N_15413,N_15165);
or U16637 (N_16637,N_14904,N_14690);
nor U16638 (N_16638,N_14430,N_15623);
and U16639 (N_16639,N_15701,N_15209);
or U16640 (N_16640,N_14330,N_15587);
or U16641 (N_16641,N_14273,N_14511);
xor U16642 (N_16642,N_15218,N_14821);
or U16643 (N_16643,N_15950,N_15470);
and U16644 (N_16644,N_14592,N_15479);
nand U16645 (N_16645,N_15488,N_14208);
nand U16646 (N_16646,N_14818,N_14080);
or U16647 (N_16647,N_15820,N_14451);
or U16648 (N_16648,N_15837,N_14952);
nor U16649 (N_16649,N_15567,N_15176);
or U16650 (N_16650,N_15750,N_15570);
nand U16651 (N_16651,N_15057,N_14094);
and U16652 (N_16652,N_15868,N_14295);
nor U16653 (N_16653,N_15109,N_15911);
or U16654 (N_16654,N_15509,N_15915);
xor U16655 (N_16655,N_14658,N_14927);
nor U16656 (N_16656,N_14934,N_14990);
nand U16657 (N_16657,N_14405,N_14869);
nand U16658 (N_16658,N_15175,N_14807);
and U16659 (N_16659,N_15117,N_15845);
xnor U16660 (N_16660,N_14660,N_14374);
nor U16661 (N_16661,N_14561,N_15597);
nor U16662 (N_16662,N_14399,N_15916);
or U16663 (N_16663,N_14015,N_15119);
nor U16664 (N_16664,N_14723,N_15673);
xnor U16665 (N_16665,N_15031,N_15664);
xor U16666 (N_16666,N_14901,N_15765);
xnor U16667 (N_16667,N_15642,N_15675);
nand U16668 (N_16668,N_14165,N_14774);
or U16669 (N_16669,N_15772,N_15128);
nand U16670 (N_16670,N_14445,N_15433);
xnor U16671 (N_16671,N_15327,N_14506);
xnor U16672 (N_16672,N_15354,N_14095);
or U16673 (N_16673,N_14239,N_15943);
nor U16674 (N_16674,N_15481,N_15410);
nor U16675 (N_16675,N_14293,N_14121);
or U16676 (N_16676,N_15834,N_15304);
or U16677 (N_16677,N_15162,N_15299);
or U16678 (N_16678,N_15760,N_15519);
nor U16679 (N_16679,N_14321,N_15424);
xnor U16680 (N_16680,N_14161,N_15170);
nand U16681 (N_16681,N_14300,N_14579);
xnor U16682 (N_16682,N_14006,N_14678);
xnor U16683 (N_16683,N_15335,N_15207);
or U16684 (N_16684,N_15790,N_15850);
or U16685 (N_16685,N_14444,N_14750);
xnor U16686 (N_16686,N_15906,N_14827);
nor U16687 (N_16687,N_15441,N_14510);
xor U16688 (N_16688,N_15849,N_15653);
xnor U16689 (N_16689,N_14758,N_15313);
nand U16690 (N_16690,N_15227,N_15247);
or U16691 (N_16691,N_14623,N_15665);
or U16692 (N_16692,N_15134,N_14687);
xnor U16693 (N_16693,N_15877,N_15362);
xor U16694 (N_16694,N_15348,N_14317);
or U16695 (N_16695,N_15187,N_14456);
nor U16696 (N_16696,N_15177,N_15088);
nor U16697 (N_16697,N_15281,N_15708);
nor U16698 (N_16698,N_14308,N_14882);
and U16699 (N_16699,N_15490,N_15608);
and U16700 (N_16700,N_15537,N_14524);
nand U16701 (N_16701,N_15796,N_14442);
and U16702 (N_16702,N_14423,N_14909);
nand U16703 (N_16703,N_14700,N_15173);
and U16704 (N_16704,N_15843,N_15279);
nand U16705 (N_16705,N_14088,N_15026);
nand U16706 (N_16706,N_14123,N_15270);
nor U16707 (N_16707,N_14222,N_14254);
nor U16708 (N_16708,N_14871,N_15953);
nor U16709 (N_16709,N_15860,N_14848);
nor U16710 (N_16710,N_14914,N_15545);
nor U16711 (N_16711,N_14027,N_15387);
nand U16712 (N_16712,N_14092,N_14686);
nor U16713 (N_16713,N_14650,N_14500);
or U16714 (N_16714,N_14432,N_14298);
and U16715 (N_16715,N_15210,N_15272);
nor U16716 (N_16716,N_14303,N_15262);
nand U16717 (N_16717,N_14621,N_15006);
xor U16718 (N_16718,N_15613,N_15951);
xnor U16719 (N_16719,N_15334,N_15996);
nand U16720 (N_16720,N_14684,N_15003);
and U16721 (N_16721,N_14142,N_14210);
nor U16722 (N_16722,N_15028,N_15216);
nand U16723 (N_16723,N_14044,N_14345);
nor U16724 (N_16724,N_14936,N_14799);
nor U16725 (N_16725,N_15314,N_15259);
and U16726 (N_16726,N_14248,N_14371);
xnor U16727 (N_16727,N_15056,N_14148);
nand U16728 (N_16728,N_14529,N_14997);
nor U16729 (N_16729,N_15577,N_14025);
and U16730 (N_16730,N_14048,N_15551);
nand U16731 (N_16731,N_14928,N_15744);
nand U16732 (N_16732,N_15078,N_14326);
nand U16733 (N_16733,N_15044,N_15172);
xor U16734 (N_16734,N_14569,N_15440);
and U16735 (N_16735,N_15403,N_15626);
nand U16736 (N_16736,N_15869,N_14380);
and U16737 (N_16737,N_15396,N_15239);
nand U16738 (N_16738,N_14522,N_14264);
nand U16739 (N_16739,N_15912,N_15113);
xnor U16740 (N_16740,N_14665,N_15337);
or U16741 (N_16741,N_14002,N_14501);
nor U16742 (N_16742,N_14508,N_15556);
xor U16743 (N_16743,N_15936,N_14649);
or U16744 (N_16744,N_15451,N_14829);
and U16745 (N_16745,N_14160,N_15199);
or U16746 (N_16746,N_15521,N_14902);
xnor U16747 (N_16747,N_15417,N_14467);
nand U16748 (N_16748,N_15483,N_14810);
and U16749 (N_16749,N_14305,N_15051);
nand U16750 (N_16750,N_15147,N_14290);
nor U16751 (N_16751,N_15371,N_14339);
nand U16752 (N_16752,N_15822,N_15138);
xnor U16753 (N_16753,N_14624,N_14096);
xor U16754 (N_16754,N_14789,N_14247);
xnor U16755 (N_16755,N_15499,N_15131);
nor U16756 (N_16756,N_15036,N_14498);
or U16757 (N_16757,N_14667,N_15217);
nand U16758 (N_16758,N_14884,N_14120);
xor U16759 (N_16759,N_15151,N_14779);
xnor U16760 (N_16760,N_14404,N_14856);
or U16761 (N_16761,N_14229,N_15339);
xnor U16762 (N_16762,N_14000,N_15872);
nor U16763 (N_16763,N_15069,N_14318);
xor U16764 (N_16764,N_14948,N_15461);
nor U16765 (N_16765,N_14146,N_14415);
and U16766 (N_16766,N_15497,N_14693);
nor U16767 (N_16767,N_15516,N_15699);
xor U16768 (N_16768,N_15222,N_15386);
or U16769 (N_16769,N_14857,N_14916);
nand U16770 (N_16770,N_15450,N_15021);
xnor U16771 (N_16771,N_15168,N_15400);
or U16772 (N_16772,N_14625,N_14780);
and U16773 (N_16773,N_14334,N_14691);
xnor U16774 (N_16774,N_15254,N_15243);
nor U16775 (N_16775,N_14104,N_14488);
xnor U16776 (N_16776,N_15972,N_14331);
nor U16777 (N_16777,N_14324,N_15298);
nand U16778 (N_16778,N_15985,N_14643);
nand U16779 (N_16779,N_14932,N_15856);
xnor U16780 (N_16780,N_14757,N_14603);
xnor U16781 (N_16781,N_14356,N_15885);
and U16782 (N_16782,N_14013,N_15366);
and U16783 (N_16783,N_14846,N_15346);
nor U16784 (N_16784,N_15973,N_15408);
nor U16785 (N_16785,N_14979,N_14734);
or U16786 (N_16786,N_14543,N_15703);
nand U16787 (N_16787,N_14941,N_14265);
and U16788 (N_16788,N_15195,N_14076);
xnor U16789 (N_16789,N_15746,N_15309);
nor U16790 (N_16790,N_14494,N_14396);
and U16791 (N_16791,N_15278,N_15007);
nand U16792 (N_16792,N_15798,N_15183);
or U16793 (N_16793,N_14915,N_15466);
nor U16794 (N_16794,N_14134,N_14833);
nor U16795 (N_16795,N_15861,N_15121);
nand U16796 (N_16796,N_14629,N_14875);
or U16797 (N_16797,N_15315,N_14243);
or U16798 (N_16798,N_14852,N_14800);
nand U16799 (N_16799,N_15774,N_14075);
nor U16800 (N_16800,N_15565,N_15918);
or U16801 (N_16801,N_14093,N_15782);
xor U16802 (N_16802,N_14409,N_14156);
nor U16803 (N_16803,N_14659,N_14296);
or U16804 (N_16804,N_15416,N_15874);
nor U16805 (N_16805,N_15374,N_14541);
nor U16806 (N_16806,N_14394,N_14046);
xnor U16807 (N_16807,N_15349,N_14628);
or U16808 (N_16808,N_14109,N_15306);
and U16809 (N_16809,N_14689,N_15496);
nand U16810 (N_16810,N_15815,N_15946);
nor U16811 (N_16811,N_14843,N_14116);
nor U16812 (N_16812,N_15290,N_15025);
or U16813 (N_16813,N_14447,N_15878);
nor U16814 (N_16814,N_15472,N_15089);
xnor U16815 (N_16815,N_14573,N_15237);
and U16816 (N_16816,N_14100,N_15316);
xor U16817 (N_16817,N_15542,N_14438);
nor U16818 (N_16818,N_14521,N_15695);
or U16819 (N_16819,N_14164,N_14038);
or U16820 (N_16820,N_14766,N_15090);
and U16821 (N_16821,N_15206,N_14059);
and U16822 (N_16822,N_15464,N_14889);
xnor U16823 (N_16823,N_15889,N_14482);
or U16824 (N_16824,N_14141,N_15378);
nor U16825 (N_16825,N_14090,N_15873);
nand U16826 (N_16826,N_15196,N_14261);
xnor U16827 (N_16827,N_14512,N_15840);
nand U16828 (N_16828,N_14718,N_15557);
xnor U16829 (N_16829,N_15305,N_14382);
and U16830 (N_16830,N_15365,N_14926);
or U16831 (N_16831,N_15097,N_14738);
or U16832 (N_16832,N_15976,N_14347);
and U16833 (N_16833,N_15677,N_14646);
or U16834 (N_16834,N_14202,N_14642);
xnor U16835 (N_16835,N_15372,N_15657);
xor U16836 (N_16836,N_15949,N_15425);
xor U16837 (N_16837,N_14234,N_14450);
nor U16838 (N_16838,N_15508,N_14349);
nor U16839 (N_16839,N_14014,N_15639);
and U16840 (N_16840,N_15970,N_14507);
nor U16841 (N_16841,N_14381,N_14037);
or U16842 (N_16842,N_14877,N_15230);
or U16843 (N_16843,N_14259,N_14523);
xor U16844 (N_16844,N_15476,N_15564);
and U16845 (N_16845,N_14099,N_14701);
nand U16846 (N_16846,N_14644,N_14836);
or U16847 (N_16847,N_14580,N_15550);
nand U16848 (N_16848,N_15618,N_14436);
xor U16849 (N_16849,N_14289,N_15133);
xnor U16850 (N_16850,N_14283,N_15727);
or U16851 (N_16851,N_14971,N_15093);
nand U16852 (N_16852,N_14314,N_15539);
xnor U16853 (N_16853,N_15726,N_14127);
xnor U16854 (N_16854,N_15604,N_15426);
nand U16855 (N_16855,N_15631,N_15507);
and U16856 (N_16856,N_14069,N_15459);
nand U16857 (N_16857,N_14237,N_15641);
and U16858 (N_16858,N_15904,N_15040);
nor U16859 (N_16859,N_15223,N_15559);
or U16860 (N_16860,N_14572,N_15428);
and U16861 (N_16861,N_15434,N_14937);
and U16862 (N_16862,N_15271,N_15369);
nand U16863 (N_16863,N_14947,N_14721);
xnor U16864 (N_16864,N_14615,N_14468);
xnor U16865 (N_16865,N_15802,N_14899);
or U16866 (N_16866,N_15118,N_15194);
and U16867 (N_16867,N_14209,N_15504);
nand U16868 (N_16868,N_14365,N_14003);
nor U16869 (N_16869,N_15409,N_15598);
xor U16870 (N_16870,N_14344,N_15636);
nand U16871 (N_16871,N_14777,N_14194);
nor U16872 (N_16872,N_15724,N_14808);
xor U16873 (N_16873,N_15333,N_14668);
nor U16874 (N_16874,N_14648,N_14631);
nand U16875 (N_16875,N_15759,N_15854);
or U16876 (N_16876,N_14007,N_15609);
xor U16877 (N_16877,N_14064,N_15518);
nand U16878 (N_16878,N_15345,N_14960);
and U16879 (N_16879,N_14490,N_15283);
nor U16880 (N_16880,N_15810,N_14792);
xnor U16881 (N_16881,N_15899,N_14921);
or U16882 (N_16882,N_15896,N_14032);
nand U16883 (N_16883,N_15739,N_15033);
nand U16884 (N_16884,N_15692,N_15236);
xor U16885 (N_16885,N_14223,N_14389);
and U16886 (N_16886,N_14945,N_14275);
and U16887 (N_16887,N_15819,N_15908);
nor U16888 (N_16888,N_14372,N_15108);
and U16889 (N_16889,N_14666,N_15331);
nor U16890 (N_16890,N_14375,N_14555);
nor U16891 (N_16891,N_15302,N_15668);
or U16892 (N_16892,N_15534,N_15029);
nor U16893 (N_16893,N_15821,N_15852);
or U16894 (N_16894,N_14688,N_14049);
xor U16895 (N_16895,N_14563,N_14426);
and U16896 (N_16896,N_14607,N_14866);
and U16897 (N_16897,N_15494,N_14459);
xnor U16898 (N_16898,N_15444,N_15807);
or U16899 (N_16899,N_15957,N_14477);
xnor U16900 (N_16900,N_14139,N_15777);
nand U16901 (N_16901,N_14353,N_15487);
xor U16902 (N_16902,N_15431,N_15373);
and U16903 (N_16903,N_15449,N_15616);
nand U16904 (N_16904,N_15526,N_15467);
and U16905 (N_16905,N_14397,N_15190);
and U16906 (N_16906,N_15307,N_14029);
and U16907 (N_16907,N_15619,N_15881);
xor U16908 (N_16908,N_14602,N_15800);
xor U16909 (N_16909,N_14183,N_15388);
nor U16910 (N_16910,N_15880,N_15406);
nand U16911 (N_16911,N_14638,N_15788);
xor U16912 (N_16912,N_15455,N_14867);
nor U16913 (N_16913,N_14943,N_15977);
xor U16914 (N_16914,N_14129,N_14513);
xor U16915 (N_16915,N_14878,N_15323);
nor U16916 (N_16916,N_15273,N_14452);
xnor U16917 (N_16917,N_14425,N_15294);
xor U16918 (N_16918,N_15181,N_15146);
xor U16919 (N_16919,N_14737,N_15961);
xnor U16920 (N_16920,N_14804,N_15382);
nor U16921 (N_16921,N_15831,N_14343);
xnor U16922 (N_16922,N_15573,N_14144);
nor U16923 (N_16923,N_14610,N_15375);
xor U16924 (N_16924,N_15419,N_15846);
nand U16925 (N_16925,N_15546,N_15538);
and U16926 (N_16926,N_15414,N_14266);
nor U16927 (N_16927,N_14954,N_15022);
nor U16928 (N_16928,N_15617,N_15105);
nand U16929 (N_16929,N_15792,N_15308);
nand U16930 (N_16930,N_14022,N_15189);
or U16931 (N_16931,N_15432,N_14858);
or U16932 (N_16932,N_14743,N_14695);
and U16933 (N_16933,N_15234,N_14269);
and U16934 (N_16934,N_15103,N_15394);
and U16935 (N_16935,N_14824,N_14162);
or U16936 (N_16936,N_15143,N_14835);
xor U16937 (N_16937,N_14154,N_15702);
nor U16938 (N_16938,N_15120,N_14364);
xnor U16939 (N_16939,N_14320,N_15027);
xnor U16940 (N_16940,N_14105,N_15489);
nor U16941 (N_16941,N_15710,N_14895);
xor U16942 (N_16942,N_15884,N_14126);
or U16943 (N_16943,N_14406,N_15685);
or U16944 (N_16944,N_15091,N_15697);
nor U16945 (N_16945,N_14010,N_15046);
and U16946 (N_16946,N_14338,N_14462);
and U16947 (N_16947,N_15932,N_14578);
xnor U16948 (N_16948,N_14228,N_15804);
nand U16949 (N_16949,N_14823,N_14886);
nand U16950 (N_16950,N_15280,N_14352);
xnor U16951 (N_16951,N_15799,N_14706);
and U16952 (N_16952,N_15865,N_14717);
nor U16953 (N_16953,N_15019,N_14355);
or U16954 (N_16954,N_15232,N_15420);
and U16955 (N_16955,N_15100,N_15193);
xor U16956 (N_16956,N_15553,N_14434);
and U16957 (N_16957,N_15640,N_15411);
and U16958 (N_16958,N_14539,N_14143);
nand U16959 (N_16959,N_15124,N_14270);
or U16960 (N_16960,N_14519,N_15625);
nor U16961 (N_16961,N_14705,N_15644);
nand U16962 (N_16962,N_14486,N_14282);
xnor U16963 (N_16963,N_15638,N_15111);
nand U16964 (N_16964,N_15329,N_14913);
nand U16965 (N_16965,N_15982,N_15628);
and U16966 (N_16966,N_14439,N_14335);
nor U16967 (N_16967,N_14128,N_14855);
xor U16968 (N_16968,N_15442,N_15667);
nand U16969 (N_16969,N_14745,N_15691);
and U16970 (N_16970,N_15405,N_14145);
nand U16971 (N_16971,N_15292,N_14370);
nor U16972 (N_16972,N_14626,N_15389);
xor U16973 (N_16973,N_14530,N_14492);
nor U16974 (N_16974,N_15448,N_14980);
nor U16975 (N_16975,N_15087,N_14598);
xnor U16976 (N_16976,N_14089,N_15447);
and U16977 (N_16977,N_15999,N_15773);
xor U16978 (N_16978,N_14974,N_14584);
xnor U16979 (N_16979,N_15185,N_14939);
or U16980 (N_16980,N_15495,N_14017);
xnor U16981 (N_16981,N_15979,N_15688);
xor U16982 (N_16982,N_15501,N_14072);
nand U16983 (N_16983,N_14192,N_15689);
and U16984 (N_16984,N_15785,N_14656);
nor U16985 (N_16985,N_14900,N_15552);
xor U16986 (N_16986,N_15150,N_14753);
nor U16987 (N_16987,N_15813,N_15008);
xor U16988 (N_16988,N_14885,N_14390);
or U16989 (N_16989,N_14333,N_14577);
nand U16990 (N_16990,N_15719,N_15717);
or U16991 (N_16991,N_14337,N_14950);
or U16992 (N_16992,N_15094,N_15721);
xor U16993 (N_16993,N_14203,N_14132);
nand U16994 (N_16994,N_15213,N_14747);
or U16995 (N_16995,N_14063,N_15740);
or U16996 (N_16996,N_14673,N_15620);
and U16997 (N_16997,N_15700,N_14113);
nor U16998 (N_16998,N_14796,N_15264);
or U16999 (N_16999,N_15220,N_15445);
nor U17000 (N_17000,N_14596,N_15435);
and U17001 (N_17001,N_14351,N_15254);
xnor U17002 (N_17002,N_14845,N_14240);
and U17003 (N_17003,N_15719,N_15567);
nand U17004 (N_17004,N_15844,N_15350);
nor U17005 (N_17005,N_14486,N_14928);
nand U17006 (N_17006,N_14036,N_14440);
or U17007 (N_17007,N_15131,N_15068);
xnor U17008 (N_17008,N_15607,N_14765);
and U17009 (N_17009,N_14068,N_14996);
nor U17010 (N_17010,N_14184,N_14633);
nand U17011 (N_17011,N_14894,N_15323);
nor U17012 (N_17012,N_15546,N_15778);
or U17013 (N_17013,N_14895,N_15735);
and U17014 (N_17014,N_14989,N_15250);
nor U17015 (N_17015,N_15073,N_15753);
or U17016 (N_17016,N_14622,N_15529);
nor U17017 (N_17017,N_14446,N_15490);
and U17018 (N_17018,N_15339,N_14072);
nor U17019 (N_17019,N_15639,N_15120);
nand U17020 (N_17020,N_15746,N_14107);
nor U17021 (N_17021,N_14453,N_15821);
nand U17022 (N_17022,N_14439,N_14052);
and U17023 (N_17023,N_15927,N_14538);
nand U17024 (N_17024,N_15376,N_15919);
nand U17025 (N_17025,N_15647,N_14167);
and U17026 (N_17026,N_15660,N_15990);
or U17027 (N_17027,N_15421,N_15813);
or U17028 (N_17028,N_15809,N_14410);
or U17029 (N_17029,N_14240,N_15278);
nor U17030 (N_17030,N_14532,N_14870);
nand U17031 (N_17031,N_14276,N_14382);
nor U17032 (N_17032,N_15958,N_14460);
xor U17033 (N_17033,N_14631,N_14863);
nand U17034 (N_17034,N_15613,N_15427);
xor U17035 (N_17035,N_14789,N_14108);
or U17036 (N_17036,N_14297,N_15256);
nor U17037 (N_17037,N_15630,N_14564);
xor U17038 (N_17038,N_14579,N_15282);
or U17039 (N_17039,N_15722,N_14450);
xnor U17040 (N_17040,N_14402,N_14955);
nand U17041 (N_17041,N_14785,N_15634);
xnor U17042 (N_17042,N_15987,N_15490);
or U17043 (N_17043,N_14589,N_14193);
nand U17044 (N_17044,N_14673,N_15305);
nand U17045 (N_17045,N_15777,N_15619);
or U17046 (N_17046,N_14530,N_14655);
nand U17047 (N_17047,N_14609,N_15542);
nor U17048 (N_17048,N_15193,N_14537);
xnor U17049 (N_17049,N_15243,N_15117);
nor U17050 (N_17050,N_14218,N_15156);
xor U17051 (N_17051,N_14948,N_15780);
or U17052 (N_17052,N_15969,N_15202);
and U17053 (N_17053,N_15083,N_15829);
and U17054 (N_17054,N_15496,N_14369);
xor U17055 (N_17055,N_14962,N_15053);
nand U17056 (N_17056,N_15183,N_15164);
xor U17057 (N_17057,N_15624,N_14033);
and U17058 (N_17058,N_14592,N_15714);
nor U17059 (N_17059,N_14010,N_14479);
or U17060 (N_17060,N_15389,N_14180);
or U17061 (N_17061,N_15534,N_15175);
xor U17062 (N_17062,N_14398,N_15807);
nand U17063 (N_17063,N_15067,N_15319);
nor U17064 (N_17064,N_14137,N_15031);
or U17065 (N_17065,N_14524,N_14977);
nor U17066 (N_17066,N_15807,N_14417);
nor U17067 (N_17067,N_15329,N_14960);
nand U17068 (N_17068,N_14330,N_15067);
or U17069 (N_17069,N_15349,N_15976);
or U17070 (N_17070,N_14891,N_14834);
nand U17071 (N_17071,N_14596,N_15221);
nand U17072 (N_17072,N_14284,N_14889);
or U17073 (N_17073,N_15905,N_14263);
nor U17074 (N_17074,N_15468,N_15176);
or U17075 (N_17075,N_15843,N_15210);
and U17076 (N_17076,N_14257,N_15612);
or U17077 (N_17077,N_15514,N_15735);
xor U17078 (N_17078,N_15645,N_15871);
nand U17079 (N_17079,N_15689,N_15971);
and U17080 (N_17080,N_15937,N_15447);
xor U17081 (N_17081,N_14408,N_14329);
xnor U17082 (N_17082,N_15974,N_15004);
nand U17083 (N_17083,N_14922,N_15034);
nor U17084 (N_17084,N_15131,N_14991);
or U17085 (N_17085,N_14935,N_15401);
nor U17086 (N_17086,N_15236,N_14137);
nor U17087 (N_17087,N_14784,N_15470);
and U17088 (N_17088,N_14609,N_14665);
and U17089 (N_17089,N_14170,N_15403);
nor U17090 (N_17090,N_15930,N_14731);
nor U17091 (N_17091,N_15219,N_14071);
xor U17092 (N_17092,N_14952,N_14528);
nor U17093 (N_17093,N_14689,N_15498);
nor U17094 (N_17094,N_14134,N_14950);
or U17095 (N_17095,N_14077,N_15832);
nand U17096 (N_17096,N_15803,N_15249);
nor U17097 (N_17097,N_14905,N_14777);
nand U17098 (N_17098,N_14471,N_15702);
or U17099 (N_17099,N_14012,N_15919);
xnor U17100 (N_17100,N_14642,N_15273);
nor U17101 (N_17101,N_14429,N_14058);
nor U17102 (N_17102,N_14786,N_14087);
xnor U17103 (N_17103,N_14386,N_14795);
nor U17104 (N_17104,N_15754,N_14780);
and U17105 (N_17105,N_15165,N_15911);
nor U17106 (N_17106,N_15475,N_14695);
nor U17107 (N_17107,N_14137,N_15193);
nand U17108 (N_17108,N_14305,N_15682);
nor U17109 (N_17109,N_15878,N_14398);
or U17110 (N_17110,N_15932,N_14038);
nand U17111 (N_17111,N_14811,N_14571);
nor U17112 (N_17112,N_14455,N_15010);
nand U17113 (N_17113,N_14535,N_14337);
nor U17114 (N_17114,N_15967,N_15583);
xnor U17115 (N_17115,N_14446,N_14611);
or U17116 (N_17116,N_15289,N_14816);
or U17117 (N_17117,N_15202,N_14352);
nor U17118 (N_17118,N_14728,N_15045);
nor U17119 (N_17119,N_15071,N_14886);
xnor U17120 (N_17120,N_14880,N_15561);
xnor U17121 (N_17121,N_15381,N_15293);
xnor U17122 (N_17122,N_15272,N_15593);
nor U17123 (N_17123,N_14844,N_14860);
or U17124 (N_17124,N_14219,N_15567);
and U17125 (N_17125,N_14999,N_15643);
and U17126 (N_17126,N_14234,N_14321);
nand U17127 (N_17127,N_14589,N_14410);
xor U17128 (N_17128,N_14389,N_14876);
nand U17129 (N_17129,N_15210,N_15610);
nor U17130 (N_17130,N_14216,N_14152);
xnor U17131 (N_17131,N_14613,N_15538);
nand U17132 (N_17132,N_15914,N_14637);
nor U17133 (N_17133,N_14305,N_14853);
or U17134 (N_17134,N_14036,N_15823);
and U17135 (N_17135,N_15047,N_15732);
xnor U17136 (N_17136,N_15462,N_14041);
nand U17137 (N_17137,N_14475,N_14685);
nand U17138 (N_17138,N_14621,N_14459);
or U17139 (N_17139,N_15842,N_14001);
nor U17140 (N_17140,N_14059,N_14602);
xnor U17141 (N_17141,N_15405,N_15599);
or U17142 (N_17142,N_15373,N_14508);
xnor U17143 (N_17143,N_14044,N_15443);
or U17144 (N_17144,N_15283,N_14720);
nor U17145 (N_17145,N_15311,N_15052);
and U17146 (N_17146,N_14530,N_15401);
or U17147 (N_17147,N_14234,N_14600);
xnor U17148 (N_17148,N_14731,N_15434);
nand U17149 (N_17149,N_15104,N_15364);
nand U17150 (N_17150,N_14385,N_14709);
nand U17151 (N_17151,N_14356,N_14185);
xor U17152 (N_17152,N_14002,N_14256);
nor U17153 (N_17153,N_14152,N_15401);
nand U17154 (N_17154,N_14470,N_15446);
xor U17155 (N_17155,N_14004,N_15420);
and U17156 (N_17156,N_15916,N_15354);
or U17157 (N_17157,N_14527,N_14779);
or U17158 (N_17158,N_14348,N_15995);
xor U17159 (N_17159,N_15529,N_15989);
or U17160 (N_17160,N_15165,N_14609);
or U17161 (N_17161,N_15444,N_15507);
or U17162 (N_17162,N_14167,N_14391);
or U17163 (N_17163,N_15057,N_14327);
and U17164 (N_17164,N_14018,N_14594);
xnor U17165 (N_17165,N_14804,N_14909);
xor U17166 (N_17166,N_15351,N_15859);
nor U17167 (N_17167,N_15572,N_15475);
or U17168 (N_17168,N_15092,N_15412);
nand U17169 (N_17169,N_14201,N_14724);
and U17170 (N_17170,N_15936,N_14068);
xor U17171 (N_17171,N_15787,N_15410);
xor U17172 (N_17172,N_15745,N_14929);
and U17173 (N_17173,N_14823,N_14030);
xor U17174 (N_17174,N_15657,N_15355);
xnor U17175 (N_17175,N_14757,N_14284);
xnor U17176 (N_17176,N_14557,N_14796);
and U17177 (N_17177,N_14613,N_14913);
or U17178 (N_17178,N_14761,N_14859);
and U17179 (N_17179,N_14227,N_15591);
nor U17180 (N_17180,N_15868,N_14158);
or U17181 (N_17181,N_15265,N_15728);
nor U17182 (N_17182,N_15649,N_14690);
and U17183 (N_17183,N_15853,N_14665);
or U17184 (N_17184,N_14493,N_15826);
or U17185 (N_17185,N_14329,N_14272);
or U17186 (N_17186,N_15394,N_15892);
xnor U17187 (N_17187,N_14906,N_14039);
xor U17188 (N_17188,N_15347,N_15384);
xor U17189 (N_17189,N_15937,N_14336);
nand U17190 (N_17190,N_15126,N_14861);
xnor U17191 (N_17191,N_14994,N_14526);
and U17192 (N_17192,N_14409,N_15350);
and U17193 (N_17193,N_14144,N_14793);
nand U17194 (N_17194,N_15720,N_14098);
and U17195 (N_17195,N_14201,N_14589);
or U17196 (N_17196,N_15659,N_14551);
nor U17197 (N_17197,N_14251,N_15367);
nand U17198 (N_17198,N_15521,N_15465);
and U17199 (N_17199,N_15136,N_14187);
and U17200 (N_17200,N_15551,N_15330);
or U17201 (N_17201,N_15364,N_14694);
nand U17202 (N_17202,N_15365,N_14762);
and U17203 (N_17203,N_14502,N_14084);
nand U17204 (N_17204,N_14621,N_14842);
nand U17205 (N_17205,N_15619,N_14434);
or U17206 (N_17206,N_14286,N_14037);
and U17207 (N_17207,N_14938,N_15071);
or U17208 (N_17208,N_14290,N_15835);
nand U17209 (N_17209,N_14164,N_15470);
nor U17210 (N_17210,N_15219,N_14254);
nor U17211 (N_17211,N_15353,N_15822);
nand U17212 (N_17212,N_14992,N_14003);
or U17213 (N_17213,N_15488,N_14807);
xor U17214 (N_17214,N_14242,N_14359);
nand U17215 (N_17215,N_14720,N_15231);
xnor U17216 (N_17216,N_15697,N_15480);
and U17217 (N_17217,N_14722,N_15321);
nand U17218 (N_17218,N_14206,N_15573);
nand U17219 (N_17219,N_14629,N_14779);
and U17220 (N_17220,N_14057,N_15775);
and U17221 (N_17221,N_15226,N_14017);
nand U17222 (N_17222,N_14174,N_14835);
nor U17223 (N_17223,N_14689,N_15582);
nand U17224 (N_17224,N_15263,N_15562);
xor U17225 (N_17225,N_14270,N_14618);
or U17226 (N_17226,N_15798,N_15194);
nor U17227 (N_17227,N_14986,N_15789);
nand U17228 (N_17228,N_14744,N_15594);
or U17229 (N_17229,N_15946,N_14857);
or U17230 (N_17230,N_14463,N_14541);
xor U17231 (N_17231,N_15752,N_15595);
and U17232 (N_17232,N_14481,N_14676);
xnor U17233 (N_17233,N_15083,N_15407);
and U17234 (N_17234,N_14199,N_14206);
or U17235 (N_17235,N_14543,N_15371);
or U17236 (N_17236,N_14137,N_15944);
nor U17237 (N_17237,N_14994,N_15730);
nand U17238 (N_17238,N_14082,N_15146);
xnor U17239 (N_17239,N_15399,N_14037);
or U17240 (N_17240,N_14964,N_14907);
xnor U17241 (N_17241,N_15202,N_14867);
nand U17242 (N_17242,N_15599,N_15372);
xnor U17243 (N_17243,N_15192,N_15054);
nor U17244 (N_17244,N_15159,N_15446);
nand U17245 (N_17245,N_14601,N_15020);
xor U17246 (N_17246,N_15368,N_15134);
xnor U17247 (N_17247,N_15445,N_14712);
nand U17248 (N_17248,N_15164,N_15613);
nor U17249 (N_17249,N_14294,N_15668);
xnor U17250 (N_17250,N_15403,N_15474);
xor U17251 (N_17251,N_15526,N_15964);
nor U17252 (N_17252,N_15288,N_15599);
nand U17253 (N_17253,N_15321,N_15475);
or U17254 (N_17254,N_14261,N_15619);
or U17255 (N_17255,N_15568,N_15428);
and U17256 (N_17256,N_14785,N_14577);
nor U17257 (N_17257,N_15930,N_15273);
nand U17258 (N_17258,N_15958,N_14768);
or U17259 (N_17259,N_14996,N_15206);
and U17260 (N_17260,N_15491,N_14316);
or U17261 (N_17261,N_14379,N_15114);
and U17262 (N_17262,N_15074,N_14620);
nand U17263 (N_17263,N_15367,N_15279);
xnor U17264 (N_17264,N_15086,N_14220);
nor U17265 (N_17265,N_14429,N_15987);
xnor U17266 (N_17266,N_15151,N_15612);
and U17267 (N_17267,N_15026,N_14650);
or U17268 (N_17268,N_15674,N_14937);
or U17269 (N_17269,N_15776,N_15224);
and U17270 (N_17270,N_15671,N_14053);
nand U17271 (N_17271,N_15702,N_14257);
or U17272 (N_17272,N_14556,N_14973);
nor U17273 (N_17273,N_15814,N_14613);
and U17274 (N_17274,N_14589,N_14928);
xnor U17275 (N_17275,N_14463,N_14445);
xnor U17276 (N_17276,N_14905,N_14602);
nand U17277 (N_17277,N_14895,N_14473);
nand U17278 (N_17278,N_14387,N_15116);
nand U17279 (N_17279,N_15603,N_15392);
xor U17280 (N_17280,N_14327,N_15450);
xnor U17281 (N_17281,N_15293,N_14021);
xnor U17282 (N_17282,N_14989,N_14120);
xnor U17283 (N_17283,N_14613,N_14837);
and U17284 (N_17284,N_15909,N_15064);
or U17285 (N_17285,N_14979,N_15476);
nand U17286 (N_17286,N_15134,N_15274);
xnor U17287 (N_17287,N_15608,N_15450);
nor U17288 (N_17288,N_15176,N_14504);
or U17289 (N_17289,N_15675,N_15546);
or U17290 (N_17290,N_14099,N_14356);
and U17291 (N_17291,N_14394,N_15919);
or U17292 (N_17292,N_14311,N_14969);
and U17293 (N_17293,N_15608,N_14447);
xnor U17294 (N_17294,N_15390,N_14438);
or U17295 (N_17295,N_14222,N_14865);
nand U17296 (N_17296,N_14898,N_14998);
xor U17297 (N_17297,N_14609,N_15321);
nor U17298 (N_17298,N_14463,N_15173);
xor U17299 (N_17299,N_14836,N_14260);
xor U17300 (N_17300,N_15548,N_14933);
nand U17301 (N_17301,N_15651,N_14060);
and U17302 (N_17302,N_15644,N_14767);
xor U17303 (N_17303,N_15168,N_14223);
or U17304 (N_17304,N_15100,N_14874);
or U17305 (N_17305,N_15223,N_14463);
or U17306 (N_17306,N_15498,N_14435);
nor U17307 (N_17307,N_14826,N_14882);
and U17308 (N_17308,N_14731,N_15594);
nor U17309 (N_17309,N_15765,N_14835);
nor U17310 (N_17310,N_15405,N_15607);
or U17311 (N_17311,N_14563,N_15867);
nand U17312 (N_17312,N_15806,N_15316);
xor U17313 (N_17313,N_14106,N_15371);
nor U17314 (N_17314,N_15172,N_14630);
nand U17315 (N_17315,N_15829,N_14176);
nor U17316 (N_17316,N_15271,N_15628);
and U17317 (N_17317,N_14910,N_15268);
nor U17318 (N_17318,N_14400,N_14477);
nor U17319 (N_17319,N_14223,N_15802);
nand U17320 (N_17320,N_15520,N_15804);
nor U17321 (N_17321,N_15918,N_14762);
nand U17322 (N_17322,N_14080,N_15000);
nor U17323 (N_17323,N_15442,N_14705);
nor U17324 (N_17324,N_15389,N_14461);
or U17325 (N_17325,N_14945,N_14460);
nor U17326 (N_17326,N_15318,N_14711);
and U17327 (N_17327,N_14239,N_15291);
and U17328 (N_17328,N_14149,N_14873);
and U17329 (N_17329,N_14329,N_15388);
nor U17330 (N_17330,N_15243,N_15461);
nor U17331 (N_17331,N_15466,N_14346);
and U17332 (N_17332,N_15001,N_14822);
nand U17333 (N_17333,N_14338,N_14645);
and U17334 (N_17334,N_14769,N_14917);
nand U17335 (N_17335,N_14485,N_15626);
or U17336 (N_17336,N_14722,N_14161);
or U17337 (N_17337,N_14097,N_15526);
nand U17338 (N_17338,N_14357,N_15363);
and U17339 (N_17339,N_14886,N_14694);
nand U17340 (N_17340,N_14280,N_14746);
xor U17341 (N_17341,N_15319,N_15498);
nand U17342 (N_17342,N_15910,N_15231);
and U17343 (N_17343,N_15207,N_14514);
or U17344 (N_17344,N_14432,N_14301);
nor U17345 (N_17345,N_15808,N_15829);
nand U17346 (N_17346,N_15418,N_14635);
nand U17347 (N_17347,N_15501,N_15027);
nor U17348 (N_17348,N_15593,N_15874);
and U17349 (N_17349,N_15677,N_15931);
and U17350 (N_17350,N_15224,N_14186);
nand U17351 (N_17351,N_14113,N_14762);
nand U17352 (N_17352,N_15759,N_15575);
or U17353 (N_17353,N_15536,N_15002);
xnor U17354 (N_17354,N_14983,N_14488);
xor U17355 (N_17355,N_15852,N_14782);
nand U17356 (N_17356,N_15820,N_15036);
nor U17357 (N_17357,N_14089,N_14947);
nand U17358 (N_17358,N_15867,N_15937);
nor U17359 (N_17359,N_14253,N_15172);
xor U17360 (N_17360,N_15815,N_15552);
xnor U17361 (N_17361,N_14836,N_15827);
nor U17362 (N_17362,N_14806,N_15065);
or U17363 (N_17363,N_14840,N_15413);
or U17364 (N_17364,N_14453,N_14825);
nand U17365 (N_17365,N_14252,N_14987);
and U17366 (N_17366,N_14473,N_15202);
nand U17367 (N_17367,N_14803,N_14049);
or U17368 (N_17368,N_14778,N_15002);
nand U17369 (N_17369,N_15130,N_15368);
or U17370 (N_17370,N_15601,N_15948);
nand U17371 (N_17371,N_14319,N_14361);
xnor U17372 (N_17372,N_15526,N_14509);
xor U17373 (N_17373,N_14881,N_14921);
nor U17374 (N_17374,N_15623,N_15224);
nand U17375 (N_17375,N_15376,N_15624);
and U17376 (N_17376,N_14183,N_14176);
or U17377 (N_17377,N_14596,N_14178);
nand U17378 (N_17378,N_15952,N_15412);
xnor U17379 (N_17379,N_15733,N_15582);
or U17380 (N_17380,N_15829,N_15178);
xnor U17381 (N_17381,N_15584,N_15129);
or U17382 (N_17382,N_14068,N_15871);
or U17383 (N_17383,N_15417,N_14202);
xor U17384 (N_17384,N_14874,N_15436);
xor U17385 (N_17385,N_15253,N_14336);
or U17386 (N_17386,N_15272,N_15694);
nand U17387 (N_17387,N_14443,N_14405);
or U17388 (N_17388,N_15743,N_14567);
and U17389 (N_17389,N_14664,N_15105);
nor U17390 (N_17390,N_15717,N_14556);
or U17391 (N_17391,N_15930,N_14702);
nor U17392 (N_17392,N_15304,N_14098);
or U17393 (N_17393,N_15467,N_14667);
nand U17394 (N_17394,N_14666,N_14018);
or U17395 (N_17395,N_15742,N_14896);
or U17396 (N_17396,N_14653,N_15317);
xor U17397 (N_17397,N_15350,N_14851);
or U17398 (N_17398,N_14019,N_14847);
nor U17399 (N_17399,N_15328,N_15196);
or U17400 (N_17400,N_15225,N_15474);
nand U17401 (N_17401,N_14675,N_14859);
xnor U17402 (N_17402,N_14274,N_14317);
and U17403 (N_17403,N_14196,N_15211);
nand U17404 (N_17404,N_15480,N_14420);
or U17405 (N_17405,N_15689,N_15188);
nand U17406 (N_17406,N_14126,N_14012);
nor U17407 (N_17407,N_15642,N_15214);
xor U17408 (N_17408,N_15711,N_15198);
nor U17409 (N_17409,N_15640,N_14004);
nand U17410 (N_17410,N_14331,N_14943);
nand U17411 (N_17411,N_15303,N_15861);
xnor U17412 (N_17412,N_15867,N_15152);
nand U17413 (N_17413,N_15402,N_15855);
nor U17414 (N_17414,N_15746,N_15594);
or U17415 (N_17415,N_15869,N_14978);
or U17416 (N_17416,N_15795,N_14812);
or U17417 (N_17417,N_15707,N_15108);
nor U17418 (N_17418,N_15980,N_14151);
nor U17419 (N_17419,N_14149,N_14902);
or U17420 (N_17420,N_14451,N_15456);
or U17421 (N_17421,N_15633,N_15611);
or U17422 (N_17422,N_14798,N_15455);
xor U17423 (N_17423,N_14249,N_15251);
nor U17424 (N_17424,N_14321,N_14967);
and U17425 (N_17425,N_15962,N_14803);
nor U17426 (N_17426,N_14526,N_15061);
and U17427 (N_17427,N_14217,N_14003);
xor U17428 (N_17428,N_15430,N_14619);
or U17429 (N_17429,N_15427,N_14090);
nor U17430 (N_17430,N_15803,N_14792);
or U17431 (N_17431,N_15597,N_15487);
and U17432 (N_17432,N_14569,N_15904);
xnor U17433 (N_17433,N_14034,N_15196);
xnor U17434 (N_17434,N_14576,N_15566);
or U17435 (N_17435,N_15516,N_14046);
or U17436 (N_17436,N_14232,N_14355);
nor U17437 (N_17437,N_14352,N_14557);
or U17438 (N_17438,N_14262,N_14371);
nand U17439 (N_17439,N_14120,N_15639);
and U17440 (N_17440,N_14728,N_15053);
nor U17441 (N_17441,N_14643,N_14115);
and U17442 (N_17442,N_15362,N_14955);
nand U17443 (N_17443,N_14093,N_14949);
nand U17444 (N_17444,N_14565,N_14101);
nand U17445 (N_17445,N_14994,N_14848);
and U17446 (N_17446,N_14864,N_15483);
xor U17447 (N_17447,N_14960,N_14426);
nand U17448 (N_17448,N_15745,N_14857);
nor U17449 (N_17449,N_15336,N_14816);
nand U17450 (N_17450,N_14459,N_15647);
xnor U17451 (N_17451,N_14148,N_14260);
xor U17452 (N_17452,N_14828,N_15668);
and U17453 (N_17453,N_14652,N_15829);
xnor U17454 (N_17454,N_15136,N_14024);
nand U17455 (N_17455,N_14666,N_15901);
xnor U17456 (N_17456,N_15683,N_15955);
nand U17457 (N_17457,N_14988,N_15269);
or U17458 (N_17458,N_14787,N_15708);
xnor U17459 (N_17459,N_15998,N_14151);
or U17460 (N_17460,N_14674,N_15447);
and U17461 (N_17461,N_15101,N_15501);
or U17462 (N_17462,N_14663,N_15900);
xnor U17463 (N_17463,N_14160,N_15544);
nand U17464 (N_17464,N_14799,N_14995);
nand U17465 (N_17465,N_15529,N_15651);
xnor U17466 (N_17466,N_14518,N_14727);
or U17467 (N_17467,N_14662,N_15336);
nor U17468 (N_17468,N_14453,N_14717);
xnor U17469 (N_17469,N_14517,N_15888);
and U17470 (N_17470,N_15756,N_14394);
or U17471 (N_17471,N_14537,N_14091);
or U17472 (N_17472,N_15922,N_15106);
and U17473 (N_17473,N_14737,N_15052);
nand U17474 (N_17474,N_15899,N_14548);
and U17475 (N_17475,N_15371,N_15982);
and U17476 (N_17476,N_14391,N_15081);
nand U17477 (N_17477,N_15104,N_14441);
xor U17478 (N_17478,N_15606,N_15466);
or U17479 (N_17479,N_14200,N_15738);
and U17480 (N_17480,N_15283,N_14786);
xor U17481 (N_17481,N_14533,N_15646);
and U17482 (N_17482,N_14055,N_14628);
nand U17483 (N_17483,N_14260,N_15395);
nand U17484 (N_17484,N_15973,N_15011);
or U17485 (N_17485,N_14238,N_14901);
nand U17486 (N_17486,N_14662,N_15167);
and U17487 (N_17487,N_15598,N_14712);
nand U17488 (N_17488,N_15868,N_15248);
and U17489 (N_17489,N_15895,N_14015);
nor U17490 (N_17490,N_14252,N_14321);
and U17491 (N_17491,N_14238,N_15097);
xnor U17492 (N_17492,N_15528,N_14633);
nor U17493 (N_17493,N_14095,N_15947);
or U17494 (N_17494,N_14625,N_14614);
and U17495 (N_17495,N_15385,N_14911);
nand U17496 (N_17496,N_14061,N_14875);
nand U17497 (N_17497,N_14913,N_14895);
or U17498 (N_17498,N_14619,N_14004);
and U17499 (N_17499,N_15318,N_15825);
xor U17500 (N_17500,N_15260,N_15867);
and U17501 (N_17501,N_14254,N_14267);
and U17502 (N_17502,N_15947,N_15932);
and U17503 (N_17503,N_14062,N_15005);
and U17504 (N_17504,N_14086,N_15518);
xor U17505 (N_17505,N_14118,N_14071);
nor U17506 (N_17506,N_14442,N_14650);
and U17507 (N_17507,N_14247,N_15865);
and U17508 (N_17508,N_15559,N_14294);
or U17509 (N_17509,N_15374,N_15022);
nor U17510 (N_17510,N_15403,N_15113);
nand U17511 (N_17511,N_15938,N_15597);
xor U17512 (N_17512,N_15298,N_15643);
nor U17513 (N_17513,N_15672,N_15478);
xnor U17514 (N_17514,N_14065,N_15078);
nand U17515 (N_17515,N_15685,N_15652);
xor U17516 (N_17516,N_14556,N_15885);
nor U17517 (N_17517,N_15097,N_15032);
and U17518 (N_17518,N_15201,N_15273);
and U17519 (N_17519,N_15948,N_14461);
or U17520 (N_17520,N_14686,N_14714);
nand U17521 (N_17521,N_15649,N_14567);
xor U17522 (N_17522,N_14174,N_15551);
or U17523 (N_17523,N_15651,N_14821);
xnor U17524 (N_17524,N_14865,N_14946);
xor U17525 (N_17525,N_14206,N_15216);
xor U17526 (N_17526,N_14606,N_14950);
nor U17527 (N_17527,N_14229,N_15529);
or U17528 (N_17528,N_14219,N_15584);
and U17529 (N_17529,N_14603,N_15618);
and U17530 (N_17530,N_15543,N_14198);
nor U17531 (N_17531,N_15047,N_15050);
and U17532 (N_17532,N_14151,N_15568);
xor U17533 (N_17533,N_15057,N_15355);
or U17534 (N_17534,N_14162,N_15876);
nand U17535 (N_17535,N_14276,N_14645);
or U17536 (N_17536,N_14986,N_15500);
nor U17537 (N_17537,N_15740,N_15550);
xor U17538 (N_17538,N_14988,N_14207);
and U17539 (N_17539,N_15260,N_15835);
nor U17540 (N_17540,N_14203,N_14943);
and U17541 (N_17541,N_14318,N_14643);
and U17542 (N_17542,N_15050,N_15243);
and U17543 (N_17543,N_15802,N_15758);
nor U17544 (N_17544,N_15920,N_14187);
nor U17545 (N_17545,N_15274,N_15548);
and U17546 (N_17546,N_14788,N_15062);
xor U17547 (N_17547,N_14278,N_15024);
xor U17548 (N_17548,N_14498,N_14119);
or U17549 (N_17549,N_14174,N_15267);
and U17550 (N_17550,N_14663,N_15654);
nor U17551 (N_17551,N_15025,N_15206);
nand U17552 (N_17552,N_15708,N_14837);
nand U17553 (N_17553,N_14592,N_15904);
or U17554 (N_17554,N_15720,N_14453);
xor U17555 (N_17555,N_14417,N_15764);
nand U17556 (N_17556,N_14863,N_14801);
and U17557 (N_17557,N_15701,N_15266);
or U17558 (N_17558,N_14419,N_15657);
nor U17559 (N_17559,N_14414,N_15597);
nor U17560 (N_17560,N_14582,N_14458);
nor U17561 (N_17561,N_14558,N_15191);
and U17562 (N_17562,N_15188,N_14258);
and U17563 (N_17563,N_15847,N_15579);
nor U17564 (N_17564,N_14175,N_15187);
nor U17565 (N_17565,N_15214,N_14081);
and U17566 (N_17566,N_15741,N_14270);
nor U17567 (N_17567,N_15587,N_14521);
nand U17568 (N_17568,N_14449,N_14541);
or U17569 (N_17569,N_15979,N_14244);
xnor U17570 (N_17570,N_14996,N_14189);
nand U17571 (N_17571,N_15528,N_15674);
nand U17572 (N_17572,N_14521,N_14360);
or U17573 (N_17573,N_15739,N_14114);
or U17574 (N_17574,N_15331,N_15728);
nor U17575 (N_17575,N_14016,N_14484);
nand U17576 (N_17576,N_15904,N_14119);
xor U17577 (N_17577,N_14913,N_14460);
nand U17578 (N_17578,N_15101,N_14982);
nand U17579 (N_17579,N_15886,N_14367);
or U17580 (N_17580,N_14364,N_14333);
nand U17581 (N_17581,N_14033,N_15558);
xor U17582 (N_17582,N_15462,N_15252);
nor U17583 (N_17583,N_14186,N_15096);
or U17584 (N_17584,N_14415,N_15960);
nand U17585 (N_17585,N_14488,N_14151);
nor U17586 (N_17586,N_15026,N_15773);
nor U17587 (N_17587,N_14510,N_15265);
nor U17588 (N_17588,N_14631,N_15112);
or U17589 (N_17589,N_14124,N_14203);
nor U17590 (N_17590,N_14868,N_15874);
nand U17591 (N_17591,N_15366,N_15309);
nand U17592 (N_17592,N_14354,N_15154);
and U17593 (N_17593,N_14705,N_15566);
or U17594 (N_17594,N_15816,N_15336);
nand U17595 (N_17595,N_15932,N_14147);
and U17596 (N_17596,N_15543,N_14069);
and U17597 (N_17597,N_15248,N_14800);
nor U17598 (N_17598,N_15774,N_14933);
nand U17599 (N_17599,N_15635,N_14325);
and U17600 (N_17600,N_14737,N_14798);
or U17601 (N_17601,N_14115,N_14666);
nand U17602 (N_17602,N_15152,N_14587);
and U17603 (N_17603,N_15804,N_14144);
and U17604 (N_17604,N_14213,N_15723);
or U17605 (N_17605,N_15386,N_15144);
nand U17606 (N_17606,N_14995,N_14982);
or U17607 (N_17607,N_15407,N_14609);
nor U17608 (N_17608,N_15918,N_14058);
xnor U17609 (N_17609,N_15790,N_14729);
xor U17610 (N_17610,N_15860,N_14362);
or U17611 (N_17611,N_15810,N_15001);
and U17612 (N_17612,N_15049,N_15719);
xnor U17613 (N_17613,N_14625,N_14709);
or U17614 (N_17614,N_14097,N_14857);
and U17615 (N_17615,N_14662,N_14926);
nor U17616 (N_17616,N_14901,N_15617);
xnor U17617 (N_17617,N_15237,N_14185);
and U17618 (N_17618,N_14430,N_14070);
xnor U17619 (N_17619,N_14973,N_14338);
xnor U17620 (N_17620,N_15471,N_15581);
and U17621 (N_17621,N_15325,N_15946);
nand U17622 (N_17622,N_14690,N_15883);
xnor U17623 (N_17623,N_15968,N_15352);
nand U17624 (N_17624,N_15476,N_15840);
xnor U17625 (N_17625,N_14489,N_15256);
nand U17626 (N_17626,N_15822,N_15857);
xor U17627 (N_17627,N_14211,N_15388);
nor U17628 (N_17628,N_14116,N_15464);
nor U17629 (N_17629,N_14893,N_14131);
nand U17630 (N_17630,N_14456,N_14539);
nor U17631 (N_17631,N_15331,N_14436);
and U17632 (N_17632,N_14478,N_15702);
nor U17633 (N_17633,N_15854,N_15495);
xor U17634 (N_17634,N_14900,N_14333);
nand U17635 (N_17635,N_14563,N_14286);
and U17636 (N_17636,N_14725,N_15623);
or U17637 (N_17637,N_14629,N_15617);
nand U17638 (N_17638,N_15962,N_14392);
nor U17639 (N_17639,N_14634,N_15632);
xnor U17640 (N_17640,N_15191,N_14798);
and U17641 (N_17641,N_15834,N_15509);
nor U17642 (N_17642,N_15723,N_15444);
nor U17643 (N_17643,N_14683,N_15168);
nor U17644 (N_17644,N_14666,N_14317);
nand U17645 (N_17645,N_15259,N_14148);
nand U17646 (N_17646,N_15008,N_14259);
or U17647 (N_17647,N_15332,N_14311);
xnor U17648 (N_17648,N_15509,N_15844);
nand U17649 (N_17649,N_14728,N_15920);
or U17650 (N_17650,N_14344,N_15293);
nand U17651 (N_17651,N_15369,N_15387);
or U17652 (N_17652,N_15091,N_14989);
nor U17653 (N_17653,N_15513,N_14223);
and U17654 (N_17654,N_14838,N_14674);
xnor U17655 (N_17655,N_14278,N_14863);
or U17656 (N_17656,N_14110,N_14762);
or U17657 (N_17657,N_14014,N_14922);
nor U17658 (N_17658,N_15016,N_14500);
nand U17659 (N_17659,N_15990,N_15480);
and U17660 (N_17660,N_14157,N_14395);
nor U17661 (N_17661,N_14579,N_15540);
xnor U17662 (N_17662,N_14548,N_14924);
nor U17663 (N_17663,N_14529,N_15354);
and U17664 (N_17664,N_15613,N_14577);
nand U17665 (N_17665,N_14133,N_14858);
nand U17666 (N_17666,N_15124,N_14872);
nor U17667 (N_17667,N_14308,N_15947);
or U17668 (N_17668,N_15342,N_15662);
nor U17669 (N_17669,N_14407,N_15071);
nor U17670 (N_17670,N_15383,N_15256);
nand U17671 (N_17671,N_15843,N_14714);
and U17672 (N_17672,N_15930,N_15858);
nor U17673 (N_17673,N_15808,N_14855);
nor U17674 (N_17674,N_15848,N_15627);
nor U17675 (N_17675,N_15292,N_14944);
xnor U17676 (N_17676,N_14964,N_15753);
nor U17677 (N_17677,N_15309,N_14636);
nor U17678 (N_17678,N_15715,N_15511);
nor U17679 (N_17679,N_15505,N_14310);
nand U17680 (N_17680,N_15771,N_15343);
and U17681 (N_17681,N_14157,N_15886);
nor U17682 (N_17682,N_15428,N_14074);
nand U17683 (N_17683,N_15835,N_15308);
and U17684 (N_17684,N_15608,N_14745);
xnor U17685 (N_17685,N_15860,N_14074);
xnor U17686 (N_17686,N_15267,N_14133);
nor U17687 (N_17687,N_14082,N_14749);
or U17688 (N_17688,N_14050,N_14814);
or U17689 (N_17689,N_15723,N_15882);
xnor U17690 (N_17690,N_14714,N_14043);
and U17691 (N_17691,N_14909,N_15901);
nor U17692 (N_17692,N_15343,N_15022);
nor U17693 (N_17693,N_15813,N_14994);
nand U17694 (N_17694,N_14433,N_14619);
and U17695 (N_17695,N_14344,N_14474);
and U17696 (N_17696,N_15391,N_15001);
xnor U17697 (N_17697,N_14811,N_14660);
and U17698 (N_17698,N_15624,N_14066);
nand U17699 (N_17699,N_14219,N_15147);
xnor U17700 (N_17700,N_14974,N_14587);
xnor U17701 (N_17701,N_14501,N_14085);
nand U17702 (N_17702,N_15652,N_14654);
and U17703 (N_17703,N_15642,N_14943);
xnor U17704 (N_17704,N_15063,N_15701);
xor U17705 (N_17705,N_15533,N_14987);
or U17706 (N_17706,N_14755,N_14489);
and U17707 (N_17707,N_15190,N_14172);
or U17708 (N_17708,N_15167,N_15390);
nor U17709 (N_17709,N_14234,N_15928);
nand U17710 (N_17710,N_15419,N_15359);
nor U17711 (N_17711,N_14231,N_15336);
xor U17712 (N_17712,N_14898,N_14879);
nor U17713 (N_17713,N_15795,N_15571);
and U17714 (N_17714,N_14699,N_14097);
or U17715 (N_17715,N_14329,N_15258);
or U17716 (N_17716,N_14584,N_15327);
or U17717 (N_17717,N_15859,N_15079);
nor U17718 (N_17718,N_15822,N_14389);
and U17719 (N_17719,N_15710,N_14868);
nand U17720 (N_17720,N_15961,N_15538);
nand U17721 (N_17721,N_14396,N_14591);
nor U17722 (N_17722,N_14659,N_14220);
or U17723 (N_17723,N_15314,N_14217);
nor U17724 (N_17724,N_14825,N_15174);
nor U17725 (N_17725,N_14304,N_14712);
xor U17726 (N_17726,N_14871,N_14231);
nand U17727 (N_17727,N_15647,N_15562);
nor U17728 (N_17728,N_15065,N_14680);
or U17729 (N_17729,N_14335,N_14629);
nand U17730 (N_17730,N_14716,N_14492);
or U17731 (N_17731,N_14730,N_14064);
nand U17732 (N_17732,N_15158,N_15181);
nand U17733 (N_17733,N_14175,N_14599);
or U17734 (N_17734,N_15361,N_14864);
and U17735 (N_17735,N_15444,N_15141);
or U17736 (N_17736,N_15521,N_15907);
nor U17737 (N_17737,N_15372,N_14091);
nor U17738 (N_17738,N_14068,N_14414);
nor U17739 (N_17739,N_15624,N_15175);
and U17740 (N_17740,N_15093,N_15698);
and U17741 (N_17741,N_14492,N_14574);
xor U17742 (N_17742,N_15139,N_14075);
nand U17743 (N_17743,N_15634,N_15973);
nor U17744 (N_17744,N_15970,N_15897);
nand U17745 (N_17745,N_15915,N_14525);
and U17746 (N_17746,N_14112,N_14948);
nand U17747 (N_17747,N_15940,N_14498);
nor U17748 (N_17748,N_14941,N_15558);
or U17749 (N_17749,N_15659,N_15943);
nand U17750 (N_17750,N_14280,N_15111);
nor U17751 (N_17751,N_14123,N_15943);
xnor U17752 (N_17752,N_15080,N_14259);
and U17753 (N_17753,N_15656,N_15418);
xor U17754 (N_17754,N_15552,N_15535);
nor U17755 (N_17755,N_15116,N_14108);
nor U17756 (N_17756,N_14641,N_14017);
nor U17757 (N_17757,N_15365,N_14123);
nand U17758 (N_17758,N_15435,N_15445);
or U17759 (N_17759,N_15656,N_14778);
or U17760 (N_17760,N_15189,N_15461);
or U17761 (N_17761,N_14675,N_15587);
nor U17762 (N_17762,N_15619,N_14836);
xnor U17763 (N_17763,N_15922,N_15407);
xnor U17764 (N_17764,N_14107,N_14649);
and U17765 (N_17765,N_15251,N_15146);
and U17766 (N_17766,N_15867,N_14577);
nand U17767 (N_17767,N_15044,N_15774);
nor U17768 (N_17768,N_14852,N_15155);
nand U17769 (N_17769,N_15960,N_15594);
xnor U17770 (N_17770,N_14277,N_14706);
nor U17771 (N_17771,N_15285,N_14035);
nor U17772 (N_17772,N_15645,N_14187);
xor U17773 (N_17773,N_14239,N_15359);
xnor U17774 (N_17774,N_15135,N_15774);
xnor U17775 (N_17775,N_14067,N_14765);
nand U17776 (N_17776,N_15262,N_15880);
nor U17777 (N_17777,N_14758,N_14061);
or U17778 (N_17778,N_14751,N_15686);
or U17779 (N_17779,N_15998,N_15467);
xor U17780 (N_17780,N_14338,N_14558);
nand U17781 (N_17781,N_15273,N_15066);
xor U17782 (N_17782,N_14663,N_14604);
xor U17783 (N_17783,N_15703,N_14549);
xor U17784 (N_17784,N_14192,N_15876);
nand U17785 (N_17785,N_15321,N_15579);
nand U17786 (N_17786,N_15992,N_14437);
nor U17787 (N_17787,N_14976,N_14004);
and U17788 (N_17788,N_15279,N_14627);
and U17789 (N_17789,N_15748,N_15797);
nand U17790 (N_17790,N_15458,N_15061);
or U17791 (N_17791,N_15889,N_14308);
xnor U17792 (N_17792,N_14090,N_14752);
xor U17793 (N_17793,N_15219,N_15799);
and U17794 (N_17794,N_14879,N_14341);
and U17795 (N_17795,N_14785,N_15571);
nand U17796 (N_17796,N_14108,N_15195);
or U17797 (N_17797,N_15495,N_15361);
xor U17798 (N_17798,N_14884,N_15084);
xor U17799 (N_17799,N_14015,N_15743);
xnor U17800 (N_17800,N_15231,N_14979);
nor U17801 (N_17801,N_15307,N_14422);
and U17802 (N_17802,N_14966,N_14058);
and U17803 (N_17803,N_15363,N_14455);
and U17804 (N_17804,N_14950,N_14510);
or U17805 (N_17805,N_15930,N_14979);
nand U17806 (N_17806,N_14727,N_14045);
nor U17807 (N_17807,N_15776,N_14565);
xor U17808 (N_17808,N_15673,N_15354);
nand U17809 (N_17809,N_15360,N_15039);
xnor U17810 (N_17810,N_14635,N_15159);
xor U17811 (N_17811,N_14231,N_15668);
xor U17812 (N_17812,N_14382,N_15864);
and U17813 (N_17813,N_14420,N_15689);
nand U17814 (N_17814,N_14194,N_14734);
and U17815 (N_17815,N_15994,N_15051);
xor U17816 (N_17816,N_15164,N_14333);
and U17817 (N_17817,N_14629,N_15035);
xnor U17818 (N_17818,N_15089,N_14381);
nor U17819 (N_17819,N_15386,N_14239);
or U17820 (N_17820,N_14276,N_14178);
or U17821 (N_17821,N_14921,N_15110);
nand U17822 (N_17822,N_14267,N_15229);
or U17823 (N_17823,N_15212,N_15112);
or U17824 (N_17824,N_15149,N_15040);
nand U17825 (N_17825,N_15023,N_15660);
xnor U17826 (N_17826,N_15868,N_15826);
xnor U17827 (N_17827,N_14627,N_14351);
and U17828 (N_17828,N_15133,N_15568);
nand U17829 (N_17829,N_15325,N_14920);
or U17830 (N_17830,N_14300,N_14127);
nor U17831 (N_17831,N_15851,N_15710);
nand U17832 (N_17832,N_14797,N_15693);
xor U17833 (N_17833,N_15513,N_14611);
nand U17834 (N_17834,N_14219,N_15248);
xor U17835 (N_17835,N_14178,N_15177);
nor U17836 (N_17836,N_14982,N_15894);
xnor U17837 (N_17837,N_14984,N_14215);
xor U17838 (N_17838,N_14167,N_15564);
and U17839 (N_17839,N_14867,N_15731);
nor U17840 (N_17840,N_14874,N_14916);
or U17841 (N_17841,N_15176,N_14035);
or U17842 (N_17842,N_15330,N_14381);
nand U17843 (N_17843,N_14619,N_14136);
xor U17844 (N_17844,N_14742,N_15356);
and U17845 (N_17845,N_15485,N_15923);
xnor U17846 (N_17846,N_14577,N_15931);
and U17847 (N_17847,N_14657,N_15817);
nor U17848 (N_17848,N_15551,N_15106);
or U17849 (N_17849,N_14482,N_14326);
xnor U17850 (N_17850,N_15138,N_15478);
and U17851 (N_17851,N_14434,N_15749);
and U17852 (N_17852,N_15361,N_15077);
nand U17853 (N_17853,N_15683,N_15950);
and U17854 (N_17854,N_15052,N_15758);
nand U17855 (N_17855,N_14310,N_15522);
xnor U17856 (N_17856,N_14785,N_15263);
xnor U17857 (N_17857,N_14971,N_15781);
and U17858 (N_17858,N_15164,N_15241);
nor U17859 (N_17859,N_14795,N_14150);
or U17860 (N_17860,N_14610,N_15464);
nor U17861 (N_17861,N_14993,N_14808);
or U17862 (N_17862,N_14816,N_15139);
or U17863 (N_17863,N_15425,N_15198);
nand U17864 (N_17864,N_15108,N_15336);
or U17865 (N_17865,N_14177,N_15481);
or U17866 (N_17866,N_15154,N_15905);
nand U17867 (N_17867,N_15865,N_14499);
and U17868 (N_17868,N_15190,N_15159);
or U17869 (N_17869,N_14606,N_14444);
or U17870 (N_17870,N_15476,N_14297);
nand U17871 (N_17871,N_15952,N_14544);
nand U17872 (N_17872,N_15989,N_15685);
nor U17873 (N_17873,N_14212,N_15453);
xnor U17874 (N_17874,N_14171,N_14701);
nand U17875 (N_17875,N_14889,N_14619);
xnor U17876 (N_17876,N_14539,N_14851);
or U17877 (N_17877,N_14234,N_15162);
nand U17878 (N_17878,N_14247,N_14461);
and U17879 (N_17879,N_15088,N_15495);
nand U17880 (N_17880,N_14955,N_14206);
nor U17881 (N_17881,N_14378,N_15347);
and U17882 (N_17882,N_14869,N_15294);
xor U17883 (N_17883,N_15586,N_14669);
nand U17884 (N_17884,N_14644,N_15239);
or U17885 (N_17885,N_15591,N_15389);
nand U17886 (N_17886,N_15445,N_14967);
or U17887 (N_17887,N_14699,N_15288);
nor U17888 (N_17888,N_14684,N_14668);
nand U17889 (N_17889,N_15225,N_15430);
and U17890 (N_17890,N_15464,N_14767);
xnor U17891 (N_17891,N_15782,N_15739);
and U17892 (N_17892,N_15171,N_14509);
and U17893 (N_17893,N_15587,N_14394);
or U17894 (N_17894,N_15049,N_14916);
and U17895 (N_17895,N_15362,N_14554);
nor U17896 (N_17896,N_14406,N_15496);
nor U17897 (N_17897,N_14905,N_15848);
or U17898 (N_17898,N_15167,N_15351);
nand U17899 (N_17899,N_14670,N_14783);
and U17900 (N_17900,N_14873,N_14472);
nor U17901 (N_17901,N_15728,N_14085);
or U17902 (N_17902,N_15241,N_14689);
or U17903 (N_17903,N_15954,N_15030);
xor U17904 (N_17904,N_14236,N_14799);
and U17905 (N_17905,N_14263,N_15370);
nor U17906 (N_17906,N_15760,N_15299);
xor U17907 (N_17907,N_14200,N_15827);
or U17908 (N_17908,N_14782,N_14837);
xor U17909 (N_17909,N_15561,N_15556);
nor U17910 (N_17910,N_14991,N_14307);
or U17911 (N_17911,N_15131,N_15014);
xor U17912 (N_17912,N_14798,N_15334);
nand U17913 (N_17913,N_15505,N_15161);
or U17914 (N_17914,N_14878,N_14244);
xor U17915 (N_17915,N_14332,N_14267);
and U17916 (N_17916,N_15256,N_14110);
or U17917 (N_17917,N_15947,N_14215);
xnor U17918 (N_17918,N_14034,N_14393);
nor U17919 (N_17919,N_14279,N_15692);
nor U17920 (N_17920,N_15156,N_15538);
and U17921 (N_17921,N_14514,N_14034);
and U17922 (N_17922,N_15121,N_14172);
nand U17923 (N_17923,N_15762,N_14329);
and U17924 (N_17924,N_14810,N_14431);
xnor U17925 (N_17925,N_14502,N_14139);
or U17926 (N_17926,N_15168,N_15519);
nand U17927 (N_17927,N_14998,N_15575);
xnor U17928 (N_17928,N_14528,N_14648);
xnor U17929 (N_17929,N_14561,N_15860);
nor U17930 (N_17930,N_15028,N_15909);
or U17931 (N_17931,N_15034,N_15133);
xor U17932 (N_17932,N_14287,N_14733);
nor U17933 (N_17933,N_15137,N_15488);
nand U17934 (N_17934,N_15380,N_14020);
xnor U17935 (N_17935,N_15502,N_15206);
nor U17936 (N_17936,N_14495,N_15812);
nand U17937 (N_17937,N_14598,N_15371);
xnor U17938 (N_17938,N_14948,N_15478);
or U17939 (N_17939,N_14236,N_15151);
or U17940 (N_17940,N_15292,N_14965);
nor U17941 (N_17941,N_15742,N_14386);
or U17942 (N_17942,N_15664,N_15184);
nor U17943 (N_17943,N_14342,N_15564);
nor U17944 (N_17944,N_14345,N_14663);
or U17945 (N_17945,N_14790,N_14971);
nand U17946 (N_17946,N_15124,N_15035);
and U17947 (N_17947,N_15780,N_14265);
or U17948 (N_17948,N_15144,N_14966);
xnor U17949 (N_17949,N_14583,N_14858);
and U17950 (N_17950,N_14541,N_15235);
and U17951 (N_17951,N_14010,N_15730);
or U17952 (N_17952,N_14021,N_14148);
or U17953 (N_17953,N_14105,N_14856);
nor U17954 (N_17954,N_15952,N_14363);
nor U17955 (N_17955,N_15270,N_14062);
or U17956 (N_17956,N_14540,N_14470);
xnor U17957 (N_17957,N_14104,N_15717);
or U17958 (N_17958,N_14389,N_15086);
xnor U17959 (N_17959,N_15159,N_14436);
xor U17960 (N_17960,N_14152,N_14078);
xnor U17961 (N_17961,N_14547,N_15658);
xor U17962 (N_17962,N_15710,N_15148);
xnor U17963 (N_17963,N_15822,N_15600);
xnor U17964 (N_17964,N_14343,N_15512);
xor U17965 (N_17965,N_14471,N_14322);
nand U17966 (N_17966,N_15861,N_15052);
nand U17967 (N_17967,N_15590,N_14286);
xnor U17968 (N_17968,N_15902,N_15452);
or U17969 (N_17969,N_15712,N_15132);
nand U17970 (N_17970,N_14239,N_14989);
and U17971 (N_17971,N_15503,N_14472);
xor U17972 (N_17972,N_14579,N_15732);
nand U17973 (N_17973,N_14373,N_14001);
nand U17974 (N_17974,N_15166,N_14750);
nand U17975 (N_17975,N_15381,N_15954);
or U17976 (N_17976,N_15092,N_14608);
xnor U17977 (N_17977,N_14824,N_14949);
xnor U17978 (N_17978,N_15645,N_15429);
or U17979 (N_17979,N_15480,N_15598);
or U17980 (N_17980,N_14886,N_14593);
nor U17981 (N_17981,N_14238,N_15219);
or U17982 (N_17982,N_14187,N_14528);
and U17983 (N_17983,N_14790,N_14521);
or U17984 (N_17984,N_15753,N_14847);
nand U17985 (N_17985,N_15245,N_14901);
or U17986 (N_17986,N_15836,N_15251);
nand U17987 (N_17987,N_15693,N_14056);
and U17988 (N_17988,N_15565,N_15331);
or U17989 (N_17989,N_14954,N_15654);
xor U17990 (N_17990,N_14372,N_15227);
and U17991 (N_17991,N_15478,N_14730);
xnor U17992 (N_17992,N_14298,N_14054);
nand U17993 (N_17993,N_14890,N_14150);
nand U17994 (N_17994,N_15277,N_14053);
or U17995 (N_17995,N_15594,N_15071);
and U17996 (N_17996,N_15624,N_15102);
nor U17997 (N_17997,N_15023,N_14487);
and U17998 (N_17998,N_15624,N_15353);
xor U17999 (N_17999,N_14808,N_15205);
nand U18000 (N_18000,N_16454,N_17320);
or U18001 (N_18001,N_16094,N_16451);
nor U18002 (N_18002,N_16936,N_17657);
nor U18003 (N_18003,N_17656,N_16206);
and U18004 (N_18004,N_17350,N_17321);
xnor U18005 (N_18005,N_16077,N_17278);
or U18006 (N_18006,N_17708,N_17345);
nand U18007 (N_18007,N_17033,N_16397);
or U18008 (N_18008,N_17375,N_16236);
xor U18009 (N_18009,N_17461,N_17249);
and U18010 (N_18010,N_17550,N_16685);
nand U18011 (N_18011,N_16811,N_17798);
xor U18012 (N_18012,N_17797,N_16944);
nand U18013 (N_18013,N_16486,N_16548);
nor U18014 (N_18014,N_17495,N_17447);
or U18015 (N_18015,N_17792,N_17599);
and U18016 (N_18016,N_16752,N_16097);
nand U18017 (N_18017,N_16862,N_16037);
nand U18018 (N_18018,N_17970,N_17431);
or U18019 (N_18019,N_16614,N_16759);
and U18020 (N_18020,N_16322,N_16426);
or U18021 (N_18021,N_16370,N_17411);
and U18022 (N_18022,N_17817,N_16544);
or U18023 (N_18023,N_16181,N_17303);
and U18024 (N_18024,N_17854,N_17511);
nor U18025 (N_18025,N_16976,N_16150);
nor U18026 (N_18026,N_16931,N_16139);
xnor U18027 (N_18027,N_17665,N_17347);
and U18028 (N_18028,N_16915,N_17148);
or U18029 (N_18029,N_16355,N_16443);
xor U18030 (N_18030,N_16934,N_17801);
nor U18031 (N_18031,N_17416,N_16377);
and U18032 (N_18032,N_16007,N_17327);
and U18033 (N_18033,N_16636,N_17283);
nor U18034 (N_18034,N_16885,N_17450);
nand U18035 (N_18035,N_17097,N_16802);
and U18036 (N_18036,N_16172,N_16637);
or U18037 (N_18037,N_16026,N_16252);
xor U18038 (N_18038,N_16897,N_17740);
nand U18039 (N_18039,N_17109,N_17610);
and U18040 (N_18040,N_17858,N_17679);
and U18041 (N_18041,N_16683,N_17795);
xnor U18042 (N_18042,N_17257,N_17160);
xnor U18043 (N_18043,N_16147,N_16837);
nor U18044 (N_18044,N_16553,N_17986);
nand U18045 (N_18045,N_16424,N_16599);
xor U18046 (N_18046,N_16148,N_17157);
and U18047 (N_18047,N_17448,N_16063);
nand U18048 (N_18048,N_16713,N_16048);
and U18049 (N_18049,N_16358,N_17339);
nand U18050 (N_18050,N_16843,N_17769);
and U18051 (N_18051,N_17232,N_16638);
or U18052 (N_18052,N_16894,N_16615);
xnor U18053 (N_18053,N_17721,N_17166);
or U18054 (N_18054,N_17393,N_17732);
xor U18055 (N_18055,N_17156,N_16572);
xnor U18056 (N_18056,N_16722,N_17235);
nand U18057 (N_18057,N_17548,N_17059);
and U18058 (N_18058,N_17524,N_17057);
or U18059 (N_18059,N_16753,N_16761);
xor U18060 (N_18060,N_16854,N_16482);
and U18061 (N_18061,N_17950,N_17880);
and U18062 (N_18062,N_17529,N_16167);
or U18063 (N_18063,N_16285,N_17521);
nor U18064 (N_18064,N_17125,N_17510);
and U18065 (N_18065,N_17515,N_16547);
nand U18066 (N_18066,N_16901,N_17605);
nand U18067 (N_18067,N_17389,N_17228);
and U18068 (N_18068,N_16144,N_17454);
nand U18069 (N_18069,N_17381,N_16992);
or U18070 (N_18070,N_16237,N_16771);
and U18071 (N_18071,N_16012,N_16794);
nor U18072 (N_18072,N_17026,N_16699);
or U18073 (N_18073,N_17990,N_17781);
nand U18074 (N_18074,N_16178,N_17434);
nor U18075 (N_18075,N_17113,N_16475);
nand U18076 (N_18076,N_17103,N_17341);
xor U18077 (N_18077,N_16689,N_16573);
nand U18078 (N_18078,N_16983,N_17756);
nor U18079 (N_18079,N_17982,N_17618);
or U18080 (N_18080,N_17883,N_16087);
nand U18081 (N_18081,N_16402,N_17875);
xor U18082 (N_18082,N_16390,N_16495);
or U18083 (N_18083,N_16008,N_16398);
or U18084 (N_18084,N_16265,N_17742);
xor U18085 (N_18085,N_16845,N_17567);
nor U18086 (N_18086,N_17172,N_17242);
nor U18087 (N_18087,N_16306,N_17907);
xor U18088 (N_18088,N_17972,N_16861);
nor U18089 (N_18089,N_17607,N_17908);
or U18090 (N_18090,N_17074,N_17799);
xnor U18091 (N_18091,N_17582,N_16380);
and U18092 (N_18092,N_16601,N_17004);
and U18093 (N_18093,N_16881,N_16066);
xnor U18094 (N_18094,N_17192,N_16217);
or U18095 (N_18095,N_16744,N_17762);
xor U18096 (N_18096,N_17114,N_17892);
nand U18097 (N_18097,N_16082,N_16311);
and U18098 (N_18098,N_17323,N_17037);
nor U18099 (N_18099,N_17244,N_17170);
and U18100 (N_18100,N_17851,N_16775);
nand U18101 (N_18101,N_17855,N_16704);
nor U18102 (N_18102,N_17147,N_16290);
nand U18103 (N_18103,N_16395,N_17396);
xnor U18104 (N_18104,N_16904,N_17559);
nor U18105 (N_18105,N_17934,N_16746);
nand U18106 (N_18106,N_16857,N_17534);
nand U18107 (N_18107,N_17506,N_17671);
and U18108 (N_18108,N_16820,N_17500);
nand U18109 (N_18109,N_16100,N_16198);
and U18110 (N_18110,N_17081,N_17841);
xnor U18111 (N_18111,N_16690,N_16307);
xor U18112 (N_18112,N_16581,N_17887);
or U18113 (N_18113,N_17348,N_16255);
and U18114 (N_18114,N_17065,N_17615);
nand U18115 (N_18115,N_17919,N_16118);
nand U18116 (N_18116,N_17398,N_16504);
xor U18117 (N_18117,N_17922,N_16001);
nor U18118 (N_18118,N_16863,N_17318);
and U18119 (N_18119,N_17196,N_16988);
xor U18120 (N_18120,N_17989,N_17491);
and U18121 (N_18121,N_16231,N_16348);
xnor U18122 (N_18122,N_17988,N_16764);
nand U18123 (N_18123,N_16321,N_16978);
xor U18124 (N_18124,N_17728,N_16437);
nor U18125 (N_18125,N_16565,N_17358);
nor U18126 (N_18126,N_16496,N_16392);
or U18127 (N_18127,N_16296,N_16902);
and U18128 (N_18128,N_17508,N_16073);
nor U18129 (N_18129,N_17248,N_16590);
and U18130 (N_18130,N_16661,N_17083);
nor U18131 (N_18131,N_17701,N_16175);
and U18132 (N_18132,N_17182,N_17473);
nor U18133 (N_18133,N_16790,N_16328);
nor U18134 (N_18134,N_17068,N_16877);
or U18135 (N_18135,N_16295,N_16731);
nand U18136 (N_18136,N_17173,N_16153);
and U18137 (N_18137,N_16982,N_16014);
or U18138 (N_18138,N_16228,N_17996);
xnor U18139 (N_18139,N_17675,N_16987);
xor U18140 (N_18140,N_17146,N_17682);
nor U18141 (N_18141,N_17788,N_16256);
or U18142 (N_18142,N_16546,N_17713);
or U18143 (N_18143,N_17269,N_17539);
nand U18144 (N_18144,N_16340,N_17304);
or U18145 (N_18145,N_16706,N_16937);
xor U18146 (N_18146,N_16163,N_16418);
nor U18147 (N_18147,N_16972,N_17775);
or U18148 (N_18148,N_16798,N_17296);
xnor U18149 (N_18149,N_17370,N_17415);
xnor U18150 (N_18150,N_16550,N_17429);
xnor U18151 (N_18151,N_17203,N_17642);
xor U18152 (N_18152,N_16003,N_16438);
xor U18153 (N_18153,N_17426,N_16728);
and U18154 (N_18154,N_17834,N_17308);
nand U18155 (N_18155,N_17107,N_16613);
and U18156 (N_18156,N_16433,N_17064);
or U18157 (N_18157,N_17070,N_17509);
and U18158 (N_18158,N_16520,N_16542);
nand U18159 (N_18159,N_16420,N_17806);
xnor U18160 (N_18160,N_17388,N_16021);
nor U18161 (N_18161,N_17749,N_17018);
nand U18162 (N_18162,N_17357,N_16477);
xnor U18163 (N_18163,N_16436,N_16059);
nand U18164 (N_18164,N_17791,N_16154);
xor U18165 (N_18165,N_17717,N_17758);
nor U18166 (N_18166,N_16580,N_16018);
nor U18167 (N_18167,N_17027,N_17889);
nor U18168 (N_18168,N_17284,N_16448);
nand U18169 (N_18169,N_16801,N_16812);
and U18170 (N_18170,N_17460,N_17365);
nor U18171 (N_18171,N_16170,N_16226);
or U18172 (N_18172,N_16169,N_17777);
and U18173 (N_18173,N_17367,N_16566);
xor U18174 (N_18174,N_16326,N_16359);
nand U18175 (N_18175,N_16445,N_16386);
or U18176 (N_18176,N_17119,N_16994);
or U18177 (N_18177,N_16408,N_17234);
xnor U18178 (N_18178,N_17600,N_17171);
and U18179 (N_18179,N_16027,N_17666);
nor U18180 (N_18180,N_16016,N_16062);
nor U18181 (N_18181,N_16493,N_17092);
nor U18182 (N_18182,N_16558,N_16914);
nor U18183 (N_18183,N_16109,N_16955);
or U18184 (N_18184,N_17385,N_17514);
and U18185 (N_18185,N_17723,N_17267);
or U18186 (N_18186,N_17343,N_16755);
xor U18187 (N_18187,N_17634,N_16041);
nor U18188 (N_18188,N_17476,N_16896);
or U18189 (N_18189,N_16528,N_17086);
nor U18190 (N_18190,N_16492,N_16336);
xor U18191 (N_18191,N_17127,N_16498);
nand U18192 (N_18192,N_16289,N_16060);
nand U18193 (N_18193,N_17360,N_16313);
or U18194 (N_18194,N_17702,N_16391);
nand U18195 (N_18195,N_17028,N_17819);
and U18196 (N_18196,N_17319,N_17424);
or U18197 (N_18197,N_16586,N_17977);
and U18198 (N_18198,N_16500,N_16530);
or U18199 (N_18199,N_17313,N_16072);
and U18200 (N_18200,N_17194,N_17122);
nor U18201 (N_18201,N_17457,N_16765);
xnor U18202 (N_18202,N_17686,N_16610);
and U18203 (N_18203,N_16792,N_17100);
or U18204 (N_18204,N_16521,N_17941);
nand U18205 (N_18205,N_16508,N_17289);
nand U18206 (N_18206,N_17088,N_16594);
xnor U18207 (N_18207,N_17538,N_17459);
and U18208 (N_18208,N_17593,N_17374);
and U18209 (N_18209,N_17186,N_16507);
xor U18210 (N_18210,N_16724,N_16218);
or U18211 (N_18211,N_16197,N_17525);
and U18212 (N_18212,N_17900,N_17104);
or U18213 (N_18213,N_16966,N_17685);
and U18214 (N_18214,N_17803,N_17330);
and U18215 (N_18215,N_16549,N_16184);
nor U18216 (N_18216,N_16083,N_17061);
nand U18217 (N_18217,N_17928,N_17785);
nor U18218 (N_18218,N_16560,N_16751);
or U18219 (N_18219,N_17213,N_16382);
xnor U18220 (N_18220,N_17118,N_16770);
and U18221 (N_18221,N_17418,N_16518);
and U18222 (N_18222,N_17102,N_16917);
xnor U18223 (N_18223,N_17093,N_17885);
or U18224 (N_18224,N_16168,N_17551);
nand U18225 (N_18225,N_17958,N_17456);
or U18226 (N_18226,N_16463,N_17250);
or U18227 (N_18227,N_16998,N_16005);
or U18228 (N_18228,N_16385,N_17573);
and U18229 (N_18229,N_16000,N_16241);
and U18230 (N_18230,N_16293,N_16791);
nor U18231 (N_18231,N_17453,N_16563);
xor U18232 (N_18232,N_17383,N_16160);
nand U18233 (N_18233,N_16145,N_16733);
nand U18234 (N_18234,N_17489,N_16024);
and U18235 (N_18235,N_16648,N_17487);
nand U18236 (N_18236,N_16162,N_17309);
nor U18237 (N_18237,N_17580,N_17688);
and U18238 (N_18238,N_16272,N_17240);
nand U18239 (N_18239,N_16114,N_16186);
xnor U18240 (N_18240,N_17942,N_17655);
nand U18241 (N_18241,N_16776,N_16333);
xnor U18242 (N_18242,N_17778,N_16271);
or U18243 (N_18243,N_16047,N_17690);
xnor U18244 (N_18244,N_16611,N_16387);
xnor U18245 (N_18245,N_17449,N_17625);
nand U18246 (N_18246,N_16298,N_16138);
nor U18247 (N_18247,N_16287,N_17921);
and U18248 (N_18248,N_17162,N_16253);
and U18249 (N_18249,N_17918,N_16292);
and U18250 (N_18250,N_17041,N_16585);
or U18251 (N_18251,N_16207,N_16795);
xor U18252 (N_18252,N_16876,N_17901);
or U18253 (N_18253,N_17804,N_16875);
and U18254 (N_18254,N_17532,N_17696);
xnor U18255 (N_18255,N_16803,N_17949);
nor U18256 (N_18256,N_16916,N_16105);
and U18257 (N_18257,N_17207,N_17555);
nor U18258 (N_18258,N_16129,N_16177);
and U18259 (N_18259,N_17528,N_17991);
or U18260 (N_18260,N_17470,N_17340);
and U18261 (N_18261,N_16479,N_16161);
nand U18262 (N_18262,N_17060,N_17006);
xnor U18263 (N_18263,N_16243,N_16229);
nor U18264 (N_18264,N_17346,N_16254);
or U18265 (N_18265,N_16777,N_17624);
xnor U18266 (N_18266,N_17753,N_16692);
and U18267 (N_18267,N_16165,N_17743);
nand U18268 (N_18268,N_16334,N_16095);
or U18269 (N_18269,N_16085,N_17220);
or U18270 (N_18270,N_16069,N_16928);
and U18271 (N_18271,N_17169,N_17019);
nor U18272 (N_18272,N_17905,N_16680);
or U18273 (N_18273,N_16291,N_17926);
xnor U18274 (N_18274,N_16055,N_16659);
xor U18275 (N_18275,N_17979,N_17334);
or U18276 (N_18276,N_17286,N_17992);
and U18277 (N_18277,N_16841,N_16260);
xor U18278 (N_18278,N_17277,N_17463);
nor U18279 (N_18279,N_16444,N_16946);
or U18280 (N_18280,N_17485,N_16757);
nor U18281 (N_18281,N_16848,N_17633);
or U18282 (N_18282,N_17899,N_16906);
xnor U18283 (N_18283,N_17766,N_16804);
or U18284 (N_18284,N_17189,N_17581);
xnor U18285 (N_18285,N_17324,N_17222);
nor U18286 (N_18286,N_16210,N_16609);
nand U18287 (N_18287,N_16891,N_17363);
nor U18288 (N_18288,N_17481,N_17591);
and U18289 (N_18289,N_17042,N_16376);
nor U18290 (N_18290,N_17852,N_16952);
xor U18291 (N_18291,N_17594,N_17468);
and U18292 (N_18292,N_17430,N_17748);
nor U18293 (N_18293,N_16535,N_16247);
xor U18294 (N_18294,N_16511,N_16831);
nand U18295 (N_18295,N_16742,N_17836);
nand U18296 (N_18296,N_16101,N_16384);
nor U18297 (N_18297,N_16506,N_16694);
nand U18298 (N_18298,N_16887,N_16552);
nor U18299 (N_18299,N_17126,N_16597);
xor U18300 (N_18300,N_16985,N_16209);
or U18301 (N_18301,N_17043,N_16591);
nand U18302 (N_18302,N_17054,N_17895);
and U18303 (N_18303,N_17630,N_17015);
nor U18304 (N_18304,N_16403,N_16702);
nand U18305 (N_18305,N_16275,N_17698);
or U18306 (N_18306,N_17295,N_17527);
nand U18307 (N_18307,N_16128,N_17399);
xor U18308 (N_18308,N_17705,N_17362);
or U18309 (N_18309,N_16905,N_17999);
nand U18310 (N_18310,N_17779,N_16641);
or U18311 (N_18311,N_16793,N_16244);
nand U18312 (N_18312,N_16545,N_16747);
xor U18313 (N_18313,N_17985,N_16280);
nor U18314 (N_18314,N_17075,N_17247);
nor U18315 (N_18315,N_17874,N_17782);
nor U18316 (N_18316,N_16634,N_17442);
xnor U18317 (N_18317,N_16478,N_17079);
nand U18318 (N_18318,N_17722,N_17706);
or U18319 (N_18319,N_17839,N_16400);
nor U18320 (N_18320,N_16465,N_17676);
nand U18321 (N_18321,N_17419,N_17137);
and U18322 (N_18322,N_17071,N_16423);
nand U18323 (N_18323,N_16277,N_17379);
nand U18324 (N_18324,N_16068,N_17862);
xor U18325 (N_18325,N_16709,N_17332);
or U18326 (N_18326,N_16577,N_16649);
nand U18327 (N_18327,N_17603,N_17585);
or U18328 (N_18328,N_16413,N_16338);
nand U18329 (N_18329,N_17712,N_16039);
nor U18330 (N_18330,N_17121,N_16886);
or U18331 (N_18331,N_17586,N_17281);
or U18332 (N_18332,N_16137,N_16053);
xor U18333 (N_18333,N_17554,N_17604);
and U18334 (N_18334,N_16717,N_17904);
nor U18335 (N_18335,N_16351,N_17544);
xnor U18336 (N_18336,N_16782,N_16223);
and U18337 (N_18337,N_17427,N_16199);
and U18338 (N_18338,N_17577,N_17478);
xnor U18339 (N_18339,N_17626,N_16374);
xnor U18340 (N_18340,N_17204,N_17711);
nor U18341 (N_18341,N_16971,N_17913);
nand U18342 (N_18342,N_16013,N_17155);
nor U18343 (N_18343,N_17187,N_17823);
nor U18344 (N_18344,N_16632,N_17536);
or U18345 (N_18345,N_16948,N_16625);
nor U18346 (N_18346,N_16335,N_16204);
nor U18347 (N_18347,N_16950,N_16949);
or U18348 (N_18348,N_17410,N_17215);
or U18349 (N_18349,N_17650,N_16570);
nand U18350 (N_18350,N_16503,N_16234);
or U18351 (N_18351,N_16174,N_17261);
nor U18352 (N_18352,N_17774,N_17025);
nor U18353 (N_18353,N_17565,N_16809);
nand U18354 (N_18354,N_16679,N_17499);
or U18355 (N_18355,N_17469,N_16850);
or U18356 (N_18356,N_16045,N_16404);
nand U18357 (N_18357,N_16647,N_17643);
xnor U18358 (N_18358,N_17329,N_16242);
xor U18359 (N_18359,N_17805,N_16286);
nor U18360 (N_18360,N_17387,N_16369);
or U18361 (N_18361,N_17294,N_16682);
and U18362 (N_18362,N_17667,N_16773);
or U18363 (N_18363,N_17896,N_17877);
and U18364 (N_18364,N_16633,N_16120);
xor U18365 (N_18365,N_17246,N_16180);
xor U18366 (N_18366,N_16929,N_16716);
and U18367 (N_18367,N_16650,N_16888);
nor U18368 (N_18368,N_17151,N_16619);
nor U18369 (N_18369,N_16990,N_17929);
xnor U18370 (N_18370,N_16895,N_17631);
or U18371 (N_18371,N_17110,N_17751);
nand U18372 (N_18372,N_17828,N_16079);
or U18373 (N_18373,N_17502,N_17815);
or U18374 (N_18374,N_17455,N_16074);
or U18375 (N_18375,N_17770,N_16409);
or U18376 (N_18376,N_17271,N_17552);
and U18377 (N_18377,N_16718,N_16196);
nand U18378 (N_18378,N_17307,N_16605);
and U18379 (N_18379,N_16785,N_17428);
and U18380 (N_18380,N_16526,N_17869);
or U18381 (N_18381,N_17692,N_16194);
nand U18382 (N_18382,N_16346,N_17870);
nand U18383 (N_18383,N_17953,N_17984);
nor U18384 (N_18384,N_17649,N_17820);
nor U18385 (N_18385,N_17458,N_16266);
nand U18386 (N_18386,N_17252,N_16484);
nand U18387 (N_18387,N_16968,N_16092);
nand U18388 (N_18388,N_17394,N_17161);
or U18389 (N_18389,N_16363,N_16727);
or U18390 (N_18390,N_17617,N_17969);
nor U18391 (N_18391,N_17715,N_17566);
and U18392 (N_18392,N_17446,N_16273);
nor U18393 (N_18393,N_16490,N_16668);
and U18394 (N_18394,N_16999,N_17435);
or U18395 (N_18395,N_17944,N_16980);
nand U18396 (N_18396,N_16766,N_17780);
or U18397 (N_18397,N_17653,N_16628);
nor U18398 (N_18398,N_17568,N_16838);
xor U18399 (N_18399,N_16211,N_16658);
xnor U18400 (N_18400,N_17968,N_16061);
nand U18401 (N_18401,N_17637,N_17111);
or U18402 (N_18402,N_16942,N_16378);
nor U18403 (N_18403,N_16225,N_16856);
xnor U18404 (N_18404,N_17105,N_17466);
xnor U18405 (N_18405,N_17338,N_17031);
nand U18406 (N_18406,N_16667,N_16991);
xor U18407 (N_18407,N_16527,N_16575);
nor U18408 (N_18408,N_16458,N_16921);
and U18409 (N_18409,N_17843,N_17291);
nand U18410 (N_18410,N_16935,N_17231);
xor U18411 (N_18411,N_17592,N_17597);
nand U18412 (N_18412,N_17747,N_16453);
nor U18413 (N_18413,N_17008,N_16918);
or U18414 (N_18414,N_16245,N_16612);
xnor U18415 (N_18415,N_17654,N_16367);
and U18416 (N_18416,N_16310,N_17505);
nand U18417 (N_18417,N_16783,N_17290);
xor U18418 (N_18418,N_16835,N_17245);
and U18419 (N_18419,N_16878,N_17754);
nand U18420 (N_18420,N_17965,N_16467);
nor U18421 (N_18421,N_16739,N_17523);
or U18422 (N_18422,N_16368,N_17786);
xnor U18423 (N_18423,N_16250,N_17522);
nor U18424 (N_18424,N_16556,N_17386);
nor U18425 (N_18425,N_16489,N_17336);
and U18426 (N_18426,N_16582,N_16331);
nand U18427 (N_18427,N_16587,N_17106);
and U18428 (N_18428,N_16332,N_16833);
nor U18429 (N_18429,N_16319,N_17314);
or U18430 (N_18430,N_17098,N_17498);
or U18431 (N_18431,N_16440,N_17335);
nor U18432 (N_18432,N_16561,N_16600);
nand U18433 (N_18433,N_16933,N_17793);
nor U18434 (N_18434,N_16112,N_16539);
or U18435 (N_18435,N_17226,N_17200);
nand U18436 (N_18436,N_16442,N_16462);
nand U18437 (N_18437,N_17443,N_16616);
or U18438 (N_18438,N_17516,N_17050);
nor U18439 (N_18439,N_17402,N_16604);
and U18440 (N_18440,N_16028,N_17178);
xor U18441 (N_18441,N_16571,N_16762);
nor U18442 (N_18442,N_16476,N_17371);
and U18443 (N_18443,N_17645,N_16381);
nand U18444 (N_18444,N_16815,N_17535);
xnor U18445 (N_18445,N_16951,N_17465);
nor U18446 (N_18446,N_16240,N_16674);
xor U18447 (N_18447,N_16911,N_17480);
or U18448 (N_18448,N_16134,N_16188);
or U18449 (N_18449,N_16672,N_17488);
or U18450 (N_18450,N_17438,N_16720);
and U18451 (N_18451,N_16870,N_17142);
and U18452 (N_18452,N_16763,N_16088);
or U18453 (N_18453,N_16883,N_16712);
nand U18454 (N_18454,N_16166,N_17556);
nor U18455 (N_18455,N_16703,N_16309);
xor U18456 (N_18456,N_16093,N_17983);
xor U18457 (N_18457,N_17325,N_17214);
xor U18458 (N_18458,N_16439,N_17315);
nor U18459 (N_18459,N_17811,N_17181);
and U18460 (N_18460,N_17832,N_17475);
nand U18461 (N_18461,N_17962,N_16049);
nand U18462 (N_18462,N_16559,N_16276);
or U18463 (N_18463,N_16908,N_17614);
or U18464 (N_18464,N_17451,N_17794);
and U18465 (N_18465,N_17021,N_16127);
or U18466 (N_18466,N_16574,N_16268);
nand U18467 (N_18467,N_16350,N_17693);
nor U18468 (N_18468,N_17662,N_16873);
nand U18469 (N_18469,N_16455,N_17849);
xnor U18470 (N_18470,N_16675,N_16701);
and U18471 (N_18471,N_17501,N_17726);
or U18472 (N_18472,N_16979,N_16754);
nand U18473 (N_18473,N_16461,N_17848);
and U18474 (N_18474,N_16781,N_16126);
nor U18475 (N_18475,N_17013,N_17482);
nand U18476 (N_18476,N_16646,N_16023);
nor U18477 (N_18477,N_16662,N_16688);
and U18478 (N_18478,N_17197,N_16960);
and U18479 (N_18479,N_17087,N_17917);
xnor U18480 (N_18480,N_17237,N_17714);
xnor U18481 (N_18481,N_16212,N_16447);
nand U18482 (N_18482,N_17167,N_16474);
or U18483 (N_18483,N_16515,N_16970);
and U18484 (N_18484,N_17745,N_16081);
and U18485 (N_18485,N_17462,N_17471);
nor U18486 (N_18486,N_16361,N_17300);
or U18487 (N_18487,N_17764,N_16687);
nor U18488 (N_18488,N_17420,N_17787);
and U18489 (N_18489,N_16945,N_16524);
xor U18490 (N_18490,N_16576,N_17956);
nor U18491 (N_18491,N_17725,N_17973);
nand U18492 (N_18492,N_16651,N_16954);
and U18493 (N_18493,N_17710,N_17814);
nor U18494 (N_18494,N_16173,N_16695);
xnor U18495 (N_18495,N_16136,N_17055);
nand U18496 (N_18496,N_16832,N_17354);
nand U18497 (N_18497,N_16664,N_17184);
xor U18498 (N_18498,N_16239,N_16595);
and U18499 (N_18499,N_17219,N_16974);
nor U18500 (N_18500,N_17974,N_16868);
and U18501 (N_18501,N_17078,N_16158);
nor U18502 (N_18502,N_16554,N_17752);
nor U18503 (N_18503,N_16635,N_17744);
xnor U18504 (N_18504,N_17135,N_17230);
nand U18505 (N_18505,N_16466,N_17807);
nor U18506 (N_18506,N_16555,N_17588);
and U18507 (N_18507,N_16769,N_16124);
or U18508 (N_18508,N_17616,N_16963);
and U18509 (N_18509,N_17884,N_16825);
and U18510 (N_18510,N_17397,N_16401);
and U18511 (N_18511,N_17720,N_16345);
nand U18512 (N_18512,N_17351,N_16259);
nor U18513 (N_18513,N_17763,N_17221);
and U18514 (N_18514,N_16606,N_17687);
nor U18515 (N_18515,N_17873,N_16660);
nand U18516 (N_18516,N_17262,N_17188);
and U18517 (N_18517,N_16304,N_16726);
nand U18518 (N_18518,N_16767,N_16624);
nor U18519 (N_18519,N_17238,N_16004);
and U18520 (N_18520,N_16784,N_17981);
and U18521 (N_18521,N_16091,N_16302);
nand U18522 (N_18522,N_16669,N_17030);
or U18523 (N_18523,N_17541,N_17734);
nand U18524 (N_18524,N_16509,N_17954);
and U18525 (N_18525,N_17241,N_17275);
or U18526 (N_18526,N_16089,N_16058);
or U18527 (N_18527,N_17530,N_16070);
nand U18528 (N_18528,N_17251,N_16108);
nor U18529 (N_18529,N_17727,N_16927);
or U18530 (N_18530,N_17195,N_17412);
xnor U18531 (N_18531,N_17840,N_16123);
or U18532 (N_18532,N_17808,N_16654);
nor U18533 (N_18533,N_16315,N_16622);
nor U18534 (N_18534,N_16655,N_16015);
or U18535 (N_18535,N_17349,N_17719);
xnor U18536 (N_18536,N_17995,N_17401);
and U18537 (N_18537,N_16416,N_16607);
nor U18538 (N_18538,N_16666,N_17842);
nand U18539 (N_18539,N_17209,N_16676);
nor U18540 (N_18540,N_16263,N_16925);
or U18541 (N_18541,N_17914,N_16372);
and U18542 (N_18542,N_17602,N_17570);
xor U18543 (N_18543,N_16264,N_17674);
or U18544 (N_18544,N_17683,N_17890);
xor U18545 (N_18545,N_17844,N_16269);
or U18546 (N_18546,N_16514,N_17590);
or U18547 (N_18547,N_16700,N_16882);
and U18548 (N_18548,N_17202,N_16898);
and U18549 (N_18549,N_17258,N_16312);
xor U18550 (N_18550,N_17355,N_17260);
or U18551 (N_18551,N_17916,N_16171);
xor U18552 (N_18552,N_16975,N_16029);
and U18553 (N_18553,N_16967,N_17259);
nand U18554 (N_18554,N_16957,N_17816);
or U18555 (N_18555,N_17812,N_16431);
and U18556 (N_18556,N_16711,N_17322);
nand U18557 (N_18557,N_17175,N_17560);
and U18558 (N_18558,N_17016,N_16314);
or U18559 (N_18559,N_17822,N_16141);
nor U18560 (N_18560,N_17731,N_17735);
nor U18561 (N_18561,N_17886,N_16826);
and U18562 (N_18562,N_17003,N_16989);
xor U18563 (N_18563,N_16284,N_16294);
nand U18564 (N_18564,N_17464,N_17153);
nor U18565 (N_18565,N_17518,N_17867);
and U18566 (N_18566,N_17542,N_16750);
nand U18567 (N_18567,N_16325,N_17044);
xnor U18568 (N_18568,N_16532,N_16516);
nor U18569 (N_18569,N_16691,N_16221);
and U18570 (N_18570,N_16780,N_17584);
nor U18571 (N_18571,N_17266,N_17909);
or U18572 (N_18572,N_17733,N_16693);
or U18573 (N_18573,N_16834,N_17361);
nand U18574 (N_18574,N_17878,N_17796);
xor U18575 (N_18575,N_17644,N_16730);
nand U18576 (N_18576,N_17640,N_17888);
and U18577 (N_18577,N_16959,N_16399);
and U18578 (N_18578,N_17661,N_17337);
nor U18579 (N_18579,N_17422,N_16389);
nor U18580 (N_18580,N_16602,N_17005);
nand U18581 (N_18581,N_16317,N_16419);
nand U18582 (N_18582,N_16473,N_17035);
or U18583 (N_18583,N_16623,N_17576);
nor U18584 (N_18584,N_16405,N_16288);
nor U18585 (N_18585,N_17938,N_16119);
nand U18586 (N_18586,N_16869,N_17651);
xnor U18587 (N_18587,N_16135,N_17293);
and U18588 (N_18588,N_17668,N_17163);
or U18589 (N_18589,N_17141,N_16512);
nand U18590 (N_18590,N_17276,N_16349);
or U18591 (N_18591,N_17239,N_16410);
nor U18592 (N_18592,N_17578,N_17709);
nand U18593 (N_18593,N_17229,N_16579);
xor U18594 (N_18594,N_17821,N_16441);
and U18595 (N_18595,N_16852,N_16025);
and U18596 (N_18596,N_17310,N_16233);
xnor U18597 (N_18597,N_17414,N_17789);
or U18598 (N_18598,N_16786,N_17915);
or U18599 (N_18599,N_16353,N_17218);
nor U18600 (N_18600,N_17486,N_17391);
xor U18601 (N_18601,N_17759,N_16567);
or U18602 (N_18602,N_16347,N_17612);
nor U18603 (N_18603,N_17254,N_16009);
or U18604 (N_18604,N_17316,N_16631);
nand U18605 (N_18605,N_17264,N_16116);
nand U18606 (N_18606,N_17376,N_16564);
nand U18607 (N_18607,N_17205,N_17095);
and U18608 (N_18608,N_16953,N_17622);
or U18609 (N_18609,N_17967,N_17767);
xor U18610 (N_18610,N_16107,N_16884);
nor U18611 (N_18611,N_16630,N_16362);
nand U18612 (N_18612,N_17589,N_17099);
and U18613 (N_18613,N_16456,N_17623);
and U18614 (N_18614,N_17051,N_16213);
nand U18615 (N_18615,N_17052,N_17212);
nor U18616 (N_18616,N_16740,N_16860);
and U18617 (N_18617,N_17317,N_17270);
nor U18618 (N_18618,N_17863,N_17507);
or U18619 (N_18619,N_17955,N_17694);
xnor U18620 (N_18620,N_17130,N_17574);
nor U18621 (N_18621,N_16903,N_17298);
xor U18622 (N_18622,N_17882,N_16457);
and U18623 (N_18623,N_17519,N_17150);
and U18624 (N_18624,N_16279,N_16075);
or U18625 (N_18625,N_16022,N_17467);
and U18626 (N_18626,N_16006,N_17077);
nor U18627 (N_18627,N_16435,N_16536);
nor U18628 (N_18628,N_16193,N_16301);
or U18629 (N_18629,N_16502,N_17154);
or U18630 (N_18630,N_17377,N_16714);
and U18631 (N_18631,N_16909,N_16583);
nor U18632 (N_18632,N_17180,N_16808);
nand U18633 (N_18633,N_16639,N_17898);
and U18634 (N_18634,N_16741,N_17526);
nor U18635 (N_18635,N_17768,N_16459);
nand U18636 (N_18636,N_17353,N_17621);
nand U18637 (N_18637,N_16537,N_17959);
nor U18638 (N_18638,N_16962,N_17014);
or U18639 (N_18639,N_16984,N_17067);
or U18640 (N_18640,N_16617,N_17860);
nor U18641 (N_18641,N_17437,N_16056);
and U18642 (N_18642,N_17404,N_17800);
and U18643 (N_18643,N_17145,N_16187);
and U18644 (N_18644,N_17331,N_16958);
or U18645 (N_18645,N_16828,N_16491);
nor U18646 (N_18646,N_17673,N_17306);
or U18647 (N_18647,N_17073,N_17866);
xor U18648 (N_18648,N_17833,N_16373);
xor U18649 (N_18649,N_17927,N_16743);
nor U18650 (N_18650,N_16106,N_17596);
and U18651 (N_18651,N_17143,N_16578);
or U18652 (N_18652,N_16339,N_17635);
or U18653 (N_18653,N_17066,N_17253);
or U18654 (N_18654,N_17611,N_16969);
nor U18655 (N_18655,N_16185,N_16907);
nor U18656 (N_18656,N_16749,N_16411);
nand U18657 (N_18657,N_16406,N_16480);
or U18658 (N_18658,N_16977,N_16562);
nor U18659 (N_18659,N_16485,N_16799);
or U18660 (N_18660,N_16620,N_17545);
xor U18661 (N_18661,N_17993,N_17707);
nor U18662 (N_18662,N_17129,N_16865);
nand U18663 (N_18663,N_17421,N_17703);
nor U18664 (N_18664,N_16525,N_17871);
or U18665 (N_18665,N_17975,N_17423);
and U18666 (N_18666,N_17835,N_16080);
xnor U18667 (N_18667,N_17647,N_16810);
nor U18668 (N_18668,N_16964,N_17718);
nand U18669 (N_18669,N_16657,N_16071);
and U18670 (N_18670,N_17872,N_16375);
and U18671 (N_18671,N_16822,N_17432);
xor U18672 (N_18672,N_16947,N_17140);
or U18673 (N_18673,N_17920,N_16827);
nand U18674 (N_18674,N_17032,N_16719);
nor U18675 (N_18675,N_16592,N_16760);
xnor U18676 (N_18676,N_16142,N_16745);
nor U18677 (N_18677,N_17641,N_17392);
and U18678 (N_18678,N_16468,N_17652);
nand U18679 (N_18679,N_16608,N_17826);
or U18680 (N_18680,N_16417,N_17689);
xnor U18681 (N_18681,N_17190,N_17893);
nand U18682 (N_18682,N_17930,N_16899);
or U18683 (N_18683,N_17818,N_16686);
xor U18684 (N_18684,N_16851,N_16748);
nand U18685 (N_18685,N_17211,N_16858);
nand U18686 (N_18686,N_17569,N_17952);
and U18687 (N_18687,N_17947,N_17627);
or U18688 (N_18688,N_17810,N_17206);
nand U18689 (N_18689,N_16645,N_16140);
or U18690 (N_18690,N_16330,N_16540);
or U18691 (N_18691,N_17493,N_17619);
nand U18692 (N_18692,N_17853,N_17699);
and U18693 (N_18693,N_17199,N_16656);
or U18694 (N_18694,N_17089,N_16797);
nand U18695 (N_18695,N_16412,N_16230);
nand U18696 (N_18696,N_17368,N_17124);
nand U18697 (N_18697,N_17546,N_16383);
nor U18698 (N_18698,N_16366,N_17765);
nor U18699 (N_18699,N_17233,N_16501);
and U18700 (N_18700,N_16736,N_17503);
nand U18701 (N_18701,N_17911,N_16388);
nor U18702 (N_18702,N_16830,N_17948);
xor U18703 (N_18703,N_17776,N_17755);
nand U18704 (N_18704,N_17405,N_16824);
xor U18705 (N_18705,N_16517,N_16365);
xnor U18706 (N_18706,N_17112,N_17009);
nor U18707 (N_18707,N_16603,N_16202);
or U18708 (N_18708,N_17096,N_16222);
xnor U18709 (N_18709,N_17830,N_16452);
nor U18710 (N_18710,N_17287,N_16342);
and U18711 (N_18711,N_17020,N_17159);
or U18712 (N_18712,N_16924,N_16113);
or U18713 (N_18713,N_17034,N_17062);
nor U18714 (N_18714,N_17403,N_16853);
and U18715 (N_18715,N_17494,N_16464);
nor U18716 (N_18716,N_17413,N_17531);
or U18717 (N_18717,N_16469,N_16483);
nand U18718 (N_18718,N_17101,N_16432);
nor U18719 (N_18719,N_17272,N_16159);
or U18720 (N_18720,N_16758,N_16096);
and U18721 (N_18721,N_17894,N_16665);
or U18722 (N_18722,N_17660,N_16427);
and U18723 (N_18723,N_17572,N_17730);
nor U18724 (N_18724,N_16995,N_16855);
or U18725 (N_18725,N_17784,N_17936);
nor U18726 (N_18726,N_16543,N_17695);
or U18727 (N_18727,N_16487,N_17549);
and U18728 (N_18728,N_17179,N_16787);
nand U18729 (N_18729,N_17116,N_17352);
nand U18730 (N_18730,N_17891,N_17636);
nor U18731 (N_18731,N_17865,N_16364);
and U18732 (N_18732,N_16930,N_16893);
nand U18733 (N_18733,N_17932,N_17609);
or U18734 (N_18734,N_16874,N_17094);
xnor U18735 (N_18735,N_17408,N_17216);
or U18736 (N_18736,N_16033,N_17390);
nor U18737 (N_18737,N_17208,N_16122);
nand U18738 (N_18738,N_16044,N_17010);
or U18739 (N_18739,N_16938,N_17857);
xor U18740 (N_18740,N_16673,N_16235);
or U18741 (N_18741,N_17282,N_16697);
or U18742 (N_18742,N_17076,N_16849);
nand U18743 (N_18743,N_17847,N_16723);
or U18744 (N_18744,N_16099,N_17380);
nand U18745 (N_18745,N_17369,N_17512);
xnor U18746 (N_18746,N_17048,N_17382);
nand U18747 (N_18747,N_16505,N_16892);
or U18748 (N_18748,N_17452,N_16670);
nand U18749 (N_18749,N_17225,N_16844);
or U18750 (N_18750,N_17445,N_16182);
nor U18751 (N_18751,N_16189,N_17716);
xnor U18752 (N_18752,N_17117,N_17305);
or U18753 (N_18753,N_17036,N_16428);
nor U18754 (N_18754,N_17971,N_17302);
xnor U18755 (N_18755,N_17739,N_16246);
or U18756 (N_18756,N_17134,N_16224);
xor U18757 (N_18757,N_16993,N_17045);
and U18758 (N_18758,N_16879,N_16407);
nor U18759 (N_18759,N_16819,N_16584);
xor U18760 (N_18760,N_17409,N_17002);
and U18761 (N_18761,N_16829,N_16497);
xor U18762 (N_18762,N_16859,N_17131);
and U18763 (N_18763,N_17557,N_17039);
nand U18764 (N_18764,N_16251,N_17069);
xnor U18765 (N_18765,N_16038,N_16104);
xor U18766 (N_18766,N_16494,N_16823);
nor U18767 (N_18767,N_17263,N_16379);
or U18768 (N_18768,N_16429,N_17943);
nand U18769 (N_18769,N_16997,N_16121);
and U18770 (N_18770,N_17937,N_16922);
xnor U18771 (N_18771,N_16588,N_17359);
or U18772 (N_18772,N_16103,N_17672);
xnor U18773 (N_18773,N_16721,N_16110);
nor U18774 (N_18774,N_16598,N_17736);
or U18775 (N_18775,N_17080,N_16840);
or U18776 (N_18776,N_16278,N_16065);
or U18777 (N_18777,N_17724,N_16778);
nand U18778 (N_18778,N_17268,N_17378);
or U18779 (N_18779,N_17910,N_16684);
nand U18780 (N_18780,N_16732,N_16920);
nor U18781 (N_18781,N_16533,N_16965);
or U18782 (N_18782,N_16806,N_17925);
and U18783 (N_18783,N_17961,N_16219);
nor U18784 (N_18784,N_17024,N_17608);
xnor U18785 (N_18785,N_17827,N_16050);
nor U18786 (N_18786,N_16052,N_16208);
or U18787 (N_18787,N_16179,N_17761);
nand U18788 (N_18788,N_17047,N_17772);
and U18789 (N_18789,N_17356,N_17176);
nor U18790 (N_18790,N_17236,N_16176);
and U18791 (N_18791,N_16796,N_16846);
and U18792 (N_18792,N_16596,N_16941);
nand U18793 (N_18793,N_16880,N_17185);
xnor U18794 (N_18794,N_17940,N_16642);
or U18795 (N_18795,N_17935,N_16205);
and U18796 (N_18796,N_17648,N_16449);
or U18797 (N_18797,N_16191,N_17831);
nand U18798 (N_18798,N_17123,N_17183);
nor U18799 (N_18799,N_17670,N_16117);
or U18800 (N_18800,N_16890,N_17704);
nand U18801 (N_18801,N_17023,N_17746);
or U18802 (N_18802,N_17441,N_16300);
nand U18803 (N_18803,N_17861,N_16324);
nand U18804 (N_18804,N_17613,N_17436);
xnor U18805 (N_18805,N_17902,N_17224);
nand U18806 (N_18806,N_16078,N_17056);
and U18807 (N_18807,N_17802,N_16522);
or U18808 (N_18808,N_16913,N_17809);
nand U18809 (N_18809,N_16111,N_16011);
nor U18810 (N_18810,N_17120,N_16867);
xor U18811 (N_18811,N_17504,N_16337);
nor U18812 (N_18812,N_17440,N_17691);
or U18813 (N_18813,N_16267,N_16513);
nor U18814 (N_18814,N_16046,N_17737);
or U18815 (N_18815,N_16472,N_17168);
or U18816 (N_18816,N_16541,N_16568);
nand U18817 (N_18817,N_16618,N_16203);
and U18818 (N_18818,N_16460,N_17285);
xor U18819 (N_18819,N_16030,N_17773);
nor U18820 (N_18820,N_17311,N_17939);
nand U18821 (N_18821,N_17760,N_17193);
nor U18822 (N_18822,N_17628,N_16677);
nand U18823 (N_18823,N_17966,N_16531);
xor U18824 (N_18824,N_17537,N_16422);
nand U18825 (N_18825,N_16816,N_17312);
xnor U18826 (N_18826,N_16130,N_17483);
nand U18827 (N_18827,N_17658,N_17144);
nor U18828 (N_18828,N_16471,N_16538);
xor U18829 (N_18829,N_17158,N_16220);
nor U18830 (N_18830,N_17980,N_17923);
nand U18831 (N_18831,N_17472,N_17837);
nor U18832 (N_18832,N_17680,N_17174);
and U18833 (N_18833,N_16032,N_17001);
nor U18834 (N_18834,N_16621,N_17868);
and U18835 (N_18835,N_16020,N_16681);
xnor U18836 (N_18836,N_17017,N_17407);
or U18837 (N_18837,N_17274,N_16923);
or U18838 (N_18838,N_17575,N_17177);
or U18839 (N_18839,N_17433,N_17227);
or U18840 (N_18840,N_16653,N_16297);
and U18841 (N_18841,N_17165,N_16864);
nand U18842 (N_18842,N_16996,N_16248);
or U18843 (N_18843,N_17912,N_17049);
nor U18844 (N_18844,N_16034,N_16215);
and U18845 (N_18845,N_16839,N_17829);
nand U18846 (N_18846,N_17444,N_16788);
nand U18847 (N_18847,N_17946,N_17587);
nor U18848 (N_18848,N_16354,N_17133);
or U18849 (N_18849,N_16707,N_17366);
nand U18850 (N_18850,N_17813,N_17217);
nand U18851 (N_18851,N_16010,N_17333);
xor U18852 (N_18852,N_17598,N_17838);
and U18853 (N_18853,N_17000,N_16090);
xor U18854 (N_18854,N_17223,N_17297);
and U18855 (N_18855,N_17063,N_16629);
nand U18856 (N_18856,N_17011,N_16814);
and U18857 (N_18857,N_17479,N_16756);
nand U18858 (N_18858,N_17164,N_16735);
nor U18859 (N_18859,N_17639,N_16900);
nor U18860 (N_18860,N_17342,N_17072);
nand U18861 (N_18861,N_16190,N_17620);
or U18862 (N_18862,N_17540,N_17963);
xor U18863 (N_18863,N_16981,N_17629);
nand U18864 (N_18864,N_16705,N_16036);
nor U18865 (N_18865,N_16813,N_17562);
and U18866 (N_18866,N_17520,N_17957);
or U18867 (N_18867,N_17395,N_16274);
nand U18868 (N_18868,N_16652,N_16261);
nand U18869 (N_18869,N_17964,N_16371);
nand U18870 (N_18870,N_16238,N_16125);
or U18871 (N_18871,N_16214,N_17864);
nand U18872 (N_18872,N_17945,N_17497);
and U18873 (N_18873,N_16216,N_16064);
or U18874 (N_18874,N_17876,N_17669);
and U18875 (N_18875,N_17053,N_17960);
and U18876 (N_18876,N_16357,N_16499);
xnor U18877 (N_18877,N_16149,N_17856);
nor U18878 (N_18878,N_16308,N_16772);
nand U18879 (N_18879,N_17879,N_16067);
nand U18880 (N_18880,N_17998,N_17646);
nand U18881 (N_18881,N_17563,N_16352);
xor U18882 (N_18882,N_17659,N_17663);
or U18883 (N_18883,N_17547,N_16551);
xnor U18884 (N_18884,N_17344,N_16042);
and U18885 (N_18885,N_16643,N_17517);
or U18886 (N_18886,N_16519,N_17738);
and U18887 (N_18887,N_16316,N_16866);
xnor U18888 (N_18888,N_16644,N_17243);
nor U18889 (N_18889,N_17558,N_16098);
and U18890 (N_18890,N_17632,N_17090);
xnor U18891 (N_18891,N_17477,N_17601);
nor U18892 (N_18892,N_16523,N_17484);
or U18893 (N_18893,N_17128,N_17136);
nor U18894 (N_18894,N_16035,N_17824);
nand U18895 (N_18895,N_16872,N_16283);
xnor U18896 (N_18896,N_16696,N_17678);
xnor U18897 (N_18897,N_16305,N_16593);
and U18898 (N_18898,N_17881,N_17677);
and U18899 (N_18899,N_16708,N_17425);
xnor U18900 (N_18900,N_16926,N_16725);
and U18901 (N_18901,N_17400,N_16394);
nand U18902 (N_18902,N_17741,N_16329);
xor U18903 (N_18903,N_17490,N_17492);
xnor U18904 (N_18904,N_17771,N_17951);
nor U18905 (N_18905,N_17553,N_16737);
nor U18906 (N_18906,N_17022,N_17897);
or U18907 (N_18907,N_17664,N_17638);
nand U18908 (N_18908,N_17007,N_16054);
xor U18909 (N_18909,N_17976,N_17987);
nor U18910 (N_18910,N_17579,N_16262);
and U18911 (N_18911,N_17931,N_17288);
and U18912 (N_18912,N_16710,N_17326);
nor U18913 (N_18913,N_17684,N_16152);
nor U18914 (N_18914,N_17084,N_16131);
or U18915 (N_18915,N_17108,N_17046);
nand U18916 (N_18916,N_17058,N_16678);
nor U18917 (N_18917,N_16232,N_17681);
and U18918 (N_18918,N_16281,N_16450);
nor U18919 (N_18919,N_17700,N_16663);
nand U18920 (N_18920,N_16146,N_16557);
nand U18921 (N_18921,N_16343,N_16817);
nand U18922 (N_18922,N_17859,N_17406);
and U18923 (N_18923,N_16510,N_17790);
nor U18924 (N_18924,N_17997,N_16076);
or U18925 (N_18925,N_17850,N_16534);
and U18926 (N_18926,N_17571,N_16257);
or U18927 (N_18927,N_17384,N_16956);
nand U18928 (N_18928,N_16939,N_17906);
and U18929 (N_18929,N_16057,N_16470);
xnor U18930 (N_18930,N_16698,N_17301);
nand U18931 (N_18931,N_17256,N_16821);
or U18932 (N_18932,N_16943,N_16847);
xnor U18933 (N_18933,N_17292,N_16143);
xnor U18934 (N_18934,N_16155,N_17091);
and U18935 (N_18935,N_17255,N_16344);
and U18936 (N_18936,N_17533,N_17299);
xnor U18937 (N_18937,N_16282,N_17757);
nor U18938 (N_18938,N_16019,N_16156);
nor U18939 (N_18939,N_16434,N_16183);
xor U18940 (N_18940,N_16415,N_17265);
and U18941 (N_18941,N_16910,N_16299);
and U18942 (N_18942,N_17138,N_17564);
and U18943 (N_18943,N_16818,N_16481);
or U18944 (N_18944,N_17012,N_17845);
nor U18945 (N_18945,N_17697,N_16086);
or U18946 (N_18946,N_16040,N_16164);
and U18947 (N_18947,N_16715,N_16446);
and U18948 (N_18948,N_16626,N_17994);
nand U18949 (N_18949,N_16488,N_17040);
xor U18950 (N_18950,N_16842,N_17115);
nor U18951 (N_18951,N_16807,N_16919);
and U18952 (N_18952,N_16132,N_17825);
nor U18953 (N_18953,N_17198,N_16360);
or U18954 (N_18954,N_16421,N_16986);
nand U18955 (N_18955,N_16973,N_16430);
xnor U18956 (N_18956,N_17038,N_17191);
nor U18957 (N_18957,N_16323,N_17417);
or U18958 (N_18958,N_16115,N_16320);
or U18959 (N_18959,N_17328,N_16396);
nor U18960 (N_18960,N_16738,N_17210);
or U18961 (N_18961,N_17201,N_17903);
nor U18962 (N_18962,N_17978,N_17924);
nor U18963 (N_18963,N_17474,N_16414);
and U18964 (N_18964,N_17279,N_17583);
or U18965 (N_18965,N_16671,N_16002);
or U18966 (N_18966,N_16327,N_16836);
nand U18967 (N_18967,N_17543,N_17082);
xor U18968 (N_18968,N_17373,N_16303);
xor U18969 (N_18969,N_16774,N_16341);
or U18970 (N_18970,N_17149,N_16031);
nand U18971 (N_18971,N_16195,N_17029);
or U18972 (N_18972,N_17085,N_16192);
nand U18973 (N_18973,N_16258,N_17729);
nor U18974 (N_18974,N_17750,N_16425);
nand U18975 (N_18975,N_17364,N_16051);
xnor U18976 (N_18976,N_17561,N_16912);
or U18977 (N_18977,N_16589,N_16569);
nor U18978 (N_18978,N_17152,N_17595);
nand U18979 (N_18979,N_16393,N_16789);
and U18980 (N_18980,N_16043,N_16102);
xor U18981 (N_18981,N_16627,N_16734);
and U18982 (N_18982,N_16157,N_17496);
or U18983 (N_18983,N_17139,N_17933);
or U18984 (N_18984,N_17132,N_16017);
xor U18985 (N_18985,N_16800,N_16889);
or U18986 (N_18986,N_16729,N_16961);
or U18987 (N_18987,N_16871,N_16151);
and U18988 (N_18988,N_16932,N_16227);
nor U18989 (N_18989,N_16270,N_16779);
or U18990 (N_18990,N_16940,N_16356);
nor U18991 (N_18991,N_16084,N_17783);
or U18992 (N_18992,N_16133,N_17273);
xor U18993 (N_18993,N_17513,N_17846);
nor U18994 (N_18994,N_16805,N_17439);
xor U18995 (N_18995,N_16529,N_17372);
nor U18996 (N_18996,N_17280,N_16201);
nand U18997 (N_18997,N_16768,N_16249);
and U18998 (N_18998,N_16318,N_16640);
and U18999 (N_18999,N_17606,N_16200);
nor U19000 (N_19000,N_16722,N_16759);
or U19001 (N_19001,N_17946,N_17345);
nand U19002 (N_19002,N_17457,N_17099);
and U19003 (N_19003,N_17201,N_17226);
and U19004 (N_19004,N_16887,N_16287);
nand U19005 (N_19005,N_17986,N_17052);
nor U19006 (N_19006,N_16302,N_17042);
and U19007 (N_19007,N_17631,N_17849);
and U19008 (N_19008,N_17369,N_16921);
xor U19009 (N_19009,N_17204,N_16273);
or U19010 (N_19010,N_17882,N_17186);
or U19011 (N_19011,N_16519,N_17691);
nand U19012 (N_19012,N_17396,N_16466);
nor U19013 (N_19013,N_16876,N_16659);
or U19014 (N_19014,N_16968,N_17952);
xnor U19015 (N_19015,N_16611,N_17127);
nand U19016 (N_19016,N_16047,N_16674);
or U19017 (N_19017,N_17876,N_16482);
or U19018 (N_19018,N_17693,N_17227);
nand U19019 (N_19019,N_16022,N_17619);
xor U19020 (N_19020,N_17727,N_17988);
nand U19021 (N_19021,N_17659,N_17342);
nand U19022 (N_19022,N_16232,N_17991);
or U19023 (N_19023,N_17019,N_17502);
nor U19024 (N_19024,N_16628,N_17340);
and U19025 (N_19025,N_16048,N_17667);
nand U19026 (N_19026,N_17176,N_17191);
xor U19027 (N_19027,N_17124,N_16833);
and U19028 (N_19028,N_16940,N_16612);
nor U19029 (N_19029,N_17386,N_17072);
or U19030 (N_19030,N_16914,N_16635);
and U19031 (N_19031,N_16009,N_16431);
xor U19032 (N_19032,N_17808,N_16020);
or U19033 (N_19033,N_17200,N_16094);
or U19034 (N_19034,N_16646,N_16994);
xor U19035 (N_19035,N_16029,N_17248);
nand U19036 (N_19036,N_16177,N_16018);
nand U19037 (N_19037,N_17239,N_16833);
xor U19038 (N_19038,N_17641,N_16172);
xor U19039 (N_19039,N_17545,N_17444);
nand U19040 (N_19040,N_16812,N_17841);
nand U19041 (N_19041,N_16502,N_16629);
nand U19042 (N_19042,N_17204,N_16408);
nor U19043 (N_19043,N_17583,N_16599);
xor U19044 (N_19044,N_17754,N_17489);
nand U19045 (N_19045,N_16370,N_16961);
or U19046 (N_19046,N_17825,N_17649);
xor U19047 (N_19047,N_16450,N_17742);
nand U19048 (N_19048,N_16497,N_17699);
xor U19049 (N_19049,N_17441,N_17685);
nand U19050 (N_19050,N_17224,N_17916);
and U19051 (N_19051,N_17843,N_16264);
nor U19052 (N_19052,N_17049,N_16057);
or U19053 (N_19053,N_17509,N_16066);
nor U19054 (N_19054,N_17230,N_16394);
xnor U19055 (N_19055,N_17779,N_16799);
or U19056 (N_19056,N_16681,N_16240);
or U19057 (N_19057,N_17111,N_16518);
or U19058 (N_19058,N_16023,N_17633);
xor U19059 (N_19059,N_16787,N_17530);
nor U19060 (N_19060,N_16485,N_17202);
and U19061 (N_19061,N_16794,N_17370);
nand U19062 (N_19062,N_16207,N_16478);
nand U19063 (N_19063,N_16412,N_17317);
nor U19064 (N_19064,N_16546,N_17473);
nand U19065 (N_19065,N_17990,N_17236);
nand U19066 (N_19066,N_17117,N_16595);
and U19067 (N_19067,N_17883,N_17145);
or U19068 (N_19068,N_16202,N_16441);
and U19069 (N_19069,N_16320,N_17065);
nor U19070 (N_19070,N_17979,N_16827);
xor U19071 (N_19071,N_16612,N_17413);
or U19072 (N_19072,N_17284,N_17222);
and U19073 (N_19073,N_16653,N_17221);
xnor U19074 (N_19074,N_17456,N_16447);
xnor U19075 (N_19075,N_16745,N_16905);
and U19076 (N_19076,N_16213,N_17288);
and U19077 (N_19077,N_17580,N_16221);
nor U19078 (N_19078,N_17768,N_16346);
and U19079 (N_19079,N_17293,N_17340);
or U19080 (N_19080,N_16028,N_17017);
nand U19081 (N_19081,N_17157,N_17973);
and U19082 (N_19082,N_16946,N_17439);
nor U19083 (N_19083,N_16792,N_17217);
or U19084 (N_19084,N_17387,N_16697);
nand U19085 (N_19085,N_17074,N_16974);
and U19086 (N_19086,N_17704,N_16901);
nand U19087 (N_19087,N_17359,N_17875);
nor U19088 (N_19088,N_16565,N_16784);
and U19089 (N_19089,N_16120,N_16889);
nand U19090 (N_19090,N_17458,N_17518);
nor U19091 (N_19091,N_16284,N_17301);
and U19092 (N_19092,N_17967,N_17490);
and U19093 (N_19093,N_16725,N_17523);
nand U19094 (N_19094,N_16183,N_17528);
nor U19095 (N_19095,N_17518,N_16910);
nand U19096 (N_19096,N_17673,N_17293);
or U19097 (N_19097,N_16418,N_17483);
and U19098 (N_19098,N_17600,N_16375);
xor U19099 (N_19099,N_16280,N_17768);
or U19100 (N_19100,N_16211,N_17300);
or U19101 (N_19101,N_16657,N_16653);
xnor U19102 (N_19102,N_16030,N_17616);
and U19103 (N_19103,N_16798,N_16753);
nand U19104 (N_19104,N_16162,N_17017);
and U19105 (N_19105,N_16929,N_17478);
and U19106 (N_19106,N_16134,N_17362);
or U19107 (N_19107,N_16229,N_17736);
or U19108 (N_19108,N_17509,N_17281);
nor U19109 (N_19109,N_16067,N_16875);
nand U19110 (N_19110,N_16671,N_17310);
nand U19111 (N_19111,N_16506,N_16516);
nor U19112 (N_19112,N_17872,N_17948);
or U19113 (N_19113,N_16115,N_17668);
xnor U19114 (N_19114,N_17352,N_16578);
or U19115 (N_19115,N_16163,N_16506);
nand U19116 (N_19116,N_17184,N_16742);
nor U19117 (N_19117,N_17746,N_17353);
nand U19118 (N_19118,N_17004,N_17997);
nor U19119 (N_19119,N_16210,N_16393);
nand U19120 (N_19120,N_17573,N_16564);
or U19121 (N_19121,N_17146,N_17318);
or U19122 (N_19122,N_16378,N_17721);
and U19123 (N_19123,N_16280,N_17806);
nand U19124 (N_19124,N_17259,N_17962);
xor U19125 (N_19125,N_16839,N_16885);
nor U19126 (N_19126,N_17646,N_17776);
nand U19127 (N_19127,N_16730,N_16560);
or U19128 (N_19128,N_17353,N_16040);
xnor U19129 (N_19129,N_17192,N_17511);
or U19130 (N_19130,N_17945,N_16595);
nand U19131 (N_19131,N_17324,N_17235);
xnor U19132 (N_19132,N_16020,N_16023);
xor U19133 (N_19133,N_16852,N_17151);
xor U19134 (N_19134,N_17120,N_16757);
and U19135 (N_19135,N_17764,N_17273);
or U19136 (N_19136,N_16274,N_17141);
nor U19137 (N_19137,N_17935,N_16954);
or U19138 (N_19138,N_16142,N_17554);
or U19139 (N_19139,N_16848,N_16142);
xor U19140 (N_19140,N_16941,N_16377);
or U19141 (N_19141,N_17385,N_17954);
and U19142 (N_19142,N_17675,N_17524);
or U19143 (N_19143,N_16584,N_17461);
xor U19144 (N_19144,N_17541,N_16949);
xor U19145 (N_19145,N_16488,N_16228);
xor U19146 (N_19146,N_16245,N_17079);
or U19147 (N_19147,N_17493,N_16143);
xor U19148 (N_19148,N_16050,N_17001);
nand U19149 (N_19149,N_17028,N_17158);
and U19150 (N_19150,N_17315,N_17189);
or U19151 (N_19151,N_17124,N_16135);
or U19152 (N_19152,N_16554,N_16111);
nor U19153 (N_19153,N_17431,N_17612);
xor U19154 (N_19154,N_17264,N_16522);
and U19155 (N_19155,N_17858,N_16923);
nand U19156 (N_19156,N_17736,N_17112);
nor U19157 (N_19157,N_16518,N_17334);
or U19158 (N_19158,N_16707,N_17007);
xor U19159 (N_19159,N_16926,N_16946);
xor U19160 (N_19160,N_17653,N_16533);
nand U19161 (N_19161,N_16852,N_16199);
nor U19162 (N_19162,N_17007,N_17194);
nand U19163 (N_19163,N_17307,N_16782);
xnor U19164 (N_19164,N_16799,N_17862);
or U19165 (N_19165,N_17329,N_17739);
and U19166 (N_19166,N_17592,N_16798);
nand U19167 (N_19167,N_17722,N_17763);
xor U19168 (N_19168,N_17960,N_16895);
xor U19169 (N_19169,N_16706,N_16268);
xor U19170 (N_19170,N_16844,N_17574);
and U19171 (N_19171,N_17494,N_16483);
and U19172 (N_19172,N_17723,N_17175);
nand U19173 (N_19173,N_16886,N_16829);
nand U19174 (N_19174,N_17073,N_16439);
or U19175 (N_19175,N_17810,N_17469);
nand U19176 (N_19176,N_17976,N_16261);
nand U19177 (N_19177,N_17472,N_16569);
xnor U19178 (N_19178,N_17137,N_17645);
and U19179 (N_19179,N_17719,N_17511);
xor U19180 (N_19180,N_17760,N_16321);
nor U19181 (N_19181,N_16301,N_17926);
nor U19182 (N_19182,N_16391,N_16368);
nor U19183 (N_19183,N_16262,N_17308);
or U19184 (N_19184,N_16962,N_16986);
nor U19185 (N_19185,N_17716,N_16622);
or U19186 (N_19186,N_17249,N_16903);
or U19187 (N_19187,N_17583,N_17714);
xnor U19188 (N_19188,N_17237,N_17512);
nand U19189 (N_19189,N_16303,N_17462);
nor U19190 (N_19190,N_16121,N_17961);
and U19191 (N_19191,N_16415,N_17523);
or U19192 (N_19192,N_17907,N_16486);
or U19193 (N_19193,N_16269,N_17579);
or U19194 (N_19194,N_16332,N_16965);
nor U19195 (N_19195,N_17848,N_16898);
xnor U19196 (N_19196,N_16511,N_17119);
and U19197 (N_19197,N_17660,N_16573);
and U19198 (N_19198,N_16311,N_17132);
and U19199 (N_19199,N_16814,N_17547);
nand U19200 (N_19200,N_17744,N_16293);
or U19201 (N_19201,N_16648,N_17344);
or U19202 (N_19202,N_17739,N_17351);
or U19203 (N_19203,N_17258,N_16429);
nand U19204 (N_19204,N_17225,N_17205);
or U19205 (N_19205,N_17662,N_16137);
and U19206 (N_19206,N_17960,N_17634);
nand U19207 (N_19207,N_17292,N_17929);
nor U19208 (N_19208,N_17484,N_16696);
or U19209 (N_19209,N_17404,N_17798);
or U19210 (N_19210,N_17539,N_16758);
nand U19211 (N_19211,N_17072,N_17193);
and U19212 (N_19212,N_17132,N_16105);
or U19213 (N_19213,N_16474,N_17473);
and U19214 (N_19214,N_16570,N_16571);
nand U19215 (N_19215,N_16149,N_17804);
xnor U19216 (N_19216,N_16102,N_16455);
and U19217 (N_19217,N_16002,N_17038);
nand U19218 (N_19218,N_17320,N_17588);
nor U19219 (N_19219,N_17033,N_17927);
nand U19220 (N_19220,N_17227,N_17549);
nand U19221 (N_19221,N_17970,N_16979);
nor U19222 (N_19222,N_17832,N_16544);
nand U19223 (N_19223,N_17583,N_16716);
and U19224 (N_19224,N_17543,N_16524);
xnor U19225 (N_19225,N_17534,N_16813);
nand U19226 (N_19226,N_17381,N_16247);
nand U19227 (N_19227,N_17963,N_17209);
and U19228 (N_19228,N_17368,N_17798);
and U19229 (N_19229,N_17438,N_16077);
xnor U19230 (N_19230,N_16768,N_16436);
and U19231 (N_19231,N_16155,N_16904);
nand U19232 (N_19232,N_16460,N_16279);
nor U19233 (N_19233,N_16676,N_16490);
nand U19234 (N_19234,N_16396,N_16156);
nand U19235 (N_19235,N_17077,N_17711);
nor U19236 (N_19236,N_16001,N_16548);
and U19237 (N_19237,N_17477,N_16155);
xor U19238 (N_19238,N_16703,N_16944);
nand U19239 (N_19239,N_16290,N_16265);
or U19240 (N_19240,N_17262,N_16013);
nor U19241 (N_19241,N_16249,N_16304);
nor U19242 (N_19242,N_16293,N_16712);
xor U19243 (N_19243,N_17791,N_17685);
nor U19244 (N_19244,N_16809,N_16179);
xnor U19245 (N_19245,N_17153,N_16654);
and U19246 (N_19246,N_17171,N_16084);
xor U19247 (N_19247,N_17191,N_17845);
or U19248 (N_19248,N_16069,N_16549);
or U19249 (N_19249,N_16872,N_17497);
xnor U19250 (N_19250,N_17516,N_16629);
nor U19251 (N_19251,N_16004,N_16947);
nand U19252 (N_19252,N_16862,N_16606);
nor U19253 (N_19253,N_17198,N_16629);
nand U19254 (N_19254,N_16704,N_17730);
xor U19255 (N_19255,N_17787,N_16595);
nor U19256 (N_19256,N_17899,N_17951);
or U19257 (N_19257,N_17813,N_16706);
and U19258 (N_19258,N_17736,N_16020);
xor U19259 (N_19259,N_16357,N_17790);
nand U19260 (N_19260,N_16725,N_17124);
xor U19261 (N_19261,N_16088,N_17565);
or U19262 (N_19262,N_17244,N_17697);
nand U19263 (N_19263,N_17234,N_16733);
xnor U19264 (N_19264,N_16830,N_17410);
nand U19265 (N_19265,N_17191,N_17202);
and U19266 (N_19266,N_17919,N_16212);
and U19267 (N_19267,N_16181,N_16989);
and U19268 (N_19268,N_17246,N_16431);
nand U19269 (N_19269,N_17784,N_16834);
nand U19270 (N_19270,N_17066,N_16897);
and U19271 (N_19271,N_16091,N_17837);
xor U19272 (N_19272,N_16237,N_17234);
nand U19273 (N_19273,N_16491,N_16858);
and U19274 (N_19274,N_17762,N_17371);
nand U19275 (N_19275,N_17782,N_16459);
or U19276 (N_19276,N_17852,N_17664);
or U19277 (N_19277,N_16747,N_17914);
or U19278 (N_19278,N_17734,N_17239);
xnor U19279 (N_19279,N_16356,N_16951);
nor U19280 (N_19280,N_17010,N_16531);
or U19281 (N_19281,N_16068,N_17334);
and U19282 (N_19282,N_16728,N_17823);
nand U19283 (N_19283,N_17838,N_16643);
or U19284 (N_19284,N_17256,N_17481);
or U19285 (N_19285,N_16105,N_16315);
and U19286 (N_19286,N_17530,N_17352);
and U19287 (N_19287,N_16584,N_17625);
and U19288 (N_19288,N_16473,N_17484);
nand U19289 (N_19289,N_16147,N_16886);
nand U19290 (N_19290,N_16141,N_16635);
or U19291 (N_19291,N_16315,N_17589);
or U19292 (N_19292,N_16524,N_17532);
xnor U19293 (N_19293,N_16796,N_16262);
and U19294 (N_19294,N_17613,N_16575);
xor U19295 (N_19295,N_17813,N_17068);
nand U19296 (N_19296,N_17576,N_17160);
nand U19297 (N_19297,N_17839,N_16750);
or U19298 (N_19298,N_17785,N_17968);
xnor U19299 (N_19299,N_16549,N_17373);
nor U19300 (N_19300,N_17091,N_16185);
or U19301 (N_19301,N_17783,N_16438);
nor U19302 (N_19302,N_16616,N_16506);
xor U19303 (N_19303,N_17220,N_16243);
and U19304 (N_19304,N_17053,N_17373);
nand U19305 (N_19305,N_17157,N_17067);
or U19306 (N_19306,N_16385,N_16633);
or U19307 (N_19307,N_16844,N_16172);
xnor U19308 (N_19308,N_16191,N_16824);
nand U19309 (N_19309,N_17092,N_16260);
or U19310 (N_19310,N_17773,N_16601);
nand U19311 (N_19311,N_16965,N_17752);
nor U19312 (N_19312,N_16772,N_17496);
xnor U19313 (N_19313,N_17391,N_16878);
nor U19314 (N_19314,N_16447,N_16880);
nand U19315 (N_19315,N_16555,N_16814);
and U19316 (N_19316,N_17058,N_16495);
nand U19317 (N_19317,N_16276,N_17190);
or U19318 (N_19318,N_17145,N_16196);
and U19319 (N_19319,N_17217,N_16991);
or U19320 (N_19320,N_16780,N_16540);
or U19321 (N_19321,N_17112,N_16246);
xnor U19322 (N_19322,N_17350,N_16167);
nor U19323 (N_19323,N_16601,N_16017);
and U19324 (N_19324,N_16650,N_16975);
or U19325 (N_19325,N_16499,N_16643);
and U19326 (N_19326,N_16530,N_17279);
and U19327 (N_19327,N_16564,N_16900);
or U19328 (N_19328,N_17864,N_16108);
or U19329 (N_19329,N_17316,N_16869);
and U19330 (N_19330,N_16870,N_16880);
and U19331 (N_19331,N_17076,N_16930);
xor U19332 (N_19332,N_16448,N_16494);
nand U19333 (N_19333,N_16401,N_17144);
xor U19334 (N_19334,N_17980,N_17402);
and U19335 (N_19335,N_16935,N_17621);
xnor U19336 (N_19336,N_17001,N_17244);
nand U19337 (N_19337,N_16408,N_16523);
nand U19338 (N_19338,N_16656,N_17993);
nand U19339 (N_19339,N_17890,N_16317);
nand U19340 (N_19340,N_17294,N_16071);
and U19341 (N_19341,N_17322,N_16375);
or U19342 (N_19342,N_17250,N_17120);
nor U19343 (N_19343,N_17709,N_16368);
or U19344 (N_19344,N_17967,N_17792);
and U19345 (N_19345,N_17647,N_17392);
or U19346 (N_19346,N_17526,N_16343);
xor U19347 (N_19347,N_16600,N_17998);
and U19348 (N_19348,N_17653,N_17828);
nand U19349 (N_19349,N_16264,N_16503);
or U19350 (N_19350,N_17473,N_17355);
nand U19351 (N_19351,N_16827,N_17640);
xnor U19352 (N_19352,N_16790,N_16123);
nand U19353 (N_19353,N_17214,N_17697);
nand U19354 (N_19354,N_17844,N_16718);
nand U19355 (N_19355,N_16974,N_16240);
or U19356 (N_19356,N_17508,N_16621);
or U19357 (N_19357,N_17620,N_17442);
nand U19358 (N_19358,N_16484,N_17092);
nand U19359 (N_19359,N_16892,N_16809);
or U19360 (N_19360,N_17100,N_17594);
and U19361 (N_19361,N_16558,N_17028);
and U19362 (N_19362,N_16040,N_17893);
and U19363 (N_19363,N_16121,N_16567);
xor U19364 (N_19364,N_16519,N_17468);
nand U19365 (N_19365,N_17407,N_16923);
and U19366 (N_19366,N_16106,N_17090);
nand U19367 (N_19367,N_16034,N_16785);
nand U19368 (N_19368,N_16007,N_16010);
or U19369 (N_19369,N_17644,N_17074);
nand U19370 (N_19370,N_17538,N_17529);
xor U19371 (N_19371,N_16573,N_16853);
xor U19372 (N_19372,N_17893,N_17398);
nand U19373 (N_19373,N_16552,N_17835);
and U19374 (N_19374,N_16349,N_16234);
nor U19375 (N_19375,N_17046,N_16486);
and U19376 (N_19376,N_17127,N_16575);
or U19377 (N_19377,N_17154,N_17731);
and U19378 (N_19378,N_16954,N_16781);
xor U19379 (N_19379,N_16895,N_16322);
or U19380 (N_19380,N_17931,N_17488);
nor U19381 (N_19381,N_17148,N_17402);
nor U19382 (N_19382,N_17726,N_16171);
nor U19383 (N_19383,N_17923,N_16149);
and U19384 (N_19384,N_16184,N_17613);
xnor U19385 (N_19385,N_17072,N_16365);
and U19386 (N_19386,N_17219,N_16551);
and U19387 (N_19387,N_16396,N_17260);
and U19388 (N_19388,N_17217,N_17033);
xnor U19389 (N_19389,N_16931,N_16799);
nand U19390 (N_19390,N_16135,N_17095);
and U19391 (N_19391,N_16937,N_17018);
nor U19392 (N_19392,N_17781,N_17220);
and U19393 (N_19393,N_16371,N_16873);
nor U19394 (N_19394,N_16087,N_17711);
xnor U19395 (N_19395,N_16340,N_16420);
nand U19396 (N_19396,N_16147,N_16383);
and U19397 (N_19397,N_17357,N_16056);
and U19398 (N_19398,N_16350,N_17712);
or U19399 (N_19399,N_17531,N_17891);
nand U19400 (N_19400,N_17457,N_16456);
xor U19401 (N_19401,N_17293,N_16841);
and U19402 (N_19402,N_17977,N_17510);
nand U19403 (N_19403,N_17232,N_17594);
nand U19404 (N_19404,N_17248,N_16712);
xor U19405 (N_19405,N_16555,N_17004);
xnor U19406 (N_19406,N_17136,N_16089);
nor U19407 (N_19407,N_17022,N_17499);
or U19408 (N_19408,N_16129,N_16754);
nand U19409 (N_19409,N_17387,N_17354);
xnor U19410 (N_19410,N_16722,N_17023);
xor U19411 (N_19411,N_17569,N_16936);
nand U19412 (N_19412,N_16932,N_16300);
and U19413 (N_19413,N_16481,N_17455);
or U19414 (N_19414,N_16781,N_16339);
nand U19415 (N_19415,N_16198,N_16449);
xnor U19416 (N_19416,N_17043,N_17243);
nor U19417 (N_19417,N_16945,N_17534);
nor U19418 (N_19418,N_17199,N_16774);
and U19419 (N_19419,N_17836,N_17848);
xnor U19420 (N_19420,N_17043,N_16558);
xnor U19421 (N_19421,N_17343,N_16091);
and U19422 (N_19422,N_17100,N_17374);
xor U19423 (N_19423,N_16690,N_17564);
or U19424 (N_19424,N_16383,N_16385);
xor U19425 (N_19425,N_16011,N_16196);
xnor U19426 (N_19426,N_17686,N_17334);
xnor U19427 (N_19427,N_17853,N_16709);
nand U19428 (N_19428,N_16820,N_17718);
nor U19429 (N_19429,N_16583,N_17934);
and U19430 (N_19430,N_17514,N_17058);
xor U19431 (N_19431,N_16350,N_17420);
nor U19432 (N_19432,N_16244,N_16810);
or U19433 (N_19433,N_17608,N_17255);
nor U19434 (N_19434,N_16055,N_16011);
nor U19435 (N_19435,N_16343,N_16358);
xnor U19436 (N_19436,N_16054,N_16924);
nor U19437 (N_19437,N_16419,N_17094);
and U19438 (N_19438,N_17277,N_16269);
xnor U19439 (N_19439,N_16462,N_16729);
nand U19440 (N_19440,N_17971,N_16804);
nor U19441 (N_19441,N_17343,N_17209);
xnor U19442 (N_19442,N_17620,N_16252);
xnor U19443 (N_19443,N_17617,N_17767);
or U19444 (N_19444,N_16016,N_16955);
or U19445 (N_19445,N_16065,N_17857);
and U19446 (N_19446,N_16475,N_17325);
or U19447 (N_19447,N_16068,N_16233);
nand U19448 (N_19448,N_16448,N_16768);
nand U19449 (N_19449,N_16394,N_17727);
xor U19450 (N_19450,N_16651,N_17823);
nand U19451 (N_19451,N_16413,N_16024);
or U19452 (N_19452,N_17131,N_17786);
nand U19453 (N_19453,N_16381,N_17840);
nor U19454 (N_19454,N_17492,N_16092);
xor U19455 (N_19455,N_17190,N_16163);
or U19456 (N_19456,N_16178,N_17888);
nor U19457 (N_19457,N_16614,N_16540);
nand U19458 (N_19458,N_17118,N_16701);
or U19459 (N_19459,N_16624,N_17621);
nor U19460 (N_19460,N_16506,N_17967);
or U19461 (N_19461,N_16269,N_16757);
xor U19462 (N_19462,N_17101,N_17731);
nand U19463 (N_19463,N_17714,N_16550);
xnor U19464 (N_19464,N_16839,N_16671);
or U19465 (N_19465,N_16362,N_16002);
nor U19466 (N_19466,N_16487,N_17042);
nor U19467 (N_19467,N_16073,N_17306);
nor U19468 (N_19468,N_17034,N_16808);
nand U19469 (N_19469,N_17800,N_16709);
and U19470 (N_19470,N_16311,N_16489);
nand U19471 (N_19471,N_17743,N_16865);
xor U19472 (N_19472,N_17758,N_16843);
xnor U19473 (N_19473,N_17622,N_16644);
nor U19474 (N_19474,N_17327,N_16332);
and U19475 (N_19475,N_16282,N_17207);
nand U19476 (N_19476,N_17732,N_16011);
nor U19477 (N_19477,N_16195,N_17546);
and U19478 (N_19478,N_17933,N_17308);
or U19479 (N_19479,N_17282,N_17834);
xor U19480 (N_19480,N_16558,N_17370);
nand U19481 (N_19481,N_16678,N_17796);
xnor U19482 (N_19482,N_17087,N_16880);
xnor U19483 (N_19483,N_17132,N_16525);
and U19484 (N_19484,N_16004,N_16769);
nor U19485 (N_19485,N_17477,N_16567);
nand U19486 (N_19486,N_16166,N_16734);
and U19487 (N_19487,N_16726,N_17977);
xnor U19488 (N_19488,N_16430,N_16631);
nor U19489 (N_19489,N_17145,N_16933);
xnor U19490 (N_19490,N_16890,N_17857);
or U19491 (N_19491,N_17320,N_16151);
and U19492 (N_19492,N_16039,N_16564);
nor U19493 (N_19493,N_17613,N_16176);
xor U19494 (N_19494,N_17874,N_16938);
xnor U19495 (N_19495,N_16390,N_17844);
or U19496 (N_19496,N_16607,N_17608);
nor U19497 (N_19497,N_16729,N_16364);
xnor U19498 (N_19498,N_17752,N_16053);
and U19499 (N_19499,N_16906,N_16100);
xor U19500 (N_19500,N_16810,N_17723);
xnor U19501 (N_19501,N_16891,N_16986);
or U19502 (N_19502,N_17147,N_16897);
xor U19503 (N_19503,N_16307,N_17640);
xor U19504 (N_19504,N_17901,N_17428);
nor U19505 (N_19505,N_16350,N_16281);
xnor U19506 (N_19506,N_16157,N_17490);
nand U19507 (N_19507,N_16214,N_16719);
or U19508 (N_19508,N_16612,N_16130);
nand U19509 (N_19509,N_17063,N_16831);
or U19510 (N_19510,N_16228,N_16527);
and U19511 (N_19511,N_17024,N_17757);
nand U19512 (N_19512,N_16893,N_17686);
nor U19513 (N_19513,N_17930,N_16289);
or U19514 (N_19514,N_17103,N_17874);
and U19515 (N_19515,N_17232,N_17715);
nor U19516 (N_19516,N_17924,N_17222);
nand U19517 (N_19517,N_16058,N_17755);
nor U19518 (N_19518,N_16689,N_16621);
nand U19519 (N_19519,N_16016,N_16353);
and U19520 (N_19520,N_16567,N_16749);
and U19521 (N_19521,N_16617,N_17538);
nor U19522 (N_19522,N_16053,N_16693);
nor U19523 (N_19523,N_16166,N_17299);
xnor U19524 (N_19524,N_17906,N_16902);
or U19525 (N_19525,N_17573,N_16991);
nor U19526 (N_19526,N_16468,N_16300);
and U19527 (N_19527,N_16704,N_16866);
nand U19528 (N_19528,N_17081,N_17433);
nor U19529 (N_19529,N_16676,N_16035);
or U19530 (N_19530,N_16760,N_17110);
nand U19531 (N_19531,N_16555,N_16785);
and U19532 (N_19532,N_17310,N_16665);
nor U19533 (N_19533,N_17090,N_17993);
or U19534 (N_19534,N_16589,N_17841);
xnor U19535 (N_19535,N_16248,N_16924);
nor U19536 (N_19536,N_16511,N_16281);
nand U19537 (N_19537,N_16706,N_17617);
or U19538 (N_19538,N_16487,N_16588);
or U19539 (N_19539,N_16980,N_17343);
nor U19540 (N_19540,N_17355,N_17339);
nor U19541 (N_19541,N_17657,N_16218);
nand U19542 (N_19542,N_16497,N_16515);
xor U19543 (N_19543,N_16294,N_17780);
nand U19544 (N_19544,N_16989,N_17367);
or U19545 (N_19545,N_16236,N_16073);
nor U19546 (N_19546,N_16858,N_17779);
nand U19547 (N_19547,N_17273,N_16450);
nor U19548 (N_19548,N_16609,N_16714);
nand U19549 (N_19549,N_16462,N_16489);
nor U19550 (N_19550,N_17222,N_17212);
nor U19551 (N_19551,N_17578,N_17742);
and U19552 (N_19552,N_16721,N_16129);
nor U19553 (N_19553,N_17629,N_17497);
nor U19554 (N_19554,N_17505,N_16747);
or U19555 (N_19555,N_17849,N_16284);
xnor U19556 (N_19556,N_16728,N_17103);
nor U19557 (N_19557,N_17223,N_17950);
nor U19558 (N_19558,N_16645,N_17517);
or U19559 (N_19559,N_16120,N_16736);
nand U19560 (N_19560,N_16166,N_17707);
and U19561 (N_19561,N_16924,N_17445);
and U19562 (N_19562,N_16519,N_16524);
xor U19563 (N_19563,N_17958,N_16312);
nand U19564 (N_19564,N_16386,N_17946);
and U19565 (N_19565,N_16147,N_17155);
and U19566 (N_19566,N_17957,N_16249);
or U19567 (N_19567,N_16726,N_16904);
xor U19568 (N_19568,N_16509,N_17356);
xnor U19569 (N_19569,N_16341,N_17466);
nand U19570 (N_19570,N_16681,N_16950);
nor U19571 (N_19571,N_17043,N_16704);
or U19572 (N_19572,N_17790,N_16011);
nand U19573 (N_19573,N_16324,N_16833);
xor U19574 (N_19574,N_17944,N_17252);
nor U19575 (N_19575,N_17042,N_17276);
and U19576 (N_19576,N_17118,N_16395);
and U19577 (N_19577,N_17604,N_16001);
nand U19578 (N_19578,N_16146,N_16124);
and U19579 (N_19579,N_17973,N_16510);
or U19580 (N_19580,N_16654,N_17806);
nor U19581 (N_19581,N_16431,N_16610);
nor U19582 (N_19582,N_16552,N_16901);
nor U19583 (N_19583,N_16553,N_17166);
or U19584 (N_19584,N_17831,N_16002);
or U19585 (N_19585,N_16723,N_17153);
xnor U19586 (N_19586,N_16213,N_17461);
and U19587 (N_19587,N_16537,N_16880);
nor U19588 (N_19588,N_17936,N_17659);
xnor U19589 (N_19589,N_17692,N_16048);
or U19590 (N_19590,N_17016,N_17941);
xor U19591 (N_19591,N_17604,N_16090);
and U19592 (N_19592,N_16801,N_17672);
xnor U19593 (N_19593,N_17273,N_17015);
nand U19594 (N_19594,N_16274,N_16446);
nand U19595 (N_19595,N_16369,N_16153);
xor U19596 (N_19596,N_16239,N_16015);
nand U19597 (N_19597,N_17904,N_17607);
or U19598 (N_19598,N_16647,N_17655);
xor U19599 (N_19599,N_17807,N_16636);
nor U19600 (N_19600,N_16839,N_17686);
and U19601 (N_19601,N_17990,N_16668);
xor U19602 (N_19602,N_17359,N_16225);
xnor U19603 (N_19603,N_16655,N_17035);
nand U19604 (N_19604,N_17302,N_17702);
nand U19605 (N_19605,N_17054,N_17082);
and U19606 (N_19606,N_16888,N_16346);
xnor U19607 (N_19607,N_17601,N_16842);
nor U19608 (N_19608,N_16110,N_16720);
nand U19609 (N_19609,N_17204,N_16246);
or U19610 (N_19610,N_17490,N_16922);
and U19611 (N_19611,N_17441,N_16311);
xor U19612 (N_19612,N_17742,N_16798);
or U19613 (N_19613,N_17372,N_17660);
xnor U19614 (N_19614,N_17269,N_16403);
nand U19615 (N_19615,N_16651,N_17100);
and U19616 (N_19616,N_17220,N_17577);
xnor U19617 (N_19617,N_16250,N_17670);
and U19618 (N_19618,N_16789,N_17033);
and U19619 (N_19619,N_17461,N_17860);
and U19620 (N_19620,N_16111,N_17867);
or U19621 (N_19621,N_17725,N_17121);
nor U19622 (N_19622,N_17186,N_16201);
xor U19623 (N_19623,N_17740,N_17157);
xor U19624 (N_19624,N_16705,N_17200);
xnor U19625 (N_19625,N_17350,N_17399);
xnor U19626 (N_19626,N_16454,N_16438);
xor U19627 (N_19627,N_16324,N_17155);
or U19628 (N_19628,N_17954,N_16336);
and U19629 (N_19629,N_16392,N_17160);
xor U19630 (N_19630,N_17840,N_16440);
xor U19631 (N_19631,N_16934,N_16338);
nand U19632 (N_19632,N_17786,N_17764);
and U19633 (N_19633,N_17966,N_16207);
nand U19634 (N_19634,N_17940,N_16627);
nand U19635 (N_19635,N_17260,N_16092);
nor U19636 (N_19636,N_16629,N_17492);
nand U19637 (N_19637,N_17111,N_17993);
nor U19638 (N_19638,N_17723,N_17979);
nand U19639 (N_19639,N_17993,N_17822);
or U19640 (N_19640,N_17756,N_16380);
xor U19641 (N_19641,N_16359,N_17373);
and U19642 (N_19642,N_17311,N_16706);
nand U19643 (N_19643,N_17300,N_16800);
nand U19644 (N_19644,N_16239,N_17205);
or U19645 (N_19645,N_16627,N_17755);
nand U19646 (N_19646,N_16749,N_16279);
and U19647 (N_19647,N_17647,N_17646);
xor U19648 (N_19648,N_17601,N_16655);
nor U19649 (N_19649,N_16358,N_17249);
nor U19650 (N_19650,N_17073,N_17370);
nor U19651 (N_19651,N_17521,N_17298);
nand U19652 (N_19652,N_17049,N_17271);
xnor U19653 (N_19653,N_17251,N_17594);
xor U19654 (N_19654,N_17978,N_17509);
or U19655 (N_19655,N_16791,N_17255);
nand U19656 (N_19656,N_17826,N_17653);
nor U19657 (N_19657,N_16302,N_17939);
xnor U19658 (N_19658,N_16918,N_16230);
nor U19659 (N_19659,N_17710,N_17869);
nor U19660 (N_19660,N_16101,N_17487);
nor U19661 (N_19661,N_16849,N_17731);
nand U19662 (N_19662,N_16580,N_16041);
nand U19663 (N_19663,N_17883,N_17449);
or U19664 (N_19664,N_16150,N_17722);
nand U19665 (N_19665,N_17862,N_17701);
nand U19666 (N_19666,N_16639,N_17948);
xnor U19667 (N_19667,N_16692,N_17948);
nand U19668 (N_19668,N_16335,N_16457);
or U19669 (N_19669,N_17249,N_16572);
nand U19670 (N_19670,N_17835,N_17485);
xnor U19671 (N_19671,N_16043,N_16624);
and U19672 (N_19672,N_17174,N_17640);
or U19673 (N_19673,N_16511,N_17820);
nor U19674 (N_19674,N_17277,N_17768);
xnor U19675 (N_19675,N_16037,N_17748);
and U19676 (N_19676,N_17682,N_16382);
xnor U19677 (N_19677,N_17339,N_17595);
xnor U19678 (N_19678,N_17149,N_17900);
nand U19679 (N_19679,N_16155,N_17513);
nand U19680 (N_19680,N_16415,N_17830);
nor U19681 (N_19681,N_17627,N_16404);
xnor U19682 (N_19682,N_16024,N_17470);
and U19683 (N_19683,N_16494,N_17654);
xnor U19684 (N_19684,N_17207,N_16295);
nand U19685 (N_19685,N_17584,N_17266);
and U19686 (N_19686,N_17584,N_17134);
and U19687 (N_19687,N_17421,N_16786);
or U19688 (N_19688,N_17532,N_16712);
xnor U19689 (N_19689,N_17663,N_17275);
and U19690 (N_19690,N_16887,N_16660);
nor U19691 (N_19691,N_16149,N_17552);
or U19692 (N_19692,N_17411,N_16330);
nand U19693 (N_19693,N_16580,N_17012);
nor U19694 (N_19694,N_16038,N_17339);
or U19695 (N_19695,N_16013,N_17353);
nand U19696 (N_19696,N_16399,N_16746);
nand U19697 (N_19697,N_16015,N_16683);
nor U19698 (N_19698,N_17077,N_16624);
nand U19699 (N_19699,N_16283,N_16048);
and U19700 (N_19700,N_17735,N_16887);
or U19701 (N_19701,N_16263,N_17788);
nor U19702 (N_19702,N_16134,N_16957);
nand U19703 (N_19703,N_17071,N_16509);
nand U19704 (N_19704,N_17637,N_17233);
nand U19705 (N_19705,N_16714,N_16981);
or U19706 (N_19706,N_17281,N_16106);
or U19707 (N_19707,N_17607,N_17654);
xor U19708 (N_19708,N_16956,N_16603);
and U19709 (N_19709,N_16374,N_17273);
nor U19710 (N_19710,N_16030,N_16010);
nor U19711 (N_19711,N_17909,N_16998);
nand U19712 (N_19712,N_16751,N_16534);
or U19713 (N_19713,N_16273,N_17685);
or U19714 (N_19714,N_16914,N_17583);
nand U19715 (N_19715,N_17000,N_16344);
nor U19716 (N_19716,N_17978,N_16352);
and U19717 (N_19717,N_16092,N_16584);
and U19718 (N_19718,N_17988,N_17721);
xnor U19719 (N_19719,N_16215,N_16126);
nor U19720 (N_19720,N_17255,N_17390);
xor U19721 (N_19721,N_17256,N_17764);
and U19722 (N_19722,N_16552,N_16645);
xor U19723 (N_19723,N_16776,N_17924);
xor U19724 (N_19724,N_16427,N_17180);
and U19725 (N_19725,N_17599,N_17864);
nand U19726 (N_19726,N_16995,N_16195);
nor U19727 (N_19727,N_16946,N_17115);
or U19728 (N_19728,N_16832,N_16671);
or U19729 (N_19729,N_17733,N_16646);
or U19730 (N_19730,N_17338,N_17445);
or U19731 (N_19731,N_17618,N_17978);
and U19732 (N_19732,N_16733,N_16037);
or U19733 (N_19733,N_17406,N_16396);
nor U19734 (N_19734,N_17442,N_16664);
or U19735 (N_19735,N_16922,N_16973);
and U19736 (N_19736,N_16846,N_17898);
and U19737 (N_19737,N_17417,N_16882);
nand U19738 (N_19738,N_16317,N_17611);
and U19739 (N_19739,N_16667,N_16612);
nand U19740 (N_19740,N_16788,N_17212);
nor U19741 (N_19741,N_17321,N_17283);
xor U19742 (N_19742,N_16838,N_17483);
and U19743 (N_19743,N_17436,N_16431);
and U19744 (N_19744,N_17945,N_17830);
and U19745 (N_19745,N_16674,N_16724);
nor U19746 (N_19746,N_16759,N_17148);
nand U19747 (N_19747,N_17217,N_16343);
xnor U19748 (N_19748,N_16880,N_16022);
and U19749 (N_19749,N_17954,N_17882);
xnor U19750 (N_19750,N_17511,N_17907);
xor U19751 (N_19751,N_16284,N_17471);
or U19752 (N_19752,N_16730,N_17634);
nand U19753 (N_19753,N_17125,N_16054);
or U19754 (N_19754,N_17689,N_16965);
nand U19755 (N_19755,N_17070,N_16824);
nand U19756 (N_19756,N_17094,N_16501);
nand U19757 (N_19757,N_16793,N_16911);
or U19758 (N_19758,N_16392,N_17737);
nor U19759 (N_19759,N_16407,N_17596);
or U19760 (N_19760,N_16648,N_16108);
or U19761 (N_19761,N_16900,N_17948);
nand U19762 (N_19762,N_16769,N_17207);
nor U19763 (N_19763,N_17417,N_16871);
and U19764 (N_19764,N_16937,N_17826);
or U19765 (N_19765,N_17814,N_16057);
and U19766 (N_19766,N_17149,N_17053);
nand U19767 (N_19767,N_16876,N_17238);
or U19768 (N_19768,N_16485,N_16178);
and U19769 (N_19769,N_16186,N_16413);
and U19770 (N_19770,N_16884,N_17248);
or U19771 (N_19771,N_17578,N_16248);
nor U19772 (N_19772,N_17077,N_17525);
or U19773 (N_19773,N_16204,N_17106);
or U19774 (N_19774,N_16226,N_16914);
or U19775 (N_19775,N_16150,N_16311);
nor U19776 (N_19776,N_16300,N_16306);
nand U19777 (N_19777,N_16793,N_16609);
and U19778 (N_19778,N_16452,N_16145);
and U19779 (N_19779,N_16206,N_17855);
xor U19780 (N_19780,N_16196,N_17757);
xor U19781 (N_19781,N_17482,N_16954);
nor U19782 (N_19782,N_16852,N_16672);
xor U19783 (N_19783,N_16688,N_17443);
or U19784 (N_19784,N_16135,N_17751);
and U19785 (N_19785,N_17213,N_17865);
nor U19786 (N_19786,N_17408,N_17089);
and U19787 (N_19787,N_17709,N_17123);
xnor U19788 (N_19788,N_16138,N_16784);
or U19789 (N_19789,N_17303,N_16310);
nand U19790 (N_19790,N_17836,N_17498);
or U19791 (N_19791,N_16566,N_16421);
and U19792 (N_19792,N_16218,N_16801);
xnor U19793 (N_19793,N_17576,N_17195);
and U19794 (N_19794,N_16543,N_16615);
nand U19795 (N_19795,N_17744,N_16989);
nor U19796 (N_19796,N_17396,N_17478);
or U19797 (N_19797,N_16104,N_17990);
or U19798 (N_19798,N_16956,N_17563);
nor U19799 (N_19799,N_16144,N_17712);
or U19800 (N_19800,N_16682,N_16908);
or U19801 (N_19801,N_17709,N_16297);
xnor U19802 (N_19802,N_17953,N_16542);
nor U19803 (N_19803,N_17389,N_16114);
and U19804 (N_19804,N_17180,N_17487);
nand U19805 (N_19805,N_17732,N_17892);
xor U19806 (N_19806,N_17739,N_16443);
xnor U19807 (N_19807,N_16287,N_16558);
xor U19808 (N_19808,N_16283,N_16474);
nor U19809 (N_19809,N_16528,N_17242);
or U19810 (N_19810,N_16394,N_16025);
and U19811 (N_19811,N_17501,N_17835);
nand U19812 (N_19812,N_17180,N_16335);
or U19813 (N_19813,N_16966,N_16426);
and U19814 (N_19814,N_16338,N_17016);
or U19815 (N_19815,N_16221,N_17530);
xor U19816 (N_19816,N_17008,N_16876);
and U19817 (N_19817,N_16790,N_16891);
nor U19818 (N_19818,N_17861,N_16187);
xnor U19819 (N_19819,N_16743,N_17722);
and U19820 (N_19820,N_17645,N_17994);
nand U19821 (N_19821,N_17150,N_16444);
or U19822 (N_19822,N_16488,N_17595);
nand U19823 (N_19823,N_17771,N_16086);
and U19824 (N_19824,N_16365,N_17581);
nor U19825 (N_19825,N_16443,N_16622);
nor U19826 (N_19826,N_16836,N_16311);
or U19827 (N_19827,N_17567,N_17487);
nor U19828 (N_19828,N_17462,N_16771);
nand U19829 (N_19829,N_17249,N_17319);
and U19830 (N_19830,N_16371,N_17849);
nor U19831 (N_19831,N_17771,N_17011);
xor U19832 (N_19832,N_17020,N_17740);
or U19833 (N_19833,N_17899,N_16088);
xor U19834 (N_19834,N_16310,N_16525);
or U19835 (N_19835,N_17931,N_16430);
or U19836 (N_19836,N_16249,N_17323);
and U19837 (N_19837,N_17078,N_16540);
or U19838 (N_19838,N_17737,N_17703);
or U19839 (N_19839,N_17010,N_16375);
nor U19840 (N_19840,N_17027,N_16259);
and U19841 (N_19841,N_17239,N_17849);
nand U19842 (N_19842,N_17204,N_17079);
nand U19843 (N_19843,N_17373,N_17934);
and U19844 (N_19844,N_17940,N_16093);
nor U19845 (N_19845,N_16026,N_17945);
xnor U19846 (N_19846,N_16631,N_16573);
nor U19847 (N_19847,N_16457,N_16390);
nand U19848 (N_19848,N_17922,N_16709);
and U19849 (N_19849,N_16499,N_17905);
and U19850 (N_19850,N_17228,N_17345);
nor U19851 (N_19851,N_16886,N_17854);
or U19852 (N_19852,N_17704,N_17007);
or U19853 (N_19853,N_16135,N_17765);
nand U19854 (N_19854,N_16167,N_17721);
and U19855 (N_19855,N_16382,N_16359);
xor U19856 (N_19856,N_17576,N_17435);
or U19857 (N_19857,N_16072,N_17495);
xor U19858 (N_19858,N_17063,N_16254);
or U19859 (N_19859,N_16835,N_17097);
or U19860 (N_19860,N_16222,N_16901);
nand U19861 (N_19861,N_17167,N_16162);
nand U19862 (N_19862,N_17781,N_16066);
xnor U19863 (N_19863,N_16729,N_16618);
and U19864 (N_19864,N_17052,N_16912);
or U19865 (N_19865,N_17451,N_16017);
or U19866 (N_19866,N_17716,N_17432);
nand U19867 (N_19867,N_16943,N_16302);
xor U19868 (N_19868,N_16694,N_17479);
nor U19869 (N_19869,N_17280,N_17581);
or U19870 (N_19870,N_16781,N_17989);
or U19871 (N_19871,N_16951,N_17545);
nand U19872 (N_19872,N_16282,N_16509);
nor U19873 (N_19873,N_16145,N_17740);
nand U19874 (N_19874,N_16967,N_16291);
nor U19875 (N_19875,N_16596,N_17130);
nand U19876 (N_19876,N_17532,N_17869);
nand U19877 (N_19877,N_17175,N_17527);
xor U19878 (N_19878,N_16864,N_16377);
nor U19879 (N_19879,N_17607,N_17052);
or U19880 (N_19880,N_17481,N_17885);
or U19881 (N_19881,N_17216,N_16517);
nor U19882 (N_19882,N_16410,N_16377);
nand U19883 (N_19883,N_17894,N_16526);
or U19884 (N_19884,N_17979,N_17293);
nand U19885 (N_19885,N_16423,N_16266);
or U19886 (N_19886,N_17128,N_17306);
nor U19887 (N_19887,N_16599,N_16329);
and U19888 (N_19888,N_17122,N_16255);
xnor U19889 (N_19889,N_17357,N_16486);
and U19890 (N_19890,N_16612,N_17792);
nand U19891 (N_19891,N_16261,N_16804);
or U19892 (N_19892,N_17453,N_16595);
xor U19893 (N_19893,N_16405,N_17368);
nand U19894 (N_19894,N_16812,N_17215);
nand U19895 (N_19895,N_16469,N_16471);
nand U19896 (N_19896,N_17445,N_16671);
and U19897 (N_19897,N_17031,N_16800);
nand U19898 (N_19898,N_17446,N_16081);
xor U19899 (N_19899,N_16997,N_17325);
nor U19900 (N_19900,N_16344,N_16463);
and U19901 (N_19901,N_17881,N_17555);
xnor U19902 (N_19902,N_17776,N_16685);
and U19903 (N_19903,N_17102,N_16027);
and U19904 (N_19904,N_16392,N_17563);
nor U19905 (N_19905,N_17506,N_17693);
nor U19906 (N_19906,N_17579,N_17416);
or U19907 (N_19907,N_16121,N_17139);
or U19908 (N_19908,N_16426,N_16256);
and U19909 (N_19909,N_16724,N_16259);
xnor U19910 (N_19910,N_16501,N_17243);
nand U19911 (N_19911,N_16597,N_17241);
xnor U19912 (N_19912,N_17368,N_16074);
and U19913 (N_19913,N_17567,N_17387);
nand U19914 (N_19914,N_16113,N_17132);
xor U19915 (N_19915,N_16849,N_17650);
and U19916 (N_19916,N_16866,N_16571);
or U19917 (N_19917,N_17753,N_16103);
nand U19918 (N_19918,N_17382,N_16876);
or U19919 (N_19919,N_17321,N_16589);
xor U19920 (N_19920,N_16407,N_16948);
and U19921 (N_19921,N_17774,N_16398);
or U19922 (N_19922,N_17144,N_17290);
or U19923 (N_19923,N_16215,N_16360);
nand U19924 (N_19924,N_17159,N_16318);
and U19925 (N_19925,N_17403,N_16513);
or U19926 (N_19926,N_16477,N_16099);
nand U19927 (N_19927,N_16264,N_16100);
nor U19928 (N_19928,N_16023,N_16316);
nor U19929 (N_19929,N_17232,N_16330);
nand U19930 (N_19930,N_16521,N_16676);
nor U19931 (N_19931,N_16851,N_17665);
nor U19932 (N_19932,N_16923,N_17025);
nor U19933 (N_19933,N_16919,N_16960);
and U19934 (N_19934,N_16587,N_16760);
nand U19935 (N_19935,N_17507,N_16235);
or U19936 (N_19936,N_17844,N_17886);
or U19937 (N_19937,N_17969,N_16598);
nand U19938 (N_19938,N_17942,N_17523);
nand U19939 (N_19939,N_16171,N_17516);
xnor U19940 (N_19940,N_16740,N_17993);
or U19941 (N_19941,N_17751,N_17560);
xor U19942 (N_19942,N_17196,N_16944);
or U19943 (N_19943,N_17279,N_17072);
nand U19944 (N_19944,N_17573,N_17941);
nand U19945 (N_19945,N_16444,N_16360);
nor U19946 (N_19946,N_16666,N_17075);
or U19947 (N_19947,N_17928,N_17002);
nand U19948 (N_19948,N_17835,N_16661);
nand U19949 (N_19949,N_16377,N_16888);
nand U19950 (N_19950,N_16552,N_16077);
or U19951 (N_19951,N_17766,N_16322);
xor U19952 (N_19952,N_17220,N_16195);
nor U19953 (N_19953,N_16570,N_17612);
and U19954 (N_19954,N_16678,N_17579);
nand U19955 (N_19955,N_16221,N_16601);
nand U19956 (N_19956,N_17873,N_16506);
and U19957 (N_19957,N_16393,N_17615);
xnor U19958 (N_19958,N_17789,N_17492);
xor U19959 (N_19959,N_17952,N_16039);
nand U19960 (N_19960,N_17930,N_17577);
and U19961 (N_19961,N_17317,N_16181);
and U19962 (N_19962,N_16174,N_17487);
and U19963 (N_19963,N_16717,N_16223);
xnor U19964 (N_19964,N_17629,N_17365);
nand U19965 (N_19965,N_16147,N_16270);
nand U19966 (N_19966,N_17483,N_16752);
or U19967 (N_19967,N_16595,N_16860);
xnor U19968 (N_19968,N_16481,N_17429);
or U19969 (N_19969,N_17614,N_16186);
xnor U19970 (N_19970,N_16555,N_16983);
nor U19971 (N_19971,N_17051,N_16563);
nor U19972 (N_19972,N_17550,N_16458);
and U19973 (N_19973,N_17356,N_17308);
and U19974 (N_19974,N_17051,N_17532);
nor U19975 (N_19975,N_17580,N_16127);
xnor U19976 (N_19976,N_16395,N_16656);
and U19977 (N_19977,N_17913,N_17293);
nand U19978 (N_19978,N_16599,N_17372);
or U19979 (N_19979,N_17715,N_17117);
nor U19980 (N_19980,N_17239,N_16861);
and U19981 (N_19981,N_17297,N_17001);
xor U19982 (N_19982,N_17365,N_17856);
nor U19983 (N_19983,N_17198,N_16372);
xor U19984 (N_19984,N_16951,N_17593);
xor U19985 (N_19985,N_17466,N_16604);
xnor U19986 (N_19986,N_16484,N_16491);
nand U19987 (N_19987,N_16321,N_17090);
and U19988 (N_19988,N_17067,N_16902);
and U19989 (N_19989,N_16073,N_17925);
xor U19990 (N_19990,N_16386,N_17008);
nand U19991 (N_19991,N_16976,N_16776);
xnor U19992 (N_19992,N_17858,N_16034);
and U19993 (N_19993,N_17652,N_16327);
nand U19994 (N_19994,N_16443,N_16874);
nor U19995 (N_19995,N_16071,N_17286);
or U19996 (N_19996,N_17870,N_17461);
nor U19997 (N_19997,N_17499,N_17077);
or U19998 (N_19998,N_17832,N_16069);
xnor U19999 (N_19999,N_16444,N_17930);
and U20000 (N_20000,N_19761,N_18825);
xnor U20001 (N_20001,N_19343,N_19482);
nand U20002 (N_20002,N_19471,N_18397);
nand U20003 (N_20003,N_18837,N_18316);
xnor U20004 (N_20004,N_19551,N_19206);
xnor U20005 (N_20005,N_18019,N_19142);
or U20006 (N_20006,N_18456,N_18520);
nor U20007 (N_20007,N_19659,N_18741);
or U20008 (N_20008,N_19284,N_19825);
nor U20009 (N_20009,N_19481,N_19261);
and U20010 (N_20010,N_19915,N_19675);
nor U20011 (N_20011,N_19706,N_18766);
nor U20012 (N_20012,N_19589,N_18988);
nand U20013 (N_20013,N_19328,N_19297);
nor U20014 (N_20014,N_19055,N_18812);
or U20015 (N_20015,N_19906,N_19337);
nor U20016 (N_20016,N_19074,N_19145);
nor U20017 (N_20017,N_18166,N_18896);
or U20018 (N_20018,N_18755,N_19827);
or U20019 (N_20019,N_18479,N_18150);
xor U20020 (N_20020,N_19548,N_19900);
nand U20021 (N_20021,N_18453,N_18518);
and U20022 (N_20022,N_19495,N_18129);
or U20023 (N_20023,N_19193,N_19536);
nor U20024 (N_20024,N_18650,N_19355);
nand U20025 (N_20025,N_19568,N_19350);
and U20026 (N_20026,N_18949,N_18685);
or U20027 (N_20027,N_19034,N_19505);
xor U20028 (N_20028,N_18757,N_19420);
or U20029 (N_20029,N_18279,N_18818);
and U20030 (N_20030,N_18706,N_18032);
and U20031 (N_20031,N_18756,N_19773);
nand U20032 (N_20032,N_18596,N_18199);
and U20033 (N_20033,N_19741,N_18508);
and U20034 (N_20034,N_18249,N_18463);
and U20035 (N_20035,N_18382,N_19131);
xor U20036 (N_20036,N_18945,N_18370);
and U20037 (N_20037,N_19240,N_19744);
nor U20038 (N_20038,N_19704,N_19690);
xor U20039 (N_20039,N_18295,N_18233);
and U20040 (N_20040,N_18272,N_19214);
nand U20041 (N_20041,N_18388,N_18642);
nor U20042 (N_20042,N_18220,N_19517);
and U20043 (N_20043,N_18428,N_18173);
nor U20044 (N_20044,N_19788,N_18708);
and U20045 (N_20045,N_19533,N_19671);
nand U20046 (N_20046,N_19263,N_18012);
nand U20047 (N_20047,N_18512,N_18466);
and U20048 (N_20048,N_19160,N_18528);
and U20049 (N_20049,N_18513,N_18696);
xnor U20050 (N_20050,N_18433,N_18779);
and U20051 (N_20051,N_18865,N_19040);
nor U20052 (N_20052,N_19881,N_18728);
xnor U20053 (N_20053,N_18114,N_19324);
or U20054 (N_20054,N_19635,N_18355);
nand U20055 (N_20055,N_18315,N_19114);
or U20056 (N_20056,N_18634,N_18296);
nand U20057 (N_20057,N_19331,N_19384);
nand U20058 (N_20058,N_19856,N_18658);
or U20059 (N_20059,N_19338,N_18432);
xor U20060 (N_20060,N_19645,N_19027);
or U20061 (N_20061,N_19001,N_19200);
and U20062 (N_20062,N_19751,N_18835);
nand U20063 (N_20063,N_18345,N_18711);
or U20064 (N_20064,N_18498,N_18243);
xor U20065 (N_20065,N_19219,N_18346);
or U20066 (N_20066,N_18516,N_18142);
nand U20067 (N_20067,N_18123,N_18542);
nand U20068 (N_20068,N_18308,N_19208);
nand U20069 (N_20069,N_19466,N_19388);
or U20070 (N_20070,N_18043,N_18965);
nor U20071 (N_20071,N_18935,N_18442);
and U20072 (N_20072,N_19380,N_18020);
and U20073 (N_20073,N_19873,N_18703);
or U20074 (N_20074,N_18098,N_18564);
nor U20075 (N_20075,N_18917,N_19707);
nor U20076 (N_20076,N_19258,N_18833);
nand U20077 (N_20077,N_19799,N_19248);
xor U20078 (N_20078,N_19766,N_18876);
nand U20079 (N_20079,N_19362,N_18036);
nand U20080 (N_20080,N_18499,N_18090);
nand U20081 (N_20081,N_19941,N_19436);
nand U20082 (N_20082,N_19912,N_19394);
nor U20083 (N_20083,N_18571,N_19299);
nor U20084 (N_20084,N_18033,N_19419);
xor U20085 (N_20085,N_18301,N_18413);
or U20086 (N_20086,N_18152,N_18104);
nand U20087 (N_20087,N_19479,N_19218);
nor U20088 (N_20088,N_18930,N_18815);
and U20089 (N_20089,N_18053,N_18964);
nor U20090 (N_20090,N_19532,N_18938);
nor U20091 (N_20091,N_18656,N_18067);
and U20092 (N_20092,N_18664,N_19545);
xnor U20093 (N_20093,N_19884,N_19181);
nor U20094 (N_20094,N_18377,N_18080);
xnor U20095 (N_20095,N_19192,N_19225);
and U20096 (N_20096,N_19801,N_18344);
nor U20097 (N_20097,N_18335,N_18286);
nand U20098 (N_20098,N_19427,N_19168);
nor U20099 (N_20099,N_18726,N_18869);
nand U20100 (N_20100,N_19603,N_18532);
or U20101 (N_20101,N_19846,N_19991);
and U20102 (N_20102,N_19796,N_19425);
or U20103 (N_20103,N_18617,N_18806);
nor U20104 (N_20104,N_18995,N_18299);
nand U20105 (N_20105,N_18076,N_18576);
nand U20106 (N_20106,N_19945,N_19819);
xnor U20107 (N_20107,N_18115,N_19512);
nor U20108 (N_20108,N_18899,N_19893);
nor U20109 (N_20109,N_18572,N_18647);
xor U20110 (N_20110,N_19389,N_19653);
nor U20111 (N_20111,N_18278,N_18409);
or U20112 (N_20112,N_18385,N_18307);
xnor U20113 (N_20113,N_18934,N_19021);
and U20114 (N_20114,N_19600,N_18188);
nand U20115 (N_20115,N_19951,N_19584);
nand U20116 (N_20116,N_18901,N_18170);
and U20117 (N_20117,N_19919,N_18544);
or U20118 (N_20118,N_18100,N_18585);
and U20119 (N_20119,N_19238,N_19890);
nand U20120 (N_20120,N_18419,N_19613);
or U20121 (N_20121,N_18798,N_19958);
xnor U20122 (N_20122,N_18514,N_18963);
or U20123 (N_20123,N_18029,N_18954);
xnor U20124 (N_20124,N_18288,N_19469);
nor U20125 (N_20125,N_19336,N_18530);
nand U20126 (N_20126,N_18410,N_18504);
nand U20127 (N_20127,N_18027,N_19026);
xor U20128 (N_20128,N_19538,N_18582);
and U20129 (N_20129,N_19360,N_19904);
nand U20130 (N_20130,N_19777,N_18169);
nand U20131 (N_20131,N_18007,N_19562);
xnor U20132 (N_20132,N_18439,N_18016);
and U20133 (N_20133,N_18776,N_18636);
nand U20134 (N_20134,N_19046,N_18805);
and U20135 (N_20135,N_19174,N_18045);
xor U20136 (N_20136,N_18227,N_19000);
or U20137 (N_20137,N_19073,N_19230);
or U20138 (N_20138,N_19688,N_18823);
and U20139 (N_20139,N_19296,N_18222);
nor U20140 (N_20140,N_18905,N_18376);
xor U20141 (N_20141,N_19746,N_19334);
nand U20142 (N_20142,N_18488,N_18049);
and U20143 (N_20143,N_18167,N_19062);
nor U20144 (N_20144,N_18487,N_19226);
or U20145 (N_20145,N_19935,N_18793);
nand U20146 (N_20146,N_19699,N_18135);
or U20147 (N_20147,N_18782,N_18883);
and U20148 (N_20148,N_18729,N_19647);
xnor U20149 (N_20149,N_18481,N_18071);
nor U20150 (N_20150,N_18072,N_19433);
nand U20151 (N_20151,N_18662,N_18052);
nor U20152 (N_20152,N_19292,N_18446);
nor U20153 (N_20153,N_18816,N_19458);
nor U20154 (N_20154,N_18490,N_18943);
nand U20155 (N_20155,N_19866,N_19447);
or U20156 (N_20156,N_18610,N_18213);
nor U20157 (N_20157,N_18799,N_19249);
or U20158 (N_20158,N_19088,N_19477);
and U20159 (N_20159,N_18602,N_19685);
nand U20160 (N_20160,N_18615,N_18004);
and U20161 (N_20161,N_18984,N_18986);
nand U20162 (N_20162,N_18834,N_19570);
and U20163 (N_20163,N_19408,N_18452);
and U20164 (N_20164,N_18441,N_18973);
xnor U20165 (N_20165,N_18753,N_19998);
xnor U20166 (N_20166,N_19378,N_19182);
and U20167 (N_20167,N_18342,N_19438);
xor U20168 (N_20168,N_19674,N_19937);
xnor U20169 (N_20169,N_18219,N_19515);
and U20170 (N_20170,N_19139,N_19076);
xnor U20171 (N_20171,N_18113,N_19845);
or U20172 (N_20172,N_19332,N_18786);
nand U20173 (N_20173,N_18593,N_19650);
and U20174 (N_20174,N_19767,N_18525);
nor U20175 (N_20175,N_18125,N_18721);
nor U20176 (N_20176,N_18624,N_18009);
nand U20177 (N_20177,N_18160,N_18505);
nor U20178 (N_20178,N_19004,N_18074);
and U20179 (N_20179,N_19883,N_19453);
xnor U20180 (N_20180,N_18886,N_19760);
nand U20181 (N_20181,N_18861,N_18948);
nand U20182 (N_20182,N_19109,N_18124);
or U20183 (N_20183,N_18459,N_18569);
nand U20184 (N_20184,N_18814,N_18822);
or U20185 (N_20185,N_19785,N_18797);
and U20186 (N_20186,N_19141,N_18700);
nor U20187 (N_20187,N_18655,N_19493);
nand U20188 (N_20188,N_18083,N_19916);
nor U20189 (N_20189,N_19780,N_18095);
or U20190 (N_20190,N_18214,N_18399);
nand U20191 (N_20191,N_18707,N_19103);
xnor U20192 (N_20192,N_18749,N_19606);
nand U20193 (N_20193,N_19198,N_18063);
and U20194 (N_20194,N_18827,N_18107);
or U20195 (N_20195,N_18851,N_18185);
nor U20196 (N_20196,N_19499,N_18578);
nor U20197 (N_20197,N_19352,N_18174);
nand U20198 (N_20198,N_19676,N_18946);
xor U20199 (N_20199,N_18875,N_19740);
and U20200 (N_20200,N_18927,N_18191);
or U20201 (N_20201,N_19077,N_18130);
nor U20202 (N_20202,N_18681,N_19490);
nor U20203 (N_20203,N_19692,N_18939);
nand U20204 (N_20204,N_19700,N_19564);
xor U20205 (N_20205,N_18400,N_18161);
nand U20206 (N_20206,N_18424,N_19423);
xnor U20207 (N_20207,N_19960,N_18319);
and U20208 (N_20208,N_19483,N_19223);
nand U20209 (N_20209,N_19289,N_18715);
xor U20210 (N_20210,N_18506,N_18637);
nand U20211 (N_20211,N_18180,N_18772);
nor U20212 (N_20212,N_18341,N_18343);
or U20213 (N_20213,N_18443,N_19455);
or U20214 (N_20214,N_18960,N_18491);
and U20215 (N_20215,N_18678,N_18460);
xnor U20216 (N_20216,N_19013,N_19311);
nand U20217 (N_20217,N_18641,N_18751);
and U20218 (N_20218,N_19014,N_19898);
and U20219 (N_20219,N_19537,N_18712);
nor U20220 (N_20220,N_18752,N_18181);
xor U20221 (N_20221,N_18689,N_19146);
nand U20222 (N_20222,N_18607,N_19778);
nor U20223 (N_20223,N_18122,N_19703);
nor U20224 (N_20224,N_18110,N_18131);
nor U20225 (N_20225,N_18415,N_18209);
nor U20226 (N_20226,N_19376,N_18334);
or U20227 (N_20227,N_18026,N_19309);
nor U20228 (N_20228,N_19303,N_19640);
or U20229 (N_20229,N_19179,N_18785);
and U20230 (N_20230,N_19984,N_19725);
xnor U20231 (N_20231,N_18897,N_19059);
nand U20232 (N_20232,N_19604,N_18257);
nand U20233 (N_20233,N_19968,N_19401);
or U20234 (N_20234,N_18620,N_18325);
xnor U20235 (N_20235,N_18966,N_18489);
nor U20236 (N_20236,N_18760,N_19122);
or U20237 (N_20237,N_18193,N_18811);
xor U20238 (N_20238,N_19136,N_19670);
nand U20239 (N_20239,N_18884,N_19366);
and U20240 (N_20240,N_18105,N_19615);
nand U20241 (N_20241,N_19201,N_18872);
xnor U20242 (N_20242,N_19634,N_19468);
nand U20243 (N_20243,N_18991,N_18612);
nand U20244 (N_20244,N_18996,N_18575);
nand U20245 (N_20245,N_18839,N_19057);
and U20246 (N_20246,N_18163,N_18015);
nor U20247 (N_20247,N_19246,N_19903);
nand U20248 (N_20248,N_18900,N_18970);
or U20249 (N_20249,N_19070,N_19185);
nor U20250 (N_20250,N_19843,N_19730);
and U20251 (N_20251,N_19295,N_19421);
and U20252 (N_20252,N_19178,N_18842);
and U20253 (N_20253,N_19112,N_19808);
nand U20254 (N_20254,N_19979,N_19925);
nor U20255 (N_20255,N_19478,N_18549);
nand U20256 (N_20256,N_19702,N_18294);
or U20257 (N_20257,N_18724,N_19552);
xor U20258 (N_20258,N_18248,N_19412);
xnor U20259 (N_20259,N_18064,N_18661);
and U20260 (N_20260,N_18195,N_18788);
nand U20261 (N_20261,N_18849,N_19508);
or U20262 (N_20262,N_19871,N_18857);
xor U20263 (N_20263,N_19831,N_18539);
nand U20264 (N_20264,N_19115,N_19535);
nor U20265 (N_20265,N_18373,N_19099);
or U20266 (N_20266,N_18958,N_19422);
nand U20267 (N_20267,N_19762,N_19771);
nor U20268 (N_20268,N_19449,N_18175);
or U20269 (N_20269,N_18137,N_18298);
nor U20270 (N_20270,N_18482,N_19528);
nand U20271 (N_20271,N_19267,N_19863);
nor U20272 (N_20272,N_18402,N_19180);
xnor U20273 (N_20273,N_19460,N_18186);
xnor U20274 (N_20274,N_18024,N_18116);
xor U20275 (N_20275,N_18283,N_19577);
and U20276 (N_20276,N_19934,N_18030);
and U20277 (N_20277,N_19559,N_19134);
nor U20278 (N_20278,N_19504,N_18391);
nand U20279 (N_20279,N_18077,N_18312);
nand U20280 (N_20280,N_19498,N_19853);
or U20281 (N_20281,N_19723,N_18903);
and U20282 (N_20282,N_19291,N_18465);
nand U20283 (N_20283,N_19092,N_19591);
or U20284 (N_20284,N_19507,N_19812);
and U20285 (N_20285,N_19339,N_19015);
nand U20286 (N_20286,N_19789,N_18885);
nand U20287 (N_20287,N_18727,N_18062);
nand U20288 (N_20288,N_18500,N_19541);
and U20289 (N_20289,N_18638,N_18533);
nand U20290 (N_20290,N_18944,N_19031);
nand U20291 (N_20291,N_19410,N_18853);
nand U20292 (N_20292,N_18523,N_18069);
or U20293 (N_20293,N_19628,N_18709);
nand U20294 (N_20294,N_19855,N_18234);
and U20295 (N_20295,N_18338,N_19260);
and U20296 (N_20296,N_18055,N_18867);
and U20297 (N_20297,N_18092,N_19278);
and U20298 (N_20298,N_18556,N_19983);
xnor U20299 (N_20299,N_19834,N_18239);
or U20300 (N_20300,N_19071,N_19089);
nor U20301 (N_20301,N_19156,N_18980);
or U20302 (N_20302,N_19082,N_19413);
or U20303 (N_20303,N_18494,N_18887);
and U20304 (N_20304,N_18652,N_18144);
nor U20305 (N_20305,N_19739,N_19795);
nand U20306 (N_20306,N_18739,N_18282);
and U20307 (N_20307,N_18522,N_19157);
and U20308 (N_20308,N_18651,N_19164);
xnor U20309 (N_20309,N_19665,N_19727);
xnor U20310 (N_20310,N_18371,N_19110);
nand U20311 (N_20311,N_19068,N_19287);
nand U20312 (N_20312,N_19682,N_18904);
nand U20313 (N_20313,N_19529,N_19784);
nor U20314 (N_20314,N_19794,N_18543);
and U20315 (N_20315,N_18224,N_18425);
nand U20316 (N_20316,N_19555,N_18691);
nor U20317 (N_20317,N_19901,N_19828);
and U20318 (N_20318,N_19631,N_18380);
or U20319 (N_20319,N_19921,N_19950);
and U20320 (N_20320,N_18770,N_18235);
nand U20321 (N_20321,N_18117,N_19010);
and U20322 (N_20322,N_19032,N_19143);
or U20323 (N_20323,N_19657,N_19609);
nor U20324 (N_20324,N_19569,N_19188);
xnor U20325 (N_20325,N_18390,N_18916);
and U20326 (N_20326,N_18293,N_18644);
xor U20327 (N_20327,N_19470,N_18746);
xnor U20328 (N_20328,N_18720,N_18046);
xnor U20329 (N_20329,N_19837,N_19851);
xor U20330 (N_20330,N_18372,N_19683);
nor U20331 (N_20331,N_18127,N_18730);
xnor U20332 (N_20332,N_18541,N_19752);
nor U20333 (N_20333,N_18606,N_19830);
xor U20334 (N_20334,N_19839,N_19779);
xnor U20335 (N_20335,N_19043,N_19662);
nor U20336 (N_20336,N_19572,N_18919);
nand U20337 (N_20337,N_18592,N_19868);
and U20338 (N_20338,N_18416,N_19877);
or U20339 (N_20339,N_19909,N_19158);
or U20340 (N_20340,N_18737,N_18665);
or U20341 (N_20341,N_19587,N_19857);
nor U20342 (N_20342,N_19583,N_18982);
nor U20343 (N_20343,N_19372,N_19588);
nor U20344 (N_20344,N_18354,N_18314);
and U20345 (N_20345,N_19905,N_19742);
or U20346 (N_20346,N_18616,N_19215);
xnor U20347 (N_20347,N_18601,N_18112);
xor U20348 (N_20348,N_19244,N_19306);
nand U20349 (N_20349,N_18281,N_18526);
xor U20350 (N_20350,N_19502,N_19733);
xor U20351 (N_20351,N_18898,N_19140);
and U20352 (N_20352,N_19133,N_19993);
and U20353 (N_20353,N_19988,N_19654);
nor U20354 (N_20354,N_18566,N_19045);
nand U20355 (N_20355,N_19687,N_19861);
or U20356 (N_20356,N_19323,N_18438);
nor U20357 (N_20357,N_19017,N_18947);
nand U20358 (N_20358,N_19491,N_18686);
nor U20359 (N_20359,N_18826,N_19966);
or U20360 (N_20360,N_18629,N_18363);
xor U20361 (N_20361,N_18829,N_18205);
or U20362 (N_20362,N_18471,N_19847);
xnor U20363 (N_20363,N_19667,N_19571);
and U20364 (N_20364,N_18436,N_18990);
nand U20365 (N_20365,N_19041,N_18396);
nor U20366 (N_20366,N_19770,N_19550);
nand U20367 (N_20367,N_19203,N_19177);
nand U20368 (N_20368,N_19279,N_19149);
nor U20369 (N_20369,N_19818,N_19910);
and U20370 (N_20370,N_18577,N_19629);
or U20371 (N_20371,N_18676,N_19756);
nand U20372 (N_20372,N_19623,N_18042);
or U20373 (N_20373,N_19930,N_19269);
xnor U20374 (N_20374,N_19633,N_19123);
xor U20375 (N_20375,N_19975,N_19962);
xnor U20376 (N_20376,N_19037,N_18911);
nor U20377 (N_20377,N_18061,N_18977);
nor U20378 (N_20378,N_18058,N_19035);
nand U20379 (N_20379,N_19409,N_18418);
xor U20380 (N_20380,N_18010,N_19353);
nor U20381 (N_20381,N_19186,N_19902);
and U20382 (N_20382,N_18177,N_18111);
xnor U20383 (N_20383,N_18734,N_18747);
nor U20384 (N_20384,N_18736,N_19716);
nor U20385 (N_20385,N_18987,N_19227);
xnor U20386 (N_20386,N_18365,N_18368);
or U20387 (N_20387,N_19245,N_19152);
or U20388 (N_20388,N_18744,N_18348);
xnor U20389 (N_20389,N_19250,N_19982);
nor U20390 (N_20390,N_19737,N_19549);
and U20391 (N_20391,N_19989,N_19257);
xnor U20392 (N_20392,N_18232,N_18820);
or U20393 (N_20393,N_18358,N_19184);
nand U20394 (N_20394,N_18262,N_18059);
or U20395 (N_20395,N_19300,N_19557);
or U20396 (N_20396,N_18978,N_18565);
and U20397 (N_20397,N_18581,N_19663);
nand U20398 (N_20398,N_19308,N_18657);
or U20399 (N_20399,N_19803,N_18017);
and U20400 (N_20400,N_19660,N_18289);
nor U20401 (N_20401,N_19882,N_19539);
and U20402 (N_20402,N_18194,N_19524);
nor U20403 (N_20403,N_18156,N_18492);
xnor U20404 (N_20404,N_19724,N_18484);
and U20405 (N_20405,N_18604,N_19302);
xnor U20406 (N_20406,N_18969,N_19170);
xnor U20407 (N_20407,N_19695,N_18961);
or U20408 (N_20408,N_19363,N_18226);
xnor U20409 (N_20409,N_19457,N_18085);
and U20410 (N_20410,N_19116,N_18777);
and U20411 (N_20411,N_18906,N_19063);
and U20412 (N_20412,N_19321,N_18773);
nand U20413 (N_20413,N_19393,N_18732);
nand U20414 (N_20414,N_18480,N_18750);
or U20415 (N_20415,N_19519,N_18132);
nor U20416 (N_20416,N_19987,N_18268);
nand U20417 (N_20417,N_19782,N_18445);
nor U20418 (N_20418,N_19494,N_18557);
and U20419 (N_20419,N_19165,N_19025);
nor U20420 (N_20420,N_18148,N_19052);
xnor U20421 (N_20421,N_19084,N_19439);
nand U20422 (N_20422,N_18364,N_18051);
nand U20423 (N_20423,N_18347,N_19642);
xor U20424 (N_20424,N_19392,N_19500);
nand U20425 (N_20425,N_19585,N_18369);
nor U20426 (N_20426,N_19897,N_19224);
xnor U20427 (N_20427,N_18225,N_19486);
nand U20428 (N_20428,N_19108,N_19632);
and U20429 (N_20429,N_18863,N_18472);
or U20430 (N_20430,N_18192,N_18457);
and U20431 (N_20431,N_19820,N_19489);
nand U20432 (N_20432,N_18120,N_19608);
and U20433 (N_20433,N_18423,N_19416);
xor U20434 (N_20434,N_18240,N_18168);
or U20435 (N_20435,N_19829,N_18710);
or U20436 (N_20436,N_19908,N_19712);
or U20437 (N_20437,N_19042,N_19672);
xnor U20438 (N_20438,N_19102,N_19781);
nand U20439 (N_20439,N_18183,N_18246);
nor U20440 (N_20440,N_18450,N_18337);
nand U20441 (N_20441,N_18992,N_18803);
nor U20442 (N_20442,N_19621,N_19996);
or U20443 (N_20443,N_19816,N_18824);
nand U20444 (N_20444,N_19199,N_18221);
nand U20445 (N_20445,N_18999,N_19617);
or U20446 (N_20446,N_18014,N_19256);
or U20447 (N_20447,N_19889,N_18748);
or U20448 (N_20448,N_18204,N_19277);
nand U20449 (N_20449,N_19920,N_19605);
nor U20450 (N_20450,N_19128,N_18106);
xor U20451 (N_20451,N_18646,N_18599);
or U20452 (N_20452,N_18890,N_19560);
and U20453 (N_20453,N_18360,N_18159);
nand U20454 (N_20454,N_18412,N_18587);
xnor U20455 (N_20455,N_18340,N_19811);
nor U20456 (N_20456,N_19440,N_18972);
nor U20457 (N_20457,N_18554,N_18109);
or U20458 (N_20458,N_18623,N_19774);
or U20459 (N_20459,N_18379,N_18197);
or U20460 (N_20460,N_18330,N_18807);
and U20461 (N_20461,N_18912,N_18780);
and U20462 (N_20462,N_18247,N_18942);
nor U20463 (N_20463,N_18073,N_19406);
or U20464 (N_20464,N_18395,N_19121);
and U20465 (N_20465,N_19511,N_19862);
and U20466 (N_20466,N_19091,N_18324);
xor U20467 (N_20467,N_18719,N_19018);
nor U20468 (N_20468,N_19253,N_19161);
and U20469 (N_20469,N_18006,N_18202);
and U20470 (N_20470,N_18447,N_19361);
nor U20471 (N_20471,N_19558,N_19262);
or U20472 (N_20472,N_18769,N_19776);
or U20473 (N_20473,N_18800,N_19579);
nor U20474 (N_20474,N_19317,N_18787);
xnor U20475 (N_20475,N_18091,N_18429);
or U20476 (N_20476,N_19636,N_18403);
nor U20477 (N_20477,N_19722,N_18626);
nor U20478 (N_20478,N_19876,N_19163);
nor U20479 (N_20479,N_18189,N_19807);
nand U20480 (N_20480,N_19484,N_18310);
nand U20481 (N_20481,N_19333,N_18795);
xnor U20482 (N_20482,N_19233,N_18796);
nor U20483 (N_20483,N_18553,N_19620);
and U20484 (N_20484,N_18555,N_19171);
nor U20485 (N_20485,N_18044,N_18094);
or U20486 (N_20486,N_18690,N_18630);
and U20487 (N_20487,N_19802,N_18420);
nor U20488 (N_20488,N_19094,N_18668);
nor U20489 (N_20489,N_18493,N_19150);
xor U20490 (N_20490,N_19415,N_19607);
nand U20491 (N_20491,N_19405,N_19117);
or U20492 (N_20492,N_18361,N_19044);
nand U20493 (N_20493,N_19923,N_18790);
nor U20494 (N_20494,N_18603,N_19106);
or U20495 (N_20495,N_19213,N_18745);
nor U20496 (N_20496,N_18473,N_18392);
nand U20497 (N_20497,N_19349,N_19891);
xor U20498 (N_20498,N_19735,N_18635);
or U20499 (N_20499,N_19154,N_18187);
nor U20500 (N_20500,N_18983,N_19518);
xnor U20501 (N_20501,N_18831,N_18099);
nor U20502 (N_20502,N_18041,N_19849);
xnor U20503 (N_20503,N_19053,N_19793);
nor U20504 (N_20504,N_18464,N_19243);
xnor U20505 (N_20505,N_19973,N_19124);
and U20506 (N_20506,N_19093,N_18065);
xor U20507 (N_20507,N_19974,N_19467);
nand U20508 (N_20508,N_18843,N_18921);
xnor U20509 (N_20509,N_19701,N_19473);
or U20510 (N_20510,N_19516,N_18147);
and U20511 (N_20511,N_18317,N_18519);
and U20512 (N_20512,N_18674,N_18529);
xor U20513 (N_20513,N_19926,N_19651);
or U20514 (N_20514,N_19946,N_18216);
and U20515 (N_20515,N_18366,N_19813);
nand U20516 (N_20516,N_18735,N_19720);
xor U20517 (N_20517,N_19948,N_18375);
nand U20518 (N_20518,N_18266,N_18922);
nor U20519 (N_20519,N_19036,N_19643);
or U20520 (N_20520,N_19325,N_18877);
xnor U20521 (N_20521,N_19242,N_19932);
and U20522 (N_20522,N_19060,N_19576);
and U20523 (N_20523,N_19971,N_18121);
or U20524 (N_20524,N_19750,N_18672);
or U20525 (N_20525,N_18190,N_19451);
nand U20526 (N_20526,N_19590,N_19288);
nor U20527 (N_20527,N_19228,N_19497);
xor U20528 (N_20528,N_18475,N_19790);
nor U20529 (N_20529,N_18448,N_18435);
and U20530 (N_20530,N_18667,N_19523);
xor U20531 (N_20531,N_19083,N_19972);
nand U20532 (N_20532,N_18979,N_18868);
and U20533 (N_20533,N_18230,N_19918);
nor U20534 (N_20534,N_19952,N_18567);
nor U20535 (N_20535,N_19356,N_19506);
xnor U20536 (N_20536,N_18840,N_19999);
or U20537 (N_20537,N_19953,N_18427);
and U20538 (N_20538,N_19978,N_18149);
nand U20539 (N_20539,N_19681,N_18684);
or U20540 (N_20540,N_19475,N_19664);
and U20541 (N_20541,N_19009,N_18879);
nor U20542 (N_20542,N_19315,N_18039);
and U20543 (N_20543,N_18619,N_19397);
or U20544 (N_20544,N_19748,N_18300);
and U20545 (N_20545,N_18929,N_18210);
xor U20546 (N_20546,N_18931,N_18430);
xnor U20547 (N_20547,N_19581,N_18251);
nor U20548 (N_20548,N_18588,N_19622);
nand U20549 (N_20549,N_19835,N_18962);
xor U20550 (N_20550,N_19379,N_19661);
nor U20551 (N_20551,N_19434,N_19574);
nand U20552 (N_20552,N_19282,N_19765);
and U20553 (N_20553,N_18218,N_19673);
xor U20554 (N_20554,N_18932,N_18146);
nor U20555 (N_20555,N_18495,N_18666);
or U20556 (N_20556,N_18066,N_19592);
nand U20557 (N_20557,N_18383,N_19254);
nor U20558 (N_20558,N_19342,N_18697);
and U20559 (N_20559,N_19326,N_19020);
nor U20560 (N_20560,N_18951,N_19313);
nand U20561 (N_20561,N_18040,N_18968);
xnor U20562 (N_20562,N_19899,N_18950);
and U20563 (N_20563,N_19721,N_19189);
nand U20564 (N_20564,N_18001,N_19067);
or U20565 (N_20565,N_19236,N_19575);
xnor U20566 (N_20566,N_18421,N_19307);
or U20567 (N_20567,N_18631,N_18359);
or U20568 (N_20568,N_19066,N_18303);
or U20569 (N_20569,N_19867,N_19879);
nand U20570 (N_20570,N_18694,N_19832);
xnor U20571 (N_20571,N_18290,N_18386);
xor U20572 (N_20572,N_19369,N_18184);
nand U20573 (N_20573,N_19459,N_19922);
xor U20574 (N_20574,N_18546,N_19514);
xor U20575 (N_20575,N_18398,N_19414);
nand U20576 (N_20576,N_18614,N_19431);
and U20577 (N_20577,N_18524,N_19387);
xnor U20578 (N_20578,N_19065,N_19016);
nor U20579 (N_20579,N_19464,N_18570);
xor U20580 (N_20580,N_18406,N_19864);
and U20581 (N_20581,N_18873,N_18659);
or U20582 (N_20582,N_18352,N_18705);
and U20583 (N_20583,N_19119,N_18971);
and U20584 (N_20584,N_19865,N_19521);
nand U20585 (N_20585,N_18817,N_19513);
nor U20586 (N_20586,N_19810,N_18118);
xnor U20587 (N_20587,N_19544,N_19275);
xor U20588 (N_20588,N_19652,N_18154);
nand U20589 (N_20589,N_19990,N_19522);
xnor U20590 (N_20590,N_19602,N_19169);
and U20591 (N_20591,N_19098,N_19463);
or U20592 (N_20592,N_18079,N_19527);
nand U20593 (N_20593,N_18075,N_18362);
or U20594 (N_20594,N_19496,N_19693);
nor U20595 (N_20595,N_19713,N_18993);
and U20596 (N_20596,N_18444,N_18483);
xnor U20597 (N_20597,N_18236,N_19395);
and U20598 (N_20598,N_19312,N_18178);
nand U20599 (N_20599,N_18321,N_18633);
nand U20600 (N_20600,N_18537,N_18561);
nor U20601 (N_20601,N_19113,N_19492);
nor U20602 (N_20602,N_19929,N_19896);
xor U20603 (N_20603,N_18411,N_18560);
nor U20604 (N_20604,N_18910,N_18208);
and U20605 (N_20605,N_19085,N_18153);
xor U20606 (N_20606,N_18468,N_18759);
and U20607 (N_20607,N_19358,N_18309);
or U20608 (N_20608,N_19424,N_19530);
and U20609 (N_20609,N_19407,N_18196);
and U20610 (N_20610,N_18176,N_18384);
nor U20611 (N_20611,N_19656,N_19173);
nor U20612 (N_20612,N_18654,N_19259);
or U20613 (N_20613,N_19894,N_19194);
nand U20614 (N_20614,N_18622,N_19265);
xor U20615 (N_20615,N_18139,N_19126);
and U20616 (N_20616,N_18378,N_18941);
nor U20617 (N_20617,N_18573,N_18864);
and U20618 (N_20618,N_18056,N_18967);
or U20619 (N_20619,N_19969,N_18809);
nand U20620 (N_20620,N_19520,N_18260);
nand U20621 (N_20621,N_19383,N_18791);
nand U20622 (N_20622,N_18164,N_19429);
and U20623 (N_20623,N_19050,N_19005);
nand U20624 (N_20624,N_19344,N_19273);
nand U20625 (N_20625,N_18401,N_18957);
nand U20626 (N_20626,N_18761,N_18021);
and U20627 (N_20627,N_18141,N_19708);
or U20628 (N_20628,N_18847,N_19854);
and U20629 (N_20629,N_18171,N_18552);
xnor U20630 (N_20630,N_19710,N_19054);
nand U20631 (N_20631,N_19627,N_18848);
nand U20632 (N_20632,N_19954,N_18742);
and U20633 (N_20633,N_19276,N_19485);
xnor U20634 (N_20634,N_19705,N_19578);
xnor U20635 (N_20635,N_19697,N_19456);
nand U20636 (N_20636,N_18828,N_19107);
and U20637 (N_20637,N_19399,N_19911);
xnor U20638 (N_20638,N_19619,N_19446);
and U20639 (N_20639,N_18627,N_18253);
and U20640 (N_20640,N_19135,N_18136);
xnor U20641 (N_20641,N_19480,N_18496);
nand U20642 (N_20642,N_18538,N_18830);
nor U20643 (N_20643,N_19209,N_18273);
nor U20644 (N_20644,N_18680,N_18304);
xor U20645 (N_20645,N_18874,N_18394);
nor U20646 (N_20646,N_18461,N_19365);
xnor U20647 (N_20647,N_19939,N_19105);
xor U20648 (N_20648,N_18937,N_18005);
or U20649 (N_20649,N_18804,N_19285);
nor U20650 (N_20650,N_18060,N_19554);
or U20651 (N_20651,N_18449,N_18455);
and U20652 (N_20652,N_19743,N_19526);
and U20653 (N_20653,N_18259,N_19869);
nor U20654 (N_20654,N_18975,N_18928);
and U20655 (N_20655,N_18200,N_18086);
xnor U20656 (N_20656,N_19049,N_18351);
nor U20657 (N_20657,N_18808,N_19775);
nor U20658 (N_20658,N_18598,N_19913);
xnor U20659 (N_20659,N_18702,N_19985);
xnor U20660 (N_20660,N_19058,N_19561);
nor U20661 (N_20661,N_18521,N_19138);
and U20662 (N_20662,N_19402,N_19211);
nor U20663 (N_20663,N_18920,N_19709);
xnor U20664 (N_20664,N_18859,N_18434);
or U20665 (N_20665,N_19728,N_19241);
nor U20666 (N_20666,N_19942,N_19732);
and U20667 (N_20667,N_19281,N_18589);
xor U20668 (N_20668,N_19069,N_18306);
and U20669 (N_20669,N_18437,N_19593);
xnor U20670 (N_20670,N_19474,N_18892);
nor U20671 (N_20671,N_19805,N_19196);
and U20672 (N_20672,N_18002,N_19007);
nor U20673 (N_20673,N_19826,N_19327);
or U20674 (N_20674,N_18918,N_19204);
xor U20675 (N_20675,N_19417,N_18323);
nand U20676 (N_20676,N_18718,N_19994);
nand U20677 (N_20677,N_18211,N_19210);
and U20678 (N_20678,N_19764,N_18648);
or U20679 (N_20679,N_18801,N_19612);
and U20680 (N_20680,N_19745,N_18908);
and U20681 (N_20681,N_19023,N_19679);
or U20682 (N_20682,N_18695,N_19207);
nand U20683 (N_20683,N_19137,N_18936);
and U20684 (N_20684,N_19172,N_19823);
or U20685 (N_20685,N_19354,N_18836);
nor U20686 (N_20686,N_19127,N_19822);
or U20687 (N_20687,N_19445,N_18893);
nor U20688 (N_20688,N_18203,N_18841);
nor U20689 (N_20689,N_19101,N_19095);
or U20690 (N_20690,N_19783,N_18670);
or U20691 (N_20691,N_18895,N_18215);
xnor U20692 (N_20692,N_19582,N_19019);
nor U20693 (N_20693,N_19833,N_19270);
xor U20694 (N_20694,N_18998,N_18716);
and U20695 (N_20695,N_19283,N_18590);
xnor U20696 (N_20696,N_18832,N_18653);
or U20697 (N_20697,N_19543,N_18802);
and U20698 (N_20698,N_18102,N_18485);
or U20699 (N_20699,N_18784,N_18870);
and U20700 (N_20700,N_18547,N_18902);
or U20701 (N_20701,N_18688,N_18474);
nor U20702 (N_20702,N_19375,N_19144);
or U20703 (N_20703,N_18959,N_19870);
nand U20704 (N_20704,N_19028,N_19729);
xnor U20705 (N_20705,N_18926,N_19648);
nand U20706 (N_20706,N_19821,N_19995);
and U20707 (N_20707,N_18155,N_18733);
and U20708 (N_20708,N_18502,N_19231);
xnor U20709 (N_20709,N_19759,N_18789);
nand U20710 (N_20710,N_18454,N_18274);
nor U20711 (N_20711,N_19510,N_19318);
nor U20712 (N_20712,N_18503,N_18591);
or U20713 (N_20713,N_19809,N_19450);
xor U20714 (N_20714,N_18008,N_19677);
nand U20715 (N_20715,N_18440,N_18140);
or U20716 (N_20716,N_19398,N_18198);
nor U20717 (N_20717,N_19887,N_19970);
nand U20718 (N_20718,N_19222,N_19197);
or U20719 (N_20719,N_19255,N_19166);
or U20720 (N_20720,N_19221,N_19618);
or U20721 (N_20721,N_19329,N_18540);
and U20722 (N_20722,N_18275,N_18731);
xnor U20723 (N_20723,N_19090,N_19237);
or U20724 (N_20724,N_18597,N_19111);
and U20725 (N_20725,N_19928,N_18357);
and U20726 (N_20726,N_18740,N_19509);
xnor U20727 (N_20727,N_19195,N_19462);
xor U20728 (N_20728,N_18649,N_19875);
xnor U20729 (N_20729,N_19914,N_19817);
and U20730 (N_20730,N_19319,N_19646);
xnor U20731 (N_20731,N_18108,N_18333);
nor U20732 (N_20732,N_19432,N_19787);
or U20733 (N_20733,N_18862,N_19151);
and U20734 (N_20734,N_18469,N_18758);
xor U20735 (N_20735,N_18924,N_19757);
or U20736 (N_20736,N_19340,N_18426);
or U20737 (N_20737,N_18261,N_19487);
nand U20738 (N_20738,N_19370,N_19411);
xor U20739 (N_20739,N_19980,N_18022);
nor U20740 (N_20740,N_19003,N_18088);
nand U20741 (N_20741,N_19033,N_19594);
nor U20742 (N_20742,N_19048,N_18866);
and U20743 (N_20743,N_19335,N_19531);
and U20744 (N_20744,N_19461,N_19159);
and U20745 (N_20745,N_19454,N_19949);
nor U20746 (N_20746,N_19611,N_19874);
xnor U20747 (N_20747,N_19373,N_19167);
nand U20748 (N_20748,N_19792,N_18250);
nand U20749 (N_20749,N_18011,N_19357);
xor U20750 (N_20750,N_18813,N_19125);
nand U20751 (N_20751,N_18671,N_18878);
nor U20752 (N_20752,N_19763,N_18034);
nor U20753 (N_20753,N_19341,N_19556);
xor U20754 (N_20754,N_19814,N_19997);
xor U20755 (N_20755,N_18701,N_18374);
or U20756 (N_20756,N_19268,N_19717);
nor U20757 (N_20757,N_18145,N_18608);
nand U20758 (N_20758,N_18517,N_18367);
xnor U20759 (N_20759,N_18417,N_19191);
nor U20760 (N_20760,N_18018,N_19087);
or U20761 (N_20761,N_19155,N_18763);
nand U20762 (N_20762,N_18350,N_18501);
nor U20763 (N_20763,N_19251,N_18302);
and U20764 (N_20764,N_19118,N_19738);
xor U20765 (N_20765,N_19029,N_18256);
xor U20766 (N_20766,N_19859,N_19301);
or U20767 (N_20767,N_19305,N_18414);
and U20768 (N_20768,N_18258,N_19364);
nor U20769 (N_20769,N_19965,N_18477);
xor U20770 (N_20770,N_18128,N_19540);
nand U20771 (N_20771,N_18704,N_19736);
nand U20772 (N_20772,N_19426,N_19658);
nor U20773 (N_20773,N_19888,N_19320);
xor U20774 (N_20774,N_19878,N_18913);
and U20775 (N_20775,N_18618,N_19992);
or U20776 (N_20776,N_18327,N_19981);
nand U20777 (N_20777,N_19931,N_18328);
nand U20778 (N_20778,N_18254,N_18754);
or U20779 (N_20779,N_19595,N_18550);
nand U20780 (N_20780,N_19944,N_18850);
nor U20781 (N_20781,N_18511,N_18771);
nand U20782 (N_20782,N_19836,N_18265);
xnor U20783 (N_20783,N_19924,N_18087);
nor U20784 (N_20784,N_19061,N_19964);
nor U20785 (N_20785,N_18852,N_18119);
or U20786 (N_20786,N_19678,N_18134);
nor U20787 (N_20787,N_19566,N_19239);
xnor U20788 (N_20788,N_19064,N_18625);
nor U20789 (N_20789,N_19002,N_18510);
nand U20790 (N_20790,N_18103,N_18660);
and U20791 (N_20791,N_19755,N_18028);
or U20792 (N_20792,N_18252,N_18238);
xnor U20793 (N_20793,N_18981,N_18269);
and U20794 (N_20794,N_18687,N_19234);
xnor U20795 (N_20795,N_19596,N_19669);
and U20796 (N_20796,N_18003,N_19022);
nand U20797 (N_20797,N_18284,N_18563);
xnor U20798 (N_20798,N_18158,N_19147);
nand U20799 (N_20799,N_18579,N_19860);
nand U20800 (N_20800,N_18639,N_19120);
and U20801 (N_20801,N_18515,N_19444);
nor U20802 (N_20802,N_18621,N_18329);
nor U20803 (N_20803,N_19649,N_18280);
nand U20804 (N_20804,N_18891,N_18698);
and U20805 (N_20805,N_19938,N_18765);
xor U20806 (N_20806,N_18605,N_18548);
nand U20807 (N_20807,N_18332,N_19382);
or U20808 (N_20808,N_18287,N_18387);
and U20809 (N_20809,N_19598,N_18693);
nor U20810 (N_20810,N_18914,N_19346);
xor U20811 (N_20811,N_18404,N_18909);
xnor U20812 (N_20812,N_18889,N_19625);
nand U20813 (N_20813,N_19404,N_19747);
nand U20814 (N_20814,N_18458,N_18267);
xor U20815 (N_20815,N_18940,N_18985);
or U20816 (N_20816,N_18509,N_18923);
xor U20817 (N_20817,N_19842,N_18381);
or U20818 (N_20818,N_18182,N_19100);
or U20819 (N_20819,N_18486,N_19153);
and U20820 (N_20820,N_19310,N_18078);
and U20821 (N_20821,N_18860,N_19686);
nand U20822 (N_20822,N_18682,N_18206);
nand U20823 (N_20823,N_19441,N_18070);
nor U20824 (N_20824,N_19374,N_19465);
and U20825 (N_20825,N_18527,N_19976);
nand U20826 (N_20826,N_18207,N_19086);
xnor U20827 (N_20827,N_18133,N_19488);
nor U20828 (N_20828,N_19216,N_19148);
nand U20829 (N_20829,N_18699,N_19694);
nand U20830 (N_20830,N_18138,N_19428);
xnor U20831 (N_20831,N_18956,N_18047);
nand U20832 (N_20832,N_18212,N_19472);
xor U20833 (N_20833,N_19501,N_18407);
xnor U20834 (N_20834,N_19959,N_18038);
xor U20835 (N_20835,N_18580,N_19711);
nand U20836 (N_20836,N_19205,N_19666);
xnor U20837 (N_20837,N_18462,N_19852);
and U20838 (N_20838,N_18497,N_18143);
and U20839 (N_20839,N_18476,N_18783);
or U20840 (N_20840,N_18881,N_19396);
or U20841 (N_20841,N_18764,N_18393);
nand U20842 (N_20842,N_18792,N_19553);
nor U20843 (N_20843,N_19047,N_19314);
or U20844 (N_20844,N_19104,N_19129);
and U20845 (N_20845,N_19266,N_19437);
or U20846 (N_20846,N_19391,N_19933);
nor U20847 (N_20847,N_18609,N_19271);
and U20848 (N_20848,N_18507,N_19038);
nand U20849 (N_20849,N_19293,N_19655);
nand U20850 (N_20850,N_19290,N_18339);
nand U20851 (N_20851,N_19078,N_18677);
nor U20852 (N_20852,N_19726,N_18349);
nor U20853 (N_20853,N_18632,N_18583);
nor U20854 (N_20854,N_19345,N_18389);
nand U20855 (N_20855,N_19080,N_18068);
and U20856 (N_20856,N_18405,N_18774);
xor U20857 (N_20857,N_18353,N_18050);
nand U20858 (N_20858,N_18242,N_18531);
or U20859 (N_20859,N_19274,N_19547);
or U20860 (N_20860,N_18536,N_19280);
and U20861 (N_20861,N_18331,N_19626);
xnor U20862 (N_20862,N_18692,N_19232);
nand U20863 (N_20863,N_18933,N_18318);
nand U20864 (N_20864,N_18880,N_19714);
or U20865 (N_20865,N_19917,N_19217);
and U20866 (N_20866,N_18326,N_18013);
nand U20867 (N_20867,N_19386,N_18451);
and U20868 (N_20868,N_18534,N_18229);
xor U20869 (N_20869,N_19006,N_18467);
nor U20870 (N_20870,N_19754,N_19986);
or U20871 (N_20871,N_19848,N_19039);
nor U20872 (N_20872,N_18322,N_18285);
nor U20873 (N_20873,N_18856,N_19075);
nand U20874 (N_20874,N_18952,N_19639);
xnor U20875 (N_20875,N_18775,N_18422);
nand U20876 (N_20876,N_19322,N_19542);
and U20877 (N_20877,N_18611,N_18025);
and U20878 (N_20878,N_18974,N_19691);
and U20879 (N_20879,N_18725,N_18640);
nor U20880 (N_20880,N_18297,N_19565);
nand U20881 (N_20881,N_19886,N_19359);
and U20882 (N_20882,N_19844,N_18217);
nand U20883 (N_20883,N_18821,N_19907);
nor U20884 (N_20884,N_18551,N_18157);
nand U20885 (N_20885,N_19024,N_18255);
nor U20886 (N_20886,N_19668,N_18264);
nand U20887 (N_20887,N_19316,N_18955);
nor U20888 (N_20888,N_18925,N_18613);
and U20889 (N_20889,N_19400,N_19132);
nor U20890 (N_20890,N_18762,N_18535);
xnor U20891 (N_20891,N_19008,N_19698);
nor U20892 (N_20892,N_19381,N_19546);
nand U20893 (N_20893,N_19097,N_19264);
xor U20894 (N_20894,N_19418,N_18084);
nand U20895 (N_20895,N_19011,N_18778);
or U20896 (N_20896,N_18478,N_19850);
nand U20897 (N_20897,N_19563,N_19624);
xnor U20898 (N_20898,N_18276,N_18431);
xnor U20899 (N_20899,N_18035,N_19580);
and U20900 (N_20900,N_18245,N_19967);
and U20901 (N_20901,N_19130,N_18584);
or U20902 (N_20902,N_19286,N_18356);
nor U20903 (N_20903,N_19797,N_19749);
nand U20904 (N_20904,N_18679,N_19079);
or U20905 (N_20905,N_18855,N_18722);
and U20906 (N_20906,N_18023,N_18738);
nor U20907 (N_20907,N_19630,N_18000);
xor U20908 (N_20908,N_18819,N_18096);
nand U20909 (N_20909,N_19442,N_19476);
nand U20910 (N_20910,N_19272,N_18717);
nand U20911 (N_20911,N_18558,N_19371);
xnor U20912 (N_20912,N_19503,N_19838);
or U20913 (N_20913,N_19304,N_18645);
xor U20914 (N_20914,N_19936,N_19162);
and U20915 (N_20915,N_18277,N_19927);
nand U20916 (N_20916,N_19885,N_19586);
nand U20917 (N_20917,N_19385,N_18057);
or U20918 (N_20918,N_19403,N_19880);
xnor U20919 (N_20919,N_18470,N_19443);
xnor U20920 (N_20920,N_18336,N_18101);
xor U20921 (N_20921,N_18997,N_19956);
xnor U20922 (N_20922,N_18663,N_19892);
or U20923 (N_20923,N_18082,N_19943);
xor U20924 (N_20924,N_19947,N_18545);
nor U20925 (N_20925,N_18408,N_18320);
xor U20926 (N_20926,N_19212,N_19601);
or U20927 (N_20927,N_19183,N_18767);
nor U20928 (N_20928,N_19815,N_18291);
nor U20929 (N_20929,N_18845,N_18594);
or U20930 (N_20930,N_18894,N_19638);
and U20931 (N_20931,N_19715,N_19719);
nand U20932 (N_20932,N_18311,N_19348);
nand U20933 (N_20933,N_18151,N_18237);
nand U20934 (N_20934,N_18846,N_19351);
or U20935 (N_20935,N_18048,N_19798);
nand U20936 (N_20936,N_18643,N_19734);
nor U20937 (N_20937,N_18714,N_19330);
nand U20938 (N_20938,N_19644,N_19806);
and U20939 (N_20939,N_18162,N_18562);
nor U20940 (N_20940,N_18781,N_18231);
xor U20941 (N_20941,N_19573,N_19298);
nand U20942 (N_20942,N_19448,N_18172);
and U20943 (N_20943,N_19758,N_18907);
nor U20944 (N_20944,N_18810,N_18223);
xnor U20945 (N_20945,N_18673,N_18713);
nand U20946 (N_20946,N_18768,N_19187);
xor U20947 (N_20947,N_18595,N_19824);
nand U20948 (N_20948,N_19347,N_18600);
xor U20949 (N_20949,N_19696,N_18093);
xnor U20950 (N_20950,N_19800,N_19753);
and U20951 (N_20951,N_19977,N_18675);
xnor U20952 (N_20952,N_18271,N_19610);
xor U20953 (N_20953,N_19963,N_19567);
and U20954 (N_20954,N_18097,N_19791);
or U20955 (N_20955,N_19430,N_19840);
and U20956 (N_20956,N_19294,N_18270);
and U20957 (N_20957,N_18244,N_18305);
or U20958 (N_20958,N_18858,N_19895);
nand U20959 (N_20959,N_19452,N_18844);
and U20960 (N_20960,N_19804,N_18574);
nand U20961 (N_20961,N_18871,N_19841);
nor U20962 (N_20962,N_19768,N_19614);
or U20963 (N_20963,N_18559,N_18054);
nor U20964 (N_20964,N_19731,N_19872);
nand U20965 (N_20965,N_19858,N_19051);
and U20966 (N_20966,N_18126,N_18568);
and U20967 (N_20967,N_19252,N_18179);
and U20968 (N_20968,N_18628,N_19368);
nor U20969 (N_20969,N_18031,N_19190);
xnor U20970 (N_20970,N_19030,N_18037);
nand U20971 (N_20971,N_19718,N_18989);
and U20972 (N_20972,N_18089,N_19072);
and U20973 (N_20973,N_19247,N_18228);
nor U20974 (N_20974,N_19175,N_18081);
xnor U20975 (N_20975,N_19202,N_19772);
nor U20976 (N_20976,N_19081,N_19176);
and U20977 (N_20977,N_18241,N_19096);
or U20978 (N_20978,N_18976,N_19435);
nand U20979 (N_20979,N_19786,N_18743);
and U20980 (N_20980,N_19955,N_19641);
nand U20981 (N_20981,N_18838,N_19637);
nand U20982 (N_20982,N_19940,N_18263);
or U20983 (N_20983,N_19684,N_18683);
and U20984 (N_20984,N_19012,N_18669);
nor U20985 (N_20985,N_18854,N_19680);
xor U20986 (N_20986,N_18882,N_18723);
and U20987 (N_20987,N_18888,N_19220);
nor U20988 (N_20988,N_19534,N_19367);
or U20989 (N_20989,N_19616,N_19525);
xor U20990 (N_20990,N_18794,N_18586);
or U20991 (N_20991,N_19377,N_18292);
and U20992 (N_20992,N_19229,N_18313);
nand U20993 (N_20993,N_18165,N_19056);
nor U20994 (N_20994,N_19769,N_19961);
nand U20995 (N_20995,N_19597,N_18953);
xor U20996 (N_20996,N_19957,N_18994);
nor U20997 (N_20997,N_19599,N_19235);
nand U20998 (N_20998,N_18915,N_19689);
nand U20999 (N_20999,N_19390,N_18201);
nand U21000 (N_21000,N_19839,N_19240);
nand U21001 (N_21001,N_18391,N_19672);
xor U21002 (N_21002,N_18871,N_18733);
and U21003 (N_21003,N_19964,N_18133);
or U21004 (N_21004,N_19999,N_18154);
xnor U21005 (N_21005,N_19771,N_19130);
nor U21006 (N_21006,N_19456,N_19063);
xor U21007 (N_21007,N_19945,N_18837);
xnor U21008 (N_21008,N_18056,N_19533);
and U21009 (N_21009,N_18509,N_19126);
and U21010 (N_21010,N_19553,N_19926);
and U21011 (N_21011,N_19450,N_18929);
xor U21012 (N_21012,N_18131,N_19656);
nand U21013 (N_21013,N_19549,N_19193);
or U21014 (N_21014,N_19959,N_19990);
nand U21015 (N_21015,N_19362,N_18262);
or U21016 (N_21016,N_19110,N_18662);
and U21017 (N_21017,N_19042,N_18373);
or U21018 (N_21018,N_19813,N_18145);
nor U21019 (N_21019,N_18537,N_19037);
and U21020 (N_21020,N_18306,N_19255);
and U21021 (N_21021,N_19684,N_19838);
nor U21022 (N_21022,N_18975,N_18331);
and U21023 (N_21023,N_18032,N_19011);
or U21024 (N_21024,N_19462,N_18285);
xnor U21025 (N_21025,N_18652,N_19208);
and U21026 (N_21026,N_18470,N_19229);
or U21027 (N_21027,N_18849,N_19085);
nand U21028 (N_21028,N_18323,N_19232);
nand U21029 (N_21029,N_18880,N_18726);
nand U21030 (N_21030,N_19648,N_19771);
xnor U21031 (N_21031,N_19606,N_18557);
nand U21032 (N_21032,N_19162,N_19208);
xnor U21033 (N_21033,N_19685,N_19664);
and U21034 (N_21034,N_19909,N_18458);
xor U21035 (N_21035,N_18879,N_19011);
nand U21036 (N_21036,N_19493,N_19950);
or U21037 (N_21037,N_18266,N_18182);
nor U21038 (N_21038,N_19640,N_19710);
and U21039 (N_21039,N_19894,N_19793);
xor U21040 (N_21040,N_18958,N_18185);
xor U21041 (N_21041,N_18680,N_19424);
nand U21042 (N_21042,N_19774,N_18577);
nand U21043 (N_21043,N_19054,N_18559);
or U21044 (N_21044,N_19924,N_18430);
nor U21045 (N_21045,N_18020,N_19934);
xnor U21046 (N_21046,N_18340,N_19332);
and U21047 (N_21047,N_19461,N_18960);
nor U21048 (N_21048,N_19719,N_19454);
nor U21049 (N_21049,N_19571,N_19221);
xor U21050 (N_21050,N_18271,N_18373);
and U21051 (N_21051,N_18032,N_19957);
nand U21052 (N_21052,N_19946,N_18726);
nand U21053 (N_21053,N_19504,N_19851);
xnor U21054 (N_21054,N_18089,N_19735);
nand U21055 (N_21055,N_19927,N_18348);
or U21056 (N_21056,N_19314,N_19391);
and U21057 (N_21057,N_18479,N_18891);
nor U21058 (N_21058,N_19713,N_19575);
nand U21059 (N_21059,N_18687,N_19538);
nand U21060 (N_21060,N_18151,N_18497);
nand U21061 (N_21061,N_18053,N_19552);
or U21062 (N_21062,N_19984,N_18418);
and U21063 (N_21063,N_19234,N_19373);
or U21064 (N_21064,N_18983,N_18967);
or U21065 (N_21065,N_18014,N_19377);
nor U21066 (N_21066,N_18287,N_19719);
nor U21067 (N_21067,N_18832,N_19982);
nor U21068 (N_21068,N_18247,N_18180);
nand U21069 (N_21069,N_19861,N_18589);
nand U21070 (N_21070,N_19471,N_19283);
xnor U21071 (N_21071,N_19975,N_19034);
or U21072 (N_21072,N_18032,N_18340);
and U21073 (N_21073,N_18161,N_18346);
and U21074 (N_21074,N_19696,N_18257);
and U21075 (N_21075,N_19781,N_19447);
nand U21076 (N_21076,N_19583,N_18389);
or U21077 (N_21077,N_18605,N_18081);
nand U21078 (N_21078,N_18979,N_19061);
or U21079 (N_21079,N_19832,N_18687);
xnor U21080 (N_21080,N_18065,N_19428);
nand U21081 (N_21081,N_18902,N_19991);
xor U21082 (N_21082,N_19786,N_18546);
and U21083 (N_21083,N_19633,N_18484);
nor U21084 (N_21084,N_19107,N_19881);
xnor U21085 (N_21085,N_19050,N_19424);
nand U21086 (N_21086,N_18032,N_18562);
and U21087 (N_21087,N_19412,N_19113);
nor U21088 (N_21088,N_19992,N_18093);
nand U21089 (N_21089,N_18569,N_18735);
and U21090 (N_21090,N_18109,N_19161);
or U21091 (N_21091,N_19776,N_18682);
nand U21092 (N_21092,N_19840,N_18098);
or U21093 (N_21093,N_19198,N_19881);
nor U21094 (N_21094,N_18388,N_18697);
nor U21095 (N_21095,N_19596,N_18592);
nor U21096 (N_21096,N_19680,N_18901);
xnor U21097 (N_21097,N_18911,N_19644);
and U21098 (N_21098,N_18133,N_18183);
xnor U21099 (N_21099,N_18154,N_19093);
and U21100 (N_21100,N_18009,N_18167);
and U21101 (N_21101,N_18954,N_18850);
xor U21102 (N_21102,N_18476,N_19982);
nand U21103 (N_21103,N_18257,N_18926);
and U21104 (N_21104,N_19907,N_18725);
nand U21105 (N_21105,N_18735,N_19658);
or U21106 (N_21106,N_18547,N_18927);
nor U21107 (N_21107,N_19960,N_18734);
or U21108 (N_21108,N_18347,N_19505);
nand U21109 (N_21109,N_18333,N_19086);
xor U21110 (N_21110,N_19217,N_18931);
or U21111 (N_21111,N_18121,N_18657);
nor U21112 (N_21112,N_18050,N_18909);
and U21113 (N_21113,N_18972,N_18012);
and U21114 (N_21114,N_19153,N_19415);
nor U21115 (N_21115,N_18046,N_18629);
xor U21116 (N_21116,N_19631,N_19207);
or U21117 (N_21117,N_18113,N_19495);
and U21118 (N_21118,N_19220,N_19011);
xor U21119 (N_21119,N_19679,N_19837);
and U21120 (N_21120,N_19642,N_18392);
xnor U21121 (N_21121,N_18164,N_19577);
xor U21122 (N_21122,N_18515,N_18226);
or U21123 (N_21123,N_19166,N_19539);
or U21124 (N_21124,N_19426,N_18376);
or U21125 (N_21125,N_18776,N_18867);
or U21126 (N_21126,N_19071,N_18597);
xnor U21127 (N_21127,N_19619,N_18919);
nor U21128 (N_21128,N_19881,N_18554);
or U21129 (N_21129,N_18660,N_18983);
nor U21130 (N_21130,N_18503,N_19628);
nand U21131 (N_21131,N_18139,N_19384);
or U21132 (N_21132,N_19859,N_19919);
xnor U21133 (N_21133,N_18055,N_18507);
xnor U21134 (N_21134,N_19590,N_19382);
or U21135 (N_21135,N_18473,N_18105);
xnor U21136 (N_21136,N_19480,N_18848);
nor U21137 (N_21137,N_19450,N_18541);
or U21138 (N_21138,N_18917,N_18444);
or U21139 (N_21139,N_18578,N_19104);
nand U21140 (N_21140,N_19934,N_18736);
nor U21141 (N_21141,N_19822,N_19068);
xor U21142 (N_21142,N_18566,N_19983);
xor U21143 (N_21143,N_19575,N_18515);
or U21144 (N_21144,N_19687,N_18084);
and U21145 (N_21145,N_19690,N_18607);
nand U21146 (N_21146,N_19346,N_18227);
xnor U21147 (N_21147,N_18869,N_18268);
nand U21148 (N_21148,N_19775,N_18191);
or U21149 (N_21149,N_18595,N_18961);
nor U21150 (N_21150,N_19149,N_18143);
nand U21151 (N_21151,N_19663,N_18340);
nand U21152 (N_21152,N_18326,N_19322);
nand U21153 (N_21153,N_19259,N_18298);
nand U21154 (N_21154,N_18354,N_18865);
xor U21155 (N_21155,N_19012,N_18131);
and U21156 (N_21156,N_18830,N_19295);
or U21157 (N_21157,N_19497,N_19403);
xnor U21158 (N_21158,N_18715,N_18323);
or U21159 (N_21159,N_18040,N_19137);
nand U21160 (N_21160,N_19236,N_19553);
and U21161 (N_21161,N_18088,N_18797);
or U21162 (N_21162,N_19548,N_18149);
nand U21163 (N_21163,N_18274,N_19449);
and U21164 (N_21164,N_18699,N_18064);
nand U21165 (N_21165,N_18973,N_19286);
or U21166 (N_21166,N_19541,N_19803);
nand U21167 (N_21167,N_19056,N_18279);
xor U21168 (N_21168,N_19217,N_18857);
nand U21169 (N_21169,N_18808,N_19787);
or U21170 (N_21170,N_19812,N_18940);
and U21171 (N_21171,N_18833,N_19043);
or U21172 (N_21172,N_18967,N_19899);
nor U21173 (N_21173,N_19005,N_19062);
and U21174 (N_21174,N_19618,N_19232);
or U21175 (N_21175,N_18547,N_19965);
nor U21176 (N_21176,N_18046,N_18114);
or U21177 (N_21177,N_18819,N_18720);
nand U21178 (N_21178,N_18108,N_18606);
or U21179 (N_21179,N_19430,N_19828);
nor U21180 (N_21180,N_19798,N_19387);
nor U21181 (N_21181,N_18252,N_18175);
nand U21182 (N_21182,N_18559,N_19798);
xor U21183 (N_21183,N_18094,N_19373);
nand U21184 (N_21184,N_19836,N_18685);
and U21185 (N_21185,N_18194,N_19255);
or U21186 (N_21186,N_19161,N_18684);
or U21187 (N_21187,N_18784,N_19011);
nor U21188 (N_21188,N_18926,N_19396);
nor U21189 (N_21189,N_18427,N_19084);
nor U21190 (N_21190,N_19784,N_19566);
and U21191 (N_21191,N_19309,N_19400);
nand U21192 (N_21192,N_18096,N_19036);
nand U21193 (N_21193,N_18692,N_18487);
or U21194 (N_21194,N_19592,N_19948);
nor U21195 (N_21195,N_18940,N_19326);
and U21196 (N_21196,N_18043,N_19166);
and U21197 (N_21197,N_18147,N_18480);
xnor U21198 (N_21198,N_18341,N_19938);
nand U21199 (N_21199,N_19783,N_18010);
nor U21200 (N_21200,N_19112,N_19483);
or U21201 (N_21201,N_18479,N_19179);
or U21202 (N_21202,N_19489,N_19685);
xor U21203 (N_21203,N_18908,N_19498);
xor U21204 (N_21204,N_19393,N_19890);
xnor U21205 (N_21205,N_18661,N_19812);
and U21206 (N_21206,N_19097,N_19729);
and U21207 (N_21207,N_18702,N_19083);
nor U21208 (N_21208,N_19668,N_18243);
and U21209 (N_21209,N_19097,N_19281);
nor U21210 (N_21210,N_18952,N_18297);
xor U21211 (N_21211,N_19555,N_19608);
nand U21212 (N_21212,N_19674,N_18481);
xor U21213 (N_21213,N_18083,N_18807);
and U21214 (N_21214,N_18308,N_19079);
nand U21215 (N_21215,N_18921,N_18191);
xnor U21216 (N_21216,N_18975,N_18239);
and U21217 (N_21217,N_18186,N_18661);
nor U21218 (N_21218,N_19044,N_19259);
xor U21219 (N_21219,N_18882,N_19921);
nor U21220 (N_21220,N_19836,N_18889);
nor U21221 (N_21221,N_18283,N_18267);
xor U21222 (N_21222,N_18769,N_18153);
or U21223 (N_21223,N_18215,N_19239);
or U21224 (N_21224,N_18169,N_18380);
nand U21225 (N_21225,N_18287,N_19312);
or U21226 (N_21226,N_18968,N_19032);
xor U21227 (N_21227,N_19121,N_18851);
xor U21228 (N_21228,N_19303,N_19260);
and U21229 (N_21229,N_19443,N_19696);
and U21230 (N_21230,N_19050,N_18201);
nand U21231 (N_21231,N_19684,N_18973);
nor U21232 (N_21232,N_19274,N_18111);
or U21233 (N_21233,N_19861,N_19938);
xnor U21234 (N_21234,N_19587,N_19259);
nand U21235 (N_21235,N_19388,N_19410);
and U21236 (N_21236,N_18845,N_19186);
xor U21237 (N_21237,N_18024,N_19369);
nand U21238 (N_21238,N_19981,N_19901);
xor U21239 (N_21239,N_18804,N_19181);
xor U21240 (N_21240,N_18791,N_19944);
nor U21241 (N_21241,N_19109,N_18322);
nor U21242 (N_21242,N_19413,N_18583);
xnor U21243 (N_21243,N_19092,N_18971);
or U21244 (N_21244,N_19549,N_18995);
and U21245 (N_21245,N_18889,N_19557);
and U21246 (N_21246,N_19918,N_18021);
nand U21247 (N_21247,N_19926,N_18316);
nor U21248 (N_21248,N_18058,N_19512);
xor U21249 (N_21249,N_18486,N_19990);
nor U21250 (N_21250,N_19310,N_19792);
and U21251 (N_21251,N_19187,N_18901);
nor U21252 (N_21252,N_19551,N_19401);
nor U21253 (N_21253,N_19693,N_19532);
or U21254 (N_21254,N_18267,N_18780);
xnor U21255 (N_21255,N_19161,N_19272);
xor U21256 (N_21256,N_19871,N_19156);
nand U21257 (N_21257,N_19509,N_18224);
nand U21258 (N_21258,N_18448,N_18682);
or U21259 (N_21259,N_18661,N_18513);
xor U21260 (N_21260,N_19551,N_18670);
nor U21261 (N_21261,N_19000,N_18950);
and U21262 (N_21262,N_19441,N_19113);
and U21263 (N_21263,N_19220,N_19603);
nor U21264 (N_21264,N_18918,N_18387);
xnor U21265 (N_21265,N_19098,N_18366);
xnor U21266 (N_21266,N_19072,N_19719);
xnor U21267 (N_21267,N_19020,N_19691);
nor U21268 (N_21268,N_19523,N_18922);
xor U21269 (N_21269,N_19084,N_18006);
nand U21270 (N_21270,N_19217,N_19712);
xor U21271 (N_21271,N_19100,N_19371);
and U21272 (N_21272,N_18754,N_19810);
nor U21273 (N_21273,N_19502,N_18912);
or U21274 (N_21274,N_18422,N_18237);
nor U21275 (N_21275,N_19134,N_19867);
or U21276 (N_21276,N_19129,N_18211);
xor U21277 (N_21277,N_18725,N_19187);
nand U21278 (N_21278,N_18872,N_19935);
nand U21279 (N_21279,N_18774,N_18050);
nand U21280 (N_21280,N_19300,N_19661);
and U21281 (N_21281,N_18989,N_18027);
nor U21282 (N_21282,N_18211,N_19828);
nand U21283 (N_21283,N_19929,N_18139);
or U21284 (N_21284,N_18154,N_18808);
nand U21285 (N_21285,N_19981,N_19341);
or U21286 (N_21286,N_19420,N_18897);
and U21287 (N_21287,N_18912,N_19662);
nand U21288 (N_21288,N_18256,N_19404);
nor U21289 (N_21289,N_19167,N_18425);
nor U21290 (N_21290,N_19181,N_18523);
nor U21291 (N_21291,N_19060,N_19008);
and U21292 (N_21292,N_19000,N_18302);
and U21293 (N_21293,N_18746,N_19215);
or U21294 (N_21294,N_18268,N_19668);
and U21295 (N_21295,N_19075,N_19428);
and U21296 (N_21296,N_19102,N_18152);
xor U21297 (N_21297,N_19213,N_19856);
and U21298 (N_21298,N_19528,N_18268);
nor U21299 (N_21299,N_18293,N_19764);
nor U21300 (N_21300,N_19237,N_19600);
nor U21301 (N_21301,N_19571,N_18261);
xor U21302 (N_21302,N_18814,N_18586);
nor U21303 (N_21303,N_19811,N_18521);
or U21304 (N_21304,N_18337,N_18058);
and U21305 (N_21305,N_19345,N_19692);
or U21306 (N_21306,N_19930,N_18672);
nand U21307 (N_21307,N_18488,N_19381);
and U21308 (N_21308,N_19343,N_19145);
and U21309 (N_21309,N_18113,N_19236);
or U21310 (N_21310,N_19475,N_18655);
nand U21311 (N_21311,N_18068,N_18984);
nor U21312 (N_21312,N_19757,N_18548);
and U21313 (N_21313,N_18368,N_19431);
nand U21314 (N_21314,N_18091,N_19698);
and U21315 (N_21315,N_19675,N_19876);
nand U21316 (N_21316,N_19256,N_19652);
xnor U21317 (N_21317,N_18929,N_18069);
and U21318 (N_21318,N_18671,N_19865);
xnor U21319 (N_21319,N_18590,N_18253);
and U21320 (N_21320,N_18344,N_19524);
or U21321 (N_21321,N_19470,N_19056);
xnor U21322 (N_21322,N_19694,N_18956);
or U21323 (N_21323,N_19865,N_18515);
xnor U21324 (N_21324,N_19468,N_19035);
nand U21325 (N_21325,N_18645,N_19621);
or U21326 (N_21326,N_18700,N_18901);
or U21327 (N_21327,N_19569,N_19198);
nor U21328 (N_21328,N_19572,N_19354);
or U21329 (N_21329,N_19514,N_19561);
nand U21330 (N_21330,N_18061,N_19503);
nor U21331 (N_21331,N_19566,N_18447);
nand U21332 (N_21332,N_19929,N_18217);
or U21333 (N_21333,N_18697,N_18981);
nand U21334 (N_21334,N_19330,N_18849);
or U21335 (N_21335,N_18302,N_18137);
nor U21336 (N_21336,N_18688,N_18586);
xor U21337 (N_21337,N_19459,N_19145);
xnor U21338 (N_21338,N_19020,N_18738);
nor U21339 (N_21339,N_19109,N_19689);
nor U21340 (N_21340,N_19238,N_19787);
and U21341 (N_21341,N_19832,N_19788);
nor U21342 (N_21342,N_18405,N_18816);
nor U21343 (N_21343,N_19507,N_18843);
or U21344 (N_21344,N_19358,N_19266);
xor U21345 (N_21345,N_19622,N_19632);
nand U21346 (N_21346,N_18717,N_19393);
or U21347 (N_21347,N_18689,N_18548);
and U21348 (N_21348,N_19973,N_18822);
and U21349 (N_21349,N_18832,N_18248);
xor U21350 (N_21350,N_19376,N_19605);
xnor U21351 (N_21351,N_19279,N_19259);
nor U21352 (N_21352,N_18963,N_19931);
or U21353 (N_21353,N_18554,N_18843);
or U21354 (N_21354,N_19314,N_19424);
nand U21355 (N_21355,N_19262,N_18087);
xnor U21356 (N_21356,N_18006,N_18098);
nand U21357 (N_21357,N_19440,N_19303);
xor U21358 (N_21358,N_19989,N_18030);
nand U21359 (N_21359,N_19433,N_19747);
and U21360 (N_21360,N_19277,N_19065);
or U21361 (N_21361,N_19586,N_18139);
or U21362 (N_21362,N_19350,N_18154);
nor U21363 (N_21363,N_19430,N_18616);
xnor U21364 (N_21364,N_19199,N_18492);
xnor U21365 (N_21365,N_18464,N_19752);
or U21366 (N_21366,N_19554,N_18289);
and U21367 (N_21367,N_19008,N_18357);
or U21368 (N_21368,N_18202,N_19672);
xnor U21369 (N_21369,N_18737,N_19267);
nand U21370 (N_21370,N_18699,N_18880);
nand U21371 (N_21371,N_18874,N_19756);
xor U21372 (N_21372,N_19051,N_18530);
xnor U21373 (N_21373,N_19175,N_19369);
and U21374 (N_21374,N_18028,N_18159);
and U21375 (N_21375,N_18564,N_19507);
xor U21376 (N_21376,N_19291,N_18778);
and U21377 (N_21377,N_19523,N_19874);
and U21378 (N_21378,N_19198,N_19670);
and U21379 (N_21379,N_18283,N_19734);
xor U21380 (N_21380,N_19093,N_18926);
or U21381 (N_21381,N_19402,N_19599);
xnor U21382 (N_21382,N_19255,N_19164);
nand U21383 (N_21383,N_19881,N_18273);
and U21384 (N_21384,N_18782,N_19765);
nor U21385 (N_21385,N_19276,N_18063);
nor U21386 (N_21386,N_18648,N_19565);
xor U21387 (N_21387,N_19216,N_19000);
or U21388 (N_21388,N_19968,N_19379);
xor U21389 (N_21389,N_18025,N_18482);
and U21390 (N_21390,N_19190,N_18182);
and U21391 (N_21391,N_18668,N_18780);
or U21392 (N_21392,N_18514,N_18460);
nor U21393 (N_21393,N_19413,N_18274);
nand U21394 (N_21394,N_19997,N_19126);
or U21395 (N_21395,N_19491,N_19720);
and U21396 (N_21396,N_19467,N_18051);
nor U21397 (N_21397,N_18436,N_19312);
xor U21398 (N_21398,N_19163,N_18563);
or U21399 (N_21399,N_18150,N_19235);
nand U21400 (N_21400,N_18096,N_18128);
nor U21401 (N_21401,N_18000,N_18104);
and U21402 (N_21402,N_19283,N_18441);
xor U21403 (N_21403,N_18014,N_18273);
nor U21404 (N_21404,N_19103,N_18785);
or U21405 (N_21405,N_18928,N_18128);
xor U21406 (N_21406,N_19705,N_18413);
xnor U21407 (N_21407,N_19489,N_19770);
or U21408 (N_21408,N_18822,N_19868);
xnor U21409 (N_21409,N_18711,N_18729);
nor U21410 (N_21410,N_19559,N_19087);
nor U21411 (N_21411,N_18630,N_18133);
nor U21412 (N_21412,N_19868,N_19468);
nor U21413 (N_21413,N_19371,N_19543);
or U21414 (N_21414,N_19367,N_19401);
xor U21415 (N_21415,N_18982,N_18673);
and U21416 (N_21416,N_18857,N_19013);
or U21417 (N_21417,N_18309,N_18485);
nand U21418 (N_21418,N_18044,N_18579);
or U21419 (N_21419,N_18758,N_19548);
nor U21420 (N_21420,N_19050,N_18965);
nand U21421 (N_21421,N_19864,N_19883);
and U21422 (N_21422,N_19847,N_18946);
nor U21423 (N_21423,N_19719,N_19156);
and U21424 (N_21424,N_18317,N_19427);
and U21425 (N_21425,N_19939,N_18764);
xnor U21426 (N_21426,N_19654,N_19877);
and U21427 (N_21427,N_19467,N_18502);
or U21428 (N_21428,N_18744,N_19760);
and U21429 (N_21429,N_19060,N_19061);
or U21430 (N_21430,N_19513,N_19326);
or U21431 (N_21431,N_19154,N_19352);
and U21432 (N_21432,N_19657,N_19420);
xnor U21433 (N_21433,N_19391,N_19805);
nand U21434 (N_21434,N_19380,N_19042);
nand U21435 (N_21435,N_19028,N_19424);
nor U21436 (N_21436,N_19914,N_19805);
or U21437 (N_21437,N_18022,N_18869);
and U21438 (N_21438,N_19587,N_18533);
and U21439 (N_21439,N_18303,N_18593);
nor U21440 (N_21440,N_18158,N_18614);
or U21441 (N_21441,N_19188,N_18685);
xnor U21442 (N_21442,N_18462,N_18347);
xor U21443 (N_21443,N_18901,N_19627);
and U21444 (N_21444,N_19868,N_18640);
and U21445 (N_21445,N_19384,N_19994);
xor U21446 (N_21446,N_19075,N_19688);
xor U21447 (N_21447,N_19161,N_19447);
xor U21448 (N_21448,N_19619,N_18820);
nand U21449 (N_21449,N_18314,N_18156);
xnor U21450 (N_21450,N_18713,N_18560);
nand U21451 (N_21451,N_18760,N_18627);
or U21452 (N_21452,N_18122,N_19435);
nand U21453 (N_21453,N_19265,N_18806);
and U21454 (N_21454,N_18123,N_19615);
nand U21455 (N_21455,N_18649,N_19904);
and U21456 (N_21456,N_18917,N_18298);
and U21457 (N_21457,N_19553,N_18729);
nor U21458 (N_21458,N_19433,N_18906);
and U21459 (N_21459,N_19170,N_19285);
nor U21460 (N_21460,N_19735,N_18049);
and U21461 (N_21461,N_18822,N_18621);
nand U21462 (N_21462,N_18548,N_18241);
and U21463 (N_21463,N_19539,N_18257);
nand U21464 (N_21464,N_19694,N_19254);
or U21465 (N_21465,N_19134,N_19362);
nor U21466 (N_21466,N_18827,N_19529);
and U21467 (N_21467,N_18768,N_19919);
or U21468 (N_21468,N_19427,N_19406);
nor U21469 (N_21469,N_19556,N_18073);
and U21470 (N_21470,N_18910,N_18608);
nand U21471 (N_21471,N_19636,N_19182);
or U21472 (N_21472,N_19677,N_18908);
nand U21473 (N_21473,N_19704,N_18506);
xnor U21474 (N_21474,N_18295,N_19805);
nor U21475 (N_21475,N_18295,N_19485);
or U21476 (N_21476,N_19190,N_18405);
nand U21477 (N_21477,N_18680,N_18632);
nand U21478 (N_21478,N_18024,N_19459);
or U21479 (N_21479,N_18072,N_19495);
xor U21480 (N_21480,N_18169,N_19202);
nor U21481 (N_21481,N_19074,N_19417);
nand U21482 (N_21482,N_18969,N_19295);
nor U21483 (N_21483,N_18251,N_19227);
nor U21484 (N_21484,N_19026,N_19622);
nor U21485 (N_21485,N_19536,N_19415);
or U21486 (N_21486,N_18405,N_19035);
and U21487 (N_21487,N_18118,N_18103);
xor U21488 (N_21488,N_19232,N_18844);
nor U21489 (N_21489,N_19035,N_19866);
nand U21490 (N_21490,N_18667,N_18080);
and U21491 (N_21491,N_19173,N_19150);
nor U21492 (N_21492,N_18353,N_18154);
and U21493 (N_21493,N_19594,N_19874);
and U21494 (N_21494,N_19248,N_18359);
or U21495 (N_21495,N_18889,N_18176);
nand U21496 (N_21496,N_19081,N_18063);
nand U21497 (N_21497,N_18817,N_19585);
xor U21498 (N_21498,N_19064,N_18591);
nor U21499 (N_21499,N_18250,N_18274);
or U21500 (N_21500,N_18579,N_19512);
nor U21501 (N_21501,N_18397,N_19479);
and U21502 (N_21502,N_19027,N_18960);
xnor U21503 (N_21503,N_19539,N_19052);
nand U21504 (N_21504,N_19074,N_19723);
xnor U21505 (N_21505,N_18501,N_18686);
xor U21506 (N_21506,N_19954,N_18513);
nand U21507 (N_21507,N_18417,N_19523);
nor U21508 (N_21508,N_18689,N_19105);
nor U21509 (N_21509,N_19541,N_18302);
xor U21510 (N_21510,N_19798,N_18425);
and U21511 (N_21511,N_18113,N_19522);
nor U21512 (N_21512,N_19498,N_19448);
nor U21513 (N_21513,N_18546,N_19697);
nor U21514 (N_21514,N_19070,N_19673);
nand U21515 (N_21515,N_18983,N_19634);
xor U21516 (N_21516,N_18031,N_18736);
and U21517 (N_21517,N_18267,N_18460);
xnor U21518 (N_21518,N_19094,N_18446);
nor U21519 (N_21519,N_19327,N_19568);
and U21520 (N_21520,N_18743,N_18441);
nand U21521 (N_21521,N_18975,N_18605);
nor U21522 (N_21522,N_18994,N_19000);
nor U21523 (N_21523,N_19796,N_19711);
nand U21524 (N_21524,N_19783,N_19965);
and U21525 (N_21525,N_18709,N_18508);
xor U21526 (N_21526,N_18613,N_18832);
nand U21527 (N_21527,N_19957,N_19008);
and U21528 (N_21528,N_19363,N_19958);
xnor U21529 (N_21529,N_19669,N_19895);
or U21530 (N_21530,N_19076,N_18236);
nand U21531 (N_21531,N_19092,N_18260);
nor U21532 (N_21532,N_18258,N_19903);
xor U21533 (N_21533,N_18021,N_19581);
nand U21534 (N_21534,N_18565,N_19611);
or U21535 (N_21535,N_19407,N_19011);
or U21536 (N_21536,N_19690,N_19278);
xnor U21537 (N_21537,N_19821,N_18237);
and U21538 (N_21538,N_19261,N_19114);
and U21539 (N_21539,N_18068,N_18965);
or U21540 (N_21540,N_18166,N_19982);
xnor U21541 (N_21541,N_18294,N_18992);
or U21542 (N_21542,N_18221,N_18296);
and U21543 (N_21543,N_19511,N_19220);
and U21544 (N_21544,N_18285,N_18690);
nand U21545 (N_21545,N_19338,N_18730);
and U21546 (N_21546,N_18544,N_18341);
nand U21547 (N_21547,N_19961,N_18391);
nand U21548 (N_21548,N_19707,N_18314);
nand U21549 (N_21549,N_18152,N_18507);
and U21550 (N_21550,N_18954,N_18085);
and U21551 (N_21551,N_18081,N_19605);
and U21552 (N_21552,N_19093,N_18889);
nor U21553 (N_21553,N_18925,N_18800);
and U21554 (N_21554,N_18743,N_18781);
xnor U21555 (N_21555,N_18729,N_18599);
nand U21556 (N_21556,N_19068,N_19174);
and U21557 (N_21557,N_18399,N_18466);
and U21558 (N_21558,N_18917,N_19464);
or U21559 (N_21559,N_18165,N_19628);
or U21560 (N_21560,N_19533,N_19398);
xnor U21561 (N_21561,N_19056,N_18164);
and U21562 (N_21562,N_19476,N_18546);
and U21563 (N_21563,N_19540,N_19024);
nand U21564 (N_21564,N_19175,N_19430);
nand U21565 (N_21565,N_19255,N_19081);
nor U21566 (N_21566,N_19652,N_19853);
or U21567 (N_21567,N_19494,N_18105);
nor U21568 (N_21568,N_18981,N_19616);
nor U21569 (N_21569,N_18837,N_18240);
and U21570 (N_21570,N_18247,N_18767);
nor U21571 (N_21571,N_18510,N_18495);
and U21572 (N_21572,N_18175,N_19539);
nand U21573 (N_21573,N_19438,N_19713);
or U21574 (N_21574,N_19431,N_19219);
nand U21575 (N_21575,N_19156,N_19595);
or U21576 (N_21576,N_19344,N_19910);
or U21577 (N_21577,N_18003,N_19522);
and U21578 (N_21578,N_18113,N_19965);
nor U21579 (N_21579,N_18783,N_19872);
nand U21580 (N_21580,N_18492,N_19435);
nand U21581 (N_21581,N_18796,N_18581);
xor U21582 (N_21582,N_18989,N_18541);
nor U21583 (N_21583,N_18653,N_18072);
nor U21584 (N_21584,N_18196,N_19395);
xor U21585 (N_21585,N_19366,N_18879);
xor U21586 (N_21586,N_19528,N_19840);
xor U21587 (N_21587,N_19959,N_18302);
or U21588 (N_21588,N_18618,N_19939);
nor U21589 (N_21589,N_18369,N_18970);
and U21590 (N_21590,N_19331,N_19860);
and U21591 (N_21591,N_19020,N_19663);
or U21592 (N_21592,N_18078,N_19218);
xor U21593 (N_21593,N_19716,N_19517);
and U21594 (N_21594,N_19988,N_19808);
xor U21595 (N_21595,N_19025,N_19755);
or U21596 (N_21596,N_18746,N_19257);
nor U21597 (N_21597,N_19407,N_18003);
or U21598 (N_21598,N_19164,N_19146);
xnor U21599 (N_21599,N_19512,N_19747);
xor U21600 (N_21600,N_18780,N_18223);
nor U21601 (N_21601,N_18860,N_18394);
nor U21602 (N_21602,N_19021,N_18555);
nand U21603 (N_21603,N_19121,N_19088);
xor U21604 (N_21604,N_18706,N_18195);
or U21605 (N_21605,N_18012,N_18537);
nor U21606 (N_21606,N_18908,N_19451);
or U21607 (N_21607,N_19578,N_18123);
xnor U21608 (N_21608,N_19141,N_19991);
or U21609 (N_21609,N_19690,N_18308);
nand U21610 (N_21610,N_18045,N_18166);
xnor U21611 (N_21611,N_19863,N_19951);
and U21612 (N_21612,N_19686,N_19099);
xor U21613 (N_21613,N_19498,N_19941);
and U21614 (N_21614,N_19166,N_18769);
and U21615 (N_21615,N_19864,N_18291);
or U21616 (N_21616,N_18343,N_19496);
or U21617 (N_21617,N_18847,N_19457);
nand U21618 (N_21618,N_19184,N_19433);
nand U21619 (N_21619,N_19941,N_18602);
or U21620 (N_21620,N_19768,N_19394);
nor U21621 (N_21621,N_19486,N_19598);
and U21622 (N_21622,N_18726,N_18141);
nor U21623 (N_21623,N_18545,N_18577);
or U21624 (N_21624,N_19335,N_18519);
nand U21625 (N_21625,N_19865,N_19482);
nor U21626 (N_21626,N_19144,N_18708);
nand U21627 (N_21627,N_18822,N_18739);
and U21628 (N_21628,N_18568,N_19223);
and U21629 (N_21629,N_18976,N_19928);
and U21630 (N_21630,N_18578,N_18656);
xor U21631 (N_21631,N_18094,N_18255);
xor U21632 (N_21632,N_18923,N_18456);
nor U21633 (N_21633,N_18787,N_19461);
or U21634 (N_21634,N_18934,N_18793);
nand U21635 (N_21635,N_18153,N_19241);
nor U21636 (N_21636,N_19364,N_18489);
nand U21637 (N_21637,N_19980,N_18193);
nand U21638 (N_21638,N_19605,N_18096);
and U21639 (N_21639,N_19518,N_19763);
xor U21640 (N_21640,N_18243,N_18477);
nand U21641 (N_21641,N_18194,N_18369);
and U21642 (N_21642,N_18727,N_19609);
xor U21643 (N_21643,N_19360,N_19058);
nor U21644 (N_21644,N_19363,N_18413);
nor U21645 (N_21645,N_18010,N_19717);
xnor U21646 (N_21646,N_19388,N_18270);
nand U21647 (N_21647,N_18124,N_18427);
nand U21648 (N_21648,N_19201,N_19418);
nor U21649 (N_21649,N_19378,N_18016);
or U21650 (N_21650,N_18314,N_19933);
or U21651 (N_21651,N_19520,N_18097);
nand U21652 (N_21652,N_18024,N_19942);
or U21653 (N_21653,N_19394,N_19601);
and U21654 (N_21654,N_19913,N_18945);
xor U21655 (N_21655,N_18748,N_19558);
nor U21656 (N_21656,N_19755,N_19977);
and U21657 (N_21657,N_19518,N_18171);
nor U21658 (N_21658,N_19140,N_18712);
or U21659 (N_21659,N_18163,N_18740);
nand U21660 (N_21660,N_18217,N_19202);
xor U21661 (N_21661,N_18119,N_19014);
or U21662 (N_21662,N_18216,N_19445);
nor U21663 (N_21663,N_18198,N_18443);
and U21664 (N_21664,N_19345,N_18323);
nand U21665 (N_21665,N_18128,N_18651);
or U21666 (N_21666,N_18905,N_18828);
xnor U21667 (N_21667,N_18434,N_19094);
or U21668 (N_21668,N_18967,N_18990);
xnor U21669 (N_21669,N_18966,N_19259);
nand U21670 (N_21670,N_18246,N_18652);
nor U21671 (N_21671,N_18727,N_18338);
xnor U21672 (N_21672,N_18476,N_18992);
xor U21673 (N_21673,N_19817,N_18069);
xnor U21674 (N_21674,N_18584,N_19641);
and U21675 (N_21675,N_18146,N_19290);
or U21676 (N_21676,N_18421,N_18123);
nand U21677 (N_21677,N_19996,N_19428);
and U21678 (N_21678,N_19330,N_19737);
and U21679 (N_21679,N_18711,N_18087);
xor U21680 (N_21680,N_18444,N_18454);
or U21681 (N_21681,N_18986,N_18084);
or U21682 (N_21682,N_18305,N_19427);
nand U21683 (N_21683,N_19200,N_19618);
nor U21684 (N_21684,N_18013,N_18300);
xnor U21685 (N_21685,N_19014,N_19364);
nand U21686 (N_21686,N_19765,N_18137);
nand U21687 (N_21687,N_19964,N_18372);
nor U21688 (N_21688,N_18336,N_19192);
nor U21689 (N_21689,N_19116,N_18140);
nand U21690 (N_21690,N_18178,N_19225);
or U21691 (N_21691,N_18138,N_18890);
and U21692 (N_21692,N_19573,N_19818);
nand U21693 (N_21693,N_18880,N_18787);
xor U21694 (N_21694,N_18737,N_19547);
nand U21695 (N_21695,N_19350,N_19121);
xor U21696 (N_21696,N_18041,N_19974);
nand U21697 (N_21697,N_19610,N_18017);
and U21698 (N_21698,N_19072,N_19050);
xnor U21699 (N_21699,N_18932,N_18576);
and U21700 (N_21700,N_19446,N_19899);
or U21701 (N_21701,N_18553,N_19045);
nor U21702 (N_21702,N_19642,N_18959);
nand U21703 (N_21703,N_19409,N_18658);
or U21704 (N_21704,N_19463,N_19954);
nand U21705 (N_21705,N_19516,N_19112);
or U21706 (N_21706,N_19821,N_18103);
and U21707 (N_21707,N_18826,N_18848);
nor U21708 (N_21708,N_19294,N_18334);
and U21709 (N_21709,N_19514,N_19760);
nand U21710 (N_21710,N_19400,N_19500);
and U21711 (N_21711,N_18154,N_18980);
nand U21712 (N_21712,N_18425,N_18350);
and U21713 (N_21713,N_19724,N_19290);
xor U21714 (N_21714,N_18630,N_18093);
nand U21715 (N_21715,N_18525,N_18511);
xor U21716 (N_21716,N_18526,N_18559);
and U21717 (N_21717,N_18854,N_19487);
nand U21718 (N_21718,N_19227,N_18800);
xnor U21719 (N_21719,N_19956,N_18942);
nand U21720 (N_21720,N_19190,N_18364);
xor U21721 (N_21721,N_19272,N_19944);
and U21722 (N_21722,N_18318,N_19939);
nand U21723 (N_21723,N_18029,N_18448);
xnor U21724 (N_21724,N_19206,N_18061);
or U21725 (N_21725,N_19523,N_18937);
xor U21726 (N_21726,N_19476,N_19753);
and U21727 (N_21727,N_18655,N_18513);
and U21728 (N_21728,N_19441,N_19282);
nor U21729 (N_21729,N_18803,N_19846);
and U21730 (N_21730,N_19812,N_19608);
and U21731 (N_21731,N_19005,N_19917);
nor U21732 (N_21732,N_19381,N_19521);
nor U21733 (N_21733,N_18425,N_19457);
nand U21734 (N_21734,N_18140,N_18073);
xor U21735 (N_21735,N_18219,N_19702);
xnor U21736 (N_21736,N_18082,N_19749);
xnor U21737 (N_21737,N_19055,N_18359);
nand U21738 (N_21738,N_19018,N_18167);
nor U21739 (N_21739,N_18080,N_19979);
or U21740 (N_21740,N_19421,N_19564);
or U21741 (N_21741,N_19320,N_19300);
or U21742 (N_21742,N_18289,N_18922);
nand U21743 (N_21743,N_18551,N_18359);
nand U21744 (N_21744,N_19778,N_18421);
and U21745 (N_21745,N_19612,N_18326);
nand U21746 (N_21746,N_19425,N_18256);
xnor U21747 (N_21747,N_18958,N_18818);
nand U21748 (N_21748,N_19297,N_18236);
or U21749 (N_21749,N_19330,N_18516);
and U21750 (N_21750,N_18310,N_19213);
and U21751 (N_21751,N_19169,N_18218);
and U21752 (N_21752,N_19948,N_18081);
and U21753 (N_21753,N_19599,N_19970);
xor U21754 (N_21754,N_18834,N_19438);
nor U21755 (N_21755,N_18740,N_18283);
nor U21756 (N_21756,N_19630,N_19036);
xnor U21757 (N_21757,N_18159,N_18907);
xor U21758 (N_21758,N_19183,N_18852);
and U21759 (N_21759,N_19743,N_19659);
nor U21760 (N_21760,N_19255,N_18846);
or U21761 (N_21761,N_18890,N_18905);
nor U21762 (N_21762,N_18981,N_19206);
nor U21763 (N_21763,N_18736,N_18085);
nand U21764 (N_21764,N_19720,N_18238);
and U21765 (N_21765,N_18471,N_18314);
nor U21766 (N_21766,N_18467,N_19580);
or U21767 (N_21767,N_19405,N_18067);
xnor U21768 (N_21768,N_19249,N_18577);
nand U21769 (N_21769,N_19836,N_19742);
nand U21770 (N_21770,N_19757,N_19622);
and U21771 (N_21771,N_18838,N_18359);
nor U21772 (N_21772,N_18321,N_19309);
and U21773 (N_21773,N_19044,N_18729);
or U21774 (N_21774,N_19696,N_18866);
and U21775 (N_21775,N_19188,N_18663);
and U21776 (N_21776,N_18284,N_19516);
xnor U21777 (N_21777,N_19356,N_19133);
xnor U21778 (N_21778,N_19609,N_18378);
and U21779 (N_21779,N_19095,N_18173);
nand U21780 (N_21780,N_19411,N_19103);
or U21781 (N_21781,N_18086,N_19456);
xnor U21782 (N_21782,N_19242,N_18674);
and U21783 (N_21783,N_18994,N_19649);
nor U21784 (N_21784,N_18370,N_19437);
and U21785 (N_21785,N_18659,N_18180);
nand U21786 (N_21786,N_19002,N_19195);
and U21787 (N_21787,N_18760,N_18899);
xnor U21788 (N_21788,N_19610,N_19893);
xor U21789 (N_21789,N_19057,N_19124);
nand U21790 (N_21790,N_19627,N_19098);
and U21791 (N_21791,N_18521,N_19466);
nor U21792 (N_21792,N_19065,N_19726);
nand U21793 (N_21793,N_19737,N_19388);
and U21794 (N_21794,N_18245,N_18481);
xor U21795 (N_21795,N_18580,N_18621);
or U21796 (N_21796,N_19333,N_19810);
nor U21797 (N_21797,N_18250,N_19935);
and U21798 (N_21798,N_19614,N_19931);
xor U21799 (N_21799,N_18009,N_18952);
nand U21800 (N_21800,N_18607,N_18683);
nand U21801 (N_21801,N_18106,N_19775);
nand U21802 (N_21802,N_19282,N_18500);
and U21803 (N_21803,N_18716,N_18461);
nand U21804 (N_21804,N_19177,N_18255);
nor U21805 (N_21805,N_18888,N_18821);
or U21806 (N_21806,N_18331,N_19850);
or U21807 (N_21807,N_18892,N_18213);
xnor U21808 (N_21808,N_18946,N_19589);
and U21809 (N_21809,N_18736,N_18655);
nand U21810 (N_21810,N_18111,N_18743);
xor U21811 (N_21811,N_19717,N_19176);
or U21812 (N_21812,N_19903,N_18832);
and U21813 (N_21813,N_18916,N_18471);
and U21814 (N_21814,N_19609,N_18506);
nor U21815 (N_21815,N_19719,N_18949);
nor U21816 (N_21816,N_19616,N_19956);
xor U21817 (N_21817,N_19437,N_18525);
and U21818 (N_21818,N_19768,N_19252);
nor U21819 (N_21819,N_18550,N_19268);
or U21820 (N_21820,N_19196,N_18904);
and U21821 (N_21821,N_18940,N_19686);
nor U21822 (N_21822,N_18799,N_18010);
nor U21823 (N_21823,N_19837,N_18992);
nand U21824 (N_21824,N_19946,N_18560);
xnor U21825 (N_21825,N_18773,N_18482);
nand U21826 (N_21826,N_18686,N_19384);
and U21827 (N_21827,N_19709,N_18624);
and U21828 (N_21828,N_19052,N_18572);
xor U21829 (N_21829,N_18090,N_18801);
or U21830 (N_21830,N_19964,N_18089);
and U21831 (N_21831,N_18647,N_19878);
xnor U21832 (N_21832,N_19231,N_19253);
nand U21833 (N_21833,N_19178,N_18309);
nor U21834 (N_21834,N_19987,N_19804);
and U21835 (N_21835,N_19768,N_19265);
nand U21836 (N_21836,N_19537,N_19657);
nor U21837 (N_21837,N_19461,N_18841);
nand U21838 (N_21838,N_19139,N_18603);
or U21839 (N_21839,N_19525,N_19853);
nor U21840 (N_21840,N_18496,N_18344);
nor U21841 (N_21841,N_18314,N_19074);
nand U21842 (N_21842,N_19374,N_18420);
and U21843 (N_21843,N_18550,N_18157);
or U21844 (N_21844,N_19786,N_18193);
xnor U21845 (N_21845,N_18675,N_19988);
or U21846 (N_21846,N_18243,N_19542);
xnor U21847 (N_21847,N_19886,N_18143);
and U21848 (N_21848,N_19626,N_18012);
or U21849 (N_21849,N_19106,N_19839);
nand U21850 (N_21850,N_19081,N_19896);
nand U21851 (N_21851,N_18160,N_18633);
nor U21852 (N_21852,N_18131,N_19774);
or U21853 (N_21853,N_18171,N_18944);
xor U21854 (N_21854,N_18709,N_19333);
xnor U21855 (N_21855,N_18210,N_18665);
xor U21856 (N_21856,N_18651,N_18522);
xor U21857 (N_21857,N_18722,N_19453);
nand U21858 (N_21858,N_18351,N_19931);
xor U21859 (N_21859,N_19704,N_19142);
or U21860 (N_21860,N_18393,N_19158);
and U21861 (N_21861,N_18248,N_19988);
xnor U21862 (N_21862,N_19215,N_18989);
nand U21863 (N_21863,N_18779,N_18062);
nor U21864 (N_21864,N_19210,N_18607);
nand U21865 (N_21865,N_19454,N_18945);
or U21866 (N_21866,N_18096,N_19606);
xnor U21867 (N_21867,N_19019,N_18934);
nand U21868 (N_21868,N_18160,N_19710);
nor U21869 (N_21869,N_18761,N_19684);
nor U21870 (N_21870,N_19187,N_18958);
and U21871 (N_21871,N_19655,N_18912);
nor U21872 (N_21872,N_19091,N_18970);
nand U21873 (N_21873,N_18835,N_19413);
nand U21874 (N_21874,N_18658,N_19842);
xor U21875 (N_21875,N_19967,N_19140);
nor U21876 (N_21876,N_18450,N_18344);
and U21877 (N_21877,N_19900,N_18018);
or U21878 (N_21878,N_19611,N_18108);
nand U21879 (N_21879,N_18761,N_19543);
nand U21880 (N_21880,N_19391,N_19138);
nand U21881 (N_21881,N_18939,N_18061);
nand U21882 (N_21882,N_19228,N_19609);
nand U21883 (N_21883,N_19413,N_18425);
and U21884 (N_21884,N_18826,N_19543);
nand U21885 (N_21885,N_19476,N_18612);
or U21886 (N_21886,N_19397,N_19413);
nand U21887 (N_21887,N_18401,N_18706);
or U21888 (N_21888,N_18828,N_18283);
xnor U21889 (N_21889,N_18650,N_18285);
or U21890 (N_21890,N_18674,N_18450);
or U21891 (N_21891,N_18310,N_19072);
and U21892 (N_21892,N_18088,N_18450);
nand U21893 (N_21893,N_18127,N_19345);
and U21894 (N_21894,N_19356,N_19655);
nor U21895 (N_21895,N_18837,N_18783);
nand U21896 (N_21896,N_19380,N_18466);
nor U21897 (N_21897,N_18304,N_19679);
or U21898 (N_21898,N_18138,N_19953);
nor U21899 (N_21899,N_19614,N_18296);
xor U21900 (N_21900,N_18387,N_18990);
nor U21901 (N_21901,N_19639,N_19016);
xnor U21902 (N_21902,N_19689,N_18483);
xor U21903 (N_21903,N_19915,N_18777);
xnor U21904 (N_21904,N_19351,N_19225);
or U21905 (N_21905,N_18207,N_19149);
nand U21906 (N_21906,N_19184,N_19344);
nor U21907 (N_21907,N_19576,N_19997);
nor U21908 (N_21908,N_18269,N_19712);
xnor U21909 (N_21909,N_19065,N_18913);
or U21910 (N_21910,N_18316,N_19278);
or U21911 (N_21911,N_18309,N_18273);
nor U21912 (N_21912,N_18277,N_19967);
and U21913 (N_21913,N_18203,N_18192);
and U21914 (N_21914,N_19076,N_18289);
or U21915 (N_21915,N_18638,N_18024);
and U21916 (N_21916,N_18945,N_18246);
nand U21917 (N_21917,N_19288,N_19372);
nand U21918 (N_21918,N_18923,N_18780);
or U21919 (N_21919,N_18592,N_18757);
xor U21920 (N_21920,N_19195,N_19142);
or U21921 (N_21921,N_19315,N_19850);
xnor U21922 (N_21922,N_19694,N_18023);
nand U21923 (N_21923,N_18207,N_19376);
nand U21924 (N_21924,N_18145,N_19718);
and U21925 (N_21925,N_19134,N_19572);
and U21926 (N_21926,N_19628,N_18885);
nand U21927 (N_21927,N_19907,N_19336);
nand U21928 (N_21928,N_19299,N_19867);
or U21929 (N_21929,N_19921,N_18061);
nand U21930 (N_21930,N_18813,N_18186);
and U21931 (N_21931,N_19789,N_18458);
and U21932 (N_21932,N_19410,N_19667);
and U21933 (N_21933,N_19211,N_19538);
and U21934 (N_21934,N_18832,N_18450);
xnor U21935 (N_21935,N_18736,N_19551);
nand U21936 (N_21936,N_19536,N_18308);
or U21937 (N_21937,N_18318,N_18488);
nand U21938 (N_21938,N_18512,N_19179);
and U21939 (N_21939,N_19662,N_19624);
xor U21940 (N_21940,N_18618,N_19022);
nor U21941 (N_21941,N_18803,N_19543);
and U21942 (N_21942,N_19876,N_18704);
nor U21943 (N_21943,N_18597,N_19358);
xnor U21944 (N_21944,N_19698,N_18780);
xor U21945 (N_21945,N_18710,N_19025);
nand U21946 (N_21946,N_18065,N_18362);
xnor U21947 (N_21947,N_19910,N_19357);
xnor U21948 (N_21948,N_19796,N_19259);
nand U21949 (N_21949,N_19539,N_19350);
or U21950 (N_21950,N_18237,N_18803);
and U21951 (N_21951,N_18807,N_18750);
nand U21952 (N_21952,N_19871,N_18409);
and U21953 (N_21953,N_19641,N_18114);
and U21954 (N_21954,N_19273,N_18383);
or U21955 (N_21955,N_18809,N_19308);
nand U21956 (N_21956,N_19215,N_19803);
xnor U21957 (N_21957,N_18426,N_19159);
xor U21958 (N_21958,N_18590,N_19901);
nand U21959 (N_21959,N_18583,N_19360);
and U21960 (N_21960,N_19149,N_18738);
xnor U21961 (N_21961,N_19759,N_18170);
nand U21962 (N_21962,N_19122,N_18145);
and U21963 (N_21963,N_18954,N_18672);
and U21964 (N_21964,N_18932,N_19065);
nor U21965 (N_21965,N_18047,N_18974);
or U21966 (N_21966,N_18528,N_19575);
and U21967 (N_21967,N_19866,N_18784);
or U21968 (N_21968,N_18409,N_18476);
nor U21969 (N_21969,N_18513,N_19360);
nand U21970 (N_21970,N_18677,N_19972);
nand U21971 (N_21971,N_18197,N_19131);
and U21972 (N_21972,N_18952,N_19374);
xnor U21973 (N_21973,N_18479,N_18402);
nor U21974 (N_21974,N_19975,N_19756);
and U21975 (N_21975,N_18787,N_19226);
or U21976 (N_21976,N_18973,N_19840);
or U21977 (N_21977,N_18035,N_19619);
nor U21978 (N_21978,N_18471,N_19566);
or U21979 (N_21979,N_19010,N_18978);
or U21980 (N_21980,N_18205,N_18053);
xnor U21981 (N_21981,N_18693,N_18489);
xnor U21982 (N_21982,N_19081,N_18738);
nor U21983 (N_21983,N_18341,N_18240);
nor U21984 (N_21984,N_18423,N_18050);
xnor U21985 (N_21985,N_18519,N_19199);
nand U21986 (N_21986,N_19207,N_19988);
nor U21987 (N_21987,N_19547,N_18458);
nor U21988 (N_21988,N_18711,N_19288);
nor U21989 (N_21989,N_19530,N_19141);
nor U21990 (N_21990,N_18407,N_18065);
xor U21991 (N_21991,N_18920,N_19275);
or U21992 (N_21992,N_19048,N_19657);
xnor U21993 (N_21993,N_19601,N_18458);
nor U21994 (N_21994,N_18048,N_18868);
and U21995 (N_21995,N_18437,N_18392);
xor U21996 (N_21996,N_19356,N_19394);
or U21997 (N_21997,N_18367,N_18872);
nor U21998 (N_21998,N_18498,N_19099);
or U21999 (N_21999,N_18981,N_18565);
and U22000 (N_22000,N_21734,N_20438);
nor U22001 (N_22001,N_20887,N_21123);
nand U22002 (N_22002,N_20322,N_21494);
and U22003 (N_22003,N_20090,N_21896);
or U22004 (N_22004,N_20633,N_21650);
xor U22005 (N_22005,N_21897,N_21413);
nor U22006 (N_22006,N_20965,N_21879);
or U22007 (N_22007,N_21213,N_20646);
nand U22008 (N_22008,N_20132,N_21893);
or U22009 (N_22009,N_20597,N_20666);
xor U22010 (N_22010,N_20324,N_20863);
xor U22011 (N_22011,N_21041,N_20535);
or U22012 (N_22012,N_20081,N_20546);
nor U22013 (N_22013,N_21304,N_20967);
xor U22014 (N_22014,N_21515,N_20102);
or U22015 (N_22015,N_21699,N_21384);
or U22016 (N_22016,N_20695,N_21627);
nor U22017 (N_22017,N_21722,N_21560);
nor U22018 (N_22018,N_20983,N_21276);
xor U22019 (N_22019,N_21605,N_21505);
and U22020 (N_22020,N_20248,N_21883);
or U22021 (N_22021,N_21323,N_21656);
nor U22022 (N_22022,N_21755,N_21575);
xor U22023 (N_22023,N_20408,N_20947);
and U22024 (N_22024,N_21369,N_20083);
nand U22025 (N_22025,N_21490,N_20871);
and U22026 (N_22026,N_21001,N_21710);
nand U22027 (N_22027,N_20714,N_20501);
xnor U22028 (N_22028,N_20037,N_21085);
xnor U22029 (N_22029,N_20593,N_21353);
or U22030 (N_22030,N_21137,N_21887);
nor U22031 (N_22031,N_21818,N_20832);
xor U22032 (N_22032,N_20946,N_20620);
nand U22033 (N_22033,N_20259,N_21367);
and U22034 (N_22034,N_20054,N_20909);
nand U22035 (N_22035,N_20530,N_21519);
nand U22036 (N_22036,N_20139,N_21685);
nand U22037 (N_22037,N_20389,N_20064);
and U22038 (N_22038,N_21581,N_21923);
nand U22039 (N_22039,N_21348,N_20131);
nand U22040 (N_22040,N_20708,N_20249);
nor U22041 (N_22041,N_20799,N_20920);
nor U22042 (N_22042,N_21529,N_20932);
and U22043 (N_22043,N_20521,N_20686);
and U22044 (N_22044,N_20532,N_21217);
xnor U22045 (N_22045,N_20283,N_20464);
or U22046 (N_22046,N_21791,N_20097);
xor U22047 (N_22047,N_20539,N_21470);
or U22048 (N_22048,N_21872,N_21527);
nand U22049 (N_22049,N_21174,N_21767);
and U22050 (N_22050,N_21759,N_20450);
nand U22051 (N_22051,N_21107,N_20281);
or U22052 (N_22052,N_20527,N_21064);
nor U22053 (N_22053,N_20637,N_21951);
and U22054 (N_22054,N_21315,N_21044);
nand U22055 (N_22055,N_21545,N_20827);
or U22056 (N_22056,N_20570,N_20246);
and U22057 (N_22057,N_20219,N_20505);
nand U22058 (N_22058,N_21007,N_21212);
xor U22059 (N_22059,N_20923,N_20460);
or U22060 (N_22060,N_20895,N_21956);
xor U22061 (N_22061,N_20301,N_20892);
xnor U22062 (N_22062,N_20373,N_20607);
or U22063 (N_22063,N_20158,N_21113);
and U22064 (N_22064,N_20021,N_20228);
xnor U22065 (N_22065,N_21145,N_20297);
nand U22066 (N_22066,N_21664,N_21018);
nor U22067 (N_22067,N_21160,N_21294);
or U22068 (N_22068,N_20344,N_21155);
nor U22069 (N_22069,N_20733,N_21378);
nor U22070 (N_22070,N_21686,N_21124);
nor U22071 (N_22071,N_21610,N_20856);
xor U22072 (N_22072,N_20067,N_21130);
xnor U22073 (N_22073,N_21885,N_21537);
and U22074 (N_22074,N_20626,N_21719);
nand U22075 (N_22075,N_21478,N_21332);
nor U22076 (N_22076,N_20578,N_21159);
xnor U22077 (N_22077,N_21894,N_20515);
nand U22078 (N_22078,N_21031,N_21059);
or U22079 (N_22079,N_20769,N_21015);
xnor U22080 (N_22080,N_21587,N_21307);
nand U22081 (N_22081,N_20512,N_20860);
nand U22082 (N_22082,N_20970,N_21637);
nor U22083 (N_22083,N_20365,N_21356);
xor U22084 (N_22084,N_21850,N_21943);
or U22085 (N_22085,N_20788,N_20013);
xor U22086 (N_22086,N_20968,N_20507);
nor U22087 (N_22087,N_20017,N_21114);
nor U22088 (N_22088,N_20142,N_21436);
or U22089 (N_22089,N_21689,N_21225);
xnor U22090 (N_22090,N_20767,N_20332);
xnor U22091 (N_22091,N_21272,N_20598);
and U22092 (N_22092,N_21981,N_21659);
or U22093 (N_22093,N_21351,N_20615);
and U22094 (N_22094,N_20202,N_21401);
or U22095 (N_22095,N_21669,N_21028);
or U22096 (N_22096,N_20234,N_21405);
xor U22097 (N_22097,N_21191,N_21034);
or U22098 (N_22098,N_20904,N_21100);
or U22099 (N_22099,N_20777,N_20200);
nor U22100 (N_22100,N_20048,N_21329);
nor U22101 (N_22101,N_21717,N_20729);
and U22102 (N_22102,N_21520,N_21625);
nor U22103 (N_22103,N_20610,N_21188);
xnor U22104 (N_22104,N_21649,N_20979);
nor U22105 (N_22105,N_20541,N_21565);
xnor U22106 (N_22106,N_20095,N_21492);
or U22107 (N_22107,N_21542,N_21088);
xor U22108 (N_22108,N_21810,N_21877);
and U22109 (N_22109,N_21864,N_20263);
and U22110 (N_22110,N_21517,N_20785);
nor U22111 (N_22111,N_20820,N_20872);
xor U22112 (N_22112,N_21661,N_20543);
nor U22113 (N_22113,N_20415,N_20999);
nand U22114 (N_22114,N_20053,N_20227);
nand U22115 (N_22115,N_21021,N_20596);
or U22116 (N_22116,N_20542,N_20986);
and U22117 (N_22117,N_20492,N_21042);
or U22118 (N_22118,N_21309,N_21909);
nor U22119 (N_22119,N_20191,N_21381);
xor U22120 (N_22120,N_20295,N_21093);
xnor U22121 (N_22121,N_20477,N_20052);
xnor U22122 (N_22122,N_21508,N_21603);
and U22123 (N_22123,N_21800,N_20351);
nand U22124 (N_22124,N_21804,N_20183);
nand U22125 (N_22125,N_20068,N_20341);
or U22126 (N_22126,N_21534,N_21974);
and U22127 (N_22127,N_20199,N_20148);
xnor U22128 (N_22128,N_21697,N_21814);
nor U22129 (N_22129,N_21091,N_20943);
nor U22130 (N_22130,N_21870,N_20412);
and U22131 (N_22131,N_20724,N_21579);
and U22132 (N_22132,N_20153,N_21533);
and U22133 (N_22133,N_21148,N_21119);
xor U22134 (N_22134,N_20796,N_21540);
or U22135 (N_22135,N_20896,N_20122);
and U22136 (N_22136,N_20135,N_20220);
xnor U22137 (N_22137,N_20027,N_20647);
nand U22138 (N_22138,N_21944,N_20078);
nor U22139 (N_22139,N_21694,N_21189);
and U22140 (N_22140,N_21360,N_21097);
or U22141 (N_22141,N_21498,N_20185);
nor U22142 (N_22142,N_21173,N_20380);
xnor U22143 (N_22143,N_20124,N_21501);
xor U22144 (N_22144,N_20944,N_21884);
or U22145 (N_22145,N_20743,N_21695);
or U22146 (N_22146,N_21840,N_21516);
and U22147 (N_22147,N_20243,N_20712);
nor U22148 (N_22148,N_21852,N_20406);
nand U22149 (N_22149,N_20993,N_21257);
xnor U22150 (N_22150,N_21999,N_20163);
and U22151 (N_22151,N_21448,N_21256);
nand U22152 (N_22152,N_21428,N_20302);
xnor U22153 (N_22153,N_21180,N_21102);
or U22154 (N_22154,N_21241,N_21795);
xnor U22155 (N_22155,N_20573,N_20602);
nor U22156 (N_22156,N_20239,N_20293);
nand U22157 (N_22157,N_21047,N_21248);
and U22158 (N_22158,N_20485,N_20959);
and U22159 (N_22159,N_21115,N_20008);
nand U22160 (N_22160,N_21777,N_20910);
nor U22161 (N_22161,N_20256,N_21132);
nand U22162 (N_22162,N_21237,N_20024);
nor U22163 (N_22163,N_20493,N_20118);
xnor U22164 (N_22164,N_21046,N_20608);
xnor U22165 (N_22165,N_20671,N_21403);
xor U22166 (N_22166,N_21429,N_20244);
nor U22167 (N_22167,N_20016,N_21539);
nor U22168 (N_22168,N_20452,N_20662);
nand U22169 (N_22169,N_21720,N_20687);
nand U22170 (N_22170,N_20852,N_21615);
nor U22171 (N_22171,N_20367,N_21580);
xor U22172 (N_22172,N_20441,N_20640);
or U22173 (N_22173,N_20446,N_21701);
nor U22174 (N_22174,N_21484,N_21099);
nor U22175 (N_22175,N_20981,N_20399);
nor U22176 (N_22176,N_21254,N_20557);
nand U22177 (N_22177,N_20329,N_21196);
and U22178 (N_22178,N_21960,N_20804);
nand U22179 (N_22179,N_21161,N_21440);
nor U22180 (N_22180,N_21952,N_21535);
xor U22181 (N_22181,N_21301,N_20349);
nand U22182 (N_22182,N_20416,N_20739);
and U22183 (N_22183,N_21375,N_21039);
xor U22184 (N_22184,N_21101,N_20877);
xnor U22185 (N_22185,N_20069,N_21321);
nor U22186 (N_22186,N_20437,N_21946);
and U22187 (N_22187,N_21013,N_21392);
xnor U22188 (N_22188,N_20825,N_21339);
nor U22189 (N_22189,N_21947,N_20560);
or U22190 (N_22190,N_20326,N_20960);
or U22191 (N_22191,N_20591,N_20681);
or U22192 (N_22192,N_21288,N_21350);
nand U22193 (N_22193,N_20606,N_21022);
or U22194 (N_22194,N_20942,N_21730);
xnor U22195 (N_22195,N_21293,N_21144);
nand U22196 (N_22196,N_21616,N_21192);
or U22197 (N_22197,N_20042,N_20426);
nor U22198 (N_22198,N_20663,N_20801);
xnor U22199 (N_22199,N_20758,N_20179);
and U22200 (N_22200,N_20823,N_20624);
nand U22201 (N_22201,N_21712,N_20985);
and U22202 (N_22202,N_21891,N_20652);
nand U22203 (N_22203,N_21541,N_20980);
xnor U22204 (N_22204,N_20945,N_21128);
nand U22205 (N_22205,N_21333,N_20298);
nor U22206 (N_22206,N_21993,N_20092);
nand U22207 (N_22207,N_20616,N_20203);
and U22208 (N_22208,N_20716,N_21546);
or U22209 (N_22209,N_20525,N_21917);
and U22210 (N_22210,N_20574,N_20818);
or U22211 (N_22211,N_21290,N_20144);
nor U22212 (N_22212,N_21434,N_21316);
or U22213 (N_22213,N_21338,N_20674);
nor U22214 (N_22214,N_21950,N_21666);
nand U22215 (N_22215,N_21980,N_21570);
or U22216 (N_22216,N_20178,N_21780);
nand U22217 (N_22217,N_21715,N_21831);
or U22218 (N_22218,N_21766,N_21142);
or U22219 (N_22219,N_20831,N_20996);
or U22220 (N_22220,N_20814,N_21679);
nand U22221 (N_22221,N_21286,N_20056);
nor U22222 (N_22222,N_21503,N_20390);
nor U22223 (N_22223,N_21589,N_21030);
xor U22224 (N_22224,N_20731,N_21585);
nand U22225 (N_22225,N_20693,N_20360);
xnor U22226 (N_22226,N_21383,N_21170);
xnor U22227 (N_22227,N_21104,N_20270);
nand U22228 (N_22228,N_21978,N_20563);
xnor U22229 (N_22229,N_20212,N_21549);
xor U22230 (N_22230,N_20269,N_21373);
xor U22231 (N_22231,N_21010,N_21349);
or U22232 (N_22232,N_20665,N_21558);
xor U22233 (N_22233,N_20523,N_20311);
nand U22234 (N_22234,N_21716,N_20723);
nand U22235 (N_22235,N_21738,N_20342);
or U22236 (N_22236,N_21583,N_20489);
or U22237 (N_22237,N_21439,N_20421);
nand U22238 (N_22238,N_20372,N_21108);
nor U22239 (N_22239,N_21745,N_20888);
nand U22240 (N_22240,N_20235,N_20274);
nor U22241 (N_22241,N_20838,N_20700);
nor U22242 (N_22242,N_21274,N_20843);
xnor U22243 (N_22243,N_20376,N_21236);
and U22244 (N_22244,N_20014,N_21149);
nand U22245 (N_22245,N_21255,N_21851);
nor U22246 (N_22246,N_20356,N_21502);
and U22247 (N_22247,N_21991,N_21606);
nand U22248 (N_22248,N_20196,N_20461);
xnor U22249 (N_22249,N_21920,N_20549);
nand U22250 (N_22250,N_20976,N_21480);
and U22251 (N_22251,N_21929,N_21382);
nand U22252 (N_22252,N_21823,N_20783);
or U22253 (N_22253,N_20740,N_21684);
xor U22254 (N_22254,N_21222,N_21076);
and U22255 (N_22255,N_21345,N_21068);
nor U22256 (N_22256,N_21963,N_20066);
or U22257 (N_22257,N_21045,N_20728);
xor U22258 (N_22258,N_20292,N_20023);
nor U22259 (N_22259,N_21675,N_21836);
and U22260 (N_22260,N_20459,N_20676);
xor U22261 (N_22261,N_21997,N_20881);
nand U22262 (N_22262,N_20961,N_21908);
nand U22263 (N_22263,N_20701,N_21479);
nand U22264 (N_22264,N_20669,N_20319);
xor U22265 (N_22265,N_20222,N_20899);
nor U22266 (N_22266,N_21753,N_21476);
nor U22267 (N_22267,N_20759,N_21230);
nand U22268 (N_22268,N_20868,N_20273);
xor U22269 (N_22269,N_20009,N_21658);
nor U22270 (N_22270,N_21857,N_20581);
nor U22271 (N_22271,N_20345,N_20171);
nand U22272 (N_22272,N_20405,N_21925);
xnor U22273 (N_22273,N_20684,N_21049);
and U22274 (N_22274,N_21326,N_20388);
xor U22275 (N_22275,N_20140,N_20382);
or U22276 (N_22276,N_21156,N_21750);
nor U22277 (N_22277,N_21597,N_21739);
xor U22278 (N_22278,N_21399,N_21521);
and U22279 (N_22279,N_20327,N_21166);
nand U22280 (N_22280,N_20201,N_20705);
nand U22281 (N_22281,N_20245,N_21444);
nand U22282 (N_22282,N_20966,N_20738);
xnor U22283 (N_22283,N_20396,N_21138);
or U22284 (N_22284,N_21233,N_20147);
or U22285 (N_22285,N_21906,N_21298);
xnor U22286 (N_22286,N_21229,N_21312);
nand U22287 (N_22287,N_21690,N_20497);
and U22288 (N_22288,N_20003,N_20821);
or U22289 (N_22289,N_21017,N_21234);
and U22290 (N_22290,N_21320,N_21463);
nand U22291 (N_22291,N_21735,N_21569);
and U22292 (N_22292,N_20514,N_21855);
or U22293 (N_22293,N_20328,N_20619);
nand U22294 (N_22294,N_21355,N_20395);
or U22295 (N_22295,N_21873,N_20924);
nor U22296 (N_22296,N_20043,N_20850);
and U22297 (N_22297,N_20490,N_21904);
nand U22298 (N_22298,N_21024,N_21201);
xnor U22299 (N_22299,N_21131,N_21133);
nand U22300 (N_22300,N_20696,N_20126);
xor U22301 (N_22301,N_20190,N_20706);
xor U22302 (N_22302,N_21670,N_20173);
xor U22303 (N_22303,N_20186,N_21127);
nor U22304 (N_22304,N_20371,N_20305);
nand U22305 (N_22305,N_21211,N_20779);
or U22306 (N_22306,N_21393,N_20134);
nand U22307 (N_22307,N_21958,N_21740);
or U22308 (N_22308,N_20407,N_21143);
xor U22309 (N_22309,N_20879,N_21964);
nor U22310 (N_22310,N_20154,N_21388);
xor U22311 (N_22311,N_20278,N_20076);
nand U22312 (N_22312,N_21763,N_20928);
nand U22313 (N_22313,N_20275,N_20346);
nand U22314 (N_22314,N_20660,N_21424);
nand U22315 (N_22315,N_21949,N_21450);
nor U22316 (N_22316,N_20774,N_21644);
nor U22317 (N_22317,N_21518,N_21566);
xor U22318 (N_22318,N_21308,N_20240);
nor U22319 (N_22319,N_21206,N_20473);
xor U22320 (N_22320,N_21325,N_20468);
nand U22321 (N_22321,N_20953,N_21249);
xnor U22322 (N_22322,N_21147,N_20104);
and U22323 (N_22323,N_21486,N_21086);
and U22324 (N_22324,N_20379,N_20160);
and U22325 (N_22325,N_20839,N_21460);
and U22326 (N_22326,N_21074,N_21151);
nand U22327 (N_22327,N_20718,N_21862);
xor U22328 (N_22328,N_21698,N_20431);
nor U22329 (N_22329,N_21402,N_20075);
nor U22330 (N_22330,N_21749,N_21988);
nor U22331 (N_22331,N_21837,N_20350);
nor U22332 (N_22332,N_21523,N_21344);
or U22333 (N_22333,N_21187,N_21871);
nor U22334 (N_22334,N_20262,N_21930);
and U22335 (N_22335,N_21921,N_21331);
and U22336 (N_22336,N_20933,N_21667);
or U22337 (N_22337,N_21250,N_20418);
nand U22338 (N_22338,N_20257,N_20339);
and U22339 (N_22339,N_20802,N_21512);
nor U22340 (N_22340,N_21171,N_20300);
xnor U22341 (N_22341,N_21397,N_20479);
xnor U22342 (N_22342,N_21544,N_21477);
xnor U22343 (N_22343,N_20642,N_21487);
and U22344 (N_22344,N_20517,N_21688);
or U22345 (N_22345,N_21496,N_20001);
nand U22346 (N_22346,N_21861,N_21263);
and U22347 (N_22347,N_20120,N_21227);
and U22348 (N_22348,N_20562,N_21754);
nand U22349 (N_22349,N_21696,N_21500);
xor U22350 (N_22350,N_20580,N_21591);
nand U22351 (N_22351,N_21961,N_21404);
xor U22352 (N_22352,N_20564,N_21833);
and U22353 (N_22353,N_20994,N_20434);
and U22354 (N_22354,N_20130,N_20595);
or U22355 (N_22355,N_20429,N_21182);
xor U22356 (N_22356,N_20475,N_21577);
nor U22357 (N_22357,N_21281,N_20629);
or U22358 (N_22358,N_21185,N_20002);
nand U22359 (N_22359,N_21646,N_21297);
nand U22360 (N_22360,N_20934,N_20841);
or U22361 (N_22361,N_21183,N_21370);
nand U22362 (N_22362,N_20150,N_20781);
nand U22363 (N_22363,N_21945,N_20890);
and U22364 (N_22364,N_21866,N_20484);
nor U22365 (N_22365,N_20699,N_20764);
nand U22366 (N_22366,N_20471,N_20138);
and U22367 (N_22367,N_21336,N_20025);
or U22368 (N_22368,N_20834,N_21802);
xor U22369 (N_22369,N_20030,N_21202);
or U22370 (N_22370,N_20455,N_20251);
xnor U22371 (N_22371,N_20997,N_21736);
nor U22372 (N_22372,N_21292,N_20209);
nand U22373 (N_22373,N_20604,N_21604);
or U22374 (N_22374,N_21072,N_20366);
xnor U22375 (N_22375,N_20091,N_20206);
and U22376 (N_22376,N_20093,N_20088);
xnor U22377 (N_22377,N_20636,N_20260);
xnor U22378 (N_22378,N_21311,N_21758);
nor U22379 (N_22379,N_21655,N_20451);
xor U22380 (N_22380,N_20233,N_21362);
and U22381 (N_22381,N_21761,N_21054);
and U22382 (N_22382,N_21733,N_21340);
nand U22383 (N_22383,N_21922,N_20058);
xnor U22384 (N_22384,N_21083,N_20713);
nor U22385 (N_22385,N_20538,N_20208);
xor U22386 (N_22386,N_20678,N_20704);
or U22387 (N_22387,N_20112,N_21445);
nor U22388 (N_22388,N_21441,N_20726);
nand U22389 (N_22389,N_21959,N_21955);
nand U22390 (N_22390,N_20355,N_20231);
nor U22391 (N_22391,N_21458,N_20184);
nor U22392 (N_22392,N_20588,N_20383);
or U22393 (N_22393,N_21430,N_21279);
xor U22394 (N_22394,N_21343,N_20972);
nor U22395 (N_22395,N_21391,N_20105);
xnor U22396 (N_22396,N_21358,N_21238);
or U22397 (N_22397,N_20012,N_20285);
and U22398 (N_22398,N_20544,N_20252);
and U22399 (N_22399,N_20116,N_21617);
and U22400 (N_22400,N_21938,N_21177);
xor U22401 (N_22401,N_20569,N_20844);
and U22402 (N_22402,N_21576,N_20623);
and U22403 (N_22403,N_20392,N_20855);
nor U22404 (N_22404,N_20710,N_20427);
nand U22405 (N_22405,N_20498,N_21285);
nand U22406 (N_22406,N_21079,N_20742);
nand U22407 (N_22407,N_21654,N_21040);
and U22408 (N_22408,N_20664,N_21240);
nand U22409 (N_22409,N_20987,N_20129);
xnor U22410 (N_22410,N_21619,N_21036);
or U22411 (N_22411,N_20922,N_21630);
nor U22412 (N_22412,N_21582,N_20268);
nand U22413 (N_22413,N_20603,N_21648);
nor U22414 (N_22414,N_21251,N_20157);
and U22415 (N_22415,N_20982,N_20145);
or U22416 (N_22416,N_20555,N_21966);
nand U22417 (N_22417,N_20938,N_21481);
and U22418 (N_22418,N_21798,N_20100);
or U22419 (N_22419,N_21788,N_21681);
or U22420 (N_22420,N_20237,N_21218);
xor U22421 (N_22421,N_20151,N_21965);
xor U22422 (N_22422,N_20170,N_21522);
or U22423 (N_22423,N_21412,N_21379);
or U22424 (N_22424,N_20331,N_20526);
nand U22425 (N_22425,N_20404,N_20826);
xnor U22426 (N_22426,N_21284,N_20658);
and U22427 (N_22427,N_20502,N_21858);
nand U22428 (N_22428,N_20780,N_21751);
and U22429 (N_22429,N_20417,N_21359);
nand U22430 (N_22430,N_21095,N_20359);
nand U22431 (N_22431,N_20086,N_21310);
or U22432 (N_22432,N_21158,N_21106);
or U22433 (N_22433,N_20749,N_21979);
nand U22434 (N_22434,N_20703,N_20625);
nor U22435 (N_22435,N_20026,N_20230);
and U22436 (N_22436,N_21346,N_21726);
or U22437 (N_22437,N_20509,N_20661);
xnor U22438 (N_22438,N_20414,N_20884);
and U22439 (N_22439,N_21414,N_21426);
nand U22440 (N_22440,N_21411,N_20931);
nor U22441 (N_22441,N_20108,N_20644);
nor U22442 (N_22442,N_20921,N_20751);
and U22443 (N_22443,N_20004,N_21806);
xor U22444 (N_22444,N_20337,N_21942);
nor U22445 (N_22445,N_20187,N_20478);
xor U22446 (N_22446,N_21613,N_21692);
xor U22447 (N_22447,N_21226,N_21609);
nand U22448 (N_22448,N_21216,N_20254);
nand U22449 (N_22449,N_20435,N_20534);
and U22450 (N_22450,N_20065,N_21179);
xor U22451 (N_22451,N_21557,N_21014);
and U22452 (N_22452,N_21469,N_20089);
xor U22453 (N_22453,N_21731,N_21398);
and U22454 (N_22454,N_21706,N_21258);
xnor U22455 (N_22455,N_21299,N_20762);
and U22456 (N_22456,N_20015,N_20152);
nor U22457 (N_22457,N_21260,N_21796);
xor U22458 (N_22458,N_21623,N_21005);
and U22459 (N_22459,N_21728,N_20384);
nor U22460 (N_22460,N_21936,N_20677);
xor U22461 (N_22461,N_21742,N_21832);
nor U22462 (N_22462,N_21640,N_20467);
nand U22463 (N_22463,N_21636,N_21771);
xor U22464 (N_22464,N_21289,N_20503);
or U22465 (N_22465,N_20746,N_20572);
nand U22466 (N_22466,N_21317,N_21772);
xnor U22467 (N_22467,N_21626,N_21817);
nor U22468 (N_22468,N_21052,N_20221);
or U22469 (N_22469,N_20167,N_21809);
and U22470 (N_22470,N_21437,N_20299);
or U22471 (N_22471,N_21056,N_20210);
and U22472 (N_22472,N_21683,N_20568);
nor U22473 (N_22473,N_20165,N_20977);
nand U22474 (N_22474,N_20627,N_21483);
or U22475 (N_22475,N_20159,N_21531);
xor U22476 (N_22476,N_21680,N_20486);
and U22477 (N_22477,N_21446,N_20592);
and U22478 (N_22478,N_20436,N_21867);
and U22479 (N_22479,N_21888,N_20071);
xor U22480 (N_22480,N_20812,N_21970);
and U22481 (N_22481,N_21075,N_21900);
or U22482 (N_22482,N_20935,N_21801);
and U22483 (N_22483,N_20031,N_20320);
nand U22484 (N_22484,N_21807,N_20628);
and U22485 (N_22485,N_20306,N_20400);
nor U22486 (N_22486,N_20853,N_20858);
or U22487 (N_22487,N_20730,N_20368);
xor U22488 (N_22488,N_21525,N_21794);
nand U22489 (N_22489,N_21889,N_21874);
and U22490 (N_22490,N_21563,N_21578);
and U22491 (N_22491,N_21208,N_20833);
or U22492 (N_22492,N_21524,N_20304);
and U22493 (N_22493,N_21586,N_20794);
nor U22494 (N_22494,N_21327,N_21080);
or U22495 (N_22495,N_21792,N_21057);
and U22496 (N_22496,N_21342,N_21427);
nand U22497 (N_22497,N_20035,N_20028);
nor U22498 (N_22498,N_21975,N_21934);
and U22499 (N_22499,N_21094,N_20466);
xnor U22500 (N_22500,N_20491,N_21475);
xor U22501 (N_22501,N_20842,N_21070);
nand U22502 (N_22502,N_20470,N_20137);
or U22503 (N_22503,N_21628,N_21528);
nor U22504 (N_22504,N_20049,N_21651);
xnor U22505 (N_22505,N_20864,N_20756);
nor U22506 (N_22506,N_21457,N_20271);
xnor U22507 (N_22507,N_21396,N_21197);
nand U22508 (N_22508,N_21176,N_20668);
xor U22509 (N_22509,N_21747,N_20114);
nand U22510 (N_22510,N_21620,N_21117);
xor U22511 (N_22511,N_20576,N_21553);
or U22512 (N_22512,N_21065,N_21488);
nor U22513 (N_22513,N_20387,N_21456);
nor U22514 (N_22514,N_21555,N_20018);
and U22515 (N_22515,N_21860,N_21668);
xor U22516 (N_22516,N_20386,N_20732);
and U22517 (N_22517,N_20101,N_20448);
and U22518 (N_22518,N_21341,N_20287);
nand U22519 (N_22519,N_20975,N_20223);
and U22520 (N_22520,N_21677,N_21507);
and U22521 (N_22521,N_21195,N_20760);
and U22522 (N_22522,N_20867,N_20672);
or U22523 (N_22523,N_20641,N_20791);
and U22524 (N_22524,N_20343,N_20115);
nand U22525 (N_22525,N_21053,N_20917);
nand U22526 (N_22526,N_21574,N_21592);
nand U22527 (N_22527,N_20106,N_20815);
nor U22528 (N_22528,N_21116,N_20411);
nor U22529 (N_22529,N_20317,N_21983);
nor U22530 (N_22530,N_20198,N_21154);
nor U22531 (N_22531,N_21595,N_21305);
nor U22532 (N_22532,N_21495,N_21568);
xor U22533 (N_22533,N_20819,N_21693);
and U22534 (N_22534,N_20529,N_21366);
nor U22535 (N_22535,N_20715,N_20600);
nand U22536 (N_22536,N_21868,N_21971);
nand U22537 (N_22537,N_21313,N_21998);
and U22538 (N_22538,N_21678,N_20226);
nor U22539 (N_22539,N_20800,N_20599);
xnor U22540 (N_22540,N_20340,N_20321);
or U22541 (N_22541,N_20717,N_21687);
and U22542 (N_22542,N_20481,N_21050);
nand U22543 (N_22543,N_21911,N_20537);
nor U22544 (N_22544,N_21423,N_20377);
and U22545 (N_22545,N_20121,N_20401);
nand U22546 (N_22546,N_20655,N_21665);
or U22547 (N_22547,N_21624,N_21785);
or U22548 (N_22548,N_20719,N_20074);
or U22549 (N_22549,N_20419,N_20207);
nor U22550 (N_22550,N_21590,N_20458);
or U22551 (N_22551,N_21509,N_21702);
xor U22552 (N_22552,N_20241,N_21663);
nor U22553 (N_22553,N_20929,N_20561);
or U22554 (N_22554,N_21886,N_21210);
and U22555 (N_22555,N_21207,N_20482);
xnor U22556 (N_22556,N_20589,N_21926);
nor U22557 (N_22557,N_20720,N_21322);
or U22558 (N_22558,N_20238,N_21084);
nor U22559 (N_22559,N_21764,N_20680);
nand U22560 (N_22560,N_21813,N_21672);
or U22561 (N_22561,N_20631,N_21572);
xor U22562 (N_22562,N_21618,N_21253);
and U22563 (N_22563,N_21394,N_21432);
or U22564 (N_22564,N_21387,N_20005);
and U22565 (N_22565,N_21768,N_20019);
nand U22566 (N_22566,N_20309,N_21016);
xnor U22567 (N_22567,N_21368,N_21006);
nand U22568 (N_22568,N_20956,N_20754);
and U22569 (N_22569,N_21385,N_21567);
nand U22570 (N_22570,N_20989,N_20062);
xnor U22571 (N_22571,N_21536,N_20795);
or U22572 (N_22572,N_20736,N_20859);
nor U22573 (N_22573,N_20483,N_20897);
xnor U22574 (N_22574,N_20984,N_20784);
nand U22575 (N_22575,N_21357,N_21976);
xor U22576 (N_22576,N_20613,N_21811);
or U22577 (N_22577,N_20916,N_21198);
nor U22578 (N_22578,N_20957,N_20265);
or U22579 (N_22579,N_20070,N_21854);
nand U22580 (N_22580,N_21474,N_21822);
nand U22581 (N_22581,N_21773,N_21704);
and U22582 (N_22582,N_21002,N_21571);
nand U22583 (N_22583,N_20524,N_21573);
xnor U22584 (N_22584,N_20992,N_20889);
nor U22585 (N_22585,N_21602,N_21493);
xor U22586 (N_22586,N_20782,N_20725);
and U22587 (N_22587,N_20381,N_20808);
xor U22588 (N_22588,N_20480,N_20099);
xnor U22589 (N_22589,N_21638,N_21652);
xnor U22590 (N_22590,N_21869,N_21614);
nand U22591 (N_22591,N_20870,N_21037);
or U22592 (N_22592,N_20143,N_20775);
or U22593 (N_22593,N_20348,N_21032);
or U22594 (N_22594,N_20667,N_20194);
or U22595 (N_22595,N_20551,N_20084);
nor U22596 (N_22596,N_20255,N_21550);
nand U22597 (N_22597,N_20772,N_20894);
nor U22598 (N_22598,N_21984,N_21532);
nor U22599 (N_22599,N_20303,N_20585);
nand U22600 (N_22600,N_20874,N_21721);
or U22601 (N_22601,N_20176,N_21554);
xnor U22602 (N_22602,N_21835,N_20177);
or U22603 (N_22603,N_20296,N_20694);
nand U22604 (N_22604,N_21087,N_20689);
and U22605 (N_22605,N_20605,N_21136);
and U22606 (N_22606,N_20528,N_20047);
and U22607 (N_22607,N_21718,N_21600);
or U22608 (N_22608,N_21491,N_21364);
nor U22609 (N_22609,N_21135,N_20188);
nor U22610 (N_22610,N_21892,N_20995);
xor U22611 (N_22611,N_21821,N_20805);
nor U22612 (N_22612,N_21442,N_20548);
or U22613 (N_22613,N_21676,N_20045);
nand U22614 (N_22614,N_21895,N_20639);
xnor U22615 (N_22615,N_20063,N_21239);
xnor U22616 (N_22616,N_20744,N_20919);
nor U22617 (N_22617,N_20500,N_21903);
or U22618 (N_22618,N_21556,N_21181);
and U22619 (N_22619,N_20651,N_20893);
nand U22620 (N_22620,N_21447,N_21029);
xor U22621 (N_22621,N_20952,N_21330);
xor U22622 (N_22622,N_21838,N_20809);
or U22623 (N_22623,N_21789,N_21186);
xor U22624 (N_22624,N_21221,N_20522);
nor U22625 (N_22625,N_21657,N_21011);
xnor U22626 (N_22626,N_21103,N_21653);
nand U22627 (N_22627,N_21482,N_21842);
xor U22628 (N_22628,N_20279,N_21214);
nor U22629 (N_22629,N_20745,N_20432);
xor U22630 (N_22630,N_21765,N_21547);
and U22631 (N_22631,N_20830,N_20051);
or U22632 (N_22632,N_21756,N_20683);
nor U22633 (N_22633,N_21283,N_20288);
nand U22634 (N_22634,N_20236,N_21781);
xor U22635 (N_22635,N_20583,N_21259);
nor U22636 (N_22636,N_20873,N_21878);
or U22637 (N_22637,N_21377,N_20875);
xor U22638 (N_22638,N_20902,N_20582);
or U22639 (N_22639,N_21709,N_21551);
nand U22640 (N_22640,N_21118,N_20193);
nand U22641 (N_22641,N_21361,N_20622);
and U22642 (N_22642,N_20828,N_21601);
xnor U22643 (N_22643,N_20939,N_20033);
nor U22644 (N_22644,N_20964,N_20266);
nor U22645 (N_22645,N_20558,N_20456);
and U22646 (N_22646,N_20217,N_21380);
or U22647 (N_22647,N_21141,N_21916);
nor U22648 (N_22648,N_21844,N_21641);
and U22649 (N_22649,N_21912,N_20333);
nor U22650 (N_22650,N_21467,N_21770);
or U22651 (N_22651,N_21846,N_21264);
and U22652 (N_22652,N_20307,N_21918);
nor U22653 (N_22653,N_20516,N_21242);
nor U22654 (N_22654,N_20648,N_20883);
xnor U22655 (N_22655,N_20204,N_21438);
nand U22656 (N_22656,N_21839,N_20409);
xor U22657 (N_22657,N_20232,N_20567);
and U22658 (N_22658,N_21337,N_20156);
nand U22659 (N_22659,N_21856,N_21098);
nor U22660 (N_22660,N_21875,N_20282);
nand U22661 (N_22661,N_20155,N_21732);
nor U22662 (N_22662,N_21073,N_20469);
nor U22663 (N_22663,N_20166,N_20798);
xnor U22664 (N_22664,N_20849,N_20611);
nand U22665 (N_22665,N_20374,N_20218);
and U22666 (N_22666,N_21407,N_21713);
nand U22667 (N_22667,N_21419,N_20082);
and U22668 (N_22668,N_21167,N_20508);
xor U22669 (N_22669,N_20445,N_20403);
xnor U22670 (N_22670,N_20192,N_20722);
or U22671 (N_22671,N_20213,N_21816);
and U22672 (N_22672,N_21853,N_21061);
or U22673 (N_22673,N_20442,N_20164);
xor U22674 (N_22674,N_21270,N_21596);
or U22675 (N_22675,N_21621,N_21278);
and U22676 (N_22676,N_20353,N_21793);
or U22677 (N_22677,N_20136,N_20913);
and U22678 (N_22678,N_21561,N_20630);
xor U22679 (N_22679,N_21000,N_20261);
nor U22680 (N_22680,N_21435,N_21244);
nand U22681 (N_22681,N_21431,N_20793);
and U22682 (N_22682,N_20653,N_20457);
and U22683 (N_22683,N_21631,N_21082);
nand U22684 (N_22684,N_21306,N_21220);
nand U22685 (N_22685,N_20635,N_20901);
nand U22686 (N_22686,N_21612,N_21209);
nor U22687 (N_22687,N_21164,N_20840);
or U22688 (N_22688,N_21295,N_20378);
and U22689 (N_22689,N_21826,N_21165);
nand U22690 (N_22690,N_21422,N_20229);
xnor U22691 (N_22691,N_20638,N_20545);
nand U22692 (N_22692,N_21905,N_20954);
nor U22693 (N_22693,N_21829,N_21635);
nand U22694 (N_22694,N_21433,N_20520);
nor U22695 (N_22695,N_21224,N_21787);
xnor U22696 (N_22696,N_21593,N_21849);
nor U22697 (N_22697,N_20413,N_20499);
nor U22698 (N_22698,N_20181,N_20951);
or U22699 (N_22699,N_21465,N_21268);
nand U22700 (N_22700,N_20752,N_20750);
nor U22701 (N_22701,N_20128,N_20836);
and U22702 (N_22702,N_20038,N_20290);
and U22703 (N_22703,N_21703,N_20865);
or U22704 (N_22704,N_21957,N_20654);
nand U22705 (N_22705,N_21935,N_20385);
or U22706 (N_22706,N_21200,N_21269);
and U22707 (N_22707,N_20496,N_20778);
xnor U22708 (N_22708,N_20707,N_21707);
or U22709 (N_22709,N_21033,N_21996);
nand U22710 (N_22710,N_20552,N_20926);
or U22711 (N_22711,N_21594,N_20352);
or U22712 (N_22712,N_20361,N_21449);
and U22713 (N_22713,N_21245,N_20941);
nand U22714 (N_22714,N_21243,N_20272);
nor U22715 (N_22715,N_21365,N_20363);
or U22716 (N_22716,N_20318,N_21634);
nor U22717 (N_22717,N_20022,N_21643);
nor U22718 (N_22718,N_20488,N_20990);
and U22719 (N_22719,N_21485,N_21468);
nor U22720 (N_22720,N_20866,N_20851);
and U22721 (N_22721,N_20963,N_21009);
or U22722 (N_22722,N_20962,N_21662);
nor U22723 (N_22723,N_20590,N_20685);
nand U22724 (N_22724,N_21962,N_21043);
nor U22725 (N_22725,N_21287,N_20790);
nand U22726 (N_22726,N_20579,N_21277);
or U22727 (N_22727,N_20057,N_21865);
and U22728 (N_22728,N_21303,N_20918);
xor U22729 (N_22729,N_21729,N_21111);
nor U22730 (N_22730,N_21231,N_21275);
xor U22731 (N_22731,N_20721,N_21815);
and U22732 (N_22732,N_21389,N_20553);
nor U22733 (N_22733,N_20085,N_21881);
or U22734 (N_22734,N_21417,N_20766);
or U22735 (N_22735,N_21090,N_20632);
xnor U22736 (N_22736,N_20978,N_21880);
nand U22737 (N_22737,N_21977,N_20430);
and U22738 (N_22738,N_20146,N_20375);
nand U22739 (N_22739,N_21193,N_20643);
and U22740 (N_22740,N_20697,N_21363);
nor U22741 (N_22741,N_20109,N_21409);
nand U22742 (N_22742,N_20362,N_21737);
and U22743 (N_22743,N_21882,N_20747);
xor U22744 (N_22744,N_20291,N_20657);
nand U22745 (N_22745,N_20770,N_21538);
or U22746 (N_22746,N_21744,N_21622);
and U22747 (N_22747,N_21919,N_21125);
and U22748 (N_22748,N_20449,N_20908);
nor U22749 (N_22749,N_20675,N_20511);
nand U22750 (N_22750,N_20659,N_20495);
nand U22751 (N_22751,N_20903,N_21232);
xor U22752 (N_22752,N_21415,N_20690);
nor U22753 (N_22753,N_20811,N_20540);
xor U22754 (N_22754,N_20253,N_20397);
and U22755 (N_22755,N_20077,N_20991);
and U22756 (N_22756,N_21092,N_21691);
xor U22757 (N_22757,N_21985,N_21647);
or U22758 (N_22758,N_20927,N_21205);
xnor U22759 (N_22759,N_21588,N_20789);
or U22760 (N_22760,N_20797,N_21723);
or U22761 (N_22761,N_20950,N_21543);
and U22762 (N_22762,N_20476,N_20829);
or U22763 (N_22763,N_20402,N_20175);
xnor U22764 (N_22764,N_20338,N_20565);
xor U22765 (N_22765,N_21954,N_20205);
and U22766 (N_22766,N_20891,N_20006);
and U22767 (N_22767,N_21982,N_21089);
xnor U22768 (N_22768,N_20472,N_20310);
nor U22769 (N_22769,N_20810,N_20010);
and U22770 (N_22770,N_20440,N_21940);
or U22771 (N_22771,N_20172,N_21058);
and U22772 (N_22772,N_20656,N_20837);
or U22773 (N_22773,N_20692,N_21741);
xor U22774 (N_22774,N_20267,N_21968);
and U22775 (N_22775,N_21762,N_21109);
nand U22776 (N_22776,N_21453,N_21700);
and U22777 (N_22777,N_20900,N_21421);
nor U22778 (N_22778,N_20314,N_21526);
or U22779 (N_22779,N_21608,N_21499);
and U22780 (N_22780,N_20727,N_20771);
or U22781 (N_22781,N_21335,N_21914);
nand U22782 (N_22782,N_21808,N_20487);
xnor U22783 (N_22783,N_20673,N_21410);
nor U22784 (N_22784,N_21629,N_21012);
and U22785 (N_22785,N_20741,N_21828);
xnor U22786 (N_22786,N_20315,N_21066);
and U22787 (N_22787,N_21462,N_21121);
or U22788 (N_22788,N_21972,N_21902);
nor U22789 (N_22789,N_21126,N_20912);
nand U22790 (N_22790,N_20566,N_20098);
nand U22791 (N_22791,N_20614,N_20617);
nand U22792 (N_22792,N_20559,N_21055);
nand U22793 (N_22793,N_21472,N_21352);
or U22794 (N_22794,N_21078,N_20474);
xor U22795 (N_22795,N_20649,N_20586);
nand U22796 (N_22796,N_21927,N_21513);
and U22797 (N_22797,N_21708,N_20776);
or U22798 (N_22798,N_21530,N_20393);
or U22799 (N_22799,N_21937,N_20264);
nand U22800 (N_22800,N_21163,N_20876);
nand U22801 (N_22801,N_20059,N_20734);
xnor U22802 (N_22802,N_21372,N_21261);
nor U22803 (N_22803,N_21711,N_20556);
nand U22804 (N_22804,N_21157,N_21673);
nor U22805 (N_22805,N_21783,N_21035);
nor U22806 (N_22806,N_21008,N_21633);
or U22807 (N_22807,N_21986,N_20061);
and U22808 (N_22808,N_21992,N_20369);
nand U22809 (N_22809,N_21724,N_21062);
xnor U22810 (N_22810,N_21025,N_20803);
xor U22811 (N_22811,N_21347,N_21296);
or U22812 (N_22812,N_21139,N_21146);
nand U22813 (N_22813,N_20465,N_20974);
nand U22814 (N_22814,N_20645,N_21995);
or U22815 (N_22815,N_20763,N_21899);
and U22816 (N_22816,N_21262,N_20197);
nor U22817 (N_22817,N_20691,N_20958);
or U22818 (N_22818,N_20587,N_21824);
nand U22819 (N_22819,N_20948,N_21319);
xor U22820 (N_22820,N_21812,N_20915);
nor U22821 (N_22821,N_20753,N_20162);
nor U22822 (N_22822,N_21847,N_20513);
and U22823 (N_22823,N_21928,N_21228);
or U22824 (N_22824,N_21510,N_21611);
nor U22825 (N_22825,N_20787,N_21152);
nand U22826 (N_22826,N_21803,N_21153);
xnor U22827 (N_22827,N_20087,N_20550);
nand U22828 (N_22828,N_21948,N_20141);
xnor U22829 (N_22829,N_21120,N_21907);
and U22830 (N_22830,N_20755,N_20242);
nor U22831 (N_22831,N_21776,N_20336);
or U22832 (N_22832,N_20073,N_21471);
nor U22833 (N_22833,N_21026,N_21506);
nand U22834 (N_22834,N_21019,N_21390);
nand U22835 (N_22835,N_21280,N_21416);
or U22836 (N_22836,N_21150,N_21354);
nand U22837 (N_22837,N_20313,N_20354);
nand U22838 (N_22838,N_20594,N_20050);
nand U22839 (N_22839,N_20123,N_20316);
and U22840 (N_22840,N_20041,N_20425);
and U22841 (N_22841,N_21790,N_20334);
or U22842 (N_22842,N_20161,N_21671);
nor U22843 (N_22843,N_20504,N_21805);
or U22844 (N_22844,N_21096,N_20973);
xnor U22845 (N_22845,N_20612,N_20174);
nor U22846 (N_22846,N_20133,N_20711);
and U22847 (N_22847,N_20211,N_21459);
or U22848 (N_22848,N_20861,N_21859);
nand U22849 (N_22849,N_20454,N_21775);
and U22850 (N_22850,N_20835,N_20806);
or U22851 (N_22851,N_21063,N_20533);
nor U22852 (N_22852,N_21110,N_21408);
xnor U22853 (N_22853,N_21910,N_21376);
xnor U22854 (N_22854,N_21461,N_21941);
xor U22855 (N_22855,N_21769,N_20907);
nor U22856 (N_22856,N_20905,N_20335);
and U22857 (N_22857,N_20096,N_20792);
and U22858 (N_22858,N_21223,N_20280);
and U22859 (N_22859,N_20634,N_21455);
nor U22860 (N_22860,N_21843,N_20169);
xnor U22861 (N_22861,N_21235,N_20463);
or U22862 (N_22862,N_20127,N_21266);
nand U22863 (N_22863,N_21466,N_20930);
and U22864 (N_22864,N_20702,N_20813);
xnor U22865 (N_22865,N_21443,N_20289);
xnor U22866 (N_22866,N_21987,N_20046);
and U22867 (N_22867,N_21933,N_20554);
nand U22868 (N_22868,N_20936,N_21282);
or U22869 (N_22869,N_21129,N_20444);
and U22870 (N_22870,N_21819,N_20682);
or U22871 (N_22871,N_20518,N_20168);
nand U22872 (N_22872,N_21834,N_20577);
or U22873 (N_22873,N_20845,N_20737);
xnor U22874 (N_22874,N_21172,N_20250);
and U22875 (N_22875,N_21564,N_20906);
or U22876 (N_22876,N_21552,N_21077);
nand U22877 (N_22877,N_20761,N_20325);
and U22878 (N_22878,N_20103,N_21425);
nor U22879 (N_22879,N_20391,N_21913);
or U22880 (N_22880,N_21863,N_21112);
and U22881 (N_22881,N_20195,N_21973);
and U22882 (N_22882,N_21267,N_20650);
nand U22883 (N_22883,N_21924,N_21071);
xnor U22884 (N_22884,N_20536,N_21060);
or U22885 (N_22885,N_21175,N_20735);
nor U22886 (N_22886,N_21464,N_20420);
nor U22887 (N_22887,N_21271,N_20020);
or U22888 (N_22888,N_20039,N_20807);
nand U22889 (N_22889,N_20215,N_21489);
or U22890 (N_22890,N_21386,N_20410);
nand U22891 (N_22891,N_21989,N_20308);
nor U22892 (N_22892,N_20971,N_21645);
or U22893 (N_22893,N_21252,N_21178);
nor U22894 (N_22894,N_21931,N_20225);
and U22895 (N_22895,N_21023,N_20698);
xnor U22896 (N_22896,N_21051,N_20998);
and U22897 (N_22897,N_20312,N_21607);
and U22898 (N_22898,N_21273,N_21140);
xor U22899 (N_22899,N_20688,N_21830);
nor U22900 (N_22900,N_20277,N_21748);
and U22901 (N_22901,N_21452,N_20357);
xnor U22902 (N_22902,N_20584,N_20914);
and U22903 (N_22903,N_21632,N_21048);
nor U22904 (N_22904,N_21639,N_21497);
nor U22905 (N_22905,N_21584,N_20055);
and U22906 (N_22906,N_21514,N_20462);
xor U22907 (N_22907,N_20224,N_20898);
xnor U22908 (N_22908,N_20119,N_20862);
xnor U22909 (N_22909,N_20824,N_20547);
nor U22910 (N_22910,N_20094,N_20453);
or U22911 (N_22911,N_21901,N_20878);
nand U22912 (N_22912,N_20394,N_21219);
nor U22913 (N_22913,N_20848,N_21020);
nand U22914 (N_22914,N_20748,N_20107);
xnor U22915 (N_22915,N_20180,N_21827);
or U22916 (N_22916,N_21598,N_20709);
xnor U22917 (N_22917,N_21559,N_20370);
xor U22918 (N_22918,N_21548,N_20885);
and U22919 (N_22919,N_20060,N_20925);
nand U22920 (N_22920,N_20822,N_20117);
nor U22921 (N_22921,N_20080,N_21400);
nor U22922 (N_22922,N_20773,N_20189);
xnor U22923 (N_22923,N_20768,N_21784);
or U22924 (N_22924,N_20817,N_20854);
nand U22925 (N_22925,N_20113,N_21069);
nand U22926 (N_22926,N_21194,N_21038);
and U22927 (N_22927,N_20011,N_21841);
nand U22928 (N_22928,N_20036,N_20422);
and U22929 (N_22929,N_21334,N_21660);
nor U22930 (N_22930,N_20424,N_20847);
nand U22931 (N_22931,N_21752,N_20149);
or U22932 (N_22932,N_20816,N_20040);
and U22933 (N_22933,N_21395,N_21184);
and U22934 (N_22934,N_20447,N_20940);
and U22935 (N_22935,N_21727,N_21504);
xor U22936 (N_22936,N_20258,N_21247);
or U22937 (N_22937,N_20079,N_21451);
or U22938 (N_22938,N_20765,N_21774);
xnor U22939 (N_22939,N_20757,N_21371);
nand U22940 (N_22940,N_21473,N_20072);
nand U22941 (N_22941,N_20044,N_20428);
nand U22942 (N_22942,N_20506,N_21746);
or U22943 (N_22943,N_20007,N_21169);
and U22944 (N_22944,N_20000,N_20575);
nor U22945 (N_22945,N_20286,N_21003);
and U22946 (N_22946,N_21324,N_20571);
nand U22947 (N_22947,N_21705,N_20347);
nand U22948 (N_22948,N_21797,N_21318);
or U22949 (N_22949,N_20214,N_21953);
or U22950 (N_22950,N_21328,N_20443);
or U22951 (N_22951,N_21067,N_21939);
or U22952 (N_22952,N_20882,N_21725);
and U22953 (N_22953,N_21203,N_21374);
nor U22954 (N_22954,N_21134,N_20519);
or U22955 (N_22955,N_20969,N_21599);
or U22956 (N_22956,N_21743,N_21848);
nand U22957 (N_22957,N_21511,N_20358);
xnor U22958 (N_22958,N_20276,N_20247);
nor U22959 (N_22959,N_21682,N_20886);
or U22960 (N_22960,N_20216,N_21454);
and U22961 (N_22961,N_21199,N_21406);
or U22962 (N_22962,N_20330,N_20786);
or U22963 (N_22963,N_21799,N_20670);
or U22964 (N_22964,N_21004,N_21105);
nand U22965 (N_22965,N_20618,N_20423);
and U22966 (N_22966,N_20609,N_21967);
and U22967 (N_22967,N_20857,N_21122);
or U22968 (N_22968,N_21714,N_21420);
or U22969 (N_22969,N_21782,N_21760);
nand U22970 (N_22970,N_21418,N_21915);
xnor U22971 (N_22971,N_20439,N_20111);
nor U22972 (N_22972,N_20110,N_21876);
nor U22973 (N_22973,N_21204,N_21081);
and U22974 (N_22974,N_21562,N_21778);
nor U22975 (N_22975,N_20182,N_21990);
nor U22976 (N_22976,N_21845,N_21969);
and U22977 (N_22977,N_20364,N_21168);
and U22978 (N_22978,N_20510,N_21820);
nand U22979 (N_22979,N_21779,N_20955);
and U22980 (N_22980,N_21190,N_20433);
nand U22981 (N_22981,N_21890,N_20846);
and U22982 (N_22982,N_21162,N_20531);
nor U22983 (N_22983,N_20284,N_21302);
nor U22984 (N_22984,N_21994,N_20679);
and U22985 (N_22985,N_20494,N_20323);
nand U22986 (N_22986,N_20034,N_21674);
nor U22987 (N_22987,N_20911,N_20937);
and U22988 (N_22988,N_21825,N_20029);
nor U22989 (N_22989,N_21265,N_20398);
and U22990 (N_22990,N_21215,N_20949);
or U22991 (N_22991,N_21300,N_21757);
xor U22992 (N_22992,N_20125,N_21786);
or U22993 (N_22993,N_20869,N_21932);
or U22994 (N_22994,N_20032,N_20621);
nor U22995 (N_22995,N_21314,N_20880);
nand U22996 (N_22996,N_20601,N_20294);
or U22997 (N_22997,N_21642,N_21898);
xnor U22998 (N_22998,N_21246,N_21027);
nand U22999 (N_22999,N_21291,N_20988);
nor U23000 (N_23000,N_21051,N_21201);
nand U23001 (N_23001,N_21545,N_20824);
nand U23002 (N_23002,N_20229,N_21289);
nand U23003 (N_23003,N_21657,N_21756);
nor U23004 (N_23004,N_21080,N_20728);
nand U23005 (N_23005,N_21430,N_21239);
nand U23006 (N_23006,N_21640,N_20099);
xor U23007 (N_23007,N_20334,N_21439);
or U23008 (N_23008,N_21789,N_20992);
nand U23009 (N_23009,N_20795,N_20608);
nand U23010 (N_23010,N_20801,N_20936);
or U23011 (N_23011,N_20409,N_21332);
nor U23012 (N_23012,N_20821,N_21538);
nand U23013 (N_23013,N_20186,N_20343);
and U23014 (N_23014,N_20091,N_21596);
and U23015 (N_23015,N_21852,N_21833);
or U23016 (N_23016,N_20404,N_20530);
xnor U23017 (N_23017,N_20892,N_21560);
nand U23018 (N_23018,N_20853,N_20594);
or U23019 (N_23019,N_20057,N_20265);
nand U23020 (N_23020,N_20917,N_20182);
or U23021 (N_23021,N_21717,N_20870);
or U23022 (N_23022,N_20482,N_21255);
xnor U23023 (N_23023,N_21943,N_21141);
nand U23024 (N_23024,N_21899,N_21925);
nor U23025 (N_23025,N_21462,N_21692);
xor U23026 (N_23026,N_21447,N_21752);
or U23027 (N_23027,N_21190,N_20253);
xor U23028 (N_23028,N_21904,N_20765);
and U23029 (N_23029,N_21203,N_21359);
nor U23030 (N_23030,N_21491,N_21247);
nor U23031 (N_23031,N_20645,N_20610);
nand U23032 (N_23032,N_21867,N_21480);
and U23033 (N_23033,N_20465,N_21915);
or U23034 (N_23034,N_20796,N_20754);
and U23035 (N_23035,N_21463,N_20589);
xor U23036 (N_23036,N_20289,N_21145);
xor U23037 (N_23037,N_20204,N_20968);
or U23038 (N_23038,N_20261,N_21026);
or U23039 (N_23039,N_20085,N_21670);
or U23040 (N_23040,N_21216,N_21021);
nor U23041 (N_23041,N_20760,N_20862);
and U23042 (N_23042,N_20320,N_20019);
nor U23043 (N_23043,N_21818,N_20626);
nor U23044 (N_23044,N_20925,N_20870);
or U23045 (N_23045,N_20430,N_21271);
and U23046 (N_23046,N_21400,N_20155);
nand U23047 (N_23047,N_21114,N_21640);
xor U23048 (N_23048,N_20035,N_20095);
or U23049 (N_23049,N_21955,N_20546);
and U23050 (N_23050,N_21415,N_20282);
and U23051 (N_23051,N_20967,N_21800);
or U23052 (N_23052,N_20260,N_20378);
or U23053 (N_23053,N_20899,N_21210);
xnor U23054 (N_23054,N_20641,N_21510);
nand U23055 (N_23055,N_20700,N_21864);
nand U23056 (N_23056,N_21363,N_21521);
nor U23057 (N_23057,N_20991,N_21430);
nor U23058 (N_23058,N_20865,N_20401);
nand U23059 (N_23059,N_20036,N_20346);
nand U23060 (N_23060,N_21802,N_20951);
nand U23061 (N_23061,N_20246,N_20861);
or U23062 (N_23062,N_21811,N_20028);
nor U23063 (N_23063,N_20737,N_21827);
and U23064 (N_23064,N_20831,N_20953);
nand U23065 (N_23065,N_21679,N_21897);
and U23066 (N_23066,N_20835,N_21572);
and U23067 (N_23067,N_21568,N_21565);
or U23068 (N_23068,N_21226,N_20931);
nand U23069 (N_23069,N_21291,N_20742);
and U23070 (N_23070,N_20178,N_20365);
nand U23071 (N_23071,N_20448,N_20146);
or U23072 (N_23072,N_21407,N_20906);
or U23073 (N_23073,N_21242,N_21839);
and U23074 (N_23074,N_20529,N_21935);
or U23075 (N_23075,N_21150,N_20574);
xnor U23076 (N_23076,N_20894,N_21905);
nor U23077 (N_23077,N_21548,N_20122);
or U23078 (N_23078,N_20577,N_20910);
xor U23079 (N_23079,N_21836,N_21917);
and U23080 (N_23080,N_20800,N_20219);
or U23081 (N_23081,N_20008,N_20220);
nor U23082 (N_23082,N_21216,N_21116);
nor U23083 (N_23083,N_21613,N_20860);
xnor U23084 (N_23084,N_21462,N_20784);
and U23085 (N_23085,N_20702,N_21427);
xnor U23086 (N_23086,N_21280,N_21007);
nor U23087 (N_23087,N_20488,N_21875);
or U23088 (N_23088,N_20246,N_21279);
or U23089 (N_23089,N_20736,N_20673);
and U23090 (N_23090,N_21020,N_20554);
and U23091 (N_23091,N_20326,N_20217);
or U23092 (N_23092,N_21371,N_20251);
and U23093 (N_23093,N_21127,N_21626);
and U23094 (N_23094,N_20920,N_20147);
nand U23095 (N_23095,N_20325,N_20550);
nor U23096 (N_23096,N_21525,N_20030);
nand U23097 (N_23097,N_20717,N_21517);
or U23098 (N_23098,N_20149,N_21599);
xor U23099 (N_23099,N_21164,N_21978);
or U23100 (N_23100,N_20206,N_20981);
xor U23101 (N_23101,N_20483,N_21206);
nor U23102 (N_23102,N_20601,N_21682);
and U23103 (N_23103,N_20909,N_20377);
or U23104 (N_23104,N_21823,N_21446);
and U23105 (N_23105,N_21437,N_20918);
nand U23106 (N_23106,N_21111,N_20356);
xor U23107 (N_23107,N_21636,N_20476);
nor U23108 (N_23108,N_20826,N_21690);
nand U23109 (N_23109,N_21751,N_21278);
or U23110 (N_23110,N_21519,N_20074);
nand U23111 (N_23111,N_20735,N_20434);
nor U23112 (N_23112,N_20963,N_20825);
nor U23113 (N_23113,N_20246,N_20494);
and U23114 (N_23114,N_21762,N_20231);
or U23115 (N_23115,N_21266,N_20278);
xnor U23116 (N_23116,N_21975,N_20258);
nor U23117 (N_23117,N_20627,N_21024);
and U23118 (N_23118,N_21332,N_20551);
nand U23119 (N_23119,N_20800,N_20508);
nor U23120 (N_23120,N_20610,N_21055);
or U23121 (N_23121,N_20612,N_20874);
xor U23122 (N_23122,N_21167,N_20552);
and U23123 (N_23123,N_20682,N_21504);
nor U23124 (N_23124,N_20174,N_21410);
nand U23125 (N_23125,N_21942,N_21117);
xor U23126 (N_23126,N_21453,N_20768);
or U23127 (N_23127,N_20763,N_21081);
nand U23128 (N_23128,N_20053,N_21618);
or U23129 (N_23129,N_20276,N_20971);
nor U23130 (N_23130,N_20549,N_21454);
or U23131 (N_23131,N_21517,N_20274);
nand U23132 (N_23132,N_20720,N_20070);
or U23133 (N_23133,N_20581,N_21875);
nor U23134 (N_23134,N_20075,N_20221);
nand U23135 (N_23135,N_21928,N_20656);
xnor U23136 (N_23136,N_21799,N_20565);
or U23137 (N_23137,N_21604,N_21817);
nor U23138 (N_23138,N_21645,N_21257);
and U23139 (N_23139,N_20610,N_20619);
and U23140 (N_23140,N_20386,N_20845);
xnor U23141 (N_23141,N_20303,N_21621);
xnor U23142 (N_23142,N_20255,N_21424);
nand U23143 (N_23143,N_21923,N_20158);
or U23144 (N_23144,N_20204,N_21738);
nand U23145 (N_23145,N_21431,N_20772);
xor U23146 (N_23146,N_20254,N_21974);
nand U23147 (N_23147,N_20641,N_20581);
and U23148 (N_23148,N_21286,N_21361);
nand U23149 (N_23149,N_20526,N_21761);
nand U23150 (N_23150,N_20996,N_21323);
or U23151 (N_23151,N_21399,N_20974);
nor U23152 (N_23152,N_21311,N_20644);
and U23153 (N_23153,N_20105,N_21091);
nor U23154 (N_23154,N_20682,N_21267);
or U23155 (N_23155,N_20111,N_20156);
and U23156 (N_23156,N_20229,N_20180);
and U23157 (N_23157,N_21730,N_20567);
or U23158 (N_23158,N_20546,N_20194);
or U23159 (N_23159,N_20216,N_21964);
nand U23160 (N_23160,N_21023,N_20429);
nor U23161 (N_23161,N_21809,N_21191);
or U23162 (N_23162,N_20585,N_20284);
or U23163 (N_23163,N_20120,N_21624);
and U23164 (N_23164,N_21373,N_21391);
or U23165 (N_23165,N_21555,N_21485);
xor U23166 (N_23166,N_20222,N_21457);
nor U23167 (N_23167,N_20397,N_20682);
and U23168 (N_23168,N_20825,N_21005);
or U23169 (N_23169,N_21425,N_21941);
nand U23170 (N_23170,N_20312,N_21702);
nand U23171 (N_23171,N_20660,N_21294);
nand U23172 (N_23172,N_20964,N_20986);
or U23173 (N_23173,N_20228,N_21226);
and U23174 (N_23174,N_20652,N_20426);
or U23175 (N_23175,N_20089,N_20052);
nor U23176 (N_23176,N_21868,N_20546);
or U23177 (N_23177,N_20065,N_21554);
and U23178 (N_23178,N_21768,N_20160);
and U23179 (N_23179,N_20172,N_20624);
nor U23180 (N_23180,N_20139,N_21744);
xnor U23181 (N_23181,N_20043,N_21022);
xor U23182 (N_23182,N_20963,N_20799);
xor U23183 (N_23183,N_21800,N_20928);
xnor U23184 (N_23184,N_21901,N_20657);
or U23185 (N_23185,N_21871,N_20854);
nand U23186 (N_23186,N_21386,N_21674);
nor U23187 (N_23187,N_21146,N_20804);
nand U23188 (N_23188,N_20225,N_21745);
nor U23189 (N_23189,N_20779,N_20381);
nand U23190 (N_23190,N_21985,N_20041);
xnor U23191 (N_23191,N_20662,N_21504);
xnor U23192 (N_23192,N_20196,N_21734);
and U23193 (N_23193,N_20711,N_21977);
nor U23194 (N_23194,N_20357,N_21251);
or U23195 (N_23195,N_21626,N_21952);
nor U23196 (N_23196,N_21410,N_20017);
and U23197 (N_23197,N_20178,N_20366);
xor U23198 (N_23198,N_20266,N_20688);
nor U23199 (N_23199,N_21512,N_21838);
nand U23200 (N_23200,N_20489,N_21764);
and U23201 (N_23201,N_21415,N_20268);
nor U23202 (N_23202,N_20897,N_20995);
or U23203 (N_23203,N_20834,N_21490);
or U23204 (N_23204,N_21142,N_20657);
nand U23205 (N_23205,N_20216,N_21938);
nand U23206 (N_23206,N_20961,N_21727);
nor U23207 (N_23207,N_20718,N_21422);
or U23208 (N_23208,N_21706,N_20514);
xor U23209 (N_23209,N_20743,N_21814);
or U23210 (N_23210,N_20614,N_21606);
xnor U23211 (N_23211,N_20540,N_21430);
or U23212 (N_23212,N_20255,N_20053);
nor U23213 (N_23213,N_20465,N_20395);
or U23214 (N_23214,N_20683,N_21121);
nor U23215 (N_23215,N_20154,N_21802);
and U23216 (N_23216,N_20616,N_20944);
or U23217 (N_23217,N_21196,N_21486);
nand U23218 (N_23218,N_21840,N_21331);
xor U23219 (N_23219,N_21716,N_21785);
or U23220 (N_23220,N_20477,N_20995);
and U23221 (N_23221,N_20779,N_21199);
nand U23222 (N_23222,N_21110,N_20700);
nand U23223 (N_23223,N_20137,N_20811);
and U23224 (N_23224,N_20350,N_20019);
or U23225 (N_23225,N_21714,N_21696);
nor U23226 (N_23226,N_21344,N_20572);
and U23227 (N_23227,N_21524,N_20191);
nand U23228 (N_23228,N_21335,N_20315);
nor U23229 (N_23229,N_21626,N_21566);
nand U23230 (N_23230,N_20586,N_20058);
nand U23231 (N_23231,N_21664,N_21828);
and U23232 (N_23232,N_21353,N_21056);
nand U23233 (N_23233,N_21557,N_20193);
nand U23234 (N_23234,N_20059,N_21574);
nand U23235 (N_23235,N_20996,N_21080);
or U23236 (N_23236,N_21745,N_21496);
nor U23237 (N_23237,N_21447,N_21498);
or U23238 (N_23238,N_20455,N_21399);
nor U23239 (N_23239,N_21742,N_20734);
nand U23240 (N_23240,N_20303,N_21960);
or U23241 (N_23241,N_20082,N_20534);
nor U23242 (N_23242,N_20953,N_21905);
nand U23243 (N_23243,N_21555,N_20454);
xor U23244 (N_23244,N_21058,N_21536);
and U23245 (N_23245,N_20894,N_21941);
nor U23246 (N_23246,N_20947,N_20130);
nor U23247 (N_23247,N_20015,N_21153);
or U23248 (N_23248,N_21535,N_20913);
xnor U23249 (N_23249,N_21689,N_20300);
xor U23250 (N_23250,N_20115,N_20087);
or U23251 (N_23251,N_21968,N_21991);
and U23252 (N_23252,N_20940,N_20421);
nor U23253 (N_23253,N_21068,N_21422);
or U23254 (N_23254,N_21504,N_20381);
nor U23255 (N_23255,N_20708,N_20129);
xor U23256 (N_23256,N_20204,N_21270);
nor U23257 (N_23257,N_21065,N_20856);
and U23258 (N_23258,N_21088,N_20841);
and U23259 (N_23259,N_20127,N_21453);
or U23260 (N_23260,N_20304,N_20892);
or U23261 (N_23261,N_21589,N_20069);
nor U23262 (N_23262,N_20932,N_20740);
or U23263 (N_23263,N_21023,N_20110);
xor U23264 (N_23264,N_20950,N_20014);
or U23265 (N_23265,N_20260,N_20471);
xor U23266 (N_23266,N_21305,N_21953);
and U23267 (N_23267,N_20090,N_20524);
nand U23268 (N_23268,N_20143,N_21141);
or U23269 (N_23269,N_21678,N_20444);
nand U23270 (N_23270,N_20252,N_20328);
and U23271 (N_23271,N_20737,N_21397);
and U23272 (N_23272,N_20086,N_20407);
nand U23273 (N_23273,N_21261,N_20100);
nand U23274 (N_23274,N_21932,N_20855);
nor U23275 (N_23275,N_21263,N_21584);
and U23276 (N_23276,N_20443,N_20310);
or U23277 (N_23277,N_21643,N_20470);
xor U23278 (N_23278,N_20497,N_20042);
nand U23279 (N_23279,N_21495,N_21623);
and U23280 (N_23280,N_20197,N_20987);
xnor U23281 (N_23281,N_21497,N_21005);
nand U23282 (N_23282,N_20855,N_20073);
xor U23283 (N_23283,N_21563,N_21663);
or U23284 (N_23284,N_21350,N_20767);
and U23285 (N_23285,N_20696,N_21778);
nand U23286 (N_23286,N_21714,N_20660);
xor U23287 (N_23287,N_21804,N_20738);
or U23288 (N_23288,N_20093,N_21814);
or U23289 (N_23289,N_20374,N_20043);
or U23290 (N_23290,N_20349,N_20958);
nor U23291 (N_23291,N_21158,N_20533);
nor U23292 (N_23292,N_21998,N_20483);
xnor U23293 (N_23293,N_21604,N_20441);
nand U23294 (N_23294,N_21697,N_20443);
and U23295 (N_23295,N_21922,N_20366);
and U23296 (N_23296,N_20965,N_20114);
nand U23297 (N_23297,N_21238,N_20123);
or U23298 (N_23298,N_21773,N_21898);
or U23299 (N_23299,N_20270,N_20414);
xor U23300 (N_23300,N_20760,N_21974);
and U23301 (N_23301,N_21642,N_20408);
xor U23302 (N_23302,N_20281,N_20056);
nor U23303 (N_23303,N_20824,N_20420);
nor U23304 (N_23304,N_20038,N_20089);
xor U23305 (N_23305,N_20782,N_21638);
nand U23306 (N_23306,N_20818,N_21252);
nand U23307 (N_23307,N_20787,N_20556);
nand U23308 (N_23308,N_20009,N_21906);
or U23309 (N_23309,N_20699,N_21860);
nand U23310 (N_23310,N_20598,N_21472);
and U23311 (N_23311,N_21722,N_21637);
nor U23312 (N_23312,N_21430,N_20590);
nand U23313 (N_23313,N_20392,N_20902);
and U23314 (N_23314,N_21911,N_21492);
and U23315 (N_23315,N_20073,N_21642);
or U23316 (N_23316,N_21043,N_20834);
xnor U23317 (N_23317,N_20874,N_20804);
nand U23318 (N_23318,N_20827,N_21298);
nor U23319 (N_23319,N_20271,N_20206);
xnor U23320 (N_23320,N_21981,N_20254);
and U23321 (N_23321,N_21188,N_21025);
xor U23322 (N_23322,N_20815,N_20054);
nand U23323 (N_23323,N_20328,N_21333);
nor U23324 (N_23324,N_21363,N_21970);
or U23325 (N_23325,N_20519,N_20454);
nor U23326 (N_23326,N_21528,N_20791);
and U23327 (N_23327,N_20922,N_21006);
nor U23328 (N_23328,N_21048,N_20553);
nor U23329 (N_23329,N_21441,N_20076);
xor U23330 (N_23330,N_21213,N_20205);
nand U23331 (N_23331,N_20209,N_20145);
or U23332 (N_23332,N_20682,N_20370);
nor U23333 (N_23333,N_20979,N_20594);
or U23334 (N_23334,N_21753,N_20608);
or U23335 (N_23335,N_21640,N_20754);
nor U23336 (N_23336,N_21022,N_21760);
and U23337 (N_23337,N_21004,N_20866);
nand U23338 (N_23338,N_21369,N_21473);
or U23339 (N_23339,N_21799,N_20722);
nor U23340 (N_23340,N_20192,N_20172);
or U23341 (N_23341,N_21282,N_20042);
or U23342 (N_23342,N_20220,N_21803);
nand U23343 (N_23343,N_20655,N_20574);
or U23344 (N_23344,N_21619,N_20404);
and U23345 (N_23345,N_21998,N_20927);
xor U23346 (N_23346,N_20767,N_21946);
and U23347 (N_23347,N_21453,N_21547);
and U23348 (N_23348,N_21888,N_20145);
nand U23349 (N_23349,N_20142,N_20983);
nor U23350 (N_23350,N_20897,N_21765);
nor U23351 (N_23351,N_21028,N_20942);
or U23352 (N_23352,N_21677,N_20372);
nand U23353 (N_23353,N_20301,N_21106);
nand U23354 (N_23354,N_20219,N_21282);
xnor U23355 (N_23355,N_21975,N_20975);
xnor U23356 (N_23356,N_21941,N_20724);
nor U23357 (N_23357,N_21487,N_21567);
and U23358 (N_23358,N_20606,N_20304);
xor U23359 (N_23359,N_20860,N_20821);
nand U23360 (N_23360,N_21511,N_21492);
nor U23361 (N_23361,N_21021,N_20659);
nor U23362 (N_23362,N_21842,N_20635);
nor U23363 (N_23363,N_20570,N_21389);
nand U23364 (N_23364,N_20735,N_21856);
nand U23365 (N_23365,N_20706,N_20227);
or U23366 (N_23366,N_21131,N_20738);
nand U23367 (N_23367,N_21508,N_21309);
nand U23368 (N_23368,N_21740,N_20246);
nand U23369 (N_23369,N_20664,N_20793);
xnor U23370 (N_23370,N_21995,N_20722);
and U23371 (N_23371,N_21747,N_21797);
xor U23372 (N_23372,N_20633,N_21658);
xor U23373 (N_23373,N_20456,N_20543);
nand U23374 (N_23374,N_21949,N_21296);
nor U23375 (N_23375,N_21821,N_21097);
and U23376 (N_23376,N_21077,N_21026);
nor U23377 (N_23377,N_20497,N_20445);
or U23378 (N_23378,N_20490,N_20552);
xor U23379 (N_23379,N_20947,N_21298);
or U23380 (N_23380,N_20911,N_20657);
and U23381 (N_23381,N_21036,N_21395);
and U23382 (N_23382,N_20524,N_20226);
and U23383 (N_23383,N_21468,N_20038);
nand U23384 (N_23384,N_20112,N_21426);
nand U23385 (N_23385,N_21787,N_20936);
xor U23386 (N_23386,N_20373,N_20089);
or U23387 (N_23387,N_20274,N_21173);
xor U23388 (N_23388,N_21517,N_20747);
or U23389 (N_23389,N_21330,N_21652);
and U23390 (N_23390,N_21180,N_20374);
xor U23391 (N_23391,N_21615,N_20314);
nand U23392 (N_23392,N_20948,N_20832);
and U23393 (N_23393,N_20593,N_20133);
nor U23394 (N_23394,N_21253,N_20008);
and U23395 (N_23395,N_21144,N_20785);
and U23396 (N_23396,N_21983,N_21276);
or U23397 (N_23397,N_21387,N_21926);
nand U23398 (N_23398,N_21619,N_21725);
or U23399 (N_23399,N_21698,N_20728);
nor U23400 (N_23400,N_20854,N_21579);
nor U23401 (N_23401,N_21105,N_21802);
xor U23402 (N_23402,N_20162,N_21230);
xnor U23403 (N_23403,N_21720,N_20494);
nand U23404 (N_23404,N_21233,N_21855);
nor U23405 (N_23405,N_20505,N_21227);
and U23406 (N_23406,N_21323,N_20663);
and U23407 (N_23407,N_20533,N_20523);
and U23408 (N_23408,N_21316,N_21614);
xor U23409 (N_23409,N_21160,N_21318);
nor U23410 (N_23410,N_21257,N_20852);
and U23411 (N_23411,N_20035,N_21075);
and U23412 (N_23412,N_21717,N_20971);
nand U23413 (N_23413,N_21993,N_20922);
nor U23414 (N_23414,N_20390,N_21443);
xnor U23415 (N_23415,N_20915,N_20867);
and U23416 (N_23416,N_20576,N_21164);
xor U23417 (N_23417,N_20660,N_21905);
nand U23418 (N_23418,N_21060,N_20860);
nand U23419 (N_23419,N_21500,N_21990);
nor U23420 (N_23420,N_20584,N_20815);
and U23421 (N_23421,N_20630,N_21772);
xor U23422 (N_23422,N_21081,N_20797);
nand U23423 (N_23423,N_20967,N_21465);
xor U23424 (N_23424,N_20518,N_21018);
nor U23425 (N_23425,N_20852,N_20378);
and U23426 (N_23426,N_20056,N_20152);
and U23427 (N_23427,N_21101,N_21995);
and U23428 (N_23428,N_20730,N_20344);
xor U23429 (N_23429,N_20896,N_20870);
and U23430 (N_23430,N_20035,N_21916);
nor U23431 (N_23431,N_21574,N_21559);
xnor U23432 (N_23432,N_20367,N_20825);
xnor U23433 (N_23433,N_21264,N_21521);
xor U23434 (N_23434,N_21894,N_20425);
nor U23435 (N_23435,N_20859,N_20204);
nand U23436 (N_23436,N_20025,N_21844);
and U23437 (N_23437,N_21924,N_21145);
nand U23438 (N_23438,N_20153,N_21616);
xnor U23439 (N_23439,N_21509,N_20972);
or U23440 (N_23440,N_20313,N_20834);
xor U23441 (N_23441,N_21028,N_20061);
xor U23442 (N_23442,N_20183,N_21290);
or U23443 (N_23443,N_21068,N_21723);
xor U23444 (N_23444,N_20448,N_20956);
or U23445 (N_23445,N_20838,N_20058);
and U23446 (N_23446,N_20045,N_21068);
nand U23447 (N_23447,N_21250,N_20005);
or U23448 (N_23448,N_21993,N_21772);
nand U23449 (N_23449,N_21704,N_20966);
or U23450 (N_23450,N_21786,N_21551);
xor U23451 (N_23451,N_21804,N_20480);
xnor U23452 (N_23452,N_21232,N_21005);
and U23453 (N_23453,N_20885,N_20192);
nor U23454 (N_23454,N_21075,N_20830);
or U23455 (N_23455,N_21795,N_20223);
or U23456 (N_23456,N_20990,N_21714);
and U23457 (N_23457,N_21911,N_21182);
xnor U23458 (N_23458,N_21233,N_21806);
xor U23459 (N_23459,N_20716,N_20800);
and U23460 (N_23460,N_20599,N_21329);
nand U23461 (N_23461,N_20714,N_20014);
or U23462 (N_23462,N_20555,N_21636);
or U23463 (N_23463,N_21216,N_21520);
xnor U23464 (N_23464,N_21437,N_21132);
nor U23465 (N_23465,N_20893,N_21009);
or U23466 (N_23466,N_21682,N_20130);
and U23467 (N_23467,N_20582,N_20364);
xnor U23468 (N_23468,N_20117,N_20478);
nor U23469 (N_23469,N_20296,N_21032);
nor U23470 (N_23470,N_20884,N_20901);
nor U23471 (N_23471,N_20333,N_20302);
or U23472 (N_23472,N_20022,N_21760);
nand U23473 (N_23473,N_20719,N_21794);
nand U23474 (N_23474,N_20445,N_21054);
xnor U23475 (N_23475,N_21688,N_20955);
and U23476 (N_23476,N_20163,N_20790);
nand U23477 (N_23477,N_21352,N_20182);
and U23478 (N_23478,N_21542,N_20950);
xnor U23479 (N_23479,N_20083,N_20023);
nand U23480 (N_23480,N_21819,N_21270);
nor U23481 (N_23481,N_20931,N_21881);
or U23482 (N_23482,N_21235,N_21581);
nor U23483 (N_23483,N_21900,N_20718);
nand U23484 (N_23484,N_21772,N_21698);
and U23485 (N_23485,N_20246,N_20330);
nor U23486 (N_23486,N_21993,N_20204);
and U23487 (N_23487,N_21321,N_20250);
or U23488 (N_23488,N_21750,N_20935);
and U23489 (N_23489,N_21838,N_20672);
or U23490 (N_23490,N_21917,N_21919);
and U23491 (N_23491,N_21959,N_20208);
or U23492 (N_23492,N_21849,N_20824);
nor U23493 (N_23493,N_21466,N_21371);
and U23494 (N_23494,N_20669,N_20571);
nand U23495 (N_23495,N_20549,N_20971);
or U23496 (N_23496,N_21823,N_21245);
nor U23497 (N_23497,N_20010,N_20966);
nor U23498 (N_23498,N_20797,N_21753);
and U23499 (N_23499,N_20830,N_21202);
and U23500 (N_23500,N_21080,N_20725);
xor U23501 (N_23501,N_21726,N_20553);
nand U23502 (N_23502,N_21160,N_20600);
or U23503 (N_23503,N_21668,N_20159);
and U23504 (N_23504,N_20421,N_20995);
nand U23505 (N_23505,N_21803,N_21901);
xor U23506 (N_23506,N_20444,N_20178);
nor U23507 (N_23507,N_20208,N_21747);
nand U23508 (N_23508,N_21181,N_20959);
xor U23509 (N_23509,N_20646,N_20071);
or U23510 (N_23510,N_20738,N_20596);
or U23511 (N_23511,N_21605,N_20459);
nor U23512 (N_23512,N_21413,N_20064);
nand U23513 (N_23513,N_20619,N_20120);
and U23514 (N_23514,N_21885,N_20833);
xor U23515 (N_23515,N_21765,N_20123);
nand U23516 (N_23516,N_20265,N_21846);
nor U23517 (N_23517,N_20881,N_21012);
nand U23518 (N_23518,N_21634,N_21183);
nand U23519 (N_23519,N_21608,N_21143);
and U23520 (N_23520,N_20231,N_21064);
nand U23521 (N_23521,N_20738,N_21891);
nand U23522 (N_23522,N_21714,N_21021);
nor U23523 (N_23523,N_20008,N_21447);
or U23524 (N_23524,N_20391,N_20880);
nand U23525 (N_23525,N_20532,N_21152);
nor U23526 (N_23526,N_21500,N_21523);
and U23527 (N_23527,N_21351,N_21474);
or U23528 (N_23528,N_20628,N_20594);
or U23529 (N_23529,N_21099,N_21401);
nor U23530 (N_23530,N_20499,N_21831);
and U23531 (N_23531,N_20276,N_21690);
nand U23532 (N_23532,N_20543,N_21131);
nand U23533 (N_23533,N_21947,N_21662);
and U23534 (N_23534,N_20725,N_21046);
xnor U23535 (N_23535,N_20617,N_20439);
and U23536 (N_23536,N_20420,N_20746);
and U23537 (N_23537,N_21283,N_21109);
xor U23538 (N_23538,N_21821,N_20233);
nand U23539 (N_23539,N_20951,N_20770);
or U23540 (N_23540,N_20138,N_20873);
or U23541 (N_23541,N_20600,N_20907);
nor U23542 (N_23542,N_21200,N_21266);
and U23543 (N_23543,N_20844,N_21302);
nor U23544 (N_23544,N_20434,N_20277);
nor U23545 (N_23545,N_21642,N_20926);
and U23546 (N_23546,N_20071,N_20047);
nand U23547 (N_23547,N_21895,N_20324);
nand U23548 (N_23548,N_20827,N_20987);
or U23549 (N_23549,N_21303,N_20244);
nor U23550 (N_23550,N_21396,N_20739);
nand U23551 (N_23551,N_21790,N_20137);
nor U23552 (N_23552,N_21293,N_21027);
nand U23553 (N_23553,N_21843,N_21381);
and U23554 (N_23554,N_21767,N_20852);
or U23555 (N_23555,N_20469,N_20522);
or U23556 (N_23556,N_20732,N_21432);
and U23557 (N_23557,N_20447,N_21660);
xor U23558 (N_23558,N_20264,N_20508);
or U23559 (N_23559,N_21355,N_20938);
xnor U23560 (N_23560,N_21358,N_21038);
or U23561 (N_23561,N_20311,N_21230);
or U23562 (N_23562,N_21001,N_20878);
nor U23563 (N_23563,N_20569,N_21261);
nand U23564 (N_23564,N_20026,N_20070);
and U23565 (N_23565,N_20026,N_20030);
nor U23566 (N_23566,N_21070,N_21107);
nand U23567 (N_23567,N_21116,N_21850);
xnor U23568 (N_23568,N_20718,N_21611);
or U23569 (N_23569,N_21637,N_20395);
nor U23570 (N_23570,N_21867,N_21968);
and U23571 (N_23571,N_20702,N_21388);
and U23572 (N_23572,N_21015,N_20912);
or U23573 (N_23573,N_21892,N_20555);
xnor U23574 (N_23574,N_21726,N_20366);
nand U23575 (N_23575,N_20228,N_20550);
or U23576 (N_23576,N_20290,N_21945);
nand U23577 (N_23577,N_21863,N_21279);
nand U23578 (N_23578,N_20509,N_20020);
xnor U23579 (N_23579,N_20554,N_20875);
nand U23580 (N_23580,N_20125,N_21733);
nor U23581 (N_23581,N_21061,N_21519);
or U23582 (N_23582,N_21876,N_21589);
xnor U23583 (N_23583,N_21463,N_21275);
nand U23584 (N_23584,N_21866,N_21559);
nor U23585 (N_23585,N_20929,N_20822);
or U23586 (N_23586,N_20475,N_21585);
or U23587 (N_23587,N_21906,N_20757);
and U23588 (N_23588,N_20082,N_21326);
nand U23589 (N_23589,N_21899,N_20137);
xor U23590 (N_23590,N_21184,N_20105);
nor U23591 (N_23591,N_21924,N_21295);
nand U23592 (N_23592,N_20114,N_21443);
nor U23593 (N_23593,N_21242,N_21434);
xor U23594 (N_23594,N_20049,N_21523);
nor U23595 (N_23595,N_20523,N_20306);
nor U23596 (N_23596,N_21609,N_20916);
nand U23597 (N_23597,N_20864,N_21038);
nand U23598 (N_23598,N_20447,N_21512);
and U23599 (N_23599,N_21309,N_20118);
nand U23600 (N_23600,N_21226,N_20378);
and U23601 (N_23601,N_21770,N_20378);
nand U23602 (N_23602,N_20634,N_21249);
nor U23603 (N_23603,N_20444,N_21324);
xnor U23604 (N_23604,N_20918,N_20034);
xor U23605 (N_23605,N_21435,N_21495);
xor U23606 (N_23606,N_20835,N_21462);
nor U23607 (N_23607,N_21177,N_20020);
nor U23608 (N_23608,N_21157,N_21159);
xnor U23609 (N_23609,N_20474,N_21656);
and U23610 (N_23610,N_20173,N_20139);
nor U23611 (N_23611,N_21580,N_20766);
nor U23612 (N_23612,N_20132,N_20406);
nor U23613 (N_23613,N_20302,N_21879);
or U23614 (N_23614,N_21547,N_20178);
nand U23615 (N_23615,N_20666,N_20861);
and U23616 (N_23616,N_21268,N_21296);
nor U23617 (N_23617,N_21615,N_21835);
nand U23618 (N_23618,N_20854,N_20271);
nor U23619 (N_23619,N_21206,N_20852);
nand U23620 (N_23620,N_21915,N_20908);
nand U23621 (N_23621,N_21747,N_21530);
nor U23622 (N_23622,N_20032,N_21704);
and U23623 (N_23623,N_21701,N_20347);
nor U23624 (N_23624,N_20293,N_20397);
nor U23625 (N_23625,N_20509,N_20983);
and U23626 (N_23626,N_21791,N_20612);
nand U23627 (N_23627,N_21213,N_20309);
xor U23628 (N_23628,N_20737,N_21559);
or U23629 (N_23629,N_21268,N_21978);
nor U23630 (N_23630,N_20336,N_20243);
or U23631 (N_23631,N_20259,N_20281);
xnor U23632 (N_23632,N_20030,N_20528);
or U23633 (N_23633,N_21609,N_20654);
xnor U23634 (N_23634,N_21184,N_20733);
nor U23635 (N_23635,N_20745,N_21397);
and U23636 (N_23636,N_20087,N_21798);
nor U23637 (N_23637,N_21225,N_20470);
xnor U23638 (N_23638,N_21673,N_21284);
nor U23639 (N_23639,N_20377,N_20226);
nor U23640 (N_23640,N_20986,N_20271);
nand U23641 (N_23641,N_21637,N_20662);
nand U23642 (N_23642,N_21907,N_21214);
nand U23643 (N_23643,N_21498,N_20014);
xnor U23644 (N_23644,N_20021,N_21330);
nor U23645 (N_23645,N_20149,N_20077);
nor U23646 (N_23646,N_20567,N_21112);
and U23647 (N_23647,N_21679,N_20649);
and U23648 (N_23648,N_20597,N_20199);
and U23649 (N_23649,N_21843,N_20295);
or U23650 (N_23650,N_21450,N_20057);
and U23651 (N_23651,N_20527,N_21040);
nor U23652 (N_23652,N_21407,N_20733);
and U23653 (N_23653,N_21561,N_21811);
xor U23654 (N_23654,N_20063,N_21514);
nor U23655 (N_23655,N_20665,N_20915);
nor U23656 (N_23656,N_20470,N_20976);
xor U23657 (N_23657,N_21702,N_20353);
xor U23658 (N_23658,N_21854,N_20702);
and U23659 (N_23659,N_21375,N_20834);
nor U23660 (N_23660,N_21175,N_20979);
or U23661 (N_23661,N_20768,N_21248);
xnor U23662 (N_23662,N_20005,N_20812);
or U23663 (N_23663,N_21799,N_20503);
nor U23664 (N_23664,N_20566,N_20725);
nor U23665 (N_23665,N_21703,N_20465);
nand U23666 (N_23666,N_21230,N_20959);
and U23667 (N_23667,N_20642,N_20504);
or U23668 (N_23668,N_20024,N_21360);
nand U23669 (N_23669,N_20567,N_20031);
nor U23670 (N_23670,N_21180,N_20760);
nor U23671 (N_23671,N_21171,N_20666);
and U23672 (N_23672,N_20630,N_20384);
nor U23673 (N_23673,N_20793,N_21801);
and U23674 (N_23674,N_20068,N_21931);
xor U23675 (N_23675,N_21485,N_21916);
and U23676 (N_23676,N_20938,N_20463);
xor U23677 (N_23677,N_20776,N_21377);
nand U23678 (N_23678,N_20630,N_21752);
or U23679 (N_23679,N_20742,N_20764);
nor U23680 (N_23680,N_20462,N_20870);
xnor U23681 (N_23681,N_21950,N_20297);
xor U23682 (N_23682,N_21247,N_21456);
or U23683 (N_23683,N_20314,N_21733);
or U23684 (N_23684,N_21914,N_20296);
nor U23685 (N_23685,N_20121,N_20036);
nor U23686 (N_23686,N_21078,N_21964);
xor U23687 (N_23687,N_20062,N_20958);
nand U23688 (N_23688,N_21027,N_21077);
nand U23689 (N_23689,N_20666,N_20081);
nand U23690 (N_23690,N_20688,N_21640);
and U23691 (N_23691,N_20705,N_21902);
xor U23692 (N_23692,N_20525,N_21701);
and U23693 (N_23693,N_21420,N_21597);
and U23694 (N_23694,N_20640,N_20422);
and U23695 (N_23695,N_21267,N_20493);
xnor U23696 (N_23696,N_20008,N_20893);
xnor U23697 (N_23697,N_21812,N_21423);
nand U23698 (N_23698,N_20054,N_20027);
or U23699 (N_23699,N_21494,N_20317);
nor U23700 (N_23700,N_20756,N_20484);
nor U23701 (N_23701,N_20878,N_21627);
and U23702 (N_23702,N_20481,N_20353);
nand U23703 (N_23703,N_21592,N_20411);
nand U23704 (N_23704,N_21990,N_21460);
nor U23705 (N_23705,N_20693,N_20675);
nand U23706 (N_23706,N_21700,N_20214);
or U23707 (N_23707,N_20471,N_21707);
and U23708 (N_23708,N_21773,N_21318);
nor U23709 (N_23709,N_21526,N_21938);
nand U23710 (N_23710,N_20565,N_21006);
nand U23711 (N_23711,N_21202,N_21860);
and U23712 (N_23712,N_21185,N_21902);
or U23713 (N_23713,N_21422,N_21130);
nor U23714 (N_23714,N_20434,N_21408);
or U23715 (N_23715,N_21946,N_20777);
nor U23716 (N_23716,N_20304,N_20253);
xnor U23717 (N_23717,N_20092,N_20611);
or U23718 (N_23718,N_20572,N_21420);
or U23719 (N_23719,N_20240,N_20211);
nand U23720 (N_23720,N_21164,N_21979);
or U23721 (N_23721,N_20783,N_20651);
nor U23722 (N_23722,N_20469,N_21558);
nor U23723 (N_23723,N_20800,N_20084);
nor U23724 (N_23724,N_20314,N_21247);
xor U23725 (N_23725,N_20010,N_20098);
or U23726 (N_23726,N_20207,N_21788);
and U23727 (N_23727,N_20750,N_21960);
nor U23728 (N_23728,N_20488,N_20161);
nor U23729 (N_23729,N_21822,N_21919);
or U23730 (N_23730,N_20939,N_21419);
nand U23731 (N_23731,N_21265,N_21066);
nor U23732 (N_23732,N_20957,N_20339);
xor U23733 (N_23733,N_21803,N_20132);
nand U23734 (N_23734,N_21290,N_21421);
and U23735 (N_23735,N_20403,N_21232);
xnor U23736 (N_23736,N_21599,N_21093);
nand U23737 (N_23737,N_20460,N_21950);
or U23738 (N_23738,N_20282,N_21805);
nor U23739 (N_23739,N_21819,N_20631);
and U23740 (N_23740,N_20664,N_20566);
xor U23741 (N_23741,N_20231,N_20341);
nor U23742 (N_23742,N_20120,N_20385);
nor U23743 (N_23743,N_20248,N_21307);
xor U23744 (N_23744,N_21246,N_21186);
xor U23745 (N_23745,N_20239,N_21540);
nand U23746 (N_23746,N_21478,N_21179);
nor U23747 (N_23747,N_20428,N_21351);
nor U23748 (N_23748,N_21370,N_21415);
or U23749 (N_23749,N_20355,N_21021);
nand U23750 (N_23750,N_21645,N_21037);
nor U23751 (N_23751,N_21001,N_20955);
or U23752 (N_23752,N_20551,N_21360);
xnor U23753 (N_23753,N_20014,N_20245);
nand U23754 (N_23754,N_20845,N_21429);
nor U23755 (N_23755,N_21955,N_21061);
nor U23756 (N_23756,N_20133,N_21864);
and U23757 (N_23757,N_21725,N_20023);
nor U23758 (N_23758,N_20522,N_21907);
nand U23759 (N_23759,N_20050,N_20544);
and U23760 (N_23760,N_20650,N_21099);
xor U23761 (N_23761,N_20433,N_20613);
or U23762 (N_23762,N_21149,N_20920);
or U23763 (N_23763,N_21105,N_21831);
nor U23764 (N_23764,N_21856,N_20635);
nor U23765 (N_23765,N_21408,N_21484);
or U23766 (N_23766,N_21852,N_20737);
and U23767 (N_23767,N_20411,N_21947);
and U23768 (N_23768,N_20997,N_20085);
and U23769 (N_23769,N_20920,N_20414);
or U23770 (N_23770,N_21717,N_20454);
nor U23771 (N_23771,N_21153,N_21484);
nand U23772 (N_23772,N_21094,N_20125);
xnor U23773 (N_23773,N_20247,N_20202);
or U23774 (N_23774,N_21316,N_20392);
nor U23775 (N_23775,N_20002,N_21608);
and U23776 (N_23776,N_20909,N_20203);
xor U23777 (N_23777,N_20103,N_21237);
or U23778 (N_23778,N_20453,N_21447);
xnor U23779 (N_23779,N_21573,N_20116);
and U23780 (N_23780,N_21182,N_20080);
or U23781 (N_23781,N_21032,N_21171);
nand U23782 (N_23782,N_21460,N_20219);
nor U23783 (N_23783,N_21331,N_20426);
xor U23784 (N_23784,N_21991,N_20400);
xor U23785 (N_23785,N_20655,N_21223);
nand U23786 (N_23786,N_21515,N_20565);
or U23787 (N_23787,N_21183,N_20615);
nand U23788 (N_23788,N_20201,N_20671);
nand U23789 (N_23789,N_20728,N_20627);
nor U23790 (N_23790,N_20662,N_20774);
nand U23791 (N_23791,N_21850,N_20549);
and U23792 (N_23792,N_20208,N_20193);
nand U23793 (N_23793,N_21451,N_21428);
nand U23794 (N_23794,N_21629,N_20774);
or U23795 (N_23795,N_20858,N_20621);
or U23796 (N_23796,N_20432,N_21306);
nor U23797 (N_23797,N_21977,N_20599);
xor U23798 (N_23798,N_20001,N_21256);
and U23799 (N_23799,N_21660,N_20637);
xor U23800 (N_23800,N_20099,N_20285);
nand U23801 (N_23801,N_20771,N_20424);
nor U23802 (N_23802,N_21651,N_21824);
and U23803 (N_23803,N_20777,N_20876);
or U23804 (N_23804,N_21528,N_20495);
and U23805 (N_23805,N_21958,N_20156);
xnor U23806 (N_23806,N_20692,N_20771);
or U23807 (N_23807,N_21826,N_20311);
and U23808 (N_23808,N_21609,N_21668);
nand U23809 (N_23809,N_21610,N_20220);
nand U23810 (N_23810,N_21883,N_21024);
and U23811 (N_23811,N_21906,N_20577);
and U23812 (N_23812,N_20393,N_20382);
nand U23813 (N_23813,N_20265,N_21331);
or U23814 (N_23814,N_20279,N_20564);
nand U23815 (N_23815,N_20348,N_20197);
and U23816 (N_23816,N_20729,N_21814);
xor U23817 (N_23817,N_21855,N_21482);
xnor U23818 (N_23818,N_21461,N_20145);
xnor U23819 (N_23819,N_20539,N_21572);
nand U23820 (N_23820,N_20379,N_20881);
or U23821 (N_23821,N_20469,N_20272);
xnor U23822 (N_23822,N_20375,N_21955);
nor U23823 (N_23823,N_20990,N_20231);
xor U23824 (N_23824,N_21997,N_21982);
and U23825 (N_23825,N_21102,N_21195);
nor U23826 (N_23826,N_20399,N_20702);
or U23827 (N_23827,N_20737,N_20606);
or U23828 (N_23828,N_20934,N_21630);
nand U23829 (N_23829,N_20332,N_20535);
nor U23830 (N_23830,N_21479,N_21260);
and U23831 (N_23831,N_21411,N_21179);
nand U23832 (N_23832,N_20843,N_21154);
nor U23833 (N_23833,N_21371,N_20049);
nor U23834 (N_23834,N_20272,N_20967);
or U23835 (N_23835,N_21016,N_20067);
or U23836 (N_23836,N_21096,N_21626);
and U23837 (N_23837,N_20395,N_21315);
or U23838 (N_23838,N_21912,N_21937);
or U23839 (N_23839,N_21650,N_21112);
nand U23840 (N_23840,N_20612,N_21356);
and U23841 (N_23841,N_20019,N_20437);
nand U23842 (N_23842,N_21114,N_21903);
nor U23843 (N_23843,N_20892,N_21831);
and U23844 (N_23844,N_21892,N_21468);
nand U23845 (N_23845,N_21393,N_20329);
and U23846 (N_23846,N_21028,N_21509);
and U23847 (N_23847,N_21217,N_20236);
and U23848 (N_23848,N_21495,N_20744);
nor U23849 (N_23849,N_21732,N_20577);
nor U23850 (N_23850,N_21130,N_20218);
xor U23851 (N_23851,N_20768,N_20597);
nor U23852 (N_23852,N_21616,N_21651);
and U23853 (N_23853,N_21232,N_21174);
and U23854 (N_23854,N_20228,N_21954);
xnor U23855 (N_23855,N_20920,N_20215);
nor U23856 (N_23856,N_20027,N_20966);
nor U23857 (N_23857,N_20554,N_21048);
nand U23858 (N_23858,N_20965,N_21245);
xnor U23859 (N_23859,N_20121,N_21405);
xor U23860 (N_23860,N_20174,N_20111);
or U23861 (N_23861,N_20112,N_20875);
and U23862 (N_23862,N_21853,N_20221);
nand U23863 (N_23863,N_20944,N_21909);
and U23864 (N_23864,N_21000,N_20862);
xor U23865 (N_23865,N_20772,N_21830);
or U23866 (N_23866,N_20351,N_20266);
and U23867 (N_23867,N_21230,N_21801);
xor U23868 (N_23868,N_21903,N_20195);
nor U23869 (N_23869,N_21975,N_20795);
and U23870 (N_23870,N_21934,N_20824);
nand U23871 (N_23871,N_21845,N_20282);
nand U23872 (N_23872,N_21176,N_21605);
nand U23873 (N_23873,N_21419,N_20946);
or U23874 (N_23874,N_21056,N_21603);
xnor U23875 (N_23875,N_20730,N_21187);
or U23876 (N_23876,N_21723,N_21492);
nor U23877 (N_23877,N_21253,N_21550);
nor U23878 (N_23878,N_21889,N_21826);
nor U23879 (N_23879,N_20781,N_21339);
nand U23880 (N_23880,N_21488,N_20203);
or U23881 (N_23881,N_20138,N_20785);
xnor U23882 (N_23882,N_20439,N_21141);
and U23883 (N_23883,N_21817,N_20953);
nand U23884 (N_23884,N_20998,N_21242);
and U23885 (N_23885,N_20170,N_21701);
nor U23886 (N_23886,N_21943,N_20397);
or U23887 (N_23887,N_21054,N_20690);
and U23888 (N_23888,N_20362,N_21517);
nor U23889 (N_23889,N_21256,N_20924);
nor U23890 (N_23890,N_20349,N_21579);
nor U23891 (N_23891,N_20548,N_20033);
and U23892 (N_23892,N_20084,N_21655);
or U23893 (N_23893,N_20903,N_21526);
nand U23894 (N_23894,N_21990,N_21196);
nor U23895 (N_23895,N_20075,N_21148);
or U23896 (N_23896,N_21994,N_20048);
xnor U23897 (N_23897,N_20972,N_21450);
xnor U23898 (N_23898,N_21630,N_20208);
xnor U23899 (N_23899,N_21430,N_20492);
and U23900 (N_23900,N_21636,N_21286);
xnor U23901 (N_23901,N_21488,N_21997);
nand U23902 (N_23902,N_20658,N_20577);
or U23903 (N_23903,N_20386,N_21526);
nand U23904 (N_23904,N_21541,N_20081);
nor U23905 (N_23905,N_20448,N_21977);
and U23906 (N_23906,N_20769,N_20334);
nand U23907 (N_23907,N_21524,N_21306);
nor U23908 (N_23908,N_20938,N_21206);
xnor U23909 (N_23909,N_21488,N_21224);
nor U23910 (N_23910,N_20033,N_21777);
xnor U23911 (N_23911,N_20203,N_20307);
nor U23912 (N_23912,N_20842,N_21894);
nor U23913 (N_23913,N_21447,N_21485);
xor U23914 (N_23914,N_20991,N_20951);
xnor U23915 (N_23915,N_20228,N_20728);
or U23916 (N_23916,N_21736,N_21916);
nor U23917 (N_23917,N_20254,N_20877);
nor U23918 (N_23918,N_21736,N_20762);
nor U23919 (N_23919,N_20882,N_21975);
xnor U23920 (N_23920,N_20564,N_20057);
and U23921 (N_23921,N_21111,N_21269);
nor U23922 (N_23922,N_20446,N_21729);
xor U23923 (N_23923,N_21222,N_20316);
nand U23924 (N_23924,N_21713,N_20398);
or U23925 (N_23925,N_21127,N_21052);
or U23926 (N_23926,N_21325,N_21186);
nor U23927 (N_23927,N_21784,N_20011);
nor U23928 (N_23928,N_20957,N_20252);
or U23929 (N_23929,N_20616,N_20230);
or U23930 (N_23930,N_20469,N_20219);
xnor U23931 (N_23931,N_21843,N_20676);
and U23932 (N_23932,N_20576,N_20322);
or U23933 (N_23933,N_20169,N_20058);
nand U23934 (N_23934,N_20177,N_20205);
xnor U23935 (N_23935,N_21257,N_20356);
and U23936 (N_23936,N_20029,N_21120);
nor U23937 (N_23937,N_20518,N_21341);
xnor U23938 (N_23938,N_20142,N_21601);
and U23939 (N_23939,N_20431,N_21780);
nand U23940 (N_23940,N_20013,N_20204);
and U23941 (N_23941,N_21781,N_21546);
or U23942 (N_23942,N_21619,N_20017);
and U23943 (N_23943,N_21809,N_21318);
nor U23944 (N_23944,N_20271,N_20188);
nor U23945 (N_23945,N_20089,N_20853);
or U23946 (N_23946,N_21454,N_20473);
or U23947 (N_23947,N_20268,N_20895);
or U23948 (N_23948,N_21175,N_20872);
xnor U23949 (N_23949,N_20355,N_20516);
nor U23950 (N_23950,N_21188,N_21435);
nor U23951 (N_23951,N_20866,N_20123);
or U23952 (N_23952,N_21217,N_21350);
and U23953 (N_23953,N_20889,N_21272);
nor U23954 (N_23954,N_20031,N_20076);
or U23955 (N_23955,N_20515,N_20882);
nand U23956 (N_23956,N_20805,N_20610);
and U23957 (N_23957,N_21753,N_20832);
and U23958 (N_23958,N_21536,N_20677);
nor U23959 (N_23959,N_20472,N_20727);
or U23960 (N_23960,N_21065,N_21618);
or U23961 (N_23961,N_20686,N_20108);
nor U23962 (N_23962,N_21458,N_21831);
and U23963 (N_23963,N_21386,N_21453);
nand U23964 (N_23964,N_20892,N_20026);
nor U23965 (N_23965,N_21805,N_20185);
or U23966 (N_23966,N_20642,N_21755);
xor U23967 (N_23967,N_20571,N_20429);
nand U23968 (N_23968,N_20076,N_21975);
nor U23969 (N_23969,N_20492,N_20269);
nand U23970 (N_23970,N_20124,N_20902);
or U23971 (N_23971,N_21163,N_20000);
or U23972 (N_23972,N_21476,N_21243);
or U23973 (N_23973,N_21332,N_21458);
nand U23974 (N_23974,N_20383,N_20877);
nand U23975 (N_23975,N_21083,N_20747);
or U23976 (N_23976,N_21579,N_20141);
or U23977 (N_23977,N_21514,N_20536);
nor U23978 (N_23978,N_21537,N_21393);
or U23979 (N_23979,N_20929,N_20221);
nand U23980 (N_23980,N_21793,N_21715);
and U23981 (N_23981,N_20510,N_20952);
and U23982 (N_23982,N_21978,N_21135);
nor U23983 (N_23983,N_20070,N_21904);
and U23984 (N_23984,N_21815,N_20200);
nor U23985 (N_23985,N_21374,N_21316);
nand U23986 (N_23986,N_21169,N_20685);
nor U23987 (N_23987,N_20494,N_21220);
or U23988 (N_23988,N_21487,N_21731);
and U23989 (N_23989,N_21746,N_20018);
and U23990 (N_23990,N_21669,N_20562);
and U23991 (N_23991,N_20157,N_21386);
xor U23992 (N_23992,N_21608,N_21616);
xnor U23993 (N_23993,N_20574,N_21250);
or U23994 (N_23994,N_21860,N_20863);
nand U23995 (N_23995,N_21806,N_21323);
nand U23996 (N_23996,N_20016,N_20681);
nor U23997 (N_23997,N_21508,N_20706);
or U23998 (N_23998,N_20827,N_20532);
or U23999 (N_23999,N_21308,N_21100);
xor U24000 (N_24000,N_23785,N_23742);
and U24001 (N_24001,N_23935,N_23452);
or U24002 (N_24002,N_22636,N_22379);
or U24003 (N_24003,N_23947,N_23889);
and U24004 (N_24004,N_23199,N_22580);
nand U24005 (N_24005,N_23324,N_23024);
nor U24006 (N_24006,N_22256,N_22598);
and U24007 (N_24007,N_23458,N_23266);
xnor U24008 (N_24008,N_22676,N_22761);
nand U24009 (N_24009,N_23915,N_23920);
xnor U24010 (N_24010,N_22563,N_23527);
nand U24011 (N_24011,N_23558,N_22036);
xnor U24012 (N_24012,N_23321,N_23862);
and U24013 (N_24013,N_23313,N_22618);
and U24014 (N_24014,N_23428,N_23007);
or U24015 (N_24015,N_23547,N_23532);
and U24016 (N_24016,N_23339,N_23178);
xor U24017 (N_24017,N_23934,N_23939);
or U24018 (N_24018,N_23474,N_22467);
xor U24019 (N_24019,N_22791,N_22503);
nand U24020 (N_24020,N_23437,N_23460);
or U24021 (N_24021,N_22799,N_23447);
or U24022 (N_24022,N_23867,N_22183);
nor U24023 (N_24023,N_23316,N_23948);
nor U24024 (N_24024,N_22737,N_23227);
xor U24025 (N_24025,N_23264,N_22307);
nand U24026 (N_24026,N_23223,N_22170);
and U24027 (N_24027,N_23820,N_23666);
and U24028 (N_24028,N_23743,N_23591);
or U24029 (N_24029,N_22728,N_23769);
and U24030 (N_24030,N_22508,N_23149);
nor U24031 (N_24031,N_22510,N_23026);
and U24032 (N_24032,N_22306,N_22238);
nor U24033 (N_24033,N_22884,N_22140);
nand U24034 (N_24034,N_23354,N_22518);
and U24035 (N_24035,N_22611,N_22829);
and U24036 (N_24036,N_22371,N_23563);
nor U24037 (N_24037,N_23086,N_22608);
and U24038 (N_24038,N_22020,N_23125);
or U24039 (N_24039,N_23749,N_23622);
nor U24040 (N_24040,N_23551,N_22187);
or U24041 (N_24041,N_22412,N_22346);
xor U24042 (N_24042,N_22076,N_22858);
or U24043 (N_24043,N_23176,N_22182);
nor U24044 (N_24044,N_23422,N_22871);
nand U24045 (N_24045,N_23260,N_22910);
nor U24046 (N_24046,N_22119,N_22311);
nand U24047 (N_24047,N_22203,N_22367);
nor U24048 (N_24048,N_22021,N_23728);
nor U24049 (N_24049,N_22493,N_23475);
and U24050 (N_24050,N_23393,N_22414);
nand U24051 (N_24051,N_23231,N_23943);
xnor U24052 (N_24052,N_23353,N_22305);
or U24053 (N_24053,N_22572,N_22186);
xnor U24054 (N_24054,N_22616,N_22952);
nor U24055 (N_24055,N_22396,N_22250);
or U24056 (N_24056,N_23689,N_23120);
and U24057 (N_24057,N_22835,N_23841);
xnor U24058 (N_24058,N_23850,N_22294);
xnor U24059 (N_24059,N_23955,N_23601);
nand U24060 (N_24060,N_23617,N_23959);
nand U24061 (N_24061,N_22716,N_22751);
or U24062 (N_24062,N_22524,N_22339);
nand U24063 (N_24063,N_22115,N_22504);
xnor U24064 (N_24064,N_22885,N_23992);
nand U24065 (N_24065,N_23792,N_22255);
and U24066 (N_24066,N_23216,N_23465);
and U24067 (N_24067,N_22805,N_22803);
xor U24068 (N_24068,N_23006,N_23750);
nor U24069 (N_24069,N_23982,N_23213);
or U24070 (N_24070,N_23800,N_23188);
nand U24071 (N_24071,N_23413,N_23357);
or U24072 (N_24072,N_22681,N_22543);
nand U24073 (N_24073,N_23745,N_22513);
xnor U24074 (N_24074,N_22351,N_22141);
nor U24075 (N_24075,N_22784,N_23654);
nor U24076 (N_24076,N_22614,N_23277);
and U24077 (N_24077,N_23259,N_22623);
xor U24078 (N_24078,N_23294,N_22825);
nor U24079 (N_24079,N_22559,N_22961);
nor U24080 (N_24080,N_22837,N_22477);
and U24081 (N_24081,N_23767,N_23166);
or U24082 (N_24082,N_22804,N_22642);
xnor U24083 (N_24083,N_22533,N_22487);
nand U24084 (N_24084,N_23197,N_22447);
nor U24085 (N_24085,N_22499,N_23950);
nor U24086 (N_24086,N_23423,N_22318);
xnor U24087 (N_24087,N_23190,N_23506);
nand U24088 (N_24088,N_23242,N_23013);
and U24089 (N_24089,N_22286,N_23416);
nor U24090 (N_24090,N_22735,N_23234);
and U24091 (N_24091,N_23185,N_22989);
nand U24092 (N_24092,N_22770,N_23191);
and U24093 (N_24093,N_23719,N_23675);
xnor U24094 (N_24094,N_23008,N_23297);
and U24095 (N_24095,N_23840,N_22029);
nor U24096 (N_24096,N_23420,N_23431);
xor U24097 (N_24097,N_23633,N_23479);
and U24098 (N_24098,N_22104,N_22857);
or U24099 (N_24099,N_23523,N_23516);
xnor U24100 (N_24100,N_22360,N_23442);
xnor U24101 (N_24101,N_23912,N_23187);
and U24102 (N_24102,N_22356,N_22413);
or U24103 (N_24103,N_23363,N_22683);
or U24104 (N_24104,N_23502,N_23031);
nand U24105 (N_24105,N_22887,N_23146);
nor U24106 (N_24106,N_23459,N_22970);
nand U24107 (N_24107,N_23916,N_22401);
xnor U24108 (N_24108,N_23898,N_22303);
nand U24109 (N_24109,N_23468,N_23969);
nor U24110 (N_24110,N_22004,N_22529);
or U24111 (N_24111,N_22423,N_22484);
and U24112 (N_24112,N_22842,N_22832);
and U24113 (N_24113,N_23366,N_22122);
or U24114 (N_24114,N_23695,N_22348);
nor U24115 (N_24115,N_22913,N_22922);
or U24116 (N_24116,N_22968,N_23441);
xor U24117 (N_24117,N_23782,N_23524);
nor U24118 (N_24118,N_23195,N_23741);
or U24119 (N_24119,N_23789,N_22344);
or U24120 (N_24120,N_22750,N_22295);
xnor U24121 (N_24121,N_22710,N_23685);
nand U24122 (N_24122,N_22098,N_22424);
xnor U24123 (N_24123,N_23609,N_22908);
xor U24124 (N_24124,N_22596,N_22852);
and U24125 (N_24125,N_23011,N_22662);
nand U24126 (N_24126,N_23057,N_22117);
xnor U24127 (N_24127,N_22497,N_23905);
nor U24128 (N_24128,N_22022,N_22181);
nand U24129 (N_24129,N_23847,N_23001);
xnor U24130 (N_24130,N_23148,N_23257);
xnor U24131 (N_24131,N_23530,N_23069);
and U24132 (N_24132,N_23746,N_22382);
or U24133 (N_24133,N_23074,N_22925);
and U24134 (N_24134,N_22836,N_22519);
xor U24135 (N_24135,N_22395,N_22840);
and U24136 (N_24136,N_22815,N_22127);
or U24137 (N_24137,N_22979,N_22478);
nand U24138 (N_24138,N_22025,N_23845);
nor U24139 (N_24139,N_22560,N_22156);
and U24140 (N_24140,N_22998,N_22262);
nand U24141 (N_24141,N_23127,N_22700);
and U24142 (N_24142,N_23981,N_23499);
nor U24143 (N_24143,N_23846,N_23970);
or U24144 (N_24144,N_22648,N_22637);
nor U24145 (N_24145,N_22350,N_22381);
xnor U24146 (N_24146,N_22934,N_22860);
nor U24147 (N_24147,N_22765,N_23508);
nand U24148 (N_24148,N_22530,N_22121);
nand U24149 (N_24149,N_23207,N_23583);
nor U24150 (N_24150,N_23809,N_22577);
or U24151 (N_24151,N_22668,N_23937);
or U24152 (N_24152,N_22509,N_23710);
or U24153 (N_24153,N_23173,N_22341);
or U24154 (N_24154,N_22912,N_22292);
xor U24155 (N_24155,N_22599,N_23725);
nor U24156 (N_24156,N_22253,N_23070);
nand U24157 (N_24157,N_23993,N_23112);
nor U24158 (N_24158,N_23483,N_22366);
or U24159 (N_24159,N_23359,N_22859);
xor U24160 (N_24160,N_23559,N_22853);
xnor U24161 (N_24161,N_22139,N_22012);
and U24162 (N_24162,N_22595,N_23117);
nand U24163 (N_24163,N_22663,N_23880);
xor U24164 (N_24164,N_23630,N_23844);
or U24165 (N_24165,N_22528,N_22643);
nor U24166 (N_24166,N_22236,N_22847);
or U24167 (N_24167,N_22212,N_23635);
nand U24168 (N_24168,N_23106,N_22581);
xor U24169 (N_24169,N_22031,N_23881);
nand U24170 (N_24170,N_22694,N_22748);
or U24171 (N_24171,N_22387,N_23812);
and U24172 (N_24172,N_23778,N_23930);
xnor U24173 (N_24173,N_23625,N_23752);
nor U24174 (N_24174,N_23080,N_23453);
and U24175 (N_24175,N_22613,N_22445);
or U24176 (N_24176,N_22196,N_23748);
and U24177 (N_24177,N_23519,N_23537);
and U24178 (N_24178,N_23803,N_22277);
and U24179 (N_24179,N_22715,N_23744);
and U24180 (N_24180,N_22450,N_23376);
or U24181 (N_24181,N_22045,N_22909);
nor U24182 (N_24182,N_22352,N_22856);
and U24183 (N_24183,N_22693,N_23075);
or U24184 (N_24184,N_22354,N_23713);
and U24185 (N_24185,N_22762,N_22438);
nor U24186 (N_24186,N_22105,N_23957);
or U24187 (N_24187,N_23214,N_23571);
xor U24188 (N_24188,N_23680,N_22574);
xnor U24189 (N_24189,N_22875,N_23588);
xnor U24190 (N_24190,N_23758,N_23281);
xor U24191 (N_24191,N_22023,N_22435);
nand U24192 (N_24192,N_22687,N_23462);
nand U24193 (N_24193,N_23342,N_22824);
or U24194 (N_24194,N_22557,N_22327);
nand U24195 (N_24195,N_23068,N_23918);
or U24196 (N_24196,N_22271,N_23320);
nand U24197 (N_24197,N_23640,N_23333);
or U24198 (N_24198,N_22163,N_23379);
nand U24199 (N_24199,N_23501,N_23433);
or U24200 (N_24200,N_22848,N_22289);
nor U24201 (N_24201,N_23550,N_23585);
xor U24202 (N_24202,N_22850,N_22521);
xor U24203 (N_24203,N_23830,N_22464);
xor U24204 (N_24204,N_22343,N_23271);
nor U24205 (N_24205,N_22434,N_23407);
nor U24206 (N_24206,N_23664,N_23842);
nor U24207 (N_24207,N_22627,N_23765);
and U24208 (N_24208,N_22915,N_23102);
and U24209 (N_24209,N_22874,N_22601);
nor U24210 (N_24210,N_23819,N_23312);
or U24211 (N_24211,N_22746,N_23626);
and U24212 (N_24212,N_23810,N_23595);
nand U24213 (N_24213,N_22780,N_22778);
xor U24214 (N_24214,N_23738,N_23619);
and U24215 (N_24215,N_22077,N_23647);
nor U24216 (N_24216,N_22674,N_22368);
and U24217 (N_24217,N_23072,N_23562);
nand U24218 (N_24218,N_23050,N_22633);
nand U24219 (N_24219,N_22759,N_22719);
nand U24220 (N_24220,N_23720,N_22554);
nand U24221 (N_24221,N_22777,N_22834);
nor U24222 (N_24222,N_23557,N_23781);
or U24223 (N_24223,N_22034,N_22767);
or U24224 (N_24224,N_23855,N_23065);
and U24225 (N_24225,N_23799,N_22763);
nor U24226 (N_24226,N_22193,N_22906);
nand U24227 (N_24227,N_22245,N_23470);
xor U24228 (N_24228,N_23087,N_23497);
xnor U24229 (N_24229,N_22612,N_22609);
and U24230 (N_24230,N_23764,N_23409);
nor U24231 (N_24231,N_22669,N_22891);
nand U24232 (N_24232,N_23730,N_22749);
and U24233 (N_24233,N_23747,N_22760);
nor U24234 (N_24234,N_22461,N_22699);
nand U24235 (N_24235,N_22514,N_23651);
nor U24236 (N_24236,N_22280,N_23184);
nor U24237 (N_24237,N_23674,N_22455);
and U24238 (N_24238,N_23410,N_22702);
nor U24239 (N_24239,N_23139,N_22332);
nor U24240 (N_24240,N_22657,N_22112);
nor U24241 (N_24241,N_22326,N_23568);
and U24242 (N_24242,N_22526,N_23427);
nand U24243 (N_24243,N_23477,N_22442);
nand U24244 (N_24244,N_22838,N_23894);
nor U24245 (N_24245,N_23882,N_23079);
nand U24246 (N_24246,N_23295,N_22392);
or U24247 (N_24247,N_22130,N_23945);
nand U24248 (N_24248,N_23384,N_23977);
nor U24249 (N_24249,N_23949,N_22254);
or U24250 (N_24250,N_23656,N_23122);
xnor U24251 (N_24251,N_23099,N_22177);
nand U24252 (N_24252,N_22083,N_22325);
xor U24253 (N_24253,N_22172,N_22708);
nor U24254 (N_24254,N_23902,N_22224);
and U24255 (N_24255,N_22606,N_23404);
and U24256 (N_24256,N_23472,N_23552);
nor U24257 (N_24257,N_22607,N_23715);
nor U24258 (N_24258,N_23017,N_22818);
nor U24259 (N_24259,N_22188,N_22391);
and U24260 (N_24260,N_22474,N_23192);
or U24261 (N_24261,N_23703,N_23440);
nand U24262 (N_24262,N_23267,N_23135);
and U24263 (N_24263,N_23972,N_22027);
or U24264 (N_24264,N_23144,N_22243);
nor U24265 (N_24265,N_22417,N_23953);
nor U24266 (N_24266,N_22788,N_23283);
and U24267 (N_24267,N_22864,N_23340);
xor U24268 (N_24268,N_23700,N_22877);
nor U24269 (N_24269,N_22619,N_22285);
xnor U24270 (N_24270,N_22397,N_22429);
nor U24271 (N_24271,N_23999,N_22666);
and U24272 (N_24272,N_22895,N_22373);
and U24273 (N_24273,N_22407,N_22394);
and U24274 (N_24274,N_23940,N_23158);
and U24275 (N_24275,N_23167,N_22399);
xnor U24276 (N_24276,N_23318,N_22667);
nand U24277 (N_24277,N_23131,N_22334);
nor U24278 (N_24278,N_23151,N_23244);
or U24279 (N_24279,N_22873,N_23729);
and U24280 (N_24280,N_23150,N_23771);
nand U24281 (N_24281,N_22492,N_23761);
nor U24282 (N_24282,N_23291,N_22201);
nand U24283 (N_24283,N_22209,N_22592);
xor U24284 (N_24284,N_22812,N_23786);
nand U24285 (N_24285,N_22135,N_22570);
nand U24286 (N_24286,N_22386,N_23143);
and U24287 (N_24287,N_22491,N_22960);
nand U24288 (N_24288,N_23642,N_23589);
or U24289 (N_24289,N_22195,N_22422);
or U24290 (N_24290,N_22428,N_23966);
nor U24291 (N_24291,N_22248,N_22703);
and U24292 (N_24292,N_23067,N_23757);
xnor U24293 (N_24293,N_23309,N_23186);
nor U24294 (N_24294,N_23274,N_22276);
nand U24295 (N_24295,N_23218,N_23514);
and U24296 (N_24296,N_23066,N_23751);
or U24297 (N_24297,N_22591,N_23358);
xnor U24298 (N_24298,N_22639,N_22260);
or U24299 (N_24299,N_23119,N_22535);
nor U24300 (N_24300,N_22846,N_23372);
nor U24301 (N_24301,N_23023,N_22030);
or U24302 (N_24302,N_22481,N_23027);
and U24303 (N_24303,N_23206,N_22174);
and U24304 (N_24304,N_23263,N_22880);
nand U24305 (N_24305,N_22907,N_23138);
and U24306 (N_24306,N_23314,N_23702);
and U24307 (N_24307,N_23322,N_22109);
nor U24308 (N_24308,N_22655,N_22349);
and U24309 (N_24309,N_23852,N_22009);
xor U24310 (N_24310,N_22890,N_23991);
nor U24311 (N_24311,N_23181,N_23913);
and U24312 (N_24312,N_23798,N_23971);
xor U24313 (N_24313,N_22977,N_23145);
nand U24314 (N_24314,N_23606,N_23451);
nand U24315 (N_24315,N_22126,N_23289);
nor U24316 (N_24316,N_22019,N_22107);
nor U24317 (N_24317,N_23003,N_22615);
nand U24318 (N_24318,N_22309,N_22830);
nand U24319 (N_24319,N_23539,N_22975);
xnor U24320 (N_24320,N_23543,N_23432);
xnor U24321 (N_24321,N_23317,N_23860);
xor U24322 (N_24322,N_23929,N_23247);
xor U24323 (N_24323,N_23018,N_22133);
nor U24324 (N_24324,N_23927,N_22649);
or U24325 (N_24325,N_23723,N_22073);
nor U24326 (N_24326,N_22789,N_22820);
xnor U24327 (N_24327,N_23893,N_22766);
xor U24328 (N_24328,N_23476,N_22957);
nand U24329 (N_24329,N_23641,N_23323);
and U24330 (N_24330,N_22816,N_22000);
and U24331 (N_24331,N_23132,N_22550);
xor U24332 (N_24332,N_23446,N_23667);
or U24333 (N_24333,N_22995,N_22866);
nor U24334 (N_24334,N_23964,N_22734);
nand U24335 (N_24335,N_23096,N_23212);
or U24336 (N_24336,N_23693,N_23136);
nand U24337 (N_24337,N_22670,N_23464);
and U24338 (N_24338,N_22604,N_23296);
nand U24339 (N_24339,N_23444,N_22774);
or U24340 (N_24340,N_23859,N_23019);
nand U24341 (N_24341,N_22056,N_23368);
nand U24342 (N_24342,N_23574,N_23361);
xnor U24343 (N_24343,N_23076,N_22929);
or U24344 (N_24344,N_22390,N_22498);
nor U24345 (N_24345,N_22963,N_22568);
or U24346 (N_24346,N_23756,N_23721);
nor U24347 (N_24347,N_22213,N_22164);
nand U24348 (N_24348,N_22831,N_22179);
nand U24349 (N_24349,N_23512,N_22316);
nand U24350 (N_24350,N_23224,N_22720);
and U24351 (N_24351,N_22582,N_22567);
nor U24352 (N_24352,N_23718,N_23620);
nor U24353 (N_24353,N_22240,N_23034);
nand U24354 (N_24354,N_23285,N_22002);
nor U24355 (N_24355,N_22380,N_23327);
or U24356 (N_24356,N_22257,N_23804);
nand U24357 (N_24357,N_22549,N_23010);
or U24358 (N_24358,N_22152,N_22166);
xor U24359 (N_24359,N_23240,N_22071);
nand U24360 (N_24360,N_23660,N_22544);
or U24361 (N_24361,N_23770,N_22333);
and U24362 (N_24362,N_22267,N_22771);
and U24363 (N_24363,N_22755,N_23485);
or U24364 (N_24364,N_23225,N_22132);
nor U24365 (N_24365,N_23994,N_22764);
or U24366 (N_24366,N_22093,N_22270);
and U24367 (N_24367,N_23042,N_23596);
nand U24368 (N_24368,N_23374,N_22185);
nor U24369 (N_24369,N_23838,N_22947);
or U24370 (N_24370,N_23403,N_22261);
or U24371 (N_24371,N_23717,N_22610);
or U24372 (N_24372,N_23863,N_23033);
nand U24373 (N_24373,N_23534,N_22843);
nor U24374 (N_24374,N_23137,N_23036);
nor U24375 (N_24375,N_22078,N_22990);
and U24376 (N_24376,N_22787,N_22473);
or U24377 (N_24377,N_22718,N_22103);
and U24378 (N_24378,N_22226,N_22219);
nor U24379 (N_24379,N_23714,N_23597);
nor U24380 (N_24380,N_22108,N_22042);
nand U24381 (N_24381,N_22128,N_22015);
nand U24382 (N_24382,N_23973,N_23396);
nand U24383 (N_24383,N_22851,N_22650);
nor U24384 (N_24384,N_23513,N_23293);
or U24385 (N_24385,N_22129,N_22779);
and U24386 (N_24386,N_22018,N_23967);
nor U24387 (N_24387,N_23021,N_22299);
and U24388 (N_24388,N_22551,N_22040);
nor U24389 (N_24389,N_23627,N_23215);
xor U24390 (N_24390,N_22232,N_23044);
or U24391 (N_24391,N_23375,N_22279);
nand U24392 (N_24392,N_22652,N_23835);
and U24393 (N_24393,N_23888,N_23351);
xnor U24394 (N_24394,N_23579,N_23473);
and U24395 (N_24395,N_23343,N_22897);
nand U24396 (N_24396,N_23790,N_23794);
nor U24397 (N_24397,N_23836,N_23286);
or U24398 (N_24398,N_22819,N_22208);
nor U24399 (N_24399,N_23592,N_23997);
nor U24400 (N_24400,N_22684,N_22426);
or U24401 (N_24401,N_23854,N_22162);
nand U24402 (N_24402,N_22051,N_23892);
nor U24403 (N_24403,N_22336,N_22849);
nand U24404 (N_24404,N_23503,N_22060);
nor U24405 (N_24405,N_23832,N_22597);
nor U24406 (N_24406,N_22986,N_23088);
nand U24407 (N_24407,N_23634,N_23153);
nor U24408 (N_24408,N_22796,N_22939);
nand U24409 (N_24409,N_23039,N_23435);
nand U24410 (N_24410,N_22211,N_22446);
xor U24411 (N_24411,N_22867,N_22403);
xor U24412 (N_24412,N_22100,N_22006);
and U24413 (N_24413,N_23663,N_23616);
or U24414 (N_24414,N_23933,N_22587);
and U24415 (N_24415,N_23163,N_23690);
nand U24416 (N_24416,N_23275,N_23356);
nand U24417 (N_24417,N_23914,N_22089);
or U24418 (N_24418,N_22793,N_22338);
nand U24419 (N_24419,N_22756,N_23009);
nor U24420 (N_24420,N_23910,N_23335);
and U24421 (N_24421,N_23208,N_22502);
nor U24422 (N_24422,N_22335,N_23142);
nor U24423 (N_24423,N_22010,N_23360);
nor U24424 (N_24424,N_23670,N_22297);
nand U24425 (N_24425,N_22096,N_23676);
xnor U24426 (N_24426,N_22808,N_23114);
xnor U24427 (N_24427,N_22246,N_22082);
or U24428 (N_24428,N_23491,N_22290);
xnor U24429 (N_24429,N_23907,N_23268);
and U24430 (N_24430,N_23421,N_23716);
and U24431 (N_24431,N_22039,N_23974);
xor U24432 (N_24432,N_23531,N_23678);
and U24433 (N_24433,N_23418,N_23600);
xor U24434 (N_24434,N_23529,N_22944);
and U24435 (N_24435,N_23254,N_22026);
and U24436 (N_24436,N_23346,N_23487);
nand U24437 (N_24437,N_23874,N_23813);
nor U24438 (N_24438,N_22106,N_23107);
xnor U24439 (N_24439,N_22889,N_22966);
or U24440 (N_24440,N_22199,N_23201);
xnor U24441 (N_24441,N_22085,N_23498);
and U24442 (N_24442,N_23347,N_22994);
xor U24443 (N_24443,N_22449,N_22090);
and U24444 (N_24444,N_23928,N_23671);
nor U24445 (N_24445,N_22754,N_23038);
and U24446 (N_24446,N_23696,N_22483);
xor U24447 (N_24447,N_22558,N_23900);
nor U24448 (N_24448,N_23390,N_22631);
nor U24449 (N_24449,N_22638,N_22151);
or U24450 (N_24450,N_22878,N_23657);
xnor U24451 (N_24451,N_22538,N_23652);
xnor U24452 (N_24452,N_23814,N_23662);
xnor U24453 (N_24453,N_23326,N_22137);
xnor U24454 (N_24454,N_22190,N_23791);
xor U24455 (N_24455,N_22724,N_23015);
xnor U24456 (N_24456,N_22237,N_22537);
nor U24457 (N_24457,N_23046,N_23304);
nor U24458 (N_24458,N_23113,N_22712);
nand U24459 (N_24459,N_22458,N_22173);
xor U24460 (N_24460,N_23486,N_22893);
nand U24461 (N_24461,N_22987,N_22923);
nand U24462 (N_24462,N_22008,N_22532);
and U24463 (N_24463,N_22328,N_23364);
xnor U24464 (N_24464,N_22041,N_23480);
xor U24465 (N_24465,N_23735,N_22941);
nor U24466 (N_24466,N_22782,N_23397);
xnor U24467 (N_24467,N_22244,N_23891);
or U24468 (N_24468,N_22383,N_23989);
nand U24469 (N_24469,N_22340,N_23707);
or U24470 (N_24470,N_22204,N_22772);
xnor U24471 (N_24471,N_23946,N_23202);
xor U24472 (N_24472,N_23580,N_22634);
nand U24473 (N_24473,N_23545,N_23164);
and U24474 (N_24474,N_23668,N_23536);
and U24475 (N_24475,N_23909,N_22753);
xor U24476 (N_24476,N_23560,N_22953);
nand U24477 (N_24477,N_22679,N_23586);
and U24478 (N_24478,N_22622,N_23236);
or U24479 (N_24479,N_23084,N_22659);
nand U24480 (N_24480,N_22523,N_23526);
xnor U24481 (N_24481,N_23613,N_22485);
nand U24482 (N_24482,N_22672,N_22827);
nor U24483 (N_24483,N_22274,N_23637);
xor U24484 (N_24484,N_23241,N_23848);
and U24485 (N_24485,N_23706,N_22826);
nor U24486 (N_24486,N_23694,N_23533);
xor U24487 (N_24487,N_22635,N_23302);
nor U24488 (N_24488,N_23521,N_23279);
or U24489 (N_24489,N_23439,N_22628);
xor U24490 (N_24490,N_23724,N_23684);
or U24491 (N_24491,N_23762,N_22223);
and U24492 (N_24492,N_22421,N_23699);
nor U24493 (N_24493,N_23976,N_22564);
and U24494 (N_24494,N_22926,N_23448);
nor U24495 (N_24495,N_23051,N_23352);
and U24496 (N_24496,N_23865,N_23869);
nand U24497 (N_24497,N_22677,N_22653);
or U24498 (N_24498,N_23053,N_22575);
xor U24499 (N_24499,N_23002,N_23180);
xor U24500 (N_24500,N_22522,N_23573);
or U24501 (N_24501,N_23825,N_23331);
and U24502 (N_24502,N_22411,N_22807);
nor U24503 (N_24503,N_22822,N_23570);
or U24504 (N_24504,N_23398,N_23525);
and U24505 (N_24505,N_22512,N_23116);
nand U24506 (N_24506,N_23329,N_23030);
or U24507 (N_24507,N_23556,N_22589);
xnor U24508 (N_24508,N_23064,N_23877);
nor U24509 (N_24509,N_23917,N_22374);
nor U24510 (N_24510,N_22415,N_23430);
nor U24511 (N_24511,N_23436,N_23906);
and U24512 (N_24512,N_22942,N_23055);
xor U24513 (N_24513,N_23885,N_22490);
and U24514 (N_24514,N_23091,N_23170);
and U24515 (N_24515,N_22323,N_22016);
nand U24516 (N_24516,N_23179,N_22283);
nand U24517 (N_24517,N_23338,N_23124);
nand U24518 (N_24518,N_22313,N_23219);
nor U24519 (N_24519,N_22259,N_22661);
nor U24520 (N_24520,N_22745,N_22969);
and U24521 (N_24521,N_22099,N_22281);
nor U24522 (N_24522,N_22817,N_23155);
and U24523 (N_24523,N_22408,N_22888);
and U24524 (N_24524,N_23371,N_22301);
and U24525 (N_24525,N_23837,N_22839);
xnor U24526 (N_24526,N_22420,N_23824);
xnor U24527 (N_24527,N_22911,N_23577);
xnor U24528 (N_24528,N_22233,N_22378);
xor U24529 (N_24529,N_22542,N_22854);
xnor U24530 (N_24530,N_22741,N_23779);
nand U24531 (N_24531,N_23542,N_22116);
and U24532 (N_24532,N_22123,N_22917);
nor U24533 (N_24533,N_23990,N_22752);
xor U24534 (N_24534,N_23203,N_22217);
and U24535 (N_24535,N_23105,N_23061);
or U24536 (N_24536,N_22235,N_23092);
and U24537 (N_24537,N_23232,N_22358);
and U24538 (N_24538,N_23141,N_22014);
or U24539 (N_24539,N_23020,N_23211);
or U24540 (N_24540,N_22673,N_22409);
and U24541 (N_24541,N_23337,N_22959);
nor U24542 (N_24542,N_22302,N_23424);
nor U24543 (N_24543,N_23901,N_22017);
or U24544 (N_24544,N_23054,N_23755);
nand U24545 (N_24545,N_22158,N_22087);
nor U24546 (N_24546,N_23063,N_23461);
nor U24547 (N_24547,N_23209,N_22656);
or U24548 (N_24548,N_23012,N_22184);
nor U24549 (N_24549,N_23029,N_22239);
nor U24550 (N_24550,N_22978,N_23833);
nand U24551 (N_24551,N_22928,N_23237);
nor U24552 (N_24552,N_23123,N_23478);
or U24553 (N_24553,N_22320,N_22932);
or U24554 (N_24554,N_22377,N_23658);
nor U24555 (N_24555,N_22419,N_23768);
nor U24556 (N_24556,N_22962,N_22050);
nor U24557 (N_24557,N_23307,N_23248);
xor U24558 (N_24558,N_23911,N_23932);
nand U24559 (N_24559,N_23490,N_23697);
or U24560 (N_24560,N_23687,N_22427);
xnor U24561 (N_24561,N_22971,N_23639);
xnor U24562 (N_24562,N_23886,N_23849);
nand U24563 (N_24563,N_22479,N_23968);
xnor U24564 (N_24564,N_22322,N_23871);
xor U24565 (N_24565,N_22058,N_22388);
xor U24566 (N_24566,N_22949,N_22937);
and U24567 (N_24567,N_23336,N_23594);
or U24568 (N_24568,N_23417,N_23344);
nor U24569 (N_24569,N_23082,N_23306);
nand U24570 (N_24570,N_23367,N_23636);
nor U24571 (N_24571,N_22101,N_22258);
and U24572 (N_24572,N_22697,N_22293);
xor U24573 (N_24573,N_23382,N_23960);
nand U24574 (N_24574,N_23400,N_23156);
or U24575 (N_24575,N_23045,N_22583);
nor U24576 (N_24576,N_23505,N_23772);
or U24577 (N_24577,N_23827,N_22319);
nor U24578 (N_24578,N_23466,N_22918);
or U24579 (N_24579,N_22773,N_22561);
xor U24580 (N_24580,N_22973,N_22393);
and U24581 (N_24581,N_23040,N_22471);
nor U24582 (N_24582,N_22153,N_22324);
xor U24583 (N_24583,N_23310,N_23904);
nor U24584 (N_24584,N_23249,N_23884);
nand U24585 (N_24585,N_23807,N_23806);
and U24586 (N_24586,N_22363,N_22505);
xor U24587 (N_24587,N_22221,N_22171);
nor U24588 (N_24588,N_22097,N_23041);
and U24589 (N_24589,N_23683,N_22730);
or U24590 (N_24590,N_23873,N_23655);
and U24591 (N_24591,N_23645,N_22230);
xnor U24592 (N_24592,N_23649,N_22312);
nor U24593 (N_24593,N_23160,N_23165);
and U24594 (N_24594,N_23089,N_23705);
nand U24595 (N_24595,N_23035,N_22144);
or U24596 (N_24596,N_22743,N_23518);
nor U24597 (N_24597,N_23822,N_22143);
xnor U24598 (N_24598,N_23722,N_23821);
nand U24599 (N_24599,N_22147,N_22146);
xor U24600 (N_24600,N_23152,N_22469);
xor U24601 (N_24601,N_23047,N_22974);
xor U24602 (N_24602,N_23049,N_23575);
xor U24603 (N_24603,N_22198,N_22855);
or U24604 (N_24604,N_22882,N_22861);
or U24605 (N_24605,N_23604,N_23956);
nor U24606 (N_24606,N_23456,N_23270);
or U24607 (N_24607,N_23408,N_23037);
nand U24608 (N_24608,N_23987,N_22562);
or U24609 (N_24609,N_23454,N_23607);
nand U24610 (N_24610,N_22956,N_22114);
nand U24611 (N_24611,N_23290,N_22222);
nor U24612 (N_24612,N_22689,N_22470);
and U24613 (N_24613,N_22933,N_23100);
nor U24614 (N_24614,N_23134,N_23921);
nand U24615 (N_24615,N_22296,N_22207);
or U24616 (N_24616,N_23426,N_22288);
nand U24617 (N_24617,N_23816,N_22717);
xnor U24618 (N_24618,N_23183,N_23878);
nand U24619 (N_24619,N_22310,N_23692);
nor U24620 (N_24620,N_23000,N_22950);
and U24621 (N_24621,N_22520,N_22459);
xnor U24622 (N_24622,N_23387,N_23818);
and U24623 (N_24623,N_22282,N_22525);
and U24624 (N_24624,N_23980,N_23605);
and U24625 (N_24625,N_22456,N_23093);
nand U24626 (N_24626,N_22468,N_23984);
and U24627 (N_24627,N_23238,N_23278);
or U24628 (N_24628,N_22714,N_22935);
nand U24629 (N_24629,N_23853,N_22475);
or U24630 (N_24630,N_23194,N_23887);
or U24631 (N_24631,N_23315,N_22821);
nor U24632 (N_24632,N_22886,N_22736);
nand U24633 (N_24633,N_22566,N_22794);
or U24634 (N_24634,N_23546,N_22632);
or U24635 (N_24635,N_22496,N_23004);
nand U24636 (N_24636,N_23052,N_22876);
and U24637 (N_24637,N_22534,N_22321);
and U24638 (N_24638,N_22783,N_22043);
nand U24639 (N_24639,N_22870,N_23979);
xor U24640 (N_24640,N_22265,N_22287);
and U24641 (N_24641,N_23805,N_23412);
or U24642 (N_24642,N_23282,N_23128);
and U24643 (N_24643,N_22180,N_23130);
nand U24644 (N_24644,N_22234,N_23938);
xnor U24645 (N_24645,N_22920,N_22900);
xnor U24646 (N_24646,N_23083,N_23425);
xor U24647 (N_24647,N_22902,N_22118);
or U24648 (N_24648,N_22433,N_22790);
nor U24649 (N_24649,N_23796,N_22047);
and U24650 (N_24650,N_23760,N_22161);
xnor U24651 (N_24651,N_23540,N_22489);
and U24652 (N_24652,N_22624,N_22938);
and U24653 (N_24653,N_22731,N_22406);
xor U24654 (N_24654,N_22068,N_23507);
xor U24655 (N_24655,N_23252,N_22569);
nor U24656 (N_24656,N_22691,N_23712);
nor U24657 (N_24657,N_23221,N_23883);
or U24658 (N_24658,N_22785,N_22263);
xor U24659 (N_24659,N_23392,N_23005);
and U24660 (N_24660,N_23661,N_23961);
nand U24661 (N_24661,N_23496,N_22062);
or U24662 (N_24662,N_23492,N_23565);
nor U24663 (N_24663,N_22013,N_22066);
nor U24664 (N_24664,N_22038,N_23828);
and U24665 (N_24665,N_23405,N_23787);
nor U24666 (N_24666,N_22930,N_23298);
xor U24667 (N_24667,N_23071,N_22278);
and U24668 (N_24668,N_23235,N_22862);
or U24669 (N_24669,N_23058,N_22032);
or U24670 (N_24670,N_23463,N_22868);
or U24671 (N_24671,N_23590,N_23549);
nand U24672 (N_24672,N_23121,N_22571);
xnor U24673 (N_24673,N_22416,N_22626);
or U24674 (N_24674,N_22630,N_23305);
xor U24675 (N_24675,N_22869,N_23797);
nand U24676 (N_24676,N_23890,N_22814);
xnor U24677 (N_24677,N_22067,N_23509);
or U24678 (N_24678,N_22410,N_22733);
and U24679 (N_24679,N_23253,N_23157);
or U24680 (N_24680,N_23233,N_22094);
and U24681 (N_24681,N_22228,N_22365);
xor U24682 (N_24682,N_22154,N_23250);
or U24683 (N_24683,N_22758,N_22149);
nor U24684 (N_24684,N_23829,N_22722);
or U24685 (N_24685,N_23922,N_23098);
nor U24686 (N_24686,N_22586,N_23555);
or U24687 (N_24687,N_23727,N_22625);
nand U24688 (N_24688,N_22167,N_23056);
and U24689 (N_24689,N_22665,N_23612);
nand U24690 (N_24690,N_22113,N_23857);
xor U24691 (N_24691,N_22092,N_22268);
nand U24692 (N_24692,N_22594,N_22776);
nand U24693 (N_24693,N_22317,N_22931);
nand U24694 (N_24694,N_22229,N_22726);
nand U24695 (N_24695,N_22454,N_22048);
and U24696 (N_24696,N_23048,N_22206);
nand U24697 (N_24697,N_23553,N_22664);
and U24698 (N_24698,N_23783,N_23147);
nor U24699 (N_24699,N_23245,N_23383);
and U24700 (N_24700,N_22813,N_22298);
nor U24701 (N_24701,N_23510,N_23815);
nand U24702 (N_24702,N_22747,N_23851);
xnor U24703 (N_24703,N_23638,N_22495);
xnor U24704 (N_24704,N_23951,N_23587);
xor U24705 (N_24705,N_22033,N_23265);
nand U24706 (N_24706,N_23520,N_23406);
nor U24707 (N_24707,N_22345,N_23826);
nor U24708 (N_24708,N_22355,N_22801);
and U24709 (N_24709,N_22192,N_23133);
or U24710 (N_24710,N_22342,N_22531);
nor U24711 (N_24711,N_22466,N_22647);
nand U24712 (N_24712,N_23032,N_22688);
or U24713 (N_24713,N_23926,N_23062);
nand U24714 (N_24714,N_22500,N_23377);
nor U24715 (N_24715,N_22145,N_23517);
and U24716 (N_24716,N_22792,N_22727);
xnor U24717 (N_24717,N_23401,N_23355);
nor U24718 (N_24718,N_22671,N_22964);
xnor U24719 (N_24719,N_23226,N_23578);
and U24720 (N_24720,N_23965,N_22865);
nand U24721 (N_24721,N_22740,N_23109);
or U24722 (N_24722,N_23691,N_23766);
nor U24723 (N_24723,N_22081,N_23434);
xnor U24724 (N_24724,N_22802,N_23025);
xnor U24725 (N_24725,N_22585,N_22160);
and U24726 (N_24726,N_23108,N_22095);
nor U24727 (N_24727,N_23488,N_22757);
or U24728 (N_24728,N_22965,N_23776);
nor U24729 (N_24729,N_23734,N_22996);
nor U24730 (N_24730,N_22565,N_23801);
or U24731 (N_24731,N_23172,N_23808);
xor U24732 (N_24732,N_22621,N_23411);
xor U24733 (N_24733,N_22028,N_23154);
nand U24734 (N_24734,N_23414,N_23896);
or U24735 (N_24735,N_23220,N_23897);
xnor U24736 (N_24736,N_23711,N_23349);
and U24737 (N_24737,N_22052,N_23471);
nand U24738 (N_24738,N_22178,N_23538);
or U24739 (N_24739,N_22400,N_22125);
nand U24740 (N_24740,N_23217,N_23174);
nand U24741 (N_24741,N_22330,N_22111);
and U24742 (N_24742,N_23582,N_22894);
or U24743 (N_24743,N_22227,N_22972);
and U24744 (N_24744,N_23500,N_22451);
or U24745 (N_24745,N_23511,N_23101);
or U24746 (N_24746,N_23541,N_23864);
and U24747 (N_24747,N_23362,N_22482);
and U24748 (N_24748,N_23350,N_23394);
nand U24749 (N_24749,N_22175,N_22059);
xor U24750 (N_24750,N_22769,N_23126);
nor U24751 (N_24751,N_23073,N_23060);
or U24752 (N_24752,N_23733,N_23944);
xnor U24753 (N_24753,N_22225,N_22197);
and U24754 (N_24754,N_23104,N_22065);
nand U24755 (N_24755,N_23875,N_22102);
nor U24756 (N_24756,N_22357,N_23081);
xor U24757 (N_24757,N_23481,N_22696);
or U24758 (N_24758,N_23988,N_23115);
nor U24759 (N_24759,N_22061,N_22005);
nand U24760 (N_24760,N_22361,N_23731);
nor U24761 (N_24761,N_23584,N_22120);
nand U24762 (N_24762,N_23482,N_22686);
nand U24763 (N_24763,N_22645,N_23610);
or U24764 (N_24764,N_22629,N_22863);
or U24765 (N_24765,N_22883,N_22084);
nand U24766 (N_24766,N_22903,N_22809);
nor U24767 (N_24767,N_22053,N_23095);
xnor U24768 (N_24768,N_22441,N_23239);
or U24769 (N_24769,N_22600,N_22879);
xor U24770 (N_24770,N_22713,N_23548);
or U24771 (N_24771,N_22946,N_22359);
nor U24772 (N_24772,N_23515,N_23484);
and U24773 (N_24773,N_23941,N_22806);
and U24774 (N_24774,N_23643,N_23261);
xnor U24775 (N_24775,N_22329,N_23924);
nor U24776 (N_24776,N_23777,N_22064);
nand U24777 (N_24777,N_23457,N_23954);
and U24778 (N_24778,N_23111,N_22220);
xor U24779 (N_24779,N_23544,N_22480);
xor U24780 (N_24780,N_23229,N_23090);
nor U24781 (N_24781,N_23169,N_22536);
nand U24782 (N_24782,N_22304,N_22690);
nand U24783 (N_24783,N_22376,N_22742);
xor U24784 (N_24784,N_23494,N_23171);
nor U24785 (N_24785,N_23843,N_22247);
nand U24786 (N_24786,N_23564,N_22984);
or U24787 (N_24787,N_23443,N_23567);
nand U24788 (N_24788,N_23196,N_22138);
nor U24789 (N_24789,N_22210,N_23256);
and U24790 (N_24790,N_22202,N_23650);
or U24791 (N_24791,N_22725,N_23341);
or U24792 (N_24792,N_22658,N_22506);
nor U24793 (N_24793,N_23292,N_22899);
xor U24794 (N_24794,N_23726,N_23962);
nor U24795 (N_24795,N_23739,N_23059);
nand U24796 (N_24796,N_23569,N_23028);
and U24797 (N_24797,N_23467,N_23861);
or U24798 (N_24798,N_22744,N_23923);
nor U24799 (N_24799,N_23784,N_22692);
nand U24800 (N_24800,N_22833,N_23672);
or U24801 (N_24801,N_23985,N_22721);
xnor U24802 (N_24802,N_22556,N_22982);
nand U24803 (N_24803,N_23308,N_22516);
nand U24804 (N_24804,N_22091,N_22545);
and U24805 (N_24805,N_23614,N_22511);
nand U24806 (N_24806,N_22914,N_23872);
nor U24807 (N_24807,N_22993,N_22675);
xor U24808 (N_24808,N_22131,N_23866);
xnor U24809 (N_24809,N_22588,N_22405);
or U24810 (N_24810,N_23996,N_23615);
nor U24811 (N_24811,N_22418,N_23942);
and U24812 (N_24812,N_22431,N_22054);
nor U24813 (N_24813,N_23385,N_23686);
nor U24814 (N_24814,N_23328,N_23653);
nor U24815 (N_24815,N_22951,N_22216);
or U24816 (N_24816,N_22579,N_22603);
and U24817 (N_24817,N_22548,N_23795);
nand U24818 (N_24818,N_22157,N_22948);
nor U24819 (N_24819,N_23817,N_22057);
and U24820 (N_24820,N_22781,N_23016);
xnor U24821 (N_24821,N_22460,N_22881);
nor U24822 (N_24822,N_23269,N_22905);
or U24823 (N_24823,N_23319,N_23831);
and U24824 (N_24824,N_22704,N_22300);
nor U24825 (N_24825,N_22362,N_23334);
nand U24826 (N_24826,N_23262,N_22711);
nor U24827 (N_24827,N_22916,N_22110);
and U24828 (N_24828,N_22798,N_23182);
nand U24829 (N_24829,N_23773,N_22823);
nor U24830 (N_24830,N_22252,N_23879);
nand U24831 (N_24831,N_23572,N_23273);
xor U24832 (N_24832,N_23399,N_23618);
and U24833 (N_24833,N_22462,N_23210);
and U24834 (N_24834,N_23763,N_22024);
or U24835 (N_24835,N_23759,N_23834);
or U24836 (N_24836,N_22457,N_23774);
or U24837 (N_24837,N_23246,N_23228);
nor U24838 (N_24838,N_23701,N_23698);
xnor U24839 (N_24839,N_23876,N_22845);
and U24840 (N_24840,N_22983,N_22353);
and U24841 (N_24841,N_23489,N_23775);
nor U24842 (N_24842,N_22786,N_22375);
or U24843 (N_24843,N_22644,N_22685);
and U24844 (N_24844,N_22515,N_22011);
or U24845 (N_24845,N_22646,N_22828);
xnor U24846 (N_24846,N_22169,N_23276);
xor U24847 (N_24847,N_22682,N_22620);
or U24848 (N_24848,N_22841,N_22465);
or U24849 (N_24849,N_23402,N_23952);
nand U24850 (N_24850,N_22981,N_23665);
nor U24851 (N_24851,N_22584,N_22425);
nor U24852 (N_24852,N_23682,N_23598);
nand U24853 (N_24853,N_23608,N_23856);
xnor U24854 (N_24854,N_23022,N_22308);
nand U24855 (N_24855,N_23709,N_22698);
nor U24856 (N_24856,N_22640,N_22988);
or U24857 (N_24857,N_22284,N_22501);
nor U24858 (N_24858,N_23118,N_23632);
nand U24859 (N_24859,N_22275,N_22150);
or U24860 (N_24860,N_23624,N_22486);
or U24861 (N_24861,N_22370,N_22576);
and U24862 (N_24862,N_22680,N_22001);
or U24863 (N_24863,N_22476,N_22892);
nor U24864 (N_24864,N_23679,N_22732);
or U24865 (N_24865,N_23272,N_23373);
nor U24866 (N_24866,N_23998,N_22527);
nand U24867 (N_24867,N_23386,N_23535);
or U24868 (N_24868,N_22546,N_23611);
nand U24869 (N_24869,N_22453,N_23681);
and U24870 (N_24870,N_22555,N_23129);
nand U24871 (N_24871,N_22539,N_22552);
or U24872 (N_24872,N_23200,N_22337);
xor U24873 (N_24873,N_23858,N_23975);
and U24874 (N_24874,N_23995,N_23243);
nor U24875 (N_24875,N_22432,N_23175);
xor U24876 (N_24876,N_23753,N_22660);
nor U24877 (N_24877,N_23280,N_22775);
nand U24878 (N_24878,N_22936,N_22218);
xor U24879 (N_24879,N_23870,N_23103);
and U24880 (N_24880,N_23078,N_23162);
and U24881 (N_24881,N_23811,N_23868);
and U24882 (N_24882,N_23793,N_23648);
and U24883 (N_24883,N_23623,N_22768);
nand U24884 (N_24884,N_23450,N_22124);
xnor U24885 (N_24885,N_23895,N_22904);
nor U24886 (N_24886,N_23963,N_23380);
and U24887 (N_24887,N_23449,N_23311);
nand U24888 (N_24888,N_23576,N_23378);
nand U24889 (N_24889,N_23899,N_22007);
or U24890 (N_24890,N_23097,N_23330);
nor U24891 (N_24891,N_23085,N_23177);
or U24892 (N_24892,N_23732,N_23919);
nand U24893 (N_24893,N_23205,N_22134);
nor U24894 (N_24894,N_22999,N_22602);
xnor U24895 (N_24895,N_23631,N_22439);
nor U24896 (N_24896,N_23986,N_23736);
or U24897 (N_24897,N_22189,N_23189);
nor U24898 (N_24898,N_22641,N_23554);
or U24899 (N_24899,N_23369,N_23593);
or U24900 (N_24900,N_22086,N_23198);
xor U24901 (N_24901,N_22070,N_23602);
xor U24902 (N_24902,N_22242,N_22898);
nand U24903 (N_24903,N_23566,N_23255);
and U24904 (N_24904,N_22231,N_22709);
and U24905 (N_24905,N_22678,N_23230);
and U24906 (N_24906,N_23788,N_22273);
nor U24907 (N_24907,N_23522,N_22729);
nand U24908 (N_24908,N_22436,N_22088);
and U24909 (N_24909,N_22992,N_22430);
or U24910 (N_24910,N_22517,N_22404);
nand U24911 (N_24911,N_23628,N_23258);
xnor U24912 (N_24912,N_22958,N_22046);
or U24913 (N_24913,N_22507,N_23603);
or U24914 (N_24914,N_22991,N_22955);
and U24915 (N_24915,N_23903,N_23599);
nand U24916 (N_24916,N_23395,N_23737);
nor U24917 (N_24917,N_23381,N_22494);
and U24918 (N_24918,N_23688,N_22940);
and U24919 (N_24919,N_22063,N_23300);
xor U24920 (N_24920,N_23621,N_22266);
nand U24921 (N_24921,N_23429,N_23504);
nand U24922 (N_24922,N_23677,N_23754);
nor U24923 (N_24923,N_23740,N_23222);
or U24924 (N_24924,N_22739,N_23094);
xnor U24925 (N_24925,N_22921,N_23958);
nor U24926 (N_24926,N_22472,N_23495);
and U24927 (N_24927,N_22980,N_22707);
and U24928 (N_24928,N_23561,N_23159);
nor U24929 (N_24929,N_23014,N_23043);
nor U24930 (N_24930,N_22148,N_22049);
or U24931 (N_24931,N_23673,N_23391);
and U24932 (N_24932,N_22452,N_23287);
nor U24933 (N_24933,N_23325,N_22810);
or U24934 (N_24934,N_22593,N_22437);
and U24935 (N_24935,N_23839,N_22738);
or U24936 (N_24936,N_23646,N_22448);
or U24937 (N_24937,N_22003,N_22331);
nand U24938 (N_24938,N_22590,N_23708);
xor U24939 (N_24939,N_22214,N_22385);
nor U24940 (N_24940,N_22795,N_23168);
nor U24941 (N_24941,N_22291,N_22251);
and U24942 (N_24942,N_22723,N_23389);
nor U24943 (N_24943,N_22398,N_22200);
xor U24944 (N_24944,N_22919,N_23669);
and U24945 (N_24945,N_22943,N_22927);
nor U24946 (N_24946,N_22055,N_22079);
or U24947 (N_24947,N_22080,N_22264);
and U24948 (N_24948,N_23140,N_22695);
xor U24949 (N_24949,N_23345,N_22997);
xor U24950 (N_24950,N_22074,N_22072);
xnor U24951 (N_24951,N_22444,N_23659);
or U24952 (N_24952,N_22844,N_22389);
nor U24953 (N_24953,N_23288,N_22901);
nor U24954 (N_24954,N_22578,N_22573);
and U24955 (N_24955,N_22954,N_22985);
or U24956 (N_24956,N_22924,N_23493);
xnor U24957 (N_24957,N_22553,N_23204);
nand U24958 (N_24958,N_23823,N_23301);
or U24959 (N_24959,N_22372,N_22800);
nand U24960 (N_24960,N_22651,N_23978);
nor U24961 (N_24961,N_22191,N_23251);
nor U24962 (N_24962,N_23419,N_22136);
nand U24963 (N_24963,N_23438,N_23704);
xnor U24964 (N_24964,N_23161,N_23780);
nand U24965 (N_24965,N_23348,N_22155);
or U24966 (N_24966,N_23077,N_23193);
xor U24967 (N_24967,N_22364,N_22811);
nor U24968 (N_24968,N_23303,N_23983);
and U24969 (N_24969,N_22945,N_22347);
nand U24970 (N_24970,N_23644,N_22142);
or U24971 (N_24971,N_22194,N_22605);
or U24972 (N_24972,N_22176,N_22701);
nor U24973 (N_24973,N_22976,N_23370);
and U24974 (N_24974,N_22269,N_23528);
nor U24975 (N_24975,N_23936,N_22205);
nand U24976 (N_24976,N_22315,N_23908);
xor U24977 (N_24977,N_22463,N_22044);
xor U24978 (N_24978,N_23925,N_23581);
and U24979 (N_24979,N_22075,N_23415);
nor U24980 (N_24980,N_22797,N_23332);
nand U24981 (N_24981,N_22037,N_22165);
and U24982 (N_24982,N_23629,N_22654);
xor U24983 (N_24983,N_22967,N_22706);
and U24984 (N_24984,N_23455,N_22069);
and U24985 (N_24985,N_23931,N_23284);
or U24986 (N_24986,N_22705,N_23469);
nand U24987 (N_24987,N_22617,N_22215);
and U24988 (N_24988,N_23445,N_22159);
xnor U24989 (N_24989,N_22369,N_23365);
or U24990 (N_24990,N_22035,N_22249);
xnor U24991 (N_24991,N_22488,N_22384);
xor U24992 (N_24992,N_23299,N_23110);
nand U24993 (N_24993,N_22872,N_22168);
or U24994 (N_24994,N_22547,N_22314);
nand U24995 (N_24995,N_22241,N_22272);
or U24996 (N_24996,N_22443,N_22541);
nor U24997 (N_24997,N_22440,N_23388);
nor U24998 (N_24998,N_23802,N_22540);
xnor U24999 (N_24999,N_22896,N_22402);
nor U25000 (N_25000,N_23927,N_22442);
nor U25001 (N_25001,N_23929,N_23833);
nand U25002 (N_25002,N_23065,N_22403);
nor U25003 (N_25003,N_22771,N_22471);
nand U25004 (N_25004,N_22689,N_23230);
xor U25005 (N_25005,N_22398,N_23365);
nand U25006 (N_25006,N_23643,N_22171);
xnor U25007 (N_25007,N_23357,N_22027);
xor U25008 (N_25008,N_22099,N_23536);
and U25009 (N_25009,N_23085,N_22192);
xor U25010 (N_25010,N_23719,N_23006);
nand U25011 (N_25011,N_23678,N_22429);
or U25012 (N_25012,N_23487,N_23960);
or U25013 (N_25013,N_22425,N_23064);
nor U25014 (N_25014,N_23512,N_22935);
nand U25015 (N_25015,N_22289,N_23252);
xnor U25016 (N_25016,N_22432,N_23027);
nand U25017 (N_25017,N_23113,N_22294);
or U25018 (N_25018,N_23427,N_23708);
nor U25019 (N_25019,N_22023,N_23045);
xnor U25020 (N_25020,N_22776,N_23309);
or U25021 (N_25021,N_23002,N_23883);
nor U25022 (N_25022,N_22213,N_22465);
nand U25023 (N_25023,N_22388,N_23664);
or U25024 (N_25024,N_22842,N_23431);
xnor U25025 (N_25025,N_22273,N_23000);
nor U25026 (N_25026,N_23335,N_22418);
and U25027 (N_25027,N_23586,N_23432);
xor U25028 (N_25028,N_22690,N_22955);
nor U25029 (N_25029,N_22447,N_23016);
and U25030 (N_25030,N_22359,N_23127);
nor U25031 (N_25031,N_23572,N_23441);
and U25032 (N_25032,N_23711,N_22710);
nand U25033 (N_25033,N_22102,N_22183);
xor U25034 (N_25034,N_23415,N_23505);
nor U25035 (N_25035,N_22942,N_23509);
and U25036 (N_25036,N_22165,N_22949);
xnor U25037 (N_25037,N_23592,N_22835);
nand U25038 (N_25038,N_22259,N_22996);
and U25039 (N_25039,N_23256,N_23075);
or U25040 (N_25040,N_23682,N_23971);
or U25041 (N_25041,N_23093,N_23446);
xnor U25042 (N_25042,N_23367,N_23810);
and U25043 (N_25043,N_23656,N_22128);
nor U25044 (N_25044,N_22381,N_23703);
nand U25045 (N_25045,N_22660,N_23843);
xnor U25046 (N_25046,N_23337,N_22084);
nor U25047 (N_25047,N_23903,N_22320);
nor U25048 (N_25048,N_22231,N_23956);
nand U25049 (N_25049,N_22639,N_22072);
nand U25050 (N_25050,N_23615,N_23770);
or U25051 (N_25051,N_23272,N_23855);
and U25052 (N_25052,N_23291,N_23967);
nor U25053 (N_25053,N_23774,N_22519);
nand U25054 (N_25054,N_22198,N_23713);
or U25055 (N_25055,N_23310,N_23298);
xor U25056 (N_25056,N_23287,N_23325);
nor U25057 (N_25057,N_23043,N_22517);
and U25058 (N_25058,N_23252,N_22235);
xnor U25059 (N_25059,N_23709,N_23625);
and U25060 (N_25060,N_23036,N_22660);
nand U25061 (N_25061,N_22951,N_23062);
or U25062 (N_25062,N_22318,N_22006);
nand U25063 (N_25063,N_23367,N_23294);
or U25064 (N_25064,N_23852,N_23253);
nand U25065 (N_25065,N_22224,N_23177);
nor U25066 (N_25066,N_23342,N_22652);
and U25067 (N_25067,N_22186,N_22325);
or U25068 (N_25068,N_22948,N_22225);
xnor U25069 (N_25069,N_22066,N_22813);
xor U25070 (N_25070,N_22379,N_22131);
nor U25071 (N_25071,N_23209,N_22840);
and U25072 (N_25072,N_22356,N_22389);
nand U25073 (N_25073,N_23414,N_22520);
xor U25074 (N_25074,N_22888,N_23150);
nor U25075 (N_25075,N_22069,N_22780);
and U25076 (N_25076,N_23195,N_23113);
or U25077 (N_25077,N_23258,N_23461);
nor U25078 (N_25078,N_22375,N_23977);
or U25079 (N_25079,N_23165,N_22735);
and U25080 (N_25080,N_23575,N_22128);
and U25081 (N_25081,N_23315,N_23262);
nand U25082 (N_25082,N_22225,N_22187);
nor U25083 (N_25083,N_22363,N_23915);
or U25084 (N_25084,N_22429,N_23590);
and U25085 (N_25085,N_23055,N_22794);
and U25086 (N_25086,N_22171,N_23928);
nor U25087 (N_25087,N_22922,N_22011);
and U25088 (N_25088,N_23591,N_22719);
nand U25089 (N_25089,N_23892,N_23294);
or U25090 (N_25090,N_23124,N_22196);
xnor U25091 (N_25091,N_22620,N_22569);
and U25092 (N_25092,N_23817,N_22574);
nor U25093 (N_25093,N_23521,N_22601);
or U25094 (N_25094,N_22745,N_22608);
nand U25095 (N_25095,N_22433,N_22277);
and U25096 (N_25096,N_22289,N_23629);
and U25097 (N_25097,N_22998,N_22684);
nand U25098 (N_25098,N_22450,N_22490);
nand U25099 (N_25099,N_22283,N_23399);
or U25100 (N_25100,N_22360,N_23278);
nand U25101 (N_25101,N_22362,N_22338);
xor U25102 (N_25102,N_22040,N_23966);
or U25103 (N_25103,N_22384,N_22894);
nand U25104 (N_25104,N_22308,N_23680);
nand U25105 (N_25105,N_22645,N_23903);
nand U25106 (N_25106,N_22902,N_22268);
nor U25107 (N_25107,N_23831,N_22281);
nand U25108 (N_25108,N_22811,N_23107);
or U25109 (N_25109,N_23371,N_22572);
nor U25110 (N_25110,N_23817,N_22797);
xnor U25111 (N_25111,N_23653,N_22959);
or U25112 (N_25112,N_23295,N_22318);
or U25113 (N_25113,N_23889,N_22300);
or U25114 (N_25114,N_22706,N_23230);
nor U25115 (N_25115,N_22503,N_22419);
or U25116 (N_25116,N_23876,N_22881);
nand U25117 (N_25117,N_22835,N_23467);
nor U25118 (N_25118,N_23360,N_23325);
or U25119 (N_25119,N_22955,N_23100);
or U25120 (N_25120,N_23917,N_23192);
nor U25121 (N_25121,N_23451,N_22475);
and U25122 (N_25122,N_23012,N_23234);
xnor U25123 (N_25123,N_23202,N_22172);
nand U25124 (N_25124,N_22816,N_22684);
and U25125 (N_25125,N_23511,N_22080);
nor U25126 (N_25126,N_23299,N_23680);
or U25127 (N_25127,N_22298,N_22329);
nor U25128 (N_25128,N_22279,N_23856);
and U25129 (N_25129,N_22678,N_23254);
and U25130 (N_25130,N_22583,N_22881);
or U25131 (N_25131,N_22549,N_22315);
nor U25132 (N_25132,N_23300,N_23325);
or U25133 (N_25133,N_22511,N_22736);
and U25134 (N_25134,N_23866,N_23480);
nor U25135 (N_25135,N_23679,N_23959);
xnor U25136 (N_25136,N_22731,N_22733);
and U25137 (N_25137,N_22118,N_22317);
and U25138 (N_25138,N_23955,N_23714);
nand U25139 (N_25139,N_22850,N_22899);
nor U25140 (N_25140,N_22777,N_23305);
xor U25141 (N_25141,N_22215,N_22558);
and U25142 (N_25142,N_22871,N_22677);
nor U25143 (N_25143,N_22585,N_22091);
xnor U25144 (N_25144,N_23807,N_22683);
or U25145 (N_25145,N_22116,N_23532);
or U25146 (N_25146,N_22322,N_23274);
xnor U25147 (N_25147,N_22082,N_22042);
nor U25148 (N_25148,N_22722,N_23444);
nor U25149 (N_25149,N_23339,N_22656);
xor U25150 (N_25150,N_22395,N_22873);
or U25151 (N_25151,N_23314,N_22337);
nor U25152 (N_25152,N_23986,N_23517);
nand U25153 (N_25153,N_23393,N_23129);
nor U25154 (N_25154,N_22466,N_23404);
nand U25155 (N_25155,N_22016,N_22043);
nand U25156 (N_25156,N_23155,N_23466);
nor U25157 (N_25157,N_22032,N_22702);
nor U25158 (N_25158,N_23304,N_23764);
nand U25159 (N_25159,N_23328,N_23860);
or U25160 (N_25160,N_22737,N_22262);
and U25161 (N_25161,N_22528,N_22536);
xnor U25162 (N_25162,N_23310,N_22489);
or U25163 (N_25163,N_22139,N_22190);
nand U25164 (N_25164,N_22222,N_23782);
nor U25165 (N_25165,N_22915,N_23179);
xor U25166 (N_25166,N_23077,N_23925);
nand U25167 (N_25167,N_23922,N_22875);
nand U25168 (N_25168,N_22214,N_23656);
or U25169 (N_25169,N_22145,N_22000);
xor U25170 (N_25170,N_23001,N_23245);
xnor U25171 (N_25171,N_22058,N_23446);
or U25172 (N_25172,N_22238,N_23643);
or U25173 (N_25173,N_22415,N_22505);
xnor U25174 (N_25174,N_23556,N_23286);
xnor U25175 (N_25175,N_23098,N_22667);
or U25176 (N_25176,N_23690,N_22681);
nor U25177 (N_25177,N_22391,N_23153);
xor U25178 (N_25178,N_22505,N_22924);
nor U25179 (N_25179,N_23512,N_23371);
nand U25180 (N_25180,N_23560,N_23864);
xor U25181 (N_25181,N_23445,N_23563);
xor U25182 (N_25182,N_22389,N_22865);
nor U25183 (N_25183,N_23721,N_22504);
and U25184 (N_25184,N_23143,N_23275);
nand U25185 (N_25185,N_23022,N_23224);
nand U25186 (N_25186,N_23451,N_22034);
nor U25187 (N_25187,N_23631,N_22510);
xor U25188 (N_25188,N_22779,N_23927);
and U25189 (N_25189,N_23608,N_22374);
and U25190 (N_25190,N_22028,N_23843);
nand U25191 (N_25191,N_23232,N_23140);
nand U25192 (N_25192,N_22365,N_23045);
nor U25193 (N_25193,N_23305,N_22254);
xnor U25194 (N_25194,N_23010,N_23617);
nand U25195 (N_25195,N_23428,N_22317);
nor U25196 (N_25196,N_22437,N_22761);
nor U25197 (N_25197,N_23902,N_23114);
and U25198 (N_25198,N_22813,N_22593);
xor U25199 (N_25199,N_22654,N_22333);
and U25200 (N_25200,N_23126,N_22287);
nor U25201 (N_25201,N_23858,N_22778);
nor U25202 (N_25202,N_22244,N_23907);
and U25203 (N_25203,N_22968,N_22238);
xor U25204 (N_25204,N_22213,N_23951);
and U25205 (N_25205,N_23626,N_22161);
and U25206 (N_25206,N_23148,N_22310);
or U25207 (N_25207,N_23913,N_22640);
and U25208 (N_25208,N_23287,N_23432);
or U25209 (N_25209,N_23204,N_23049);
xor U25210 (N_25210,N_23474,N_22692);
nand U25211 (N_25211,N_22047,N_22984);
nor U25212 (N_25212,N_23994,N_23836);
nor U25213 (N_25213,N_23192,N_23902);
nor U25214 (N_25214,N_23732,N_22311);
xnor U25215 (N_25215,N_22862,N_23559);
or U25216 (N_25216,N_22524,N_23295);
or U25217 (N_25217,N_22683,N_23542);
xnor U25218 (N_25218,N_23731,N_22671);
and U25219 (N_25219,N_23930,N_22267);
nor U25220 (N_25220,N_22224,N_23322);
or U25221 (N_25221,N_23932,N_22711);
nand U25222 (N_25222,N_23625,N_23066);
xor U25223 (N_25223,N_23651,N_23932);
nand U25224 (N_25224,N_22008,N_22416);
xor U25225 (N_25225,N_23551,N_22076);
and U25226 (N_25226,N_22320,N_23035);
nand U25227 (N_25227,N_22889,N_22234);
nand U25228 (N_25228,N_22148,N_23685);
or U25229 (N_25229,N_23744,N_22401);
xor U25230 (N_25230,N_22252,N_23479);
or U25231 (N_25231,N_23675,N_23003);
nand U25232 (N_25232,N_23320,N_23519);
xor U25233 (N_25233,N_23216,N_23331);
and U25234 (N_25234,N_22906,N_22871);
nor U25235 (N_25235,N_22367,N_22852);
xor U25236 (N_25236,N_22481,N_23796);
nand U25237 (N_25237,N_22912,N_22587);
or U25238 (N_25238,N_22366,N_22633);
or U25239 (N_25239,N_22906,N_23401);
and U25240 (N_25240,N_22799,N_22697);
nand U25241 (N_25241,N_23760,N_22703);
or U25242 (N_25242,N_22330,N_23631);
xnor U25243 (N_25243,N_23469,N_23901);
nand U25244 (N_25244,N_22011,N_22829);
or U25245 (N_25245,N_23626,N_22403);
nor U25246 (N_25246,N_23050,N_22886);
or U25247 (N_25247,N_23776,N_23281);
or U25248 (N_25248,N_23565,N_23189);
xor U25249 (N_25249,N_22017,N_22319);
and U25250 (N_25250,N_22326,N_22131);
or U25251 (N_25251,N_23924,N_23147);
nand U25252 (N_25252,N_22263,N_22744);
or U25253 (N_25253,N_22629,N_22274);
or U25254 (N_25254,N_23014,N_23805);
or U25255 (N_25255,N_22728,N_23725);
or U25256 (N_25256,N_23679,N_23754);
and U25257 (N_25257,N_22820,N_23658);
nor U25258 (N_25258,N_23295,N_22093);
or U25259 (N_25259,N_23185,N_22058);
nand U25260 (N_25260,N_22297,N_22832);
or U25261 (N_25261,N_23075,N_23081);
or U25262 (N_25262,N_23213,N_22107);
and U25263 (N_25263,N_22569,N_23055);
or U25264 (N_25264,N_22794,N_22646);
or U25265 (N_25265,N_23651,N_22305);
and U25266 (N_25266,N_23717,N_22795);
or U25267 (N_25267,N_23638,N_22327);
xor U25268 (N_25268,N_22354,N_22570);
or U25269 (N_25269,N_23629,N_22134);
nand U25270 (N_25270,N_23507,N_22862);
and U25271 (N_25271,N_22600,N_23263);
and U25272 (N_25272,N_22328,N_22770);
nand U25273 (N_25273,N_22343,N_22916);
or U25274 (N_25274,N_23977,N_22586);
and U25275 (N_25275,N_23601,N_22247);
nand U25276 (N_25276,N_22236,N_22798);
nand U25277 (N_25277,N_22020,N_23483);
nor U25278 (N_25278,N_23972,N_23520);
xnor U25279 (N_25279,N_22429,N_23534);
nand U25280 (N_25280,N_23324,N_23853);
and U25281 (N_25281,N_22134,N_23291);
xnor U25282 (N_25282,N_23588,N_23315);
nand U25283 (N_25283,N_23042,N_22676);
or U25284 (N_25284,N_23871,N_23762);
nand U25285 (N_25285,N_23400,N_22337);
nor U25286 (N_25286,N_23473,N_23838);
or U25287 (N_25287,N_23936,N_23098);
nand U25288 (N_25288,N_22856,N_23444);
nor U25289 (N_25289,N_22314,N_23723);
and U25290 (N_25290,N_22344,N_23841);
or U25291 (N_25291,N_23757,N_23898);
nand U25292 (N_25292,N_23412,N_22721);
or U25293 (N_25293,N_22494,N_22474);
xnor U25294 (N_25294,N_22872,N_22472);
and U25295 (N_25295,N_23556,N_23629);
and U25296 (N_25296,N_22527,N_22605);
nor U25297 (N_25297,N_23716,N_23584);
nor U25298 (N_25298,N_22396,N_23503);
nor U25299 (N_25299,N_23980,N_22093);
nor U25300 (N_25300,N_23100,N_22771);
or U25301 (N_25301,N_22101,N_22561);
or U25302 (N_25302,N_23931,N_23161);
and U25303 (N_25303,N_22697,N_22188);
and U25304 (N_25304,N_22251,N_22745);
and U25305 (N_25305,N_22449,N_22244);
nor U25306 (N_25306,N_23656,N_22588);
nor U25307 (N_25307,N_23828,N_22668);
nor U25308 (N_25308,N_22613,N_22795);
nor U25309 (N_25309,N_22126,N_23928);
nand U25310 (N_25310,N_23047,N_23839);
nand U25311 (N_25311,N_23685,N_23912);
or U25312 (N_25312,N_22721,N_23013);
xnor U25313 (N_25313,N_22370,N_23495);
and U25314 (N_25314,N_23186,N_22457);
or U25315 (N_25315,N_22733,N_22965);
xnor U25316 (N_25316,N_22427,N_23389);
xnor U25317 (N_25317,N_23100,N_22113);
nor U25318 (N_25318,N_23304,N_22485);
nand U25319 (N_25319,N_22362,N_23093);
or U25320 (N_25320,N_22846,N_22477);
nor U25321 (N_25321,N_22213,N_22022);
xnor U25322 (N_25322,N_22822,N_22192);
xnor U25323 (N_25323,N_22748,N_23646);
nor U25324 (N_25324,N_22741,N_22514);
or U25325 (N_25325,N_23045,N_22534);
xor U25326 (N_25326,N_22265,N_22267);
or U25327 (N_25327,N_23365,N_23393);
or U25328 (N_25328,N_22103,N_23377);
xnor U25329 (N_25329,N_23017,N_23772);
and U25330 (N_25330,N_22398,N_22716);
nor U25331 (N_25331,N_23982,N_23215);
or U25332 (N_25332,N_23416,N_23868);
and U25333 (N_25333,N_23179,N_22009);
and U25334 (N_25334,N_22740,N_22115);
nand U25335 (N_25335,N_22569,N_22342);
nor U25336 (N_25336,N_22846,N_22639);
or U25337 (N_25337,N_22060,N_22006);
xnor U25338 (N_25338,N_23126,N_22280);
and U25339 (N_25339,N_22705,N_22262);
nand U25340 (N_25340,N_23883,N_23030);
nand U25341 (N_25341,N_22974,N_22519);
nand U25342 (N_25342,N_22044,N_23316);
xor U25343 (N_25343,N_23599,N_23556);
nand U25344 (N_25344,N_23211,N_23840);
and U25345 (N_25345,N_23025,N_23725);
xnor U25346 (N_25346,N_23298,N_23284);
xor U25347 (N_25347,N_22784,N_23833);
and U25348 (N_25348,N_22840,N_22766);
and U25349 (N_25349,N_23911,N_23538);
and U25350 (N_25350,N_23055,N_22307);
nor U25351 (N_25351,N_23691,N_22834);
nand U25352 (N_25352,N_22206,N_23225);
nand U25353 (N_25353,N_23812,N_22414);
or U25354 (N_25354,N_23634,N_23491);
nor U25355 (N_25355,N_23656,N_22459);
or U25356 (N_25356,N_23862,N_23265);
nor U25357 (N_25357,N_23194,N_23088);
and U25358 (N_25358,N_23780,N_23654);
and U25359 (N_25359,N_23326,N_23435);
and U25360 (N_25360,N_22286,N_22148);
or U25361 (N_25361,N_22890,N_23809);
xnor U25362 (N_25362,N_23830,N_22468);
nor U25363 (N_25363,N_22908,N_22253);
or U25364 (N_25364,N_22686,N_22061);
nor U25365 (N_25365,N_23104,N_22069);
nand U25366 (N_25366,N_23132,N_22925);
nand U25367 (N_25367,N_23305,N_23926);
or U25368 (N_25368,N_23773,N_22985);
nor U25369 (N_25369,N_23939,N_22708);
and U25370 (N_25370,N_22857,N_23064);
nand U25371 (N_25371,N_23843,N_22959);
nand U25372 (N_25372,N_23575,N_23439);
nor U25373 (N_25373,N_23709,N_23050);
nand U25374 (N_25374,N_22451,N_22298);
xor U25375 (N_25375,N_22361,N_23603);
nand U25376 (N_25376,N_23364,N_22511);
or U25377 (N_25377,N_23015,N_22213);
nand U25378 (N_25378,N_22919,N_23881);
nor U25379 (N_25379,N_22598,N_23586);
nor U25380 (N_25380,N_23433,N_23044);
xor U25381 (N_25381,N_22062,N_22815);
nor U25382 (N_25382,N_23441,N_22331);
and U25383 (N_25383,N_22672,N_23415);
xor U25384 (N_25384,N_23721,N_23295);
nand U25385 (N_25385,N_23417,N_23710);
and U25386 (N_25386,N_23742,N_23006);
nand U25387 (N_25387,N_23780,N_22794);
xnor U25388 (N_25388,N_22971,N_22079);
and U25389 (N_25389,N_22065,N_23356);
or U25390 (N_25390,N_22831,N_22460);
or U25391 (N_25391,N_22909,N_22795);
xnor U25392 (N_25392,N_22269,N_22253);
xnor U25393 (N_25393,N_23121,N_22958);
nor U25394 (N_25394,N_22172,N_23987);
xnor U25395 (N_25395,N_23740,N_23686);
xor U25396 (N_25396,N_22813,N_23099);
nor U25397 (N_25397,N_22761,N_22882);
nand U25398 (N_25398,N_23815,N_22332);
and U25399 (N_25399,N_22466,N_23841);
nor U25400 (N_25400,N_22601,N_22432);
or U25401 (N_25401,N_22708,N_23178);
or U25402 (N_25402,N_22838,N_22675);
and U25403 (N_25403,N_23948,N_23609);
or U25404 (N_25404,N_22805,N_22949);
and U25405 (N_25405,N_23322,N_22981);
xnor U25406 (N_25406,N_23586,N_22562);
xor U25407 (N_25407,N_23329,N_23351);
and U25408 (N_25408,N_22777,N_23187);
xor U25409 (N_25409,N_22241,N_22019);
nand U25410 (N_25410,N_23463,N_22388);
nor U25411 (N_25411,N_22420,N_23042);
and U25412 (N_25412,N_22233,N_22530);
nor U25413 (N_25413,N_22808,N_22260);
xnor U25414 (N_25414,N_22462,N_22475);
nand U25415 (N_25415,N_22709,N_22221);
xor U25416 (N_25416,N_22013,N_22144);
or U25417 (N_25417,N_23858,N_22507);
nand U25418 (N_25418,N_23615,N_22774);
and U25419 (N_25419,N_23176,N_23720);
nand U25420 (N_25420,N_23663,N_22702);
nor U25421 (N_25421,N_22334,N_22364);
nor U25422 (N_25422,N_23245,N_23368);
xor U25423 (N_25423,N_22254,N_22296);
nand U25424 (N_25424,N_22338,N_22980);
nor U25425 (N_25425,N_23542,N_23296);
xnor U25426 (N_25426,N_22906,N_23300);
or U25427 (N_25427,N_22922,N_22719);
nor U25428 (N_25428,N_22438,N_23505);
nand U25429 (N_25429,N_23202,N_22178);
nand U25430 (N_25430,N_22285,N_23618);
or U25431 (N_25431,N_23279,N_23476);
and U25432 (N_25432,N_23661,N_23297);
or U25433 (N_25433,N_22878,N_23890);
nor U25434 (N_25434,N_22306,N_22712);
and U25435 (N_25435,N_22971,N_23199);
nand U25436 (N_25436,N_23051,N_23426);
and U25437 (N_25437,N_23991,N_22569);
nor U25438 (N_25438,N_23676,N_22506);
nor U25439 (N_25439,N_23581,N_23521);
or U25440 (N_25440,N_22984,N_22884);
nand U25441 (N_25441,N_22533,N_22427);
or U25442 (N_25442,N_22155,N_23408);
xnor U25443 (N_25443,N_22649,N_22972);
nor U25444 (N_25444,N_22722,N_23963);
and U25445 (N_25445,N_23613,N_23727);
xnor U25446 (N_25446,N_23706,N_23332);
nor U25447 (N_25447,N_22027,N_22276);
nor U25448 (N_25448,N_22205,N_22689);
or U25449 (N_25449,N_23799,N_22187);
xnor U25450 (N_25450,N_23447,N_22214);
and U25451 (N_25451,N_23352,N_23375);
or U25452 (N_25452,N_22100,N_22975);
nor U25453 (N_25453,N_22447,N_23040);
xnor U25454 (N_25454,N_22120,N_22139);
or U25455 (N_25455,N_22303,N_22307);
or U25456 (N_25456,N_22656,N_23537);
xnor U25457 (N_25457,N_23124,N_23343);
and U25458 (N_25458,N_22402,N_23739);
xor U25459 (N_25459,N_23269,N_23166);
and U25460 (N_25460,N_22394,N_23983);
xor U25461 (N_25461,N_22781,N_23068);
or U25462 (N_25462,N_22146,N_23930);
nand U25463 (N_25463,N_23686,N_22240);
nor U25464 (N_25464,N_23211,N_22665);
nor U25465 (N_25465,N_23013,N_22991);
nor U25466 (N_25466,N_22057,N_23926);
xor U25467 (N_25467,N_23210,N_22869);
and U25468 (N_25468,N_22334,N_23524);
or U25469 (N_25469,N_22366,N_22435);
and U25470 (N_25470,N_23404,N_23190);
xor U25471 (N_25471,N_22117,N_23667);
xnor U25472 (N_25472,N_23650,N_22180);
or U25473 (N_25473,N_22405,N_22823);
or U25474 (N_25474,N_22831,N_23360);
xnor U25475 (N_25475,N_22903,N_22040);
nor U25476 (N_25476,N_23448,N_23147);
nor U25477 (N_25477,N_23286,N_22696);
nor U25478 (N_25478,N_23374,N_23749);
xor U25479 (N_25479,N_22381,N_23135);
nor U25480 (N_25480,N_23690,N_23107);
nor U25481 (N_25481,N_23988,N_23860);
nor U25482 (N_25482,N_22582,N_22765);
nor U25483 (N_25483,N_22973,N_23095);
nand U25484 (N_25484,N_23380,N_23973);
and U25485 (N_25485,N_22905,N_22955);
nand U25486 (N_25486,N_23870,N_23680);
nor U25487 (N_25487,N_22567,N_23501);
and U25488 (N_25488,N_23898,N_23986);
nor U25489 (N_25489,N_22253,N_23894);
xor U25490 (N_25490,N_22851,N_23479);
or U25491 (N_25491,N_23372,N_22084);
xnor U25492 (N_25492,N_22420,N_23379);
nand U25493 (N_25493,N_22680,N_23223);
or U25494 (N_25494,N_22760,N_23080);
xnor U25495 (N_25495,N_23652,N_23502);
nand U25496 (N_25496,N_23850,N_22730);
or U25497 (N_25497,N_23666,N_22065);
nand U25498 (N_25498,N_23136,N_23079);
nor U25499 (N_25499,N_23793,N_22292);
or U25500 (N_25500,N_22722,N_22762);
nor U25501 (N_25501,N_22690,N_22282);
and U25502 (N_25502,N_23058,N_23497);
and U25503 (N_25503,N_22466,N_22912);
xnor U25504 (N_25504,N_22650,N_23253);
nor U25505 (N_25505,N_23837,N_23182);
xnor U25506 (N_25506,N_22648,N_22609);
and U25507 (N_25507,N_23941,N_22160);
nand U25508 (N_25508,N_22200,N_23045);
and U25509 (N_25509,N_22462,N_22182);
and U25510 (N_25510,N_23027,N_22243);
or U25511 (N_25511,N_23148,N_22407);
xnor U25512 (N_25512,N_22116,N_22374);
nor U25513 (N_25513,N_23032,N_23802);
nand U25514 (N_25514,N_22646,N_22778);
nor U25515 (N_25515,N_22161,N_23571);
xor U25516 (N_25516,N_23709,N_22091);
nor U25517 (N_25517,N_22457,N_22575);
nor U25518 (N_25518,N_23589,N_22475);
nand U25519 (N_25519,N_23400,N_23065);
nor U25520 (N_25520,N_23502,N_22688);
xnor U25521 (N_25521,N_23153,N_23182);
nand U25522 (N_25522,N_23930,N_22726);
and U25523 (N_25523,N_23199,N_22921);
nor U25524 (N_25524,N_23411,N_22146);
or U25525 (N_25525,N_23131,N_22274);
or U25526 (N_25526,N_23267,N_22221);
nor U25527 (N_25527,N_22075,N_22261);
nand U25528 (N_25528,N_23532,N_23291);
nand U25529 (N_25529,N_23876,N_22465);
and U25530 (N_25530,N_23654,N_23085);
and U25531 (N_25531,N_22398,N_22748);
xnor U25532 (N_25532,N_23316,N_22122);
or U25533 (N_25533,N_23260,N_23171);
nor U25534 (N_25534,N_22104,N_23193);
nand U25535 (N_25535,N_22749,N_23169);
xnor U25536 (N_25536,N_22496,N_22038);
nor U25537 (N_25537,N_22521,N_23893);
or U25538 (N_25538,N_22657,N_23211);
and U25539 (N_25539,N_23155,N_23661);
nand U25540 (N_25540,N_23483,N_22693);
nor U25541 (N_25541,N_22338,N_23514);
and U25542 (N_25542,N_22701,N_23524);
and U25543 (N_25543,N_23548,N_22837);
and U25544 (N_25544,N_23704,N_23864);
xnor U25545 (N_25545,N_22422,N_23715);
or U25546 (N_25546,N_23564,N_23522);
nor U25547 (N_25547,N_23378,N_22145);
xnor U25548 (N_25548,N_22913,N_23972);
or U25549 (N_25549,N_22156,N_22348);
xnor U25550 (N_25550,N_23237,N_22869);
nor U25551 (N_25551,N_23395,N_23384);
and U25552 (N_25552,N_23847,N_22437);
nor U25553 (N_25553,N_23561,N_22116);
and U25554 (N_25554,N_22159,N_22975);
nor U25555 (N_25555,N_23172,N_22927);
nor U25556 (N_25556,N_23412,N_23633);
and U25557 (N_25557,N_23120,N_23531);
or U25558 (N_25558,N_22734,N_22416);
xnor U25559 (N_25559,N_23093,N_23670);
xor U25560 (N_25560,N_23801,N_23240);
and U25561 (N_25561,N_22729,N_23153);
or U25562 (N_25562,N_22396,N_23016);
and U25563 (N_25563,N_23157,N_23413);
nor U25564 (N_25564,N_23423,N_22507);
or U25565 (N_25565,N_22976,N_23709);
nand U25566 (N_25566,N_22749,N_22952);
xor U25567 (N_25567,N_22889,N_22956);
xor U25568 (N_25568,N_22888,N_23512);
nor U25569 (N_25569,N_22195,N_23631);
and U25570 (N_25570,N_23417,N_23095);
xor U25571 (N_25571,N_23772,N_22493);
nand U25572 (N_25572,N_23394,N_22107);
or U25573 (N_25573,N_22355,N_22171);
and U25574 (N_25574,N_22419,N_23319);
nor U25575 (N_25575,N_22162,N_23636);
or U25576 (N_25576,N_22267,N_22886);
nand U25577 (N_25577,N_23715,N_22456);
nand U25578 (N_25578,N_23461,N_23995);
or U25579 (N_25579,N_23117,N_22131);
xor U25580 (N_25580,N_22574,N_23646);
or U25581 (N_25581,N_22134,N_22028);
nand U25582 (N_25582,N_22533,N_23240);
nand U25583 (N_25583,N_23361,N_23369);
and U25584 (N_25584,N_22023,N_22820);
or U25585 (N_25585,N_23864,N_23625);
and U25586 (N_25586,N_23314,N_22069);
xnor U25587 (N_25587,N_23928,N_22356);
or U25588 (N_25588,N_22438,N_22221);
nand U25589 (N_25589,N_22230,N_23074);
xnor U25590 (N_25590,N_23683,N_22179);
or U25591 (N_25591,N_22543,N_23284);
nand U25592 (N_25592,N_23072,N_22162);
or U25593 (N_25593,N_22825,N_23370);
or U25594 (N_25594,N_23774,N_23565);
or U25595 (N_25595,N_23030,N_23984);
and U25596 (N_25596,N_23896,N_23764);
and U25597 (N_25597,N_22238,N_22741);
nor U25598 (N_25598,N_22691,N_23250);
and U25599 (N_25599,N_22974,N_23917);
nor U25600 (N_25600,N_23131,N_23010);
nor U25601 (N_25601,N_23579,N_22471);
and U25602 (N_25602,N_23204,N_23262);
or U25603 (N_25603,N_22034,N_22721);
or U25604 (N_25604,N_23297,N_23058);
nor U25605 (N_25605,N_23006,N_22793);
or U25606 (N_25606,N_22976,N_22515);
or U25607 (N_25607,N_22636,N_22203);
or U25608 (N_25608,N_23697,N_23397);
nor U25609 (N_25609,N_22790,N_23645);
nor U25610 (N_25610,N_22201,N_22253);
nand U25611 (N_25611,N_23834,N_22634);
and U25612 (N_25612,N_23457,N_23615);
xnor U25613 (N_25613,N_23208,N_22292);
xor U25614 (N_25614,N_22684,N_22570);
and U25615 (N_25615,N_23584,N_22629);
xnor U25616 (N_25616,N_23264,N_22080);
or U25617 (N_25617,N_22839,N_22160);
or U25618 (N_25618,N_23168,N_23614);
or U25619 (N_25619,N_23524,N_22685);
nand U25620 (N_25620,N_22821,N_23805);
and U25621 (N_25621,N_22291,N_23610);
or U25622 (N_25622,N_22928,N_23330);
nand U25623 (N_25623,N_22722,N_22832);
and U25624 (N_25624,N_22858,N_22407);
nand U25625 (N_25625,N_23545,N_22888);
or U25626 (N_25626,N_23971,N_23311);
nand U25627 (N_25627,N_23011,N_22409);
and U25628 (N_25628,N_22173,N_22434);
or U25629 (N_25629,N_22786,N_22487);
nand U25630 (N_25630,N_23338,N_22492);
nor U25631 (N_25631,N_22138,N_22783);
nor U25632 (N_25632,N_22624,N_22007);
or U25633 (N_25633,N_22434,N_23189);
and U25634 (N_25634,N_22040,N_23962);
or U25635 (N_25635,N_22723,N_22325);
xnor U25636 (N_25636,N_23741,N_22881);
or U25637 (N_25637,N_23104,N_23622);
or U25638 (N_25638,N_22943,N_23885);
or U25639 (N_25639,N_22392,N_23688);
and U25640 (N_25640,N_22406,N_23691);
or U25641 (N_25641,N_22371,N_22310);
nor U25642 (N_25642,N_23458,N_22811);
nand U25643 (N_25643,N_22271,N_22161);
and U25644 (N_25644,N_23774,N_23820);
and U25645 (N_25645,N_23489,N_23650);
nand U25646 (N_25646,N_22007,N_23689);
or U25647 (N_25647,N_22699,N_22848);
nand U25648 (N_25648,N_22314,N_23380);
or U25649 (N_25649,N_22120,N_23297);
nor U25650 (N_25650,N_22490,N_22809);
and U25651 (N_25651,N_23765,N_23277);
nand U25652 (N_25652,N_22029,N_22560);
xnor U25653 (N_25653,N_23334,N_23043);
and U25654 (N_25654,N_22225,N_23502);
nand U25655 (N_25655,N_23982,N_23323);
nand U25656 (N_25656,N_22046,N_23674);
or U25657 (N_25657,N_23480,N_23959);
nor U25658 (N_25658,N_23810,N_22117);
nand U25659 (N_25659,N_23651,N_22070);
nor U25660 (N_25660,N_22393,N_22748);
nor U25661 (N_25661,N_22535,N_22728);
or U25662 (N_25662,N_22409,N_23731);
or U25663 (N_25663,N_22197,N_22520);
nor U25664 (N_25664,N_23008,N_22596);
and U25665 (N_25665,N_22150,N_23838);
and U25666 (N_25666,N_22361,N_23235);
and U25667 (N_25667,N_22451,N_23566);
nor U25668 (N_25668,N_22766,N_22429);
nor U25669 (N_25669,N_22481,N_22765);
or U25670 (N_25670,N_22062,N_22352);
nand U25671 (N_25671,N_23140,N_22503);
or U25672 (N_25672,N_22376,N_23535);
and U25673 (N_25673,N_23371,N_23080);
nand U25674 (N_25674,N_23538,N_22369);
and U25675 (N_25675,N_23522,N_23560);
nor U25676 (N_25676,N_23300,N_22910);
nand U25677 (N_25677,N_22462,N_23082);
and U25678 (N_25678,N_22097,N_23434);
nor U25679 (N_25679,N_22923,N_23622);
xnor U25680 (N_25680,N_23856,N_23618);
nand U25681 (N_25681,N_23773,N_22947);
and U25682 (N_25682,N_23737,N_23929);
and U25683 (N_25683,N_22895,N_22521);
or U25684 (N_25684,N_23094,N_22220);
nand U25685 (N_25685,N_22100,N_22710);
xor U25686 (N_25686,N_22259,N_22506);
xor U25687 (N_25687,N_23760,N_23036);
nand U25688 (N_25688,N_22261,N_22246);
nand U25689 (N_25689,N_22380,N_22580);
nand U25690 (N_25690,N_22831,N_22397);
nand U25691 (N_25691,N_23383,N_23283);
nand U25692 (N_25692,N_22628,N_23008);
xor U25693 (N_25693,N_23365,N_22666);
nand U25694 (N_25694,N_23323,N_23278);
and U25695 (N_25695,N_23803,N_23700);
and U25696 (N_25696,N_22943,N_22577);
xnor U25697 (N_25697,N_23769,N_23086);
and U25698 (N_25698,N_22408,N_23089);
nor U25699 (N_25699,N_23472,N_23517);
or U25700 (N_25700,N_22281,N_23759);
and U25701 (N_25701,N_23256,N_23319);
and U25702 (N_25702,N_23574,N_22391);
or U25703 (N_25703,N_22190,N_22591);
nor U25704 (N_25704,N_22874,N_22634);
nand U25705 (N_25705,N_23725,N_22891);
or U25706 (N_25706,N_22070,N_22845);
nand U25707 (N_25707,N_23947,N_22158);
or U25708 (N_25708,N_23311,N_22962);
and U25709 (N_25709,N_22278,N_22636);
or U25710 (N_25710,N_23869,N_22678);
and U25711 (N_25711,N_23700,N_22224);
nand U25712 (N_25712,N_23689,N_22906);
nand U25713 (N_25713,N_23527,N_23872);
or U25714 (N_25714,N_23733,N_23176);
or U25715 (N_25715,N_23604,N_23376);
nand U25716 (N_25716,N_23095,N_23035);
nand U25717 (N_25717,N_22705,N_23029);
and U25718 (N_25718,N_23159,N_22485);
or U25719 (N_25719,N_22415,N_22608);
nand U25720 (N_25720,N_23745,N_23758);
nor U25721 (N_25721,N_22999,N_22031);
xor U25722 (N_25722,N_23238,N_23093);
nand U25723 (N_25723,N_23330,N_23918);
or U25724 (N_25724,N_22402,N_23237);
xnor U25725 (N_25725,N_23551,N_23350);
xor U25726 (N_25726,N_22664,N_23957);
and U25727 (N_25727,N_23680,N_22043);
nand U25728 (N_25728,N_22352,N_23819);
nand U25729 (N_25729,N_22746,N_22017);
nor U25730 (N_25730,N_23090,N_22112);
and U25731 (N_25731,N_22083,N_23400);
and U25732 (N_25732,N_22365,N_23796);
and U25733 (N_25733,N_22610,N_23957);
xor U25734 (N_25734,N_23800,N_22202);
nor U25735 (N_25735,N_22507,N_22261);
xnor U25736 (N_25736,N_23444,N_22151);
xor U25737 (N_25737,N_22760,N_22517);
and U25738 (N_25738,N_22721,N_22728);
and U25739 (N_25739,N_22054,N_23074);
or U25740 (N_25740,N_23149,N_22166);
xnor U25741 (N_25741,N_22586,N_23117);
or U25742 (N_25742,N_22320,N_22035);
and U25743 (N_25743,N_23402,N_22230);
nand U25744 (N_25744,N_23398,N_22419);
or U25745 (N_25745,N_23662,N_22724);
and U25746 (N_25746,N_23789,N_22597);
and U25747 (N_25747,N_23651,N_22176);
and U25748 (N_25748,N_22929,N_22939);
xor U25749 (N_25749,N_22345,N_22966);
and U25750 (N_25750,N_23515,N_23901);
and U25751 (N_25751,N_23107,N_22231);
and U25752 (N_25752,N_22255,N_22910);
nand U25753 (N_25753,N_23656,N_23026);
nor U25754 (N_25754,N_22708,N_22515);
xor U25755 (N_25755,N_22358,N_22028);
xnor U25756 (N_25756,N_23043,N_22553);
nor U25757 (N_25757,N_22577,N_22285);
or U25758 (N_25758,N_22330,N_23333);
nand U25759 (N_25759,N_22301,N_23112);
or U25760 (N_25760,N_22941,N_23984);
nand U25761 (N_25761,N_23117,N_23471);
nor U25762 (N_25762,N_22063,N_22995);
and U25763 (N_25763,N_22238,N_23683);
nand U25764 (N_25764,N_23329,N_23242);
and U25765 (N_25765,N_22540,N_23968);
nand U25766 (N_25766,N_23999,N_22135);
and U25767 (N_25767,N_22043,N_23561);
xnor U25768 (N_25768,N_22499,N_23609);
nand U25769 (N_25769,N_23608,N_22370);
nor U25770 (N_25770,N_22387,N_23407);
xor U25771 (N_25771,N_22554,N_22185);
xor U25772 (N_25772,N_23942,N_22123);
or U25773 (N_25773,N_22454,N_23912);
and U25774 (N_25774,N_23640,N_23345);
and U25775 (N_25775,N_22004,N_23213);
or U25776 (N_25776,N_23428,N_22449);
xnor U25777 (N_25777,N_23395,N_22489);
xor U25778 (N_25778,N_22950,N_23029);
xnor U25779 (N_25779,N_23783,N_23160);
nand U25780 (N_25780,N_23756,N_23100);
nor U25781 (N_25781,N_23484,N_23966);
and U25782 (N_25782,N_23766,N_23659);
xnor U25783 (N_25783,N_23624,N_22097);
nand U25784 (N_25784,N_23122,N_23783);
and U25785 (N_25785,N_23584,N_23258);
or U25786 (N_25786,N_22587,N_22764);
or U25787 (N_25787,N_23059,N_23531);
or U25788 (N_25788,N_22627,N_22064);
or U25789 (N_25789,N_23126,N_23773);
nor U25790 (N_25790,N_22109,N_23655);
nand U25791 (N_25791,N_23339,N_22147);
or U25792 (N_25792,N_23549,N_23515);
or U25793 (N_25793,N_23329,N_22815);
nor U25794 (N_25794,N_22533,N_23417);
xor U25795 (N_25795,N_22413,N_22888);
and U25796 (N_25796,N_23210,N_22621);
or U25797 (N_25797,N_23724,N_22717);
and U25798 (N_25798,N_22366,N_22147);
nor U25799 (N_25799,N_22685,N_23235);
and U25800 (N_25800,N_23969,N_23486);
and U25801 (N_25801,N_22525,N_23401);
xor U25802 (N_25802,N_23410,N_22179);
xor U25803 (N_25803,N_23405,N_22792);
nand U25804 (N_25804,N_23925,N_23957);
or U25805 (N_25805,N_23544,N_23741);
xor U25806 (N_25806,N_23844,N_22090);
and U25807 (N_25807,N_23805,N_22763);
and U25808 (N_25808,N_23918,N_22442);
nor U25809 (N_25809,N_23781,N_23047);
and U25810 (N_25810,N_23714,N_22579);
and U25811 (N_25811,N_23662,N_22426);
nand U25812 (N_25812,N_22799,N_23359);
and U25813 (N_25813,N_22557,N_23136);
nor U25814 (N_25814,N_22493,N_23807);
or U25815 (N_25815,N_23270,N_22807);
nand U25816 (N_25816,N_22777,N_23693);
and U25817 (N_25817,N_22615,N_22617);
and U25818 (N_25818,N_22739,N_22076);
nor U25819 (N_25819,N_23665,N_23698);
nand U25820 (N_25820,N_23000,N_22131);
nor U25821 (N_25821,N_22550,N_23892);
and U25822 (N_25822,N_22363,N_23117);
nand U25823 (N_25823,N_23195,N_22767);
nor U25824 (N_25824,N_22421,N_22473);
nand U25825 (N_25825,N_23310,N_23952);
xnor U25826 (N_25826,N_23925,N_23360);
nand U25827 (N_25827,N_22174,N_23084);
and U25828 (N_25828,N_23611,N_22363);
or U25829 (N_25829,N_22963,N_23095);
or U25830 (N_25830,N_22141,N_22970);
xor U25831 (N_25831,N_23867,N_22278);
nand U25832 (N_25832,N_23942,N_23525);
nor U25833 (N_25833,N_22115,N_23516);
and U25834 (N_25834,N_23783,N_22158);
xnor U25835 (N_25835,N_23519,N_23491);
and U25836 (N_25836,N_22557,N_22593);
xnor U25837 (N_25837,N_23082,N_23115);
nand U25838 (N_25838,N_23110,N_23919);
nor U25839 (N_25839,N_23541,N_22540);
nand U25840 (N_25840,N_22515,N_23651);
and U25841 (N_25841,N_23293,N_23638);
xnor U25842 (N_25842,N_22067,N_22143);
or U25843 (N_25843,N_23409,N_22572);
and U25844 (N_25844,N_23737,N_22813);
xnor U25845 (N_25845,N_22225,N_22682);
and U25846 (N_25846,N_23725,N_22919);
and U25847 (N_25847,N_22358,N_22554);
xnor U25848 (N_25848,N_22163,N_23780);
nor U25849 (N_25849,N_22433,N_23133);
nand U25850 (N_25850,N_22265,N_22787);
and U25851 (N_25851,N_23474,N_23566);
xnor U25852 (N_25852,N_22079,N_22308);
or U25853 (N_25853,N_22366,N_22542);
nor U25854 (N_25854,N_22952,N_22869);
nor U25855 (N_25855,N_22280,N_23622);
or U25856 (N_25856,N_23761,N_22103);
xor U25857 (N_25857,N_22612,N_22850);
xor U25858 (N_25858,N_23799,N_23701);
nor U25859 (N_25859,N_23765,N_22086);
nand U25860 (N_25860,N_22320,N_22687);
nor U25861 (N_25861,N_22789,N_22493);
xor U25862 (N_25862,N_22632,N_23964);
and U25863 (N_25863,N_23469,N_22886);
nand U25864 (N_25864,N_22029,N_22552);
nor U25865 (N_25865,N_22957,N_22346);
and U25866 (N_25866,N_22611,N_22688);
nand U25867 (N_25867,N_23687,N_22944);
nand U25868 (N_25868,N_22154,N_22591);
nor U25869 (N_25869,N_23067,N_22811);
nand U25870 (N_25870,N_22599,N_23743);
nor U25871 (N_25871,N_23047,N_22310);
and U25872 (N_25872,N_22469,N_23917);
xor U25873 (N_25873,N_22016,N_23142);
nand U25874 (N_25874,N_22466,N_22503);
nor U25875 (N_25875,N_23220,N_23017);
nor U25876 (N_25876,N_22617,N_23569);
xor U25877 (N_25877,N_23467,N_22444);
or U25878 (N_25878,N_23318,N_23118);
nor U25879 (N_25879,N_23225,N_23805);
nand U25880 (N_25880,N_23973,N_22688);
nand U25881 (N_25881,N_22929,N_22715);
nor U25882 (N_25882,N_23629,N_22576);
xnor U25883 (N_25883,N_22788,N_23227);
and U25884 (N_25884,N_22349,N_23800);
or U25885 (N_25885,N_23304,N_23666);
or U25886 (N_25886,N_22361,N_22450);
or U25887 (N_25887,N_23163,N_23314);
nand U25888 (N_25888,N_22428,N_23933);
nand U25889 (N_25889,N_23430,N_23028);
xnor U25890 (N_25890,N_23968,N_23349);
and U25891 (N_25891,N_22795,N_23068);
xnor U25892 (N_25892,N_23788,N_22873);
nand U25893 (N_25893,N_22308,N_23352);
and U25894 (N_25894,N_23651,N_23304);
and U25895 (N_25895,N_22856,N_22965);
xor U25896 (N_25896,N_23749,N_23475);
or U25897 (N_25897,N_23213,N_22907);
nand U25898 (N_25898,N_23561,N_22755);
nor U25899 (N_25899,N_23546,N_23913);
nand U25900 (N_25900,N_23211,N_22772);
nand U25901 (N_25901,N_22689,N_23012);
xnor U25902 (N_25902,N_22435,N_23632);
xor U25903 (N_25903,N_22052,N_22062);
or U25904 (N_25904,N_22260,N_23198);
nand U25905 (N_25905,N_23943,N_22985);
and U25906 (N_25906,N_23308,N_22587);
or U25907 (N_25907,N_23047,N_23200);
and U25908 (N_25908,N_22099,N_23932);
xnor U25909 (N_25909,N_23913,N_22067);
or U25910 (N_25910,N_23353,N_23392);
and U25911 (N_25911,N_22835,N_22138);
xor U25912 (N_25912,N_23659,N_23775);
nand U25913 (N_25913,N_22500,N_22832);
or U25914 (N_25914,N_22314,N_23010);
or U25915 (N_25915,N_23448,N_23034);
nand U25916 (N_25916,N_23989,N_22179);
or U25917 (N_25917,N_22669,N_22430);
and U25918 (N_25918,N_23660,N_23748);
nand U25919 (N_25919,N_22096,N_23635);
nand U25920 (N_25920,N_23716,N_23600);
nor U25921 (N_25921,N_22279,N_23070);
or U25922 (N_25922,N_22595,N_23717);
nand U25923 (N_25923,N_23496,N_22438);
nand U25924 (N_25924,N_23503,N_22265);
or U25925 (N_25925,N_22179,N_22975);
nor U25926 (N_25926,N_22053,N_23190);
or U25927 (N_25927,N_22269,N_22589);
nor U25928 (N_25928,N_22405,N_23264);
or U25929 (N_25929,N_22159,N_22815);
nor U25930 (N_25930,N_23165,N_22280);
nand U25931 (N_25931,N_23624,N_22284);
or U25932 (N_25932,N_22371,N_22077);
and U25933 (N_25933,N_22858,N_22824);
nor U25934 (N_25934,N_23074,N_23564);
and U25935 (N_25935,N_23645,N_23955);
or U25936 (N_25936,N_22410,N_23500);
and U25937 (N_25937,N_23028,N_22062);
or U25938 (N_25938,N_22545,N_23352);
or U25939 (N_25939,N_23071,N_23761);
xor U25940 (N_25940,N_23131,N_23099);
xnor U25941 (N_25941,N_23831,N_23814);
and U25942 (N_25942,N_23782,N_22209);
nor U25943 (N_25943,N_23181,N_23921);
nand U25944 (N_25944,N_22691,N_23187);
xor U25945 (N_25945,N_22473,N_22166);
or U25946 (N_25946,N_23883,N_23583);
xnor U25947 (N_25947,N_23405,N_22380);
and U25948 (N_25948,N_22482,N_22377);
xnor U25949 (N_25949,N_23284,N_23130);
nor U25950 (N_25950,N_23659,N_23924);
or U25951 (N_25951,N_22914,N_23651);
xnor U25952 (N_25952,N_22432,N_22600);
nand U25953 (N_25953,N_22963,N_22359);
and U25954 (N_25954,N_23327,N_23751);
nor U25955 (N_25955,N_23768,N_22940);
nor U25956 (N_25956,N_23251,N_22570);
or U25957 (N_25957,N_23398,N_22892);
and U25958 (N_25958,N_23811,N_22740);
nand U25959 (N_25959,N_22359,N_23297);
xnor U25960 (N_25960,N_22184,N_23922);
or U25961 (N_25961,N_22643,N_22927);
nand U25962 (N_25962,N_22555,N_23037);
nor U25963 (N_25963,N_22754,N_22173);
nor U25964 (N_25964,N_22195,N_23393);
or U25965 (N_25965,N_22064,N_22511);
and U25966 (N_25966,N_22903,N_23467);
or U25967 (N_25967,N_23615,N_23378);
xnor U25968 (N_25968,N_22688,N_22294);
nor U25969 (N_25969,N_23928,N_22651);
nor U25970 (N_25970,N_22290,N_23686);
xnor U25971 (N_25971,N_23074,N_23387);
and U25972 (N_25972,N_22402,N_22838);
and U25973 (N_25973,N_22786,N_23246);
nand U25974 (N_25974,N_22430,N_23894);
and U25975 (N_25975,N_23879,N_22462);
xor U25976 (N_25976,N_22079,N_23802);
or U25977 (N_25977,N_23420,N_23768);
and U25978 (N_25978,N_23102,N_22126);
and U25979 (N_25979,N_22280,N_23434);
or U25980 (N_25980,N_22191,N_22086);
and U25981 (N_25981,N_22969,N_22167);
or U25982 (N_25982,N_22765,N_22529);
xor U25983 (N_25983,N_23088,N_22634);
or U25984 (N_25984,N_23917,N_23364);
nand U25985 (N_25985,N_23701,N_23444);
or U25986 (N_25986,N_22122,N_23999);
nor U25987 (N_25987,N_23341,N_23809);
nor U25988 (N_25988,N_23076,N_22678);
or U25989 (N_25989,N_23958,N_22869);
or U25990 (N_25990,N_23114,N_22338);
or U25991 (N_25991,N_23088,N_22861);
nand U25992 (N_25992,N_22886,N_23407);
xor U25993 (N_25993,N_22962,N_22820);
and U25994 (N_25994,N_22272,N_23047);
or U25995 (N_25995,N_22477,N_22203);
nor U25996 (N_25996,N_23414,N_23931);
and U25997 (N_25997,N_22679,N_22471);
or U25998 (N_25998,N_23960,N_23480);
xor U25999 (N_25999,N_22940,N_23151);
xor U26000 (N_26000,N_24102,N_25904);
xor U26001 (N_26001,N_24128,N_24124);
xnor U26002 (N_26002,N_25137,N_24225);
xnor U26003 (N_26003,N_24652,N_24272);
nor U26004 (N_26004,N_24570,N_25639);
nor U26005 (N_26005,N_24065,N_25252);
and U26006 (N_26006,N_24839,N_25077);
xor U26007 (N_26007,N_25426,N_24253);
nand U26008 (N_26008,N_24997,N_24478);
nand U26009 (N_26009,N_25795,N_25185);
and U26010 (N_26010,N_25199,N_25523);
nor U26011 (N_26011,N_25746,N_24567);
xor U26012 (N_26012,N_25057,N_25111);
nand U26013 (N_26013,N_24313,N_24336);
nand U26014 (N_26014,N_25240,N_25178);
xor U26015 (N_26015,N_25419,N_25549);
xor U26016 (N_26016,N_24142,N_24176);
nor U26017 (N_26017,N_25263,N_24003);
or U26018 (N_26018,N_24943,N_24671);
and U26019 (N_26019,N_25308,N_24091);
xor U26020 (N_26020,N_24936,N_24180);
nand U26021 (N_26021,N_24677,N_25075);
nor U26022 (N_26022,N_24165,N_25021);
and U26023 (N_26023,N_24487,N_24910);
nor U26024 (N_26024,N_25382,N_25787);
and U26025 (N_26025,N_24799,N_25157);
and U26026 (N_26026,N_24739,N_25964);
and U26027 (N_26027,N_24971,N_25878);
and U26028 (N_26028,N_24451,N_24236);
and U26029 (N_26029,N_24851,N_25899);
or U26030 (N_26030,N_25464,N_25242);
or U26031 (N_26031,N_25329,N_24160);
and U26032 (N_26032,N_25020,N_25003);
or U26033 (N_26033,N_25640,N_24070);
nand U26034 (N_26034,N_25414,N_25445);
and U26035 (N_26035,N_24712,N_25209);
xnor U26036 (N_26036,N_24682,N_24257);
xnor U26037 (N_26037,N_24542,N_24561);
nor U26038 (N_26038,N_25771,N_25732);
and U26039 (N_26039,N_25365,N_24885);
nor U26040 (N_26040,N_25337,N_24442);
or U26041 (N_26041,N_25662,N_25811);
or U26042 (N_26042,N_25692,N_25429);
and U26043 (N_26043,N_24945,N_25074);
and U26044 (N_26044,N_24144,N_24310);
and U26045 (N_26045,N_24378,N_24098);
nand U26046 (N_26046,N_24828,N_24927);
or U26047 (N_26047,N_24007,N_24448);
xor U26048 (N_26048,N_25257,N_25764);
nand U26049 (N_26049,N_24551,N_24982);
xnor U26050 (N_26050,N_25092,N_24486);
nand U26051 (N_26051,N_25495,N_24089);
nor U26052 (N_26052,N_25600,N_25163);
xnor U26053 (N_26053,N_25475,N_24887);
nor U26054 (N_26054,N_24625,N_24443);
xor U26055 (N_26055,N_24299,N_24857);
or U26056 (N_26056,N_25520,N_25061);
xor U26057 (N_26057,N_24428,N_24988);
nand U26058 (N_26058,N_24362,N_24341);
and U26059 (N_26059,N_24019,N_25581);
or U26060 (N_26060,N_24800,N_25428);
and U26061 (N_26061,N_25601,N_25848);
or U26062 (N_26062,N_24740,N_25224);
nor U26063 (N_26063,N_25299,N_25897);
and U26064 (N_26064,N_24447,N_25786);
nand U26065 (N_26065,N_24632,N_25970);
nor U26066 (N_26066,N_25915,N_25181);
or U26067 (N_26067,N_25867,N_25238);
nor U26068 (N_26068,N_24889,N_24888);
xor U26069 (N_26069,N_24500,N_25589);
and U26070 (N_26070,N_25922,N_24370);
nor U26071 (N_26071,N_25695,N_25822);
or U26072 (N_26072,N_25369,N_24396);
xor U26073 (N_26073,N_25876,N_25352);
and U26074 (N_26074,N_25696,N_24169);
and U26075 (N_26075,N_24177,N_25576);
nand U26076 (N_26076,N_24568,N_25836);
or U26077 (N_26077,N_24059,N_25345);
nor U26078 (N_26078,N_25260,N_24516);
and U26079 (N_26079,N_24733,N_24001);
or U26080 (N_26080,N_25540,N_25205);
nor U26081 (N_26081,N_25743,N_24806);
nand U26082 (N_26082,N_24491,N_25951);
or U26083 (N_26083,N_24154,N_25854);
or U26084 (N_26084,N_24690,N_25927);
nor U26085 (N_26085,N_24414,N_24787);
nand U26086 (N_26086,N_24620,N_25239);
and U26087 (N_26087,N_25539,N_24217);
and U26088 (N_26088,N_25585,N_25504);
xor U26089 (N_26089,N_25104,N_25816);
nor U26090 (N_26090,N_25674,N_24520);
or U26091 (N_26091,N_25071,N_24657);
or U26092 (N_26092,N_25596,N_25525);
xor U26093 (N_26093,N_25268,N_24139);
nand U26094 (N_26094,N_25647,N_24467);
xnor U26095 (N_26095,N_24668,N_24832);
or U26096 (N_26096,N_24840,N_25318);
nand U26097 (N_26097,N_24711,N_25992);
xor U26098 (N_26098,N_25358,N_25877);
xnor U26099 (N_26099,N_24347,N_24864);
or U26100 (N_26100,N_25605,N_24320);
nand U26101 (N_26101,N_24902,N_25142);
nor U26102 (N_26102,N_25655,N_24265);
or U26103 (N_26103,N_24781,N_24494);
xnor U26104 (N_26104,N_24614,N_24726);
or U26105 (N_26105,N_24539,N_24928);
nand U26106 (N_26106,N_24084,N_25166);
or U26107 (N_26107,N_24793,N_24323);
xor U26108 (N_26108,N_25776,N_24817);
xor U26109 (N_26109,N_24786,N_25863);
nor U26110 (N_26110,N_24771,N_25254);
nand U26111 (N_26111,N_24528,N_25672);
and U26112 (N_26112,N_25582,N_25486);
xor U26113 (N_26113,N_25131,N_24940);
xor U26114 (N_26114,N_25511,N_25593);
nor U26115 (N_26115,N_25431,N_25411);
nor U26116 (N_26116,N_25135,N_25757);
xor U26117 (N_26117,N_24496,N_24464);
nand U26118 (N_26118,N_25261,N_24314);
and U26119 (N_26119,N_24201,N_25957);
xnor U26120 (N_26120,N_25241,N_24812);
and U26121 (N_26121,N_25779,N_24758);
nor U26122 (N_26122,N_24004,N_24530);
nand U26123 (N_26123,N_25105,N_25643);
nor U26124 (N_26124,N_24452,N_25530);
or U26125 (N_26125,N_24942,N_25499);
nor U26126 (N_26126,N_24855,N_25186);
and U26127 (N_26127,N_25890,N_25212);
or U26128 (N_26128,N_25911,N_24078);
and U26129 (N_26129,N_25841,N_25051);
or U26130 (N_26130,N_24660,N_24244);
nand U26131 (N_26131,N_24510,N_25860);
or U26132 (N_26132,N_24006,N_24643);
or U26133 (N_26133,N_24790,N_24183);
nor U26134 (N_26134,N_25620,N_24878);
xor U26135 (N_26135,N_25487,N_25637);
and U26136 (N_26136,N_24756,N_25862);
or U26137 (N_26137,N_24205,N_25085);
and U26138 (N_26138,N_25140,N_24699);
or U26139 (N_26139,N_24986,N_24387);
and U26140 (N_26140,N_24120,N_25264);
nor U26141 (N_26141,N_24178,N_24663);
xnor U26142 (N_26142,N_24095,N_25990);
xor U26143 (N_26143,N_24251,N_24619);
xnor U26144 (N_26144,N_24955,N_24805);
and U26145 (N_26145,N_25128,N_25782);
or U26146 (N_26146,N_24705,N_24723);
xor U26147 (N_26147,N_24952,N_25281);
and U26148 (N_26148,N_25235,N_25792);
and U26149 (N_26149,N_24852,N_25587);
or U26150 (N_26150,N_24794,N_25227);
xor U26151 (N_26151,N_25680,N_24750);
or U26152 (N_26152,N_25461,N_24288);
xor U26153 (N_26153,N_24992,N_25468);
xnor U26154 (N_26154,N_24164,N_24687);
nor U26155 (N_26155,N_25283,N_25229);
xnor U26156 (N_26156,N_25024,N_24416);
xor U26157 (N_26157,N_25619,N_25577);
xor U26158 (N_26158,N_24117,N_25706);
and U26159 (N_26159,N_24363,N_24572);
or U26160 (N_26160,N_25032,N_25328);
xor U26161 (N_26161,N_24025,N_25825);
nand U26162 (N_26162,N_24290,N_24100);
xnor U26163 (N_26163,N_24718,N_24651);
nor U26164 (N_26164,N_25673,N_24669);
and U26165 (N_26165,N_24135,N_25381);
nand U26166 (N_26166,N_25002,N_25538);
or U26167 (N_26167,N_24770,N_24961);
nand U26168 (N_26168,N_25125,N_24335);
or U26169 (N_26169,N_24742,N_25439);
nor U26170 (N_26170,N_24247,N_25819);
and U26171 (N_26171,N_25331,N_25519);
nor U26172 (N_26172,N_25107,N_24188);
nor U26173 (N_26173,N_24905,N_25987);
or U26174 (N_26174,N_24819,N_24939);
xor U26175 (N_26175,N_24576,N_25083);
xnor U26176 (N_26176,N_24404,N_25847);
nand U26177 (N_26177,N_24693,N_24147);
xor U26178 (N_26178,N_25873,N_25798);
xnor U26179 (N_26179,N_24399,N_25668);
nor U26180 (N_26180,N_25670,N_25768);
xor U26181 (N_26181,N_25944,N_24836);
nand U26182 (N_26182,N_24623,N_24175);
or U26183 (N_26183,N_24611,N_25516);
or U26184 (N_26184,N_25366,N_25386);
nor U26185 (N_26185,N_24874,N_25949);
nand U26186 (N_26186,N_25820,N_24366);
nor U26187 (N_26187,N_25962,N_24951);
xor U26188 (N_26188,N_24460,N_25517);
nor U26189 (N_26189,N_25451,N_24903);
or U26190 (N_26190,N_24907,N_24655);
or U26191 (N_26191,N_25629,N_25658);
and U26192 (N_26192,N_24810,N_24618);
nor U26193 (N_26193,N_25344,N_25245);
nor U26194 (N_26194,N_25467,N_24064);
and U26195 (N_26195,N_25286,N_25446);
xor U26196 (N_26196,N_25543,N_25558);
xnor U26197 (N_26197,N_24246,N_24985);
nand U26198 (N_26198,N_24929,N_25682);
nor U26199 (N_26199,N_25925,N_24999);
and U26200 (N_26200,N_24316,N_25720);
or U26201 (N_26201,N_24615,N_25697);
nand U26202 (N_26202,N_24104,N_25652);
nand U26203 (N_26203,N_25374,N_25007);
xor U26204 (N_26204,N_25404,N_25684);
nor U26205 (N_26205,N_25055,N_24697);
xnor U26206 (N_26206,N_25733,N_24213);
and U26207 (N_26207,N_24987,N_24196);
or U26208 (N_26208,N_24879,N_25972);
and U26209 (N_26209,N_25592,N_25127);
and U26210 (N_26210,N_25955,N_25430);
and U26211 (N_26211,N_24191,N_25183);
and U26212 (N_26212,N_24681,N_25282);
and U26213 (N_26213,N_24161,N_25714);
nand U26214 (N_26214,N_25929,N_25579);
or U26215 (N_26215,N_24538,N_24242);
nor U26216 (N_26216,N_25572,N_25853);
xnor U26217 (N_26217,N_25718,N_25053);
and U26218 (N_26218,N_24710,N_24368);
and U26219 (N_26219,N_25722,N_24882);
nor U26220 (N_26220,N_25028,N_24604);
nor U26221 (N_26221,N_25029,N_25700);
nand U26222 (N_26222,N_25500,N_25698);
and U26223 (N_26223,N_25588,N_25801);
nor U26224 (N_26224,N_25785,N_25638);
xor U26225 (N_26225,N_24748,N_25541);
nand U26226 (N_26226,N_25594,N_25703);
nor U26227 (N_26227,N_24360,N_25044);
xor U26228 (N_26228,N_24862,N_24186);
and U26229 (N_26229,N_24397,N_25158);
xnor U26230 (N_26230,N_24359,N_24248);
or U26231 (N_26231,N_25918,N_24014);
xor U26232 (N_26232,N_25221,N_24689);
nor U26233 (N_26233,N_24113,N_24779);
or U26234 (N_26234,N_25995,N_24593);
or U26235 (N_26235,N_25067,N_24010);
or U26236 (N_26236,N_25300,N_24297);
nor U26237 (N_26237,N_24484,N_24527);
nor U26238 (N_26238,N_25512,N_24085);
or U26239 (N_26239,N_25646,N_25472);
nand U26240 (N_26240,N_25206,N_25749);
xnor U26241 (N_26241,N_24371,N_25406);
nor U26242 (N_26242,N_24934,N_24911);
nor U26243 (N_26243,N_25770,N_24277);
and U26244 (N_26244,N_24476,N_24002);
and U26245 (N_26245,N_24340,N_25121);
nand U26246 (N_26246,N_25409,N_25452);
or U26247 (N_26247,N_25740,N_25350);
nand U26248 (N_26248,N_24173,N_24018);
nor U26249 (N_26249,N_25978,N_24743);
nand U26250 (N_26250,N_24716,N_24591);
xnor U26251 (N_26251,N_25815,N_24958);
nand U26252 (N_26252,N_25326,N_24184);
xor U26253 (N_26253,N_24410,N_25171);
nor U26254 (N_26254,N_25490,N_24262);
nor U26255 (N_26255,N_25980,N_24369);
xor U26256 (N_26256,N_25156,N_24055);
or U26257 (N_26257,N_24092,N_24259);
xnor U26258 (N_26258,N_25433,N_24264);
or U26259 (N_26259,N_25296,N_24497);
nand U26260 (N_26260,N_24269,N_25947);
and U26261 (N_26261,N_24645,N_24079);
nor U26262 (N_26262,N_24924,N_24588);
nand U26263 (N_26263,N_25902,N_24458);
xnor U26264 (N_26264,N_24168,N_24913);
nand U26265 (N_26265,N_24093,N_24768);
xor U26266 (N_26266,N_25561,N_25072);
or U26267 (N_26267,N_25315,N_24504);
xor U26268 (N_26268,N_25859,N_24848);
nand U26269 (N_26269,N_24675,N_25159);
xor U26270 (N_26270,N_25755,N_24330);
xor U26271 (N_26271,N_25336,N_25609);
and U26272 (N_26272,N_24754,N_25542);
or U26273 (N_26273,N_24221,N_25138);
nand U26274 (N_26274,N_24532,N_25086);
xnor U26275 (N_26275,N_25050,N_25591);
nand U26276 (N_26276,N_25810,N_24067);
nand U26277 (N_26277,N_24577,N_24881);
xor U26278 (N_26278,N_25642,N_25388);
and U26279 (N_26279,N_25341,N_25800);
and U26280 (N_26280,N_25334,N_24134);
nand U26281 (N_26281,N_24233,N_24445);
and U26282 (N_26282,N_24775,N_25040);
nand U26283 (N_26283,N_24920,N_25378);
nor U26284 (N_26284,N_25338,N_24495);
xnor U26285 (N_26285,N_24899,N_25496);
nor U26286 (N_26286,N_25685,N_25113);
xor U26287 (N_26287,N_25317,N_24569);
and U26288 (N_26288,N_24607,N_24110);
or U26289 (N_26289,N_25501,N_24630);
xor U26290 (N_26290,N_24937,N_25146);
and U26291 (N_26291,N_25396,N_24275);
and U26292 (N_26292,N_24082,N_25834);
and U26293 (N_26293,N_24040,N_24015);
or U26294 (N_26294,N_24385,N_25874);
or U26295 (N_26295,N_25442,N_24769);
or U26296 (N_26296,N_25249,N_24749);
or U26297 (N_26297,N_25139,N_24146);
and U26298 (N_26298,N_24586,N_25748);
or U26299 (N_26299,N_25780,N_24271);
and U26300 (N_26300,N_24738,N_24389);
xnor U26301 (N_26301,N_24865,N_25560);
nor U26302 (N_26302,N_25923,N_24580);
nand U26303 (N_26303,N_24140,N_25744);
and U26304 (N_26304,N_24274,N_25194);
nor U26305 (N_26305,N_24054,N_25935);
or U26306 (N_26306,N_24112,N_25364);
nand U26307 (N_26307,N_24296,N_25371);
and U26308 (N_26308,N_25228,N_25099);
nand U26309 (N_26309,N_25025,N_24254);
or U26310 (N_26310,N_24890,N_25231);
or U26311 (N_26311,N_25750,N_24240);
nor U26312 (N_26312,N_25351,N_24755);
xor U26313 (N_26313,N_25034,N_25650);
and U26314 (N_26314,N_25781,N_24052);
or U26315 (N_26315,N_24692,N_25043);
or U26316 (N_26316,N_25457,N_25705);
nand U26317 (N_26317,N_24706,N_25598);
nand U26318 (N_26318,N_25958,N_25463);
nand U26319 (N_26319,N_25310,N_24212);
nor U26320 (N_26320,N_25389,N_25546);
nand U26321 (N_26321,N_24933,N_25444);
or U26322 (N_26322,N_25656,N_24801);
nor U26323 (N_26323,N_24617,N_25006);
nand U26324 (N_26324,N_24959,N_24229);
nand U26325 (N_26325,N_25115,N_25711);
nand U26326 (N_26326,N_25023,N_24980);
and U26327 (N_26327,N_25521,N_24342);
nand U26328 (N_26328,N_25522,N_24115);
or U26329 (N_26329,N_24114,N_25362);
nand U26330 (N_26330,N_25702,N_25886);
nor U26331 (N_26331,N_25660,N_25928);
and U26332 (N_26332,N_25736,N_25109);
xor U26333 (N_26333,N_25954,N_24914);
or U26334 (N_26334,N_25934,N_24037);
or U26335 (N_26335,N_25041,N_24796);
or U26336 (N_26336,N_25207,N_25564);
or U26337 (N_26337,N_25208,N_25909);
and U26338 (N_26338,N_25665,N_24908);
nand U26339 (N_26339,N_25160,N_25996);
xnor U26340 (N_26340,N_24305,N_25731);
xor U26341 (N_26341,N_24960,N_25030);
nand U26342 (N_26342,N_24734,N_25641);
or U26343 (N_26343,N_24802,N_24393);
or U26344 (N_26344,N_25399,N_24373);
and U26345 (N_26345,N_25628,N_25611);
nor U26346 (N_26346,N_24546,N_25590);
nand U26347 (N_26347,N_25998,N_24485);
or U26348 (N_26348,N_25751,N_24715);
or U26349 (N_26349,N_24919,N_24667);
and U26350 (N_26350,N_24422,N_25797);
nor U26351 (N_26351,N_24856,N_24127);
and U26352 (N_26352,N_24587,N_25844);
nand U26353 (N_26353,N_24838,N_25271);
nor U26354 (N_26354,N_24735,N_24076);
or U26355 (N_26355,N_24818,N_25091);
nor U26356 (N_26356,N_25884,N_24599);
or U26357 (N_26357,N_24600,N_25676);
nor U26358 (N_26358,N_24461,N_24954);
or U26359 (N_26359,N_25942,N_25881);
xor U26360 (N_26360,N_24099,N_24598);
and U26361 (N_26361,N_25737,N_25031);
and U26362 (N_26362,N_24167,N_24249);
or U26363 (N_26363,N_24270,N_25566);
nand U26364 (N_26364,N_24592,N_24821);
nor U26365 (N_26365,N_24732,N_25190);
nand U26366 (N_26366,N_24867,N_25427);
nor U26367 (N_26367,N_25574,N_24590);
nand U26368 (N_26368,N_24087,N_25627);
and U26369 (N_26369,N_24814,N_25154);
or U26370 (N_26370,N_24398,N_25545);
nor U26371 (N_26371,N_24747,N_25173);
nor U26372 (N_26372,N_25307,N_24627);
nor U26373 (N_26373,N_24302,N_24798);
xnor U26374 (N_26374,N_25112,N_24631);
nand U26375 (N_26375,N_24647,N_24823);
nor U26376 (N_26376,N_24068,N_24379);
xor U26377 (N_26377,N_24629,N_24023);
or U26378 (N_26378,N_24352,N_25037);
xnor U26379 (N_26379,N_25165,N_25959);
nor U26380 (N_26380,N_25060,N_25269);
nand U26381 (N_26381,N_25394,N_24382);
nor U26382 (N_26382,N_24553,N_24543);
and U26383 (N_26383,N_25355,N_25657);
or U26384 (N_26384,N_25952,N_24315);
nor U26385 (N_26385,N_25387,N_24766);
and U26386 (N_26386,N_25237,N_24941);
and U26387 (N_26387,N_24195,N_25913);
nor U26388 (N_26388,N_24597,N_24778);
and U26389 (N_26389,N_24343,N_24462);
nand U26390 (N_26390,N_25681,N_25480);
nand U26391 (N_26391,N_24189,N_24482);
xor U26392 (N_26392,N_25536,N_24883);
or U26393 (N_26393,N_25989,N_25636);
nor U26394 (N_26394,N_24993,N_24412);
nor U26395 (N_26395,N_24143,N_24956);
or U26396 (N_26396,N_25289,N_25195);
or U26397 (N_26397,N_24622,N_25089);
xor U26398 (N_26398,N_24376,N_24815);
nor U26399 (N_26399,N_25827,N_25912);
nand U26400 (N_26400,N_24536,N_24944);
nor U26401 (N_26401,N_25994,N_24489);
or U26402 (N_26402,N_25547,N_24822);
xnor U26403 (N_26403,N_25460,N_25484);
xor U26404 (N_26404,N_25405,N_24900);
and U26405 (N_26405,N_24638,N_24050);
xor U26406 (N_26406,N_25979,N_24132);
nand U26407 (N_26407,N_25941,N_25494);
or U26408 (N_26408,N_24268,N_25174);
nor U26409 (N_26409,N_25568,N_24153);
nand U26410 (N_26410,N_24051,N_24273);
nor U26411 (N_26411,N_25274,N_24833);
nor U26412 (N_26412,N_24250,N_25901);
or U26413 (N_26413,N_24728,N_25356);
or U26414 (N_26414,N_25882,N_25313);
xor U26415 (N_26415,N_24921,N_24721);
or U26416 (N_26416,N_24071,N_24408);
xor U26417 (N_26417,N_24654,N_25491);
xor U26418 (N_26418,N_24574,N_24130);
and U26419 (N_26419,N_24190,N_24602);
xnor U26420 (N_26420,N_25891,N_25838);
nand U26421 (N_26421,N_24608,N_24306);
or U26422 (N_26422,N_25965,N_24309);
nand U26423 (N_26423,N_25664,N_24585);
xor U26424 (N_26424,N_25624,N_24395);
nor U26425 (N_26425,N_25288,N_24056);
nand U26426 (N_26426,N_24245,N_25895);
or U26427 (N_26427,N_25384,N_24372);
nand U26428 (N_26428,N_24166,N_25839);
xnor U26429 (N_26429,N_25790,N_25689);
nor U26430 (N_26430,N_25514,N_25136);
or U26431 (N_26431,N_24641,N_25869);
and U26432 (N_26432,N_25508,N_25435);
nor U26433 (N_26433,N_24694,N_24519);
nand U26434 (N_26434,N_24328,N_25339);
or U26435 (N_26435,N_24116,N_24024);
nand U26436 (N_26436,N_25470,N_24243);
xor U26437 (N_26437,N_25395,N_24226);
and U26438 (N_26438,N_24884,N_25936);
nor U26439 (N_26439,N_25218,N_24463);
nor U26440 (N_26440,N_25971,N_24179);
or U26441 (N_26441,N_24891,N_25728);
nor U26442 (N_26442,N_25907,N_24946);
or U26443 (N_26443,N_24503,N_25476);
or U26444 (N_26444,N_25407,N_24628);
nand U26445 (N_26445,N_25210,N_25082);
nand U26446 (N_26446,N_25130,N_24736);
xor U26447 (N_26447,N_24034,N_25932);
nor U26448 (N_26448,N_25222,N_25571);
and U26449 (N_26449,N_25778,N_25986);
nor U26450 (N_26450,N_25462,N_25230);
nor U26451 (N_26451,N_24918,N_24912);
nor U26452 (N_26452,N_25898,N_25946);
nand U26453 (N_26453,N_25554,N_24234);
nor U26454 (N_26454,N_25035,N_25379);
nor U26455 (N_26455,N_24744,N_24774);
nand U26456 (N_26456,N_25709,N_24998);
nand U26457 (N_26457,N_25976,N_25595);
or U26458 (N_26458,N_25280,N_25515);
or U26459 (N_26459,N_25769,N_24198);
xor U26460 (N_26460,N_24375,N_25567);
or U26461 (N_26461,N_25416,N_25048);
nand U26462 (N_26462,N_24820,N_24957);
xnor U26463 (N_26463,N_25919,N_25621);
or U26464 (N_26464,N_24119,N_25065);
or U26465 (N_26465,N_25708,N_24322);
xor U26466 (N_26466,N_24702,N_24696);
or U26467 (N_26467,N_25380,N_24214);
nor U26468 (N_26468,N_24317,N_24187);
or U26469 (N_26469,N_25250,N_25532);
nor U26470 (N_26470,N_24081,N_25651);
xnor U26471 (N_26471,N_24717,N_24664);
or U26472 (N_26472,N_25933,N_25747);
xnor U26473 (N_26473,N_25533,N_24991);
nand U26474 (N_26474,N_25011,N_25726);
nand U26475 (N_26475,N_25648,N_24549);
or U26476 (N_26476,N_25794,N_25122);
xor U26477 (N_26477,N_25087,N_24219);
or U26478 (N_26478,N_24058,N_24468);
xnor U26479 (N_26479,N_24291,N_25415);
nor U26480 (N_26480,N_24639,N_24384);
nor U26481 (N_26481,N_24009,N_25833);
or U26482 (N_26482,N_24996,N_24809);
xor U26483 (N_26483,N_25828,N_24541);
xor U26484 (N_26484,N_24182,N_25458);
nor U26485 (N_26485,N_25872,N_24624);
nand U26486 (N_26486,N_25513,N_24125);
nor U26487 (N_26487,N_25064,N_25447);
nand U26488 (N_26488,N_25565,N_24401);
nor U26489 (N_26489,N_25906,N_24492);
or U26490 (N_26490,N_25049,N_24318);
xor U26491 (N_26491,N_24752,N_24803);
and U26492 (N_26492,N_24086,N_25016);
and U26493 (N_26493,N_25550,N_24152);
xnor U26494 (N_26494,N_24223,N_25583);
or U26495 (N_26495,N_25715,N_25556);
or U26496 (N_26496,N_24041,N_25840);
nor U26497 (N_26497,N_24479,N_25575);
or U26498 (N_26498,N_24162,N_24995);
xor U26499 (N_26499,N_24043,N_24895);
or U26500 (N_26500,N_24870,N_25214);
and U26501 (N_26501,N_25701,N_25359);
or U26502 (N_26502,N_25143,N_25991);
or U26503 (N_26503,N_24737,N_24480);
xnor U26504 (N_26504,N_24674,N_24656);
xnor U26505 (N_26505,N_24424,N_25046);
nor U26506 (N_26506,N_24044,N_24804);
nand U26507 (N_26507,N_24901,N_24374);
and U26508 (N_26508,N_24831,N_25679);
nand U26509 (N_26509,N_24501,N_24292);
or U26510 (N_26510,N_25303,N_25124);
nor U26511 (N_26511,N_24454,N_24419);
xnor U26512 (N_26512,N_25287,N_24057);
nand U26513 (N_26513,N_25098,N_25100);
or U26514 (N_26514,N_25483,N_25390);
nand U26515 (N_26515,N_25772,N_25632);
nor U26516 (N_26516,N_24906,N_25983);
and U26517 (N_26517,N_24028,N_25666);
nor U26518 (N_26518,N_25443,N_24030);
nand U26519 (N_26519,N_24045,N_24194);
and U26520 (N_26520,N_25108,N_25080);
nor U26521 (N_26521,N_24261,N_25056);
nand U26522 (N_26522,N_24473,N_24791);
nor U26523 (N_26523,N_25385,N_25402);
and U26524 (N_26524,N_24897,N_25868);
or U26525 (N_26525,N_25526,N_24465);
nand U26526 (N_26526,N_24459,N_24108);
nor U26527 (N_26527,N_25058,N_25188);
or U26528 (N_26528,N_25295,N_24616);
xor U26529 (N_26529,N_25805,N_25826);
xnor U26530 (N_26530,N_24021,N_24145);
and U26531 (N_26531,N_25320,N_25015);
nand U26532 (N_26532,N_24601,N_25622);
xor U26533 (N_26533,N_24472,N_25169);
and U26534 (N_26534,N_25292,N_25845);
and U26535 (N_26535,N_25145,N_24612);
nor U26536 (N_26536,N_25905,N_24210);
and U26537 (N_26537,N_24773,N_24441);
and U26538 (N_26538,N_25346,N_25001);
xor U26539 (N_26539,N_25870,N_25290);
and U26540 (N_26540,N_25319,N_24263);
nand U26541 (N_26541,N_24968,N_25789);
nand U26542 (N_26542,N_24427,N_25896);
xnor U26543 (N_26543,N_25277,N_24537);
xnor U26544 (N_26544,N_25553,N_25943);
nand U26545 (N_26545,N_25861,N_24613);
nand U26546 (N_26546,N_25161,N_24197);
nor U26547 (N_26547,N_24808,N_24406);
nor U26548 (N_26548,N_25265,N_25477);
nand U26549 (N_26549,N_24192,N_24293);
or U26550 (N_26550,N_24830,N_25975);
xor U26551 (N_26551,N_25644,N_25489);
nand U26552 (N_26552,N_25956,N_24853);
nor U26553 (N_26553,N_25401,N_25042);
nor U26554 (N_26554,N_24994,N_24565);
nand U26555 (N_26555,N_25730,N_25607);
or U26556 (N_26556,N_25783,N_25803);
xor U26557 (N_26557,N_25094,N_24579);
and U26558 (N_26558,N_24141,N_25977);
nor U26559 (N_26559,N_24383,N_25272);
or U26560 (N_26560,N_25004,N_25234);
or U26561 (N_26561,N_25634,N_24727);
and U26562 (N_26562,N_24966,N_25686);
or U26563 (N_26563,N_25802,N_25586);
or U26564 (N_26564,N_25019,N_24970);
and U26565 (N_26565,N_25855,N_24122);
nor U26566 (N_26566,N_24512,N_25930);
xor U26567 (N_26567,N_24827,N_25332);
nor U26568 (N_26568,N_24540,N_25478);
and U26569 (N_26569,N_25403,N_25182);
nand U26570 (N_26570,N_24842,N_25368);
or U26571 (N_26571,N_25552,N_24475);
and U26572 (N_26572,N_24636,N_25937);
nor U26573 (N_26573,N_24469,N_25373);
nor U26574 (N_26574,N_24915,N_24873);
or U26575 (N_26575,N_24337,N_25916);
xor U26576 (N_26576,N_25119,N_25106);
nand U26577 (N_26577,N_24193,N_24326);
xor U26578 (N_26578,N_25302,N_25885);
xor U26579 (N_26579,N_25817,N_24016);
or U26580 (N_26580,N_24894,N_25537);
and U26581 (N_26581,N_25298,N_25858);
and U26582 (N_26582,N_24730,N_25367);
or U26583 (N_26583,N_24981,N_24013);
nand U26584 (N_26584,N_24522,N_25917);
nand U26585 (N_26585,N_25311,N_24849);
or U26586 (N_26586,N_25293,N_24158);
and U26587 (N_26587,N_25713,N_24367);
nor U26588 (N_26588,N_24515,N_24121);
nand U26589 (N_26589,N_24118,N_25233);
and U26590 (N_26590,N_24642,N_24518);
nor U26591 (N_26591,N_25727,N_25162);
and U26592 (N_26592,N_24148,N_24423);
nor U26593 (N_26593,N_25220,N_24077);
or U26594 (N_26594,N_24953,N_25485);
xnor U26595 (N_26595,N_24312,N_25738);
nor U26596 (N_26596,N_24972,N_24824);
nand U26597 (N_26597,N_24923,N_25712);
xor U26598 (N_26598,N_25544,N_25654);
xnor U26599 (N_26599,N_25196,N_25661);
nand U26600 (N_26600,N_24595,N_24227);
xor U26601 (N_26601,N_25309,N_25184);
nor U26602 (N_26602,N_24826,N_24767);
xor U26603 (N_26603,N_24255,N_25070);
and U26604 (N_26604,N_24633,N_25377);
nand U26605 (N_26605,N_24666,N_25424);
or U26606 (N_26606,N_24332,N_24950);
nor U26607 (N_26607,N_25534,N_25850);
xor U26608 (N_26608,N_25699,N_24431);
and U26609 (N_26609,N_24757,N_25066);
or U26610 (N_26610,N_24026,N_24653);
nor U26611 (N_26611,N_24129,N_24218);
and U26612 (N_26612,N_25999,N_24505);
or U26613 (N_26613,N_24353,N_24807);
nor U26614 (N_26614,N_25316,N_24321);
xor U26615 (N_26615,N_24560,N_25097);
nand U26616 (N_26616,N_24429,N_25232);
xor U26617 (N_26617,N_24436,N_24224);
and U26618 (N_26618,N_25133,N_24324);
nand U26619 (N_26619,N_25791,N_25626);
xor U26620 (N_26620,N_25777,N_24813);
nor U26621 (N_26621,N_25413,N_25569);
and U26622 (N_26622,N_25920,N_24477);
nand U26623 (N_26623,N_24344,N_25843);
nor U26624 (N_26624,N_24386,N_25814);
nand U26625 (N_26625,N_24241,N_25223);
nor U26626 (N_26626,N_24783,N_24232);
nand U26627 (N_26627,N_25081,N_25570);
and U26628 (N_26628,N_25759,N_24858);
or U26629 (N_26629,N_25948,N_24380);
nand U26630 (N_26630,N_25408,N_24185);
xor U26631 (N_26631,N_24453,N_25437);
or U26632 (N_26632,N_24782,N_24101);
xnor U26633 (N_26633,N_24967,N_25469);
or U26634 (N_26634,N_24400,N_25678);
xnor U26635 (N_26635,N_24931,N_24969);
nor U26636 (N_26636,N_24073,N_25215);
xnor U26637 (N_26637,N_25323,N_25704);
or U26638 (N_26638,N_24837,N_25398);
and U26639 (N_26639,N_25118,N_25134);
and U26640 (N_26640,N_24346,N_24507);
nor U26641 (N_26641,N_25864,N_24686);
nor U26642 (N_26642,N_24049,N_25236);
or U26643 (N_26643,N_25518,N_25555);
xor U26644 (N_26644,N_24975,N_24714);
nor U26645 (N_26645,N_24136,N_25246);
xnor U26646 (N_26646,N_24533,N_25149);
nand U26647 (N_26647,N_25312,N_25150);
or U26648 (N_26648,N_24381,N_24877);
xnor U26649 (N_26649,N_25096,N_24547);
nor U26650 (N_26650,N_25481,N_24843);
xnor U26651 (N_26651,N_25479,N_24875);
nor U26652 (N_26652,N_24157,N_24564);
nand U26653 (N_26653,N_25120,N_25434);
xor U26654 (N_26654,N_25322,N_25333);
or U26655 (N_26655,N_25063,N_25423);
or U26656 (N_26656,N_25363,N_25953);
or U26657 (N_26657,N_25846,N_25524);
and U26658 (N_26658,N_25614,N_25410);
nor U26659 (N_26659,N_24072,N_24029);
and U26660 (N_26660,N_25507,N_24763);
or U26661 (N_26661,N_25618,N_24150);
xnor U26662 (N_26662,N_25285,N_25875);
and U26663 (N_26663,N_24673,N_25659);
xor U26664 (N_26664,N_25270,N_24304);
or U26665 (N_26665,N_25717,N_24964);
or U26666 (N_26666,N_24835,N_25988);
nand U26667 (N_26667,N_24207,N_25335);
nand U26668 (N_26668,N_24238,N_24871);
nand U26669 (N_26669,N_25967,N_24080);
and U26670 (N_26670,N_24863,N_25033);
or U26671 (N_26671,N_25259,N_25510);
xor U26672 (N_26672,N_24133,N_24350);
nand U26673 (N_26673,N_25529,N_25775);
and U26674 (N_26674,N_25391,N_24075);
nand U26675 (N_26675,N_25506,N_25027);
xor U26676 (N_26676,N_24759,N_24228);
or U26677 (N_26677,N_24554,N_25758);
nand U26678 (N_26678,N_24825,N_25347);
nor U26679 (N_26679,N_25683,N_24047);
nor U26680 (N_26680,N_25009,N_24984);
or U26681 (N_26681,N_24670,N_24276);
or U26682 (N_26682,N_24027,N_25425);
nand U26683 (N_26683,N_24535,N_25017);
and U26684 (N_26684,N_25551,N_25191);
or U26685 (N_26685,N_24256,N_25725);
and U26686 (N_26686,N_24295,N_24444);
and U26687 (N_26687,N_25921,N_25255);
and U26688 (N_26688,N_25950,N_24658);
and U26689 (N_26689,N_25441,N_25739);
or U26690 (N_26690,N_25806,N_24976);
or U26691 (N_26691,N_24816,N_25440);
xor U26692 (N_26692,N_24012,N_25729);
nand U26693 (N_26693,N_24609,N_25093);
nor U26694 (N_26694,N_24648,N_24345);
xor U26695 (N_26695,N_24680,N_24502);
or U26696 (N_26696,N_25849,N_24220);
nand U26697 (N_26697,N_24392,N_25008);
and U26698 (N_26698,N_25606,N_24349);
and U26699 (N_26699,N_25735,N_25649);
xor U26700 (N_26700,N_25123,N_25456);
xor U26701 (N_26701,N_24938,N_25509);
xnor U26702 (N_26702,N_25026,N_25631);
nor U26703 (N_26703,N_24287,N_24017);
or U26704 (N_26704,N_24977,N_25103);
nand U26705 (N_26705,N_25073,N_25625);
or U26706 (N_26706,N_24989,N_25327);
xnor U26707 (N_26707,N_25502,N_25164);
nand U26708 (N_26708,N_24449,N_24634);
or U26709 (N_26709,N_24278,N_24083);
nand U26710 (N_26710,N_24090,N_25273);
and U26711 (N_26711,N_24637,N_24635);
nand U26712 (N_26712,N_24701,N_24418);
xor U26713 (N_26713,N_25014,N_24425);
or U26714 (N_26714,N_24589,N_24008);
nor U26715 (N_26715,N_24646,N_25047);
nand U26716 (N_26716,N_24596,N_25559);
xor U26717 (N_26717,N_25604,N_25914);
nand U26718 (N_26718,N_25253,N_25753);
or U26719 (N_26719,N_24760,N_25793);
and U26720 (N_26720,N_24439,N_24437);
xor U26721 (N_26721,N_24231,N_25370);
nand U26722 (N_26722,N_25774,N_25459);
xor U26723 (N_26723,N_25557,N_25584);
nand U26724 (N_26724,N_24559,N_25488);
or U26725 (N_26725,N_24765,N_25038);
and U26726 (N_26726,N_25694,N_25866);
nand U26727 (N_26727,N_25330,N_24123);
or U26728 (N_26728,N_25095,N_25612);
and U26729 (N_26729,N_24672,N_24206);
nor U26730 (N_26730,N_25742,N_24284);
xnor U26731 (N_26731,N_24209,N_24685);
nor U26732 (N_26732,N_25760,N_25448);
or U26733 (N_26733,N_25852,N_24695);
nand U26734 (N_26734,N_25667,N_25301);
xor U26735 (N_26735,N_25392,N_25059);
or U26736 (N_26736,N_25203,N_25531);
or U26737 (N_26737,N_24181,N_24731);
nand U26738 (N_26738,N_24426,N_24105);
nor U26739 (N_26739,N_24949,N_24298);
xor U26740 (N_26740,N_24513,N_24904);
nor U26741 (N_26741,N_25818,N_25498);
and U26742 (N_26742,N_24785,N_24402);
nor U26743 (N_26743,N_24042,N_25968);
nor U26744 (N_26744,N_25756,N_24725);
and U26745 (N_26745,N_24688,N_24708);
or U26746 (N_26746,N_24061,N_24171);
nor U26747 (N_26747,N_24719,N_25900);
or U26748 (N_26748,N_25132,N_25454);
or U26749 (N_26749,N_25353,N_25879);
nor U26750 (N_26750,N_24048,N_24792);
nor U26751 (N_26751,N_24239,N_24850);
or U26752 (N_26752,N_24300,N_25278);
xnor U26753 (N_26753,N_25116,N_24252);
and U26754 (N_26754,N_25492,N_25808);
nor U26755 (N_26755,N_24354,N_25603);
and U26756 (N_26756,N_24107,N_24498);
nor U26757 (N_26757,N_25707,N_24935);
and U26758 (N_26758,N_25482,N_24650);
nor U26759 (N_26759,N_24435,N_25342);
xnor U26760 (N_26760,N_25832,N_24649);
and U26761 (N_26761,N_25835,N_25324);
or U26762 (N_26762,N_24474,N_25630);
xnor U26763 (N_26763,N_25653,N_24490);
and U26764 (N_26764,N_25449,N_25204);
or U26765 (N_26765,N_24713,N_25824);
and U26766 (N_26766,N_25170,N_25393);
or U26767 (N_26767,N_24096,N_24069);
xnor U26768 (N_26768,N_25418,N_24151);
nor U26769 (N_26769,N_25608,N_24301);
nand U26770 (N_26770,N_25716,N_24333);
nor U26771 (N_26771,N_24741,N_24170);
xor U26772 (N_26772,N_24797,N_25155);
nor U26773 (N_26773,N_24066,N_25767);
nor U26774 (N_26774,N_25788,N_24279);
xnor U26775 (N_26775,N_24526,N_25256);
or U26776 (N_26776,N_25079,N_25198);
xnor U26777 (N_26777,N_24764,N_24529);
xor U26778 (N_26778,N_24922,N_25180);
nand U26779 (N_26779,N_24662,N_24552);
nor U26780 (N_26780,N_25691,N_25247);
nor U26781 (N_26781,N_25052,N_25039);
and U26782 (N_26782,N_25361,N_25548);
nor U26783 (N_26783,N_24260,N_25745);
nand U26784 (N_26784,N_25076,N_25216);
xnor U26785 (N_26785,N_24415,N_24280);
or U26786 (N_26786,N_25633,N_24319);
nand U26787 (N_26787,N_24000,N_24644);
xnor U26788 (N_26788,N_25036,N_24390);
xor U26789 (N_26789,N_24094,N_24200);
xor U26790 (N_26790,N_25724,N_25267);
or U26791 (N_26791,N_24683,N_25580);
or U26792 (N_26792,N_24917,N_24215);
xnor U26793 (N_26793,N_25306,N_24216);
nor U26794 (N_26794,N_25243,N_24571);
nor U26795 (N_26795,N_25823,N_24046);
nor U26796 (N_26796,N_25961,N_25527);
xor U26797 (N_26797,N_25754,N_25372);
or U26798 (N_26798,N_24325,N_24062);
or U26799 (N_26799,N_24294,N_25602);
nand U26800 (N_26800,N_25721,N_25741);
or U26801 (N_26801,N_24962,N_25279);
nor U26802 (N_26802,N_24762,N_24514);
and U26803 (N_26803,N_25821,N_24558);
and U26804 (N_26804,N_25432,N_25796);
nor U26805 (N_26805,N_24355,N_25723);
nor U26806 (N_26806,N_25809,N_24729);
nor U26807 (N_26807,N_24303,N_24011);
xor U26808 (N_26808,N_24403,N_24471);
and U26809 (N_26809,N_24456,N_25615);
or U26810 (N_26810,N_25400,N_24348);
xor U26811 (N_26811,N_24534,N_25022);
and U26812 (N_26812,N_24509,N_24909);
nand U26813 (N_26813,N_25012,N_24876);
nand U26814 (N_26814,N_24097,N_25784);
nor U26815 (N_26815,N_24434,N_25193);
nor U26816 (N_26816,N_25669,N_25938);
xor U26817 (N_26817,N_24364,N_24022);
xnor U26818 (N_26818,N_25981,N_25528);
nor U26819 (N_26819,N_25305,N_25168);
nor U26820 (N_26820,N_25973,N_24784);
nand U26821 (N_26821,N_25997,N_24841);
and U26822 (N_26822,N_25421,N_24031);
xnor U26823 (N_26823,N_25192,N_25354);
and U26824 (N_26824,N_24388,N_25291);
and U26825 (N_26825,N_24703,N_25675);
and U26826 (N_26826,N_25473,N_24776);
or U26827 (N_26827,N_24557,N_24483);
and U26828 (N_26828,N_24088,N_25304);
xnor U26829 (N_26829,N_24893,N_25766);
nor U26830 (N_26830,N_24777,N_24457);
nand U26831 (N_26831,N_24357,N_25893);
or U26832 (N_26832,N_25172,N_25960);
xnor U26833 (N_26833,N_24795,N_25880);
nand U26834 (N_26834,N_24640,N_25799);
or U26835 (N_26835,N_25455,N_24556);
nand U26836 (N_26836,N_25201,N_24433);
xnor U26837 (N_26837,N_24684,N_25857);
or U26838 (N_26838,N_24032,N_24772);
nand U26839 (N_26839,N_25213,N_24573);
nand U26840 (N_26840,N_25578,N_25321);
xor U26841 (N_26841,N_25144,N_24455);
xnor U26842 (N_26842,N_24751,N_24761);
or U26843 (N_26843,N_24581,N_25851);
or U26844 (N_26844,N_25804,N_24466);
nand U26845 (N_26845,N_25314,N_24438);
or U26846 (N_26846,N_25348,N_24811);
nand U26847 (N_26847,N_24545,N_24411);
or U26848 (N_26848,N_24869,N_25417);
or U26849 (N_26849,N_24720,N_25474);
and U26850 (N_26850,N_25297,N_25141);
xnor U26851 (N_26851,N_24523,N_24063);
nor U26852 (N_26852,N_24679,N_24339);
xnor U26853 (N_26853,N_24155,N_24446);
xnor U26854 (N_26854,N_24338,N_24409);
nor U26855 (N_26855,N_25493,N_24420);
nand U26856 (N_26856,N_24531,N_24103);
nor U26857 (N_26857,N_25325,N_24285);
nor U26858 (N_26858,N_24508,N_24351);
and U26859 (N_26859,N_24430,N_24610);
and U26860 (N_26860,N_25262,N_24211);
nor U26861 (N_26861,N_25226,N_25719);
xnor U26862 (N_26862,N_25752,N_25993);
xnor U26863 (N_26863,N_24659,N_24665);
nand U26864 (N_26864,N_24230,N_24880);
xnor U26865 (N_26865,N_25153,N_24331);
or U26866 (N_26866,N_25147,N_25466);
xnor U26867 (N_26867,N_24407,N_24704);
nor U26868 (N_26868,N_25275,N_25101);
or U26869 (N_26869,N_24413,N_24709);
xor U26870 (N_26870,N_25175,N_25645);
and U26871 (N_26871,N_25677,N_24440);
nand U26872 (N_26872,N_25812,N_24973);
nand U26873 (N_26873,N_24035,N_25187);
nand U26874 (N_26874,N_25383,N_24159);
or U26875 (N_26875,N_25663,N_25635);
nor U26876 (N_26876,N_25152,N_24990);
or U26877 (N_26877,N_24282,N_24947);
and U26878 (N_26878,N_25167,N_24308);
nor U26879 (N_26879,N_24979,N_24930);
nand U26880 (N_26880,N_24208,N_25436);
nor U26881 (N_26881,N_24038,N_25813);
or U26882 (N_26882,N_24896,N_25102);
and U26883 (N_26883,N_25939,N_24521);
nand U26884 (N_26884,N_24237,N_25599);
xnor U26885 (N_26885,N_24548,N_24860);
or U26886 (N_26886,N_25687,N_24978);
nand U26887 (N_26887,N_24307,N_24847);
xor U26888 (N_26888,N_25438,N_24780);
nor U26889 (N_26889,N_24965,N_24606);
nor U26890 (N_26890,N_25450,N_24202);
nand U26891 (N_26891,N_25910,N_24974);
or U26892 (N_26892,N_25693,N_24594);
xnor U26893 (N_26893,N_25865,N_25807);
nand U26894 (N_26894,N_24131,N_25343);
nand U26895 (N_26895,N_24493,N_25117);
nand U26896 (N_26896,N_24137,N_25761);
xnor U26897 (N_26897,N_24235,N_24417);
and U26898 (N_26898,N_24405,N_24861);
nand U26899 (N_26899,N_25453,N_25903);
or U26900 (N_26900,N_24266,N_25276);
xnor U26901 (N_26901,N_25258,N_24499);
or U26902 (N_26902,N_24963,N_24365);
nor U26903 (N_26903,N_24789,N_24327);
xor U26904 (N_26904,N_25503,N_25573);
nor U26905 (N_26905,N_25151,N_24584);
nor U26906 (N_26906,N_24698,N_24517);
or U26907 (N_26907,N_24421,N_25671);
nand U26908 (N_26908,N_24481,N_24156);
nand U26909 (N_26909,N_25090,N_25148);
nand U26910 (N_26910,N_25266,N_25856);
and U26911 (N_26911,N_25068,N_25177);
xnor U26912 (N_26912,N_24678,N_24033);
xnor U26913 (N_26913,N_24074,N_24626);
xnor U26914 (N_26914,N_24707,N_24281);
and U26915 (N_26915,N_24329,N_25360);
nor U26916 (N_26916,N_25610,N_25985);
and U26917 (N_26917,N_25688,N_24746);
nand U26918 (N_26918,N_24676,N_24544);
and U26919 (N_26919,N_24983,N_25837);
nand U26920 (N_26920,N_24566,N_24289);
and U26921 (N_26921,N_24361,N_24550);
xnor U26922 (N_26922,N_24394,N_25924);
xnor U26923 (N_26923,N_25762,N_25984);
xnor U26924 (N_26924,N_25926,N_24582);
nor U26925 (N_26925,N_25189,N_24700);
nand U26926 (N_26926,N_25497,N_25690);
nand U26927 (N_26927,N_24722,N_24925);
nor U26928 (N_26928,N_25613,N_25054);
nand U26929 (N_26929,N_25969,N_25340);
xor U26930 (N_26930,N_25200,N_25505);
or U26931 (N_26931,N_25088,N_24060);
xor U26932 (N_26932,N_25773,N_24258);
nor U26933 (N_26933,N_24583,N_25217);
nor U26934 (N_26934,N_25062,N_25562);
and U26935 (N_26935,N_24605,N_24834);
or U26936 (N_26936,N_24829,N_25963);
or U26937 (N_26937,N_24859,N_25211);
xnor U26938 (N_26938,N_24563,N_24872);
nor U26939 (N_26939,N_24172,N_24844);
nand U26940 (N_26940,N_24745,N_24691);
or U26941 (N_26941,N_24036,N_25110);
nor U26942 (N_26942,N_25202,N_24916);
and U26943 (N_26943,N_25831,N_24286);
and U26944 (N_26944,N_24575,N_24163);
and U26945 (N_26945,N_25765,N_25908);
nand U26946 (N_26946,N_24525,N_24898);
or U26947 (N_26947,N_25251,N_25889);
nor U26948 (N_26948,N_25940,N_24788);
or U26949 (N_26949,N_24358,N_24174);
or U26950 (N_26950,N_25179,N_25045);
and U26951 (N_26951,N_24886,N_24199);
and U26952 (N_26952,N_24204,N_24126);
nand U26953 (N_26953,N_24109,N_25888);
nor U26954 (N_26954,N_24053,N_25894);
and U26955 (N_26955,N_25535,N_24111);
nor U26956 (N_26956,N_25982,N_24377);
xor U26957 (N_26957,N_25248,N_24948);
or U26958 (N_26958,N_24138,N_25623);
xor U26959 (N_26959,N_24356,N_24868);
xnor U26960 (N_26960,N_25078,N_25294);
and U26961 (N_26961,N_25763,N_24311);
nor U26962 (N_26962,N_25412,N_25931);
or U26963 (N_26963,N_24020,N_24488);
nor U26964 (N_26964,N_25010,N_24149);
or U26965 (N_26965,N_25420,N_24866);
and U26966 (N_26966,N_25376,N_24932);
or U26967 (N_26967,N_24578,N_25945);
nand U26968 (N_26968,N_24283,N_24470);
and U26969 (N_26969,N_25563,N_25013);
nand U26970 (N_26970,N_25974,N_25966);
nand U26971 (N_26971,N_25225,N_24334);
and U26972 (N_26972,N_24562,N_24603);
xnor U26973 (N_26973,N_25710,N_25375);
nand U26974 (N_26974,N_24845,N_25883);
nand U26975 (N_26975,N_25219,N_25842);
or U26976 (N_26976,N_24621,N_24724);
or U26977 (N_26977,N_24555,N_24661);
nor U26978 (N_26978,N_24753,N_25734);
or U26979 (N_26979,N_24267,N_25114);
nor U26980 (N_26980,N_25084,N_25126);
xor U26981 (N_26981,N_25005,N_24926);
xnor U26982 (N_26982,N_25871,N_24892);
or U26983 (N_26983,N_25069,N_25892);
or U26984 (N_26984,N_25829,N_25397);
nor U26985 (N_26985,N_25597,N_24846);
nor U26986 (N_26986,N_24106,N_24511);
nor U26987 (N_26987,N_25349,N_25284);
xor U26988 (N_26988,N_24203,N_24039);
and U26989 (N_26989,N_25244,N_25616);
or U26990 (N_26990,N_24432,N_25357);
xor U26991 (N_26991,N_24506,N_25176);
xnor U26992 (N_26992,N_25422,N_25617);
nand U26993 (N_26993,N_25471,N_25018);
and U26994 (N_26994,N_25465,N_25887);
nand U26995 (N_26995,N_24524,N_25197);
and U26996 (N_26996,N_25830,N_24450);
nand U26997 (N_26997,N_24222,N_24005);
and U26998 (N_26998,N_24854,N_24391);
nand U26999 (N_26999,N_25000,N_25129);
and U27000 (N_27000,N_25210,N_24833);
nand U27001 (N_27001,N_24045,N_24447);
nor U27002 (N_27002,N_25078,N_24616);
nor U27003 (N_27003,N_25539,N_25815);
nor U27004 (N_27004,N_24563,N_25268);
or U27005 (N_27005,N_24987,N_25365);
nor U27006 (N_27006,N_24353,N_25159);
nand U27007 (N_27007,N_24548,N_25470);
nand U27008 (N_27008,N_24665,N_25263);
xnor U27009 (N_27009,N_24208,N_24863);
nand U27010 (N_27010,N_24908,N_25149);
or U27011 (N_27011,N_24570,N_25303);
and U27012 (N_27012,N_25892,N_25189);
nand U27013 (N_27013,N_25442,N_24766);
and U27014 (N_27014,N_25108,N_24908);
nand U27015 (N_27015,N_25472,N_24937);
nand U27016 (N_27016,N_25679,N_25395);
or U27017 (N_27017,N_25199,N_24131);
nand U27018 (N_27018,N_24225,N_25077);
xor U27019 (N_27019,N_25933,N_24487);
xor U27020 (N_27020,N_24991,N_25579);
nor U27021 (N_27021,N_25525,N_25024);
nor U27022 (N_27022,N_24934,N_25906);
and U27023 (N_27023,N_25116,N_24313);
or U27024 (N_27024,N_25718,N_25556);
and U27025 (N_27025,N_24006,N_25372);
nor U27026 (N_27026,N_24843,N_24189);
or U27027 (N_27027,N_24031,N_25145);
nand U27028 (N_27028,N_25813,N_24032);
nand U27029 (N_27029,N_24663,N_25331);
nor U27030 (N_27030,N_24203,N_25652);
nand U27031 (N_27031,N_25985,N_25558);
nor U27032 (N_27032,N_25993,N_24000);
nor U27033 (N_27033,N_24647,N_25899);
and U27034 (N_27034,N_25101,N_25829);
nand U27035 (N_27035,N_24698,N_24438);
or U27036 (N_27036,N_24083,N_25117);
nor U27037 (N_27037,N_25169,N_25809);
xor U27038 (N_27038,N_25270,N_25471);
nand U27039 (N_27039,N_25576,N_24159);
nor U27040 (N_27040,N_25126,N_25372);
xnor U27041 (N_27041,N_25088,N_25010);
or U27042 (N_27042,N_24571,N_25934);
nand U27043 (N_27043,N_24971,N_25280);
or U27044 (N_27044,N_25764,N_24399);
nand U27045 (N_27045,N_24080,N_25953);
and U27046 (N_27046,N_24699,N_24670);
and U27047 (N_27047,N_24364,N_25660);
and U27048 (N_27048,N_25368,N_24085);
xnor U27049 (N_27049,N_25412,N_24282);
nand U27050 (N_27050,N_25326,N_24084);
and U27051 (N_27051,N_25086,N_24251);
xnor U27052 (N_27052,N_24975,N_25901);
xnor U27053 (N_27053,N_24291,N_24942);
nand U27054 (N_27054,N_24624,N_25315);
or U27055 (N_27055,N_25162,N_24584);
and U27056 (N_27056,N_25429,N_24461);
or U27057 (N_27057,N_25812,N_24096);
or U27058 (N_27058,N_24333,N_24262);
and U27059 (N_27059,N_25579,N_25066);
nand U27060 (N_27060,N_24821,N_25738);
nor U27061 (N_27061,N_25271,N_24072);
xnor U27062 (N_27062,N_25009,N_25453);
and U27063 (N_27063,N_25026,N_25233);
or U27064 (N_27064,N_24678,N_25008);
nor U27065 (N_27065,N_25180,N_25331);
xor U27066 (N_27066,N_24489,N_24630);
and U27067 (N_27067,N_24401,N_24044);
xor U27068 (N_27068,N_25623,N_25316);
xor U27069 (N_27069,N_24326,N_25962);
or U27070 (N_27070,N_24908,N_25344);
nand U27071 (N_27071,N_24684,N_25130);
nand U27072 (N_27072,N_24837,N_25406);
xor U27073 (N_27073,N_25294,N_24203);
xnor U27074 (N_27074,N_24984,N_25180);
nand U27075 (N_27075,N_24572,N_25869);
or U27076 (N_27076,N_24273,N_24428);
nand U27077 (N_27077,N_24334,N_24070);
nand U27078 (N_27078,N_25749,N_24727);
and U27079 (N_27079,N_24728,N_25063);
xor U27080 (N_27080,N_25899,N_24332);
xnor U27081 (N_27081,N_24651,N_25844);
nor U27082 (N_27082,N_25983,N_25540);
and U27083 (N_27083,N_24591,N_25995);
and U27084 (N_27084,N_25722,N_25195);
or U27085 (N_27085,N_24599,N_24176);
nand U27086 (N_27086,N_25716,N_25752);
or U27087 (N_27087,N_25405,N_25683);
xnor U27088 (N_27088,N_24284,N_24162);
nand U27089 (N_27089,N_24191,N_25656);
nor U27090 (N_27090,N_24969,N_24239);
and U27091 (N_27091,N_24161,N_24734);
nand U27092 (N_27092,N_24604,N_24467);
nand U27093 (N_27093,N_24644,N_24580);
nor U27094 (N_27094,N_24932,N_24050);
nand U27095 (N_27095,N_25805,N_24953);
xor U27096 (N_27096,N_24769,N_24301);
xor U27097 (N_27097,N_24786,N_24528);
and U27098 (N_27098,N_25896,N_25410);
xnor U27099 (N_27099,N_24802,N_24498);
and U27100 (N_27100,N_24851,N_25019);
xnor U27101 (N_27101,N_25263,N_24455);
nor U27102 (N_27102,N_24292,N_24592);
and U27103 (N_27103,N_25439,N_24958);
or U27104 (N_27104,N_24764,N_25634);
nor U27105 (N_27105,N_25984,N_24018);
xnor U27106 (N_27106,N_25860,N_25954);
xor U27107 (N_27107,N_24027,N_25575);
nor U27108 (N_27108,N_25061,N_24898);
and U27109 (N_27109,N_25643,N_24621);
and U27110 (N_27110,N_24405,N_25551);
and U27111 (N_27111,N_25718,N_24280);
or U27112 (N_27112,N_24943,N_24311);
or U27113 (N_27113,N_25506,N_24223);
or U27114 (N_27114,N_24436,N_24709);
and U27115 (N_27115,N_25792,N_25545);
and U27116 (N_27116,N_24613,N_24440);
nor U27117 (N_27117,N_25640,N_25117);
or U27118 (N_27118,N_25028,N_24778);
or U27119 (N_27119,N_24818,N_24095);
nand U27120 (N_27120,N_25300,N_24854);
xnor U27121 (N_27121,N_25269,N_24717);
xnor U27122 (N_27122,N_24258,N_24119);
nor U27123 (N_27123,N_25314,N_24830);
or U27124 (N_27124,N_24149,N_25826);
and U27125 (N_27125,N_25270,N_25306);
nand U27126 (N_27126,N_25693,N_25867);
nand U27127 (N_27127,N_24121,N_25567);
nand U27128 (N_27128,N_25616,N_25317);
nand U27129 (N_27129,N_25752,N_24662);
or U27130 (N_27130,N_25575,N_24679);
or U27131 (N_27131,N_24152,N_25859);
and U27132 (N_27132,N_25050,N_24422);
and U27133 (N_27133,N_24900,N_24356);
nor U27134 (N_27134,N_24403,N_24794);
nor U27135 (N_27135,N_24066,N_25482);
nand U27136 (N_27136,N_24319,N_25706);
nand U27137 (N_27137,N_25783,N_24022);
and U27138 (N_27138,N_24924,N_24798);
nor U27139 (N_27139,N_25908,N_24932);
and U27140 (N_27140,N_24232,N_25938);
and U27141 (N_27141,N_24152,N_25526);
and U27142 (N_27142,N_24112,N_25953);
nand U27143 (N_27143,N_25997,N_25004);
and U27144 (N_27144,N_24046,N_25966);
nand U27145 (N_27145,N_25359,N_25345);
nand U27146 (N_27146,N_24757,N_24094);
or U27147 (N_27147,N_24100,N_24724);
nand U27148 (N_27148,N_25057,N_24423);
xnor U27149 (N_27149,N_24892,N_24021);
xor U27150 (N_27150,N_24763,N_25312);
xor U27151 (N_27151,N_25818,N_24955);
and U27152 (N_27152,N_24663,N_25778);
nor U27153 (N_27153,N_24034,N_24524);
or U27154 (N_27154,N_25058,N_24268);
nand U27155 (N_27155,N_25283,N_25487);
nor U27156 (N_27156,N_25298,N_24602);
and U27157 (N_27157,N_24552,N_24214);
nor U27158 (N_27158,N_25510,N_24150);
or U27159 (N_27159,N_24828,N_24576);
xnor U27160 (N_27160,N_25742,N_24489);
xnor U27161 (N_27161,N_25096,N_25381);
and U27162 (N_27162,N_25008,N_25905);
and U27163 (N_27163,N_25820,N_24021);
xnor U27164 (N_27164,N_25928,N_25738);
and U27165 (N_27165,N_24016,N_25830);
xnor U27166 (N_27166,N_25808,N_24095);
nand U27167 (N_27167,N_24920,N_25735);
or U27168 (N_27168,N_25979,N_25659);
nor U27169 (N_27169,N_25759,N_24956);
and U27170 (N_27170,N_25297,N_24326);
xor U27171 (N_27171,N_25308,N_25524);
and U27172 (N_27172,N_24191,N_25891);
nand U27173 (N_27173,N_25234,N_24661);
nor U27174 (N_27174,N_24056,N_25577);
nor U27175 (N_27175,N_24274,N_24174);
nor U27176 (N_27176,N_25647,N_24942);
and U27177 (N_27177,N_24657,N_25277);
xnor U27178 (N_27178,N_24119,N_25909);
and U27179 (N_27179,N_25636,N_25307);
nand U27180 (N_27180,N_24965,N_24377);
and U27181 (N_27181,N_24760,N_25921);
xor U27182 (N_27182,N_24639,N_25335);
nor U27183 (N_27183,N_24068,N_25183);
xor U27184 (N_27184,N_25582,N_24787);
xor U27185 (N_27185,N_24203,N_25037);
and U27186 (N_27186,N_24486,N_25230);
and U27187 (N_27187,N_24379,N_25999);
and U27188 (N_27188,N_25437,N_25182);
or U27189 (N_27189,N_25015,N_24979);
nand U27190 (N_27190,N_24586,N_24726);
and U27191 (N_27191,N_25458,N_24480);
xnor U27192 (N_27192,N_25119,N_25191);
xor U27193 (N_27193,N_24809,N_25841);
or U27194 (N_27194,N_24963,N_24287);
and U27195 (N_27195,N_24185,N_24742);
and U27196 (N_27196,N_24493,N_25500);
xor U27197 (N_27197,N_24431,N_25530);
nand U27198 (N_27198,N_25173,N_24692);
nor U27199 (N_27199,N_24892,N_25710);
xor U27200 (N_27200,N_25270,N_24038);
and U27201 (N_27201,N_25512,N_24236);
xor U27202 (N_27202,N_25546,N_24526);
nor U27203 (N_27203,N_24353,N_25655);
nor U27204 (N_27204,N_25281,N_25819);
xor U27205 (N_27205,N_24782,N_24397);
or U27206 (N_27206,N_25199,N_24343);
or U27207 (N_27207,N_25992,N_25705);
and U27208 (N_27208,N_24794,N_25512);
xor U27209 (N_27209,N_24010,N_25337);
or U27210 (N_27210,N_25548,N_24048);
nor U27211 (N_27211,N_24598,N_24703);
xnor U27212 (N_27212,N_25176,N_24299);
nand U27213 (N_27213,N_25971,N_24120);
nor U27214 (N_27214,N_25728,N_24809);
and U27215 (N_27215,N_24989,N_24148);
and U27216 (N_27216,N_24494,N_25749);
nand U27217 (N_27217,N_24075,N_25780);
or U27218 (N_27218,N_25065,N_25393);
xnor U27219 (N_27219,N_24607,N_24529);
nand U27220 (N_27220,N_25710,N_24540);
xnor U27221 (N_27221,N_24635,N_25422);
nand U27222 (N_27222,N_25890,N_24376);
or U27223 (N_27223,N_24743,N_24449);
nand U27224 (N_27224,N_24954,N_25211);
xor U27225 (N_27225,N_24686,N_25159);
nand U27226 (N_27226,N_24294,N_24247);
or U27227 (N_27227,N_25273,N_25770);
or U27228 (N_27228,N_25031,N_24811);
and U27229 (N_27229,N_25141,N_25360);
or U27230 (N_27230,N_24875,N_25963);
nand U27231 (N_27231,N_25517,N_25336);
xor U27232 (N_27232,N_24594,N_25676);
and U27233 (N_27233,N_25414,N_25462);
and U27234 (N_27234,N_24145,N_24951);
nor U27235 (N_27235,N_25264,N_24308);
nor U27236 (N_27236,N_24098,N_24838);
and U27237 (N_27237,N_24780,N_24295);
and U27238 (N_27238,N_25190,N_24728);
or U27239 (N_27239,N_24671,N_25071);
xnor U27240 (N_27240,N_24616,N_24571);
nand U27241 (N_27241,N_24596,N_25616);
nor U27242 (N_27242,N_24495,N_24083);
and U27243 (N_27243,N_24935,N_25880);
or U27244 (N_27244,N_25553,N_24614);
xnor U27245 (N_27245,N_25639,N_24468);
or U27246 (N_27246,N_25462,N_25865);
nand U27247 (N_27247,N_24152,N_25133);
and U27248 (N_27248,N_25192,N_24755);
nor U27249 (N_27249,N_24516,N_24896);
xor U27250 (N_27250,N_24564,N_25256);
or U27251 (N_27251,N_24039,N_24199);
or U27252 (N_27252,N_24275,N_24375);
and U27253 (N_27253,N_24266,N_25439);
or U27254 (N_27254,N_25896,N_24694);
and U27255 (N_27255,N_24806,N_24146);
or U27256 (N_27256,N_25985,N_24680);
and U27257 (N_27257,N_24794,N_25713);
and U27258 (N_27258,N_25810,N_24438);
nor U27259 (N_27259,N_24788,N_25069);
nor U27260 (N_27260,N_24965,N_25845);
and U27261 (N_27261,N_24600,N_24379);
nor U27262 (N_27262,N_24408,N_25679);
or U27263 (N_27263,N_25507,N_24876);
nand U27264 (N_27264,N_25340,N_24465);
nand U27265 (N_27265,N_24178,N_25357);
nor U27266 (N_27266,N_24854,N_24114);
and U27267 (N_27267,N_25006,N_24097);
nor U27268 (N_27268,N_24270,N_24532);
and U27269 (N_27269,N_24366,N_24481);
or U27270 (N_27270,N_25712,N_25656);
xnor U27271 (N_27271,N_25134,N_25590);
xnor U27272 (N_27272,N_25758,N_25387);
xor U27273 (N_27273,N_25659,N_24920);
nor U27274 (N_27274,N_24291,N_25339);
nor U27275 (N_27275,N_25479,N_25186);
nor U27276 (N_27276,N_25464,N_25535);
xnor U27277 (N_27277,N_24304,N_24163);
nand U27278 (N_27278,N_24747,N_24959);
and U27279 (N_27279,N_25257,N_25448);
or U27280 (N_27280,N_25651,N_25412);
nor U27281 (N_27281,N_25799,N_24080);
and U27282 (N_27282,N_24624,N_25667);
and U27283 (N_27283,N_24193,N_25101);
and U27284 (N_27284,N_25270,N_25410);
or U27285 (N_27285,N_25209,N_25540);
xnor U27286 (N_27286,N_25499,N_25253);
xnor U27287 (N_27287,N_24815,N_24290);
nor U27288 (N_27288,N_24516,N_25302);
or U27289 (N_27289,N_25570,N_25847);
xnor U27290 (N_27290,N_25999,N_24659);
xnor U27291 (N_27291,N_24649,N_25010);
nand U27292 (N_27292,N_24112,N_25884);
nand U27293 (N_27293,N_24942,N_25540);
or U27294 (N_27294,N_25275,N_24358);
or U27295 (N_27295,N_25020,N_24214);
or U27296 (N_27296,N_25280,N_25956);
or U27297 (N_27297,N_25734,N_25346);
and U27298 (N_27298,N_25847,N_25238);
xnor U27299 (N_27299,N_25122,N_25970);
or U27300 (N_27300,N_25026,N_24679);
or U27301 (N_27301,N_24696,N_25874);
or U27302 (N_27302,N_25647,N_25854);
and U27303 (N_27303,N_24381,N_24710);
nor U27304 (N_27304,N_24609,N_24071);
and U27305 (N_27305,N_24130,N_25619);
and U27306 (N_27306,N_25693,N_24512);
nor U27307 (N_27307,N_24720,N_25843);
and U27308 (N_27308,N_25850,N_24626);
xor U27309 (N_27309,N_24775,N_25279);
nor U27310 (N_27310,N_24984,N_25683);
or U27311 (N_27311,N_25870,N_24258);
or U27312 (N_27312,N_25507,N_24206);
or U27313 (N_27313,N_25358,N_24135);
xor U27314 (N_27314,N_24248,N_24461);
nor U27315 (N_27315,N_24374,N_25067);
nor U27316 (N_27316,N_25881,N_24873);
xor U27317 (N_27317,N_24808,N_24268);
xnor U27318 (N_27318,N_25009,N_25322);
xnor U27319 (N_27319,N_25339,N_25942);
nand U27320 (N_27320,N_24904,N_24244);
and U27321 (N_27321,N_25103,N_25578);
nand U27322 (N_27322,N_24458,N_25941);
nor U27323 (N_27323,N_25565,N_25988);
xnor U27324 (N_27324,N_25468,N_25487);
nor U27325 (N_27325,N_24778,N_25001);
or U27326 (N_27326,N_25115,N_24704);
or U27327 (N_27327,N_25253,N_25928);
nand U27328 (N_27328,N_25671,N_25158);
nor U27329 (N_27329,N_24609,N_24206);
xor U27330 (N_27330,N_24225,N_25990);
nor U27331 (N_27331,N_25553,N_25216);
nor U27332 (N_27332,N_24341,N_25819);
and U27333 (N_27333,N_25913,N_25100);
nand U27334 (N_27334,N_25399,N_25286);
xnor U27335 (N_27335,N_25421,N_24266);
and U27336 (N_27336,N_25291,N_24961);
or U27337 (N_27337,N_24744,N_24361);
nor U27338 (N_27338,N_24376,N_24708);
nor U27339 (N_27339,N_25139,N_24188);
nor U27340 (N_27340,N_24021,N_24612);
or U27341 (N_27341,N_24009,N_24530);
nor U27342 (N_27342,N_24362,N_24326);
nand U27343 (N_27343,N_24183,N_24238);
or U27344 (N_27344,N_24741,N_24643);
nand U27345 (N_27345,N_25276,N_25953);
nor U27346 (N_27346,N_25765,N_25276);
xnor U27347 (N_27347,N_25288,N_25813);
nand U27348 (N_27348,N_25731,N_24184);
nor U27349 (N_27349,N_25210,N_24714);
nor U27350 (N_27350,N_25484,N_25408);
nand U27351 (N_27351,N_25502,N_25054);
nand U27352 (N_27352,N_25214,N_24071);
and U27353 (N_27353,N_25382,N_24243);
and U27354 (N_27354,N_25495,N_24272);
or U27355 (N_27355,N_24136,N_24080);
nor U27356 (N_27356,N_25018,N_24483);
and U27357 (N_27357,N_24097,N_24784);
nor U27358 (N_27358,N_25713,N_25089);
nor U27359 (N_27359,N_24119,N_25139);
or U27360 (N_27360,N_25465,N_24430);
and U27361 (N_27361,N_24614,N_24944);
or U27362 (N_27362,N_25712,N_24050);
or U27363 (N_27363,N_25364,N_24271);
nand U27364 (N_27364,N_25153,N_25958);
xnor U27365 (N_27365,N_25269,N_25688);
nand U27366 (N_27366,N_25596,N_24585);
nand U27367 (N_27367,N_25195,N_25158);
xor U27368 (N_27368,N_25852,N_25521);
xor U27369 (N_27369,N_24667,N_24932);
and U27370 (N_27370,N_24793,N_25160);
nor U27371 (N_27371,N_25370,N_24884);
nand U27372 (N_27372,N_24686,N_24673);
nor U27373 (N_27373,N_25153,N_25477);
nor U27374 (N_27374,N_25818,N_24251);
nand U27375 (N_27375,N_24404,N_24949);
or U27376 (N_27376,N_24290,N_24887);
or U27377 (N_27377,N_24000,N_25811);
and U27378 (N_27378,N_25215,N_25690);
nor U27379 (N_27379,N_24463,N_24772);
and U27380 (N_27380,N_25909,N_25264);
nor U27381 (N_27381,N_25596,N_24379);
and U27382 (N_27382,N_25697,N_25512);
xor U27383 (N_27383,N_25941,N_24826);
and U27384 (N_27384,N_25826,N_25531);
nor U27385 (N_27385,N_25353,N_25274);
xnor U27386 (N_27386,N_24390,N_24323);
or U27387 (N_27387,N_24425,N_25065);
and U27388 (N_27388,N_25314,N_24464);
nand U27389 (N_27389,N_24900,N_24205);
nor U27390 (N_27390,N_25546,N_24633);
nor U27391 (N_27391,N_24255,N_25199);
nand U27392 (N_27392,N_24236,N_24904);
or U27393 (N_27393,N_24658,N_25577);
or U27394 (N_27394,N_24983,N_24333);
nand U27395 (N_27395,N_25796,N_24699);
xor U27396 (N_27396,N_25523,N_25413);
xnor U27397 (N_27397,N_24235,N_24949);
nand U27398 (N_27398,N_24927,N_25018);
xor U27399 (N_27399,N_24624,N_24777);
or U27400 (N_27400,N_24186,N_24618);
and U27401 (N_27401,N_24568,N_24288);
and U27402 (N_27402,N_24076,N_25570);
or U27403 (N_27403,N_25316,N_24211);
nand U27404 (N_27404,N_25805,N_25690);
and U27405 (N_27405,N_25818,N_24635);
or U27406 (N_27406,N_24171,N_24669);
nor U27407 (N_27407,N_25148,N_24960);
xor U27408 (N_27408,N_25814,N_24825);
and U27409 (N_27409,N_25839,N_24724);
xnor U27410 (N_27410,N_24151,N_24262);
and U27411 (N_27411,N_25864,N_24798);
or U27412 (N_27412,N_24229,N_25090);
nor U27413 (N_27413,N_25433,N_24864);
xnor U27414 (N_27414,N_24342,N_25987);
nor U27415 (N_27415,N_24820,N_25502);
xor U27416 (N_27416,N_25290,N_24528);
or U27417 (N_27417,N_25853,N_24634);
and U27418 (N_27418,N_25844,N_24099);
or U27419 (N_27419,N_25881,N_24111);
or U27420 (N_27420,N_25960,N_24942);
nor U27421 (N_27421,N_25562,N_24655);
and U27422 (N_27422,N_25226,N_25783);
nor U27423 (N_27423,N_25071,N_24778);
nor U27424 (N_27424,N_25747,N_25391);
and U27425 (N_27425,N_25545,N_25713);
or U27426 (N_27426,N_25005,N_24756);
or U27427 (N_27427,N_24022,N_24527);
xnor U27428 (N_27428,N_25122,N_25837);
xnor U27429 (N_27429,N_25095,N_24185);
nor U27430 (N_27430,N_25858,N_25489);
and U27431 (N_27431,N_24552,N_24866);
nand U27432 (N_27432,N_25027,N_25432);
nor U27433 (N_27433,N_24935,N_25748);
or U27434 (N_27434,N_24060,N_25887);
nand U27435 (N_27435,N_24628,N_24296);
and U27436 (N_27436,N_24577,N_25402);
nand U27437 (N_27437,N_25553,N_24829);
xnor U27438 (N_27438,N_25523,N_25814);
nand U27439 (N_27439,N_24278,N_24367);
xnor U27440 (N_27440,N_25960,N_24642);
xnor U27441 (N_27441,N_25610,N_25905);
or U27442 (N_27442,N_25605,N_25711);
nor U27443 (N_27443,N_25511,N_24462);
or U27444 (N_27444,N_24722,N_24758);
or U27445 (N_27445,N_25939,N_24503);
or U27446 (N_27446,N_25142,N_25634);
nor U27447 (N_27447,N_24616,N_24726);
nand U27448 (N_27448,N_24379,N_24764);
nor U27449 (N_27449,N_25295,N_24335);
xor U27450 (N_27450,N_24133,N_25531);
nor U27451 (N_27451,N_25200,N_24189);
and U27452 (N_27452,N_25487,N_24851);
and U27453 (N_27453,N_25253,N_25516);
or U27454 (N_27454,N_24735,N_24595);
nand U27455 (N_27455,N_24192,N_24460);
nor U27456 (N_27456,N_24089,N_24604);
or U27457 (N_27457,N_25021,N_24924);
nor U27458 (N_27458,N_24627,N_25148);
xor U27459 (N_27459,N_25566,N_25218);
nand U27460 (N_27460,N_24246,N_25464);
xnor U27461 (N_27461,N_25979,N_24968);
and U27462 (N_27462,N_24945,N_24827);
or U27463 (N_27463,N_25296,N_24616);
nand U27464 (N_27464,N_25448,N_24997);
nor U27465 (N_27465,N_25919,N_24320);
xor U27466 (N_27466,N_24505,N_25392);
or U27467 (N_27467,N_24807,N_25297);
or U27468 (N_27468,N_24686,N_25301);
nand U27469 (N_27469,N_25282,N_25359);
or U27470 (N_27470,N_25684,N_24028);
or U27471 (N_27471,N_25824,N_25374);
nor U27472 (N_27472,N_25841,N_24652);
nand U27473 (N_27473,N_24482,N_24901);
xor U27474 (N_27474,N_24457,N_25229);
nand U27475 (N_27475,N_25471,N_25945);
nor U27476 (N_27476,N_25005,N_25594);
or U27477 (N_27477,N_25645,N_25176);
xnor U27478 (N_27478,N_25235,N_25432);
nor U27479 (N_27479,N_24598,N_25634);
or U27480 (N_27480,N_24168,N_25604);
and U27481 (N_27481,N_24910,N_25042);
and U27482 (N_27482,N_24174,N_24657);
nor U27483 (N_27483,N_25731,N_24229);
xor U27484 (N_27484,N_24784,N_24228);
xor U27485 (N_27485,N_25376,N_24880);
xor U27486 (N_27486,N_25753,N_24297);
xor U27487 (N_27487,N_25315,N_24251);
nor U27488 (N_27488,N_25750,N_24331);
nand U27489 (N_27489,N_24441,N_24684);
nand U27490 (N_27490,N_25853,N_25902);
nand U27491 (N_27491,N_24443,N_25271);
xnor U27492 (N_27492,N_25942,N_25194);
nor U27493 (N_27493,N_25784,N_25767);
nor U27494 (N_27494,N_25138,N_24136);
nor U27495 (N_27495,N_24025,N_24273);
and U27496 (N_27496,N_24130,N_25023);
xor U27497 (N_27497,N_24702,N_24693);
nand U27498 (N_27498,N_25019,N_25182);
nand U27499 (N_27499,N_25573,N_24710);
nor U27500 (N_27500,N_24066,N_25823);
or U27501 (N_27501,N_25938,N_24051);
nor U27502 (N_27502,N_25246,N_25948);
nor U27503 (N_27503,N_25931,N_25582);
or U27504 (N_27504,N_25755,N_24134);
and U27505 (N_27505,N_24769,N_24703);
or U27506 (N_27506,N_25336,N_25003);
and U27507 (N_27507,N_24379,N_24003);
or U27508 (N_27508,N_25777,N_24207);
nand U27509 (N_27509,N_24457,N_25405);
or U27510 (N_27510,N_24487,N_25056);
nand U27511 (N_27511,N_25446,N_25913);
xnor U27512 (N_27512,N_25111,N_25392);
nand U27513 (N_27513,N_25682,N_25947);
and U27514 (N_27514,N_24382,N_25344);
nor U27515 (N_27515,N_25321,N_25299);
xor U27516 (N_27516,N_25960,N_24906);
or U27517 (N_27517,N_24780,N_24187);
nand U27518 (N_27518,N_24088,N_25833);
nor U27519 (N_27519,N_24187,N_25734);
nor U27520 (N_27520,N_25432,N_25487);
nand U27521 (N_27521,N_24546,N_25946);
or U27522 (N_27522,N_25628,N_24178);
and U27523 (N_27523,N_25792,N_24588);
and U27524 (N_27524,N_25413,N_25507);
xnor U27525 (N_27525,N_25636,N_24270);
or U27526 (N_27526,N_24325,N_25424);
or U27527 (N_27527,N_25420,N_24164);
xor U27528 (N_27528,N_25429,N_25378);
nand U27529 (N_27529,N_25999,N_25245);
or U27530 (N_27530,N_25470,N_24119);
nor U27531 (N_27531,N_25739,N_24203);
nand U27532 (N_27532,N_25257,N_25485);
xor U27533 (N_27533,N_24604,N_24091);
nand U27534 (N_27534,N_25794,N_24990);
and U27535 (N_27535,N_24582,N_25255);
nand U27536 (N_27536,N_24756,N_24776);
xnor U27537 (N_27537,N_25527,N_25089);
nor U27538 (N_27538,N_25404,N_25304);
and U27539 (N_27539,N_25686,N_24147);
nand U27540 (N_27540,N_25290,N_24006);
nand U27541 (N_27541,N_24598,N_24204);
nor U27542 (N_27542,N_25656,N_25852);
or U27543 (N_27543,N_25142,N_25178);
and U27544 (N_27544,N_24524,N_25366);
nor U27545 (N_27545,N_25194,N_25441);
nand U27546 (N_27546,N_24996,N_24820);
or U27547 (N_27547,N_25364,N_24456);
and U27548 (N_27548,N_25750,N_24994);
or U27549 (N_27549,N_24122,N_24273);
nor U27550 (N_27550,N_24343,N_24039);
or U27551 (N_27551,N_25598,N_24816);
xnor U27552 (N_27552,N_24386,N_25179);
xor U27553 (N_27553,N_24831,N_24729);
nor U27554 (N_27554,N_24986,N_24841);
xor U27555 (N_27555,N_24231,N_24495);
or U27556 (N_27556,N_25631,N_24483);
xor U27557 (N_27557,N_24749,N_24513);
nand U27558 (N_27558,N_24934,N_24964);
and U27559 (N_27559,N_25375,N_25235);
and U27560 (N_27560,N_24159,N_25177);
xnor U27561 (N_27561,N_24849,N_25052);
nand U27562 (N_27562,N_24669,N_25184);
nor U27563 (N_27563,N_25572,N_25292);
and U27564 (N_27564,N_24359,N_24067);
nand U27565 (N_27565,N_25491,N_24273);
nor U27566 (N_27566,N_24741,N_24067);
xor U27567 (N_27567,N_24633,N_25329);
xnor U27568 (N_27568,N_24356,N_25582);
and U27569 (N_27569,N_24309,N_25213);
xnor U27570 (N_27570,N_25547,N_24866);
or U27571 (N_27571,N_24546,N_24181);
nand U27572 (N_27572,N_25972,N_25715);
and U27573 (N_27573,N_24332,N_25379);
xor U27574 (N_27574,N_24957,N_25965);
and U27575 (N_27575,N_24484,N_25897);
or U27576 (N_27576,N_24220,N_24805);
or U27577 (N_27577,N_24862,N_25661);
nor U27578 (N_27578,N_24940,N_24749);
nand U27579 (N_27579,N_24242,N_25084);
xnor U27580 (N_27580,N_25783,N_25674);
and U27581 (N_27581,N_25876,N_24731);
nor U27582 (N_27582,N_25698,N_24354);
nand U27583 (N_27583,N_24865,N_24867);
nand U27584 (N_27584,N_25911,N_24937);
nor U27585 (N_27585,N_25844,N_25100);
nand U27586 (N_27586,N_24291,N_25721);
nand U27587 (N_27587,N_25720,N_25499);
xnor U27588 (N_27588,N_25356,N_24492);
and U27589 (N_27589,N_24099,N_24419);
nand U27590 (N_27590,N_24039,N_24427);
xnor U27591 (N_27591,N_24281,N_25220);
nand U27592 (N_27592,N_25432,N_24580);
xnor U27593 (N_27593,N_24768,N_24988);
xnor U27594 (N_27594,N_24943,N_25926);
xnor U27595 (N_27595,N_24042,N_24657);
nor U27596 (N_27596,N_25489,N_25333);
and U27597 (N_27597,N_24039,N_24857);
nor U27598 (N_27598,N_24881,N_24257);
and U27599 (N_27599,N_25809,N_24169);
nor U27600 (N_27600,N_25820,N_25865);
and U27601 (N_27601,N_25702,N_24693);
and U27602 (N_27602,N_25660,N_24950);
nor U27603 (N_27603,N_25928,N_24098);
nor U27604 (N_27604,N_24930,N_25854);
nand U27605 (N_27605,N_24358,N_24228);
xnor U27606 (N_27606,N_24629,N_24478);
or U27607 (N_27607,N_24691,N_24407);
or U27608 (N_27608,N_24443,N_25287);
nor U27609 (N_27609,N_24904,N_25122);
nand U27610 (N_27610,N_24208,N_24969);
nand U27611 (N_27611,N_24605,N_25434);
and U27612 (N_27612,N_25422,N_24642);
xor U27613 (N_27613,N_24195,N_24278);
nor U27614 (N_27614,N_24930,N_25611);
nor U27615 (N_27615,N_24855,N_25287);
xor U27616 (N_27616,N_24868,N_24100);
xnor U27617 (N_27617,N_25576,N_25589);
xor U27618 (N_27618,N_24071,N_25232);
xnor U27619 (N_27619,N_24059,N_24489);
or U27620 (N_27620,N_24607,N_25214);
nand U27621 (N_27621,N_25722,N_25190);
nand U27622 (N_27622,N_25100,N_24702);
nor U27623 (N_27623,N_25560,N_24870);
xor U27624 (N_27624,N_25889,N_25466);
xnor U27625 (N_27625,N_24205,N_25548);
or U27626 (N_27626,N_24830,N_25051);
nor U27627 (N_27627,N_24139,N_24083);
nand U27628 (N_27628,N_25374,N_25802);
nor U27629 (N_27629,N_24978,N_24715);
or U27630 (N_27630,N_25314,N_25390);
nand U27631 (N_27631,N_25619,N_25378);
and U27632 (N_27632,N_24310,N_25001);
and U27633 (N_27633,N_25613,N_25818);
xor U27634 (N_27634,N_25760,N_25477);
or U27635 (N_27635,N_24648,N_25320);
nor U27636 (N_27636,N_25010,N_25866);
and U27637 (N_27637,N_24055,N_25952);
xnor U27638 (N_27638,N_25057,N_24199);
or U27639 (N_27639,N_25879,N_25349);
and U27640 (N_27640,N_25090,N_25385);
or U27641 (N_27641,N_25990,N_24348);
nor U27642 (N_27642,N_25363,N_24413);
xnor U27643 (N_27643,N_24682,N_24191);
nand U27644 (N_27644,N_25077,N_24442);
nor U27645 (N_27645,N_24420,N_25347);
nand U27646 (N_27646,N_25933,N_24244);
or U27647 (N_27647,N_24027,N_24870);
nand U27648 (N_27648,N_24130,N_24686);
or U27649 (N_27649,N_24301,N_25522);
nand U27650 (N_27650,N_24231,N_25040);
and U27651 (N_27651,N_25247,N_24054);
or U27652 (N_27652,N_25768,N_24065);
or U27653 (N_27653,N_25656,N_25847);
nand U27654 (N_27654,N_25829,N_25848);
nand U27655 (N_27655,N_25794,N_25596);
xnor U27656 (N_27656,N_24501,N_24565);
and U27657 (N_27657,N_24979,N_25562);
nand U27658 (N_27658,N_25527,N_24485);
nand U27659 (N_27659,N_25848,N_25124);
and U27660 (N_27660,N_24924,N_25915);
or U27661 (N_27661,N_24945,N_25590);
xnor U27662 (N_27662,N_25532,N_24786);
xor U27663 (N_27663,N_25109,N_24930);
xnor U27664 (N_27664,N_24641,N_25631);
nand U27665 (N_27665,N_24029,N_24539);
and U27666 (N_27666,N_24295,N_25912);
or U27667 (N_27667,N_24599,N_25265);
and U27668 (N_27668,N_24230,N_24284);
xor U27669 (N_27669,N_25275,N_24924);
nand U27670 (N_27670,N_25379,N_24941);
or U27671 (N_27671,N_25074,N_24758);
nand U27672 (N_27672,N_25346,N_25680);
and U27673 (N_27673,N_24601,N_24753);
nand U27674 (N_27674,N_25441,N_24065);
xnor U27675 (N_27675,N_25171,N_25925);
nand U27676 (N_27676,N_25769,N_24964);
nand U27677 (N_27677,N_24753,N_24710);
nor U27678 (N_27678,N_25462,N_25712);
and U27679 (N_27679,N_24269,N_25893);
nand U27680 (N_27680,N_25527,N_24783);
nand U27681 (N_27681,N_24425,N_24617);
xnor U27682 (N_27682,N_24598,N_25320);
and U27683 (N_27683,N_24322,N_24405);
and U27684 (N_27684,N_25277,N_24369);
and U27685 (N_27685,N_24838,N_25366);
nand U27686 (N_27686,N_24862,N_24002);
nor U27687 (N_27687,N_25039,N_24448);
nand U27688 (N_27688,N_25338,N_25637);
xnor U27689 (N_27689,N_24360,N_24324);
nand U27690 (N_27690,N_24096,N_25254);
xnor U27691 (N_27691,N_25387,N_25744);
nand U27692 (N_27692,N_25820,N_24569);
xor U27693 (N_27693,N_25900,N_25429);
or U27694 (N_27694,N_25852,N_25999);
nand U27695 (N_27695,N_25544,N_24317);
nand U27696 (N_27696,N_25938,N_24292);
nor U27697 (N_27697,N_24757,N_25147);
and U27698 (N_27698,N_24520,N_25561);
nand U27699 (N_27699,N_25762,N_25536);
or U27700 (N_27700,N_25970,N_24510);
nor U27701 (N_27701,N_24576,N_25966);
nor U27702 (N_27702,N_24520,N_24131);
and U27703 (N_27703,N_24066,N_25785);
nand U27704 (N_27704,N_25677,N_25299);
xnor U27705 (N_27705,N_25617,N_25570);
and U27706 (N_27706,N_25406,N_25759);
xor U27707 (N_27707,N_24530,N_24327);
or U27708 (N_27708,N_25246,N_24480);
xnor U27709 (N_27709,N_24181,N_24523);
or U27710 (N_27710,N_25043,N_24406);
and U27711 (N_27711,N_24111,N_24443);
or U27712 (N_27712,N_25454,N_25157);
or U27713 (N_27713,N_25319,N_25084);
xor U27714 (N_27714,N_25777,N_25805);
or U27715 (N_27715,N_25633,N_25429);
and U27716 (N_27716,N_24418,N_24921);
nor U27717 (N_27717,N_24760,N_25414);
nand U27718 (N_27718,N_24879,N_25055);
nand U27719 (N_27719,N_25138,N_24479);
or U27720 (N_27720,N_25500,N_25115);
and U27721 (N_27721,N_25977,N_25281);
and U27722 (N_27722,N_25728,N_25155);
nor U27723 (N_27723,N_25529,N_25726);
nand U27724 (N_27724,N_24549,N_25552);
nor U27725 (N_27725,N_25418,N_24608);
xor U27726 (N_27726,N_25320,N_24480);
nand U27727 (N_27727,N_24211,N_24184);
and U27728 (N_27728,N_24235,N_24577);
nand U27729 (N_27729,N_24964,N_24977);
and U27730 (N_27730,N_24130,N_25066);
xnor U27731 (N_27731,N_24170,N_25367);
nand U27732 (N_27732,N_24601,N_25148);
nor U27733 (N_27733,N_24972,N_25162);
nand U27734 (N_27734,N_25051,N_25403);
nor U27735 (N_27735,N_25047,N_25440);
nand U27736 (N_27736,N_25981,N_25023);
nor U27737 (N_27737,N_24419,N_24638);
xor U27738 (N_27738,N_24563,N_25203);
or U27739 (N_27739,N_25128,N_25122);
or U27740 (N_27740,N_25686,N_24001);
xnor U27741 (N_27741,N_25676,N_24466);
xnor U27742 (N_27742,N_25721,N_24635);
nand U27743 (N_27743,N_24704,N_24766);
or U27744 (N_27744,N_25639,N_25685);
and U27745 (N_27745,N_24648,N_24106);
nor U27746 (N_27746,N_24026,N_24132);
xnor U27747 (N_27747,N_24616,N_24108);
nor U27748 (N_27748,N_25274,N_24211);
xnor U27749 (N_27749,N_25001,N_25253);
nand U27750 (N_27750,N_24489,N_24563);
or U27751 (N_27751,N_24643,N_25489);
and U27752 (N_27752,N_24860,N_24419);
and U27753 (N_27753,N_24411,N_24485);
or U27754 (N_27754,N_24291,N_25252);
and U27755 (N_27755,N_25289,N_25439);
xor U27756 (N_27756,N_24377,N_24757);
and U27757 (N_27757,N_25552,N_25424);
nor U27758 (N_27758,N_24777,N_24425);
nor U27759 (N_27759,N_24186,N_25290);
nand U27760 (N_27760,N_25188,N_25991);
and U27761 (N_27761,N_25923,N_25955);
and U27762 (N_27762,N_25477,N_25546);
or U27763 (N_27763,N_24870,N_25832);
nand U27764 (N_27764,N_24059,N_24877);
or U27765 (N_27765,N_24482,N_24699);
or U27766 (N_27766,N_25824,N_24145);
xor U27767 (N_27767,N_25514,N_25016);
nand U27768 (N_27768,N_24039,N_24699);
and U27769 (N_27769,N_25204,N_25925);
nand U27770 (N_27770,N_24023,N_25054);
or U27771 (N_27771,N_24605,N_24340);
and U27772 (N_27772,N_24591,N_24610);
nand U27773 (N_27773,N_24051,N_25958);
and U27774 (N_27774,N_24098,N_24074);
or U27775 (N_27775,N_25830,N_25254);
or U27776 (N_27776,N_25868,N_25156);
and U27777 (N_27777,N_24317,N_25590);
nand U27778 (N_27778,N_25259,N_24013);
nor U27779 (N_27779,N_25358,N_24470);
and U27780 (N_27780,N_24956,N_24641);
xnor U27781 (N_27781,N_24659,N_25403);
nand U27782 (N_27782,N_25813,N_24662);
nand U27783 (N_27783,N_24322,N_25765);
nor U27784 (N_27784,N_24450,N_24004);
nor U27785 (N_27785,N_24778,N_24483);
and U27786 (N_27786,N_25251,N_24535);
or U27787 (N_27787,N_25121,N_24144);
xnor U27788 (N_27788,N_24958,N_24953);
or U27789 (N_27789,N_25931,N_25461);
and U27790 (N_27790,N_24307,N_24560);
nor U27791 (N_27791,N_24845,N_24686);
or U27792 (N_27792,N_24859,N_24657);
xnor U27793 (N_27793,N_25460,N_24024);
or U27794 (N_27794,N_24707,N_25386);
xor U27795 (N_27795,N_25815,N_24136);
and U27796 (N_27796,N_25658,N_24585);
or U27797 (N_27797,N_24355,N_24298);
nor U27798 (N_27798,N_24610,N_25289);
or U27799 (N_27799,N_25546,N_25459);
or U27800 (N_27800,N_24239,N_24249);
and U27801 (N_27801,N_25492,N_25132);
nand U27802 (N_27802,N_25533,N_25663);
or U27803 (N_27803,N_25252,N_24109);
nand U27804 (N_27804,N_25271,N_25384);
or U27805 (N_27805,N_24502,N_24099);
and U27806 (N_27806,N_24676,N_25206);
xnor U27807 (N_27807,N_25588,N_24399);
or U27808 (N_27808,N_24478,N_24503);
nand U27809 (N_27809,N_24360,N_24471);
xor U27810 (N_27810,N_24243,N_25008);
nor U27811 (N_27811,N_24404,N_25684);
nor U27812 (N_27812,N_25052,N_25360);
nand U27813 (N_27813,N_24074,N_25824);
and U27814 (N_27814,N_24864,N_25400);
or U27815 (N_27815,N_24927,N_25474);
nand U27816 (N_27816,N_25787,N_25280);
nand U27817 (N_27817,N_24243,N_24897);
or U27818 (N_27818,N_24093,N_24942);
or U27819 (N_27819,N_24194,N_24425);
and U27820 (N_27820,N_24104,N_24400);
nor U27821 (N_27821,N_25181,N_25215);
nand U27822 (N_27822,N_25906,N_24803);
and U27823 (N_27823,N_25536,N_24704);
nor U27824 (N_27824,N_25519,N_25838);
xor U27825 (N_27825,N_25183,N_25512);
nor U27826 (N_27826,N_24638,N_25985);
and U27827 (N_27827,N_25990,N_24830);
nand U27828 (N_27828,N_25442,N_24371);
and U27829 (N_27829,N_24883,N_24338);
nor U27830 (N_27830,N_25572,N_25619);
xnor U27831 (N_27831,N_24883,N_24475);
and U27832 (N_27832,N_24763,N_24845);
and U27833 (N_27833,N_25300,N_24576);
nand U27834 (N_27834,N_24522,N_24455);
or U27835 (N_27835,N_25268,N_24165);
xnor U27836 (N_27836,N_24590,N_24482);
nor U27837 (N_27837,N_25486,N_25975);
and U27838 (N_27838,N_24813,N_25552);
nand U27839 (N_27839,N_24153,N_24490);
nor U27840 (N_27840,N_24598,N_25965);
nand U27841 (N_27841,N_25028,N_24284);
or U27842 (N_27842,N_24301,N_25349);
nor U27843 (N_27843,N_24146,N_24457);
xor U27844 (N_27844,N_24662,N_25000);
xor U27845 (N_27845,N_24503,N_24149);
or U27846 (N_27846,N_25546,N_24338);
nand U27847 (N_27847,N_25973,N_25579);
xnor U27848 (N_27848,N_25399,N_24136);
xor U27849 (N_27849,N_25861,N_25432);
nand U27850 (N_27850,N_25786,N_25886);
nor U27851 (N_27851,N_24748,N_24675);
nor U27852 (N_27852,N_24103,N_25593);
or U27853 (N_27853,N_24850,N_24449);
and U27854 (N_27854,N_24557,N_25592);
nand U27855 (N_27855,N_24398,N_25375);
and U27856 (N_27856,N_25637,N_25040);
and U27857 (N_27857,N_24659,N_25856);
or U27858 (N_27858,N_24809,N_25874);
nor U27859 (N_27859,N_24220,N_25161);
nand U27860 (N_27860,N_25378,N_24461);
or U27861 (N_27861,N_25132,N_24496);
nor U27862 (N_27862,N_25240,N_25862);
nor U27863 (N_27863,N_25768,N_25756);
and U27864 (N_27864,N_24103,N_25912);
and U27865 (N_27865,N_25829,N_25168);
xnor U27866 (N_27866,N_24787,N_25340);
nand U27867 (N_27867,N_24651,N_24318);
nand U27868 (N_27868,N_25834,N_24558);
and U27869 (N_27869,N_25764,N_25441);
xnor U27870 (N_27870,N_25995,N_25558);
and U27871 (N_27871,N_25139,N_24176);
nand U27872 (N_27872,N_24587,N_24786);
nand U27873 (N_27873,N_25355,N_25089);
xnor U27874 (N_27874,N_25807,N_25669);
nor U27875 (N_27875,N_24739,N_24807);
xor U27876 (N_27876,N_24300,N_24640);
and U27877 (N_27877,N_25555,N_25956);
or U27878 (N_27878,N_25486,N_25149);
xor U27879 (N_27879,N_24980,N_24015);
nand U27880 (N_27880,N_24752,N_25717);
or U27881 (N_27881,N_24762,N_24012);
nand U27882 (N_27882,N_24405,N_25030);
nand U27883 (N_27883,N_24133,N_24280);
or U27884 (N_27884,N_24815,N_24098);
xnor U27885 (N_27885,N_24915,N_24509);
nand U27886 (N_27886,N_25946,N_25658);
xor U27887 (N_27887,N_24955,N_24322);
xor U27888 (N_27888,N_24416,N_24115);
nand U27889 (N_27889,N_24838,N_24324);
nand U27890 (N_27890,N_25827,N_24626);
and U27891 (N_27891,N_25501,N_25503);
nor U27892 (N_27892,N_25762,N_25940);
nor U27893 (N_27893,N_24727,N_25872);
nand U27894 (N_27894,N_24693,N_25744);
nand U27895 (N_27895,N_24982,N_24489);
nand U27896 (N_27896,N_24728,N_25969);
nor U27897 (N_27897,N_24454,N_24511);
nor U27898 (N_27898,N_24346,N_24105);
nor U27899 (N_27899,N_25552,N_25272);
or U27900 (N_27900,N_24464,N_25408);
xor U27901 (N_27901,N_24841,N_25579);
xnor U27902 (N_27902,N_25265,N_24235);
and U27903 (N_27903,N_25528,N_25272);
nor U27904 (N_27904,N_24814,N_25797);
nor U27905 (N_27905,N_24206,N_24968);
nor U27906 (N_27906,N_25711,N_25820);
xor U27907 (N_27907,N_24057,N_25745);
and U27908 (N_27908,N_25308,N_25541);
nor U27909 (N_27909,N_25384,N_25292);
or U27910 (N_27910,N_25244,N_24979);
or U27911 (N_27911,N_25886,N_24754);
xor U27912 (N_27912,N_25704,N_24652);
nand U27913 (N_27913,N_25663,N_24392);
and U27914 (N_27914,N_24582,N_25729);
xnor U27915 (N_27915,N_25264,N_25752);
nor U27916 (N_27916,N_24768,N_25213);
or U27917 (N_27917,N_24680,N_24252);
nand U27918 (N_27918,N_25030,N_24513);
and U27919 (N_27919,N_25916,N_25257);
nand U27920 (N_27920,N_24480,N_25445);
or U27921 (N_27921,N_24062,N_25424);
nor U27922 (N_27922,N_24548,N_25973);
and U27923 (N_27923,N_25923,N_25483);
and U27924 (N_27924,N_25974,N_24931);
xnor U27925 (N_27925,N_24784,N_24206);
nand U27926 (N_27926,N_24964,N_24226);
nand U27927 (N_27927,N_24335,N_25017);
nand U27928 (N_27928,N_24414,N_25538);
nor U27929 (N_27929,N_24376,N_25388);
and U27930 (N_27930,N_25690,N_25218);
nand U27931 (N_27931,N_24292,N_25775);
or U27932 (N_27932,N_24964,N_24104);
nand U27933 (N_27933,N_24429,N_25272);
xor U27934 (N_27934,N_25008,N_24292);
nand U27935 (N_27935,N_24007,N_24504);
nor U27936 (N_27936,N_24574,N_25689);
xor U27937 (N_27937,N_25605,N_24738);
and U27938 (N_27938,N_24451,N_25163);
and U27939 (N_27939,N_24918,N_25239);
xor U27940 (N_27940,N_25465,N_25559);
xor U27941 (N_27941,N_25093,N_25176);
nand U27942 (N_27942,N_25522,N_25379);
or U27943 (N_27943,N_24749,N_24329);
and U27944 (N_27944,N_25711,N_24795);
xor U27945 (N_27945,N_25276,N_24991);
or U27946 (N_27946,N_25701,N_25860);
or U27947 (N_27947,N_24692,N_24201);
and U27948 (N_27948,N_25941,N_24967);
and U27949 (N_27949,N_24601,N_25343);
nand U27950 (N_27950,N_24778,N_25374);
or U27951 (N_27951,N_24814,N_25944);
xor U27952 (N_27952,N_24791,N_24386);
nand U27953 (N_27953,N_25524,N_25253);
nor U27954 (N_27954,N_25807,N_24659);
nand U27955 (N_27955,N_25196,N_24788);
xnor U27956 (N_27956,N_25510,N_24973);
nor U27957 (N_27957,N_25011,N_24261);
xnor U27958 (N_27958,N_24623,N_24209);
nand U27959 (N_27959,N_24675,N_24117);
xor U27960 (N_27960,N_25019,N_25488);
nor U27961 (N_27961,N_24435,N_25821);
nor U27962 (N_27962,N_24484,N_25517);
or U27963 (N_27963,N_24675,N_25483);
nor U27964 (N_27964,N_24331,N_25974);
or U27965 (N_27965,N_25790,N_24238);
xor U27966 (N_27966,N_25927,N_25324);
nand U27967 (N_27967,N_25107,N_25928);
nand U27968 (N_27968,N_25444,N_25682);
xor U27969 (N_27969,N_24139,N_25078);
nand U27970 (N_27970,N_25966,N_24958);
and U27971 (N_27971,N_25240,N_24308);
nor U27972 (N_27972,N_25249,N_25482);
and U27973 (N_27973,N_24491,N_24450);
and U27974 (N_27974,N_24501,N_24684);
nand U27975 (N_27975,N_24784,N_25988);
and U27976 (N_27976,N_25472,N_25339);
and U27977 (N_27977,N_24735,N_25462);
and U27978 (N_27978,N_25276,N_25679);
nand U27979 (N_27979,N_25428,N_25171);
xnor U27980 (N_27980,N_24811,N_24936);
or U27981 (N_27981,N_24459,N_25428);
or U27982 (N_27982,N_25700,N_24850);
nand U27983 (N_27983,N_24998,N_24066);
nor U27984 (N_27984,N_24822,N_24804);
nor U27985 (N_27985,N_25473,N_25942);
and U27986 (N_27986,N_25001,N_24135);
nand U27987 (N_27987,N_24266,N_25002);
and U27988 (N_27988,N_25679,N_25306);
and U27989 (N_27989,N_25877,N_25730);
nor U27990 (N_27990,N_24698,N_24167);
nor U27991 (N_27991,N_24003,N_25444);
and U27992 (N_27992,N_25922,N_25241);
xor U27993 (N_27993,N_24706,N_24452);
nor U27994 (N_27994,N_24211,N_25221);
nor U27995 (N_27995,N_25949,N_24985);
and U27996 (N_27996,N_25748,N_25871);
or U27997 (N_27997,N_24731,N_25417);
xor U27998 (N_27998,N_24845,N_24814);
nand U27999 (N_27999,N_24292,N_25602);
and U28000 (N_28000,N_26002,N_26723);
nor U28001 (N_28001,N_27460,N_26300);
xor U28002 (N_28002,N_26001,N_27702);
or U28003 (N_28003,N_26232,N_27581);
nand U28004 (N_28004,N_27769,N_27259);
nor U28005 (N_28005,N_26456,N_27246);
xor U28006 (N_28006,N_27306,N_27607);
and U28007 (N_28007,N_26139,N_26124);
nor U28008 (N_28008,N_26432,N_27036);
and U28009 (N_28009,N_27450,N_27600);
or U28010 (N_28010,N_26993,N_26659);
or U28011 (N_28011,N_27426,N_27632);
and U28012 (N_28012,N_27993,N_27336);
or U28013 (N_28013,N_27350,N_26868);
and U28014 (N_28014,N_26441,N_26648);
nand U28015 (N_28015,N_27152,N_27179);
nor U28016 (N_28016,N_26748,N_27810);
nand U28017 (N_28017,N_27269,N_26818);
or U28018 (N_28018,N_27733,N_26419);
and U28019 (N_28019,N_27054,N_27750);
nor U28020 (N_28020,N_26435,N_27801);
or U28021 (N_28021,N_27550,N_26813);
or U28022 (N_28022,N_26514,N_26422);
and U28023 (N_28023,N_26222,N_26530);
or U28024 (N_28024,N_26628,N_26753);
and U28025 (N_28025,N_26814,N_27793);
or U28026 (N_28026,N_26663,N_26021);
nand U28027 (N_28027,N_27680,N_27310);
xor U28028 (N_28028,N_26239,N_26815);
nor U28029 (N_28029,N_27156,N_27099);
or U28030 (N_28030,N_27820,N_27176);
or U28031 (N_28031,N_26086,N_26368);
xnor U28032 (N_28032,N_26824,N_26972);
nand U28033 (N_28033,N_26590,N_26043);
or U28034 (N_28034,N_27083,N_26639);
nor U28035 (N_28035,N_27468,N_26897);
and U28036 (N_28036,N_27977,N_27797);
nor U28037 (N_28037,N_26477,N_26496);
and U28038 (N_28038,N_27656,N_27491);
and U28039 (N_28039,N_26837,N_27493);
nor U28040 (N_28040,N_27481,N_26725);
nand U28041 (N_28041,N_26333,N_27606);
or U28042 (N_28042,N_26090,N_27631);
nand U28043 (N_28043,N_26073,N_26796);
and U28044 (N_28044,N_27235,N_27761);
nor U28045 (N_28045,N_27257,N_27311);
or U28046 (N_28046,N_26069,N_27555);
or U28047 (N_28047,N_27519,N_26855);
xnor U28048 (N_28048,N_27670,N_26510);
or U28049 (N_28049,N_27159,N_26996);
nor U28050 (N_28050,N_26076,N_26495);
or U28051 (N_28051,N_26729,N_26110);
xnor U28052 (N_28052,N_26632,N_27704);
xnor U28053 (N_28053,N_26025,N_27173);
nand U28054 (N_28054,N_27939,N_27330);
nand U28055 (N_28055,N_26873,N_26889);
xor U28056 (N_28056,N_26224,N_26871);
nor U28057 (N_28057,N_27506,N_27160);
or U28058 (N_28058,N_26625,N_26079);
nand U28059 (N_28059,N_26627,N_26497);
or U28060 (N_28060,N_27128,N_26881);
nor U28061 (N_28061,N_26511,N_26061);
or U28062 (N_28062,N_27957,N_27539);
xor U28063 (N_28063,N_27024,N_27105);
nor U28064 (N_28064,N_26665,N_27279);
xnor U28065 (N_28065,N_27917,N_26760);
nand U28066 (N_28066,N_26759,N_26281);
xor U28067 (N_28067,N_27467,N_27821);
nor U28068 (N_28068,N_26391,N_27743);
or U28069 (N_28069,N_26971,N_26077);
nand U28070 (N_28070,N_26877,N_27015);
or U28071 (N_28071,N_27287,N_27211);
nor U28072 (N_28072,N_26415,N_26087);
nand U28073 (N_28073,N_27465,N_27853);
nand U28074 (N_28074,N_27513,N_27408);
xor U28075 (N_28075,N_27647,N_27583);
nor U28076 (N_28076,N_27446,N_27904);
xnor U28077 (N_28077,N_27348,N_26902);
nand U28078 (N_28078,N_27428,N_26927);
nand U28079 (N_28079,N_27948,N_27209);
or U28080 (N_28080,N_26849,N_26772);
nor U28081 (N_28081,N_27574,N_26265);
xor U28082 (N_28082,N_27031,N_27537);
or U28083 (N_28083,N_26646,N_26502);
xnor U28084 (N_28084,N_27392,N_27046);
xnor U28085 (N_28085,N_27003,N_26517);
xnor U28086 (N_28086,N_26214,N_27556);
nand U28087 (N_28087,N_26385,N_26817);
xnor U28088 (N_28088,N_26982,N_27057);
or U28089 (N_28089,N_27065,N_26722);
or U28090 (N_28090,N_26893,N_27930);
nor U28091 (N_28091,N_26440,N_27849);
xnor U28092 (N_28092,N_26852,N_27261);
or U28093 (N_28093,N_26997,N_27882);
nand U28094 (N_28094,N_27742,N_27962);
and U28095 (N_28095,N_27241,N_26520);
xnor U28096 (N_28096,N_26460,N_27997);
nor U28097 (N_28097,N_26991,N_27946);
xnor U28098 (N_28098,N_27123,N_26567);
nand U28099 (N_28099,N_27779,N_26121);
and U28100 (N_28100,N_27839,N_27367);
xor U28101 (N_28101,N_27870,N_27207);
or U28102 (N_28102,N_26149,N_27604);
nand U28103 (N_28103,N_27869,N_27421);
or U28104 (N_28104,N_27187,N_27996);
nand U28105 (N_28105,N_26324,N_26271);
xor U28106 (N_28106,N_26943,N_27775);
nor U28107 (N_28107,N_27949,N_27404);
nor U28108 (N_28108,N_26891,N_26689);
xor U28109 (N_28109,N_26907,N_27541);
xnor U28110 (N_28110,N_27780,N_26336);
and U28111 (N_28111,N_26133,N_27738);
nor U28112 (N_28112,N_26490,N_27872);
xor U28113 (N_28113,N_27458,N_27055);
nor U28114 (N_28114,N_26346,N_27273);
and U28115 (N_28115,N_26535,N_27329);
nand U28116 (N_28116,N_26500,N_26052);
or U28117 (N_28117,N_26155,N_27039);
nand U28118 (N_28118,N_27825,N_26251);
or U28119 (N_28119,N_27077,N_26105);
xnor U28120 (N_28120,N_27407,N_26706);
xor U28121 (N_28121,N_27220,N_26842);
nand U28122 (N_28122,N_27727,N_27682);
nor U28123 (N_28123,N_27700,N_26274);
nand U28124 (N_28124,N_26186,N_26680);
nor U28125 (N_28125,N_27131,N_27636);
xor U28126 (N_28126,N_27461,N_27358);
or U28127 (N_28127,N_26541,N_27444);
or U28128 (N_28128,N_26505,N_27618);
nor U28129 (N_28129,N_26778,N_26499);
and U28130 (N_28130,N_27856,N_27238);
nor U28131 (N_28131,N_27122,N_26207);
xnor U28132 (N_28132,N_27121,N_27963);
nand U28133 (N_28133,N_26790,N_27877);
and U28134 (N_28134,N_26461,N_27956);
nand U28135 (N_28135,N_26801,N_27755);
and U28136 (N_28136,N_26252,N_27169);
and U28137 (N_28137,N_27371,N_26995);
xor U28138 (N_28138,N_26137,N_27067);
xor U28139 (N_28139,N_26075,N_27756);
nor U28140 (N_28140,N_27717,N_27794);
or U28141 (N_28141,N_26565,N_26536);
xor U28142 (N_28142,N_27454,N_27705);
and U28143 (N_28143,N_27014,N_27901);
nor U28144 (N_28144,N_26476,N_26805);
or U28145 (N_28145,N_27085,N_27703);
or U28146 (N_28146,N_26939,N_26766);
xnor U28147 (N_28147,N_27546,N_27969);
xnor U28148 (N_28148,N_27594,N_26914);
or U28149 (N_28149,N_27579,N_26529);
nand U28150 (N_28150,N_26594,N_26808);
nand U28151 (N_28151,N_27130,N_26022);
and U28152 (N_28152,N_26050,N_26679);
xnor U28153 (N_28153,N_27192,N_26080);
xor U28154 (N_28154,N_26373,N_26491);
and U28155 (N_28155,N_26000,N_27955);
or U28156 (N_28156,N_27406,N_27759);
nand U28157 (N_28157,N_26283,N_27573);
and U28158 (N_28158,N_27712,N_27208);
xnor U28159 (N_28159,N_27195,N_26350);
xnor U28160 (N_28160,N_26608,N_26431);
nand U28161 (N_28161,N_27599,N_26735);
nor U28162 (N_28162,N_26029,N_26135);
and U28163 (N_28163,N_26820,N_27344);
nand U28164 (N_28164,N_27567,N_27976);
or U28165 (N_28165,N_26183,N_27205);
xnor U28166 (N_28166,N_27595,N_27225);
xor U28167 (N_28167,N_27230,N_27992);
nand U28168 (N_28168,N_26141,N_26245);
nor U28169 (N_28169,N_27394,N_27924);
and U28170 (N_28170,N_26097,N_26812);
nand U28171 (N_28171,N_26323,N_26188);
or U28172 (N_28172,N_27629,N_26377);
and U28173 (N_28173,N_27353,N_27973);
and U28174 (N_28174,N_27749,N_27288);
and U28175 (N_28175,N_27982,N_26228);
and U28176 (N_28176,N_27770,N_26150);
or U28177 (N_28177,N_27224,N_26341);
or U28178 (N_28178,N_26175,N_26213);
nor U28179 (N_28179,N_26575,N_27578);
or U28180 (N_28180,N_26545,N_27832);
xnor U28181 (N_28181,N_27707,N_27304);
or U28182 (N_28182,N_27912,N_27803);
and U28183 (N_28183,N_26171,N_27613);
or U28184 (N_28184,N_27447,N_27614);
or U28185 (N_28185,N_26065,N_27229);
and U28186 (N_28186,N_26246,N_26165);
and U28187 (N_28187,N_27326,N_26003);
nand U28188 (N_28188,N_26853,N_27634);
nor U28189 (N_28189,N_26664,N_26294);
xor U28190 (N_28190,N_27369,N_27935);
and U28191 (N_28191,N_26430,N_26225);
and U28192 (N_28192,N_26785,N_26444);
xnor U28193 (N_28193,N_26508,N_26174);
and U28194 (N_28194,N_26044,N_26869);
xor U28195 (N_28195,N_27028,N_27566);
or U28196 (N_28196,N_26258,N_27154);
or U28197 (N_28197,N_26384,N_26948);
xor U28198 (N_28198,N_26969,N_26717);
or U28199 (N_28199,N_26559,N_26085);
xor U28200 (N_28200,N_26218,N_27064);
or U28201 (N_28201,N_26958,N_26311);
or U28202 (N_28202,N_27921,N_26319);
nor U28203 (N_28203,N_26795,N_27503);
nor U28204 (N_28204,N_26060,N_27814);
and U28205 (N_28205,N_26154,N_27845);
nand U28206 (N_28206,N_27037,N_26550);
or U28207 (N_28207,N_26013,N_27048);
nand U28208 (N_28208,N_27745,N_27200);
and U28209 (N_28209,N_26705,N_26697);
xnor U28210 (N_28210,N_26799,N_26249);
nand U28211 (N_28211,N_26120,N_26994);
nand U28212 (N_28212,N_26951,N_26699);
xnor U28213 (N_28213,N_26027,N_27053);
and U28214 (N_28214,N_27627,N_27931);
or U28215 (N_28215,N_26130,N_26307);
nand U28216 (N_28216,N_27170,N_26616);
and U28217 (N_28217,N_26418,N_26216);
nor U28218 (N_28218,N_26922,N_27920);
nand U28219 (N_28219,N_27817,N_27004);
nor U28220 (N_28220,N_26504,N_26942);
xnor U28221 (N_28221,N_27475,N_27741);
nand U28222 (N_28222,N_26093,N_26205);
or U28223 (N_28223,N_27619,N_26965);
or U28224 (N_28224,N_26159,N_26787);
xor U28225 (N_28225,N_26767,N_27919);
nor U28226 (N_28226,N_26533,N_27440);
and U28227 (N_28227,N_27419,N_26153);
and U28228 (N_28228,N_27012,N_26986);
nor U28229 (N_28229,N_26008,N_26660);
nor U28230 (N_28230,N_26012,N_27754);
nor U28231 (N_28231,N_26827,N_26527);
nor U28232 (N_28232,N_26976,N_26845);
nor U28233 (N_28233,N_27909,N_26472);
xnor U28234 (N_28234,N_26987,N_26931);
or U28235 (N_28235,N_27457,N_26178);
xor U28236 (N_28236,N_27927,N_26464);
xnor U28237 (N_28237,N_27274,N_26941);
nand U28238 (N_28238,N_27385,N_27325);
or U28239 (N_28239,N_26256,N_27628);
nand U28240 (N_28240,N_26666,N_26414);
nand U28241 (N_28241,N_27270,N_26102);
nor U28242 (N_28242,N_26581,N_27232);
nor U28243 (N_28243,N_27724,N_27056);
nor U28244 (N_28244,N_26146,N_26731);
and U28245 (N_28245,N_26199,N_26945);
and U28246 (N_28246,N_26091,N_26597);
nand U28247 (N_28247,N_27652,N_26194);
nand U28248 (N_28248,N_27630,N_27291);
nand U28249 (N_28249,N_26566,N_26372);
or U28250 (N_28250,N_26162,N_27806);
nand U28251 (N_28251,N_26721,N_26623);
nand U28252 (N_28252,N_26318,N_26694);
nand U28253 (N_28253,N_26624,N_27180);
nand U28254 (N_28254,N_27415,N_27812);
or U28255 (N_28255,N_26465,N_27778);
and U28256 (N_28256,N_26950,N_26313);
and U28257 (N_28257,N_27177,N_27239);
nor U28258 (N_28258,N_26574,N_26383);
xnor U28259 (N_28259,N_27850,N_26919);
xnor U28260 (N_28260,N_26645,N_26074);
xnor U28261 (N_28261,N_27459,N_27418);
nor U28262 (N_28262,N_27437,N_26552);
or U28263 (N_28263,N_26387,N_26293);
nor U28264 (N_28264,N_27504,N_27398);
and U28265 (N_28265,N_26176,N_27968);
nand U28266 (N_28266,N_27474,N_27965);
and U28267 (N_28267,N_27174,N_27861);
nand U28268 (N_28268,N_27317,N_26089);
xor U28269 (N_28269,N_26144,N_26344);
and U28270 (N_28270,N_27213,N_26872);
nand U28271 (N_28271,N_26700,N_26557);
or U28272 (N_28272,N_27134,N_27097);
and U28273 (N_28273,N_27715,N_26026);
and U28274 (N_28274,N_27718,N_26327);
and U28275 (N_28275,N_26437,N_27403);
or U28276 (N_28276,N_27782,N_27899);
xor U28277 (N_28277,N_26620,N_26047);
or U28278 (N_28278,N_27050,N_27319);
nand U28279 (N_28279,N_27767,N_27423);
xor U28280 (N_28280,N_26277,N_27874);
nor U28281 (N_28281,N_26599,N_27928);
or U28282 (N_28282,N_27366,N_26458);
or U28283 (N_28283,N_27809,N_26718);
xor U28284 (N_28284,N_27489,N_27677);
xnor U28285 (N_28285,N_27826,N_27495);
and U28286 (N_28286,N_26158,N_27837);
or U28287 (N_28287,N_26775,N_27980);
nor U28288 (N_28288,N_27683,N_26558);
nor U28289 (N_28289,N_26916,N_27332);
and U28290 (N_28290,N_27866,N_26887);
nand U28291 (N_28291,N_26197,N_26977);
nand U28292 (N_28292,N_26177,N_27744);
or U28293 (N_28293,N_26975,N_26447);
nor U28294 (N_28294,N_26935,N_26331);
nand U28295 (N_28295,N_27278,N_26899);
xor U28296 (N_28296,N_27116,N_26446);
xor U28297 (N_28297,N_27545,N_26399);
or U28298 (N_28298,N_26688,N_27896);
xnor U28299 (N_28299,N_26936,N_26841);
xnor U28300 (N_28300,N_26896,N_27219);
nor U28301 (N_28301,N_26272,N_27303);
and U28302 (N_28302,N_27271,N_27994);
or U28303 (N_28303,N_26374,N_27103);
and U28304 (N_28304,N_27362,N_26962);
nand U28305 (N_28305,N_27507,N_27747);
xnor U28306 (N_28306,N_26343,N_27710);
nor U28307 (N_28307,N_26450,N_26315);
xor U28308 (N_28308,N_27482,N_27062);
nor U28309 (N_28309,N_26874,N_26349);
nor U28310 (N_28310,N_27142,N_27783);
nand U28311 (N_28311,N_26719,N_26443);
and U28312 (N_28312,N_26782,N_27716);
or U28313 (N_28313,N_27206,N_26901);
and U28314 (N_28314,N_27068,N_27355);
nand U28315 (N_28315,N_27906,N_27844);
and U28316 (N_28316,N_27790,N_27824);
or U28317 (N_28317,N_26804,N_27049);
nor U28318 (N_28318,N_27723,N_27802);
and U28319 (N_28319,N_27530,N_27590);
nand U28320 (N_28320,N_27589,N_27301);
xnor U28321 (N_28321,N_27351,N_27038);
nand U28322 (N_28322,N_27681,N_27150);
nand U28323 (N_28323,N_27880,N_26081);
xor U28324 (N_28324,N_27252,N_27798);
nor U28325 (N_28325,N_27643,N_26764);
nor U28326 (N_28326,N_27494,N_27720);
nand U28327 (N_28327,N_26676,N_26160);
nand U28328 (N_28328,N_27961,N_26715);
nor U28329 (N_28329,N_27588,N_27751);
or U28330 (N_28330,N_26672,N_27730);
nand U28331 (N_28331,N_26032,N_27162);
nor U28332 (N_28332,N_27808,N_26789);
nor U28333 (N_28333,N_27186,N_27289);
and U28334 (N_28334,N_27911,N_26388);
and U28335 (N_28335,N_27011,N_26203);
nand U28336 (N_28336,N_27354,N_26202);
or U28337 (N_28337,N_26006,N_27891);
xnor U28338 (N_28338,N_26190,N_26304);
xnor U28339 (N_28339,N_26912,N_26644);
or U28340 (N_28340,N_27686,N_26328);
nor U28341 (N_28341,N_27445,N_26662);
xor U28342 (N_28342,N_27938,N_27971);
xor U28343 (N_28343,N_26696,N_27498);
nor U28344 (N_28344,N_27295,N_26200);
nand U28345 (N_28345,N_27540,N_27221);
and U28346 (N_28346,N_26923,N_26234);
and U28347 (N_28347,N_27079,N_27795);
or U28348 (N_28348,N_26870,N_27580);
nand U28349 (N_28349,N_26244,N_26569);
xnor U28350 (N_28350,N_27405,N_26117);
xor U28351 (N_28351,N_27214,N_26217);
and U28352 (N_28352,N_27318,N_27022);
and U28353 (N_28353,N_27093,N_27902);
and U28354 (N_28354,N_26556,N_27496);
nand U28355 (N_28355,N_27510,N_27182);
or U28356 (N_28356,N_26992,N_27649);
or U28357 (N_28357,N_27799,N_27564);
and U28358 (N_28358,N_27661,N_27210);
and U28359 (N_28359,N_27622,N_26588);
and U28360 (N_28360,N_27438,N_26985);
xnor U28361 (N_28361,N_27001,N_26786);
nand U28362 (N_28362,N_27096,N_26166);
nand U28363 (N_28363,N_26438,N_27420);
or U28364 (N_28364,N_27313,N_26636);
or U28365 (N_28365,N_26041,N_26867);
or U28366 (N_28366,N_27835,N_27163);
nor U28367 (N_28367,N_26979,N_27433);
or U28368 (N_28368,N_26904,N_27253);
or U28369 (N_28369,N_27328,N_26926);
and U28370 (N_28370,N_26051,N_27106);
nand U28371 (N_28371,N_26289,N_26800);
nor U28372 (N_28372,N_27312,N_27490);
or U28373 (N_28373,N_27222,N_27243);
nor U28374 (N_28374,N_26686,N_27098);
or U28375 (N_28375,N_27436,N_27115);
or U28376 (N_28376,N_26055,N_27544);
and U28377 (N_28377,N_27800,N_26134);
and U28378 (N_28378,N_26455,N_27719);
or U28379 (N_28379,N_27947,N_26128);
nor U28380 (N_28380,N_27841,N_27542);
nor U28381 (N_28381,N_26955,N_26921);
or U28382 (N_28382,N_27998,N_27139);
nor U28383 (N_28383,N_27178,N_26591);
xor U28384 (N_28384,N_26340,N_27082);
nand U28385 (N_28385,N_27984,N_26858);
xor U28386 (N_28386,N_27669,N_26741);
or U28387 (N_28387,N_26539,N_27675);
xnor U28388 (N_28388,N_26161,N_26809);
nor U28389 (N_28389,N_27534,N_27734);
xor U28390 (N_28390,N_26382,N_27538);
xor U28391 (N_28391,N_26727,N_27063);
nand U28392 (N_28392,N_27603,N_27847);
and U28393 (N_28393,N_27135,N_27527);
or U28394 (N_28394,N_26357,N_26685);
nor U28395 (N_28395,N_26635,N_26279);
nor U28396 (N_28396,N_27290,N_27340);
nor U28397 (N_28397,N_27929,N_27945);
and U28398 (N_28398,N_27479,N_26860);
and U28399 (N_28399,N_26521,N_27102);
nand U28400 (N_28400,N_26674,N_27425);
or U28401 (N_28401,N_26436,N_27563);
nand U28402 (N_28402,N_27157,N_27907);
xnor U28403 (N_28403,N_26449,N_27088);
nor U28404 (N_28404,N_26960,N_27245);
and U28405 (N_28405,N_27349,N_26501);
or U28406 (N_28406,N_27551,N_27836);
or U28407 (N_28407,N_26826,N_27784);
xnor U28408 (N_28408,N_27548,N_27072);
nand U28409 (N_28409,N_27343,N_26254);
xnor U28410 (N_28410,N_27878,N_27999);
xnor U28411 (N_28411,N_26732,N_26325);
and U28412 (N_28412,N_26821,N_27104);
and U28413 (N_28413,N_26811,N_26584);
nand U28414 (N_28414,N_27073,N_27827);
and U28415 (N_28415,N_27129,N_26549);
or U28416 (N_28416,N_26522,N_27089);
nor U28417 (N_28417,N_26375,N_26291);
and U28418 (N_28418,N_27897,N_26034);
xor U28419 (N_28419,N_26949,N_27549);
nand U28420 (N_28420,N_26145,N_26754);
nand U28421 (N_28421,N_26888,N_26582);
and U28422 (N_28422,N_26292,N_27693);
and U28423 (N_28423,N_26126,N_27914);
nor U28424 (N_28424,N_26698,N_26288);
nand U28425 (N_28425,N_27020,N_27164);
and U28426 (N_28426,N_26229,N_27043);
and U28427 (N_28427,N_27172,N_26320);
xor U28428 (N_28428,N_27499,N_27854);
xor U28429 (N_28429,N_27374,N_27010);
and U28430 (N_28430,N_27360,N_27523);
or U28431 (N_28431,N_26471,N_26570);
or U28432 (N_28432,N_26658,N_27903);
nand U28433 (N_28433,N_27728,N_27008);
and U28434 (N_28434,N_26125,N_26413);
nand U28435 (N_28435,N_27378,N_26580);
or U28436 (N_28436,N_27368,N_27570);
and U28437 (N_28437,N_27633,N_26185);
or U28438 (N_28438,N_26100,N_26573);
nor U28439 (N_28439,N_27396,N_27478);
nand U28440 (N_28440,N_27508,N_26308);
nand U28441 (N_28441,N_27524,N_26365);
or U28442 (N_28442,N_27789,N_26376);
nor U28443 (N_28443,N_27857,N_26462);
xor U28444 (N_28444,N_27641,N_27740);
xnor U28445 (N_28445,N_26138,N_26961);
nand U28446 (N_28446,N_27158,N_26560);
nand U28447 (N_28447,N_26538,N_27462);
and U28448 (N_28448,N_27339,N_26540);
nor U28449 (N_28449,N_27721,N_27760);
xor U28450 (N_28450,N_26371,N_26187);
and U28451 (N_28451,N_26397,N_27124);
xnor U28452 (N_28452,N_27923,N_26825);
or U28453 (N_28453,N_26682,N_27021);
or U28454 (N_28454,N_27352,N_26009);
nor U28455 (N_28455,N_27637,N_26011);
or U28456 (N_28456,N_26062,N_26776);
nand U28457 (N_28457,N_27148,N_27293);
and U28458 (N_28458,N_27708,N_27582);
nor U28459 (N_28459,N_26136,N_27608);
xor U28460 (N_28460,N_27509,N_26829);
or U28461 (N_28461,N_26847,N_27991);
nor U28462 (N_28462,N_27898,N_27226);
nor U28463 (N_28463,N_27576,N_26354);
or U28464 (N_28464,N_26525,N_26156);
xor U28465 (N_28465,N_27660,N_27375);
and U28466 (N_28466,N_26937,N_26379);
xor U28467 (N_28467,N_26605,N_26983);
and U28468 (N_28468,N_26484,N_27281);
xnor U28469 (N_28469,N_27141,N_26408);
and U28470 (N_28470,N_27218,N_27562);
nor U28471 (N_28471,N_27401,N_26929);
or U28472 (N_28472,N_26010,N_27645);
or U28473 (N_28473,N_26607,N_26938);
nand U28474 (N_28474,N_27138,N_27771);
and U28475 (N_28475,N_26763,N_27922);
xnor U28476 (N_28476,N_27616,N_27035);
nand U28477 (N_28477,N_27663,N_27117);
xor U28478 (N_28478,N_27512,N_27264);
or U28479 (N_28479,N_27331,N_26595);
and U28480 (N_28480,N_27752,N_26053);
nor U28481 (N_28481,N_26750,N_27497);
or U28482 (N_28482,N_26708,N_27476);
nand U28483 (N_28483,N_26439,N_27381);
and U28484 (N_28484,N_27047,N_26259);
and U28485 (N_28485,N_27624,N_27765);
and U28486 (N_28486,N_27959,N_26692);
nand U28487 (N_28487,N_26637,N_27691);
and U28488 (N_28488,N_26630,N_27429);
and U28489 (N_28489,N_26959,N_26192);
or U28490 (N_28490,N_27166,N_27397);
nand U28491 (N_28491,N_27697,N_27391);
nand U28492 (N_28492,N_26779,N_26369);
nand U28493 (N_28493,N_27758,N_26726);
or U28494 (N_28494,N_26098,N_26833);
nand U28495 (N_28495,N_26316,N_26233);
xnor U28496 (N_28496,N_27940,N_26395);
or U28497 (N_28497,N_27522,N_27668);
xnor U28498 (N_28498,N_26486,N_26030);
and U28499 (N_28499,N_26193,N_27823);
nand U28500 (N_28500,N_26733,N_27240);
nand U28501 (N_28501,N_27671,N_27424);
or U28502 (N_28502,N_27521,N_26167);
or U28503 (N_28503,N_26615,N_26114);
nand U28504 (N_28504,N_27086,N_26168);
and U28505 (N_28505,N_27829,N_26070);
and U28506 (N_28506,N_26033,N_26433);
nor U28507 (N_28507,N_26593,N_26297);
xnor U28508 (N_28508,N_27236,N_26014);
nand U28509 (N_28509,N_26310,N_26480);
nor U28510 (N_28510,N_26788,N_27655);
nand U28511 (N_28511,N_27687,N_27621);
xnor U28512 (N_28512,N_26335,N_27254);
xor U28513 (N_28513,N_27943,N_26119);
nor U28514 (N_28514,N_27033,N_26184);
and U28515 (N_28515,N_26568,N_26654);
and U28516 (N_28516,N_27764,N_27617);
or U28517 (N_28517,N_26780,N_27776);
nor U28518 (N_28518,N_26578,N_27714);
nand U28519 (N_28519,N_27568,N_27345);
or U28520 (N_28520,N_26363,N_27644);
nand U28521 (N_28521,N_26037,N_27612);
xor U28522 (N_28522,N_27488,N_26769);
and U28523 (N_28523,N_26451,N_27910);
nor U28524 (N_28524,N_27598,N_26427);
and U28525 (N_28525,N_26531,N_27190);
or U28526 (N_28526,N_26876,N_26403);
and U28527 (N_28527,N_27664,N_27126);
nor U28528 (N_28528,N_27074,N_27505);
or U28529 (N_28529,N_26661,N_26163);
nor U28530 (N_28530,N_27819,N_26793);
nor U28531 (N_28531,N_26211,N_26339);
xor U28532 (N_28532,N_26248,N_26851);
or U28533 (N_28533,N_26857,N_27237);
nor U28534 (N_28534,N_27873,N_27777);
or U28535 (N_28535,N_27380,N_26634);
xor U28536 (N_28536,N_26652,N_27155);
nor U28537 (N_28537,N_27596,N_26481);
nand U28538 (N_28538,N_26269,N_27746);
nor U28539 (N_28539,N_26687,N_27387);
nand U28540 (N_28540,N_27535,N_27766);
nor U28541 (N_28541,N_26338,N_27893);
and U28542 (N_28542,N_27201,N_27554);
nand U28543 (N_28543,N_27217,N_26345);
nand U28544 (N_28544,N_27094,N_27587);
and U28545 (N_28545,N_27069,N_27967);
nand U28546 (N_28546,N_27114,N_27427);
xnor U28547 (N_28547,N_26442,N_26226);
nor U28548 (N_28548,N_27646,N_27044);
and U28549 (N_28549,N_26609,N_27762);
or U28550 (N_28550,N_26619,N_27543);
and U28551 (N_28551,N_27602,N_27638);
or U28552 (N_28552,N_27119,N_26633);
xor U28553 (N_28553,N_26406,N_27492);
nor U28554 (N_28554,N_26794,N_26651);
and U28555 (N_28555,N_26264,N_27149);
nand U28556 (N_28556,N_26749,N_26906);
xor U28557 (N_28557,N_27517,N_26878);
and U28558 (N_28558,N_27422,N_26621);
and U28559 (N_28559,N_26880,N_27635);
xor U28560 (N_28560,N_26084,N_27605);
and U28561 (N_28561,N_26330,N_27547);
xnor U28562 (N_28562,N_26428,N_27772);
nand U28563 (N_28563,N_27533,N_27305);
nand U28564 (N_28564,N_26548,N_26577);
nor U28565 (N_28565,N_26737,N_26096);
or U28566 (N_28566,N_27860,N_27388);
nor U28567 (N_28567,N_27818,N_26092);
xor U28568 (N_28568,N_26610,N_27722);
and U28569 (N_28569,N_27692,N_27092);
nor U28570 (N_28570,N_26810,N_26367);
nor U28571 (N_28571,N_27597,N_26348);
or U28572 (N_28572,N_26629,N_27025);
nor U28573 (N_28573,N_26614,N_26276);
or U28574 (N_28574,N_27585,N_26806);
nand U28575 (N_28575,N_26210,N_27297);
nor U28576 (N_28576,N_26587,N_26866);
xor U28577 (N_28577,N_27653,N_27610);
nor U28578 (N_28578,N_26518,N_27852);
nor U28579 (N_28579,N_26250,N_27081);
xor U28580 (N_28580,N_26562,N_26611);
or U28581 (N_28581,N_27341,N_26004);
or U28582 (N_28582,N_27066,N_26653);
nand U28583 (N_28583,N_27449,N_26947);
xor U28584 (N_28584,N_27470,N_27501);
xor U28585 (N_28585,N_26172,N_26989);
xor U28586 (N_28586,N_27625,N_27640);
nand U28587 (N_28587,N_27672,N_26755);
nand U28588 (N_28588,N_27263,N_26555);
and U28589 (N_28589,N_27889,N_26094);
nor U28590 (N_28590,N_26057,N_27699);
and U28591 (N_28591,N_26526,N_26831);
nor U28592 (N_28592,N_27729,N_26546);
or U28593 (N_28593,N_27560,N_27112);
nand U28594 (N_28594,N_26918,N_27932);
or U28595 (N_28595,N_26492,N_27531);
or U28596 (N_28596,N_27925,N_26148);
xnor U28597 (N_28597,N_27363,N_26612);
xor U28598 (N_28598,N_27867,N_27451);
and U28599 (N_28599,N_26019,N_26774);
or U28600 (N_28600,N_27667,N_27954);
xor U28601 (N_28601,N_26756,N_26036);
or U28602 (N_28602,N_27247,N_27833);
or U28603 (N_28603,N_27272,N_27133);
nand U28604 (N_28604,N_27486,N_27838);
xor U28605 (N_28605,N_26007,N_27532);
nand U28606 (N_28606,N_26592,N_27471);
or U28607 (N_28607,N_26334,N_26934);
nor U28608 (N_28608,N_26157,N_27487);
and U28609 (N_28609,N_27933,N_27900);
or U28610 (N_28610,N_26677,N_26579);
xnor U28611 (N_28611,N_26807,N_26843);
xor U28612 (N_28612,N_27400,N_26215);
nand U28613 (N_28613,N_26059,N_26736);
or U28614 (N_28614,N_26104,N_26116);
nand U28615 (N_28615,N_27361,N_27642);
nor U28616 (N_28616,N_26745,N_26402);
or U28617 (N_28617,N_27739,N_27231);
xor U28618 (N_28618,N_26285,N_26631);
or U28619 (N_28619,N_26078,N_27032);
nand U28620 (N_28620,N_27846,N_27042);
xnor U28621 (N_28621,N_27666,N_26129);
xnor U28622 (N_28622,N_27858,N_27859);
xor U28623 (N_28623,N_26112,N_27593);
and U28624 (N_28624,N_27472,N_26201);
or U28625 (N_28625,N_27518,N_27978);
or U28626 (N_28626,N_26031,N_27153);
or U28627 (N_28627,N_27448,N_27019);
nor U28628 (N_28628,N_26152,N_26473);
nor U28629 (N_28629,N_27125,N_27515);
nor U28630 (N_28630,N_27848,N_27379);
or U28631 (N_28631,N_26396,N_27283);
or U28632 (N_28632,N_27586,N_26742);
and U28633 (N_28633,N_26695,N_27338);
nor U28634 (N_28634,N_26835,N_27485);
nor U28635 (N_28635,N_26392,N_26142);
nor U28636 (N_28636,N_26268,N_26702);
nand U28637 (N_28637,N_27689,N_26298);
and U28638 (N_28638,N_26275,N_27974);
or U28639 (N_28639,N_26890,N_27843);
nor U28640 (N_28640,N_26884,N_26115);
nand U28641 (N_28641,N_26452,N_26703);
or U28642 (N_28642,N_26143,N_27078);
xnor U28643 (N_28643,N_26675,N_27111);
or U28644 (N_28644,N_27188,N_26850);
nand U28645 (N_28645,N_27639,N_27416);
xor U28646 (N_28646,N_27774,N_26266);
and U28647 (N_28647,N_26900,N_27026);
nor U28648 (N_28648,N_26231,N_27316);
and U28649 (N_28649,N_26684,N_27315);
and U28650 (N_28650,N_26284,N_26576);
xnor U28651 (N_28651,N_26204,N_27395);
or U28652 (N_28652,N_26113,N_27888);
nand U28653 (N_28653,N_26898,N_26710);
and U28654 (N_28654,N_26257,N_27009);
nand U28655 (N_28655,N_27132,N_26421);
or U28656 (N_28656,N_26048,N_27255);
or U28657 (N_28657,N_26127,N_27185);
nor U28658 (N_28658,N_26111,N_27000);
and U28659 (N_28659,N_27146,N_27559);
nand U28660 (N_28660,N_27256,N_26784);
and U28661 (N_28661,N_27886,N_27280);
and U28662 (N_28662,N_27051,N_27431);
or U28663 (N_28663,N_27516,N_27399);
nand U28664 (N_28664,N_27198,N_27690);
or U28665 (N_28665,N_27087,N_26892);
xnor U28666 (N_28666,N_27227,N_26714);
xor U28667 (N_28667,N_27091,N_26359);
and U28668 (N_28668,N_27052,N_26895);
nor U28669 (N_28669,N_26524,N_27709);
nor U28670 (N_28670,N_27528,N_27678);
and U28671 (N_28671,N_27071,N_27650);
or U28672 (N_28672,N_26882,N_27376);
or U28673 (N_28673,N_27005,N_27007);
xnor U28674 (N_28674,N_26220,N_27990);
nand U28675 (N_28675,N_26393,N_26381);
nor U28676 (N_28676,N_26389,N_26056);
and U28677 (N_28677,N_27737,N_26740);
and U28678 (N_28678,N_27386,N_27100);
nor U28679 (N_28679,N_26863,N_27840);
xor U28680 (N_28680,N_27763,N_27575);
xnor U28681 (N_28681,N_26572,N_27075);
nor U28682 (N_28682,N_27569,N_26542);
and U28683 (N_28683,N_27500,N_27023);
or U28684 (N_28684,N_27813,N_26132);
nand U28685 (N_28685,N_27735,N_26227);
and U28686 (N_28686,N_27165,N_26498);
and U28687 (N_28687,N_26151,N_26864);
xnor U28688 (N_28688,N_26667,N_26641);
xor U28689 (N_28689,N_26650,N_27953);
or U28690 (N_28690,N_27942,N_27552);
and U28691 (N_28691,N_26238,N_26622);
nand U28692 (N_28692,N_26299,N_26083);
xor U28693 (N_28693,N_26485,N_26543);
xnor U28694 (N_28694,N_26999,N_26657);
and U28695 (N_28695,N_27855,N_27029);
and U28696 (N_28696,N_26673,N_26426);
nand U28697 (N_28697,N_26739,N_26585);
or U28698 (N_28698,N_26196,N_27785);
xnor U28699 (N_28699,N_26988,N_27414);
nor U28700 (N_28700,N_26946,N_27805);
and U28701 (N_28701,N_26409,N_27659);
nand U28702 (N_28702,N_26106,N_27324);
xnor U28703 (N_28703,N_26747,N_26836);
xnor U28704 (N_28704,N_27466,N_26240);
nand U28705 (N_28705,N_26602,N_26862);
nor U28706 (N_28706,N_26720,N_27529);
xor U28707 (N_28707,N_26838,N_26905);
xor U28708 (N_28708,N_27147,N_27109);
or U28709 (N_28709,N_27483,N_27688);
or U28710 (N_28710,N_26554,N_27662);
or U28711 (N_28711,N_27342,N_26844);
nand U28712 (N_28712,N_27307,N_26468);
nor U28713 (N_28713,N_26260,N_26713);
nor U28714 (N_28714,N_27266,N_26064);
or U28715 (N_28715,N_26886,N_27571);
and U28716 (N_28716,N_26802,N_26968);
or U28717 (N_28717,N_27875,N_27249);
and U28718 (N_28718,N_27300,N_26072);
nor U28719 (N_28719,N_26483,N_27989);
nand U28720 (N_28720,N_27885,N_26459);
xnor U28721 (N_28721,N_27411,N_26295);
nor U28722 (N_28722,N_27145,N_26980);
xor U28723 (N_28723,N_26221,N_26963);
nand U28724 (N_28724,N_26716,N_26571);
xor U28725 (N_28725,N_27988,N_26822);
xor U28726 (N_28726,N_26038,N_26405);
and U28727 (N_28727,N_26908,N_26474);
and U28728 (N_28728,N_27831,N_26879);
nand U28729 (N_28729,N_27811,N_27202);
and U28730 (N_28730,N_26478,N_26537);
and U28731 (N_28731,N_27615,N_27383);
xor U28732 (N_28732,N_27792,N_26243);
and U28733 (N_28733,N_26212,N_27477);
or U28734 (N_28734,N_26865,N_26709);
and U28735 (N_28735,N_27674,N_26681);
or U28736 (N_28736,N_27402,N_27526);
or U28737 (N_28737,N_26005,N_26670);
nand U28738 (N_28738,N_27665,N_27941);
nor U28739 (N_28739,N_26173,N_26604);
xnor U28740 (N_28740,N_27323,N_27144);
or U28741 (N_28741,N_27275,N_26600);
xnor U28742 (N_28742,N_26470,N_27196);
and U28743 (N_28743,N_27143,N_26475);
nand U28744 (N_28744,N_26503,N_26973);
xor U28745 (N_28745,N_27851,N_26770);
and U28746 (N_28746,N_26131,N_27679);
xor U28747 (N_28747,N_27309,N_27958);
nor U28748 (N_28748,N_26410,N_27657);
nand U28749 (N_28749,N_26380,N_27862);
and U28750 (N_28750,N_27908,N_26925);
xor U28751 (N_28751,N_27828,N_27684);
or U28752 (N_28752,N_27373,N_26235);
or U28753 (N_28753,N_26467,N_27572);
xnor U28754 (N_28754,N_26765,N_27565);
nor U28755 (N_28755,N_27265,N_26598);
or U28756 (N_28756,N_26523,N_26109);
nor U28757 (N_28757,N_26347,N_26329);
xor U28758 (N_28758,N_27228,N_27197);
nand U28759 (N_28759,N_26978,N_26859);
or U28760 (N_28760,N_27979,N_27654);
nand U28761 (N_28761,N_27561,N_26954);
nor U28762 (N_28762,N_27757,N_26326);
or U28763 (N_28763,N_26691,N_26797);
nand U28764 (N_28764,N_26118,N_27658);
xor U28765 (N_28765,N_26169,N_27913);
nand U28766 (N_28766,N_26875,N_27611);
and U28767 (N_28767,N_27017,N_26404);
or U28768 (N_28768,N_26832,N_27045);
xnor U28769 (N_28769,N_27673,N_26390);
nor U28770 (N_28770,N_26039,N_27892);
nor U28771 (N_28771,N_26247,N_27884);
or U28772 (N_28772,N_26454,N_26751);
nand U28773 (N_28773,N_27456,N_26262);
nand U28774 (N_28774,N_27258,N_26182);
and U28775 (N_28775,N_26618,N_27748);
nand U28776 (N_28776,N_27918,N_26424);
xnor U28777 (N_28777,N_27333,N_26219);
nor U28778 (N_28778,N_27282,N_26366);
or U28779 (N_28779,N_26309,N_26846);
nand U28780 (N_28780,N_26282,N_27262);
nor U28781 (N_28781,N_26067,N_27871);
or U28782 (N_28782,N_27732,N_26885);
or U28783 (N_28783,N_27389,N_26488);
or U28784 (N_28784,N_27514,N_27726);
nor U28785 (N_28785,N_26626,N_26683);
or U28786 (N_28786,N_27685,N_26957);
and U28787 (N_28787,N_27525,N_27432);
and U28788 (N_28788,N_26312,N_26099);
nand U28789 (N_28789,N_26828,N_27127);
or U28790 (N_28790,N_26370,N_27090);
nor U28791 (N_28791,N_27372,N_26606);
and U28792 (N_28792,N_27251,N_26834);
and U28793 (N_28793,N_26290,N_27346);
nor U28794 (N_28794,N_27781,N_26512);
nand U28795 (N_28795,N_26314,N_27113);
nor U28796 (N_28796,N_27623,N_26586);
and U28797 (N_28797,N_26270,N_27294);
and U28798 (N_28798,N_26642,N_26701);
xnor U28799 (N_28799,N_27890,N_26280);
nand U28800 (N_28800,N_26553,N_27830);
or U28801 (N_28801,N_26515,N_27108);
xnor U28802 (N_28802,N_27215,N_27260);
xnor U28803 (N_28803,N_26940,N_26332);
and U28804 (N_28804,N_27706,N_26970);
and U28805 (N_28805,N_26930,N_26924);
xnor U28806 (N_28806,N_27916,N_27084);
nor U28807 (N_28807,N_27443,N_27299);
xnor U28808 (N_28808,N_26758,N_26974);
nor U28809 (N_28809,N_26017,N_27384);
or U28810 (N_28810,N_26840,N_27327);
nor U28811 (N_28811,N_26054,N_27464);
nor U28812 (N_28812,N_27736,N_26791);
nand U28813 (N_28813,N_27442,N_27713);
xnor U28814 (N_28814,N_26487,N_27995);
or U28815 (N_28815,N_26286,N_27905);
and U28816 (N_28816,N_26123,N_26241);
nor U28817 (N_28817,N_26302,N_26668);
nor U28818 (N_28818,N_26362,N_27952);
nand U28819 (N_28819,N_26956,N_27292);
or U28820 (N_28820,N_27557,N_26416);
and U28821 (N_28821,N_26209,N_27469);
nand U28822 (N_28822,N_26223,N_26551);
nor U28823 (N_28823,N_26944,N_27193);
nor U28824 (N_28824,N_27536,N_26358);
xor U28825 (N_28825,N_26049,N_27452);
nand U28826 (N_28826,N_26045,N_27390);
nor U28827 (N_28827,N_27711,N_26296);
xnor U28828 (N_28828,N_27577,N_27701);
and U28829 (N_28829,N_27058,N_26237);
xnor U28830 (N_28830,N_26730,N_26342);
or U28831 (N_28831,N_26928,N_27592);
xnor U28832 (N_28832,N_27337,N_27002);
xnor U28833 (N_28833,N_26261,N_26773);
or U28834 (N_28834,N_27320,N_27118);
nor U28835 (N_28835,N_26933,N_26640);
nand U28836 (N_28836,N_26781,N_26998);
xor U28837 (N_28837,N_26046,N_26669);
nand U28838 (N_28838,N_27584,N_27314);
nor U28839 (N_28839,N_27430,N_26783);
nand U28840 (N_28840,N_26649,N_26170);
or U28841 (N_28841,N_26236,N_27480);
nand U28842 (N_28842,N_26671,N_27788);
nand U28843 (N_28843,N_26743,N_27435);
and U28844 (N_28844,N_26147,N_26351);
nor U28845 (N_28845,N_27881,N_27676);
nand U28846 (N_28846,N_27883,N_26434);
xor U28847 (N_28847,N_26255,N_26792);
nor U28848 (N_28848,N_27975,N_26206);
nor U28849 (N_28849,N_26655,N_27960);
or U28850 (N_28850,N_27934,N_27944);
or U28851 (N_28851,N_26561,N_27926);
nand U28852 (N_28852,N_27250,N_26020);
and U28853 (N_28853,N_26516,N_26830);
xor U28854 (N_28854,N_26920,N_27018);
and U28855 (N_28855,N_26953,N_26757);
nand U28856 (N_28856,N_27027,N_26306);
or U28857 (N_28857,N_26964,N_27040);
nor U28858 (N_28858,N_27175,N_27842);
or U28859 (N_28859,N_26353,N_27868);
nand U28860 (N_28860,N_27233,N_26107);
nand U28861 (N_28861,N_27834,N_26423);
nand U28862 (N_28862,N_26180,N_26513);
nor U28863 (N_28863,N_26803,N_27964);
nand U28864 (N_28864,N_26647,N_26601);
and U28865 (N_28865,N_27876,N_27981);
or U28866 (N_28866,N_27370,N_27248);
nand U28867 (N_28867,N_27864,N_27804);
or U28868 (N_28868,N_26122,N_26704);
and U28869 (N_28869,N_26466,N_26411);
xor U28870 (N_28870,N_27455,N_26181);
and U28871 (N_28871,N_27986,N_27463);
nor U28872 (N_28872,N_26952,N_26482);
nand U28873 (N_28873,N_26394,N_27321);
nor U28874 (N_28874,N_26453,N_27887);
and U28875 (N_28875,N_27412,N_27347);
or U28876 (N_28876,N_26448,N_26305);
and U28877 (N_28877,N_27894,N_26848);
xor U28878 (N_28878,N_27061,N_26509);
or U28879 (N_28879,N_27753,N_27951);
nand U28880 (N_28880,N_26638,N_26707);
or U28881 (N_28881,N_26738,N_27511);
nand U28882 (N_28882,N_26643,N_27787);
nor U28883 (N_28883,N_27107,N_27626);
nor U28884 (N_28884,N_26519,N_27356);
nor U28885 (N_28885,N_26752,N_27296);
or U28886 (N_28886,N_27453,N_26469);
nand U28887 (N_28887,N_27807,N_26253);
or U28888 (N_28888,N_27972,N_26042);
and U28889 (N_28889,N_27413,N_26040);
nor U28890 (N_28890,N_27006,N_26932);
and U28891 (N_28891,N_27110,N_26386);
xor U28892 (N_28892,N_27120,N_27171);
and U28893 (N_28893,N_27286,N_26839);
xnor U28894 (N_28894,N_26425,N_27013);
or U28895 (N_28895,N_26728,N_26068);
nand U28896 (N_28896,N_27181,N_26398);
nand U28897 (N_28897,N_26915,N_27816);
nand U28898 (N_28898,N_27558,N_27284);
or U28899 (N_28899,N_26364,N_27189);
or U28900 (N_28900,N_27244,N_27267);
or U28901 (N_28901,N_26273,N_26506);
xor U28902 (N_28902,N_27601,N_26082);
nor U28903 (N_28903,N_27950,N_26361);
or U28904 (N_28904,N_26534,N_27651);
nor U28905 (N_28905,N_26164,N_27484);
or U28906 (N_28906,N_26678,N_27212);
nor U28907 (N_28907,N_27199,N_26854);
or U28908 (N_28908,N_27620,N_27136);
nand U28909 (N_28909,N_27095,N_26066);
and U28910 (N_28910,N_26910,N_27377);
and U28911 (N_28911,N_26303,N_26493);
and U28912 (N_28912,N_26967,N_27695);
or U28913 (N_28913,N_27322,N_26417);
xor U28914 (N_28914,N_26613,N_26317);
nand U28915 (N_28915,N_27502,N_26544);
xnor U28916 (N_28916,N_27204,N_27137);
or U28917 (N_28917,N_26768,N_27223);
nand U28918 (N_28918,N_26195,N_27696);
nor U28919 (N_28919,N_26088,N_26494);
and U28920 (N_28920,N_27298,N_26909);
or U28921 (N_28921,N_27167,N_26617);
nor U28922 (N_28922,N_27041,N_27895);
or U28923 (N_28923,N_27030,N_27183);
nand U28924 (N_28924,N_27365,N_26035);
nor U28925 (N_28925,N_26095,N_27773);
xnor U28926 (N_28926,N_27070,N_26108);
nor U28927 (N_28927,N_26179,N_27242);
or U28928 (N_28928,N_27216,N_27609);
nor U28929 (N_28929,N_27359,N_27302);
xor U28930 (N_28930,N_27393,N_27985);
nand U28931 (N_28931,N_26894,N_26412);
xor U28932 (N_28932,N_26762,N_27434);
or U28933 (N_28933,N_27970,N_27334);
xor U28934 (N_28934,N_26603,N_27879);
xnor U28935 (N_28935,N_26208,N_26063);
nor U28936 (N_28936,N_26407,N_26071);
nor U28937 (N_28937,N_26693,N_26401);
nor U28938 (N_28938,N_26913,N_27937);
nand U28939 (N_28939,N_26356,N_26242);
and U28940 (N_28940,N_27308,N_26023);
nor U28941 (N_28941,N_27553,N_26966);
nor U28942 (N_28942,N_27441,N_26287);
nand U28943 (N_28943,N_26191,N_27768);
nor U28944 (N_28944,N_26028,N_26984);
nor U28945 (N_28945,N_27698,N_26734);
nor U28946 (N_28946,N_26400,N_26018);
xnor U28947 (N_28947,N_27335,N_27796);
nor U28948 (N_28948,N_26744,N_26429);
xor U28949 (N_28949,N_27059,N_26819);
nand U28950 (N_28950,N_27410,N_27791);
or U28951 (N_28951,N_26917,N_26656);
and U28952 (N_28952,N_27080,N_27648);
nor U28953 (N_28953,N_26547,N_26189);
nor U28954 (N_28954,N_27473,N_26463);
or U28955 (N_28955,N_27016,N_26690);
or U28956 (N_28956,N_27101,N_27865);
and U28957 (N_28957,N_26771,N_26564);
nor U28958 (N_28958,N_27786,N_26583);
or U28959 (N_28959,N_26911,N_26360);
and U28960 (N_28960,N_27591,N_26352);
or U28961 (N_28961,N_26103,N_26816);
nor U28962 (N_28962,N_27151,N_27268);
nand U28963 (N_28963,N_27822,N_26263);
nor U28964 (N_28964,N_26322,N_26489);
xnor U28965 (N_28965,N_26746,N_26355);
nor U28966 (N_28966,N_27409,N_26278);
and U28967 (N_28967,N_26457,N_26479);
nor U28968 (N_28968,N_27034,N_26724);
xnor U28969 (N_28969,N_26101,N_26058);
nand U28970 (N_28970,N_27983,N_26015);
or U28971 (N_28971,N_27234,N_27060);
and U28972 (N_28972,N_26712,N_27357);
xor U28973 (N_28973,N_26420,N_27863);
xnor U28974 (N_28974,N_27191,N_27915);
xor U28975 (N_28975,N_27417,N_26024);
nor U28976 (N_28976,N_27161,N_27076);
xor U28977 (N_28977,N_26798,N_26856);
and U28978 (N_28978,N_27203,N_26301);
or U28979 (N_28979,N_27276,N_26378);
nand U28980 (N_28980,N_27966,N_26532);
nor U28981 (N_28981,N_26761,N_27725);
nor U28982 (N_28982,N_26445,N_26563);
nand U28983 (N_28983,N_26903,N_26321);
and U28984 (N_28984,N_26981,N_26198);
nor U28985 (N_28985,N_27439,N_27987);
xnor U28986 (N_28986,N_26507,N_27140);
nand U28987 (N_28987,N_26589,N_27194);
xnor U28988 (N_28988,N_27731,N_27694);
and U28989 (N_28989,N_27520,N_26711);
nor U28990 (N_28990,N_26230,N_26337);
or U28991 (N_28991,N_26267,N_26016);
nand U28992 (N_28992,N_27168,N_26596);
and U28993 (N_28993,N_27815,N_26883);
nand U28994 (N_28994,N_26823,N_26140);
xnor U28995 (N_28995,N_27184,N_27936);
and U28996 (N_28996,N_26861,N_26777);
and U28997 (N_28997,N_26990,N_27382);
nor U28998 (N_28998,N_27277,N_27364);
or U28999 (N_28999,N_27285,N_26528);
and U29000 (N_29000,N_27737,N_26718);
nand U29001 (N_29001,N_26605,N_26195);
xor U29002 (N_29002,N_27196,N_27501);
nand U29003 (N_29003,N_26850,N_26135);
nor U29004 (N_29004,N_26242,N_26373);
and U29005 (N_29005,N_26204,N_26918);
and U29006 (N_29006,N_26977,N_27953);
xor U29007 (N_29007,N_27629,N_26481);
xor U29008 (N_29008,N_26621,N_27794);
or U29009 (N_29009,N_27556,N_27618);
xnor U29010 (N_29010,N_27959,N_27727);
and U29011 (N_29011,N_26936,N_27365);
nor U29012 (N_29012,N_27933,N_26032);
nor U29013 (N_29013,N_27743,N_27409);
nor U29014 (N_29014,N_27444,N_26255);
and U29015 (N_29015,N_27933,N_27882);
or U29016 (N_29016,N_27739,N_27296);
or U29017 (N_29017,N_26671,N_26364);
nor U29018 (N_29018,N_26415,N_26454);
xnor U29019 (N_29019,N_27483,N_27116);
nor U29020 (N_29020,N_27425,N_27125);
or U29021 (N_29021,N_26676,N_26554);
or U29022 (N_29022,N_27915,N_27274);
nor U29023 (N_29023,N_27069,N_27860);
xor U29024 (N_29024,N_27400,N_26020);
nand U29025 (N_29025,N_26790,N_26774);
or U29026 (N_29026,N_27155,N_27701);
and U29027 (N_29027,N_27441,N_27478);
and U29028 (N_29028,N_26931,N_26368);
nor U29029 (N_29029,N_27797,N_26140);
or U29030 (N_29030,N_26167,N_27620);
or U29031 (N_29031,N_27910,N_27331);
and U29032 (N_29032,N_26671,N_27033);
nand U29033 (N_29033,N_27412,N_26340);
and U29034 (N_29034,N_26254,N_27425);
nand U29035 (N_29035,N_26490,N_26119);
nor U29036 (N_29036,N_26786,N_27103);
xnor U29037 (N_29037,N_27646,N_27544);
xor U29038 (N_29038,N_26368,N_27838);
nand U29039 (N_29039,N_27575,N_27181);
nand U29040 (N_29040,N_26975,N_27292);
xor U29041 (N_29041,N_26348,N_26248);
nand U29042 (N_29042,N_27340,N_26463);
xnor U29043 (N_29043,N_26290,N_26117);
nand U29044 (N_29044,N_26392,N_26186);
xor U29045 (N_29045,N_26506,N_27446);
nor U29046 (N_29046,N_26939,N_26271);
or U29047 (N_29047,N_26306,N_26676);
and U29048 (N_29048,N_26688,N_27954);
and U29049 (N_29049,N_27758,N_26578);
or U29050 (N_29050,N_26627,N_26777);
and U29051 (N_29051,N_26437,N_26122);
and U29052 (N_29052,N_27035,N_27447);
or U29053 (N_29053,N_26828,N_27335);
xor U29054 (N_29054,N_26826,N_26549);
and U29055 (N_29055,N_26040,N_27553);
nand U29056 (N_29056,N_26823,N_27144);
nor U29057 (N_29057,N_26872,N_27592);
or U29058 (N_29058,N_26668,N_26510);
nor U29059 (N_29059,N_26585,N_27337);
or U29060 (N_29060,N_27507,N_27191);
nand U29061 (N_29061,N_27329,N_26619);
and U29062 (N_29062,N_27387,N_27356);
and U29063 (N_29063,N_26102,N_27947);
or U29064 (N_29064,N_26712,N_27474);
nor U29065 (N_29065,N_26327,N_26044);
nand U29066 (N_29066,N_26520,N_27466);
xnor U29067 (N_29067,N_27281,N_26571);
nor U29068 (N_29068,N_26964,N_27323);
nand U29069 (N_29069,N_27098,N_27985);
nand U29070 (N_29070,N_26301,N_27880);
nor U29071 (N_29071,N_27687,N_27854);
and U29072 (N_29072,N_27925,N_26966);
xor U29073 (N_29073,N_26116,N_27522);
nand U29074 (N_29074,N_26241,N_27087);
xnor U29075 (N_29075,N_26438,N_26384);
nor U29076 (N_29076,N_27788,N_27476);
and U29077 (N_29077,N_26361,N_27588);
nand U29078 (N_29078,N_26499,N_27655);
or U29079 (N_29079,N_27596,N_27227);
or U29080 (N_29080,N_27524,N_26796);
nor U29081 (N_29081,N_26343,N_26276);
xor U29082 (N_29082,N_27724,N_27767);
or U29083 (N_29083,N_26804,N_26018);
and U29084 (N_29084,N_26934,N_27024);
xnor U29085 (N_29085,N_26947,N_27276);
nor U29086 (N_29086,N_26590,N_26933);
nor U29087 (N_29087,N_26577,N_26463);
or U29088 (N_29088,N_27100,N_27782);
nand U29089 (N_29089,N_27058,N_27916);
nor U29090 (N_29090,N_26446,N_26431);
and U29091 (N_29091,N_27195,N_27019);
and U29092 (N_29092,N_26061,N_27851);
xor U29093 (N_29093,N_27362,N_26147);
xor U29094 (N_29094,N_27229,N_26731);
nor U29095 (N_29095,N_26780,N_26716);
nor U29096 (N_29096,N_26136,N_26000);
xor U29097 (N_29097,N_26480,N_27110);
and U29098 (N_29098,N_26270,N_26955);
nand U29099 (N_29099,N_26290,N_27877);
nand U29100 (N_29100,N_27112,N_26190);
nand U29101 (N_29101,N_27190,N_26316);
nor U29102 (N_29102,N_27988,N_26966);
nor U29103 (N_29103,N_26402,N_26666);
xnor U29104 (N_29104,N_26496,N_27076);
or U29105 (N_29105,N_26560,N_27671);
nand U29106 (N_29106,N_27236,N_27709);
or U29107 (N_29107,N_27780,N_26623);
and U29108 (N_29108,N_27063,N_27183);
nand U29109 (N_29109,N_27514,N_26242);
or U29110 (N_29110,N_27140,N_27977);
xor U29111 (N_29111,N_26106,N_27304);
nor U29112 (N_29112,N_27299,N_26248);
xor U29113 (N_29113,N_27163,N_26268);
or U29114 (N_29114,N_26629,N_27234);
or U29115 (N_29115,N_27949,N_26852);
and U29116 (N_29116,N_27481,N_26168);
and U29117 (N_29117,N_27865,N_27934);
nor U29118 (N_29118,N_26005,N_27388);
nor U29119 (N_29119,N_26310,N_26641);
nor U29120 (N_29120,N_27943,N_26475);
nor U29121 (N_29121,N_27952,N_27351);
nand U29122 (N_29122,N_27457,N_26164);
and U29123 (N_29123,N_27381,N_27535);
nand U29124 (N_29124,N_26176,N_27327);
nand U29125 (N_29125,N_26666,N_27680);
or U29126 (N_29126,N_26498,N_26831);
or U29127 (N_29127,N_26920,N_27177);
xor U29128 (N_29128,N_26510,N_27042);
or U29129 (N_29129,N_27432,N_26012);
nand U29130 (N_29130,N_27400,N_26459);
xor U29131 (N_29131,N_27956,N_26060);
nor U29132 (N_29132,N_26277,N_26381);
or U29133 (N_29133,N_27846,N_27124);
or U29134 (N_29134,N_27472,N_27418);
xnor U29135 (N_29135,N_27793,N_26810);
xnor U29136 (N_29136,N_26316,N_27758);
nor U29137 (N_29137,N_26495,N_27746);
nand U29138 (N_29138,N_26108,N_27699);
nor U29139 (N_29139,N_26670,N_27262);
or U29140 (N_29140,N_27978,N_27155);
nand U29141 (N_29141,N_27505,N_27216);
or U29142 (N_29142,N_26031,N_27424);
nand U29143 (N_29143,N_26684,N_26365);
nand U29144 (N_29144,N_27582,N_26539);
nor U29145 (N_29145,N_26137,N_27573);
xor U29146 (N_29146,N_26364,N_27294);
or U29147 (N_29147,N_26550,N_26184);
and U29148 (N_29148,N_26908,N_26301);
and U29149 (N_29149,N_27660,N_26543);
and U29150 (N_29150,N_27538,N_26421);
xnor U29151 (N_29151,N_26876,N_26772);
and U29152 (N_29152,N_26617,N_27597);
xor U29153 (N_29153,N_26154,N_26804);
nor U29154 (N_29154,N_27648,N_27811);
nand U29155 (N_29155,N_27273,N_26676);
or U29156 (N_29156,N_26864,N_26108);
nand U29157 (N_29157,N_26126,N_26246);
nand U29158 (N_29158,N_26793,N_26541);
and U29159 (N_29159,N_26539,N_27167);
and U29160 (N_29160,N_26745,N_26676);
xnor U29161 (N_29161,N_26602,N_26556);
or U29162 (N_29162,N_27395,N_27018);
and U29163 (N_29163,N_26619,N_27305);
nand U29164 (N_29164,N_27700,N_26107);
nand U29165 (N_29165,N_26211,N_27658);
or U29166 (N_29166,N_26868,N_26014);
and U29167 (N_29167,N_26388,N_26208);
nand U29168 (N_29168,N_27553,N_26551);
or U29169 (N_29169,N_26495,N_26850);
nor U29170 (N_29170,N_26403,N_27851);
nand U29171 (N_29171,N_26972,N_26952);
or U29172 (N_29172,N_27164,N_26930);
nand U29173 (N_29173,N_26270,N_26016);
xnor U29174 (N_29174,N_26199,N_27292);
and U29175 (N_29175,N_27658,N_26733);
and U29176 (N_29176,N_26207,N_26859);
nor U29177 (N_29177,N_26423,N_27605);
or U29178 (N_29178,N_27508,N_26805);
nand U29179 (N_29179,N_26599,N_26475);
and U29180 (N_29180,N_27964,N_27223);
or U29181 (N_29181,N_26116,N_27841);
xnor U29182 (N_29182,N_27043,N_27900);
and U29183 (N_29183,N_26034,N_27048);
xor U29184 (N_29184,N_26840,N_27014);
and U29185 (N_29185,N_27484,N_26752);
and U29186 (N_29186,N_26577,N_27022);
nor U29187 (N_29187,N_27923,N_26592);
nor U29188 (N_29188,N_27696,N_26443);
nand U29189 (N_29189,N_26509,N_26609);
nand U29190 (N_29190,N_26362,N_27650);
and U29191 (N_29191,N_26972,N_27246);
nand U29192 (N_29192,N_26305,N_26580);
or U29193 (N_29193,N_26664,N_26480);
nand U29194 (N_29194,N_26428,N_26544);
and U29195 (N_29195,N_27658,N_26361);
nand U29196 (N_29196,N_27517,N_27743);
or U29197 (N_29197,N_26367,N_27103);
or U29198 (N_29198,N_26922,N_27165);
nor U29199 (N_29199,N_27015,N_27819);
nor U29200 (N_29200,N_27793,N_26105);
nand U29201 (N_29201,N_27855,N_27368);
or U29202 (N_29202,N_26860,N_27718);
and U29203 (N_29203,N_27003,N_27996);
nand U29204 (N_29204,N_26766,N_26650);
xor U29205 (N_29205,N_27537,N_26551);
xor U29206 (N_29206,N_27753,N_26685);
and U29207 (N_29207,N_26049,N_26178);
xor U29208 (N_29208,N_26765,N_26894);
xnor U29209 (N_29209,N_27208,N_27729);
and U29210 (N_29210,N_27874,N_27999);
xor U29211 (N_29211,N_26499,N_26046);
xnor U29212 (N_29212,N_26558,N_27096);
nand U29213 (N_29213,N_26547,N_26265);
or U29214 (N_29214,N_27150,N_27992);
nor U29215 (N_29215,N_27473,N_27661);
and U29216 (N_29216,N_26959,N_27822);
and U29217 (N_29217,N_27371,N_26947);
xnor U29218 (N_29218,N_27026,N_27741);
nand U29219 (N_29219,N_27197,N_26837);
nor U29220 (N_29220,N_26140,N_26064);
nor U29221 (N_29221,N_26459,N_26254);
and U29222 (N_29222,N_27601,N_27952);
and U29223 (N_29223,N_26550,N_26079);
nand U29224 (N_29224,N_27908,N_26897);
nor U29225 (N_29225,N_27415,N_26134);
nand U29226 (N_29226,N_27613,N_27363);
nand U29227 (N_29227,N_26581,N_27571);
nand U29228 (N_29228,N_27718,N_27628);
or U29229 (N_29229,N_27115,N_26519);
xor U29230 (N_29230,N_27677,N_26886);
nand U29231 (N_29231,N_27634,N_27731);
nor U29232 (N_29232,N_27740,N_26789);
and U29233 (N_29233,N_26158,N_27715);
and U29234 (N_29234,N_26041,N_27007);
xnor U29235 (N_29235,N_26464,N_27515);
nor U29236 (N_29236,N_27592,N_27091);
or U29237 (N_29237,N_27687,N_26713);
nand U29238 (N_29238,N_26750,N_27944);
and U29239 (N_29239,N_26609,N_26916);
and U29240 (N_29240,N_26578,N_26191);
and U29241 (N_29241,N_26406,N_27657);
nand U29242 (N_29242,N_27915,N_27825);
nor U29243 (N_29243,N_27843,N_27494);
and U29244 (N_29244,N_27565,N_27801);
xnor U29245 (N_29245,N_27662,N_27908);
or U29246 (N_29246,N_27351,N_27208);
xor U29247 (N_29247,N_27079,N_27062);
xor U29248 (N_29248,N_27681,N_26354);
xor U29249 (N_29249,N_26268,N_26495);
nor U29250 (N_29250,N_27580,N_27085);
nor U29251 (N_29251,N_26296,N_26701);
and U29252 (N_29252,N_26444,N_26032);
xor U29253 (N_29253,N_27037,N_26944);
and U29254 (N_29254,N_27052,N_26988);
xnor U29255 (N_29255,N_26473,N_26404);
nor U29256 (N_29256,N_26017,N_26106);
nor U29257 (N_29257,N_26626,N_27479);
or U29258 (N_29258,N_26968,N_27630);
and U29259 (N_29259,N_27409,N_26922);
or U29260 (N_29260,N_26455,N_26351);
nor U29261 (N_29261,N_26762,N_27435);
xnor U29262 (N_29262,N_26620,N_27531);
xnor U29263 (N_29263,N_27902,N_26359);
xor U29264 (N_29264,N_27733,N_27728);
xnor U29265 (N_29265,N_27923,N_27908);
or U29266 (N_29266,N_26572,N_27996);
or U29267 (N_29267,N_26990,N_26392);
or U29268 (N_29268,N_27000,N_27345);
xor U29269 (N_29269,N_26451,N_27396);
or U29270 (N_29270,N_27961,N_26830);
or U29271 (N_29271,N_26489,N_27037);
or U29272 (N_29272,N_26842,N_26800);
or U29273 (N_29273,N_27341,N_26795);
xor U29274 (N_29274,N_27760,N_26262);
nand U29275 (N_29275,N_26582,N_26227);
and U29276 (N_29276,N_26191,N_27110);
or U29277 (N_29277,N_26483,N_26219);
and U29278 (N_29278,N_27249,N_26570);
and U29279 (N_29279,N_27515,N_27565);
nor U29280 (N_29280,N_26291,N_26677);
nor U29281 (N_29281,N_27888,N_26456);
or U29282 (N_29282,N_26087,N_27348);
and U29283 (N_29283,N_26268,N_27151);
xnor U29284 (N_29284,N_26113,N_27515);
and U29285 (N_29285,N_26037,N_26483);
nor U29286 (N_29286,N_27093,N_26807);
and U29287 (N_29287,N_27443,N_26120);
or U29288 (N_29288,N_26627,N_27352);
xnor U29289 (N_29289,N_27285,N_26791);
nand U29290 (N_29290,N_26902,N_27283);
nand U29291 (N_29291,N_27557,N_27722);
nand U29292 (N_29292,N_27382,N_26696);
nand U29293 (N_29293,N_26631,N_26215);
nor U29294 (N_29294,N_26125,N_27425);
or U29295 (N_29295,N_26213,N_26439);
nand U29296 (N_29296,N_26447,N_27112);
or U29297 (N_29297,N_27907,N_27931);
nor U29298 (N_29298,N_27423,N_27150);
nand U29299 (N_29299,N_26422,N_26601);
xnor U29300 (N_29300,N_27558,N_26307);
or U29301 (N_29301,N_26989,N_27085);
nor U29302 (N_29302,N_27222,N_27671);
nand U29303 (N_29303,N_27248,N_27597);
or U29304 (N_29304,N_26074,N_27861);
and U29305 (N_29305,N_27346,N_27762);
or U29306 (N_29306,N_26707,N_26739);
nor U29307 (N_29307,N_26370,N_26252);
nand U29308 (N_29308,N_27800,N_26800);
nor U29309 (N_29309,N_26836,N_27265);
xor U29310 (N_29310,N_26768,N_27619);
nand U29311 (N_29311,N_27555,N_26508);
or U29312 (N_29312,N_26341,N_27201);
nand U29313 (N_29313,N_27089,N_26029);
or U29314 (N_29314,N_27418,N_27849);
nor U29315 (N_29315,N_27651,N_27983);
xnor U29316 (N_29316,N_26897,N_26348);
xor U29317 (N_29317,N_27616,N_26167);
or U29318 (N_29318,N_27712,N_26726);
or U29319 (N_29319,N_27927,N_26347);
nand U29320 (N_29320,N_26815,N_26733);
nor U29321 (N_29321,N_26294,N_26891);
nand U29322 (N_29322,N_27580,N_27924);
xnor U29323 (N_29323,N_26961,N_27944);
and U29324 (N_29324,N_26215,N_27404);
xnor U29325 (N_29325,N_26875,N_26059);
nand U29326 (N_29326,N_26589,N_26482);
or U29327 (N_29327,N_27696,N_26521);
nor U29328 (N_29328,N_26377,N_26618);
nor U29329 (N_29329,N_27592,N_26290);
nand U29330 (N_29330,N_26239,N_26079);
or U29331 (N_29331,N_27481,N_26942);
nand U29332 (N_29332,N_26834,N_27808);
and U29333 (N_29333,N_27021,N_27139);
nand U29334 (N_29334,N_26265,N_27709);
nor U29335 (N_29335,N_26756,N_26076);
nand U29336 (N_29336,N_27191,N_27403);
xnor U29337 (N_29337,N_27637,N_26143);
xnor U29338 (N_29338,N_26040,N_27772);
nand U29339 (N_29339,N_26592,N_26226);
nor U29340 (N_29340,N_26220,N_27864);
and U29341 (N_29341,N_27894,N_27582);
and U29342 (N_29342,N_26152,N_26973);
and U29343 (N_29343,N_26047,N_26150);
nor U29344 (N_29344,N_27419,N_26230);
nor U29345 (N_29345,N_27990,N_26885);
or U29346 (N_29346,N_27899,N_26013);
nand U29347 (N_29347,N_27729,N_26366);
nor U29348 (N_29348,N_26226,N_27177);
nor U29349 (N_29349,N_26240,N_26770);
nand U29350 (N_29350,N_27049,N_27830);
and U29351 (N_29351,N_26943,N_27695);
nor U29352 (N_29352,N_26895,N_26268);
nand U29353 (N_29353,N_26689,N_26196);
or U29354 (N_29354,N_26693,N_26363);
or U29355 (N_29355,N_26293,N_27416);
nand U29356 (N_29356,N_26636,N_27940);
xnor U29357 (N_29357,N_26155,N_27886);
nand U29358 (N_29358,N_26491,N_27120);
nand U29359 (N_29359,N_27253,N_27665);
or U29360 (N_29360,N_26333,N_27626);
or U29361 (N_29361,N_27635,N_27985);
and U29362 (N_29362,N_27578,N_27033);
nand U29363 (N_29363,N_26549,N_26710);
xnor U29364 (N_29364,N_26639,N_26966);
or U29365 (N_29365,N_27041,N_26085);
nor U29366 (N_29366,N_27519,N_27013);
or U29367 (N_29367,N_26491,N_26157);
xnor U29368 (N_29368,N_27552,N_27269);
xor U29369 (N_29369,N_27632,N_27763);
nand U29370 (N_29370,N_26008,N_27714);
or U29371 (N_29371,N_27545,N_27952);
xnor U29372 (N_29372,N_27503,N_27751);
and U29373 (N_29373,N_26126,N_27551);
and U29374 (N_29374,N_27189,N_27836);
nand U29375 (N_29375,N_26425,N_27411);
and U29376 (N_29376,N_26012,N_27933);
nor U29377 (N_29377,N_26201,N_27753);
and U29378 (N_29378,N_27621,N_26807);
and U29379 (N_29379,N_26857,N_27348);
nor U29380 (N_29380,N_27255,N_26269);
xor U29381 (N_29381,N_26157,N_26915);
or U29382 (N_29382,N_26168,N_27258);
xnor U29383 (N_29383,N_27533,N_26689);
xnor U29384 (N_29384,N_26963,N_26519);
and U29385 (N_29385,N_27048,N_27415);
and U29386 (N_29386,N_26642,N_26634);
nor U29387 (N_29387,N_27803,N_26884);
or U29388 (N_29388,N_26362,N_27874);
or U29389 (N_29389,N_26773,N_27448);
nor U29390 (N_29390,N_27280,N_26474);
xor U29391 (N_29391,N_27795,N_27354);
nor U29392 (N_29392,N_26893,N_26029);
nand U29393 (N_29393,N_26641,N_26655);
and U29394 (N_29394,N_26949,N_26647);
and U29395 (N_29395,N_26681,N_26689);
and U29396 (N_29396,N_26297,N_27745);
nor U29397 (N_29397,N_27597,N_26093);
xor U29398 (N_29398,N_26480,N_27837);
xor U29399 (N_29399,N_27567,N_26755);
nand U29400 (N_29400,N_26112,N_26921);
and U29401 (N_29401,N_27286,N_26221);
or U29402 (N_29402,N_26855,N_26152);
nor U29403 (N_29403,N_27429,N_26631);
xor U29404 (N_29404,N_26166,N_27642);
xnor U29405 (N_29405,N_27598,N_26252);
or U29406 (N_29406,N_27800,N_26011);
xnor U29407 (N_29407,N_26563,N_26680);
xor U29408 (N_29408,N_27733,N_26882);
nand U29409 (N_29409,N_27308,N_27440);
or U29410 (N_29410,N_27008,N_27582);
and U29411 (N_29411,N_26828,N_27450);
nand U29412 (N_29412,N_27963,N_27739);
or U29413 (N_29413,N_26860,N_27729);
and U29414 (N_29414,N_27254,N_26635);
nand U29415 (N_29415,N_26649,N_27018);
nor U29416 (N_29416,N_26148,N_26585);
nor U29417 (N_29417,N_26766,N_27962);
and U29418 (N_29418,N_27492,N_27480);
or U29419 (N_29419,N_26394,N_26083);
or U29420 (N_29420,N_26285,N_26062);
nand U29421 (N_29421,N_27405,N_27986);
and U29422 (N_29422,N_26578,N_26388);
xor U29423 (N_29423,N_26063,N_27139);
xor U29424 (N_29424,N_27267,N_26545);
xor U29425 (N_29425,N_27270,N_26948);
or U29426 (N_29426,N_26216,N_27700);
nand U29427 (N_29427,N_27977,N_26312);
nor U29428 (N_29428,N_27023,N_27241);
and U29429 (N_29429,N_27079,N_27810);
and U29430 (N_29430,N_27871,N_26631);
xnor U29431 (N_29431,N_27618,N_26445);
and U29432 (N_29432,N_27387,N_27507);
nand U29433 (N_29433,N_27905,N_27083);
and U29434 (N_29434,N_26105,N_26920);
xnor U29435 (N_29435,N_27267,N_27833);
nand U29436 (N_29436,N_27368,N_27329);
and U29437 (N_29437,N_27122,N_27649);
xor U29438 (N_29438,N_27546,N_26009);
and U29439 (N_29439,N_27581,N_27050);
and U29440 (N_29440,N_27613,N_27620);
or U29441 (N_29441,N_26783,N_26135);
and U29442 (N_29442,N_27787,N_26922);
nand U29443 (N_29443,N_27916,N_26640);
nand U29444 (N_29444,N_26321,N_27754);
xor U29445 (N_29445,N_27384,N_26724);
nand U29446 (N_29446,N_27124,N_26348);
xor U29447 (N_29447,N_26269,N_26007);
xnor U29448 (N_29448,N_26467,N_26925);
nor U29449 (N_29449,N_26538,N_27651);
nand U29450 (N_29450,N_26914,N_27434);
xor U29451 (N_29451,N_27830,N_26092);
xnor U29452 (N_29452,N_26278,N_27807);
xor U29453 (N_29453,N_26221,N_26597);
or U29454 (N_29454,N_26990,N_27367);
xor U29455 (N_29455,N_26530,N_26073);
or U29456 (N_29456,N_26888,N_27010);
nand U29457 (N_29457,N_26027,N_26348);
nor U29458 (N_29458,N_26879,N_27771);
xnor U29459 (N_29459,N_26383,N_27320);
xor U29460 (N_29460,N_27916,N_26754);
xor U29461 (N_29461,N_27811,N_27262);
and U29462 (N_29462,N_26991,N_27486);
nor U29463 (N_29463,N_26450,N_26474);
nand U29464 (N_29464,N_26465,N_27650);
nand U29465 (N_29465,N_27198,N_26998);
nand U29466 (N_29466,N_27796,N_26831);
and U29467 (N_29467,N_27202,N_27580);
or U29468 (N_29468,N_26876,N_26373);
or U29469 (N_29469,N_26051,N_26624);
nand U29470 (N_29470,N_26990,N_27038);
and U29471 (N_29471,N_27622,N_26290);
nor U29472 (N_29472,N_26409,N_27648);
and U29473 (N_29473,N_26929,N_27614);
xnor U29474 (N_29474,N_27852,N_27786);
xnor U29475 (N_29475,N_27673,N_27415);
xor U29476 (N_29476,N_27391,N_26635);
and U29477 (N_29477,N_27209,N_26203);
or U29478 (N_29478,N_26067,N_26466);
or U29479 (N_29479,N_27344,N_27115);
nor U29480 (N_29480,N_26117,N_27816);
nor U29481 (N_29481,N_27845,N_27877);
xnor U29482 (N_29482,N_27225,N_26724);
or U29483 (N_29483,N_27268,N_27228);
xor U29484 (N_29484,N_27880,N_27733);
and U29485 (N_29485,N_26517,N_27499);
nand U29486 (N_29486,N_26391,N_27301);
or U29487 (N_29487,N_27466,N_27535);
xor U29488 (N_29488,N_26002,N_26630);
xnor U29489 (N_29489,N_27977,N_26706);
nor U29490 (N_29490,N_27318,N_26641);
and U29491 (N_29491,N_27609,N_27282);
and U29492 (N_29492,N_27908,N_26805);
or U29493 (N_29493,N_27556,N_26467);
nor U29494 (N_29494,N_27243,N_26100);
or U29495 (N_29495,N_27005,N_27551);
nand U29496 (N_29496,N_26323,N_27569);
and U29497 (N_29497,N_26214,N_26226);
and U29498 (N_29498,N_27518,N_27527);
nand U29499 (N_29499,N_27826,N_26958);
xor U29500 (N_29500,N_27451,N_27754);
xnor U29501 (N_29501,N_26895,N_26142);
and U29502 (N_29502,N_26459,N_27523);
or U29503 (N_29503,N_26263,N_27219);
or U29504 (N_29504,N_26715,N_27474);
and U29505 (N_29505,N_27622,N_26709);
xnor U29506 (N_29506,N_27598,N_26126);
nor U29507 (N_29507,N_27688,N_26946);
nand U29508 (N_29508,N_27506,N_26904);
nand U29509 (N_29509,N_26169,N_27206);
and U29510 (N_29510,N_27751,N_27031);
nor U29511 (N_29511,N_26966,N_27354);
nand U29512 (N_29512,N_27151,N_27285);
xor U29513 (N_29513,N_26112,N_26931);
nor U29514 (N_29514,N_27742,N_27807);
xnor U29515 (N_29515,N_26780,N_26371);
nand U29516 (N_29516,N_26860,N_26319);
and U29517 (N_29517,N_27407,N_27435);
and U29518 (N_29518,N_27664,N_27271);
nand U29519 (N_29519,N_27829,N_26032);
xnor U29520 (N_29520,N_26111,N_26651);
or U29521 (N_29521,N_27263,N_26684);
nor U29522 (N_29522,N_27023,N_27037);
nand U29523 (N_29523,N_27595,N_26772);
xnor U29524 (N_29524,N_26328,N_26905);
nand U29525 (N_29525,N_27080,N_27294);
nand U29526 (N_29526,N_27350,N_26339);
xnor U29527 (N_29527,N_27319,N_27700);
or U29528 (N_29528,N_27380,N_27532);
and U29529 (N_29529,N_27009,N_27433);
and U29530 (N_29530,N_27256,N_27219);
or U29531 (N_29531,N_27544,N_27286);
xnor U29532 (N_29532,N_27843,N_27059);
or U29533 (N_29533,N_26754,N_27545);
xnor U29534 (N_29534,N_27609,N_27553);
xnor U29535 (N_29535,N_26494,N_26814);
or U29536 (N_29536,N_27275,N_27159);
nand U29537 (N_29537,N_27017,N_26751);
or U29538 (N_29538,N_26396,N_26064);
or U29539 (N_29539,N_26197,N_26014);
nor U29540 (N_29540,N_27705,N_26797);
or U29541 (N_29541,N_26270,N_26594);
nor U29542 (N_29542,N_26944,N_27756);
nor U29543 (N_29543,N_26825,N_27444);
or U29544 (N_29544,N_26824,N_27672);
xnor U29545 (N_29545,N_26751,N_27444);
xnor U29546 (N_29546,N_27297,N_26803);
xor U29547 (N_29547,N_26463,N_27557);
nor U29548 (N_29548,N_26931,N_27471);
nand U29549 (N_29549,N_26355,N_26729);
xnor U29550 (N_29550,N_26381,N_26787);
nor U29551 (N_29551,N_27576,N_26403);
nor U29552 (N_29552,N_26042,N_26249);
xnor U29553 (N_29553,N_26776,N_27035);
and U29554 (N_29554,N_27923,N_27538);
or U29555 (N_29555,N_26149,N_26727);
xor U29556 (N_29556,N_26455,N_26438);
nand U29557 (N_29557,N_26388,N_27927);
xor U29558 (N_29558,N_27325,N_27311);
or U29559 (N_29559,N_26071,N_26112);
xnor U29560 (N_29560,N_27923,N_27963);
nor U29561 (N_29561,N_26818,N_26721);
and U29562 (N_29562,N_27631,N_27029);
nand U29563 (N_29563,N_27769,N_26403);
nand U29564 (N_29564,N_27439,N_26583);
xnor U29565 (N_29565,N_27848,N_27473);
xnor U29566 (N_29566,N_26583,N_26863);
xor U29567 (N_29567,N_26342,N_27922);
and U29568 (N_29568,N_27696,N_26940);
xor U29569 (N_29569,N_27392,N_26115);
or U29570 (N_29570,N_26744,N_26097);
xor U29571 (N_29571,N_26493,N_26242);
and U29572 (N_29572,N_26643,N_27756);
and U29573 (N_29573,N_26348,N_26145);
nor U29574 (N_29574,N_27708,N_27454);
nor U29575 (N_29575,N_27171,N_26837);
nor U29576 (N_29576,N_26931,N_27882);
or U29577 (N_29577,N_27112,N_26774);
xnor U29578 (N_29578,N_26560,N_26191);
nand U29579 (N_29579,N_26237,N_27627);
nor U29580 (N_29580,N_27344,N_26176);
nand U29581 (N_29581,N_27079,N_26825);
or U29582 (N_29582,N_27114,N_27095);
nor U29583 (N_29583,N_27949,N_27234);
xor U29584 (N_29584,N_26366,N_26595);
or U29585 (N_29585,N_26278,N_27236);
nand U29586 (N_29586,N_26652,N_27194);
or U29587 (N_29587,N_26254,N_27791);
and U29588 (N_29588,N_27095,N_26403);
xnor U29589 (N_29589,N_27051,N_27167);
xnor U29590 (N_29590,N_26265,N_26324);
or U29591 (N_29591,N_27294,N_27726);
and U29592 (N_29592,N_27226,N_26715);
xor U29593 (N_29593,N_26845,N_27515);
xor U29594 (N_29594,N_26142,N_26909);
nand U29595 (N_29595,N_26222,N_27557);
and U29596 (N_29596,N_26543,N_27569);
nor U29597 (N_29597,N_27314,N_26241);
xor U29598 (N_29598,N_26122,N_27109);
xnor U29599 (N_29599,N_26375,N_26718);
and U29600 (N_29600,N_27287,N_27514);
or U29601 (N_29601,N_27055,N_27921);
and U29602 (N_29602,N_26619,N_27334);
or U29603 (N_29603,N_27499,N_26936);
xnor U29604 (N_29604,N_27588,N_26392);
nor U29605 (N_29605,N_27665,N_26598);
nor U29606 (N_29606,N_26932,N_27803);
or U29607 (N_29607,N_27896,N_26960);
xor U29608 (N_29608,N_26365,N_26722);
xor U29609 (N_29609,N_27994,N_27926);
nand U29610 (N_29610,N_27272,N_27759);
nand U29611 (N_29611,N_27629,N_26147);
xor U29612 (N_29612,N_26539,N_27216);
or U29613 (N_29613,N_26295,N_27541);
xor U29614 (N_29614,N_27968,N_27159);
or U29615 (N_29615,N_26987,N_27859);
nor U29616 (N_29616,N_26476,N_26182);
nor U29617 (N_29617,N_26267,N_27173);
nor U29618 (N_29618,N_26814,N_27589);
and U29619 (N_29619,N_26552,N_26494);
nor U29620 (N_29620,N_26891,N_27573);
and U29621 (N_29621,N_26745,N_27127);
nor U29622 (N_29622,N_27756,N_27798);
nor U29623 (N_29623,N_27824,N_26737);
or U29624 (N_29624,N_27243,N_26258);
xnor U29625 (N_29625,N_27070,N_27286);
and U29626 (N_29626,N_26072,N_27451);
xor U29627 (N_29627,N_27217,N_27016);
nand U29628 (N_29628,N_27871,N_26660);
or U29629 (N_29629,N_27775,N_27602);
and U29630 (N_29630,N_26540,N_26707);
nand U29631 (N_29631,N_26909,N_27801);
and U29632 (N_29632,N_26552,N_26302);
xnor U29633 (N_29633,N_26197,N_26532);
xnor U29634 (N_29634,N_27716,N_27684);
nand U29635 (N_29635,N_26182,N_26169);
and U29636 (N_29636,N_27852,N_26747);
nand U29637 (N_29637,N_26153,N_26053);
nor U29638 (N_29638,N_26422,N_26879);
nand U29639 (N_29639,N_26156,N_27460);
xor U29640 (N_29640,N_26564,N_27357);
and U29641 (N_29641,N_27697,N_26123);
xor U29642 (N_29642,N_27238,N_26577);
or U29643 (N_29643,N_26278,N_27797);
nand U29644 (N_29644,N_26759,N_27251);
nand U29645 (N_29645,N_27855,N_27726);
nor U29646 (N_29646,N_27395,N_26882);
nand U29647 (N_29647,N_26627,N_27443);
nand U29648 (N_29648,N_27222,N_26875);
and U29649 (N_29649,N_27950,N_27848);
nor U29650 (N_29650,N_26252,N_26217);
and U29651 (N_29651,N_26200,N_26943);
xor U29652 (N_29652,N_27101,N_27982);
and U29653 (N_29653,N_27158,N_27000);
xor U29654 (N_29654,N_27770,N_27800);
and U29655 (N_29655,N_27684,N_26610);
and U29656 (N_29656,N_26215,N_27163);
and U29657 (N_29657,N_27192,N_27591);
nor U29658 (N_29658,N_27484,N_26742);
xor U29659 (N_29659,N_27211,N_27301);
nor U29660 (N_29660,N_27626,N_26419);
nand U29661 (N_29661,N_26556,N_26653);
nor U29662 (N_29662,N_27657,N_27439);
and U29663 (N_29663,N_26751,N_26709);
or U29664 (N_29664,N_27368,N_26918);
nor U29665 (N_29665,N_26271,N_26529);
nand U29666 (N_29666,N_27008,N_27714);
and U29667 (N_29667,N_27915,N_26396);
xnor U29668 (N_29668,N_27707,N_27458);
nor U29669 (N_29669,N_27524,N_26756);
xor U29670 (N_29670,N_26272,N_27996);
xnor U29671 (N_29671,N_26304,N_27212);
or U29672 (N_29672,N_26821,N_27250);
nand U29673 (N_29673,N_26583,N_27317);
nor U29674 (N_29674,N_27967,N_27065);
nor U29675 (N_29675,N_27639,N_27484);
or U29676 (N_29676,N_26770,N_26687);
nand U29677 (N_29677,N_26799,N_26232);
or U29678 (N_29678,N_26045,N_27668);
or U29679 (N_29679,N_27727,N_27422);
and U29680 (N_29680,N_26685,N_27141);
or U29681 (N_29681,N_27766,N_27589);
xnor U29682 (N_29682,N_27168,N_27690);
and U29683 (N_29683,N_27279,N_26011);
or U29684 (N_29684,N_27497,N_27215);
nor U29685 (N_29685,N_26773,N_26584);
nor U29686 (N_29686,N_27139,N_27381);
or U29687 (N_29687,N_26780,N_26553);
and U29688 (N_29688,N_26720,N_27068);
or U29689 (N_29689,N_27489,N_27696);
nor U29690 (N_29690,N_26382,N_27386);
or U29691 (N_29691,N_27707,N_26948);
nor U29692 (N_29692,N_27841,N_26198);
nor U29693 (N_29693,N_27242,N_26926);
nor U29694 (N_29694,N_26539,N_27476);
nand U29695 (N_29695,N_27072,N_26251);
xnor U29696 (N_29696,N_26947,N_26037);
nor U29697 (N_29697,N_26727,N_27534);
nor U29698 (N_29698,N_27562,N_26967);
xor U29699 (N_29699,N_27615,N_26110);
nor U29700 (N_29700,N_26569,N_26461);
or U29701 (N_29701,N_26283,N_26874);
nor U29702 (N_29702,N_26456,N_27546);
or U29703 (N_29703,N_26223,N_26096);
xnor U29704 (N_29704,N_26403,N_27843);
nand U29705 (N_29705,N_26314,N_27868);
and U29706 (N_29706,N_27422,N_27243);
nor U29707 (N_29707,N_27978,N_27320);
or U29708 (N_29708,N_26210,N_26823);
and U29709 (N_29709,N_26003,N_26198);
nor U29710 (N_29710,N_27175,N_27007);
nand U29711 (N_29711,N_27801,N_26309);
or U29712 (N_29712,N_26276,N_26359);
and U29713 (N_29713,N_26386,N_26621);
nor U29714 (N_29714,N_26711,N_26249);
nand U29715 (N_29715,N_26083,N_26747);
or U29716 (N_29716,N_27948,N_26436);
nor U29717 (N_29717,N_26210,N_26775);
xor U29718 (N_29718,N_26827,N_26814);
or U29719 (N_29719,N_26554,N_27079);
or U29720 (N_29720,N_26292,N_27959);
and U29721 (N_29721,N_27508,N_27130);
nor U29722 (N_29722,N_27637,N_27549);
and U29723 (N_29723,N_27535,N_27732);
and U29724 (N_29724,N_27502,N_26006);
xnor U29725 (N_29725,N_27278,N_27788);
nand U29726 (N_29726,N_27246,N_26914);
or U29727 (N_29727,N_26907,N_26100);
nor U29728 (N_29728,N_27354,N_26330);
xor U29729 (N_29729,N_26603,N_26365);
or U29730 (N_29730,N_27436,N_27959);
nor U29731 (N_29731,N_26443,N_26508);
nor U29732 (N_29732,N_27906,N_27661);
nor U29733 (N_29733,N_26784,N_27851);
nand U29734 (N_29734,N_27288,N_27032);
or U29735 (N_29735,N_27857,N_26428);
nand U29736 (N_29736,N_26506,N_26459);
xnor U29737 (N_29737,N_26756,N_26681);
nor U29738 (N_29738,N_27631,N_26927);
and U29739 (N_29739,N_26466,N_27223);
and U29740 (N_29740,N_26226,N_27135);
xnor U29741 (N_29741,N_27781,N_26684);
nand U29742 (N_29742,N_26038,N_27550);
xor U29743 (N_29743,N_26664,N_26287);
and U29744 (N_29744,N_27541,N_27824);
and U29745 (N_29745,N_27410,N_26019);
and U29746 (N_29746,N_27873,N_26097);
nand U29747 (N_29747,N_26496,N_27134);
or U29748 (N_29748,N_26441,N_27741);
nand U29749 (N_29749,N_26549,N_26187);
nand U29750 (N_29750,N_27003,N_26015);
xnor U29751 (N_29751,N_27101,N_27688);
nor U29752 (N_29752,N_27564,N_26362);
and U29753 (N_29753,N_27074,N_27124);
nor U29754 (N_29754,N_26777,N_27193);
nand U29755 (N_29755,N_27362,N_27326);
nand U29756 (N_29756,N_27043,N_26504);
nand U29757 (N_29757,N_26042,N_26476);
or U29758 (N_29758,N_27035,N_26664);
and U29759 (N_29759,N_26677,N_26005);
or U29760 (N_29760,N_26604,N_27915);
nor U29761 (N_29761,N_26047,N_27282);
nor U29762 (N_29762,N_26299,N_27480);
and U29763 (N_29763,N_27456,N_27948);
nor U29764 (N_29764,N_27737,N_26340);
or U29765 (N_29765,N_26190,N_27816);
nor U29766 (N_29766,N_26304,N_26807);
xor U29767 (N_29767,N_26005,N_26887);
nand U29768 (N_29768,N_27286,N_26309);
or U29769 (N_29769,N_26776,N_26861);
nor U29770 (N_29770,N_26764,N_26857);
and U29771 (N_29771,N_27055,N_26260);
nand U29772 (N_29772,N_27960,N_27629);
or U29773 (N_29773,N_27825,N_26016);
xnor U29774 (N_29774,N_26812,N_27398);
nor U29775 (N_29775,N_27474,N_26717);
xnor U29776 (N_29776,N_26501,N_26313);
xnor U29777 (N_29777,N_26468,N_27314);
xor U29778 (N_29778,N_26978,N_27699);
nand U29779 (N_29779,N_27312,N_27062);
nand U29780 (N_29780,N_27618,N_27389);
nand U29781 (N_29781,N_26106,N_26079);
xor U29782 (N_29782,N_27269,N_26449);
nand U29783 (N_29783,N_26428,N_27023);
and U29784 (N_29784,N_26863,N_26232);
nor U29785 (N_29785,N_27495,N_26969);
and U29786 (N_29786,N_26901,N_27558);
or U29787 (N_29787,N_27589,N_26899);
xor U29788 (N_29788,N_26524,N_27380);
nor U29789 (N_29789,N_27877,N_26408);
or U29790 (N_29790,N_27550,N_27606);
and U29791 (N_29791,N_26614,N_26295);
or U29792 (N_29792,N_26316,N_27490);
xnor U29793 (N_29793,N_27113,N_26414);
or U29794 (N_29794,N_26009,N_26180);
or U29795 (N_29795,N_26278,N_26328);
and U29796 (N_29796,N_27093,N_27301);
xnor U29797 (N_29797,N_27231,N_27608);
xor U29798 (N_29798,N_27689,N_27114);
nand U29799 (N_29799,N_27663,N_26923);
nor U29800 (N_29800,N_26451,N_27522);
nor U29801 (N_29801,N_26831,N_26910);
and U29802 (N_29802,N_26424,N_26128);
nand U29803 (N_29803,N_27318,N_26636);
nor U29804 (N_29804,N_26273,N_26622);
xnor U29805 (N_29805,N_27060,N_26796);
xnor U29806 (N_29806,N_27417,N_27985);
nand U29807 (N_29807,N_27852,N_26880);
or U29808 (N_29808,N_27937,N_26288);
and U29809 (N_29809,N_27517,N_26192);
nor U29810 (N_29810,N_26733,N_27132);
and U29811 (N_29811,N_26165,N_26427);
nand U29812 (N_29812,N_26184,N_27286);
and U29813 (N_29813,N_26481,N_27611);
nor U29814 (N_29814,N_26521,N_26143);
and U29815 (N_29815,N_26980,N_26626);
and U29816 (N_29816,N_26173,N_26347);
xnor U29817 (N_29817,N_27522,N_27925);
and U29818 (N_29818,N_27514,N_27061);
and U29819 (N_29819,N_27921,N_27544);
or U29820 (N_29820,N_27748,N_26011);
xor U29821 (N_29821,N_27819,N_26070);
and U29822 (N_29822,N_26639,N_27012);
nor U29823 (N_29823,N_26036,N_26909);
and U29824 (N_29824,N_26600,N_26924);
or U29825 (N_29825,N_27477,N_26596);
xnor U29826 (N_29826,N_27015,N_26140);
or U29827 (N_29827,N_27823,N_26211);
nor U29828 (N_29828,N_27896,N_27167);
nand U29829 (N_29829,N_26542,N_26074);
nor U29830 (N_29830,N_26693,N_26883);
and U29831 (N_29831,N_26197,N_26705);
or U29832 (N_29832,N_27715,N_27521);
or U29833 (N_29833,N_26231,N_27679);
nor U29834 (N_29834,N_27370,N_27930);
nand U29835 (N_29835,N_27223,N_26590);
or U29836 (N_29836,N_26610,N_27372);
nor U29837 (N_29837,N_27781,N_27365);
and U29838 (N_29838,N_27623,N_26986);
xnor U29839 (N_29839,N_26613,N_27886);
and U29840 (N_29840,N_27559,N_27808);
and U29841 (N_29841,N_27562,N_26393);
xnor U29842 (N_29842,N_26329,N_27288);
and U29843 (N_29843,N_26447,N_26523);
or U29844 (N_29844,N_26117,N_26827);
nand U29845 (N_29845,N_26528,N_27848);
xor U29846 (N_29846,N_26507,N_27956);
nor U29847 (N_29847,N_26207,N_26722);
nand U29848 (N_29848,N_26831,N_27676);
or U29849 (N_29849,N_26175,N_26911);
nor U29850 (N_29850,N_27463,N_27968);
xnor U29851 (N_29851,N_27787,N_26869);
or U29852 (N_29852,N_27139,N_27667);
nand U29853 (N_29853,N_27827,N_26056);
nand U29854 (N_29854,N_27577,N_26035);
xor U29855 (N_29855,N_26279,N_27046);
nand U29856 (N_29856,N_26361,N_27024);
xor U29857 (N_29857,N_27271,N_26546);
or U29858 (N_29858,N_26787,N_27624);
nor U29859 (N_29859,N_26207,N_26339);
and U29860 (N_29860,N_26937,N_27611);
xnor U29861 (N_29861,N_26153,N_26224);
xor U29862 (N_29862,N_26702,N_26026);
xnor U29863 (N_29863,N_27225,N_27052);
nand U29864 (N_29864,N_26054,N_27725);
nand U29865 (N_29865,N_26019,N_26354);
xor U29866 (N_29866,N_26117,N_27092);
xnor U29867 (N_29867,N_26274,N_27662);
xnor U29868 (N_29868,N_27784,N_27199);
xnor U29869 (N_29869,N_26785,N_26831);
xor U29870 (N_29870,N_27733,N_26478);
or U29871 (N_29871,N_26473,N_27640);
or U29872 (N_29872,N_27268,N_27366);
or U29873 (N_29873,N_27897,N_26508);
or U29874 (N_29874,N_26647,N_26091);
nand U29875 (N_29875,N_26179,N_26214);
xor U29876 (N_29876,N_26411,N_26422);
or U29877 (N_29877,N_26460,N_27343);
or U29878 (N_29878,N_26026,N_26990);
nand U29879 (N_29879,N_27807,N_26851);
and U29880 (N_29880,N_27445,N_26760);
and U29881 (N_29881,N_26560,N_27936);
xor U29882 (N_29882,N_26840,N_27911);
nand U29883 (N_29883,N_26731,N_26684);
nand U29884 (N_29884,N_27712,N_27008);
or U29885 (N_29885,N_27682,N_26157);
or U29886 (N_29886,N_27107,N_27714);
nand U29887 (N_29887,N_27553,N_26641);
and U29888 (N_29888,N_27037,N_27008);
and U29889 (N_29889,N_27432,N_26403);
nor U29890 (N_29890,N_27087,N_26530);
xnor U29891 (N_29891,N_27549,N_26617);
xnor U29892 (N_29892,N_27695,N_26745);
xnor U29893 (N_29893,N_27933,N_26176);
xnor U29894 (N_29894,N_26306,N_26428);
xor U29895 (N_29895,N_26525,N_26708);
xnor U29896 (N_29896,N_27516,N_26594);
or U29897 (N_29897,N_27567,N_26314);
and U29898 (N_29898,N_27642,N_26856);
xor U29899 (N_29899,N_26483,N_27427);
xor U29900 (N_29900,N_26418,N_27097);
and U29901 (N_29901,N_26243,N_26520);
nand U29902 (N_29902,N_27622,N_27454);
nor U29903 (N_29903,N_27327,N_26219);
and U29904 (N_29904,N_27763,N_27404);
nor U29905 (N_29905,N_26369,N_26190);
nor U29906 (N_29906,N_27679,N_27474);
xor U29907 (N_29907,N_26800,N_27084);
or U29908 (N_29908,N_26221,N_27647);
nand U29909 (N_29909,N_26297,N_26825);
nand U29910 (N_29910,N_27991,N_27681);
nor U29911 (N_29911,N_27521,N_27999);
and U29912 (N_29912,N_26580,N_26791);
and U29913 (N_29913,N_26205,N_26542);
and U29914 (N_29914,N_26761,N_27763);
xnor U29915 (N_29915,N_26450,N_27055);
nor U29916 (N_29916,N_26032,N_26518);
nand U29917 (N_29917,N_26636,N_27547);
and U29918 (N_29918,N_26778,N_26372);
nand U29919 (N_29919,N_27196,N_26159);
nand U29920 (N_29920,N_27831,N_26693);
or U29921 (N_29921,N_27275,N_27057);
nand U29922 (N_29922,N_27760,N_26786);
xor U29923 (N_29923,N_27625,N_27338);
xor U29924 (N_29924,N_26345,N_27775);
xor U29925 (N_29925,N_26144,N_27301);
xnor U29926 (N_29926,N_26495,N_26419);
and U29927 (N_29927,N_26812,N_27664);
nor U29928 (N_29928,N_27390,N_26926);
nor U29929 (N_29929,N_27468,N_27653);
nor U29930 (N_29930,N_27616,N_27208);
nand U29931 (N_29931,N_27053,N_27504);
nand U29932 (N_29932,N_26533,N_26220);
nor U29933 (N_29933,N_26881,N_26334);
and U29934 (N_29934,N_27540,N_27806);
nand U29935 (N_29935,N_26004,N_27318);
xnor U29936 (N_29936,N_26303,N_27141);
nor U29937 (N_29937,N_27456,N_26130);
nor U29938 (N_29938,N_27477,N_26613);
nor U29939 (N_29939,N_26428,N_26764);
and U29940 (N_29940,N_26372,N_26360);
nor U29941 (N_29941,N_27353,N_26715);
xor U29942 (N_29942,N_26424,N_27788);
xnor U29943 (N_29943,N_27524,N_27818);
xnor U29944 (N_29944,N_26629,N_27269);
or U29945 (N_29945,N_27253,N_27631);
nor U29946 (N_29946,N_26961,N_27447);
or U29947 (N_29947,N_26651,N_27292);
nor U29948 (N_29948,N_27106,N_27940);
and U29949 (N_29949,N_27962,N_27759);
xor U29950 (N_29950,N_27052,N_27653);
xor U29951 (N_29951,N_26997,N_26780);
nand U29952 (N_29952,N_26726,N_27271);
nand U29953 (N_29953,N_26040,N_27906);
xnor U29954 (N_29954,N_26953,N_26157);
and U29955 (N_29955,N_27717,N_26921);
xor U29956 (N_29956,N_27756,N_26560);
nor U29957 (N_29957,N_27439,N_27771);
xnor U29958 (N_29958,N_27764,N_26855);
nor U29959 (N_29959,N_26107,N_27130);
nand U29960 (N_29960,N_27724,N_26092);
or U29961 (N_29961,N_26354,N_26753);
nor U29962 (N_29962,N_26173,N_27785);
nor U29963 (N_29963,N_26172,N_27357);
nor U29964 (N_29964,N_27059,N_27441);
xnor U29965 (N_29965,N_27418,N_26300);
and U29966 (N_29966,N_26630,N_26068);
xor U29967 (N_29967,N_27407,N_26626);
xor U29968 (N_29968,N_27866,N_26235);
or U29969 (N_29969,N_27796,N_27010);
xor U29970 (N_29970,N_26815,N_27719);
nand U29971 (N_29971,N_27839,N_27172);
xnor U29972 (N_29972,N_26636,N_27244);
and U29973 (N_29973,N_27195,N_26580);
nand U29974 (N_29974,N_26361,N_26946);
nand U29975 (N_29975,N_26786,N_27050);
nor U29976 (N_29976,N_27324,N_26194);
or U29977 (N_29977,N_26954,N_26635);
nor U29978 (N_29978,N_26853,N_27788);
nor U29979 (N_29979,N_26510,N_26779);
nor U29980 (N_29980,N_27327,N_26316);
or U29981 (N_29981,N_27166,N_26353);
nor U29982 (N_29982,N_26643,N_27849);
or U29983 (N_29983,N_26621,N_27303);
and U29984 (N_29984,N_26668,N_27999);
xor U29985 (N_29985,N_26178,N_27300);
nand U29986 (N_29986,N_26757,N_26915);
or U29987 (N_29987,N_26647,N_26718);
nand U29988 (N_29988,N_26969,N_27804);
or U29989 (N_29989,N_26835,N_26959);
nor U29990 (N_29990,N_26292,N_26566);
or U29991 (N_29991,N_26971,N_26855);
or U29992 (N_29992,N_26079,N_27909);
xnor U29993 (N_29993,N_26855,N_27572);
nand U29994 (N_29994,N_27177,N_26044);
nand U29995 (N_29995,N_27911,N_27788);
nor U29996 (N_29996,N_26191,N_26441);
nand U29997 (N_29997,N_26707,N_26065);
xnor U29998 (N_29998,N_26888,N_27775);
nor U29999 (N_29999,N_27787,N_27318);
nand UO_0 (O_0,N_28979,N_29024);
xor UO_1 (O_1,N_29467,N_28772);
or UO_2 (O_2,N_29277,N_29196);
nand UO_3 (O_3,N_29661,N_28380);
nor UO_4 (O_4,N_28567,N_29838);
and UO_5 (O_5,N_29805,N_28006);
nor UO_6 (O_6,N_28737,N_28994);
nand UO_7 (O_7,N_28671,N_29137);
xor UO_8 (O_8,N_28585,N_29411);
nand UO_9 (O_9,N_29179,N_28487);
or UO_10 (O_10,N_28693,N_28414);
nor UO_11 (O_11,N_29729,N_28322);
and UO_12 (O_12,N_29256,N_28013);
nor UO_13 (O_13,N_28631,N_29380);
and UO_14 (O_14,N_29533,N_28827);
xnor UO_15 (O_15,N_29642,N_28919);
or UO_16 (O_16,N_29781,N_29594);
nor UO_17 (O_17,N_29262,N_29392);
nand UO_18 (O_18,N_28345,N_29723);
nand UO_19 (O_19,N_29051,N_29561);
or UO_20 (O_20,N_29842,N_29113);
nand UO_21 (O_21,N_29635,N_29992);
or UO_22 (O_22,N_29471,N_28929);
nor UO_23 (O_23,N_29688,N_29798);
nand UO_24 (O_24,N_29224,N_29509);
or UO_25 (O_25,N_28313,N_29824);
or UO_26 (O_26,N_29002,N_28564);
nor UO_27 (O_27,N_29271,N_29220);
and UO_28 (O_28,N_28267,N_29036);
and UO_29 (O_29,N_29765,N_28294);
nand UO_30 (O_30,N_28799,N_28166);
and UO_31 (O_31,N_29935,N_29187);
or UO_32 (O_32,N_29840,N_29858);
nand UO_33 (O_33,N_28675,N_29214);
nor UO_34 (O_34,N_28057,N_29607);
nand UO_35 (O_35,N_28682,N_28185);
xor UO_36 (O_36,N_29662,N_29861);
or UO_37 (O_37,N_28582,N_29904);
nor UO_38 (O_38,N_28477,N_28757);
or UO_39 (O_39,N_28239,N_29261);
nand UO_40 (O_40,N_29215,N_29851);
or UO_41 (O_41,N_29993,N_29229);
nand UO_42 (O_42,N_29931,N_29756);
xnor UO_43 (O_43,N_29628,N_29061);
and UO_44 (O_44,N_29343,N_29988);
and UO_45 (O_45,N_28430,N_28999);
nand UO_46 (O_46,N_28225,N_28066);
and UO_47 (O_47,N_29245,N_28077);
nor UO_48 (O_48,N_28819,N_28741);
nor UO_49 (O_49,N_28847,N_29543);
and UO_50 (O_50,N_29979,N_29048);
or UO_51 (O_51,N_28695,N_29355);
xnor UO_52 (O_52,N_29600,N_28454);
and UO_53 (O_53,N_28945,N_29735);
xnor UO_54 (O_54,N_28094,N_28424);
xnor UO_55 (O_55,N_28636,N_28968);
xnor UO_56 (O_56,N_28680,N_28546);
nand UO_57 (O_57,N_28977,N_28056);
xor UO_58 (O_58,N_29243,N_28782);
nand UO_59 (O_59,N_28502,N_28237);
xnor UO_60 (O_60,N_28998,N_28769);
nor UO_61 (O_61,N_29385,N_29717);
nand UO_62 (O_62,N_28468,N_28422);
xor UO_63 (O_63,N_29612,N_29453);
or UO_64 (O_64,N_28807,N_28788);
xor UO_65 (O_65,N_29026,N_28236);
and UO_66 (O_66,N_28025,N_28660);
and UO_67 (O_67,N_28051,N_29323);
and UO_68 (O_68,N_28561,N_28440);
nand UO_69 (O_69,N_29198,N_28831);
nor UO_70 (O_70,N_28771,N_28674);
and UO_71 (O_71,N_28640,N_28551);
and UO_72 (O_72,N_29052,N_29529);
and UO_73 (O_73,N_29225,N_29079);
xnor UO_74 (O_74,N_28939,N_29440);
or UO_75 (O_75,N_29219,N_28405);
or UO_76 (O_76,N_29035,N_29577);
xnor UO_77 (O_77,N_28230,N_29269);
nor UO_78 (O_78,N_29047,N_29917);
and UO_79 (O_79,N_29502,N_29932);
or UO_80 (O_80,N_28738,N_29918);
xnor UO_81 (O_81,N_29557,N_29313);
xnor UO_82 (O_82,N_29981,N_28492);
or UO_83 (O_83,N_29156,N_29307);
and UO_84 (O_84,N_29815,N_28453);
nand UO_85 (O_85,N_29518,N_28081);
nand UO_86 (O_86,N_28262,N_28235);
or UO_87 (O_87,N_29724,N_29574);
or UO_88 (O_88,N_28904,N_29500);
nor UO_89 (O_89,N_29360,N_28909);
nor UO_90 (O_90,N_28529,N_29673);
or UO_91 (O_91,N_29279,N_28751);
nor UO_92 (O_92,N_29701,N_29882);
and UO_93 (O_93,N_28249,N_29161);
xor UO_94 (O_94,N_28455,N_28017);
and UO_95 (O_95,N_28438,N_28285);
nand UO_96 (O_96,N_29510,N_29326);
or UO_97 (O_97,N_28877,N_28951);
nor UO_98 (O_98,N_29045,N_29758);
xor UO_99 (O_99,N_28822,N_28205);
and UO_100 (O_100,N_28961,N_28154);
nand UO_101 (O_101,N_28341,N_29439);
xor UO_102 (O_102,N_29327,N_28570);
nand UO_103 (O_103,N_29297,N_29370);
or UO_104 (O_104,N_28777,N_29081);
nor UO_105 (O_105,N_28713,N_29302);
nand UO_106 (O_106,N_28717,N_28974);
nand UO_107 (O_107,N_28645,N_28947);
nand UO_108 (O_108,N_28161,N_28656);
xor UO_109 (O_109,N_29967,N_28084);
and UO_110 (O_110,N_29421,N_28736);
xnor UO_111 (O_111,N_28203,N_28548);
and UO_112 (O_112,N_29321,N_28124);
and UO_113 (O_113,N_29725,N_28069);
xnor UO_114 (O_114,N_28036,N_28727);
xor UO_115 (O_115,N_28629,N_28557);
and UO_116 (O_116,N_29873,N_29278);
xor UO_117 (O_117,N_29328,N_29531);
nor UO_118 (O_118,N_29378,N_28890);
nand UO_119 (O_119,N_28197,N_28286);
xnor UO_120 (O_120,N_29997,N_28334);
or UO_121 (O_121,N_29076,N_29903);
or UO_122 (O_122,N_28292,N_29107);
nor UO_123 (O_123,N_29127,N_29887);
nand UO_124 (O_124,N_28490,N_28190);
or UO_125 (O_125,N_28463,N_28993);
or UO_126 (O_126,N_29120,N_29777);
nor UO_127 (O_127,N_29016,N_28129);
nor UO_128 (O_128,N_29787,N_29938);
or UO_129 (O_129,N_28307,N_29569);
nor UO_130 (O_130,N_28689,N_28633);
xor UO_131 (O_131,N_28001,N_28785);
or UO_132 (O_132,N_29912,N_29200);
nor UO_133 (O_133,N_28834,N_28789);
nor UO_134 (O_134,N_29959,N_28913);
xor UO_135 (O_135,N_28852,N_29715);
nand UO_136 (O_136,N_29428,N_28045);
or UO_137 (O_137,N_29646,N_28469);
and UO_138 (O_138,N_28532,N_28016);
nor UO_139 (O_139,N_29634,N_28378);
and UO_140 (O_140,N_28339,N_29819);
xor UO_141 (O_141,N_29627,N_29964);
xnor UO_142 (O_142,N_28940,N_29940);
or UO_143 (O_143,N_28946,N_29859);
or UO_144 (O_144,N_29828,N_29513);
nand UO_145 (O_145,N_28397,N_28506);
nand UO_146 (O_146,N_29514,N_29281);
xnor UO_147 (O_147,N_29409,N_28406);
xor UO_148 (O_148,N_28315,N_28950);
xor UO_149 (O_149,N_28958,N_28665);
xnor UO_150 (O_150,N_29915,N_29422);
xnor UO_151 (O_151,N_29177,N_29719);
nor UO_152 (O_152,N_28673,N_28677);
or UO_153 (O_153,N_29567,N_29465);
nor UO_154 (O_154,N_28253,N_29546);
xor UO_155 (O_155,N_29386,N_29306);
nor UO_156 (O_156,N_29436,N_29417);
nor UO_157 (O_157,N_28969,N_28290);
and UO_158 (O_158,N_28617,N_28716);
nor UO_159 (O_159,N_29927,N_28905);
nor UO_160 (O_160,N_29208,N_28783);
xnor UO_161 (O_161,N_28486,N_29082);
nand UO_162 (O_162,N_29119,N_29347);
xnor UO_163 (O_163,N_29951,N_28728);
nor UO_164 (O_164,N_28902,N_28120);
or UO_165 (O_165,N_29233,N_29116);
nand UO_166 (O_166,N_28810,N_29794);
nand UO_167 (O_167,N_28431,N_29153);
xnor UO_168 (O_168,N_28376,N_29970);
nor UO_169 (O_169,N_28074,N_29969);
and UO_170 (O_170,N_28357,N_29244);
and UO_171 (O_171,N_28140,N_28667);
xnor UO_172 (O_172,N_28442,N_29276);
or UO_173 (O_173,N_29021,N_28021);
nor UO_174 (O_174,N_28257,N_28752);
or UO_175 (O_175,N_28820,N_29192);
xnor UO_176 (O_176,N_28123,N_29936);
nor UO_177 (O_177,N_29638,N_29727);
and UO_178 (O_178,N_29141,N_28770);
or UO_179 (O_179,N_29665,N_29590);
nor UO_180 (O_180,N_29696,N_28155);
nand UO_181 (O_181,N_29636,N_28600);
and UO_182 (O_182,N_29772,N_28609);
xor UO_183 (O_183,N_29681,N_28372);
nor UO_184 (O_184,N_28812,N_28196);
nor UO_185 (O_185,N_29525,N_29459);
and UO_186 (O_186,N_28034,N_29318);
or UO_187 (O_187,N_28912,N_29448);
nor UO_188 (O_188,N_28112,N_28386);
and UO_189 (O_189,N_29579,N_29771);
and UO_190 (O_190,N_29041,N_29133);
xor UO_191 (O_191,N_28063,N_28152);
nor UO_192 (O_192,N_29645,N_28348);
and UO_193 (O_193,N_28476,N_29478);
and UO_194 (O_194,N_29158,N_29901);
or UO_195 (O_195,N_29913,N_28448);
nand UO_196 (O_196,N_28776,N_28275);
nor UO_197 (O_197,N_29253,N_29788);
nand UO_198 (O_198,N_28458,N_29703);
and UO_199 (O_199,N_28457,N_29864);
and UO_200 (O_200,N_28306,N_29013);
or UO_201 (O_201,N_28516,N_28061);
xor UO_202 (O_202,N_28247,N_29706);
or UO_203 (O_203,N_28841,N_28435);
xnor UO_204 (O_204,N_29697,N_29194);
nor UO_205 (O_205,N_28138,N_29548);
nor UO_206 (O_206,N_29739,N_29446);
and UO_207 (O_207,N_29713,N_28602);
nor UO_208 (O_208,N_28298,N_29989);
or UO_209 (O_209,N_28724,N_29625);
and UO_210 (O_210,N_29110,N_29080);
nand UO_211 (O_211,N_29770,N_28581);
nand UO_212 (O_212,N_29660,N_28580);
and UO_213 (O_213,N_29234,N_28542);
nor UO_214 (O_214,N_28641,N_29702);
and UO_215 (O_215,N_28355,N_29515);
or UO_216 (O_216,N_28989,N_29049);
nand UO_217 (O_217,N_28527,N_29894);
or UO_218 (O_218,N_29403,N_29804);
or UO_219 (O_219,N_29779,N_29228);
xor UO_220 (O_220,N_28917,N_28702);
and UO_221 (O_221,N_28118,N_29493);
and UO_222 (O_222,N_29068,N_29596);
nand UO_223 (O_223,N_28217,N_28343);
or UO_224 (O_224,N_29737,N_29100);
and UO_225 (O_225,N_28539,N_29260);
xor UO_226 (O_226,N_28305,N_29420);
nand UO_227 (O_227,N_28649,N_28857);
xnor UO_228 (O_228,N_29570,N_29438);
nor UO_229 (O_229,N_29868,N_29591);
and UO_230 (O_230,N_29408,N_28489);
nand UO_231 (O_231,N_28027,N_29848);
nand UO_232 (O_232,N_28743,N_28896);
nand UO_233 (O_233,N_29659,N_28279);
and UO_234 (O_234,N_28332,N_28478);
xnor UO_235 (O_235,N_29773,N_28774);
xnor UO_236 (O_236,N_29144,N_29890);
nand UO_237 (O_237,N_29267,N_28790);
nand UO_238 (O_238,N_29855,N_28050);
or UO_239 (O_239,N_28157,N_28832);
xor UO_240 (O_240,N_29980,N_28775);
xnor UO_241 (O_241,N_29352,N_29163);
or UO_242 (O_242,N_28042,N_28957);
and UO_243 (O_243,N_28591,N_28523);
and UO_244 (O_244,N_29391,N_28528);
xor UO_245 (O_245,N_28975,N_28071);
or UO_246 (O_246,N_28250,N_29248);
nor UO_247 (O_247,N_28662,N_28663);
nand UO_248 (O_248,N_28972,N_28479);
nor UO_249 (O_249,N_29810,N_29811);
nor UO_250 (O_250,N_29084,N_29022);
or UO_251 (O_251,N_29106,N_29669);
and UO_252 (O_252,N_28568,N_28171);
nor UO_253 (O_253,N_28518,N_29169);
nand UO_254 (O_254,N_28566,N_28211);
xor UO_255 (O_255,N_28657,N_29270);
xnor UO_256 (O_256,N_29695,N_28329);
nand UO_257 (O_257,N_29379,N_29841);
xnor UO_258 (O_258,N_29199,N_29476);
nor UO_259 (O_259,N_28956,N_28614);
nand UO_260 (O_260,N_29540,N_29242);
and UO_261 (O_261,N_29535,N_29926);
nand UO_262 (O_262,N_28382,N_29406);
nand UO_263 (O_263,N_28330,N_28385);
xor UO_264 (O_264,N_29733,N_29652);
nor UO_265 (O_265,N_28089,N_28098);
nor UO_266 (O_266,N_28840,N_29507);
and UO_267 (O_267,N_28366,N_28079);
or UO_268 (O_268,N_28470,N_29558);
nor UO_269 (O_269,N_28806,N_28670);
xnor UO_270 (O_270,N_28589,N_28108);
and UO_271 (O_271,N_29900,N_28874);
and UO_272 (O_272,N_28018,N_29629);
and UO_273 (O_273,N_28668,N_29497);
nor UO_274 (O_274,N_29680,N_29419);
or UO_275 (O_275,N_29221,N_28395);
nor UO_276 (O_276,N_29663,N_29206);
nor UO_277 (O_277,N_29827,N_29599);
nand UO_278 (O_278,N_28110,N_28699);
nand UO_279 (O_279,N_28525,N_28400);
nor UO_280 (O_280,N_29028,N_29223);
xnor UO_281 (O_281,N_28274,N_29875);
xnor UO_282 (O_282,N_29499,N_28630);
nor UO_283 (O_283,N_29909,N_29466);
or UO_284 (O_284,N_28714,N_29043);
xnor UO_285 (O_285,N_29552,N_28802);
xnor UO_286 (O_286,N_29232,N_29231);
nand UO_287 (O_287,N_28204,N_28418);
nor UO_288 (O_288,N_28182,N_28475);
nand UO_289 (O_289,N_28976,N_28394);
nor UO_290 (O_290,N_29132,N_29010);
and UO_291 (O_291,N_29304,N_28595);
nand UO_292 (O_292,N_28881,N_29186);
nor UO_293 (O_293,N_29424,N_28870);
or UO_294 (O_294,N_29367,N_28121);
or UO_295 (O_295,N_29519,N_28747);
nor UO_296 (O_296,N_28715,N_28535);
nor UO_297 (O_297,N_28384,N_29450);
and UO_298 (O_298,N_28579,N_29000);
xnor UO_299 (O_299,N_28359,N_29498);
nand UO_300 (O_300,N_29382,N_28613);
or UO_301 (O_301,N_29705,N_28364);
nand UO_302 (O_302,N_28371,N_29001);
nor UO_303 (O_303,N_28337,N_28555);
xnor UO_304 (O_304,N_29291,N_29009);
or UO_305 (O_305,N_28396,N_28652);
nand UO_306 (O_306,N_28268,N_29203);
xor UO_307 (O_307,N_28335,N_28748);
xnor UO_308 (O_308,N_29053,N_29290);
or UO_309 (O_309,N_29074,N_29831);
and UO_310 (O_310,N_28260,N_28611);
xnor UO_311 (O_311,N_29844,N_29822);
xor UO_312 (O_312,N_29311,N_28593);
xor UO_313 (O_313,N_29566,N_28873);
nand UO_314 (O_314,N_28970,N_28966);
xnor UO_315 (O_315,N_29331,N_28494);
nand UO_316 (O_316,N_28134,N_29397);
or UO_317 (O_317,N_28866,N_28240);
or UO_318 (O_318,N_28046,N_28472);
nor UO_319 (O_319,N_29251,N_29769);
nor UO_320 (O_320,N_29458,N_28853);
or UO_321 (O_321,N_29934,N_29835);
nor UO_322 (O_322,N_29941,N_28584);
and UO_323 (O_323,N_28503,N_29730);
nor UO_324 (O_324,N_29005,N_28035);
nor UO_325 (O_325,N_28948,N_28316);
xnor UO_326 (O_326,N_29171,N_29806);
nand UO_327 (O_327,N_29623,N_29728);
and UO_328 (O_328,N_29155,N_28449);
nor UO_329 (O_329,N_28310,N_28484);
or UO_330 (O_330,N_28924,N_29197);
or UO_331 (O_331,N_29098,N_28113);
or UO_332 (O_332,N_29309,N_28758);
nand UO_333 (O_333,N_29490,N_28280);
and UO_334 (O_334,N_28910,N_29475);
nand UO_335 (O_335,N_28003,N_28732);
nand UO_336 (O_336,N_29834,N_28465);
nor UO_337 (O_337,N_29965,N_28508);
or UO_338 (O_338,N_28511,N_28342);
and UO_339 (O_339,N_28590,N_29956);
or UO_340 (O_340,N_29172,N_28425);
or UO_341 (O_341,N_29587,N_29335);
and UO_342 (O_342,N_29626,N_29320);
or UO_343 (O_343,N_28720,N_28263);
and UO_344 (O_344,N_29897,N_29666);
nand UO_345 (O_345,N_28328,N_28963);
and UO_346 (O_346,N_28861,N_28485);
nand UO_347 (O_347,N_29040,N_29130);
nand UO_348 (O_348,N_29863,N_29886);
nand UO_349 (O_349,N_28420,N_29182);
xor UO_350 (O_350,N_28181,N_28914);
and UO_351 (O_351,N_29889,N_29978);
nand UO_352 (O_352,N_28080,N_29671);
nor UO_353 (O_353,N_28055,N_29131);
or UO_354 (O_354,N_29791,N_28272);
xor UO_355 (O_355,N_28666,N_29390);
nand UO_356 (O_356,N_29383,N_29785);
nor UO_357 (O_357,N_29204,N_29692);
nand UO_358 (O_358,N_28044,N_28314);
nor UO_359 (O_359,N_29038,N_29550);
or UO_360 (O_360,N_28706,N_28612);
xor UO_361 (O_361,N_28698,N_28090);
and UO_362 (O_362,N_28303,N_28251);
nor UO_363 (O_363,N_28596,N_29174);
nor UO_364 (O_364,N_28126,N_29945);
or UO_365 (O_365,N_29148,N_28065);
nor UO_366 (O_366,N_29126,N_29807);
xnor UO_367 (O_367,N_28628,N_29617);
nand UO_368 (O_368,N_29273,N_28928);
and UO_369 (O_369,N_28172,N_28809);
or UO_370 (O_370,N_29122,N_29150);
and UO_371 (O_371,N_28048,N_28022);
nand UO_372 (O_372,N_28558,N_28007);
or UO_373 (O_373,N_28416,N_29745);
nor UO_374 (O_374,N_28029,N_29712);
and UO_375 (O_375,N_29162,N_28773);
xor UO_376 (O_376,N_28212,N_29795);
and UO_377 (O_377,N_29991,N_28986);
nor UO_378 (O_378,N_29103,N_29504);
xor UO_379 (O_379,N_29287,N_28616);
nor UO_380 (O_380,N_29207,N_28493);
xor UO_381 (O_381,N_28004,N_29820);
nand UO_382 (O_382,N_29373,N_29305);
nor UO_383 (O_383,N_28209,N_28646);
xnor UO_384 (O_384,N_29289,N_28183);
nand UO_385 (O_385,N_28658,N_28891);
or UO_386 (O_386,N_29966,N_28199);
and UO_387 (O_387,N_28410,N_29812);
and UO_388 (O_388,N_29709,N_29093);
xor UO_389 (O_389,N_29537,N_28565);
nor UO_390 (O_390,N_29686,N_29025);
nand UO_391 (O_391,N_28606,N_29947);
and UO_392 (O_392,N_29878,N_28886);
nand UO_393 (O_393,N_29601,N_29075);
xor UO_394 (O_394,N_28892,N_29764);
nor UO_395 (O_395,N_29292,N_29799);
xnor UO_396 (O_396,N_29865,N_29974);
nor UO_397 (O_397,N_28278,N_29065);
nand UO_398 (O_398,N_29610,N_29860);
or UO_399 (O_399,N_28632,N_28935);
nand UO_400 (O_400,N_28683,N_28882);
nand UO_401 (O_401,N_29263,N_28749);
xor UO_402 (O_402,N_29029,N_29622);
nor UO_403 (O_403,N_28445,N_28547);
nand UO_404 (O_404,N_28160,N_28811);
nand UO_405 (O_405,N_28526,N_28162);
xnor UO_406 (O_406,N_29874,N_29939);
xor UO_407 (O_407,N_28839,N_28597);
nor UO_408 (O_408,N_29388,N_28026);
and UO_409 (O_409,N_29949,N_29252);
nand UO_410 (O_410,N_29374,N_28407);
or UO_411 (O_411,N_29866,N_29693);
xnor UO_412 (O_412,N_28696,N_29264);
and UO_413 (O_413,N_29255,N_28762);
nor UO_414 (O_414,N_29463,N_28638);
nor UO_415 (O_415,N_28030,N_29054);
nand UO_416 (O_416,N_29527,N_28184);
and UO_417 (O_417,N_28813,N_29030);
nand UO_418 (O_418,N_28867,N_29907);
nor UO_419 (O_419,N_29571,N_29760);
or UO_420 (O_420,N_28232,N_29325);
nand UO_421 (O_421,N_29637,N_28784);
or UO_422 (O_422,N_28605,N_28893);
xor UO_423 (O_423,N_28200,N_29451);
xor UO_424 (O_424,N_28556,N_29209);
or UO_425 (O_425,N_28571,N_28150);
and UO_426 (O_426,N_29353,N_28223);
or UO_427 (O_427,N_29145,N_29303);
nor UO_428 (O_428,N_29259,N_29412);
and UO_429 (O_429,N_29749,N_29615);
xnor UO_430 (O_430,N_29337,N_28346);
nor UO_431 (O_431,N_29598,N_29593);
xor UO_432 (O_432,N_29405,N_29096);
nand UO_433 (O_433,N_28815,N_29998);
nor UO_434 (O_434,N_29524,N_29160);
nor UO_435 (O_435,N_29586,N_28091);
nor UO_436 (O_436,N_29181,N_29797);
nand UO_437 (O_437,N_29790,N_29332);
or UO_438 (O_438,N_28973,N_28297);
nand UO_439 (O_439,N_28903,N_28655);
and UO_440 (O_440,N_29006,N_28381);
xor UO_441 (O_441,N_28889,N_28930);
nand UO_442 (O_442,N_29101,N_29619);
and UO_443 (O_443,N_28195,N_29520);
and UO_444 (O_444,N_28273,N_28745);
and UO_445 (O_445,N_28862,N_28876);
nor UO_446 (O_446,N_28587,N_29154);
and UO_447 (O_447,N_28488,N_28243);
and UO_448 (O_448,N_28133,N_28635);
nor UO_449 (O_449,N_28786,N_29694);
and UO_450 (O_450,N_29809,N_28780);
or UO_451 (O_451,N_28353,N_28433);
or UO_452 (O_452,N_28678,N_28779);
nor UO_453 (O_453,N_28869,N_29193);
xnor UO_454 (O_454,N_28988,N_28058);
or UO_455 (O_455,N_28996,N_29222);
and UO_456 (O_456,N_28039,N_28664);
nor UO_457 (O_457,N_29275,N_28684);
nor UO_458 (O_458,N_28426,N_29895);
nor UO_459 (O_459,N_28643,N_28175);
nor UO_460 (O_460,N_29672,N_28916);
and UO_461 (O_461,N_29589,N_29340);
or UO_462 (O_462,N_28710,N_29454);
nand UO_463 (O_463,N_29908,N_28146);
nand UO_464 (O_464,N_28746,N_29676);
xnor UO_465 (O_465,N_28825,N_29948);
and UO_466 (O_466,N_28049,N_29086);
nor UO_467 (O_467,N_29902,N_28644);
xor UO_468 (O_468,N_29517,N_29783);
and UO_469 (O_469,N_28377,N_29766);
nand UO_470 (O_470,N_28088,N_29891);
nand UO_471 (O_471,N_28207,N_28942);
nor UO_472 (O_472,N_28441,N_29856);
xor UO_473 (O_473,N_29286,N_29630);
nand UO_474 (O_474,N_28661,N_29432);
nand UO_475 (O_475,N_29176,N_29508);
and UO_476 (O_476,N_28742,N_29836);
and UO_477 (O_477,N_29687,N_28402);
and UO_478 (O_478,N_28792,N_28221);
nor UO_479 (O_479,N_28131,N_29070);
or UO_480 (O_480,N_29125,N_28797);
nand UO_481 (O_481,N_29711,N_28246);
nor UO_482 (O_482,N_29042,N_28214);
and UO_483 (O_483,N_28020,N_29031);
and UO_484 (O_484,N_28575,N_29872);
or UO_485 (O_485,N_28254,N_28541);
nand UO_486 (O_486,N_29962,N_29554);
or UO_487 (O_487,N_28300,N_29456);
nor UO_488 (O_488,N_28115,N_29716);
nand UO_489 (O_489,N_28639,N_28023);
xor UO_490 (O_490,N_28417,N_29722);
nor UO_491 (O_491,N_29604,N_29847);
nor UO_492 (O_492,N_28740,N_29123);
or UO_493 (O_493,N_28444,N_28829);
or UO_494 (O_494,N_28507,N_28156);
or UO_495 (O_495,N_28846,N_29410);
nor UO_496 (O_496,N_28923,N_28352);
xor UO_497 (O_497,N_29611,N_28854);
and UO_498 (O_498,N_29972,N_29892);
xnor UO_499 (O_499,N_29195,N_28293);
nor UO_500 (O_500,N_29656,N_28351);
nor UO_501 (O_501,N_28685,N_28234);
nand UO_502 (O_502,N_29977,N_29060);
and UO_503 (O_503,N_29987,N_28466);
nor UO_504 (O_504,N_28897,N_28835);
nand UO_505 (O_505,N_29862,N_28573);
nor UO_506 (O_506,N_28722,N_29315);
nand UO_507 (O_507,N_28031,N_29377);
nor UO_508 (O_508,N_28096,N_28202);
nor UO_509 (O_509,N_29914,N_29414);
xnor UO_510 (O_510,N_29653,N_28513);
nand UO_511 (O_511,N_29034,N_28875);
and UO_512 (O_512,N_29682,N_29821);
nor UO_513 (O_513,N_28075,N_29501);
or UO_514 (O_514,N_28721,N_28540);
nand UO_515 (O_515,N_28354,N_28295);
nand UO_516 (O_516,N_29565,N_28848);
xnor UO_517 (O_517,N_28533,N_29830);
nand UO_518 (O_518,N_28347,N_28145);
or UO_519 (O_519,N_28514,N_29763);
nor UO_520 (O_520,N_29376,N_29298);
and UO_521 (O_521,N_29545,N_29789);
nor UO_522 (O_522,N_28119,N_28756);
nand UO_523 (O_523,N_29995,N_28149);
xnor UO_524 (O_524,N_28317,N_29506);
or UO_525 (O_525,N_29469,N_28467);
nand UO_526 (O_526,N_28451,N_28933);
nor UO_527 (O_527,N_29679,N_29210);
nand UO_528 (O_528,N_28625,N_29039);
nor UO_529 (O_529,N_29067,N_29090);
and UO_530 (O_530,N_29633,N_28167);
nand UO_531 (O_531,N_28767,N_29272);
nand UO_532 (O_532,N_29973,N_29528);
nand UO_533 (O_533,N_29778,N_28002);
and UO_534 (O_534,N_28097,N_28550);
and UO_535 (O_535,N_29020,N_28650);
and UO_536 (O_536,N_29063,N_28830);
or UO_537 (O_537,N_29217,N_28864);
and UO_538 (O_538,N_28193,N_29944);
and UO_539 (O_539,N_28623,N_28208);
nand UO_540 (O_540,N_28281,N_28130);
nor UO_541 (O_541,N_28694,N_28955);
nand UO_542 (O_542,N_28192,N_28311);
nor UO_543 (O_543,N_28672,N_28604);
nor UO_544 (O_544,N_28858,N_28389);
or UO_545 (O_545,N_28898,N_29280);
nor UO_546 (O_546,N_28434,N_29879);
nor UO_547 (O_547,N_29460,N_29247);
nor UO_548 (O_548,N_28496,N_29108);
nor UO_549 (O_549,N_29675,N_28095);
and UO_550 (O_550,N_28911,N_29952);
or UO_551 (O_551,N_28900,N_29135);
xnor UO_552 (O_552,N_29183,N_29542);
nand UO_553 (O_553,N_29808,N_28187);
nand UO_554 (O_554,N_29818,N_28288);
or UO_555 (O_555,N_28865,N_29954);
or UO_556 (O_556,N_29293,N_28082);
or UO_557 (O_557,N_28064,N_28141);
or UO_558 (O_558,N_29971,N_28559);
or UO_559 (O_559,N_29562,N_29282);
nor UO_560 (O_560,N_29572,N_28871);
or UO_561 (O_561,N_29905,N_28367);
xor UO_562 (O_562,N_28070,N_29019);
nand UO_563 (O_563,N_29532,N_29342);
nor UO_564 (O_564,N_28087,N_29658);
or UO_565 (O_565,N_29776,N_28562);
or UO_566 (O_566,N_29556,N_28495);
nand UO_567 (O_567,N_29968,N_29404);
nand UO_568 (O_568,N_29898,N_29826);
nand UO_569 (O_569,N_28040,N_28392);
and UO_570 (O_570,N_28586,N_29761);
or UO_571 (O_571,N_28231,N_29462);
nand UO_572 (O_572,N_28104,N_29111);
nand UO_573 (O_573,N_28679,N_29151);
nand UO_574 (O_574,N_29606,N_29857);
nand UO_575 (O_575,N_29768,N_29429);
and UO_576 (O_576,N_28447,N_28015);
xnor UO_577 (O_577,N_28787,N_29316);
nor UO_578 (O_578,N_28428,N_29759);
xnor UO_579 (O_579,N_28178,N_29356);
or UO_580 (O_580,N_28860,N_29236);
xnor UO_581 (O_581,N_29365,N_29455);
xor UO_582 (O_582,N_29444,N_29592);
xor UO_583 (O_583,N_28755,N_28878);
xor UO_584 (O_584,N_28287,N_29308);
or UO_585 (O_585,N_29699,N_29829);
and UO_586 (O_586,N_28326,N_28296);
and UO_587 (O_587,N_29620,N_29505);
and UO_588 (O_588,N_29963,N_29608);
and UO_589 (O_589,N_29319,N_28062);
nand UO_590 (O_590,N_28545,N_28450);
and UO_591 (O_591,N_29387,N_28691);
and UO_592 (O_592,N_29576,N_28560);
nor UO_593 (O_593,N_29538,N_28944);
and UO_594 (O_594,N_29910,N_28608);
nor UO_595 (O_595,N_29284,N_29037);
or UO_596 (O_596,N_29984,N_29358);
xor UO_597 (O_597,N_29880,N_28325);
xor UO_598 (O_598,N_28340,N_28137);
nor UO_599 (O_599,N_29477,N_28117);
nand UO_600 (O_600,N_28304,N_29511);
nand UO_601 (O_601,N_28686,N_28333);
nor UO_602 (O_602,N_28443,N_28915);
and UO_603 (O_603,N_29689,N_29916);
nor UO_604 (O_604,N_29893,N_29354);
and UO_605 (O_605,N_29336,N_28255);
xnor UO_606 (O_606,N_29924,N_29407);
nor UO_607 (O_607,N_28116,N_28778);
nor UO_608 (O_608,N_28461,N_28992);
nor UO_609 (O_609,N_28826,N_28967);
nor UO_610 (O_610,N_29457,N_29479);
nor UO_611 (O_611,N_29146,N_28808);
nand UO_612 (O_612,N_28390,N_29014);
and UO_613 (O_613,N_28264,N_28818);
or UO_614 (O_614,N_28517,N_28164);
nand UO_615 (O_615,N_28759,N_28158);
and UO_616 (O_616,N_28086,N_28766);
nor UO_617 (O_617,N_28481,N_29597);
nor UO_618 (O_618,N_28375,N_29957);
xnor UO_619 (O_619,N_28053,N_28266);
xnor UO_620 (O_620,N_28456,N_28768);
and UO_621 (O_621,N_28987,N_29602);
nand UO_622 (O_622,N_29767,N_29568);
xnor UO_623 (O_623,N_29928,N_29003);
xnor UO_624 (O_624,N_29468,N_28114);
and UO_625 (O_625,N_28821,N_29027);
xor UO_626 (O_626,N_28159,N_29257);
nand UO_627 (O_627,N_29441,N_28926);
or UO_628 (O_628,N_28838,N_28981);
xnor UO_629 (O_629,N_28531,N_28530);
nor UO_630 (O_630,N_29464,N_29559);
nor UO_631 (O_631,N_29240,N_29227);
nor UO_632 (O_632,N_29541,N_29147);
nor UO_633 (O_633,N_28510,N_29173);
and UO_634 (O_634,N_28369,N_29551);
and UO_635 (O_635,N_29786,N_28642);
nor UO_636 (O_636,N_29560,N_29483);
nor UO_637 (O_637,N_29534,N_29942);
or UO_638 (O_638,N_28139,N_28324);
nor UO_639 (O_639,N_28588,N_29423);
xor UO_640 (O_640,N_28501,N_29226);
xor UO_641 (O_641,N_29817,N_28270);
and UO_642 (O_642,N_28219,N_28500);
and UO_643 (O_643,N_29950,N_29056);
or UO_644 (O_644,N_29474,N_28242);
nand UO_645 (O_645,N_28920,N_28599);
or UO_646 (O_646,N_29708,N_28735);
nor UO_647 (O_647,N_28959,N_28012);
nor UO_648 (O_648,N_29180,N_29780);
xnor UO_649 (O_649,N_29512,N_28932);
nor UO_650 (O_650,N_29050,N_29188);
nor UO_651 (O_651,N_28092,N_29943);
and UO_652 (O_652,N_28984,N_29563);
xnor UO_653 (O_653,N_29055,N_28291);
xor UO_654 (O_654,N_29762,N_28978);
xor UO_655 (O_655,N_29088,N_28024);
or UO_656 (O_656,N_29632,N_28754);
nand UO_657 (O_657,N_29165,N_28226);
xnor UO_658 (O_658,N_29850,N_28883);
and UO_659 (O_659,N_28879,N_29923);
xor UO_660 (O_660,N_28165,N_29544);
or UO_661 (O_661,N_29491,N_28844);
xor UO_662 (O_662,N_29294,N_28459);
or UO_663 (O_663,N_29044,N_29955);
nand UO_664 (O_664,N_29235,N_29616);
nand UO_665 (O_665,N_28085,N_28198);
nor UO_666 (O_666,N_29329,N_29792);
and UO_667 (O_667,N_29580,N_29667);
xor UO_668 (O_668,N_28460,N_29283);
nand UO_669 (O_669,N_29008,N_28360);
and UO_670 (O_670,N_29250,N_29322);
or UO_671 (O_671,N_29461,N_29721);
nor UO_672 (O_672,N_29480,N_28474);
nand UO_673 (O_673,N_29668,N_29849);
xnor UO_674 (O_674,N_28739,N_28681);
and UO_675 (O_675,N_28823,N_29684);
and UO_676 (O_676,N_29644,N_28067);
nand UO_677 (O_677,N_29876,N_29710);
nor UO_678 (O_678,N_29288,N_28010);
nor UO_679 (O_679,N_28220,N_28624);
nor UO_680 (O_680,N_28076,N_28427);
or UO_681 (O_681,N_28719,N_29846);
nor UO_682 (O_682,N_29138,N_29362);
or UO_683 (O_683,N_28906,N_29023);
xor UO_684 (O_684,N_29032,N_28796);
xnor UO_685 (O_685,N_29285,N_29105);
nor UO_686 (O_686,N_29921,N_29338);
nor UO_687 (O_687,N_29348,N_29212);
and UO_688 (O_688,N_28491,N_29738);
nor UO_689 (O_689,N_28687,N_29241);
nand UO_690 (O_690,N_28569,N_28583);
xnor UO_691 (O_691,N_29946,N_28111);
nand UO_692 (O_692,N_28761,N_28669);
nand UO_693 (O_693,N_29339,N_29521);
and UO_694 (O_694,N_28398,N_28248);
xnor UO_695 (O_695,N_29526,N_28028);
and UO_696 (O_696,N_29919,N_29609);
or UO_697 (O_697,N_29140,N_29384);
xor UO_698 (O_698,N_28990,N_28931);
and UO_699 (O_699,N_29087,N_28194);
or UO_700 (O_700,N_29089,N_28393);
and UO_701 (O_701,N_29481,N_28907);
nor UO_702 (O_702,N_28312,N_29357);
nand UO_703 (O_703,N_29062,N_29345);
nand UO_704 (O_704,N_28701,N_28801);
xor UO_705 (O_705,N_29136,N_28189);
nand UO_706 (O_706,N_28128,N_29922);
xor UO_707 (O_707,N_28805,N_29670);
and UO_708 (O_708,N_29618,N_29482);
or UO_709 (O_709,N_29522,N_29621);
xor UO_710 (O_710,N_28135,N_29832);
nor UO_711 (O_711,N_28318,N_29707);
or UO_712 (O_712,N_28804,N_29058);
xnor UO_713 (O_713,N_28509,N_29986);
and UO_714 (O_714,N_28320,N_29143);
nor UO_715 (O_715,N_29033,N_29802);
or UO_716 (O_716,N_29775,N_29539);
and UO_717 (O_717,N_29547,N_29425);
nand UO_718 (O_718,N_29443,N_28798);
and UO_719 (O_719,N_29743,N_29603);
and UO_720 (O_720,N_29300,N_28991);
and UO_721 (O_721,N_28446,N_28233);
nand UO_722 (O_722,N_28703,N_28041);
xor UO_723 (O_723,N_28621,N_28019);
xor UO_724 (O_724,N_29128,N_28148);
xor UO_725 (O_725,N_29166,N_28794);
nand UO_726 (O_726,N_28093,N_28725);
or UO_727 (O_727,N_28705,N_28421);
xnor UO_728 (O_728,N_29664,N_28188);
and UO_729 (O_729,N_28349,N_28711);
or UO_730 (O_730,N_29426,N_29361);
nor UO_731 (O_731,N_29312,N_28692);
nand UO_732 (O_732,N_29249,N_29213);
xnor UO_733 (O_733,N_29059,N_29012);
and UO_734 (O_734,N_28436,N_29418);
xnor UO_735 (O_735,N_29445,N_28651);
nand UO_736 (O_736,N_28361,N_29317);
xor UO_737 (O_737,N_29640,N_28814);
xor UO_738 (O_738,N_28960,N_28105);
or UO_739 (O_739,N_28554,N_28370);
xor UO_740 (O_740,N_28301,N_28283);
nand UO_741 (O_741,N_29157,N_28309);
and UO_742 (O_742,N_28383,N_29072);
or UO_743 (O_743,N_29185,N_28709);
nand UO_744 (O_744,N_28244,N_29296);
nor UO_745 (O_745,N_28415,N_28100);
xnor UO_746 (O_746,N_28122,N_29310);
nor UO_747 (O_747,N_28868,N_29796);
and UO_748 (O_748,N_28109,N_28008);
xor UO_749 (O_749,N_28052,N_29238);
and UO_750 (O_750,N_29351,N_28938);
or UO_751 (O_751,N_28619,N_29581);
and UO_752 (O_752,N_29985,N_29595);
xnor UO_753 (O_753,N_28522,N_29190);
nor UO_754 (O_754,N_28170,N_29246);
nand UO_755 (O_755,N_28180,N_28411);
or UO_756 (O_756,N_28578,N_29121);
and UO_757 (O_757,N_28817,N_28222);
nand UO_758 (O_758,N_29496,N_28937);
or UO_759 (O_759,N_28936,N_29726);
nand UO_760 (O_760,N_28177,N_28206);
or UO_761 (O_761,N_29333,N_28894);
xnor UO_762 (O_762,N_29793,N_29911);
nand UO_763 (O_763,N_29124,N_29641);
and UO_764 (O_764,N_29413,N_28851);
nor UO_765 (O_765,N_29714,N_28282);
nor UO_766 (O_766,N_28965,N_29452);
nor UO_767 (O_767,N_29314,N_29871);
or UO_768 (O_768,N_29395,N_29734);
nand UO_769 (O_769,N_29129,N_28563);
or UO_770 (O_770,N_28744,N_29349);
xor UO_771 (O_771,N_28437,N_28151);
nand UO_772 (O_772,N_28653,N_28849);
and UO_773 (O_773,N_28688,N_28323);
nand UO_774 (O_774,N_29394,N_28712);
and UO_775 (O_775,N_29091,N_28344);
xor UO_776 (O_776,N_28201,N_29167);
xnor UO_777 (O_777,N_28054,N_28216);
nor UO_778 (O_778,N_28368,N_28136);
nand UO_779 (O_779,N_28952,N_28549);
xor UO_780 (O_780,N_29755,N_29427);
nand UO_781 (O_781,N_29651,N_29751);
nor UO_782 (O_782,N_29752,N_28855);
xnor UO_783 (O_783,N_28391,N_29814);
nand UO_784 (O_784,N_28482,N_29643);
xor UO_785 (O_785,N_29097,N_28038);
or UO_786 (O_786,N_28229,N_29800);
nand UO_787 (O_787,N_28519,N_29268);
nand UO_788 (O_788,N_28765,N_28594);
and UO_789 (O_789,N_28592,N_28356);
and UO_790 (O_790,N_28265,N_29369);
nand UO_791 (O_791,N_28598,N_28011);
and UO_792 (O_792,N_29837,N_29085);
nand UO_793 (O_793,N_29870,N_28763);
nor UO_794 (O_794,N_29555,N_29435);
xor UO_795 (O_795,N_28127,N_28103);
or UO_796 (O_796,N_28419,N_29324);
or UO_797 (O_797,N_29258,N_28388);
xor UO_798 (O_798,N_28338,N_28014);
nor UO_799 (O_799,N_28060,N_29929);
and UO_800 (O_800,N_28163,N_28073);
or UO_801 (O_801,N_29999,N_28601);
and UO_802 (O_802,N_28439,N_29639);
and UO_803 (O_803,N_29690,N_29530);
nor UO_804 (O_804,N_29094,N_29102);
and UO_805 (O_805,N_28289,N_28409);
nand UO_806 (O_806,N_28816,N_28962);
xor UO_807 (O_807,N_28997,N_28277);
xor UO_808 (O_808,N_29488,N_28730);
nand UO_809 (O_809,N_28210,N_28791);
nand UO_810 (O_810,N_28723,N_28985);
or UO_811 (O_811,N_29523,N_28238);
and UO_812 (O_812,N_29578,N_28750);
and UO_813 (O_813,N_29803,N_28464);
or UO_814 (O_814,N_29937,N_28536);
xor UO_815 (O_815,N_28068,N_29416);
nor UO_816 (O_816,N_28704,N_28473);
nor UO_817 (O_817,N_29434,N_28336);
xnor UO_818 (O_818,N_28173,N_28971);
or UO_819 (O_819,N_28483,N_29442);
xnor UO_820 (O_820,N_28452,N_28824);
nand UO_821 (O_821,N_28980,N_28637);
nand UO_822 (O_822,N_28259,N_29990);
nor UO_823 (O_823,N_29698,N_28760);
or UO_824 (O_824,N_29516,N_28143);
nor UO_825 (O_825,N_28659,N_29486);
and UO_826 (O_826,N_28927,N_29104);
and UO_827 (O_827,N_29782,N_28276);
xnor UO_828 (O_828,N_28925,N_29437);
nor UO_829 (O_829,N_29994,N_28700);
nand UO_830 (O_830,N_29266,N_28078);
xor UO_831 (O_831,N_28899,N_29750);
or UO_832 (O_832,N_28690,N_29149);
xnor UO_833 (O_833,N_28726,N_29648);
xor UO_834 (O_834,N_28753,N_28403);
xnor UO_835 (O_835,N_29449,N_28982);
and UO_836 (O_836,N_28885,N_29099);
and UO_837 (O_837,N_28729,N_29400);
and UO_838 (O_838,N_29585,N_28618);
or UO_839 (O_839,N_28512,N_29657);
or UO_840 (O_840,N_28498,N_29433);
or UO_841 (O_841,N_28697,N_29211);
xor UO_842 (O_842,N_28627,N_29447);
or UO_843 (O_843,N_29736,N_28099);
nor UO_844 (O_844,N_29845,N_28227);
or UO_845 (O_845,N_29732,N_29114);
and UO_846 (O_846,N_28954,N_29801);
and UO_847 (O_847,N_29057,N_28901);
xor UO_848 (O_848,N_29784,N_28224);
xnor UO_849 (O_849,N_29678,N_28032);
nand UO_850 (O_850,N_29553,N_29346);
or UO_851 (O_851,N_28922,N_28520);
and UO_852 (O_852,N_29007,N_28471);
nor UO_853 (O_853,N_29920,N_28228);
nand UO_854 (O_854,N_29189,N_29896);
xor UO_855 (O_855,N_29877,N_28934);
and UO_856 (O_856,N_28828,N_29389);
xor UO_857 (O_857,N_29757,N_28102);
nand UO_858 (O_858,N_29549,N_28995);
and UO_859 (O_859,N_28949,N_28350);
and UO_860 (O_860,N_28321,N_29301);
xnor UO_861 (O_861,N_28072,N_29334);
and UO_862 (O_862,N_28107,N_29064);
nand UO_863 (O_863,N_29774,N_29078);
nand UO_864 (O_864,N_29092,N_29564);
nand UO_865 (O_865,N_29624,N_29184);
and UO_866 (O_866,N_28284,N_28731);
xor UO_867 (O_867,N_29073,N_29274);
nand UO_868 (O_868,N_29982,N_29740);
nand UO_869 (O_869,N_28374,N_28918);
xnor UO_870 (O_870,N_28404,N_28308);
nor UO_871 (O_871,N_29605,N_29674);
or UO_872 (O_872,N_29823,N_29359);
nor UO_873 (O_873,N_29492,N_28941);
and UO_874 (O_874,N_29168,N_28880);
and UO_875 (O_875,N_29396,N_28215);
or UO_876 (O_876,N_28363,N_28953);
xor UO_877 (O_877,N_29430,N_28859);
and UO_878 (O_878,N_29139,N_29218);
and UO_879 (O_879,N_29375,N_28047);
and UO_880 (O_880,N_28676,N_28964);
nand UO_881 (O_881,N_29095,N_29495);
xnor UO_882 (O_882,N_28043,N_28412);
nor UO_883 (O_883,N_29742,N_29575);
xor UO_884 (O_884,N_28622,N_28218);
nand UO_885 (O_885,N_28626,N_29906);
nand UO_886 (O_886,N_29930,N_28169);
and UO_887 (O_887,N_29746,N_28888);
xnor UO_888 (O_888,N_28781,N_28884);
or UO_889 (O_889,N_29239,N_28718);
and UO_890 (O_890,N_28908,N_29747);
xor UO_891 (O_891,N_28607,N_28634);
nor UO_892 (O_892,N_28856,N_29953);
xor UO_893 (O_893,N_29683,N_28648);
nand UO_894 (O_894,N_28538,N_29118);
xor UO_895 (O_895,N_29178,N_28795);
nor UO_896 (O_896,N_28271,N_28544);
nor UO_897 (O_897,N_28983,N_29018);
or UO_898 (O_898,N_29704,N_28707);
and UO_899 (O_899,N_29958,N_29843);
nand UO_900 (O_900,N_28147,N_28515);
xor UO_901 (O_901,N_28576,N_29854);
nand UO_902 (O_902,N_28895,N_28174);
and UO_903 (O_903,N_29205,N_29853);
or UO_904 (O_904,N_29613,N_28387);
nand UO_905 (O_905,N_28252,N_29363);
nor UO_906 (O_906,N_28572,N_28037);
and UO_907 (O_907,N_29961,N_29487);
or UO_908 (O_908,N_29485,N_29983);
nand UO_909 (O_909,N_29473,N_29115);
xnor UO_910 (O_910,N_29647,N_28191);
nand UO_911 (O_911,N_29431,N_28083);
or UO_912 (O_912,N_29833,N_29484);
nor UO_913 (O_913,N_28845,N_29117);
nor UO_914 (O_914,N_28033,N_28480);
xnor UO_915 (O_915,N_29649,N_28269);
and UO_916 (O_916,N_29112,N_29364);
or UO_917 (O_917,N_28504,N_29015);
and UO_918 (O_918,N_29884,N_28179);
nand UO_919 (O_919,N_29216,N_29077);
nand UO_920 (O_920,N_29720,N_29584);
nand UO_921 (O_921,N_28186,N_29170);
nand UO_922 (O_922,N_29341,N_28887);
and UO_923 (O_923,N_28803,N_28524);
or UO_924 (O_924,N_29588,N_28837);
or UO_925 (O_925,N_29344,N_29813);
xor UO_926 (O_926,N_28423,N_29731);
xor UO_927 (O_927,N_28327,N_28153);
xor UO_928 (O_928,N_28850,N_28299);
xor UO_929 (O_929,N_28620,N_29741);
nand UO_930 (O_930,N_29201,N_29650);
nor UO_931 (O_931,N_28521,N_28132);
xor UO_932 (O_932,N_28245,N_28553);
and UO_933 (O_933,N_29175,N_29069);
nand UO_934 (O_934,N_28603,N_29295);
nor UO_935 (O_935,N_29582,N_29996);
and UO_936 (O_936,N_29472,N_28000);
xor UO_937 (O_937,N_28842,N_29655);
nand UO_938 (O_938,N_29265,N_29393);
or UO_939 (O_939,N_29614,N_29415);
nand UO_940 (O_940,N_28872,N_28125);
xor UO_941 (O_941,N_28401,N_28943);
xor UO_942 (O_942,N_29402,N_28497);
xnor UO_943 (O_943,N_29975,N_29825);
nor UO_944 (O_944,N_28733,N_29888);
xor UO_945 (O_945,N_28399,N_29299);
and UO_946 (O_946,N_29066,N_29381);
xor UO_947 (O_947,N_28921,N_29503);
and UO_948 (O_948,N_28843,N_28009);
xor UO_949 (O_949,N_28610,N_28358);
nor UO_950 (O_950,N_29350,N_29933);
nand UO_951 (O_951,N_28302,N_28213);
nor UO_952 (O_952,N_29816,N_29869);
or UO_953 (O_953,N_29017,N_28800);
nand UO_954 (O_954,N_28432,N_28462);
or UO_955 (O_955,N_29494,N_29960);
nor UO_956 (O_956,N_28408,N_28331);
xnor UO_957 (O_957,N_28319,N_28005);
and UO_958 (O_958,N_29536,N_29011);
xnor UO_959 (O_959,N_28256,N_29134);
or UO_960 (O_960,N_28101,N_29109);
and UO_961 (O_961,N_28647,N_29691);
or UO_962 (O_962,N_29399,N_28574);
xnor UO_963 (O_963,N_29654,N_29401);
and UO_964 (O_964,N_29883,N_28059);
xor UO_965 (O_965,N_28863,N_28176);
nor UO_966 (O_966,N_29885,N_29700);
and UO_967 (O_967,N_28764,N_28654);
and UO_968 (O_968,N_29489,N_29754);
xor UO_969 (O_969,N_29202,N_28144);
nor UO_970 (O_970,N_29152,N_29881);
and UO_971 (O_971,N_29254,N_29164);
nor UO_972 (O_972,N_29744,N_28734);
nand UO_973 (O_973,N_29071,N_29573);
nor UO_974 (O_974,N_29685,N_28168);
nor UO_975 (O_975,N_28373,N_29237);
nor UO_976 (O_976,N_28499,N_29748);
and UO_977 (O_977,N_29677,N_28552);
nor UO_978 (O_978,N_29398,N_29159);
nand UO_979 (O_979,N_28379,N_29631);
xor UO_980 (O_980,N_29330,N_28241);
nand UO_981 (O_981,N_28429,N_28577);
nand UO_982 (O_982,N_28413,N_28833);
nand UO_983 (O_983,N_29366,N_28543);
nor UO_984 (O_984,N_29867,N_29083);
and UO_985 (O_985,N_29142,N_28534);
and UO_986 (O_986,N_29976,N_29046);
or UO_987 (O_987,N_29372,N_29371);
or UO_988 (O_988,N_28505,N_28537);
or UO_989 (O_989,N_28142,N_28836);
nand UO_990 (O_990,N_28793,N_29470);
nand UO_991 (O_991,N_28362,N_28615);
nor UO_992 (O_992,N_29368,N_29852);
and UO_993 (O_993,N_29004,N_28708);
xor UO_994 (O_994,N_28258,N_29839);
nor UO_995 (O_995,N_28106,N_28261);
xor UO_996 (O_996,N_29899,N_29925);
or UO_997 (O_997,N_29230,N_29718);
nor UO_998 (O_998,N_29583,N_29191);
and UO_999 (O_999,N_28365,N_29753);
nand UO_1000 (O_1000,N_29755,N_28047);
and UO_1001 (O_1001,N_29151,N_29365);
and UO_1002 (O_1002,N_29386,N_28907);
nand UO_1003 (O_1003,N_28330,N_28195);
nand UO_1004 (O_1004,N_28879,N_28682);
nand UO_1005 (O_1005,N_28207,N_29032);
xor UO_1006 (O_1006,N_29833,N_29008);
nand UO_1007 (O_1007,N_29310,N_28430);
or UO_1008 (O_1008,N_29436,N_28967);
nor UO_1009 (O_1009,N_29708,N_28312);
and UO_1010 (O_1010,N_28515,N_28326);
xor UO_1011 (O_1011,N_28190,N_28614);
or UO_1012 (O_1012,N_28900,N_29345);
xor UO_1013 (O_1013,N_29215,N_28471);
nor UO_1014 (O_1014,N_29312,N_29774);
or UO_1015 (O_1015,N_28987,N_29167);
nor UO_1016 (O_1016,N_28628,N_28584);
and UO_1017 (O_1017,N_29367,N_28088);
or UO_1018 (O_1018,N_29075,N_28119);
xnor UO_1019 (O_1019,N_28324,N_28609);
nor UO_1020 (O_1020,N_28759,N_29686);
nand UO_1021 (O_1021,N_29824,N_28065);
xor UO_1022 (O_1022,N_28573,N_29859);
xnor UO_1023 (O_1023,N_29197,N_28416);
nand UO_1024 (O_1024,N_29586,N_28350);
nand UO_1025 (O_1025,N_29647,N_29788);
and UO_1026 (O_1026,N_28213,N_28032);
or UO_1027 (O_1027,N_29244,N_28091);
nor UO_1028 (O_1028,N_28749,N_29122);
xor UO_1029 (O_1029,N_29291,N_29417);
nand UO_1030 (O_1030,N_29935,N_29142);
nor UO_1031 (O_1031,N_28137,N_28650);
and UO_1032 (O_1032,N_28202,N_29864);
or UO_1033 (O_1033,N_28408,N_28963);
nor UO_1034 (O_1034,N_29087,N_28264);
xnor UO_1035 (O_1035,N_29438,N_28273);
nor UO_1036 (O_1036,N_28989,N_28385);
xnor UO_1037 (O_1037,N_29624,N_29013);
xor UO_1038 (O_1038,N_29630,N_28791);
nand UO_1039 (O_1039,N_28963,N_28156);
and UO_1040 (O_1040,N_28236,N_29616);
nor UO_1041 (O_1041,N_28503,N_29036);
and UO_1042 (O_1042,N_29807,N_28005);
xnor UO_1043 (O_1043,N_28242,N_28285);
and UO_1044 (O_1044,N_29669,N_29779);
nand UO_1045 (O_1045,N_28537,N_29758);
or UO_1046 (O_1046,N_29558,N_28331);
nor UO_1047 (O_1047,N_28158,N_29136);
xnor UO_1048 (O_1048,N_28422,N_29841);
xnor UO_1049 (O_1049,N_28069,N_28437);
xor UO_1050 (O_1050,N_28789,N_28237);
and UO_1051 (O_1051,N_28829,N_29899);
and UO_1052 (O_1052,N_28305,N_28585);
nand UO_1053 (O_1053,N_29717,N_28190);
xor UO_1054 (O_1054,N_29894,N_29541);
or UO_1055 (O_1055,N_28696,N_28216);
nor UO_1056 (O_1056,N_28186,N_29154);
nand UO_1057 (O_1057,N_29906,N_28686);
nor UO_1058 (O_1058,N_29915,N_28031);
nor UO_1059 (O_1059,N_29489,N_29853);
nor UO_1060 (O_1060,N_28581,N_29709);
and UO_1061 (O_1061,N_28220,N_29106);
nand UO_1062 (O_1062,N_28764,N_29365);
xor UO_1063 (O_1063,N_28737,N_28740);
and UO_1064 (O_1064,N_29145,N_29663);
or UO_1065 (O_1065,N_28147,N_28391);
nor UO_1066 (O_1066,N_28806,N_29731);
xor UO_1067 (O_1067,N_29693,N_29955);
xnor UO_1068 (O_1068,N_29229,N_28255);
nand UO_1069 (O_1069,N_28752,N_28398);
or UO_1070 (O_1070,N_28726,N_29925);
or UO_1071 (O_1071,N_28658,N_29306);
nor UO_1072 (O_1072,N_29910,N_28834);
or UO_1073 (O_1073,N_29392,N_28105);
and UO_1074 (O_1074,N_28689,N_28537);
and UO_1075 (O_1075,N_29503,N_29246);
xor UO_1076 (O_1076,N_29051,N_28546);
or UO_1077 (O_1077,N_29215,N_28808);
or UO_1078 (O_1078,N_28629,N_28365);
xnor UO_1079 (O_1079,N_28698,N_28802);
and UO_1080 (O_1080,N_28659,N_29746);
nor UO_1081 (O_1081,N_29550,N_28437);
xor UO_1082 (O_1082,N_28561,N_29597);
or UO_1083 (O_1083,N_29805,N_29045);
or UO_1084 (O_1084,N_29176,N_28863);
or UO_1085 (O_1085,N_28045,N_28747);
nand UO_1086 (O_1086,N_28388,N_29451);
or UO_1087 (O_1087,N_29369,N_29026);
nand UO_1088 (O_1088,N_29681,N_29901);
nand UO_1089 (O_1089,N_29420,N_29186);
and UO_1090 (O_1090,N_28840,N_29545);
nand UO_1091 (O_1091,N_29514,N_28425);
nand UO_1092 (O_1092,N_28563,N_28680);
nor UO_1093 (O_1093,N_28868,N_28008);
nand UO_1094 (O_1094,N_29438,N_29301);
and UO_1095 (O_1095,N_29823,N_29901);
nand UO_1096 (O_1096,N_29608,N_29932);
nand UO_1097 (O_1097,N_29839,N_28301);
xnor UO_1098 (O_1098,N_29192,N_29661);
nor UO_1099 (O_1099,N_28563,N_29539);
xor UO_1100 (O_1100,N_29983,N_29759);
or UO_1101 (O_1101,N_28515,N_29958);
and UO_1102 (O_1102,N_28211,N_29956);
and UO_1103 (O_1103,N_28032,N_28630);
nor UO_1104 (O_1104,N_29840,N_29668);
and UO_1105 (O_1105,N_28083,N_28553);
or UO_1106 (O_1106,N_29873,N_28122);
xor UO_1107 (O_1107,N_29414,N_29757);
nand UO_1108 (O_1108,N_28431,N_29058);
or UO_1109 (O_1109,N_29660,N_28107);
and UO_1110 (O_1110,N_29832,N_28161);
nor UO_1111 (O_1111,N_29919,N_28206);
nand UO_1112 (O_1112,N_29915,N_28065);
nand UO_1113 (O_1113,N_28101,N_29152);
or UO_1114 (O_1114,N_28998,N_29833);
nand UO_1115 (O_1115,N_28219,N_29382);
nand UO_1116 (O_1116,N_28284,N_28378);
and UO_1117 (O_1117,N_28796,N_29556);
xnor UO_1118 (O_1118,N_28116,N_28052);
nand UO_1119 (O_1119,N_28538,N_28086);
nand UO_1120 (O_1120,N_28917,N_29672);
and UO_1121 (O_1121,N_29595,N_28628);
or UO_1122 (O_1122,N_29020,N_28063);
nor UO_1123 (O_1123,N_29363,N_29934);
nor UO_1124 (O_1124,N_28689,N_29894);
or UO_1125 (O_1125,N_28027,N_28627);
xnor UO_1126 (O_1126,N_28404,N_28107);
nor UO_1127 (O_1127,N_29367,N_28213);
or UO_1128 (O_1128,N_29437,N_29804);
and UO_1129 (O_1129,N_28073,N_28342);
and UO_1130 (O_1130,N_28318,N_28134);
xor UO_1131 (O_1131,N_28985,N_29551);
or UO_1132 (O_1132,N_28673,N_28319);
nand UO_1133 (O_1133,N_28905,N_28892);
or UO_1134 (O_1134,N_29210,N_28287);
nor UO_1135 (O_1135,N_29982,N_29420);
xor UO_1136 (O_1136,N_29647,N_29583);
nand UO_1137 (O_1137,N_29379,N_28555);
nand UO_1138 (O_1138,N_29388,N_29031);
and UO_1139 (O_1139,N_29245,N_28689);
and UO_1140 (O_1140,N_28772,N_28304);
and UO_1141 (O_1141,N_29451,N_29224);
nand UO_1142 (O_1142,N_28615,N_29855);
xor UO_1143 (O_1143,N_28207,N_28189);
nor UO_1144 (O_1144,N_29367,N_28091);
nand UO_1145 (O_1145,N_28441,N_29952);
nand UO_1146 (O_1146,N_29152,N_28555);
nor UO_1147 (O_1147,N_29990,N_29647);
nand UO_1148 (O_1148,N_29281,N_28194);
and UO_1149 (O_1149,N_28749,N_29146);
nand UO_1150 (O_1150,N_29353,N_29418);
and UO_1151 (O_1151,N_28452,N_28196);
or UO_1152 (O_1152,N_28617,N_29024);
nand UO_1153 (O_1153,N_29840,N_29240);
xor UO_1154 (O_1154,N_29053,N_28445);
nand UO_1155 (O_1155,N_28339,N_29722);
or UO_1156 (O_1156,N_28845,N_28520);
nor UO_1157 (O_1157,N_28700,N_28114);
xor UO_1158 (O_1158,N_28014,N_29430);
xnor UO_1159 (O_1159,N_28494,N_29593);
and UO_1160 (O_1160,N_28758,N_29898);
xnor UO_1161 (O_1161,N_28762,N_28342);
nand UO_1162 (O_1162,N_29662,N_29930);
or UO_1163 (O_1163,N_28287,N_29029);
nand UO_1164 (O_1164,N_29554,N_29125);
nor UO_1165 (O_1165,N_29941,N_29398);
xnor UO_1166 (O_1166,N_28775,N_28297);
and UO_1167 (O_1167,N_29142,N_29677);
nor UO_1168 (O_1168,N_29339,N_28642);
nor UO_1169 (O_1169,N_29702,N_28051);
nand UO_1170 (O_1170,N_28140,N_29695);
nand UO_1171 (O_1171,N_28724,N_28006);
nor UO_1172 (O_1172,N_29440,N_28259);
xor UO_1173 (O_1173,N_29702,N_29881);
nor UO_1174 (O_1174,N_28092,N_28113);
and UO_1175 (O_1175,N_29477,N_29336);
nand UO_1176 (O_1176,N_28759,N_29819);
nor UO_1177 (O_1177,N_28072,N_29468);
nor UO_1178 (O_1178,N_29626,N_28455);
and UO_1179 (O_1179,N_28912,N_29283);
or UO_1180 (O_1180,N_29818,N_29301);
and UO_1181 (O_1181,N_28575,N_28039);
nor UO_1182 (O_1182,N_29086,N_29351);
nor UO_1183 (O_1183,N_28774,N_29359);
or UO_1184 (O_1184,N_29303,N_28634);
and UO_1185 (O_1185,N_28004,N_29860);
xnor UO_1186 (O_1186,N_28218,N_28103);
or UO_1187 (O_1187,N_28043,N_29691);
and UO_1188 (O_1188,N_28640,N_29207);
or UO_1189 (O_1189,N_28136,N_29408);
nand UO_1190 (O_1190,N_29211,N_28062);
nand UO_1191 (O_1191,N_29189,N_28851);
xnor UO_1192 (O_1192,N_28760,N_28038);
or UO_1193 (O_1193,N_29522,N_28425);
nand UO_1194 (O_1194,N_28846,N_29006);
or UO_1195 (O_1195,N_29972,N_29081);
or UO_1196 (O_1196,N_28116,N_28366);
nand UO_1197 (O_1197,N_28764,N_29905);
nor UO_1198 (O_1198,N_29883,N_28726);
and UO_1199 (O_1199,N_29571,N_28661);
nand UO_1200 (O_1200,N_29125,N_28967);
nand UO_1201 (O_1201,N_29603,N_29771);
nor UO_1202 (O_1202,N_29459,N_28709);
or UO_1203 (O_1203,N_28757,N_28146);
and UO_1204 (O_1204,N_29185,N_28978);
xor UO_1205 (O_1205,N_28067,N_29317);
or UO_1206 (O_1206,N_29403,N_28011);
xnor UO_1207 (O_1207,N_29772,N_28407);
nand UO_1208 (O_1208,N_28607,N_28834);
and UO_1209 (O_1209,N_29770,N_29899);
and UO_1210 (O_1210,N_29702,N_29377);
xor UO_1211 (O_1211,N_29715,N_29118);
xnor UO_1212 (O_1212,N_28768,N_29564);
nor UO_1213 (O_1213,N_28583,N_28096);
or UO_1214 (O_1214,N_29311,N_29788);
or UO_1215 (O_1215,N_28201,N_29143);
or UO_1216 (O_1216,N_28285,N_29985);
and UO_1217 (O_1217,N_29659,N_28130);
xnor UO_1218 (O_1218,N_29026,N_28112);
and UO_1219 (O_1219,N_29617,N_29236);
nor UO_1220 (O_1220,N_29483,N_29259);
and UO_1221 (O_1221,N_29399,N_29204);
or UO_1222 (O_1222,N_29086,N_29392);
nand UO_1223 (O_1223,N_28112,N_28732);
or UO_1224 (O_1224,N_28317,N_29861);
and UO_1225 (O_1225,N_29530,N_29144);
xnor UO_1226 (O_1226,N_29691,N_28829);
or UO_1227 (O_1227,N_28768,N_29146);
or UO_1228 (O_1228,N_28383,N_29156);
nand UO_1229 (O_1229,N_29306,N_28098);
nor UO_1230 (O_1230,N_28190,N_29492);
and UO_1231 (O_1231,N_28522,N_29550);
xor UO_1232 (O_1232,N_28075,N_29905);
nor UO_1233 (O_1233,N_29990,N_29695);
and UO_1234 (O_1234,N_28659,N_28870);
or UO_1235 (O_1235,N_28223,N_28258);
nor UO_1236 (O_1236,N_28873,N_28463);
or UO_1237 (O_1237,N_28568,N_29050);
and UO_1238 (O_1238,N_28423,N_29358);
or UO_1239 (O_1239,N_29777,N_28658);
xor UO_1240 (O_1240,N_28994,N_29993);
or UO_1241 (O_1241,N_29499,N_29993);
xnor UO_1242 (O_1242,N_29673,N_29490);
nand UO_1243 (O_1243,N_28910,N_29000);
nor UO_1244 (O_1244,N_28265,N_28625);
or UO_1245 (O_1245,N_28968,N_28981);
nor UO_1246 (O_1246,N_29346,N_29513);
nor UO_1247 (O_1247,N_29258,N_29463);
xor UO_1248 (O_1248,N_29839,N_29474);
nor UO_1249 (O_1249,N_29306,N_29313);
nor UO_1250 (O_1250,N_29047,N_28419);
nand UO_1251 (O_1251,N_28629,N_29251);
or UO_1252 (O_1252,N_29483,N_29649);
nand UO_1253 (O_1253,N_29765,N_29176);
nand UO_1254 (O_1254,N_29074,N_29904);
or UO_1255 (O_1255,N_28817,N_28452);
nand UO_1256 (O_1256,N_28638,N_29053);
or UO_1257 (O_1257,N_29504,N_28416);
nor UO_1258 (O_1258,N_29740,N_29262);
xor UO_1259 (O_1259,N_29107,N_29945);
nor UO_1260 (O_1260,N_28603,N_29473);
xor UO_1261 (O_1261,N_29848,N_28383);
xnor UO_1262 (O_1262,N_28258,N_28314);
nor UO_1263 (O_1263,N_28315,N_29169);
and UO_1264 (O_1264,N_28833,N_29674);
nor UO_1265 (O_1265,N_28165,N_28668);
xnor UO_1266 (O_1266,N_29081,N_28939);
or UO_1267 (O_1267,N_29186,N_28717);
nand UO_1268 (O_1268,N_29221,N_29624);
nor UO_1269 (O_1269,N_29017,N_28729);
nor UO_1270 (O_1270,N_28543,N_29173);
and UO_1271 (O_1271,N_29241,N_29062);
xnor UO_1272 (O_1272,N_29051,N_29366);
nand UO_1273 (O_1273,N_29551,N_28731);
or UO_1274 (O_1274,N_28290,N_29617);
nor UO_1275 (O_1275,N_29236,N_28041);
xnor UO_1276 (O_1276,N_29443,N_28579);
nor UO_1277 (O_1277,N_28081,N_29848);
and UO_1278 (O_1278,N_28122,N_28057);
nor UO_1279 (O_1279,N_29071,N_28657);
and UO_1280 (O_1280,N_29941,N_28571);
or UO_1281 (O_1281,N_28810,N_28250);
and UO_1282 (O_1282,N_29405,N_29851);
or UO_1283 (O_1283,N_29616,N_29721);
nor UO_1284 (O_1284,N_29416,N_28871);
and UO_1285 (O_1285,N_29185,N_29509);
or UO_1286 (O_1286,N_29115,N_28590);
and UO_1287 (O_1287,N_29887,N_28866);
xnor UO_1288 (O_1288,N_28750,N_28923);
and UO_1289 (O_1289,N_28494,N_29095);
and UO_1290 (O_1290,N_29864,N_29799);
or UO_1291 (O_1291,N_29916,N_29352);
xor UO_1292 (O_1292,N_29842,N_29035);
and UO_1293 (O_1293,N_28574,N_29787);
xor UO_1294 (O_1294,N_29970,N_28999);
xor UO_1295 (O_1295,N_29683,N_29686);
or UO_1296 (O_1296,N_28545,N_28167);
and UO_1297 (O_1297,N_28805,N_28839);
xor UO_1298 (O_1298,N_29842,N_28692);
and UO_1299 (O_1299,N_28533,N_29471);
or UO_1300 (O_1300,N_28629,N_28231);
nor UO_1301 (O_1301,N_29537,N_29767);
nor UO_1302 (O_1302,N_28433,N_29583);
nand UO_1303 (O_1303,N_28730,N_29532);
or UO_1304 (O_1304,N_28058,N_29478);
nand UO_1305 (O_1305,N_29578,N_29991);
nor UO_1306 (O_1306,N_29675,N_28083);
nand UO_1307 (O_1307,N_28927,N_28604);
and UO_1308 (O_1308,N_29426,N_28417);
xor UO_1309 (O_1309,N_28639,N_28642);
xor UO_1310 (O_1310,N_28668,N_29518);
nor UO_1311 (O_1311,N_29745,N_28920);
nand UO_1312 (O_1312,N_28479,N_28992);
or UO_1313 (O_1313,N_28238,N_28227);
nand UO_1314 (O_1314,N_28201,N_28468);
xnor UO_1315 (O_1315,N_28508,N_29718);
and UO_1316 (O_1316,N_29972,N_29489);
nor UO_1317 (O_1317,N_28132,N_29452);
nor UO_1318 (O_1318,N_29880,N_28287);
nor UO_1319 (O_1319,N_29786,N_28850);
nor UO_1320 (O_1320,N_28985,N_29787);
or UO_1321 (O_1321,N_29100,N_28762);
nand UO_1322 (O_1322,N_29934,N_29471);
or UO_1323 (O_1323,N_28688,N_29825);
or UO_1324 (O_1324,N_28849,N_28211);
and UO_1325 (O_1325,N_29184,N_29618);
or UO_1326 (O_1326,N_28245,N_28594);
nand UO_1327 (O_1327,N_28904,N_28947);
nand UO_1328 (O_1328,N_28268,N_28586);
or UO_1329 (O_1329,N_28215,N_29895);
or UO_1330 (O_1330,N_28622,N_29699);
nand UO_1331 (O_1331,N_29247,N_28609);
nand UO_1332 (O_1332,N_28565,N_29902);
and UO_1333 (O_1333,N_29773,N_28665);
nand UO_1334 (O_1334,N_29963,N_28505);
or UO_1335 (O_1335,N_29572,N_28133);
nand UO_1336 (O_1336,N_28728,N_29410);
and UO_1337 (O_1337,N_29992,N_29140);
xor UO_1338 (O_1338,N_28190,N_29801);
or UO_1339 (O_1339,N_29568,N_29949);
nand UO_1340 (O_1340,N_29218,N_29832);
and UO_1341 (O_1341,N_28919,N_29823);
xnor UO_1342 (O_1342,N_29701,N_29454);
nor UO_1343 (O_1343,N_28743,N_28264);
nor UO_1344 (O_1344,N_29785,N_29050);
nand UO_1345 (O_1345,N_28696,N_29272);
nand UO_1346 (O_1346,N_29956,N_28013);
nand UO_1347 (O_1347,N_28801,N_29502);
and UO_1348 (O_1348,N_29129,N_29224);
and UO_1349 (O_1349,N_29001,N_29289);
and UO_1350 (O_1350,N_29986,N_28716);
nor UO_1351 (O_1351,N_28141,N_28652);
or UO_1352 (O_1352,N_29156,N_28255);
xnor UO_1353 (O_1353,N_28103,N_29337);
xor UO_1354 (O_1354,N_29824,N_28271);
or UO_1355 (O_1355,N_28275,N_28845);
or UO_1356 (O_1356,N_29023,N_29762);
and UO_1357 (O_1357,N_29290,N_28609);
xnor UO_1358 (O_1358,N_29647,N_28439);
nor UO_1359 (O_1359,N_28351,N_29202);
nand UO_1360 (O_1360,N_29143,N_28327);
xor UO_1361 (O_1361,N_29069,N_29770);
nor UO_1362 (O_1362,N_28594,N_28973);
xnor UO_1363 (O_1363,N_29391,N_29585);
nor UO_1364 (O_1364,N_29017,N_29384);
or UO_1365 (O_1365,N_28407,N_29156);
and UO_1366 (O_1366,N_28441,N_28990);
or UO_1367 (O_1367,N_29158,N_28590);
or UO_1368 (O_1368,N_28317,N_29644);
nor UO_1369 (O_1369,N_28227,N_29862);
nor UO_1370 (O_1370,N_29050,N_29261);
xor UO_1371 (O_1371,N_28827,N_28694);
nor UO_1372 (O_1372,N_28408,N_29381);
nor UO_1373 (O_1373,N_29704,N_29051);
nand UO_1374 (O_1374,N_29747,N_28415);
and UO_1375 (O_1375,N_29933,N_28323);
or UO_1376 (O_1376,N_29525,N_28461);
nor UO_1377 (O_1377,N_28422,N_29648);
nand UO_1378 (O_1378,N_29394,N_28651);
or UO_1379 (O_1379,N_29671,N_29993);
and UO_1380 (O_1380,N_28330,N_29278);
and UO_1381 (O_1381,N_29804,N_28719);
nor UO_1382 (O_1382,N_29086,N_29187);
nand UO_1383 (O_1383,N_28527,N_29068);
xor UO_1384 (O_1384,N_28842,N_28456);
nor UO_1385 (O_1385,N_28424,N_29824);
and UO_1386 (O_1386,N_28212,N_28867);
nor UO_1387 (O_1387,N_29176,N_28412);
and UO_1388 (O_1388,N_29255,N_28172);
xnor UO_1389 (O_1389,N_28622,N_28773);
xor UO_1390 (O_1390,N_28509,N_28932);
xor UO_1391 (O_1391,N_28477,N_29913);
or UO_1392 (O_1392,N_29863,N_29712);
and UO_1393 (O_1393,N_29694,N_29185);
xor UO_1394 (O_1394,N_29787,N_28444);
and UO_1395 (O_1395,N_28115,N_28183);
xnor UO_1396 (O_1396,N_29055,N_28945);
nand UO_1397 (O_1397,N_29054,N_28208);
nor UO_1398 (O_1398,N_29695,N_29739);
nand UO_1399 (O_1399,N_29585,N_29135);
nor UO_1400 (O_1400,N_29276,N_28447);
nand UO_1401 (O_1401,N_29007,N_28088);
nand UO_1402 (O_1402,N_29040,N_29246);
nor UO_1403 (O_1403,N_29411,N_29661);
or UO_1404 (O_1404,N_29060,N_28102);
nor UO_1405 (O_1405,N_29717,N_29113);
or UO_1406 (O_1406,N_29055,N_29443);
or UO_1407 (O_1407,N_29611,N_28258);
or UO_1408 (O_1408,N_29873,N_28998);
or UO_1409 (O_1409,N_29453,N_28295);
nor UO_1410 (O_1410,N_28257,N_29617);
nor UO_1411 (O_1411,N_28733,N_28465);
or UO_1412 (O_1412,N_29212,N_28894);
nand UO_1413 (O_1413,N_29787,N_28996);
or UO_1414 (O_1414,N_28682,N_28020);
nand UO_1415 (O_1415,N_28228,N_29012);
xor UO_1416 (O_1416,N_28559,N_28642);
or UO_1417 (O_1417,N_28246,N_29091);
nand UO_1418 (O_1418,N_28213,N_29922);
nor UO_1419 (O_1419,N_29036,N_29845);
and UO_1420 (O_1420,N_28656,N_28189);
nand UO_1421 (O_1421,N_29998,N_28681);
and UO_1422 (O_1422,N_29308,N_29017);
and UO_1423 (O_1423,N_29501,N_28122);
nor UO_1424 (O_1424,N_29621,N_29513);
and UO_1425 (O_1425,N_29448,N_28499);
nand UO_1426 (O_1426,N_28666,N_28870);
or UO_1427 (O_1427,N_29430,N_28824);
or UO_1428 (O_1428,N_29009,N_28715);
nand UO_1429 (O_1429,N_29191,N_29375);
and UO_1430 (O_1430,N_28549,N_29630);
xnor UO_1431 (O_1431,N_28316,N_29644);
nand UO_1432 (O_1432,N_29189,N_28683);
xnor UO_1433 (O_1433,N_28226,N_28056);
nand UO_1434 (O_1434,N_28930,N_29465);
or UO_1435 (O_1435,N_28415,N_29608);
nand UO_1436 (O_1436,N_29577,N_28151);
xnor UO_1437 (O_1437,N_29921,N_29837);
nand UO_1438 (O_1438,N_28877,N_29016);
nand UO_1439 (O_1439,N_29502,N_28682);
xor UO_1440 (O_1440,N_28370,N_29749);
xnor UO_1441 (O_1441,N_28082,N_29844);
nor UO_1442 (O_1442,N_29328,N_29537);
or UO_1443 (O_1443,N_28234,N_29968);
and UO_1444 (O_1444,N_28274,N_28106);
nor UO_1445 (O_1445,N_28895,N_28666);
or UO_1446 (O_1446,N_29763,N_29866);
or UO_1447 (O_1447,N_28139,N_28804);
nand UO_1448 (O_1448,N_28048,N_29419);
nand UO_1449 (O_1449,N_29342,N_29041);
xnor UO_1450 (O_1450,N_28005,N_28369);
xor UO_1451 (O_1451,N_29630,N_29345);
nor UO_1452 (O_1452,N_28072,N_28110);
or UO_1453 (O_1453,N_28713,N_29122);
nand UO_1454 (O_1454,N_28095,N_29285);
nor UO_1455 (O_1455,N_28285,N_28423);
and UO_1456 (O_1456,N_28029,N_29786);
xnor UO_1457 (O_1457,N_28177,N_28751);
nor UO_1458 (O_1458,N_28658,N_29866);
nor UO_1459 (O_1459,N_28632,N_29825);
or UO_1460 (O_1460,N_28312,N_29843);
or UO_1461 (O_1461,N_29924,N_28795);
nor UO_1462 (O_1462,N_29630,N_28502);
nand UO_1463 (O_1463,N_28771,N_28800);
or UO_1464 (O_1464,N_29022,N_28548);
nand UO_1465 (O_1465,N_28547,N_28554);
nor UO_1466 (O_1466,N_29835,N_28200);
or UO_1467 (O_1467,N_28562,N_29403);
or UO_1468 (O_1468,N_28420,N_29233);
nor UO_1469 (O_1469,N_29838,N_28897);
nor UO_1470 (O_1470,N_29173,N_29548);
and UO_1471 (O_1471,N_28362,N_28431);
nand UO_1472 (O_1472,N_28052,N_29912);
nand UO_1473 (O_1473,N_29447,N_28584);
xor UO_1474 (O_1474,N_29138,N_29462);
nand UO_1475 (O_1475,N_28801,N_28125);
or UO_1476 (O_1476,N_29449,N_29635);
xor UO_1477 (O_1477,N_29649,N_28017);
nor UO_1478 (O_1478,N_29500,N_28384);
nor UO_1479 (O_1479,N_28907,N_29753);
xnor UO_1480 (O_1480,N_29892,N_29957);
and UO_1481 (O_1481,N_28192,N_29782);
nand UO_1482 (O_1482,N_29943,N_29523);
nand UO_1483 (O_1483,N_29626,N_29607);
or UO_1484 (O_1484,N_28188,N_28966);
nand UO_1485 (O_1485,N_29037,N_29576);
or UO_1486 (O_1486,N_29804,N_28393);
xnor UO_1487 (O_1487,N_29051,N_29781);
nand UO_1488 (O_1488,N_28152,N_28577);
or UO_1489 (O_1489,N_29435,N_29361);
xnor UO_1490 (O_1490,N_29995,N_28373);
nand UO_1491 (O_1491,N_28814,N_28115);
nand UO_1492 (O_1492,N_28201,N_29780);
nor UO_1493 (O_1493,N_29272,N_28888);
nand UO_1494 (O_1494,N_29598,N_28079);
nor UO_1495 (O_1495,N_29419,N_28249);
nor UO_1496 (O_1496,N_29374,N_29977);
nor UO_1497 (O_1497,N_29327,N_28764);
and UO_1498 (O_1498,N_28847,N_29927);
or UO_1499 (O_1499,N_28538,N_28250);
or UO_1500 (O_1500,N_29744,N_28493);
xor UO_1501 (O_1501,N_28004,N_28212);
nor UO_1502 (O_1502,N_28576,N_28439);
and UO_1503 (O_1503,N_29465,N_29018);
nor UO_1504 (O_1504,N_29424,N_29976);
nor UO_1505 (O_1505,N_28770,N_28823);
xor UO_1506 (O_1506,N_29373,N_28080);
nand UO_1507 (O_1507,N_28382,N_29318);
xnor UO_1508 (O_1508,N_29481,N_28547);
and UO_1509 (O_1509,N_28283,N_28159);
or UO_1510 (O_1510,N_29832,N_28955);
xnor UO_1511 (O_1511,N_28394,N_28694);
and UO_1512 (O_1512,N_28548,N_28654);
xor UO_1513 (O_1513,N_28239,N_28391);
nor UO_1514 (O_1514,N_29610,N_28184);
or UO_1515 (O_1515,N_29459,N_29138);
or UO_1516 (O_1516,N_29073,N_29157);
nor UO_1517 (O_1517,N_29439,N_29973);
or UO_1518 (O_1518,N_28128,N_28175);
and UO_1519 (O_1519,N_29453,N_28374);
or UO_1520 (O_1520,N_28083,N_29529);
nor UO_1521 (O_1521,N_28766,N_29752);
xor UO_1522 (O_1522,N_29858,N_28408);
xnor UO_1523 (O_1523,N_29182,N_28446);
nand UO_1524 (O_1524,N_28582,N_29733);
or UO_1525 (O_1525,N_28797,N_28324);
and UO_1526 (O_1526,N_29595,N_28888);
or UO_1527 (O_1527,N_29127,N_29499);
xor UO_1528 (O_1528,N_28868,N_29632);
and UO_1529 (O_1529,N_29846,N_29296);
nor UO_1530 (O_1530,N_28913,N_28489);
xnor UO_1531 (O_1531,N_29759,N_28595);
or UO_1532 (O_1532,N_29946,N_29930);
or UO_1533 (O_1533,N_29088,N_29695);
xnor UO_1534 (O_1534,N_28356,N_29416);
and UO_1535 (O_1535,N_28959,N_28591);
nor UO_1536 (O_1536,N_28106,N_29578);
and UO_1537 (O_1537,N_29283,N_28745);
or UO_1538 (O_1538,N_29119,N_29643);
xnor UO_1539 (O_1539,N_29845,N_28751);
nor UO_1540 (O_1540,N_28612,N_28636);
xor UO_1541 (O_1541,N_28065,N_28637);
and UO_1542 (O_1542,N_28823,N_29444);
nor UO_1543 (O_1543,N_29423,N_28461);
nor UO_1544 (O_1544,N_28257,N_28481);
and UO_1545 (O_1545,N_28907,N_28323);
nand UO_1546 (O_1546,N_28978,N_29688);
xnor UO_1547 (O_1547,N_28592,N_29431);
or UO_1548 (O_1548,N_29795,N_29624);
nand UO_1549 (O_1549,N_28002,N_29223);
xnor UO_1550 (O_1550,N_29340,N_28898);
xor UO_1551 (O_1551,N_28366,N_28561);
nor UO_1552 (O_1552,N_29906,N_29704);
nand UO_1553 (O_1553,N_28055,N_28366);
or UO_1554 (O_1554,N_29030,N_28080);
nand UO_1555 (O_1555,N_28697,N_29135);
nand UO_1556 (O_1556,N_28079,N_29514);
and UO_1557 (O_1557,N_29789,N_29707);
nor UO_1558 (O_1558,N_28064,N_29189);
xor UO_1559 (O_1559,N_28144,N_29284);
or UO_1560 (O_1560,N_29404,N_28427);
nand UO_1561 (O_1561,N_29773,N_28962);
or UO_1562 (O_1562,N_28342,N_28606);
or UO_1563 (O_1563,N_29145,N_29584);
and UO_1564 (O_1564,N_29137,N_28923);
xnor UO_1565 (O_1565,N_29612,N_29893);
nor UO_1566 (O_1566,N_29729,N_29754);
nor UO_1567 (O_1567,N_29951,N_29819);
or UO_1568 (O_1568,N_29265,N_29845);
nand UO_1569 (O_1569,N_29699,N_29407);
xnor UO_1570 (O_1570,N_29461,N_29340);
or UO_1571 (O_1571,N_29635,N_29312);
nor UO_1572 (O_1572,N_28533,N_29753);
nor UO_1573 (O_1573,N_28814,N_28576);
or UO_1574 (O_1574,N_28215,N_29809);
and UO_1575 (O_1575,N_28887,N_28981);
xnor UO_1576 (O_1576,N_29964,N_29778);
or UO_1577 (O_1577,N_29962,N_28957);
xor UO_1578 (O_1578,N_29834,N_29961);
or UO_1579 (O_1579,N_28202,N_29515);
xnor UO_1580 (O_1580,N_28983,N_29032);
nand UO_1581 (O_1581,N_28811,N_28717);
and UO_1582 (O_1582,N_29587,N_28249);
xor UO_1583 (O_1583,N_28684,N_28134);
xor UO_1584 (O_1584,N_29091,N_28376);
xor UO_1585 (O_1585,N_28620,N_29020);
xor UO_1586 (O_1586,N_28083,N_29828);
or UO_1587 (O_1587,N_28527,N_28368);
and UO_1588 (O_1588,N_29773,N_29797);
nand UO_1589 (O_1589,N_29734,N_28661);
xor UO_1590 (O_1590,N_28615,N_29807);
and UO_1591 (O_1591,N_28336,N_28005);
and UO_1592 (O_1592,N_29526,N_28971);
and UO_1593 (O_1593,N_29794,N_29873);
nand UO_1594 (O_1594,N_28206,N_28812);
or UO_1595 (O_1595,N_29512,N_29607);
xor UO_1596 (O_1596,N_29269,N_28894);
or UO_1597 (O_1597,N_28456,N_28954);
and UO_1598 (O_1598,N_28244,N_28340);
nor UO_1599 (O_1599,N_29743,N_29270);
xnor UO_1600 (O_1600,N_28181,N_28861);
xnor UO_1601 (O_1601,N_28149,N_28485);
xor UO_1602 (O_1602,N_28297,N_28063);
nand UO_1603 (O_1603,N_28021,N_29239);
xor UO_1604 (O_1604,N_29901,N_29129);
nand UO_1605 (O_1605,N_29419,N_29817);
nand UO_1606 (O_1606,N_28169,N_28551);
xnor UO_1607 (O_1607,N_29688,N_28915);
nand UO_1608 (O_1608,N_29082,N_29411);
xor UO_1609 (O_1609,N_28169,N_29157);
nor UO_1610 (O_1610,N_29237,N_28647);
nor UO_1611 (O_1611,N_28291,N_29304);
nor UO_1612 (O_1612,N_28086,N_29630);
nor UO_1613 (O_1613,N_28129,N_28305);
and UO_1614 (O_1614,N_28729,N_29473);
xor UO_1615 (O_1615,N_28436,N_29359);
nor UO_1616 (O_1616,N_28512,N_29509);
xor UO_1617 (O_1617,N_28525,N_28327);
nand UO_1618 (O_1618,N_29841,N_28711);
nand UO_1619 (O_1619,N_29953,N_29231);
and UO_1620 (O_1620,N_29498,N_29872);
nand UO_1621 (O_1621,N_28826,N_28780);
nor UO_1622 (O_1622,N_28652,N_29953);
or UO_1623 (O_1623,N_29933,N_29671);
and UO_1624 (O_1624,N_29186,N_29154);
or UO_1625 (O_1625,N_29398,N_28515);
or UO_1626 (O_1626,N_29878,N_29213);
and UO_1627 (O_1627,N_28891,N_29816);
or UO_1628 (O_1628,N_28083,N_28556);
xnor UO_1629 (O_1629,N_28540,N_28386);
nor UO_1630 (O_1630,N_29263,N_28042);
or UO_1631 (O_1631,N_28072,N_28095);
nand UO_1632 (O_1632,N_29326,N_29895);
and UO_1633 (O_1633,N_28932,N_28214);
or UO_1634 (O_1634,N_28992,N_29440);
xnor UO_1635 (O_1635,N_28790,N_28415);
nand UO_1636 (O_1636,N_29451,N_28654);
xor UO_1637 (O_1637,N_29298,N_29305);
nor UO_1638 (O_1638,N_29798,N_29164);
xor UO_1639 (O_1639,N_28013,N_29148);
xnor UO_1640 (O_1640,N_29243,N_28158);
nand UO_1641 (O_1641,N_28603,N_28579);
nand UO_1642 (O_1642,N_28592,N_28805);
nor UO_1643 (O_1643,N_28573,N_28938);
xor UO_1644 (O_1644,N_29331,N_28744);
xnor UO_1645 (O_1645,N_28433,N_29488);
xnor UO_1646 (O_1646,N_28207,N_28464);
nand UO_1647 (O_1647,N_28710,N_28840);
xor UO_1648 (O_1648,N_29210,N_29852);
and UO_1649 (O_1649,N_28680,N_29336);
or UO_1650 (O_1650,N_28791,N_29948);
nand UO_1651 (O_1651,N_29700,N_28481);
or UO_1652 (O_1652,N_28635,N_29586);
and UO_1653 (O_1653,N_28539,N_29687);
or UO_1654 (O_1654,N_29472,N_29297);
nand UO_1655 (O_1655,N_29752,N_29148);
nor UO_1656 (O_1656,N_29896,N_28280);
nand UO_1657 (O_1657,N_28745,N_29960);
and UO_1658 (O_1658,N_28970,N_28046);
and UO_1659 (O_1659,N_28211,N_28939);
or UO_1660 (O_1660,N_28583,N_29500);
nor UO_1661 (O_1661,N_28409,N_29608);
nand UO_1662 (O_1662,N_28053,N_28598);
nor UO_1663 (O_1663,N_29143,N_28364);
nor UO_1664 (O_1664,N_29488,N_29306);
and UO_1665 (O_1665,N_28858,N_29968);
xnor UO_1666 (O_1666,N_28871,N_29518);
nor UO_1667 (O_1667,N_29244,N_28171);
or UO_1668 (O_1668,N_29333,N_29386);
or UO_1669 (O_1669,N_28882,N_29761);
nor UO_1670 (O_1670,N_29291,N_28673);
and UO_1671 (O_1671,N_28300,N_29569);
nor UO_1672 (O_1672,N_29770,N_29051);
nor UO_1673 (O_1673,N_28186,N_28984);
or UO_1674 (O_1674,N_29917,N_28127);
nor UO_1675 (O_1675,N_29621,N_29384);
and UO_1676 (O_1676,N_29834,N_29789);
nand UO_1677 (O_1677,N_29625,N_29930);
nor UO_1678 (O_1678,N_29567,N_29134);
nand UO_1679 (O_1679,N_28604,N_29514);
or UO_1680 (O_1680,N_28171,N_29520);
or UO_1681 (O_1681,N_28339,N_28532);
nor UO_1682 (O_1682,N_29825,N_29096);
nor UO_1683 (O_1683,N_28675,N_28620);
or UO_1684 (O_1684,N_28143,N_29631);
xnor UO_1685 (O_1685,N_29119,N_29377);
xnor UO_1686 (O_1686,N_28342,N_28688);
and UO_1687 (O_1687,N_28678,N_29328);
xor UO_1688 (O_1688,N_29097,N_28052);
xnor UO_1689 (O_1689,N_28021,N_28163);
xor UO_1690 (O_1690,N_28258,N_29033);
nor UO_1691 (O_1691,N_28254,N_29669);
or UO_1692 (O_1692,N_28319,N_29877);
nand UO_1693 (O_1693,N_28342,N_29188);
xor UO_1694 (O_1694,N_29722,N_29197);
and UO_1695 (O_1695,N_28778,N_28260);
xnor UO_1696 (O_1696,N_29570,N_28389);
xnor UO_1697 (O_1697,N_29850,N_28331);
nor UO_1698 (O_1698,N_28038,N_28976);
nand UO_1699 (O_1699,N_28500,N_29506);
and UO_1700 (O_1700,N_29392,N_28801);
xnor UO_1701 (O_1701,N_28786,N_28685);
nand UO_1702 (O_1702,N_28603,N_29419);
and UO_1703 (O_1703,N_29447,N_28054);
nand UO_1704 (O_1704,N_29154,N_29706);
and UO_1705 (O_1705,N_28111,N_29652);
nor UO_1706 (O_1706,N_29125,N_28391);
or UO_1707 (O_1707,N_28995,N_28817);
nand UO_1708 (O_1708,N_29493,N_29735);
nand UO_1709 (O_1709,N_28917,N_28489);
nor UO_1710 (O_1710,N_28371,N_28623);
and UO_1711 (O_1711,N_29167,N_28161);
nand UO_1712 (O_1712,N_28083,N_28961);
nor UO_1713 (O_1713,N_29968,N_29958);
xor UO_1714 (O_1714,N_29165,N_29499);
nor UO_1715 (O_1715,N_29850,N_28510);
nand UO_1716 (O_1716,N_29185,N_29711);
or UO_1717 (O_1717,N_28676,N_29803);
nor UO_1718 (O_1718,N_29315,N_28266);
and UO_1719 (O_1719,N_29345,N_29081);
and UO_1720 (O_1720,N_29352,N_29152);
nor UO_1721 (O_1721,N_28892,N_28085);
nand UO_1722 (O_1722,N_29499,N_29176);
and UO_1723 (O_1723,N_28603,N_29485);
xor UO_1724 (O_1724,N_28283,N_29395);
xor UO_1725 (O_1725,N_29875,N_28662);
and UO_1726 (O_1726,N_28820,N_28116);
nand UO_1727 (O_1727,N_28797,N_28049);
or UO_1728 (O_1728,N_29396,N_29952);
nand UO_1729 (O_1729,N_29584,N_28086);
xor UO_1730 (O_1730,N_28943,N_29776);
or UO_1731 (O_1731,N_29467,N_29124);
or UO_1732 (O_1732,N_28593,N_29526);
nand UO_1733 (O_1733,N_29798,N_28895);
xor UO_1734 (O_1734,N_28490,N_29348);
and UO_1735 (O_1735,N_28036,N_29271);
and UO_1736 (O_1736,N_29276,N_29765);
and UO_1737 (O_1737,N_29492,N_28449);
nand UO_1738 (O_1738,N_28035,N_28432);
and UO_1739 (O_1739,N_28740,N_29917);
and UO_1740 (O_1740,N_28897,N_28377);
nor UO_1741 (O_1741,N_28794,N_29260);
or UO_1742 (O_1742,N_29074,N_29462);
nor UO_1743 (O_1743,N_29787,N_29024);
nor UO_1744 (O_1744,N_29752,N_29279);
nor UO_1745 (O_1745,N_29955,N_29312);
and UO_1746 (O_1746,N_28262,N_29589);
or UO_1747 (O_1747,N_28387,N_28986);
nor UO_1748 (O_1748,N_28945,N_29756);
xnor UO_1749 (O_1749,N_28593,N_29848);
and UO_1750 (O_1750,N_28974,N_28159);
nor UO_1751 (O_1751,N_29054,N_28311);
or UO_1752 (O_1752,N_28580,N_29825);
or UO_1753 (O_1753,N_29186,N_29441);
xnor UO_1754 (O_1754,N_28337,N_28403);
nand UO_1755 (O_1755,N_29834,N_28350);
nand UO_1756 (O_1756,N_29894,N_28993);
nor UO_1757 (O_1757,N_28467,N_28508);
or UO_1758 (O_1758,N_28682,N_29682);
or UO_1759 (O_1759,N_29878,N_29264);
xor UO_1760 (O_1760,N_29215,N_28982);
xor UO_1761 (O_1761,N_29906,N_29356);
nor UO_1762 (O_1762,N_28886,N_28619);
xnor UO_1763 (O_1763,N_28275,N_29423);
nand UO_1764 (O_1764,N_29769,N_29670);
or UO_1765 (O_1765,N_28315,N_29775);
or UO_1766 (O_1766,N_29502,N_29385);
and UO_1767 (O_1767,N_29892,N_29292);
and UO_1768 (O_1768,N_29458,N_29802);
xnor UO_1769 (O_1769,N_28899,N_28276);
nand UO_1770 (O_1770,N_29299,N_28323);
and UO_1771 (O_1771,N_28572,N_28241);
or UO_1772 (O_1772,N_28752,N_28446);
nor UO_1773 (O_1773,N_28998,N_29880);
or UO_1774 (O_1774,N_29331,N_29444);
nand UO_1775 (O_1775,N_29413,N_28008);
nand UO_1776 (O_1776,N_29778,N_28768);
nor UO_1777 (O_1777,N_29635,N_28645);
and UO_1778 (O_1778,N_28720,N_28682);
nor UO_1779 (O_1779,N_29553,N_28214);
and UO_1780 (O_1780,N_29447,N_29629);
xor UO_1781 (O_1781,N_28526,N_28505);
and UO_1782 (O_1782,N_28166,N_28050);
xor UO_1783 (O_1783,N_28634,N_29911);
nor UO_1784 (O_1784,N_29414,N_29673);
xnor UO_1785 (O_1785,N_28896,N_28188);
nor UO_1786 (O_1786,N_28997,N_28119);
nor UO_1787 (O_1787,N_28730,N_28272);
xnor UO_1788 (O_1788,N_29886,N_28802);
nand UO_1789 (O_1789,N_29977,N_29153);
nand UO_1790 (O_1790,N_29345,N_28178);
nand UO_1791 (O_1791,N_28674,N_29989);
nor UO_1792 (O_1792,N_29548,N_28413);
xor UO_1793 (O_1793,N_29739,N_28745);
nand UO_1794 (O_1794,N_29324,N_29202);
and UO_1795 (O_1795,N_29221,N_29371);
or UO_1796 (O_1796,N_28063,N_29193);
and UO_1797 (O_1797,N_28084,N_28435);
nand UO_1798 (O_1798,N_28236,N_28172);
or UO_1799 (O_1799,N_28537,N_28005);
xor UO_1800 (O_1800,N_28105,N_29863);
nand UO_1801 (O_1801,N_29791,N_28426);
nand UO_1802 (O_1802,N_29825,N_28837);
nand UO_1803 (O_1803,N_29357,N_29547);
xor UO_1804 (O_1804,N_28473,N_29954);
and UO_1805 (O_1805,N_28923,N_28341);
nand UO_1806 (O_1806,N_29320,N_29416);
or UO_1807 (O_1807,N_29183,N_28707);
nor UO_1808 (O_1808,N_28994,N_28913);
or UO_1809 (O_1809,N_28474,N_29409);
nand UO_1810 (O_1810,N_28329,N_28062);
xor UO_1811 (O_1811,N_29281,N_28999);
and UO_1812 (O_1812,N_29162,N_29300);
nor UO_1813 (O_1813,N_28193,N_29765);
nand UO_1814 (O_1814,N_29431,N_28298);
and UO_1815 (O_1815,N_28285,N_28157);
or UO_1816 (O_1816,N_29152,N_28549);
xor UO_1817 (O_1817,N_29219,N_28244);
xnor UO_1818 (O_1818,N_28302,N_28792);
or UO_1819 (O_1819,N_28299,N_29142);
nand UO_1820 (O_1820,N_28610,N_29727);
nor UO_1821 (O_1821,N_28528,N_28201);
nand UO_1822 (O_1822,N_28925,N_28890);
xor UO_1823 (O_1823,N_29465,N_28162);
or UO_1824 (O_1824,N_28227,N_29423);
nand UO_1825 (O_1825,N_29491,N_29930);
xor UO_1826 (O_1826,N_28330,N_29661);
nor UO_1827 (O_1827,N_28198,N_29236);
or UO_1828 (O_1828,N_28517,N_29159);
or UO_1829 (O_1829,N_29842,N_29593);
xor UO_1830 (O_1830,N_29206,N_28487);
and UO_1831 (O_1831,N_28179,N_29606);
nor UO_1832 (O_1832,N_29074,N_28232);
nor UO_1833 (O_1833,N_28687,N_29375);
or UO_1834 (O_1834,N_28450,N_29487);
or UO_1835 (O_1835,N_29785,N_28866);
nor UO_1836 (O_1836,N_29220,N_29641);
nand UO_1837 (O_1837,N_29414,N_28829);
xnor UO_1838 (O_1838,N_29536,N_29209);
or UO_1839 (O_1839,N_28756,N_29088);
and UO_1840 (O_1840,N_28747,N_29804);
nand UO_1841 (O_1841,N_29047,N_28710);
xor UO_1842 (O_1842,N_29917,N_28270);
nor UO_1843 (O_1843,N_28846,N_28023);
or UO_1844 (O_1844,N_29819,N_29253);
xor UO_1845 (O_1845,N_28113,N_28905);
nand UO_1846 (O_1846,N_29697,N_28670);
xnor UO_1847 (O_1847,N_29277,N_28472);
or UO_1848 (O_1848,N_29325,N_29807);
xnor UO_1849 (O_1849,N_28453,N_29422);
and UO_1850 (O_1850,N_29822,N_29266);
nor UO_1851 (O_1851,N_28374,N_29136);
or UO_1852 (O_1852,N_29299,N_29388);
and UO_1853 (O_1853,N_29226,N_29407);
nand UO_1854 (O_1854,N_28155,N_29154);
or UO_1855 (O_1855,N_29157,N_28214);
or UO_1856 (O_1856,N_28315,N_29761);
xor UO_1857 (O_1857,N_28132,N_29921);
nor UO_1858 (O_1858,N_28225,N_28267);
nor UO_1859 (O_1859,N_28650,N_28297);
nor UO_1860 (O_1860,N_28510,N_29345);
xor UO_1861 (O_1861,N_29577,N_29598);
or UO_1862 (O_1862,N_28648,N_28193);
nor UO_1863 (O_1863,N_29200,N_29314);
nor UO_1864 (O_1864,N_28655,N_28316);
and UO_1865 (O_1865,N_29406,N_29854);
or UO_1866 (O_1866,N_29346,N_29103);
nor UO_1867 (O_1867,N_28809,N_29548);
or UO_1868 (O_1868,N_29132,N_29436);
and UO_1869 (O_1869,N_28838,N_28397);
xor UO_1870 (O_1870,N_29167,N_28109);
xnor UO_1871 (O_1871,N_28959,N_29225);
and UO_1872 (O_1872,N_29056,N_29990);
nand UO_1873 (O_1873,N_29035,N_28575);
and UO_1874 (O_1874,N_28488,N_28963);
nor UO_1875 (O_1875,N_29673,N_29547);
and UO_1876 (O_1876,N_29242,N_28016);
and UO_1877 (O_1877,N_28525,N_28304);
or UO_1878 (O_1878,N_28555,N_28020);
or UO_1879 (O_1879,N_29594,N_28294);
nand UO_1880 (O_1880,N_29624,N_28222);
nand UO_1881 (O_1881,N_29213,N_29104);
and UO_1882 (O_1882,N_28660,N_29518);
and UO_1883 (O_1883,N_29501,N_29985);
nor UO_1884 (O_1884,N_29221,N_29873);
and UO_1885 (O_1885,N_28825,N_29495);
and UO_1886 (O_1886,N_29072,N_28278);
nand UO_1887 (O_1887,N_28818,N_29870);
nand UO_1888 (O_1888,N_28466,N_29580);
xnor UO_1889 (O_1889,N_28020,N_29966);
and UO_1890 (O_1890,N_29991,N_28912);
nor UO_1891 (O_1891,N_28788,N_28165);
xnor UO_1892 (O_1892,N_29455,N_28824);
and UO_1893 (O_1893,N_29231,N_28137);
or UO_1894 (O_1894,N_29224,N_28483);
and UO_1895 (O_1895,N_29727,N_29907);
nand UO_1896 (O_1896,N_28859,N_29339);
or UO_1897 (O_1897,N_28837,N_28316);
nand UO_1898 (O_1898,N_28709,N_28810);
nor UO_1899 (O_1899,N_28747,N_28099);
nor UO_1900 (O_1900,N_28965,N_29725);
or UO_1901 (O_1901,N_29139,N_28060);
nand UO_1902 (O_1902,N_28360,N_28477);
nand UO_1903 (O_1903,N_29805,N_29607);
xnor UO_1904 (O_1904,N_29725,N_28010);
nand UO_1905 (O_1905,N_28837,N_29562);
xor UO_1906 (O_1906,N_28622,N_28735);
nor UO_1907 (O_1907,N_28594,N_29537);
xor UO_1908 (O_1908,N_29495,N_29917);
nand UO_1909 (O_1909,N_28001,N_28689);
or UO_1910 (O_1910,N_29747,N_28642);
or UO_1911 (O_1911,N_28860,N_28651);
nor UO_1912 (O_1912,N_29847,N_28414);
nor UO_1913 (O_1913,N_29271,N_28810);
xnor UO_1914 (O_1914,N_29477,N_29501);
and UO_1915 (O_1915,N_28541,N_29497);
nor UO_1916 (O_1916,N_29216,N_28351);
and UO_1917 (O_1917,N_29924,N_28628);
and UO_1918 (O_1918,N_29153,N_28998);
nand UO_1919 (O_1919,N_29724,N_28002);
nor UO_1920 (O_1920,N_28318,N_28098);
nand UO_1921 (O_1921,N_28598,N_28171);
nor UO_1922 (O_1922,N_28551,N_29929);
nor UO_1923 (O_1923,N_28064,N_28704);
nand UO_1924 (O_1924,N_29099,N_29967);
and UO_1925 (O_1925,N_29418,N_28696);
nor UO_1926 (O_1926,N_29940,N_29606);
nor UO_1927 (O_1927,N_29164,N_28300);
nand UO_1928 (O_1928,N_29476,N_29693);
nor UO_1929 (O_1929,N_28519,N_28552);
nor UO_1930 (O_1930,N_28312,N_29098);
and UO_1931 (O_1931,N_28009,N_28482);
or UO_1932 (O_1932,N_29520,N_28114);
nor UO_1933 (O_1933,N_28582,N_28780);
nand UO_1934 (O_1934,N_28776,N_28784);
nor UO_1935 (O_1935,N_28461,N_29815);
nand UO_1936 (O_1936,N_29709,N_28602);
nor UO_1937 (O_1937,N_29964,N_29155);
and UO_1938 (O_1938,N_29749,N_29754);
xor UO_1939 (O_1939,N_28728,N_29580);
or UO_1940 (O_1940,N_28069,N_28287);
nand UO_1941 (O_1941,N_29443,N_29741);
nor UO_1942 (O_1942,N_29710,N_29954);
and UO_1943 (O_1943,N_29526,N_29913);
or UO_1944 (O_1944,N_29110,N_29482);
nand UO_1945 (O_1945,N_28058,N_29082);
nor UO_1946 (O_1946,N_28544,N_29838);
or UO_1947 (O_1947,N_29200,N_28973);
and UO_1948 (O_1948,N_29432,N_29710);
or UO_1949 (O_1949,N_29976,N_29924);
nand UO_1950 (O_1950,N_29307,N_29213);
xor UO_1951 (O_1951,N_28383,N_28438);
or UO_1952 (O_1952,N_29726,N_29732);
nor UO_1953 (O_1953,N_29818,N_28368);
xor UO_1954 (O_1954,N_28822,N_28196);
nor UO_1955 (O_1955,N_28142,N_28339);
and UO_1956 (O_1956,N_28126,N_28010);
nand UO_1957 (O_1957,N_29549,N_28999);
and UO_1958 (O_1958,N_29629,N_29565);
or UO_1959 (O_1959,N_29355,N_28506);
or UO_1960 (O_1960,N_28026,N_29030);
and UO_1961 (O_1961,N_29871,N_28188);
or UO_1962 (O_1962,N_29543,N_28183);
nor UO_1963 (O_1963,N_29647,N_28294);
nor UO_1964 (O_1964,N_29451,N_28288);
or UO_1965 (O_1965,N_28537,N_29448);
nor UO_1966 (O_1966,N_28043,N_29386);
nand UO_1967 (O_1967,N_29766,N_29600);
nor UO_1968 (O_1968,N_28658,N_29735);
and UO_1969 (O_1969,N_29945,N_29623);
or UO_1970 (O_1970,N_28427,N_28723);
nand UO_1971 (O_1971,N_29194,N_28057);
nand UO_1972 (O_1972,N_28638,N_28010);
xnor UO_1973 (O_1973,N_29793,N_29558);
nor UO_1974 (O_1974,N_29866,N_29103);
or UO_1975 (O_1975,N_29375,N_29386);
xnor UO_1976 (O_1976,N_28837,N_28638);
xnor UO_1977 (O_1977,N_28196,N_29765);
nor UO_1978 (O_1978,N_28215,N_29413);
xnor UO_1979 (O_1979,N_29661,N_29508);
nand UO_1980 (O_1980,N_28370,N_29331);
xor UO_1981 (O_1981,N_28915,N_29283);
or UO_1982 (O_1982,N_28155,N_29621);
or UO_1983 (O_1983,N_28813,N_29850);
and UO_1984 (O_1984,N_28137,N_29442);
nor UO_1985 (O_1985,N_28517,N_29807);
and UO_1986 (O_1986,N_28710,N_29461);
nand UO_1987 (O_1987,N_29356,N_28363);
or UO_1988 (O_1988,N_29085,N_28974);
nand UO_1989 (O_1989,N_29938,N_29511);
nor UO_1990 (O_1990,N_28594,N_29462);
nand UO_1991 (O_1991,N_29070,N_29126);
or UO_1992 (O_1992,N_28539,N_28852);
nor UO_1993 (O_1993,N_28158,N_29348);
xor UO_1994 (O_1994,N_29552,N_29687);
nor UO_1995 (O_1995,N_29923,N_29082);
xnor UO_1996 (O_1996,N_28374,N_29451);
or UO_1997 (O_1997,N_29362,N_29040);
nand UO_1998 (O_1998,N_29399,N_29665);
nand UO_1999 (O_1999,N_28908,N_28990);
or UO_2000 (O_2000,N_28537,N_29031);
nand UO_2001 (O_2001,N_29062,N_28227);
nor UO_2002 (O_2002,N_28683,N_29986);
nand UO_2003 (O_2003,N_29468,N_28770);
nor UO_2004 (O_2004,N_29688,N_29815);
nand UO_2005 (O_2005,N_29524,N_28118);
and UO_2006 (O_2006,N_28113,N_29888);
nor UO_2007 (O_2007,N_29135,N_29994);
nor UO_2008 (O_2008,N_29846,N_28429);
nor UO_2009 (O_2009,N_29144,N_28058);
or UO_2010 (O_2010,N_28348,N_28475);
and UO_2011 (O_2011,N_29241,N_29255);
and UO_2012 (O_2012,N_29325,N_28528);
or UO_2013 (O_2013,N_29202,N_28214);
xnor UO_2014 (O_2014,N_28274,N_28303);
or UO_2015 (O_2015,N_29705,N_29429);
nor UO_2016 (O_2016,N_29005,N_29809);
nand UO_2017 (O_2017,N_28467,N_29347);
and UO_2018 (O_2018,N_29009,N_29275);
or UO_2019 (O_2019,N_28187,N_28089);
nor UO_2020 (O_2020,N_29186,N_29112);
nor UO_2021 (O_2021,N_28066,N_28172);
nand UO_2022 (O_2022,N_28956,N_29075);
nor UO_2023 (O_2023,N_28292,N_29651);
or UO_2024 (O_2024,N_28166,N_28930);
nor UO_2025 (O_2025,N_29626,N_28013);
xor UO_2026 (O_2026,N_29244,N_29695);
or UO_2027 (O_2027,N_28149,N_28587);
xnor UO_2028 (O_2028,N_29417,N_29825);
nand UO_2029 (O_2029,N_29479,N_28883);
xnor UO_2030 (O_2030,N_29404,N_28092);
nand UO_2031 (O_2031,N_29100,N_28951);
nand UO_2032 (O_2032,N_28873,N_28102);
and UO_2033 (O_2033,N_29724,N_29391);
and UO_2034 (O_2034,N_29246,N_28600);
xnor UO_2035 (O_2035,N_28617,N_29076);
xnor UO_2036 (O_2036,N_28711,N_29996);
nor UO_2037 (O_2037,N_29959,N_29779);
nand UO_2038 (O_2038,N_28304,N_28219);
nor UO_2039 (O_2039,N_29679,N_29512);
and UO_2040 (O_2040,N_28524,N_28445);
and UO_2041 (O_2041,N_29878,N_29634);
and UO_2042 (O_2042,N_28823,N_29213);
nor UO_2043 (O_2043,N_29133,N_28012);
xor UO_2044 (O_2044,N_29251,N_29044);
and UO_2045 (O_2045,N_28425,N_29949);
nand UO_2046 (O_2046,N_29415,N_28479);
nor UO_2047 (O_2047,N_29472,N_28002);
nand UO_2048 (O_2048,N_29922,N_29159);
and UO_2049 (O_2049,N_29592,N_29297);
xnor UO_2050 (O_2050,N_28002,N_29897);
nor UO_2051 (O_2051,N_28259,N_28211);
nor UO_2052 (O_2052,N_29342,N_29540);
nand UO_2053 (O_2053,N_28577,N_28819);
or UO_2054 (O_2054,N_28575,N_28633);
or UO_2055 (O_2055,N_29570,N_29382);
nand UO_2056 (O_2056,N_28700,N_28132);
xor UO_2057 (O_2057,N_29329,N_29021);
nor UO_2058 (O_2058,N_28037,N_29888);
xnor UO_2059 (O_2059,N_28621,N_28067);
xor UO_2060 (O_2060,N_28779,N_28401);
nand UO_2061 (O_2061,N_28071,N_28428);
xnor UO_2062 (O_2062,N_29103,N_29345);
nor UO_2063 (O_2063,N_29220,N_29523);
nor UO_2064 (O_2064,N_29273,N_28447);
and UO_2065 (O_2065,N_28508,N_29088);
or UO_2066 (O_2066,N_28259,N_28083);
xnor UO_2067 (O_2067,N_29469,N_28971);
nor UO_2068 (O_2068,N_28032,N_28872);
nand UO_2069 (O_2069,N_28413,N_28232);
xor UO_2070 (O_2070,N_28844,N_29744);
nor UO_2071 (O_2071,N_28822,N_28694);
or UO_2072 (O_2072,N_28187,N_29034);
and UO_2073 (O_2073,N_29575,N_29309);
and UO_2074 (O_2074,N_28943,N_29068);
or UO_2075 (O_2075,N_29456,N_28129);
and UO_2076 (O_2076,N_29151,N_28498);
nand UO_2077 (O_2077,N_28200,N_29811);
or UO_2078 (O_2078,N_28185,N_28931);
xor UO_2079 (O_2079,N_29638,N_29647);
nor UO_2080 (O_2080,N_29277,N_28105);
nor UO_2081 (O_2081,N_29516,N_28877);
or UO_2082 (O_2082,N_29527,N_29513);
nand UO_2083 (O_2083,N_28967,N_28148);
nor UO_2084 (O_2084,N_29648,N_29418);
and UO_2085 (O_2085,N_28953,N_29815);
nor UO_2086 (O_2086,N_29322,N_28775);
nor UO_2087 (O_2087,N_28280,N_29114);
nor UO_2088 (O_2088,N_29438,N_29603);
or UO_2089 (O_2089,N_29845,N_29946);
nand UO_2090 (O_2090,N_29412,N_28081);
and UO_2091 (O_2091,N_29960,N_28665);
xnor UO_2092 (O_2092,N_28964,N_29635);
or UO_2093 (O_2093,N_29142,N_29891);
or UO_2094 (O_2094,N_28432,N_29231);
nand UO_2095 (O_2095,N_29300,N_29925);
and UO_2096 (O_2096,N_29822,N_28914);
xnor UO_2097 (O_2097,N_29733,N_28388);
and UO_2098 (O_2098,N_28412,N_29975);
xor UO_2099 (O_2099,N_28606,N_28849);
nand UO_2100 (O_2100,N_29697,N_28902);
nor UO_2101 (O_2101,N_29596,N_28699);
or UO_2102 (O_2102,N_28955,N_29422);
and UO_2103 (O_2103,N_29685,N_28134);
nand UO_2104 (O_2104,N_29019,N_28042);
xor UO_2105 (O_2105,N_29395,N_29106);
nor UO_2106 (O_2106,N_28549,N_29640);
or UO_2107 (O_2107,N_28218,N_28422);
or UO_2108 (O_2108,N_28524,N_29564);
nor UO_2109 (O_2109,N_28992,N_29035);
xor UO_2110 (O_2110,N_28728,N_28191);
nor UO_2111 (O_2111,N_28147,N_29736);
xnor UO_2112 (O_2112,N_29649,N_28074);
xor UO_2113 (O_2113,N_29614,N_28694);
and UO_2114 (O_2114,N_28990,N_29511);
nor UO_2115 (O_2115,N_28670,N_28962);
nor UO_2116 (O_2116,N_28694,N_29286);
xnor UO_2117 (O_2117,N_29376,N_29539);
nand UO_2118 (O_2118,N_28296,N_29737);
nor UO_2119 (O_2119,N_28441,N_28571);
nand UO_2120 (O_2120,N_29424,N_28179);
and UO_2121 (O_2121,N_28161,N_29433);
xnor UO_2122 (O_2122,N_28258,N_28912);
nor UO_2123 (O_2123,N_28497,N_29366);
xnor UO_2124 (O_2124,N_28552,N_28222);
or UO_2125 (O_2125,N_29993,N_28172);
nor UO_2126 (O_2126,N_29971,N_29037);
and UO_2127 (O_2127,N_29379,N_29719);
and UO_2128 (O_2128,N_29840,N_28613);
nand UO_2129 (O_2129,N_28531,N_28331);
or UO_2130 (O_2130,N_28016,N_29453);
nor UO_2131 (O_2131,N_28170,N_29425);
or UO_2132 (O_2132,N_29123,N_29804);
nor UO_2133 (O_2133,N_29541,N_29888);
or UO_2134 (O_2134,N_28847,N_28820);
or UO_2135 (O_2135,N_28576,N_28643);
nor UO_2136 (O_2136,N_29189,N_28040);
and UO_2137 (O_2137,N_28520,N_29779);
nand UO_2138 (O_2138,N_29601,N_29193);
or UO_2139 (O_2139,N_28057,N_28077);
nor UO_2140 (O_2140,N_29378,N_29642);
nor UO_2141 (O_2141,N_28105,N_28265);
nor UO_2142 (O_2142,N_29579,N_29610);
nor UO_2143 (O_2143,N_29444,N_29553);
nor UO_2144 (O_2144,N_29116,N_29726);
nor UO_2145 (O_2145,N_28223,N_29087);
xnor UO_2146 (O_2146,N_28235,N_29596);
and UO_2147 (O_2147,N_29044,N_28653);
and UO_2148 (O_2148,N_28387,N_28297);
xnor UO_2149 (O_2149,N_28319,N_28996);
nor UO_2150 (O_2150,N_29213,N_29221);
nor UO_2151 (O_2151,N_28799,N_29536);
and UO_2152 (O_2152,N_29730,N_29215);
nor UO_2153 (O_2153,N_29007,N_29420);
or UO_2154 (O_2154,N_29435,N_28574);
nor UO_2155 (O_2155,N_29668,N_29282);
or UO_2156 (O_2156,N_29601,N_28520);
xor UO_2157 (O_2157,N_28662,N_28949);
nor UO_2158 (O_2158,N_28476,N_28946);
xnor UO_2159 (O_2159,N_29403,N_28211);
and UO_2160 (O_2160,N_28433,N_28383);
nor UO_2161 (O_2161,N_29686,N_28450);
xor UO_2162 (O_2162,N_28586,N_29409);
xor UO_2163 (O_2163,N_28423,N_29634);
xnor UO_2164 (O_2164,N_28768,N_28042);
or UO_2165 (O_2165,N_29270,N_29925);
or UO_2166 (O_2166,N_29504,N_28177);
and UO_2167 (O_2167,N_29514,N_28564);
nand UO_2168 (O_2168,N_29897,N_29445);
and UO_2169 (O_2169,N_28910,N_29982);
nand UO_2170 (O_2170,N_29730,N_28266);
nand UO_2171 (O_2171,N_28486,N_29667);
xnor UO_2172 (O_2172,N_28287,N_29942);
or UO_2173 (O_2173,N_29773,N_28924);
and UO_2174 (O_2174,N_28603,N_28320);
or UO_2175 (O_2175,N_28142,N_29093);
nand UO_2176 (O_2176,N_29687,N_29189);
and UO_2177 (O_2177,N_28401,N_28945);
and UO_2178 (O_2178,N_29444,N_29163);
nand UO_2179 (O_2179,N_29406,N_28468);
nand UO_2180 (O_2180,N_28761,N_29244);
nand UO_2181 (O_2181,N_28118,N_28729);
and UO_2182 (O_2182,N_28985,N_29720);
or UO_2183 (O_2183,N_29494,N_28471);
xnor UO_2184 (O_2184,N_28248,N_29093);
and UO_2185 (O_2185,N_29041,N_28620);
nor UO_2186 (O_2186,N_29165,N_29592);
and UO_2187 (O_2187,N_29647,N_28405);
nand UO_2188 (O_2188,N_28490,N_28854);
xnor UO_2189 (O_2189,N_28783,N_28304);
and UO_2190 (O_2190,N_29086,N_28328);
xor UO_2191 (O_2191,N_28128,N_28589);
nand UO_2192 (O_2192,N_28614,N_28776);
xor UO_2193 (O_2193,N_28846,N_28714);
nand UO_2194 (O_2194,N_29016,N_29721);
nand UO_2195 (O_2195,N_28980,N_28662);
nand UO_2196 (O_2196,N_28445,N_29384);
xnor UO_2197 (O_2197,N_28210,N_28925);
nor UO_2198 (O_2198,N_28174,N_29699);
and UO_2199 (O_2199,N_29967,N_29087);
and UO_2200 (O_2200,N_28745,N_28939);
xnor UO_2201 (O_2201,N_29470,N_28771);
or UO_2202 (O_2202,N_29410,N_28875);
nand UO_2203 (O_2203,N_29810,N_28370);
nor UO_2204 (O_2204,N_28490,N_29479);
or UO_2205 (O_2205,N_28655,N_29200);
nand UO_2206 (O_2206,N_29777,N_29046);
xnor UO_2207 (O_2207,N_28067,N_29873);
xor UO_2208 (O_2208,N_29816,N_29252);
and UO_2209 (O_2209,N_28241,N_29470);
xor UO_2210 (O_2210,N_29674,N_29928);
or UO_2211 (O_2211,N_28893,N_28259);
nand UO_2212 (O_2212,N_29314,N_28096);
xor UO_2213 (O_2213,N_28055,N_28997);
nand UO_2214 (O_2214,N_28965,N_28821);
xnor UO_2215 (O_2215,N_29610,N_29070);
xor UO_2216 (O_2216,N_28842,N_29349);
and UO_2217 (O_2217,N_28005,N_28445);
nor UO_2218 (O_2218,N_28230,N_29176);
nor UO_2219 (O_2219,N_28908,N_29575);
and UO_2220 (O_2220,N_29033,N_29440);
xor UO_2221 (O_2221,N_28942,N_28562);
nor UO_2222 (O_2222,N_28942,N_28480);
nor UO_2223 (O_2223,N_28431,N_28457);
nor UO_2224 (O_2224,N_28718,N_28081);
nand UO_2225 (O_2225,N_28442,N_28017);
nand UO_2226 (O_2226,N_29564,N_29506);
or UO_2227 (O_2227,N_29655,N_29822);
nand UO_2228 (O_2228,N_28533,N_28529);
and UO_2229 (O_2229,N_29374,N_29334);
or UO_2230 (O_2230,N_28218,N_28567);
and UO_2231 (O_2231,N_28077,N_28959);
and UO_2232 (O_2232,N_28726,N_29366);
or UO_2233 (O_2233,N_28994,N_28466);
nor UO_2234 (O_2234,N_28223,N_28560);
and UO_2235 (O_2235,N_29756,N_29652);
or UO_2236 (O_2236,N_28579,N_29875);
xor UO_2237 (O_2237,N_28883,N_29463);
nand UO_2238 (O_2238,N_29163,N_28576);
xnor UO_2239 (O_2239,N_28347,N_29510);
and UO_2240 (O_2240,N_28451,N_29919);
nor UO_2241 (O_2241,N_28761,N_28454);
or UO_2242 (O_2242,N_29348,N_28051);
nor UO_2243 (O_2243,N_28354,N_28536);
or UO_2244 (O_2244,N_29661,N_28022);
nor UO_2245 (O_2245,N_28789,N_29744);
nand UO_2246 (O_2246,N_29559,N_29594);
and UO_2247 (O_2247,N_28970,N_29234);
nand UO_2248 (O_2248,N_29806,N_29026);
and UO_2249 (O_2249,N_28807,N_29709);
or UO_2250 (O_2250,N_29524,N_28818);
and UO_2251 (O_2251,N_29598,N_28255);
or UO_2252 (O_2252,N_29085,N_29377);
and UO_2253 (O_2253,N_28079,N_29205);
or UO_2254 (O_2254,N_28063,N_28724);
xnor UO_2255 (O_2255,N_28712,N_29182);
and UO_2256 (O_2256,N_29923,N_28930);
or UO_2257 (O_2257,N_28874,N_29634);
and UO_2258 (O_2258,N_29370,N_29243);
nand UO_2259 (O_2259,N_28452,N_28632);
and UO_2260 (O_2260,N_29463,N_29983);
nor UO_2261 (O_2261,N_29350,N_28551);
or UO_2262 (O_2262,N_28550,N_29610);
or UO_2263 (O_2263,N_28837,N_29024);
nand UO_2264 (O_2264,N_29863,N_29356);
xor UO_2265 (O_2265,N_28946,N_29608);
nand UO_2266 (O_2266,N_29175,N_28005);
and UO_2267 (O_2267,N_29124,N_28581);
or UO_2268 (O_2268,N_28505,N_29789);
nor UO_2269 (O_2269,N_29341,N_29337);
or UO_2270 (O_2270,N_29680,N_28810);
nand UO_2271 (O_2271,N_28307,N_29458);
xnor UO_2272 (O_2272,N_29837,N_29324);
and UO_2273 (O_2273,N_28680,N_29313);
nor UO_2274 (O_2274,N_29406,N_28674);
nand UO_2275 (O_2275,N_28799,N_28792);
nand UO_2276 (O_2276,N_29975,N_29218);
nor UO_2277 (O_2277,N_28148,N_28805);
or UO_2278 (O_2278,N_28235,N_29540);
or UO_2279 (O_2279,N_29178,N_29690);
nor UO_2280 (O_2280,N_29171,N_29109);
nor UO_2281 (O_2281,N_28632,N_28532);
xor UO_2282 (O_2282,N_29342,N_28637);
xnor UO_2283 (O_2283,N_28238,N_29711);
or UO_2284 (O_2284,N_29038,N_29433);
nor UO_2285 (O_2285,N_29067,N_28309);
nand UO_2286 (O_2286,N_28858,N_29754);
xnor UO_2287 (O_2287,N_28643,N_29690);
or UO_2288 (O_2288,N_28963,N_28699);
and UO_2289 (O_2289,N_28803,N_28157);
nand UO_2290 (O_2290,N_29050,N_28842);
and UO_2291 (O_2291,N_28420,N_29169);
xnor UO_2292 (O_2292,N_28182,N_29411);
xor UO_2293 (O_2293,N_29722,N_28996);
nand UO_2294 (O_2294,N_28379,N_28468);
and UO_2295 (O_2295,N_28503,N_28844);
nand UO_2296 (O_2296,N_29001,N_29362);
and UO_2297 (O_2297,N_29790,N_29906);
xnor UO_2298 (O_2298,N_29918,N_28705);
or UO_2299 (O_2299,N_28608,N_28609);
nand UO_2300 (O_2300,N_28142,N_28225);
xnor UO_2301 (O_2301,N_28645,N_28185);
nor UO_2302 (O_2302,N_28148,N_28291);
nand UO_2303 (O_2303,N_28904,N_28465);
nand UO_2304 (O_2304,N_28612,N_29452);
xor UO_2305 (O_2305,N_28867,N_28255);
and UO_2306 (O_2306,N_28328,N_29329);
nor UO_2307 (O_2307,N_29329,N_29134);
nand UO_2308 (O_2308,N_29212,N_28183);
nor UO_2309 (O_2309,N_29174,N_28145);
and UO_2310 (O_2310,N_28861,N_28089);
nor UO_2311 (O_2311,N_29167,N_28076);
and UO_2312 (O_2312,N_29730,N_28818);
xnor UO_2313 (O_2313,N_29285,N_28004);
or UO_2314 (O_2314,N_29588,N_29682);
or UO_2315 (O_2315,N_29280,N_29240);
xnor UO_2316 (O_2316,N_28596,N_29432);
or UO_2317 (O_2317,N_29050,N_28312);
nor UO_2318 (O_2318,N_29236,N_29079);
xnor UO_2319 (O_2319,N_29033,N_29306);
nand UO_2320 (O_2320,N_29149,N_29385);
nor UO_2321 (O_2321,N_28060,N_28471);
or UO_2322 (O_2322,N_28991,N_29587);
nand UO_2323 (O_2323,N_29047,N_28079);
and UO_2324 (O_2324,N_28089,N_28009);
nor UO_2325 (O_2325,N_29604,N_28149);
or UO_2326 (O_2326,N_29160,N_29953);
xor UO_2327 (O_2327,N_29203,N_29578);
or UO_2328 (O_2328,N_29349,N_29484);
nor UO_2329 (O_2329,N_29649,N_29150);
or UO_2330 (O_2330,N_29254,N_29788);
xnor UO_2331 (O_2331,N_29835,N_29668);
or UO_2332 (O_2332,N_28705,N_28698);
nand UO_2333 (O_2333,N_28627,N_29701);
nand UO_2334 (O_2334,N_29593,N_29459);
and UO_2335 (O_2335,N_29466,N_28803);
nand UO_2336 (O_2336,N_28175,N_28051);
nand UO_2337 (O_2337,N_29198,N_28885);
or UO_2338 (O_2338,N_28315,N_29566);
nor UO_2339 (O_2339,N_29953,N_29880);
or UO_2340 (O_2340,N_28102,N_28148);
nand UO_2341 (O_2341,N_28332,N_28042);
or UO_2342 (O_2342,N_28239,N_28544);
xnor UO_2343 (O_2343,N_28586,N_29427);
nand UO_2344 (O_2344,N_28385,N_29471);
and UO_2345 (O_2345,N_29389,N_28097);
nor UO_2346 (O_2346,N_28970,N_29092);
or UO_2347 (O_2347,N_29376,N_28216);
nand UO_2348 (O_2348,N_29860,N_28193);
xnor UO_2349 (O_2349,N_28524,N_29871);
nor UO_2350 (O_2350,N_29485,N_29989);
and UO_2351 (O_2351,N_29883,N_28170);
xor UO_2352 (O_2352,N_29253,N_29806);
and UO_2353 (O_2353,N_28839,N_28165);
and UO_2354 (O_2354,N_29935,N_29706);
or UO_2355 (O_2355,N_28626,N_29514);
nand UO_2356 (O_2356,N_28779,N_28447);
xnor UO_2357 (O_2357,N_28166,N_28343);
or UO_2358 (O_2358,N_28198,N_29080);
and UO_2359 (O_2359,N_28694,N_28339);
xnor UO_2360 (O_2360,N_29293,N_29740);
or UO_2361 (O_2361,N_28996,N_29453);
nand UO_2362 (O_2362,N_28907,N_28012);
and UO_2363 (O_2363,N_28113,N_29330);
and UO_2364 (O_2364,N_28036,N_29450);
or UO_2365 (O_2365,N_29900,N_29848);
nand UO_2366 (O_2366,N_29459,N_29298);
nand UO_2367 (O_2367,N_29231,N_29519);
nand UO_2368 (O_2368,N_28289,N_29122);
and UO_2369 (O_2369,N_28053,N_28429);
nor UO_2370 (O_2370,N_29358,N_28035);
or UO_2371 (O_2371,N_28627,N_28973);
nor UO_2372 (O_2372,N_28420,N_28046);
nand UO_2373 (O_2373,N_28320,N_29492);
or UO_2374 (O_2374,N_29929,N_29412);
nor UO_2375 (O_2375,N_28003,N_29128);
nand UO_2376 (O_2376,N_28298,N_28554);
and UO_2377 (O_2377,N_29992,N_28457);
or UO_2378 (O_2378,N_29067,N_29756);
and UO_2379 (O_2379,N_29178,N_29170);
nand UO_2380 (O_2380,N_29881,N_29156);
and UO_2381 (O_2381,N_29468,N_28688);
or UO_2382 (O_2382,N_29298,N_29847);
or UO_2383 (O_2383,N_29260,N_29697);
nor UO_2384 (O_2384,N_28806,N_29200);
nor UO_2385 (O_2385,N_29622,N_29565);
nor UO_2386 (O_2386,N_28455,N_28041);
nor UO_2387 (O_2387,N_29009,N_28190);
xnor UO_2388 (O_2388,N_28561,N_28938);
and UO_2389 (O_2389,N_28271,N_29367);
nor UO_2390 (O_2390,N_28966,N_28592);
xnor UO_2391 (O_2391,N_29843,N_28909);
and UO_2392 (O_2392,N_29334,N_28338);
xnor UO_2393 (O_2393,N_28124,N_28506);
nor UO_2394 (O_2394,N_29639,N_29803);
or UO_2395 (O_2395,N_29316,N_28143);
and UO_2396 (O_2396,N_28943,N_28494);
or UO_2397 (O_2397,N_28347,N_28957);
or UO_2398 (O_2398,N_28327,N_28368);
nor UO_2399 (O_2399,N_29977,N_28714);
nor UO_2400 (O_2400,N_29780,N_29282);
nor UO_2401 (O_2401,N_29279,N_28264);
and UO_2402 (O_2402,N_28818,N_29033);
nor UO_2403 (O_2403,N_28816,N_28066);
nand UO_2404 (O_2404,N_29851,N_29580);
and UO_2405 (O_2405,N_28255,N_28625);
nor UO_2406 (O_2406,N_28148,N_28764);
and UO_2407 (O_2407,N_29625,N_28364);
and UO_2408 (O_2408,N_28436,N_28953);
and UO_2409 (O_2409,N_28950,N_28602);
nor UO_2410 (O_2410,N_28657,N_29707);
nor UO_2411 (O_2411,N_28090,N_28963);
xor UO_2412 (O_2412,N_28744,N_29979);
xor UO_2413 (O_2413,N_28868,N_29545);
xnor UO_2414 (O_2414,N_29608,N_28876);
nor UO_2415 (O_2415,N_29340,N_29979);
nand UO_2416 (O_2416,N_28934,N_29492);
nand UO_2417 (O_2417,N_28273,N_28718);
nand UO_2418 (O_2418,N_29019,N_28239);
xnor UO_2419 (O_2419,N_29921,N_28887);
or UO_2420 (O_2420,N_29635,N_28070);
nor UO_2421 (O_2421,N_29839,N_29318);
or UO_2422 (O_2422,N_29406,N_28504);
nor UO_2423 (O_2423,N_28038,N_28649);
nand UO_2424 (O_2424,N_29022,N_28427);
xor UO_2425 (O_2425,N_29890,N_29961);
and UO_2426 (O_2426,N_29323,N_28918);
or UO_2427 (O_2427,N_28606,N_29186);
and UO_2428 (O_2428,N_29395,N_29812);
nand UO_2429 (O_2429,N_29965,N_29826);
and UO_2430 (O_2430,N_29890,N_29458);
nand UO_2431 (O_2431,N_29437,N_28282);
nor UO_2432 (O_2432,N_29354,N_28767);
and UO_2433 (O_2433,N_28072,N_29090);
nand UO_2434 (O_2434,N_29762,N_28160);
or UO_2435 (O_2435,N_29490,N_28814);
nor UO_2436 (O_2436,N_28385,N_28033);
and UO_2437 (O_2437,N_29753,N_28191);
and UO_2438 (O_2438,N_29559,N_29000);
or UO_2439 (O_2439,N_29433,N_29789);
and UO_2440 (O_2440,N_29003,N_29305);
nand UO_2441 (O_2441,N_28196,N_28626);
nand UO_2442 (O_2442,N_29855,N_28870);
nand UO_2443 (O_2443,N_29530,N_28014);
xnor UO_2444 (O_2444,N_28184,N_29238);
xnor UO_2445 (O_2445,N_29392,N_28660);
xnor UO_2446 (O_2446,N_29260,N_29222);
and UO_2447 (O_2447,N_28379,N_29019);
nand UO_2448 (O_2448,N_29403,N_28980);
and UO_2449 (O_2449,N_29440,N_28984);
nor UO_2450 (O_2450,N_28954,N_29835);
xor UO_2451 (O_2451,N_28954,N_29757);
nor UO_2452 (O_2452,N_29316,N_28919);
xor UO_2453 (O_2453,N_29882,N_29380);
xnor UO_2454 (O_2454,N_28797,N_28354);
nor UO_2455 (O_2455,N_29738,N_29489);
nand UO_2456 (O_2456,N_28409,N_28346);
nor UO_2457 (O_2457,N_29639,N_29754);
xor UO_2458 (O_2458,N_29076,N_29602);
xor UO_2459 (O_2459,N_28703,N_29474);
nor UO_2460 (O_2460,N_29234,N_29512);
nand UO_2461 (O_2461,N_28627,N_28711);
xor UO_2462 (O_2462,N_29818,N_28746);
nand UO_2463 (O_2463,N_28376,N_28674);
and UO_2464 (O_2464,N_28720,N_29134);
nand UO_2465 (O_2465,N_28788,N_29880);
and UO_2466 (O_2466,N_28621,N_29322);
and UO_2467 (O_2467,N_29473,N_28171);
and UO_2468 (O_2468,N_28926,N_29959);
and UO_2469 (O_2469,N_29885,N_29530);
nor UO_2470 (O_2470,N_29081,N_28175);
and UO_2471 (O_2471,N_29550,N_29850);
and UO_2472 (O_2472,N_28230,N_29023);
xor UO_2473 (O_2473,N_29143,N_28516);
nand UO_2474 (O_2474,N_28462,N_29194);
xor UO_2475 (O_2475,N_28093,N_28875);
xor UO_2476 (O_2476,N_29949,N_29538);
or UO_2477 (O_2477,N_28106,N_29430);
and UO_2478 (O_2478,N_29968,N_29625);
or UO_2479 (O_2479,N_29769,N_29279);
nor UO_2480 (O_2480,N_29182,N_29833);
xnor UO_2481 (O_2481,N_29308,N_29141);
nand UO_2482 (O_2482,N_29297,N_29067);
xor UO_2483 (O_2483,N_28644,N_28560);
nand UO_2484 (O_2484,N_29046,N_28985);
nor UO_2485 (O_2485,N_29433,N_29938);
and UO_2486 (O_2486,N_29013,N_28165);
xor UO_2487 (O_2487,N_29321,N_29495);
and UO_2488 (O_2488,N_28813,N_28037);
or UO_2489 (O_2489,N_28682,N_28768);
or UO_2490 (O_2490,N_28901,N_28412);
and UO_2491 (O_2491,N_29648,N_28714);
or UO_2492 (O_2492,N_29300,N_29671);
nor UO_2493 (O_2493,N_28127,N_29309);
nand UO_2494 (O_2494,N_28586,N_29128);
or UO_2495 (O_2495,N_29508,N_29572);
xor UO_2496 (O_2496,N_28518,N_28182);
nor UO_2497 (O_2497,N_29393,N_29729);
nand UO_2498 (O_2498,N_28542,N_28123);
nor UO_2499 (O_2499,N_28685,N_29168);
nor UO_2500 (O_2500,N_28267,N_29318);
or UO_2501 (O_2501,N_29466,N_29540);
and UO_2502 (O_2502,N_29663,N_28772);
and UO_2503 (O_2503,N_28935,N_28601);
nand UO_2504 (O_2504,N_28542,N_28282);
nor UO_2505 (O_2505,N_29817,N_29166);
and UO_2506 (O_2506,N_28798,N_28352);
and UO_2507 (O_2507,N_28330,N_28664);
nor UO_2508 (O_2508,N_28717,N_29012);
or UO_2509 (O_2509,N_28373,N_29595);
and UO_2510 (O_2510,N_28233,N_29259);
xor UO_2511 (O_2511,N_29877,N_29178);
nand UO_2512 (O_2512,N_29975,N_28717);
nand UO_2513 (O_2513,N_29277,N_29113);
nand UO_2514 (O_2514,N_29031,N_28595);
xnor UO_2515 (O_2515,N_29887,N_28140);
or UO_2516 (O_2516,N_28022,N_28288);
and UO_2517 (O_2517,N_29091,N_28588);
and UO_2518 (O_2518,N_28233,N_29346);
xor UO_2519 (O_2519,N_29114,N_29921);
or UO_2520 (O_2520,N_28545,N_28829);
and UO_2521 (O_2521,N_29260,N_29294);
nor UO_2522 (O_2522,N_28785,N_28264);
and UO_2523 (O_2523,N_28074,N_28693);
nand UO_2524 (O_2524,N_28875,N_29103);
xnor UO_2525 (O_2525,N_28839,N_29701);
and UO_2526 (O_2526,N_29161,N_28719);
xnor UO_2527 (O_2527,N_29280,N_28262);
nand UO_2528 (O_2528,N_29168,N_29945);
nand UO_2529 (O_2529,N_28628,N_29831);
and UO_2530 (O_2530,N_28601,N_29191);
xnor UO_2531 (O_2531,N_29272,N_29931);
nand UO_2532 (O_2532,N_29528,N_29655);
nand UO_2533 (O_2533,N_28958,N_29758);
and UO_2534 (O_2534,N_28576,N_29040);
and UO_2535 (O_2535,N_29552,N_28408);
nand UO_2536 (O_2536,N_28893,N_28414);
xor UO_2537 (O_2537,N_29684,N_28740);
or UO_2538 (O_2538,N_29367,N_28988);
or UO_2539 (O_2539,N_29135,N_29613);
and UO_2540 (O_2540,N_29639,N_28184);
and UO_2541 (O_2541,N_28941,N_29917);
nor UO_2542 (O_2542,N_29520,N_29090);
nand UO_2543 (O_2543,N_28783,N_28312);
and UO_2544 (O_2544,N_29415,N_28940);
nor UO_2545 (O_2545,N_28863,N_29136);
and UO_2546 (O_2546,N_28756,N_29725);
or UO_2547 (O_2547,N_28639,N_28610);
and UO_2548 (O_2548,N_28133,N_29811);
nand UO_2549 (O_2549,N_29421,N_28406);
nor UO_2550 (O_2550,N_29087,N_28093);
and UO_2551 (O_2551,N_29676,N_29125);
nand UO_2552 (O_2552,N_29364,N_28491);
nor UO_2553 (O_2553,N_29547,N_28288);
xnor UO_2554 (O_2554,N_29300,N_29301);
nor UO_2555 (O_2555,N_29210,N_29441);
nor UO_2556 (O_2556,N_29077,N_29208);
and UO_2557 (O_2557,N_29427,N_29476);
or UO_2558 (O_2558,N_29230,N_29337);
or UO_2559 (O_2559,N_28248,N_29443);
nor UO_2560 (O_2560,N_28609,N_29258);
nand UO_2561 (O_2561,N_28150,N_29429);
xor UO_2562 (O_2562,N_29609,N_29696);
or UO_2563 (O_2563,N_29211,N_28030);
nor UO_2564 (O_2564,N_28340,N_29778);
xnor UO_2565 (O_2565,N_29490,N_29098);
or UO_2566 (O_2566,N_29953,N_29087);
nor UO_2567 (O_2567,N_29497,N_28688);
nand UO_2568 (O_2568,N_29156,N_28580);
xor UO_2569 (O_2569,N_28380,N_28666);
xor UO_2570 (O_2570,N_29536,N_28861);
nor UO_2571 (O_2571,N_29027,N_29097);
xnor UO_2572 (O_2572,N_28475,N_29535);
xor UO_2573 (O_2573,N_28469,N_29575);
and UO_2574 (O_2574,N_28616,N_29365);
xnor UO_2575 (O_2575,N_29167,N_29415);
xnor UO_2576 (O_2576,N_28172,N_28063);
nand UO_2577 (O_2577,N_28452,N_29412);
or UO_2578 (O_2578,N_28414,N_29393);
nor UO_2579 (O_2579,N_28910,N_29795);
or UO_2580 (O_2580,N_29190,N_29277);
nor UO_2581 (O_2581,N_29403,N_28495);
nor UO_2582 (O_2582,N_29728,N_28487);
nor UO_2583 (O_2583,N_28243,N_28429);
nor UO_2584 (O_2584,N_28525,N_29005);
nand UO_2585 (O_2585,N_29934,N_28727);
xnor UO_2586 (O_2586,N_29639,N_29698);
nand UO_2587 (O_2587,N_29276,N_29707);
nor UO_2588 (O_2588,N_28175,N_29528);
nand UO_2589 (O_2589,N_29752,N_29436);
xnor UO_2590 (O_2590,N_28184,N_29589);
nor UO_2591 (O_2591,N_29016,N_29491);
nand UO_2592 (O_2592,N_28776,N_28674);
xor UO_2593 (O_2593,N_28072,N_28219);
nand UO_2594 (O_2594,N_29568,N_29985);
nor UO_2595 (O_2595,N_29628,N_28931);
or UO_2596 (O_2596,N_29610,N_29655);
and UO_2597 (O_2597,N_28957,N_28584);
or UO_2598 (O_2598,N_28197,N_29692);
nand UO_2599 (O_2599,N_28323,N_28379);
and UO_2600 (O_2600,N_28830,N_28652);
and UO_2601 (O_2601,N_28712,N_29445);
or UO_2602 (O_2602,N_28689,N_28412);
or UO_2603 (O_2603,N_28182,N_29281);
nor UO_2604 (O_2604,N_28648,N_29409);
nor UO_2605 (O_2605,N_28874,N_29488);
or UO_2606 (O_2606,N_28360,N_29204);
nor UO_2607 (O_2607,N_28927,N_29960);
nand UO_2608 (O_2608,N_28701,N_28419);
nor UO_2609 (O_2609,N_29099,N_28863);
and UO_2610 (O_2610,N_28625,N_29707);
or UO_2611 (O_2611,N_29053,N_28172);
and UO_2612 (O_2612,N_28680,N_28031);
nand UO_2613 (O_2613,N_29123,N_29843);
nand UO_2614 (O_2614,N_28762,N_28808);
nor UO_2615 (O_2615,N_28172,N_29181);
xnor UO_2616 (O_2616,N_28675,N_28969);
xor UO_2617 (O_2617,N_29090,N_28054);
nand UO_2618 (O_2618,N_28283,N_29305);
xnor UO_2619 (O_2619,N_28419,N_28255);
xor UO_2620 (O_2620,N_28112,N_29602);
xnor UO_2621 (O_2621,N_29391,N_28774);
or UO_2622 (O_2622,N_29494,N_29981);
or UO_2623 (O_2623,N_29919,N_29411);
or UO_2624 (O_2624,N_28829,N_28505);
nand UO_2625 (O_2625,N_29095,N_29087);
nand UO_2626 (O_2626,N_28521,N_29512);
xnor UO_2627 (O_2627,N_28440,N_28387);
xor UO_2628 (O_2628,N_28661,N_28880);
or UO_2629 (O_2629,N_28715,N_28461);
nor UO_2630 (O_2630,N_28463,N_28162);
nor UO_2631 (O_2631,N_28639,N_29605);
or UO_2632 (O_2632,N_28672,N_28887);
nor UO_2633 (O_2633,N_28672,N_28598);
xor UO_2634 (O_2634,N_28201,N_29963);
nand UO_2635 (O_2635,N_28726,N_29053);
or UO_2636 (O_2636,N_29898,N_28490);
or UO_2637 (O_2637,N_29483,N_29555);
or UO_2638 (O_2638,N_28902,N_28131);
nand UO_2639 (O_2639,N_29998,N_29821);
nor UO_2640 (O_2640,N_29011,N_29655);
nor UO_2641 (O_2641,N_29117,N_29813);
and UO_2642 (O_2642,N_28120,N_28767);
or UO_2643 (O_2643,N_29957,N_28441);
nor UO_2644 (O_2644,N_29245,N_28382);
nand UO_2645 (O_2645,N_29142,N_28068);
or UO_2646 (O_2646,N_29734,N_29882);
xnor UO_2647 (O_2647,N_29858,N_29785);
nor UO_2648 (O_2648,N_28436,N_29522);
nand UO_2649 (O_2649,N_28690,N_29194);
xnor UO_2650 (O_2650,N_29030,N_29831);
nor UO_2651 (O_2651,N_28070,N_29719);
or UO_2652 (O_2652,N_28325,N_28966);
nand UO_2653 (O_2653,N_28998,N_28678);
nor UO_2654 (O_2654,N_28763,N_29212);
nor UO_2655 (O_2655,N_28792,N_29387);
nand UO_2656 (O_2656,N_29396,N_28609);
nand UO_2657 (O_2657,N_28658,N_28474);
xor UO_2658 (O_2658,N_28059,N_29223);
nand UO_2659 (O_2659,N_29590,N_28052);
nor UO_2660 (O_2660,N_29029,N_29101);
xnor UO_2661 (O_2661,N_29814,N_28507);
xnor UO_2662 (O_2662,N_28845,N_29548);
or UO_2663 (O_2663,N_29884,N_28684);
xor UO_2664 (O_2664,N_29615,N_29846);
xor UO_2665 (O_2665,N_28248,N_28197);
and UO_2666 (O_2666,N_28047,N_29126);
xor UO_2667 (O_2667,N_29646,N_28069);
and UO_2668 (O_2668,N_29204,N_29628);
or UO_2669 (O_2669,N_28803,N_28988);
nor UO_2670 (O_2670,N_28979,N_29643);
and UO_2671 (O_2671,N_28454,N_28922);
xnor UO_2672 (O_2672,N_29110,N_28388);
and UO_2673 (O_2673,N_28615,N_29263);
nor UO_2674 (O_2674,N_28302,N_28407);
or UO_2675 (O_2675,N_29715,N_28335);
xnor UO_2676 (O_2676,N_28312,N_29290);
xnor UO_2677 (O_2677,N_29048,N_28787);
and UO_2678 (O_2678,N_28627,N_29798);
nand UO_2679 (O_2679,N_29139,N_28092);
nor UO_2680 (O_2680,N_28263,N_28824);
and UO_2681 (O_2681,N_29313,N_28577);
nor UO_2682 (O_2682,N_28089,N_28687);
or UO_2683 (O_2683,N_28680,N_29352);
and UO_2684 (O_2684,N_28516,N_29391);
or UO_2685 (O_2685,N_29326,N_28941);
or UO_2686 (O_2686,N_28760,N_29510);
nor UO_2687 (O_2687,N_28818,N_29855);
xor UO_2688 (O_2688,N_28281,N_29837);
and UO_2689 (O_2689,N_28254,N_28842);
and UO_2690 (O_2690,N_29451,N_29140);
and UO_2691 (O_2691,N_29890,N_29130);
nand UO_2692 (O_2692,N_28069,N_28389);
and UO_2693 (O_2693,N_28619,N_28407);
or UO_2694 (O_2694,N_29594,N_29467);
or UO_2695 (O_2695,N_29692,N_29032);
nor UO_2696 (O_2696,N_28078,N_29737);
nand UO_2697 (O_2697,N_28357,N_28871);
or UO_2698 (O_2698,N_28292,N_28032);
and UO_2699 (O_2699,N_28250,N_29247);
nor UO_2700 (O_2700,N_28390,N_28657);
nand UO_2701 (O_2701,N_28393,N_28534);
and UO_2702 (O_2702,N_29868,N_29271);
nor UO_2703 (O_2703,N_29315,N_28399);
and UO_2704 (O_2704,N_28446,N_29421);
xor UO_2705 (O_2705,N_29251,N_28689);
xor UO_2706 (O_2706,N_29594,N_29928);
nor UO_2707 (O_2707,N_29602,N_28749);
xnor UO_2708 (O_2708,N_28349,N_29207);
nor UO_2709 (O_2709,N_29685,N_29887);
nand UO_2710 (O_2710,N_29649,N_29155);
xor UO_2711 (O_2711,N_29503,N_28796);
and UO_2712 (O_2712,N_28080,N_29301);
nand UO_2713 (O_2713,N_29794,N_28831);
and UO_2714 (O_2714,N_29714,N_29660);
xnor UO_2715 (O_2715,N_28093,N_29722);
xor UO_2716 (O_2716,N_29307,N_29581);
nor UO_2717 (O_2717,N_28788,N_28294);
xor UO_2718 (O_2718,N_28023,N_28247);
xor UO_2719 (O_2719,N_29132,N_29995);
or UO_2720 (O_2720,N_28329,N_29139);
nor UO_2721 (O_2721,N_28132,N_28270);
nand UO_2722 (O_2722,N_28669,N_28114);
xnor UO_2723 (O_2723,N_28932,N_29955);
and UO_2724 (O_2724,N_28266,N_29857);
nor UO_2725 (O_2725,N_29117,N_29337);
xnor UO_2726 (O_2726,N_29139,N_28565);
xor UO_2727 (O_2727,N_28249,N_29153);
or UO_2728 (O_2728,N_28840,N_29748);
or UO_2729 (O_2729,N_28928,N_29853);
nand UO_2730 (O_2730,N_28191,N_28429);
or UO_2731 (O_2731,N_29913,N_28637);
or UO_2732 (O_2732,N_29898,N_29196);
nand UO_2733 (O_2733,N_28543,N_28705);
nand UO_2734 (O_2734,N_29349,N_28975);
nand UO_2735 (O_2735,N_28919,N_28677);
xnor UO_2736 (O_2736,N_29462,N_28839);
or UO_2737 (O_2737,N_29591,N_29879);
or UO_2738 (O_2738,N_28502,N_29016);
xor UO_2739 (O_2739,N_28285,N_29267);
nand UO_2740 (O_2740,N_29883,N_28608);
nor UO_2741 (O_2741,N_28614,N_29245);
xor UO_2742 (O_2742,N_28006,N_28155);
nand UO_2743 (O_2743,N_29259,N_28108);
or UO_2744 (O_2744,N_28255,N_29418);
nand UO_2745 (O_2745,N_29180,N_28654);
and UO_2746 (O_2746,N_29153,N_29615);
or UO_2747 (O_2747,N_28060,N_28051);
nand UO_2748 (O_2748,N_28757,N_29488);
or UO_2749 (O_2749,N_28261,N_29978);
or UO_2750 (O_2750,N_29265,N_29217);
nand UO_2751 (O_2751,N_29839,N_28531);
or UO_2752 (O_2752,N_28129,N_28787);
nor UO_2753 (O_2753,N_29330,N_29626);
xnor UO_2754 (O_2754,N_29629,N_28974);
and UO_2755 (O_2755,N_29537,N_29775);
or UO_2756 (O_2756,N_29092,N_29130);
xor UO_2757 (O_2757,N_28375,N_28404);
and UO_2758 (O_2758,N_29919,N_29288);
nor UO_2759 (O_2759,N_28711,N_29103);
nor UO_2760 (O_2760,N_28659,N_29692);
nor UO_2761 (O_2761,N_29592,N_29287);
nor UO_2762 (O_2762,N_28661,N_28955);
xor UO_2763 (O_2763,N_29956,N_28567);
xor UO_2764 (O_2764,N_28926,N_28124);
or UO_2765 (O_2765,N_29041,N_28911);
nand UO_2766 (O_2766,N_29584,N_29374);
nor UO_2767 (O_2767,N_28976,N_29239);
and UO_2768 (O_2768,N_28896,N_29680);
xor UO_2769 (O_2769,N_29693,N_29087);
xor UO_2770 (O_2770,N_28758,N_28481);
nor UO_2771 (O_2771,N_28879,N_29180);
nand UO_2772 (O_2772,N_28574,N_29674);
and UO_2773 (O_2773,N_29745,N_28259);
and UO_2774 (O_2774,N_28524,N_29342);
nor UO_2775 (O_2775,N_29910,N_28109);
nor UO_2776 (O_2776,N_28744,N_29558);
xnor UO_2777 (O_2777,N_29832,N_28383);
nor UO_2778 (O_2778,N_29158,N_29513);
or UO_2779 (O_2779,N_29415,N_28945);
xnor UO_2780 (O_2780,N_29335,N_29244);
xnor UO_2781 (O_2781,N_29486,N_29866);
xnor UO_2782 (O_2782,N_29663,N_29289);
nor UO_2783 (O_2783,N_29313,N_28343);
nand UO_2784 (O_2784,N_28691,N_29333);
and UO_2785 (O_2785,N_29530,N_29506);
nand UO_2786 (O_2786,N_28986,N_29631);
nor UO_2787 (O_2787,N_28881,N_28983);
nand UO_2788 (O_2788,N_29672,N_28319);
and UO_2789 (O_2789,N_28409,N_29995);
and UO_2790 (O_2790,N_28510,N_29116);
or UO_2791 (O_2791,N_28942,N_28446);
or UO_2792 (O_2792,N_28664,N_28652);
xor UO_2793 (O_2793,N_28743,N_28899);
and UO_2794 (O_2794,N_28736,N_28551);
nand UO_2795 (O_2795,N_28225,N_29031);
and UO_2796 (O_2796,N_28500,N_28272);
xnor UO_2797 (O_2797,N_28051,N_28277);
nand UO_2798 (O_2798,N_28284,N_29689);
nor UO_2799 (O_2799,N_28094,N_29918);
nand UO_2800 (O_2800,N_29017,N_29522);
nor UO_2801 (O_2801,N_29642,N_28540);
xor UO_2802 (O_2802,N_29304,N_29366);
or UO_2803 (O_2803,N_29135,N_29833);
xnor UO_2804 (O_2804,N_28106,N_29202);
nor UO_2805 (O_2805,N_28387,N_29410);
nor UO_2806 (O_2806,N_28689,N_29532);
nand UO_2807 (O_2807,N_28032,N_28097);
nand UO_2808 (O_2808,N_29757,N_29804);
nor UO_2809 (O_2809,N_29490,N_28164);
nand UO_2810 (O_2810,N_28272,N_28904);
xnor UO_2811 (O_2811,N_29793,N_29216);
nor UO_2812 (O_2812,N_29710,N_29787);
nor UO_2813 (O_2813,N_29202,N_28940);
or UO_2814 (O_2814,N_28145,N_29091);
nor UO_2815 (O_2815,N_29707,N_28389);
nor UO_2816 (O_2816,N_29952,N_29842);
and UO_2817 (O_2817,N_29763,N_28791);
or UO_2818 (O_2818,N_28945,N_28517);
nor UO_2819 (O_2819,N_29971,N_29642);
or UO_2820 (O_2820,N_29215,N_28947);
or UO_2821 (O_2821,N_29109,N_28305);
and UO_2822 (O_2822,N_28496,N_28335);
xor UO_2823 (O_2823,N_29935,N_29402);
and UO_2824 (O_2824,N_28344,N_28834);
nor UO_2825 (O_2825,N_29339,N_28403);
and UO_2826 (O_2826,N_28397,N_29790);
xnor UO_2827 (O_2827,N_29202,N_29987);
xor UO_2828 (O_2828,N_29807,N_28210);
nand UO_2829 (O_2829,N_28536,N_28324);
xor UO_2830 (O_2830,N_28292,N_28125);
nor UO_2831 (O_2831,N_28463,N_29698);
and UO_2832 (O_2832,N_29458,N_29187);
or UO_2833 (O_2833,N_29932,N_28527);
xnor UO_2834 (O_2834,N_28851,N_28391);
and UO_2835 (O_2835,N_28038,N_28802);
xnor UO_2836 (O_2836,N_29901,N_28471);
or UO_2837 (O_2837,N_29936,N_28857);
nor UO_2838 (O_2838,N_28521,N_29372);
xor UO_2839 (O_2839,N_28009,N_28325);
xor UO_2840 (O_2840,N_29348,N_29672);
and UO_2841 (O_2841,N_28187,N_29367);
or UO_2842 (O_2842,N_28845,N_28063);
nand UO_2843 (O_2843,N_28398,N_29930);
nand UO_2844 (O_2844,N_28155,N_29461);
and UO_2845 (O_2845,N_28090,N_28053);
and UO_2846 (O_2846,N_28419,N_28473);
nand UO_2847 (O_2847,N_28389,N_29231);
nand UO_2848 (O_2848,N_29397,N_28857);
or UO_2849 (O_2849,N_29255,N_28410);
and UO_2850 (O_2850,N_29416,N_29699);
nand UO_2851 (O_2851,N_28796,N_28877);
nor UO_2852 (O_2852,N_29158,N_28985);
nor UO_2853 (O_2853,N_29912,N_29709);
nand UO_2854 (O_2854,N_28639,N_29467);
nand UO_2855 (O_2855,N_28301,N_29885);
nor UO_2856 (O_2856,N_29052,N_28224);
or UO_2857 (O_2857,N_28379,N_28585);
or UO_2858 (O_2858,N_29506,N_28146);
nor UO_2859 (O_2859,N_29742,N_29619);
xnor UO_2860 (O_2860,N_29247,N_28885);
or UO_2861 (O_2861,N_29599,N_28263);
or UO_2862 (O_2862,N_29874,N_29974);
or UO_2863 (O_2863,N_29640,N_29733);
xor UO_2864 (O_2864,N_29166,N_29777);
or UO_2865 (O_2865,N_28840,N_29028);
nor UO_2866 (O_2866,N_29916,N_29783);
xor UO_2867 (O_2867,N_29247,N_28694);
and UO_2868 (O_2868,N_29273,N_28634);
or UO_2869 (O_2869,N_29167,N_29560);
nand UO_2870 (O_2870,N_28330,N_28673);
nand UO_2871 (O_2871,N_28432,N_29464);
nor UO_2872 (O_2872,N_29453,N_28259);
and UO_2873 (O_2873,N_29091,N_29280);
xnor UO_2874 (O_2874,N_28700,N_29377);
xnor UO_2875 (O_2875,N_28772,N_29424);
and UO_2876 (O_2876,N_29431,N_29073);
and UO_2877 (O_2877,N_29403,N_29456);
nor UO_2878 (O_2878,N_28933,N_29213);
nand UO_2879 (O_2879,N_29557,N_28717);
nand UO_2880 (O_2880,N_28380,N_28419);
nor UO_2881 (O_2881,N_28067,N_28110);
nor UO_2882 (O_2882,N_29088,N_29468);
and UO_2883 (O_2883,N_28085,N_29706);
or UO_2884 (O_2884,N_29143,N_28139);
or UO_2885 (O_2885,N_29170,N_29561);
xnor UO_2886 (O_2886,N_28455,N_29382);
xnor UO_2887 (O_2887,N_28152,N_29592);
or UO_2888 (O_2888,N_29096,N_28439);
nand UO_2889 (O_2889,N_29509,N_29682);
nor UO_2890 (O_2890,N_29122,N_29072);
and UO_2891 (O_2891,N_29784,N_28559);
or UO_2892 (O_2892,N_28565,N_28323);
nor UO_2893 (O_2893,N_29347,N_28621);
or UO_2894 (O_2894,N_28397,N_28888);
and UO_2895 (O_2895,N_29281,N_28631);
xor UO_2896 (O_2896,N_28358,N_28782);
or UO_2897 (O_2897,N_28213,N_28411);
nor UO_2898 (O_2898,N_28057,N_28972);
or UO_2899 (O_2899,N_29121,N_29301);
xor UO_2900 (O_2900,N_28083,N_28125);
or UO_2901 (O_2901,N_28569,N_29401);
or UO_2902 (O_2902,N_29524,N_29868);
nand UO_2903 (O_2903,N_29373,N_28796);
nand UO_2904 (O_2904,N_29042,N_28118);
nor UO_2905 (O_2905,N_29981,N_28187);
nand UO_2906 (O_2906,N_28016,N_29971);
or UO_2907 (O_2907,N_29864,N_29494);
or UO_2908 (O_2908,N_29903,N_29124);
and UO_2909 (O_2909,N_28616,N_28855);
nand UO_2910 (O_2910,N_28184,N_29315);
nand UO_2911 (O_2911,N_29933,N_29661);
or UO_2912 (O_2912,N_28668,N_29624);
xnor UO_2913 (O_2913,N_28790,N_29535);
nand UO_2914 (O_2914,N_28854,N_28284);
nor UO_2915 (O_2915,N_28253,N_29065);
xor UO_2916 (O_2916,N_29484,N_28791);
and UO_2917 (O_2917,N_29479,N_28159);
or UO_2918 (O_2918,N_28951,N_28563);
and UO_2919 (O_2919,N_29940,N_28589);
xor UO_2920 (O_2920,N_29302,N_28477);
or UO_2921 (O_2921,N_29821,N_29178);
or UO_2922 (O_2922,N_28033,N_28197);
or UO_2923 (O_2923,N_29649,N_28473);
xor UO_2924 (O_2924,N_29204,N_29474);
xor UO_2925 (O_2925,N_29321,N_28933);
nand UO_2926 (O_2926,N_29884,N_29522);
or UO_2927 (O_2927,N_28489,N_29063);
and UO_2928 (O_2928,N_28645,N_28413);
xnor UO_2929 (O_2929,N_28690,N_29761);
or UO_2930 (O_2930,N_28462,N_28096);
nand UO_2931 (O_2931,N_28759,N_29976);
or UO_2932 (O_2932,N_29900,N_29215);
nor UO_2933 (O_2933,N_28886,N_29136);
nand UO_2934 (O_2934,N_28031,N_28690);
nor UO_2935 (O_2935,N_29713,N_28142);
xor UO_2936 (O_2936,N_28643,N_29723);
and UO_2937 (O_2937,N_28841,N_28334);
nand UO_2938 (O_2938,N_28783,N_29760);
nor UO_2939 (O_2939,N_29118,N_28913);
and UO_2940 (O_2940,N_28706,N_28297);
nor UO_2941 (O_2941,N_28914,N_28152);
nor UO_2942 (O_2942,N_28997,N_28495);
xor UO_2943 (O_2943,N_28430,N_28546);
or UO_2944 (O_2944,N_28796,N_28936);
and UO_2945 (O_2945,N_29392,N_28988);
nor UO_2946 (O_2946,N_28513,N_28735);
and UO_2947 (O_2947,N_29767,N_29347);
nand UO_2948 (O_2948,N_28854,N_28468);
and UO_2949 (O_2949,N_28336,N_29479);
and UO_2950 (O_2950,N_28075,N_28599);
or UO_2951 (O_2951,N_28538,N_29840);
or UO_2952 (O_2952,N_28204,N_29210);
xor UO_2953 (O_2953,N_29725,N_29110);
nand UO_2954 (O_2954,N_29834,N_29379);
and UO_2955 (O_2955,N_28268,N_29787);
and UO_2956 (O_2956,N_28714,N_28188);
nor UO_2957 (O_2957,N_28443,N_28929);
or UO_2958 (O_2958,N_29021,N_29831);
xnor UO_2959 (O_2959,N_29478,N_29093);
and UO_2960 (O_2960,N_29058,N_28169);
nand UO_2961 (O_2961,N_28821,N_29566);
nand UO_2962 (O_2962,N_28885,N_28693);
nor UO_2963 (O_2963,N_28752,N_29841);
or UO_2964 (O_2964,N_28485,N_28701);
nand UO_2965 (O_2965,N_28072,N_28630);
xor UO_2966 (O_2966,N_28452,N_28675);
xor UO_2967 (O_2967,N_29204,N_28514);
nor UO_2968 (O_2968,N_29306,N_28687);
nand UO_2969 (O_2969,N_28200,N_28416);
xor UO_2970 (O_2970,N_28056,N_28214);
nand UO_2971 (O_2971,N_28800,N_29031);
or UO_2972 (O_2972,N_28076,N_28173);
nor UO_2973 (O_2973,N_28380,N_29829);
nand UO_2974 (O_2974,N_29629,N_28679);
nor UO_2975 (O_2975,N_29129,N_28370);
or UO_2976 (O_2976,N_29586,N_28337);
and UO_2977 (O_2977,N_29634,N_29444);
nor UO_2978 (O_2978,N_28393,N_29688);
nand UO_2979 (O_2979,N_29427,N_29160);
and UO_2980 (O_2980,N_29843,N_29312);
and UO_2981 (O_2981,N_29454,N_29231);
nor UO_2982 (O_2982,N_29314,N_28941);
nor UO_2983 (O_2983,N_28616,N_29598);
xor UO_2984 (O_2984,N_28388,N_28769);
and UO_2985 (O_2985,N_28594,N_29045);
or UO_2986 (O_2986,N_28434,N_29635);
and UO_2987 (O_2987,N_28367,N_28729);
nand UO_2988 (O_2988,N_28237,N_29318);
and UO_2989 (O_2989,N_29491,N_29923);
or UO_2990 (O_2990,N_28633,N_29359);
xor UO_2991 (O_2991,N_28306,N_29131);
xor UO_2992 (O_2992,N_28845,N_29855);
nand UO_2993 (O_2993,N_29729,N_28516);
nor UO_2994 (O_2994,N_28514,N_29995);
xor UO_2995 (O_2995,N_28181,N_28633);
nor UO_2996 (O_2996,N_29665,N_29805);
xnor UO_2997 (O_2997,N_29181,N_28729);
xnor UO_2998 (O_2998,N_29745,N_28068);
nor UO_2999 (O_2999,N_29571,N_29807);
nand UO_3000 (O_3000,N_29367,N_28059);
and UO_3001 (O_3001,N_29043,N_29350);
xor UO_3002 (O_3002,N_29444,N_28559);
nand UO_3003 (O_3003,N_28394,N_28500);
and UO_3004 (O_3004,N_29377,N_28715);
and UO_3005 (O_3005,N_29614,N_28938);
nor UO_3006 (O_3006,N_28495,N_29496);
and UO_3007 (O_3007,N_28469,N_29984);
and UO_3008 (O_3008,N_28406,N_28032);
xnor UO_3009 (O_3009,N_28717,N_28872);
nand UO_3010 (O_3010,N_29138,N_29896);
nand UO_3011 (O_3011,N_29241,N_28545);
and UO_3012 (O_3012,N_28868,N_28553);
or UO_3013 (O_3013,N_29515,N_29175);
or UO_3014 (O_3014,N_28054,N_28413);
nand UO_3015 (O_3015,N_28884,N_28858);
nor UO_3016 (O_3016,N_29065,N_28404);
xnor UO_3017 (O_3017,N_28873,N_28462);
or UO_3018 (O_3018,N_29340,N_29685);
nor UO_3019 (O_3019,N_29008,N_29759);
nor UO_3020 (O_3020,N_28495,N_28377);
or UO_3021 (O_3021,N_28853,N_29718);
nand UO_3022 (O_3022,N_29639,N_29126);
nor UO_3023 (O_3023,N_29249,N_29138);
xnor UO_3024 (O_3024,N_29066,N_29447);
and UO_3025 (O_3025,N_28441,N_29916);
nand UO_3026 (O_3026,N_29648,N_29755);
xor UO_3027 (O_3027,N_28984,N_29023);
nor UO_3028 (O_3028,N_29212,N_29432);
or UO_3029 (O_3029,N_29547,N_28601);
nand UO_3030 (O_3030,N_29582,N_29672);
and UO_3031 (O_3031,N_28815,N_29382);
nor UO_3032 (O_3032,N_28460,N_28474);
or UO_3033 (O_3033,N_28841,N_29846);
or UO_3034 (O_3034,N_29862,N_29442);
nand UO_3035 (O_3035,N_29830,N_28930);
nand UO_3036 (O_3036,N_28034,N_29549);
or UO_3037 (O_3037,N_28439,N_29986);
and UO_3038 (O_3038,N_28558,N_28980);
nand UO_3039 (O_3039,N_28365,N_29891);
nand UO_3040 (O_3040,N_28802,N_28293);
nor UO_3041 (O_3041,N_29503,N_28277);
nor UO_3042 (O_3042,N_29718,N_29592);
or UO_3043 (O_3043,N_28948,N_28499);
xor UO_3044 (O_3044,N_29710,N_29646);
nand UO_3045 (O_3045,N_28798,N_28241);
xor UO_3046 (O_3046,N_28863,N_28858);
or UO_3047 (O_3047,N_28777,N_28239);
and UO_3048 (O_3048,N_29831,N_29309);
and UO_3049 (O_3049,N_29804,N_28980);
nor UO_3050 (O_3050,N_28622,N_28997);
nor UO_3051 (O_3051,N_29309,N_28585);
or UO_3052 (O_3052,N_29650,N_28842);
nor UO_3053 (O_3053,N_28499,N_29369);
or UO_3054 (O_3054,N_29467,N_29688);
nand UO_3055 (O_3055,N_28863,N_28233);
nor UO_3056 (O_3056,N_29366,N_29145);
nand UO_3057 (O_3057,N_29981,N_29543);
xor UO_3058 (O_3058,N_28070,N_28684);
and UO_3059 (O_3059,N_28896,N_28293);
nand UO_3060 (O_3060,N_29904,N_28047);
nor UO_3061 (O_3061,N_29817,N_28236);
nor UO_3062 (O_3062,N_29690,N_29347);
or UO_3063 (O_3063,N_29112,N_28088);
nor UO_3064 (O_3064,N_29299,N_29219);
nor UO_3065 (O_3065,N_29114,N_28079);
and UO_3066 (O_3066,N_28844,N_28891);
xor UO_3067 (O_3067,N_29438,N_28065);
xor UO_3068 (O_3068,N_28290,N_28704);
and UO_3069 (O_3069,N_28935,N_29627);
xor UO_3070 (O_3070,N_28558,N_29784);
or UO_3071 (O_3071,N_29933,N_29330);
or UO_3072 (O_3072,N_29766,N_29229);
nand UO_3073 (O_3073,N_29529,N_28559);
and UO_3074 (O_3074,N_29129,N_29598);
or UO_3075 (O_3075,N_29992,N_29119);
nand UO_3076 (O_3076,N_29927,N_29859);
and UO_3077 (O_3077,N_28385,N_29264);
xnor UO_3078 (O_3078,N_28138,N_28969);
xor UO_3079 (O_3079,N_28552,N_29595);
xnor UO_3080 (O_3080,N_29732,N_28315);
xor UO_3081 (O_3081,N_28115,N_29338);
xnor UO_3082 (O_3082,N_28063,N_28651);
and UO_3083 (O_3083,N_28067,N_28238);
xor UO_3084 (O_3084,N_28221,N_29812);
nor UO_3085 (O_3085,N_28204,N_28094);
xor UO_3086 (O_3086,N_28762,N_28455);
or UO_3087 (O_3087,N_28057,N_29619);
nor UO_3088 (O_3088,N_29429,N_29807);
nor UO_3089 (O_3089,N_28209,N_28578);
nor UO_3090 (O_3090,N_29494,N_28025);
xor UO_3091 (O_3091,N_28467,N_28518);
nand UO_3092 (O_3092,N_29091,N_28716);
nor UO_3093 (O_3093,N_29277,N_28597);
nor UO_3094 (O_3094,N_29845,N_29083);
and UO_3095 (O_3095,N_29249,N_29422);
nand UO_3096 (O_3096,N_28674,N_28044);
nand UO_3097 (O_3097,N_28844,N_28205);
nand UO_3098 (O_3098,N_28501,N_28770);
or UO_3099 (O_3099,N_28691,N_29695);
and UO_3100 (O_3100,N_28714,N_28028);
nor UO_3101 (O_3101,N_28360,N_29336);
nand UO_3102 (O_3102,N_29422,N_28255);
and UO_3103 (O_3103,N_28112,N_28783);
and UO_3104 (O_3104,N_29181,N_28131);
xor UO_3105 (O_3105,N_28013,N_28023);
and UO_3106 (O_3106,N_29420,N_28921);
xnor UO_3107 (O_3107,N_28121,N_29689);
and UO_3108 (O_3108,N_29770,N_29078);
or UO_3109 (O_3109,N_29358,N_29213);
xnor UO_3110 (O_3110,N_28708,N_29784);
and UO_3111 (O_3111,N_28498,N_29605);
xor UO_3112 (O_3112,N_29476,N_28063);
or UO_3113 (O_3113,N_29701,N_28785);
xnor UO_3114 (O_3114,N_29388,N_28259);
xnor UO_3115 (O_3115,N_28616,N_29864);
nor UO_3116 (O_3116,N_28118,N_28918);
and UO_3117 (O_3117,N_28443,N_29197);
xnor UO_3118 (O_3118,N_29937,N_29463);
and UO_3119 (O_3119,N_29758,N_29962);
or UO_3120 (O_3120,N_29905,N_29826);
and UO_3121 (O_3121,N_29332,N_28538);
or UO_3122 (O_3122,N_29915,N_28676);
nand UO_3123 (O_3123,N_28204,N_28277);
or UO_3124 (O_3124,N_29262,N_28633);
nor UO_3125 (O_3125,N_29547,N_28170);
nor UO_3126 (O_3126,N_29766,N_29795);
nor UO_3127 (O_3127,N_29969,N_28575);
xnor UO_3128 (O_3128,N_29888,N_29050);
and UO_3129 (O_3129,N_29414,N_28586);
nand UO_3130 (O_3130,N_28165,N_29443);
or UO_3131 (O_3131,N_29183,N_28724);
xor UO_3132 (O_3132,N_29739,N_29182);
nand UO_3133 (O_3133,N_29829,N_28505);
xnor UO_3134 (O_3134,N_28619,N_29276);
or UO_3135 (O_3135,N_28000,N_28299);
and UO_3136 (O_3136,N_29889,N_29420);
or UO_3137 (O_3137,N_28533,N_29211);
or UO_3138 (O_3138,N_29285,N_28410);
and UO_3139 (O_3139,N_28425,N_29173);
and UO_3140 (O_3140,N_28148,N_29856);
nor UO_3141 (O_3141,N_28111,N_28415);
and UO_3142 (O_3142,N_29098,N_28864);
or UO_3143 (O_3143,N_28801,N_28976);
nand UO_3144 (O_3144,N_29079,N_29285);
xnor UO_3145 (O_3145,N_29052,N_29653);
nor UO_3146 (O_3146,N_28784,N_28219);
xor UO_3147 (O_3147,N_29062,N_28016);
xnor UO_3148 (O_3148,N_28960,N_28270);
and UO_3149 (O_3149,N_29824,N_28311);
nand UO_3150 (O_3150,N_29162,N_29192);
nor UO_3151 (O_3151,N_29137,N_28948);
and UO_3152 (O_3152,N_28529,N_29212);
xnor UO_3153 (O_3153,N_28163,N_28733);
or UO_3154 (O_3154,N_28740,N_29269);
and UO_3155 (O_3155,N_29097,N_29587);
and UO_3156 (O_3156,N_28427,N_28116);
and UO_3157 (O_3157,N_28753,N_29918);
or UO_3158 (O_3158,N_29305,N_29594);
nand UO_3159 (O_3159,N_29307,N_28857);
or UO_3160 (O_3160,N_28135,N_29320);
and UO_3161 (O_3161,N_28695,N_28802);
nand UO_3162 (O_3162,N_29787,N_29174);
or UO_3163 (O_3163,N_29137,N_28027);
nand UO_3164 (O_3164,N_29523,N_29988);
xor UO_3165 (O_3165,N_29579,N_28491);
xor UO_3166 (O_3166,N_28004,N_29183);
and UO_3167 (O_3167,N_28530,N_29473);
or UO_3168 (O_3168,N_28330,N_28571);
and UO_3169 (O_3169,N_29294,N_28092);
or UO_3170 (O_3170,N_28047,N_28799);
and UO_3171 (O_3171,N_28713,N_28164);
xnor UO_3172 (O_3172,N_28845,N_29876);
nor UO_3173 (O_3173,N_29913,N_28419);
nand UO_3174 (O_3174,N_29580,N_29922);
nand UO_3175 (O_3175,N_28790,N_29297);
nand UO_3176 (O_3176,N_29756,N_28268);
and UO_3177 (O_3177,N_29474,N_29187);
nor UO_3178 (O_3178,N_28378,N_29430);
nand UO_3179 (O_3179,N_28845,N_28324);
nor UO_3180 (O_3180,N_28769,N_29303);
nand UO_3181 (O_3181,N_29166,N_28835);
nand UO_3182 (O_3182,N_29887,N_28638);
and UO_3183 (O_3183,N_29446,N_28298);
nand UO_3184 (O_3184,N_28446,N_29747);
nand UO_3185 (O_3185,N_28717,N_29866);
xor UO_3186 (O_3186,N_29460,N_28977);
nor UO_3187 (O_3187,N_29743,N_29576);
or UO_3188 (O_3188,N_28701,N_28848);
nand UO_3189 (O_3189,N_29898,N_28180);
and UO_3190 (O_3190,N_28264,N_29409);
xnor UO_3191 (O_3191,N_29667,N_28054);
nand UO_3192 (O_3192,N_28351,N_29295);
or UO_3193 (O_3193,N_29286,N_29815);
xnor UO_3194 (O_3194,N_29474,N_28319);
nand UO_3195 (O_3195,N_28943,N_29072);
and UO_3196 (O_3196,N_29533,N_29418);
xor UO_3197 (O_3197,N_29731,N_29385);
and UO_3198 (O_3198,N_28718,N_29072);
and UO_3199 (O_3199,N_28358,N_28275);
or UO_3200 (O_3200,N_28196,N_29639);
nor UO_3201 (O_3201,N_28738,N_28649);
nor UO_3202 (O_3202,N_29430,N_29886);
or UO_3203 (O_3203,N_29465,N_28636);
xor UO_3204 (O_3204,N_29934,N_28109);
and UO_3205 (O_3205,N_29795,N_29116);
nand UO_3206 (O_3206,N_28927,N_28523);
or UO_3207 (O_3207,N_29319,N_28378);
xnor UO_3208 (O_3208,N_29858,N_28628);
xor UO_3209 (O_3209,N_29149,N_29332);
nor UO_3210 (O_3210,N_28641,N_28160);
or UO_3211 (O_3211,N_28448,N_28744);
nor UO_3212 (O_3212,N_28281,N_28847);
or UO_3213 (O_3213,N_28824,N_28325);
nor UO_3214 (O_3214,N_28903,N_28426);
or UO_3215 (O_3215,N_28150,N_29407);
nor UO_3216 (O_3216,N_29609,N_28993);
nor UO_3217 (O_3217,N_28974,N_28485);
xnor UO_3218 (O_3218,N_28395,N_29784);
xor UO_3219 (O_3219,N_29939,N_28884);
nand UO_3220 (O_3220,N_29157,N_28849);
or UO_3221 (O_3221,N_28974,N_28378);
and UO_3222 (O_3222,N_28207,N_28443);
xnor UO_3223 (O_3223,N_29526,N_29183);
xor UO_3224 (O_3224,N_29880,N_28649);
and UO_3225 (O_3225,N_28626,N_28241);
and UO_3226 (O_3226,N_28007,N_28824);
or UO_3227 (O_3227,N_28406,N_28890);
nand UO_3228 (O_3228,N_29937,N_28175);
or UO_3229 (O_3229,N_29542,N_28206);
nor UO_3230 (O_3230,N_28296,N_29524);
and UO_3231 (O_3231,N_28336,N_28332);
nor UO_3232 (O_3232,N_28166,N_29448);
nand UO_3233 (O_3233,N_28018,N_29952);
or UO_3234 (O_3234,N_28344,N_29361);
xor UO_3235 (O_3235,N_28711,N_28715);
and UO_3236 (O_3236,N_28403,N_28389);
and UO_3237 (O_3237,N_29848,N_29675);
and UO_3238 (O_3238,N_28899,N_29438);
nand UO_3239 (O_3239,N_28741,N_28799);
or UO_3240 (O_3240,N_29737,N_29894);
xnor UO_3241 (O_3241,N_29396,N_28934);
and UO_3242 (O_3242,N_28813,N_28026);
nand UO_3243 (O_3243,N_28105,N_29765);
xnor UO_3244 (O_3244,N_28494,N_29938);
or UO_3245 (O_3245,N_28144,N_29820);
nand UO_3246 (O_3246,N_29520,N_28476);
nand UO_3247 (O_3247,N_29685,N_28359);
nand UO_3248 (O_3248,N_29562,N_29460);
xor UO_3249 (O_3249,N_29568,N_28390);
xor UO_3250 (O_3250,N_28914,N_28252);
and UO_3251 (O_3251,N_29194,N_28211);
or UO_3252 (O_3252,N_29817,N_29239);
and UO_3253 (O_3253,N_28334,N_29363);
nand UO_3254 (O_3254,N_29471,N_29011);
nand UO_3255 (O_3255,N_28462,N_28583);
or UO_3256 (O_3256,N_29944,N_29652);
nor UO_3257 (O_3257,N_28348,N_28368);
xor UO_3258 (O_3258,N_29063,N_29792);
nand UO_3259 (O_3259,N_28747,N_29789);
xor UO_3260 (O_3260,N_28769,N_28806);
nor UO_3261 (O_3261,N_29713,N_29461);
and UO_3262 (O_3262,N_29027,N_29977);
and UO_3263 (O_3263,N_28789,N_29728);
xor UO_3264 (O_3264,N_29537,N_29607);
and UO_3265 (O_3265,N_29412,N_29732);
nor UO_3266 (O_3266,N_29657,N_29977);
nor UO_3267 (O_3267,N_29562,N_29489);
or UO_3268 (O_3268,N_28941,N_28803);
or UO_3269 (O_3269,N_29643,N_28820);
nor UO_3270 (O_3270,N_29463,N_29388);
nor UO_3271 (O_3271,N_28035,N_28019);
or UO_3272 (O_3272,N_28262,N_29545);
and UO_3273 (O_3273,N_28059,N_28735);
nand UO_3274 (O_3274,N_28175,N_29227);
and UO_3275 (O_3275,N_29418,N_29856);
xor UO_3276 (O_3276,N_29505,N_28252);
nor UO_3277 (O_3277,N_28654,N_28008);
xnor UO_3278 (O_3278,N_28353,N_29757);
nand UO_3279 (O_3279,N_29410,N_29784);
nor UO_3280 (O_3280,N_29250,N_29439);
nor UO_3281 (O_3281,N_29318,N_29662);
nand UO_3282 (O_3282,N_28663,N_29796);
and UO_3283 (O_3283,N_29324,N_28283);
nand UO_3284 (O_3284,N_28742,N_29096);
or UO_3285 (O_3285,N_29182,N_28693);
or UO_3286 (O_3286,N_28533,N_28544);
nor UO_3287 (O_3287,N_29795,N_28477);
nand UO_3288 (O_3288,N_28777,N_28391);
nor UO_3289 (O_3289,N_28121,N_29617);
nand UO_3290 (O_3290,N_28608,N_28386);
and UO_3291 (O_3291,N_29842,N_28221);
and UO_3292 (O_3292,N_28481,N_29492);
xnor UO_3293 (O_3293,N_28686,N_28164);
and UO_3294 (O_3294,N_29687,N_28568);
nand UO_3295 (O_3295,N_28649,N_28921);
nand UO_3296 (O_3296,N_28156,N_29054);
and UO_3297 (O_3297,N_29980,N_28127);
and UO_3298 (O_3298,N_28945,N_28610);
and UO_3299 (O_3299,N_29186,N_29046);
nand UO_3300 (O_3300,N_29973,N_28684);
and UO_3301 (O_3301,N_29338,N_29402);
nor UO_3302 (O_3302,N_29519,N_29558);
xnor UO_3303 (O_3303,N_28668,N_29114);
or UO_3304 (O_3304,N_28378,N_28269);
nor UO_3305 (O_3305,N_28019,N_29987);
and UO_3306 (O_3306,N_29030,N_29123);
xnor UO_3307 (O_3307,N_29317,N_28142);
or UO_3308 (O_3308,N_29317,N_29835);
nand UO_3309 (O_3309,N_28729,N_28384);
nor UO_3310 (O_3310,N_29879,N_29203);
and UO_3311 (O_3311,N_29684,N_29798);
or UO_3312 (O_3312,N_28271,N_28333);
xnor UO_3313 (O_3313,N_28263,N_28000);
or UO_3314 (O_3314,N_29935,N_29051);
nor UO_3315 (O_3315,N_28745,N_28064);
and UO_3316 (O_3316,N_28492,N_29477);
xnor UO_3317 (O_3317,N_29889,N_29885);
nand UO_3318 (O_3318,N_29388,N_29922);
and UO_3319 (O_3319,N_28893,N_28891);
and UO_3320 (O_3320,N_29949,N_29849);
nand UO_3321 (O_3321,N_28693,N_29824);
or UO_3322 (O_3322,N_29883,N_29851);
nor UO_3323 (O_3323,N_28740,N_29818);
nor UO_3324 (O_3324,N_29901,N_28237);
nand UO_3325 (O_3325,N_29808,N_29991);
xnor UO_3326 (O_3326,N_29935,N_29635);
and UO_3327 (O_3327,N_29052,N_28057);
or UO_3328 (O_3328,N_28493,N_28982);
nand UO_3329 (O_3329,N_28683,N_29657);
or UO_3330 (O_3330,N_29022,N_29489);
nor UO_3331 (O_3331,N_28237,N_29466);
and UO_3332 (O_3332,N_28117,N_29488);
nand UO_3333 (O_3333,N_29825,N_29317);
nand UO_3334 (O_3334,N_28542,N_29515);
or UO_3335 (O_3335,N_28186,N_28823);
and UO_3336 (O_3336,N_28796,N_28314);
xor UO_3337 (O_3337,N_28246,N_29269);
or UO_3338 (O_3338,N_28073,N_29089);
nor UO_3339 (O_3339,N_28330,N_28953);
nor UO_3340 (O_3340,N_28749,N_29979);
and UO_3341 (O_3341,N_29102,N_28589);
and UO_3342 (O_3342,N_29528,N_29738);
xnor UO_3343 (O_3343,N_29148,N_28243);
or UO_3344 (O_3344,N_29888,N_29322);
nor UO_3345 (O_3345,N_29922,N_28389);
and UO_3346 (O_3346,N_29346,N_29990);
xor UO_3347 (O_3347,N_28989,N_28814);
xnor UO_3348 (O_3348,N_29567,N_28020);
nand UO_3349 (O_3349,N_29403,N_29598);
nor UO_3350 (O_3350,N_29991,N_29948);
and UO_3351 (O_3351,N_28578,N_29038);
nand UO_3352 (O_3352,N_29771,N_29039);
and UO_3353 (O_3353,N_28954,N_29147);
or UO_3354 (O_3354,N_29900,N_28359);
or UO_3355 (O_3355,N_29135,N_28263);
and UO_3356 (O_3356,N_28038,N_28576);
or UO_3357 (O_3357,N_29607,N_29612);
or UO_3358 (O_3358,N_29408,N_28447);
nor UO_3359 (O_3359,N_29153,N_28540);
nand UO_3360 (O_3360,N_28083,N_29945);
and UO_3361 (O_3361,N_29490,N_28331);
xnor UO_3362 (O_3362,N_28123,N_29926);
or UO_3363 (O_3363,N_28331,N_28228);
nor UO_3364 (O_3364,N_29688,N_28496);
xnor UO_3365 (O_3365,N_28241,N_28497);
nor UO_3366 (O_3366,N_28904,N_29453);
or UO_3367 (O_3367,N_28996,N_28864);
and UO_3368 (O_3368,N_29895,N_28332);
and UO_3369 (O_3369,N_29758,N_28383);
nor UO_3370 (O_3370,N_29554,N_28462);
and UO_3371 (O_3371,N_29862,N_29727);
xor UO_3372 (O_3372,N_28883,N_29262);
xor UO_3373 (O_3373,N_29758,N_28856);
or UO_3374 (O_3374,N_28194,N_28014);
nor UO_3375 (O_3375,N_28101,N_28326);
nor UO_3376 (O_3376,N_29818,N_29298);
xnor UO_3377 (O_3377,N_28984,N_28545);
nand UO_3378 (O_3378,N_28949,N_29735);
xor UO_3379 (O_3379,N_29017,N_29604);
and UO_3380 (O_3380,N_29519,N_28612);
nand UO_3381 (O_3381,N_28692,N_28020);
xor UO_3382 (O_3382,N_28413,N_29016);
nor UO_3383 (O_3383,N_28726,N_28304);
xor UO_3384 (O_3384,N_29250,N_29081);
nor UO_3385 (O_3385,N_28524,N_29750);
nor UO_3386 (O_3386,N_28216,N_28368);
nor UO_3387 (O_3387,N_28093,N_29733);
or UO_3388 (O_3388,N_28879,N_28381);
or UO_3389 (O_3389,N_28079,N_29966);
xor UO_3390 (O_3390,N_28936,N_29491);
or UO_3391 (O_3391,N_29268,N_29333);
nand UO_3392 (O_3392,N_28781,N_28146);
and UO_3393 (O_3393,N_29524,N_28977);
or UO_3394 (O_3394,N_28414,N_28344);
or UO_3395 (O_3395,N_28172,N_28407);
and UO_3396 (O_3396,N_29551,N_29039);
nand UO_3397 (O_3397,N_28989,N_28944);
nor UO_3398 (O_3398,N_29165,N_29942);
nor UO_3399 (O_3399,N_29107,N_28285);
nor UO_3400 (O_3400,N_28360,N_28739);
or UO_3401 (O_3401,N_28416,N_29002);
and UO_3402 (O_3402,N_28821,N_29339);
nor UO_3403 (O_3403,N_28861,N_29058);
and UO_3404 (O_3404,N_29645,N_29797);
xor UO_3405 (O_3405,N_28558,N_28534);
xor UO_3406 (O_3406,N_28145,N_29541);
nand UO_3407 (O_3407,N_28012,N_28064);
xnor UO_3408 (O_3408,N_28370,N_28849);
xnor UO_3409 (O_3409,N_29130,N_29247);
nor UO_3410 (O_3410,N_28607,N_29784);
xor UO_3411 (O_3411,N_28779,N_28455);
nor UO_3412 (O_3412,N_28201,N_29176);
and UO_3413 (O_3413,N_28665,N_29411);
nand UO_3414 (O_3414,N_29232,N_29861);
or UO_3415 (O_3415,N_29196,N_29140);
or UO_3416 (O_3416,N_29579,N_29166);
xor UO_3417 (O_3417,N_28071,N_29976);
nand UO_3418 (O_3418,N_29073,N_28459);
and UO_3419 (O_3419,N_29599,N_29404);
nand UO_3420 (O_3420,N_28892,N_28322);
xor UO_3421 (O_3421,N_28726,N_28623);
nand UO_3422 (O_3422,N_29166,N_28467);
nor UO_3423 (O_3423,N_29028,N_29069);
and UO_3424 (O_3424,N_28822,N_28767);
xnor UO_3425 (O_3425,N_29648,N_28830);
nor UO_3426 (O_3426,N_28689,N_29812);
or UO_3427 (O_3427,N_29967,N_29375);
nand UO_3428 (O_3428,N_29412,N_28161);
nor UO_3429 (O_3429,N_29526,N_28782);
and UO_3430 (O_3430,N_28463,N_28490);
nor UO_3431 (O_3431,N_29618,N_29347);
nor UO_3432 (O_3432,N_28377,N_29796);
and UO_3433 (O_3433,N_28470,N_28148);
or UO_3434 (O_3434,N_29485,N_28200);
or UO_3435 (O_3435,N_28085,N_28348);
and UO_3436 (O_3436,N_28179,N_28921);
xnor UO_3437 (O_3437,N_29929,N_28818);
xor UO_3438 (O_3438,N_29641,N_28342);
or UO_3439 (O_3439,N_28028,N_28761);
nand UO_3440 (O_3440,N_29586,N_29173);
or UO_3441 (O_3441,N_28315,N_28938);
and UO_3442 (O_3442,N_29941,N_28067);
and UO_3443 (O_3443,N_29027,N_28255);
or UO_3444 (O_3444,N_28463,N_28045);
xor UO_3445 (O_3445,N_28493,N_28505);
xor UO_3446 (O_3446,N_29871,N_29537);
and UO_3447 (O_3447,N_29794,N_29012);
or UO_3448 (O_3448,N_28781,N_29067);
nand UO_3449 (O_3449,N_29779,N_28866);
nand UO_3450 (O_3450,N_28070,N_28119);
nand UO_3451 (O_3451,N_29728,N_28333);
or UO_3452 (O_3452,N_28941,N_28559);
or UO_3453 (O_3453,N_28421,N_28896);
nand UO_3454 (O_3454,N_29676,N_28063);
or UO_3455 (O_3455,N_28626,N_29009);
nand UO_3456 (O_3456,N_29485,N_28839);
nor UO_3457 (O_3457,N_29784,N_28717);
xnor UO_3458 (O_3458,N_28001,N_29076);
nand UO_3459 (O_3459,N_29722,N_29097);
or UO_3460 (O_3460,N_29881,N_29084);
xnor UO_3461 (O_3461,N_29132,N_29694);
nand UO_3462 (O_3462,N_28880,N_28507);
nand UO_3463 (O_3463,N_29295,N_28556);
nand UO_3464 (O_3464,N_29758,N_28283);
nand UO_3465 (O_3465,N_29686,N_28311);
or UO_3466 (O_3466,N_29489,N_28245);
nor UO_3467 (O_3467,N_28026,N_28842);
and UO_3468 (O_3468,N_28072,N_28602);
nor UO_3469 (O_3469,N_29358,N_29968);
nor UO_3470 (O_3470,N_29432,N_29449);
or UO_3471 (O_3471,N_29573,N_28270);
or UO_3472 (O_3472,N_29648,N_28598);
and UO_3473 (O_3473,N_28259,N_28168);
or UO_3474 (O_3474,N_29082,N_28079);
nand UO_3475 (O_3475,N_28008,N_28866);
and UO_3476 (O_3476,N_28877,N_28186);
xor UO_3477 (O_3477,N_28809,N_29328);
xor UO_3478 (O_3478,N_28229,N_28712);
nand UO_3479 (O_3479,N_28513,N_28034);
and UO_3480 (O_3480,N_28494,N_28775);
nor UO_3481 (O_3481,N_28543,N_29302);
nor UO_3482 (O_3482,N_29175,N_29916);
nor UO_3483 (O_3483,N_29937,N_29010);
and UO_3484 (O_3484,N_29152,N_28953);
and UO_3485 (O_3485,N_29010,N_28570);
xor UO_3486 (O_3486,N_29895,N_28829);
nand UO_3487 (O_3487,N_28765,N_28568);
and UO_3488 (O_3488,N_28254,N_28383);
or UO_3489 (O_3489,N_29252,N_28277);
nand UO_3490 (O_3490,N_28770,N_28609);
or UO_3491 (O_3491,N_29283,N_28766);
nor UO_3492 (O_3492,N_29978,N_29573);
xor UO_3493 (O_3493,N_29315,N_29030);
or UO_3494 (O_3494,N_29076,N_28107);
xnor UO_3495 (O_3495,N_29641,N_29545);
or UO_3496 (O_3496,N_28788,N_28192);
nand UO_3497 (O_3497,N_29523,N_28671);
and UO_3498 (O_3498,N_28304,N_28409);
and UO_3499 (O_3499,N_29367,N_29528);
endmodule