module basic_500_3000_500_4_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_290,In_371);
nand U1 (N_1,In_477,In_252);
or U2 (N_2,In_118,In_77);
nand U3 (N_3,In_144,In_160);
nand U4 (N_4,In_198,In_185);
and U5 (N_5,In_132,In_136);
and U6 (N_6,In_439,In_374);
nand U7 (N_7,In_16,In_358);
and U8 (N_8,In_492,In_129);
and U9 (N_9,In_172,In_363);
or U10 (N_10,In_476,In_366);
nor U11 (N_11,In_383,In_81);
and U12 (N_12,In_458,In_285);
nor U13 (N_13,In_196,In_39);
and U14 (N_14,In_271,In_325);
and U15 (N_15,In_124,In_262);
nand U16 (N_16,In_486,In_170);
and U17 (N_17,In_48,In_121);
and U18 (N_18,In_469,In_320);
nor U19 (N_19,In_137,In_420);
nand U20 (N_20,In_108,In_222);
nor U21 (N_21,In_55,In_394);
nor U22 (N_22,In_369,In_419);
nand U23 (N_23,In_337,In_441);
nor U24 (N_24,In_219,In_207);
nand U25 (N_25,In_499,In_401);
and U26 (N_26,In_115,In_28);
nor U27 (N_27,In_94,In_155);
and U28 (N_28,In_7,In_415);
or U29 (N_29,In_334,In_447);
nand U30 (N_30,In_249,In_340);
nand U31 (N_31,In_350,In_190);
and U32 (N_32,In_86,In_430);
nand U33 (N_33,In_310,In_125);
nor U34 (N_34,In_67,In_311);
or U35 (N_35,In_326,In_82);
nor U36 (N_36,In_327,In_153);
and U37 (N_37,In_215,In_467);
and U38 (N_38,In_385,In_38);
nand U39 (N_39,In_206,In_255);
or U40 (N_40,In_445,In_264);
and U41 (N_41,In_225,In_382);
and U42 (N_42,In_6,In_83);
and U43 (N_43,In_309,In_240);
and U44 (N_44,In_328,In_31);
or U45 (N_45,In_189,In_154);
and U46 (N_46,In_301,In_332);
and U47 (N_47,In_257,In_438);
nand U48 (N_48,In_440,In_29);
nor U49 (N_49,In_140,In_58);
nand U50 (N_50,In_355,In_432);
and U51 (N_51,In_200,In_89);
or U52 (N_52,In_237,In_278);
and U53 (N_53,In_90,In_19);
or U54 (N_54,In_423,In_111);
nand U55 (N_55,In_66,In_135);
nand U56 (N_56,In_316,In_493);
or U57 (N_57,In_209,In_496);
and U58 (N_58,In_417,In_304);
nand U59 (N_59,In_450,In_21);
and U60 (N_60,In_388,In_284);
or U61 (N_61,In_442,In_459);
or U62 (N_62,In_448,In_270);
xnor U63 (N_63,In_345,In_183);
or U64 (N_64,In_169,In_180);
nand U65 (N_65,In_236,In_197);
or U66 (N_66,In_329,In_179);
nand U67 (N_67,In_474,In_147);
or U68 (N_68,In_203,In_3);
nor U69 (N_69,In_338,In_157);
nor U70 (N_70,In_79,In_102);
nand U71 (N_71,In_347,In_488);
or U72 (N_72,In_241,In_312);
nand U73 (N_73,In_12,In_1);
and U74 (N_74,In_24,In_457);
nand U75 (N_75,In_428,In_343);
or U76 (N_76,In_96,In_421);
nand U77 (N_77,In_351,In_25);
nor U78 (N_78,In_498,In_364);
nand U79 (N_79,In_379,In_230);
and U80 (N_80,In_287,In_210);
nand U81 (N_81,In_462,In_78);
or U82 (N_82,In_18,In_396);
nor U83 (N_83,In_75,In_109);
or U84 (N_84,In_391,In_71);
nor U85 (N_85,In_218,In_173);
or U86 (N_86,In_491,In_194);
and U87 (N_87,In_263,In_245);
nand U88 (N_88,In_434,In_231);
or U89 (N_89,In_335,In_489);
and U90 (N_90,In_101,In_168);
nor U91 (N_91,In_100,In_159);
nand U92 (N_92,In_251,In_306);
or U93 (N_93,In_35,In_107);
nand U94 (N_94,In_105,In_409);
and U95 (N_95,In_389,In_233);
nand U96 (N_96,In_45,In_393);
and U97 (N_97,In_289,In_177);
nand U98 (N_98,In_279,In_449);
nor U99 (N_99,In_260,In_110);
nand U100 (N_100,In_324,In_435);
nand U101 (N_101,In_20,In_384);
nor U102 (N_102,In_178,In_53);
and U103 (N_103,In_308,In_473);
and U104 (N_104,In_176,In_76);
nand U105 (N_105,In_127,In_11);
nor U106 (N_106,In_59,In_167);
or U107 (N_107,In_142,In_475);
and U108 (N_108,In_54,In_72);
nor U109 (N_109,In_483,In_214);
nand U110 (N_110,In_114,In_295);
nor U111 (N_111,In_302,In_234);
and U112 (N_112,In_166,In_134);
nor U113 (N_113,In_22,In_92);
or U114 (N_114,In_97,In_119);
or U115 (N_115,In_205,In_112);
or U116 (N_116,In_294,In_85);
nor U117 (N_117,In_162,In_51);
nor U118 (N_118,In_372,In_411);
nor U119 (N_119,In_281,In_481);
or U120 (N_120,In_258,In_2);
or U121 (N_121,In_359,In_485);
or U122 (N_122,In_80,In_116);
and U123 (N_123,In_453,In_303);
or U124 (N_124,In_227,In_288);
or U125 (N_125,In_63,In_37);
nand U126 (N_126,In_380,In_297);
xnor U127 (N_127,In_9,In_269);
nand U128 (N_128,In_201,In_348);
or U129 (N_129,In_452,In_293);
and U130 (N_130,In_305,In_139);
nor U131 (N_131,In_165,In_381);
or U132 (N_132,In_387,In_356);
nand U133 (N_133,In_370,In_199);
and U134 (N_134,In_235,In_392);
and U135 (N_135,In_192,In_26);
nand U136 (N_136,In_404,In_451);
nand U137 (N_137,In_164,In_275);
and U138 (N_138,In_151,In_331);
nand U139 (N_139,In_282,In_149);
or U140 (N_140,In_342,In_368);
and U141 (N_141,In_405,In_276);
or U142 (N_142,In_246,In_436);
nor U143 (N_143,In_454,In_99);
nor U144 (N_144,In_344,In_161);
nor U145 (N_145,In_5,In_88);
and U146 (N_146,In_472,In_175);
nor U147 (N_147,In_74,In_181);
and U148 (N_148,In_463,In_406);
nand U149 (N_149,In_73,In_33);
nand U150 (N_150,In_484,In_422);
or U151 (N_151,In_259,In_333);
or U152 (N_152,In_468,In_213);
nand U153 (N_153,In_23,In_122);
or U154 (N_154,In_182,In_87);
or U155 (N_155,In_433,In_354);
and U156 (N_156,In_283,In_367);
nand U157 (N_157,In_239,In_478);
nor U158 (N_158,In_353,In_52);
and U159 (N_159,In_131,In_70);
nor U160 (N_160,In_323,In_128);
nor U161 (N_161,In_376,In_40);
nor U162 (N_162,In_317,In_318);
nor U163 (N_163,In_130,In_229);
and U164 (N_164,In_431,In_242);
or U165 (N_165,In_98,In_400);
nor U166 (N_166,In_195,In_133);
or U167 (N_167,In_395,In_407);
nand U168 (N_168,In_261,In_8);
nand U169 (N_169,In_444,In_300);
nand U170 (N_170,In_27,In_187);
nand U171 (N_171,In_188,In_126);
nor U172 (N_172,In_408,In_298);
nor U173 (N_173,In_138,In_487);
nand U174 (N_174,In_373,In_224);
nor U175 (N_175,In_314,In_346);
nor U176 (N_176,In_336,In_60);
nand U177 (N_177,In_14,In_437);
xnor U178 (N_178,In_232,In_174);
or U179 (N_179,In_266,In_322);
and U180 (N_180,In_91,In_57);
nand U181 (N_181,In_313,In_216);
nor U182 (N_182,In_184,In_460);
nand U183 (N_183,In_41,In_455);
nor U184 (N_184,In_402,In_254);
and U185 (N_185,In_268,In_193);
and U186 (N_186,In_32,In_291);
and U187 (N_187,In_386,In_247);
nand U188 (N_188,In_141,In_339);
or U189 (N_189,In_470,In_43);
nand U190 (N_190,In_117,In_223);
nor U191 (N_191,In_123,In_471);
nor U192 (N_192,In_321,In_10);
and U193 (N_193,In_145,In_464);
nor U194 (N_194,In_265,In_0);
and U195 (N_195,In_365,In_482);
and U196 (N_196,In_418,In_106);
nand U197 (N_197,In_150,In_248);
or U198 (N_198,In_349,In_228);
nand U199 (N_199,In_62,In_34);
nor U200 (N_200,In_158,In_103);
nand U201 (N_201,In_36,In_93);
and U202 (N_202,In_480,In_42);
or U203 (N_203,In_64,In_427);
or U204 (N_204,In_148,In_113);
or U205 (N_205,In_208,In_410);
or U206 (N_206,In_497,In_211);
nand U207 (N_207,In_30,In_299);
and U208 (N_208,In_362,In_466);
nand U209 (N_209,In_250,In_120);
or U210 (N_210,In_479,In_416);
nor U211 (N_211,In_163,In_56);
and U212 (N_212,In_413,In_104);
nor U213 (N_213,In_267,In_378);
and U214 (N_214,In_49,In_465);
and U215 (N_215,In_13,In_15);
or U216 (N_216,In_244,In_273);
nand U217 (N_217,In_330,In_95);
and U218 (N_218,In_357,In_461);
and U219 (N_219,In_352,In_286);
nand U220 (N_220,In_253,In_319);
or U221 (N_221,In_84,In_204);
nand U222 (N_222,In_17,In_212);
nor U223 (N_223,In_292,In_341);
or U224 (N_224,In_47,In_429);
and U225 (N_225,In_61,In_274);
and U226 (N_226,In_307,In_146);
nor U227 (N_227,In_226,In_424);
nand U228 (N_228,In_143,In_46);
and U229 (N_229,In_217,In_272);
and U230 (N_230,In_377,In_397);
and U231 (N_231,In_296,In_202);
and U232 (N_232,In_44,In_65);
and U233 (N_233,In_375,In_156);
nand U234 (N_234,In_446,In_238);
nand U235 (N_235,In_403,In_414);
nand U236 (N_236,In_68,In_243);
or U237 (N_237,In_443,In_50);
nor U238 (N_238,In_152,In_495);
and U239 (N_239,In_426,In_277);
nand U240 (N_240,In_315,In_425);
nor U241 (N_241,In_256,In_399);
nor U242 (N_242,In_390,In_412);
and U243 (N_243,In_69,In_4);
nor U244 (N_244,In_361,In_456);
or U245 (N_245,In_186,In_171);
nand U246 (N_246,In_494,In_221);
or U247 (N_247,In_360,In_220);
and U248 (N_248,In_280,In_490);
nand U249 (N_249,In_191,In_398);
nor U250 (N_250,In_132,In_440);
or U251 (N_251,In_275,In_310);
or U252 (N_252,In_366,In_133);
and U253 (N_253,In_328,In_295);
and U254 (N_254,In_388,In_421);
and U255 (N_255,In_112,In_332);
nor U256 (N_256,In_452,In_29);
nand U257 (N_257,In_83,In_199);
nor U258 (N_258,In_46,In_481);
nor U259 (N_259,In_306,In_184);
and U260 (N_260,In_292,In_361);
nor U261 (N_261,In_234,In_158);
nand U262 (N_262,In_321,In_431);
and U263 (N_263,In_220,In_265);
nor U264 (N_264,In_32,In_262);
and U265 (N_265,In_377,In_335);
nor U266 (N_266,In_422,In_436);
nor U267 (N_267,In_377,In_275);
or U268 (N_268,In_96,In_308);
and U269 (N_269,In_486,In_412);
nand U270 (N_270,In_284,In_156);
nor U271 (N_271,In_255,In_384);
nor U272 (N_272,In_459,In_63);
and U273 (N_273,In_158,In_140);
or U274 (N_274,In_163,In_332);
or U275 (N_275,In_127,In_403);
nor U276 (N_276,In_153,In_319);
and U277 (N_277,In_101,In_143);
nand U278 (N_278,In_200,In_431);
nor U279 (N_279,In_343,In_26);
nand U280 (N_280,In_76,In_443);
and U281 (N_281,In_275,In_172);
nand U282 (N_282,In_253,In_86);
or U283 (N_283,In_333,In_405);
nor U284 (N_284,In_83,In_425);
nor U285 (N_285,In_281,In_487);
nor U286 (N_286,In_137,In_176);
nand U287 (N_287,In_35,In_322);
nand U288 (N_288,In_283,In_477);
and U289 (N_289,In_63,In_25);
nand U290 (N_290,In_498,In_331);
nor U291 (N_291,In_386,In_26);
nor U292 (N_292,In_294,In_316);
and U293 (N_293,In_359,In_93);
and U294 (N_294,In_305,In_259);
and U295 (N_295,In_360,In_259);
nand U296 (N_296,In_163,In_309);
nor U297 (N_297,In_471,In_334);
nand U298 (N_298,In_166,In_494);
or U299 (N_299,In_300,In_144);
and U300 (N_300,In_301,In_433);
or U301 (N_301,In_184,In_205);
or U302 (N_302,In_468,In_199);
or U303 (N_303,In_129,In_83);
nand U304 (N_304,In_43,In_210);
or U305 (N_305,In_436,In_240);
nand U306 (N_306,In_279,In_176);
xor U307 (N_307,In_283,In_117);
nor U308 (N_308,In_331,In_344);
nor U309 (N_309,In_359,In_112);
and U310 (N_310,In_90,In_469);
and U311 (N_311,In_162,In_44);
or U312 (N_312,In_311,In_382);
or U313 (N_313,In_475,In_456);
nand U314 (N_314,In_251,In_250);
nand U315 (N_315,In_117,In_118);
or U316 (N_316,In_373,In_390);
and U317 (N_317,In_481,In_305);
and U318 (N_318,In_334,In_121);
nor U319 (N_319,In_430,In_422);
or U320 (N_320,In_361,In_174);
nor U321 (N_321,In_29,In_164);
nand U322 (N_322,In_138,In_139);
and U323 (N_323,In_412,In_458);
nand U324 (N_324,In_10,In_268);
nor U325 (N_325,In_80,In_430);
nand U326 (N_326,In_145,In_245);
nand U327 (N_327,In_457,In_483);
or U328 (N_328,In_278,In_157);
nand U329 (N_329,In_156,In_171);
nor U330 (N_330,In_332,In_251);
nor U331 (N_331,In_40,In_111);
nor U332 (N_332,In_310,In_446);
or U333 (N_333,In_125,In_430);
or U334 (N_334,In_8,In_141);
nor U335 (N_335,In_381,In_34);
nand U336 (N_336,In_108,In_110);
nand U337 (N_337,In_378,In_93);
nand U338 (N_338,In_178,In_405);
or U339 (N_339,In_191,In_181);
or U340 (N_340,In_179,In_139);
or U341 (N_341,In_37,In_462);
or U342 (N_342,In_378,In_322);
and U343 (N_343,In_245,In_114);
nand U344 (N_344,In_110,In_434);
nor U345 (N_345,In_168,In_22);
or U346 (N_346,In_411,In_322);
nor U347 (N_347,In_345,In_356);
and U348 (N_348,In_137,In_427);
nand U349 (N_349,In_260,In_72);
and U350 (N_350,In_417,In_245);
or U351 (N_351,In_140,In_445);
nand U352 (N_352,In_255,In_498);
and U353 (N_353,In_395,In_107);
and U354 (N_354,In_243,In_212);
nor U355 (N_355,In_403,In_399);
or U356 (N_356,In_444,In_338);
nand U357 (N_357,In_324,In_268);
and U358 (N_358,In_164,In_161);
nand U359 (N_359,In_3,In_464);
and U360 (N_360,In_337,In_489);
nor U361 (N_361,In_406,In_72);
nand U362 (N_362,In_415,In_375);
nor U363 (N_363,In_405,In_23);
and U364 (N_364,In_97,In_25);
nand U365 (N_365,In_37,In_379);
and U366 (N_366,In_221,In_258);
nor U367 (N_367,In_179,In_424);
and U368 (N_368,In_274,In_72);
nand U369 (N_369,In_64,In_306);
nor U370 (N_370,In_246,In_345);
or U371 (N_371,In_118,In_367);
nor U372 (N_372,In_253,In_452);
nor U373 (N_373,In_412,In_117);
and U374 (N_374,In_7,In_64);
nand U375 (N_375,In_336,In_274);
nand U376 (N_376,In_189,In_322);
and U377 (N_377,In_148,In_391);
or U378 (N_378,In_426,In_184);
and U379 (N_379,In_103,In_333);
nand U380 (N_380,In_286,In_115);
nand U381 (N_381,In_165,In_432);
or U382 (N_382,In_372,In_239);
or U383 (N_383,In_421,In_203);
nand U384 (N_384,In_447,In_346);
or U385 (N_385,In_101,In_474);
nor U386 (N_386,In_86,In_101);
and U387 (N_387,In_28,In_201);
nand U388 (N_388,In_233,In_225);
and U389 (N_389,In_148,In_139);
nand U390 (N_390,In_494,In_191);
xnor U391 (N_391,In_104,In_473);
nand U392 (N_392,In_93,In_191);
nand U393 (N_393,In_264,In_404);
or U394 (N_394,In_439,In_201);
nand U395 (N_395,In_472,In_107);
nor U396 (N_396,In_149,In_309);
and U397 (N_397,In_82,In_224);
nand U398 (N_398,In_40,In_472);
nand U399 (N_399,In_24,In_353);
nand U400 (N_400,In_456,In_119);
and U401 (N_401,In_391,In_221);
nand U402 (N_402,In_298,In_282);
and U403 (N_403,In_363,In_153);
nor U404 (N_404,In_498,In_27);
nand U405 (N_405,In_70,In_11);
nor U406 (N_406,In_52,In_111);
and U407 (N_407,In_331,In_66);
nand U408 (N_408,In_38,In_339);
nand U409 (N_409,In_300,In_459);
nand U410 (N_410,In_477,In_141);
or U411 (N_411,In_169,In_7);
and U412 (N_412,In_438,In_84);
nand U413 (N_413,In_479,In_417);
or U414 (N_414,In_191,In_204);
nand U415 (N_415,In_451,In_143);
nor U416 (N_416,In_142,In_202);
nor U417 (N_417,In_56,In_395);
nor U418 (N_418,In_435,In_332);
nor U419 (N_419,In_451,In_495);
and U420 (N_420,In_210,In_261);
and U421 (N_421,In_326,In_12);
or U422 (N_422,In_111,In_391);
or U423 (N_423,In_268,In_170);
nor U424 (N_424,In_192,In_36);
or U425 (N_425,In_270,In_59);
and U426 (N_426,In_432,In_414);
nor U427 (N_427,In_168,In_136);
nor U428 (N_428,In_455,In_485);
and U429 (N_429,In_117,In_126);
and U430 (N_430,In_486,In_441);
nor U431 (N_431,In_58,In_192);
or U432 (N_432,In_395,In_79);
or U433 (N_433,In_64,In_135);
and U434 (N_434,In_288,In_106);
nor U435 (N_435,In_6,In_475);
or U436 (N_436,In_264,In_2);
nand U437 (N_437,In_309,In_221);
or U438 (N_438,In_403,In_383);
or U439 (N_439,In_195,In_101);
and U440 (N_440,In_474,In_437);
and U441 (N_441,In_419,In_383);
nand U442 (N_442,In_91,In_201);
nor U443 (N_443,In_92,In_458);
nand U444 (N_444,In_218,In_198);
nand U445 (N_445,In_88,In_36);
nor U446 (N_446,In_275,In_262);
nand U447 (N_447,In_229,In_55);
or U448 (N_448,In_322,In_335);
and U449 (N_449,In_307,In_196);
and U450 (N_450,In_85,In_231);
nand U451 (N_451,In_365,In_472);
nor U452 (N_452,In_238,In_422);
nand U453 (N_453,In_296,In_142);
nor U454 (N_454,In_430,In_394);
nor U455 (N_455,In_167,In_115);
or U456 (N_456,In_205,In_466);
nor U457 (N_457,In_370,In_292);
nor U458 (N_458,In_197,In_173);
nand U459 (N_459,In_312,In_373);
nor U460 (N_460,In_266,In_42);
nor U461 (N_461,In_273,In_348);
nand U462 (N_462,In_14,In_199);
nand U463 (N_463,In_28,In_209);
and U464 (N_464,In_85,In_286);
nand U465 (N_465,In_303,In_256);
nand U466 (N_466,In_200,In_477);
nor U467 (N_467,In_445,In_22);
or U468 (N_468,In_454,In_399);
nand U469 (N_469,In_66,In_330);
or U470 (N_470,In_475,In_14);
nand U471 (N_471,In_154,In_46);
nor U472 (N_472,In_0,In_346);
nand U473 (N_473,In_74,In_269);
or U474 (N_474,In_21,In_238);
nand U475 (N_475,In_21,In_341);
and U476 (N_476,In_225,In_201);
or U477 (N_477,In_272,In_297);
and U478 (N_478,In_347,In_23);
or U479 (N_479,In_176,In_2);
nand U480 (N_480,In_263,In_181);
or U481 (N_481,In_117,In_407);
or U482 (N_482,In_183,In_186);
nand U483 (N_483,In_97,In_150);
or U484 (N_484,In_312,In_498);
or U485 (N_485,In_332,In_279);
and U486 (N_486,In_382,In_171);
nor U487 (N_487,In_287,In_258);
nand U488 (N_488,In_181,In_242);
nand U489 (N_489,In_98,In_261);
nand U490 (N_490,In_455,In_184);
nand U491 (N_491,In_349,In_239);
and U492 (N_492,In_494,In_296);
xor U493 (N_493,In_353,In_94);
and U494 (N_494,In_349,In_196);
nand U495 (N_495,In_414,In_280);
or U496 (N_496,In_134,In_145);
nand U497 (N_497,In_310,In_97);
nor U498 (N_498,In_70,In_89);
nor U499 (N_499,In_196,In_249);
or U500 (N_500,In_156,In_266);
nor U501 (N_501,In_211,In_374);
and U502 (N_502,In_124,In_288);
and U503 (N_503,In_194,In_283);
and U504 (N_504,In_394,In_149);
nand U505 (N_505,In_422,In_229);
nand U506 (N_506,In_205,In_490);
or U507 (N_507,In_353,In_6);
or U508 (N_508,In_242,In_239);
and U509 (N_509,In_372,In_363);
or U510 (N_510,In_441,In_68);
and U511 (N_511,In_328,In_121);
nor U512 (N_512,In_418,In_274);
and U513 (N_513,In_70,In_114);
and U514 (N_514,In_383,In_301);
or U515 (N_515,In_48,In_41);
or U516 (N_516,In_260,In_111);
xnor U517 (N_517,In_209,In_435);
nor U518 (N_518,In_122,In_209);
nor U519 (N_519,In_462,In_160);
and U520 (N_520,In_129,In_264);
nor U521 (N_521,In_463,In_455);
nand U522 (N_522,In_184,In_112);
nand U523 (N_523,In_27,In_121);
or U524 (N_524,In_342,In_485);
nand U525 (N_525,In_260,In_418);
nor U526 (N_526,In_105,In_57);
and U527 (N_527,In_120,In_62);
and U528 (N_528,In_53,In_405);
or U529 (N_529,In_70,In_262);
nor U530 (N_530,In_151,In_275);
or U531 (N_531,In_78,In_263);
nand U532 (N_532,In_431,In_186);
or U533 (N_533,In_198,In_116);
nand U534 (N_534,In_434,In_375);
nand U535 (N_535,In_193,In_143);
nor U536 (N_536,In_303,In_207);
nand U537 (N_537,In_391,In_479);
nor U538 (N_538,In_66,In_163);
and U539 (N_539,In_185,In_104);
nand U540 (N_540,In_56,In_236);
and U541 (N_541,In_441,In_251);
nor U542 (N_542,In_226,In_303);
and U543 (N_543,In_4,In_249);
nand U544 (N_544,In_104,In_293);
nor U545 (N_545,In_359,In_12);
and U546 (N_546,In_2,In_164);
nor U547 (N_547,In_64,In_494);
xor U548 (N_548,In_14,In_364);
or U549 (N_549,In_65,In_315);
or U550 (N_550,In_499,In_43);
nor U551 (N_551,In_174,In_212);
nand U552 (N_552,In_321,In_253);
and U553 (N_553,In_407,In_177);
and U554 (N_554,In_165,In_293);
or U555 (N_555,In_116,In_306);
nor U556 (N_556,In_181,In_444);
nand U557 (N_557,In_346,In_126);
and U558 (N_558,In_23,In_50);
and U559 (N_559,In_8,In_47);
or U560 (N_560,In_42,In_73);
and U561 (N_561,In_488,In_106);
or U562 (N_562,In_56,In_11);
nand U563 (N_563,In_141,In_366);
nor U564 (N_564,In_149,In_137);
and U565 (N_565,In_244,In_187);
or U566 (N_566,In_106,In_323);
and U567 (N_567,In_404,In_341);
nor U568 (N_568,In_94,In_337);
nand U569 (N_569,In_98,In_416);
nor U570 (N_570,In_89,In_239);
nor U571 (N_571,In_245,In_146);
or U572 (N_572,In_469,In_467);
nand U573 (N_573,In_487,In_420);
nor U574 (N_574,In_388,In_177);
nor U575 (N_575,In_391,In_436);
nand U576 (N_576,In_428,In_50);
and U577 (N_577,In_27,In_46);
or U578 (N_578,In_355,In_43);
or U579 (N_579,In_88,In_26);
nor U580 (N_580,In_78,In_149);
or U581 (N_581,In_76,In_236);
or U582 (N_582,In_477,In_249);
nor U583 (N_583,In_437,In_145);
nand U584 (N_584,In_292,In_496);
nand U585 (N_585,In_102,In_324);
or U586 (N_586,In_386,In_296);
nand U587 (N_587,In_382,In_328);
nor U588 (N_588,In_293,In_493);
and U589 (N_589,In_173,In_125);
or U590 (N_590,In_436,In_340);
or U591 (N_591,In_394,In_486);
nor U592 (N_592,In_2,In_240);
nor U593 (N_593,In_431,In_454);
or U594 (N_594,In_316,In_416);
nand U595 (N_595,In_120,In_79);
nor U596 (N_596,In_498,In_128);
or U597 (N_597,In_442,In_334);
and U598 (N_598,In_121,In_160);
or U599 (N_599,In_442,In_315);
nor U600 (N_600,In_274,In_303);
nand U601 (N_601,In_98,In_366);
or U602 (N_602,In_266,In_165);
and U603 (N_603,In_376,In_282);
or U604 (N_604,In_318,In_303);
or U605 (N_605,In_335,In_326);
nor U606 (N_606,In_52,In_5);
nor U607 (N_607,In_91,In_398);
nor U608 (N_608,In_74,In_385);
nand U609 (N_609,In_446,In_296);
nor U610 (N_610,In_430,In_60);
nor U611 (N_611,In_214,In_427);
nor U612 (N_612,In_184,In_250);
nor U613 (N_613,In_453,In_369);
nand U614 (N_614,In_264,In_373);
and U615 (N_615,In_357,In_486);
nand U616 (N_616,In_438,In_128);
or U617 (N_617,In_46,In_156);
xnor U618 (N_618,In_170,In_252);
or U619 (N_619,In_404,In_280);
and U620 (N_620,In_402,In_306);
nor U621 (N_621,In_98,In_51);
or U622 (N_622,In_161,In_45);
nor U623 (N_623,In_454,In_321);
nand U624 (N_624,In_203,In_479);
or U625 (N_625,In_348,In_14);
xor U626 (N_626,In_66,In_407);
or U627 (N_627,In_201,In_147);
nor U628 (N_628,In_491,In_250);
nor U629 (N_629,In_83,In_50);
and U630 (N_630,In_340,In_73);
nor U631 (N_631,In_59,In_127);
nor U632 (N_632,In_147,In_145);
nand U633 (N_633,In_448,In_69);
and U634 (N_634,In_173,In_33);
and U635 (N_635,In_442,In_184);
or U636 (N_636,In_180,In_425);
or U637 (N_637,In_465,In_212);
and U638 (N_638,In_416,In_63);
nor U639 (N_639,In_101,In_126);
or U640 (N_640,In_333,In_46);
nand U641 (N_641,In_452,In_61);
and U642 (N_642,In_227,In_246);
nand U643 (N_643,In_95,In_278);
nand U644 (N_644,In_106,In_57);
nand U645 (N_645,In_410,In_234);
nand U646 (N_646,In_434,In_437);
nand U647 (N_647,In_39,In_402);
or U648 (N_648,In_345,In_451);
or U649 (N_649,In_35,In_104);
and U650 (N_650,In_113,In_471);
nor U651 (N_651,In_80,In_92);
nor U652 (N_652,In_412,In_155);
nor U653 (N_653,In_303,In_370);
nor U654 (N_654,In_289,In_205);
nor U655 (N_655,In_98,In_374);
or U656 (N_656,In_243,In_412);
nand U657 (N_657,In_484,In_457);
or U658 (N_658,In_13,In_307);
and U659 (N_659,In_64,In_219);
nand U660 (N_660,In_298,In_422);
and U661 (N_661,In_390,In_243);
nand U662 (N_662,In_356,In_13);
nand U663 (N_663,In_467,In_184);
nand U664 (N_664,In_356,In_474);
nand U665 (N_665,In_15,In_81);
or U666 (N_666,In_254,In_490);
or U667 (N_667,In_446,In_54);
nor U668 (N_668,In_231,In_191);
or U669 (N_669,In_335,In_446);
nand U670 (N_670,In_171,In_195);
nor U671 (N_671,In_37,In_240);
nor U672 (N_672,In_145,In_307);
or U673 (N_673,In_267,In_7);
nor U674 (N_674,In_404,In_395);
or U675 (N_675,In_416,In_214);
or U676 (N_676,In_245,In_140);
nand U677 (N_677,In_225,In_303);
or U678 (N_678,In_38,In_120);
or U679 (N_679,In_298,In_358);
nor U680 (N_680,In_160,In_69);
nand U681 (N_681,In_218,In_442);
nand U682 (N_682,In_362,In_103);
nor U683 (N_683,In_335,In_275);
and U684 (N_684,In_105,In_106);
and U685 (N_685,In_61,In_436);
and U686 (N_686,In_137,In_411);
nor U687 (N_687,In_67,In_390);
nor U688 (N_688,In_245,In_7);
and U689 (N_689,In_146,In_493);
nor U690 (N_690,In_233,In_304);
nand U691 (N_691,In_229,In_342);
nor U692 (N_692,In_124,In_68);
nand U693 (N_693,In_6,In_389);
nor U694 (N_694,In_41,In_157);
or U695 (N_695,In_47,In_141);
nor U696 (N_696,In_169,In_267);
or U697 (N_697,In_303,In_28);
and U698 (N_698,In_425,In_155);
nor U699 (N_699,In_12,In_442);
nor U700 (N_700,In_391,In_266);
and U701 (N_701,In_84,In_162);
and U702 (N_702,In_333,In_189);
or U703 (N_703,In_455,In_116);
nand U704 (N_704,In_423,In_484);
nor U705 (N_705,In_474,In_163);
nor U706 (N_706,In_295,In_281);
or U707 (N_707,In_488,In_356);
and U708 (N_708,In_229,In_49);
nand U709 (N_709,In_238,In_305);
or U710 (N_710,In_53,In_431);
or U711 (N_711,In_386,In_39);
nor U712 (N_712,In_137,In_362);
or U713 (N_713,In_401,In_32);
nand U714 (N_714,In_197,In_468);
or U715 (N_715,In_126,In_184);
or U716 (N_716,In_81,In_146);
nand U717 (N_717,In_462,In_127);
nand U718 (N_718,In_25,In_227);
or U719 (N_719,In_445,In_325);
nor U720 (N_720,In_454,In_417);
nand U721 (N_721,In_359,In_274);
or U722 (N_722,In_155,In_441);
or U723 (N_723,In_49,In_257);
or U724 (N_724,In_291,In_42);
or U725 (N_725,In_180,In_9);
nor U726 (N_726,In_8,In_51);
or U727 (N_727,In_193,In_277);
nand U728 (N_728,In_402,In_325);
and U729 (N_729,In_34,In_417);
and U730 (N_730,In_132,In_122);
and U731 (N_731,In_403,In_478);
or U732 (N_732,In_183,In_50);
nand U733 (N_733,In_324,In_245);
or U734 (N_734,In_136,In_157);
and U735 (N_735,In_168,In_226);
or U736 (N_736,In_191,In_461);
or U737 (N_737,In_387,In_292);
nand U738 (N_738,In_438,In_132);
nand U739 (N_739,In_186,In_40);
or U740 (N_740,In_20,In_372);
and U741 (N_741,In_5,In_289);
nor U742 (N_742,In_305,In_218);
nor U743 (N_743,In_131,In_151);
nor U744 (N_744,In_380,In_315);
nor U745 (N_745,In_86,In_88);
nor U746 (N_746,In_92,In_96);
or U747 (N_747,In_0,In_68);
and U748 (N_748,In_195,In_151);
nor U749 (N_749,In_430,In_140);
nor U750 (N_750,N_538,N_202);
nor U751 (N_751,N_490,N_59);
nor U752 (N_752,N_470,N_55);
nor U753 (N_753,N_38,N_484);
and U754 (N_754,N_270,N_647);
nand U755 (N_755,N_672,N_707);
and U756 (N_756,N_366,N_521);
or U757 (N_757,N_548,N_455);
and U758 (N_758,N_699,N_730);
or U759 (N_759,N_466,N_279);
or U760 (N_760,N_680,N_549);
nand U761 (N_761,N_284,N_423);
nor U762 (N_762,N_507,N_329);
and U763 (N_763,N_495,N_491);
or U764 (N_764,N_666,N_583);
or U765 (N_765,N_518,N_163);
nor U766 (N_766,N_693,N_531);
xnor U767 (N_767,N_453,N_405);
nand U768 (N_768,N_736,N_432);
and U769 (N_769,N_170,N_90);
nor U770 (N_770,N_537,N_221);
and U771 (N_771,N_683,N_635);
nor U772 (N_772,N_649,N_522);
nor U773 (N_773,N_558,N_586);
and U774 (N_774,N_665,N_189);
nor U775 (N_775,N_724,N_261);
or U776 (N_776,N_344,N_91);
and U777 (N_777,N_292,N_361);
nor U778 (N_778,N_323,N_76);
or U779 (N_779,N_561,N_438);
or U780 (N_780,N_158,N_420);
nor U781 (N_781,N_121,N_543);
nand U782 (N_782,N_81,N_689);
nor U783 (N_783,N_267,N_749);
and U784 (N_784,N_424,N_360);
and U785 (N_785,N_480,N_479);
xor U786 (N_786,N_728,N_464);
nand U787 (N_787,N_550,N_618);
or U788 (N_788,N_250,N_732);
nand U789 (N_789,N_0,N_118);
and U790 (N_790,N_153,N_726);
or U791 (N_791,N_311,N_238);
nand U792 (N_792,N_51,N_98);
or U793 (N_793,N_79,N_559);
nor U794 (N_794,N_717,N_129);
and U795 (N_795,N_474,N_700);
nand U796 (N_796,N_506,N_535);
nand U797 (N_797,N_191,N_27);
or U798 (N_798,N_530,N_504);
or U799 (N_799,N_166,N_723);
or U800 (N_800,N_540,N_727);
or U801 (N_801,N_290,N_579);
and U802 (N_802,N_572,N_454);
or U803 (N_803,N_46,N_78);
nor U804 (N_804,N_255,N_167);
or U805 (N_805,N_607,N_89);
nand U806 (N_806,N_557,N_513);
or U807 (N_807,N_140,N_379);
and U808 (N_808,N_519,N_492);
nand U809 (N_809,N_678,N_65);
nand U810 (N_810,N_425,N_375);
nor U811 (N_811,N_141,N_355);
or U812 (N_812,N_475,N_539);
nand U813 (N_813,N_211,N_112);
or U814 (N_814,N_239,N_62);
and U815 (N_815,N_199,N_485);
nor U816 (N_816,N_127,N_315);
nor U817 (N_817,N_263,N_101);
and U818 (N_818,N_12,N_372);
and U819 (N_819,N_251,N_87);
or U820 (N_820,N_57,N_23);
or U821 (N_821,N_264,N_482);
or U822 (N_822,N_247,N_578);
nor U823 (N_823,N_354,N_88);
and U824 (N_824,N_456,N_103);
nand U825 (N_825,N_526,N_5);
or U826 (N_826,N_402,N_676);
and U827 (N_827,N_532,N_681);
or U828 (N_828,N_658,N_622);
nand U829 (N_829,N_407,N_256);
and U830 (N_830,N_688,N_626);
nand U831 (N_831,N_444,N_210);
nor U832 (N_832,N_100,N_515);
nor U833 (N_833,N_242,N_204);
nor U834 (N_834,N_75,N_660);
or U835 (N_835,N_745,N_68);
nand U836 (N_836,N_613,N_185);
or U837 (N_837,N_54,N_184);
or U838 (N_838,N_725,N_157);
nor U839 (N_839,N_107,N_236);
xnor U840 (N_840,N_505,N_708);
or U841 (N_841,N_556,N_640);
nor U842 (N_842,N_226,N_419);
nand U843 (N_843,N_368,N_350);
or U844 (N_844,N_536,N_294);
nor U845 (N_845,N_9,N_437);
nor U846 (N_846,N_188,N_318);
nand U847 (N_847,N_327,N_70);
nand U848 (N_848,N_664,N_394);
and U849 (N_849,N_200,N_661);
or U850 (N_850,N_308,N_174);
or U851 (N_851,N_194,N_214);
and U852 (N_852,N_377,N_248);
or U853 (N_853,N_254,N_671);
xor U854 (N_854,N_276,N_60);
or U855 (N_855,N_400,N_509);
nand U856 (N_856,N_47,N_147);
nand U857 (N_857,N_443,N_172);
nor U858 (N_858,N_614,N_123);
and U859 (N_859,N_703,N_348);
or U860 (N_860,N_209,N_48);
or U861 (N_861,N_326,N_392);
and U862 (N_862,N_77,N_159);
or U863 (N_863,N_208,N_523);
nor U864 (N_864,N_654,N_351);
nor U865 (N_865,N_233,N_342);
and U866 (N_866,N_566,N_670);
nand U867 (N_867,N_334,N_748);
and U868 (N_868,N_577,N_310);
nor U869 (N_869,N_300,N_501);
and U870 (N_870,N_154,N_84);
nand U871 (N_871,N_656,N_487);
and U872 (N_872,N_554,N_29);
or U873 (N_873,N_97,N_207);
nor U874 (N_874,N_24,N_620);
and U875 (N_875,N_374,N_731);
and U876 (N_876,N_94,N_433);
or U877 (N_877,N_85,N_388);
nor U878 (N_878,N_391,N_738);
nand U879 (N_879,N_600,N_674);
nand U880 (N_880,N_232,N_186);
and U881 (N_881,N_410,N_369);
nand U882 (N_882,N_376,N_52);
or U883 (N_883,N_150,N_692);
and U884 (N_884,N_499,N_469);
nand U885 (N_885,N_219,N_713);
nor U886 (N_886,N_357,N_220);
nor U887 (N_887,N_393,N_295);
and U888 (N_888,N_177,N_687);
and U889 (N_889,N_50,N_213);
nor U890 (N_890,N_414,N_293);
nand U891 (N_891,N_546,N_152);
nor U892 (N_892,N_337,N_603);
or U893 (N_893,N_216,N_462);
or U894 (N_894,N_581,N_698);
and U895 (N_895,N_445,N_307);
and U896 (N_896,N_222,N_229);
or U897 (N_897,N_696,N_472);
nor U898 (N_898,N_710,N_215);
or U899 (N_899,N_584,N_631);
and U900 (N_900,N_356,N_109);
and U901 (N_901,N_133,N_195);
or U902 (N_902,N_468,N_347);
nand U903 (N_903,N_162,N_134);
nand U904 (N_904,N_440,N_244);
nor U905 (N_905,N_64,N_617);
nor U906 (N_906,N_695,N_234);
nor U907 (N_907,N_471,N_714);
nand U908 (N_908,N_639,N_137);
or U909 (N_909,N_616,N_381);
nor U910 (N_910,N_142,N_49);
or U911 (N_911,N_42,N_227);
nor U912 (N_912,N_161,N_26);
or U913 (N_913,N_297,N_431);
and U914 (N_914,N_534,N_585);
nor U915 (N_915,N_573,N_225);
nor U916 (N_916,N_608,N_320);
and U917 (N_917,N_179,N_733);
nand U918 (N_918,N_183,N_588);
nand U919 (N_919,N_319,N_739);
nor U920 (N_920,N_458,N_31);
and U921 (N_921,N_44,N_675);
nor U922 (N_922,N_359,N_593);
or U923 (N_923,N_570,N_669);
nand U924 (N_924,N_612,N_529);
and U925 (N_925,N_596,N_429);
or U926 (N_926,N_571,N_122);
and U927 (N_927,N_560,N_637);
and U928 (N_928,N_110,N_190);
and U929 (N_929,N_321,N_69);
nor U930 (N_930,N_569,N_230);
and U931 (N_931,N_605,N_168);
and U932 (N_932,N_14,N_217);
and U933 (N_933,N_690,N_564);
and U934 (N_934,N_58,N_17);
nor U935 (N_935,N_32,N_131);
nor U936 (N_936,N_511,N_611);
and U937 (N_937,N_16,N_604);
nand U938 (N_938,N_340,N_349);
and U939 (N_939,N_187,N_35);
or U940 (N_940,N_587,N_173);
or U941 (N_941,N_63,N_231);
and U942 (N_942,N_574,N_237);
and U943 (N_943,N_117,N_61);
nand U944 (N_944,N_737,N_503);
nand U945 (N_945,N_599,N_332);
and U946 (N_946,N_144,N_324);
nand U947 (N_947,N_746,N_408);
or U948 (N_948,N_205,N_165);
nand U949 (N_949,N_104,N_288);
nor U950 (N_950,N_642,N_274);
and U951 (N_951,N_615,N_95);
and U952 (N_952,N_312,N_448);
nor U953 (N_953,N_22,N_113);
nor U954 (N_954,N_296,N_386);
nor U955 (N_955,N_404,N_592);
nand U956 (N_956,N_673,N_528);
nand U957 (N_957,N_459,N_245);
nor U958 (N_958,N_457,N_668);
nand U959 (N_959,N_304,N_151);
or U960 (N_960,N_363,N_335);
or U961 (N_961,N_228,N_265);
nand U962 (N_962,N_426,N_260);
nor U963 (N_963,N_744,N_353);
nor U964 (N_964,N_650,N_175);
and U965 (N_965,N_281,N_533);
and U966 (N_966,N_275,N_662);
nand U967 (N_967,N_120,N_269);
nand U968 (N_968,N_148,N_544);
or U969 (N_969,N_277,N_625);
or U970 (N_970,N_145,N_115);
nand U971 (N_971,N_383,N_253);
and U972 (N_972,N_271,N_206);
and U973 (N_973,N_380,N_126);
and U974 (N_974,N_305,N_2);
nand U975 (N_975,N_385,N_715);
or U976 (N_976,N_378,N_447);
nor U977 (N_977,N_346,N_283);
or U978 (N_978,N_677,N_56);
or U979 (N_979,N_13,N_125);
and U980 (N_980,N_705,N_412);
nand U981 (N_981,N_33,N_11);
nor U982 (N_982,N_246,N_352);
and U983 (N_983,N_224,N_73);
and U984 (N_984,N_439,N_72);
or U985 (N_985,N_436,N_709);
xor U986 (N_986,N_461,N_20);
nor U987 (N_987,N_657,N_694);
and U988 (N_988,N_644,N_465);
nand U989 (N_989,N_590,N_718);
nor U990 (N_990,N_623,N_740);
nor U991 (N_991,N_496,N_362);
nor U992 (N_992,N_476,N_735);
nand U993 (N_993,N_146,N_595);
and U994 (N_994,N_358,N_1);
nand U995 (N_995,N_80,N_446);
or U996 (N_996,N_627,N_132);
or U997 (N_997,N_712,N_638);
nor U998 (N_998,N_435,N_527);
nand U999 (N_999,N_682,N_336);
nor U1000 (N_1000,N_367,N_428);
or U1001 (N_1001,N_92,N_629);
nand U1002 (N_1002,N_430,N_542);
or U1003 (N_1003,N_169,N_96);
or U1004 (N_1004,N_413,N_722);
nor U1005 (N_1005,N_82,N_520);
or U1006 (N_1006,N_258,N_602);
nand U1007 (N_1007,N_494,N_299);
and U1008 (N_1008,N_401,N_636);
or U1009 (N_1009,N_719,N_711);
or U1010 (N_1010,N_164,N_619);
nor U1011 (N_1011,N_382,N_450);
and U1012 (N_1012,N_39,N_365);
nor U1013 (N_1013,N_734,N_591);
nand U1014 (N_1014,N_241,N_411);
nand U1015 (N_1015,N_317,N_697);
or U1016 (N_1016,N_309,N_30);
or U1017 (N_1017,N_742,N_373);
nor U1018 (N_1018,N_743,N_314);
and U1019 (N_1019,N_272,N_93);
nand U1020 (N_1020,N_67,N_741);
nand U1021 (N_1021,N_403,N_40);
or U1022 (N_1022,N_316,N_66);
nand U1023 (N_1023,N_567,N_524);
and U1024 (N_1024,N_510,N_328);
nand U1025 (N_1025,N_701,N_514);
nor U1026 (N_1026,N_291,N_325);
or U1027 (N_1027,N_278,N_83);
xor U1028 (N_1028,N_124,N_679);
and U1029 (N_1029,N_597,N_306);
and U1030 (N_1030,N_641,N_562);
and U1031 (N_1031,N_384,N_45);
and U1032 (N_1032,N_171,N_86);
and U1033 (N_1033,N_111,N_4);
nor U1034 (N_1034,N_156,N_243);
nand U1035 (N_1035,N_181,N_116);
or U1036 (N_1036,N_398,N_193);
or U1037 (N_1037,N_601,N_286);
nand U1038 (N_1038,N_552,N_481);
nand U1039 (N_1039,N_551,N_582);
nor U1040 (N_1040,N_331,N_409);
or U1041 (N_1041,N_345,N_37);
nor U1042 (N_1042,N_624,N_280);
and U1043 (N_1043,N_452,N_339);
or U1044 (N_1044,N_106,N_8);
xnor U1045 (N_1045,N_415,N_488);
or U1046 (N_1046,N_203,N_212);
nor U1047 (N_1047,N_74,N_160);
and U1048 (N_1048,N_545,N_223);
nand U1049 (N_1049,N_180,N_463);
nand U1050 (N_1050,N_10,N_397);
nand U1051 (N_1051,N_301,N_720);
nand U1052 (N_1052,N_621,N_442);
nor U1053 (N_1053,N_418,N_395);
and U1054 (N_1054,N_547,N_706);
or U1055 (N_1055,N_632,N_630);
nand U1056 (N_1056,N_7,N_218);
or U1057 (N_1057,N_303,N_628);
or U1058 (N_1058,N_441,N_196);
and U1059 (N_1059,N_493,N_6);
and U1060 (N_1060,N_36,N_512);
nor U1061 (N_1061,N_282,N_178);
nor U1062 (N_1062,N_338,N_201);
and U1063 (N_1063,N_473,N_262);
and U1064 (N_1064,N_149,N_130);
nor U1065 (N_1065,N_119,N_43);
or U1066 (N_1066,N_322,N_285);
nor U1067 (N_1067,N_176,N_500);
or U1068 (N_1068,N_553,N_135);
or U1069 (N_1069,N_287,N_105);
nand U1070 (N_1070,N_396,N_477);
and U1071 (N_1071,N_747,N_663);
nand U1072 (N_1072,N_155,N_114);
xnor U1073 (N_1073,N_598,N_252);
or U1074 (N_1074,N_502,N_28);
nor U1075 (N_1075,N_497,N_704);
nand U1076 (N_1076,N_298,N_53);
nor U1077 (N_1077,N_3,N_268);
nand U1078 (N_1078,N_555,N_525);
xnor U1079 (N_1079,N_370,N_449);
nor U1080 (N_1080,N_341,N_646);
nand U1081 (N_1081,N_330,N_333);
xnor U1082 (N_1082,N_406,N_659);
nor U1083 (N_1083,N_580,N_302);
nand U1084 (N_1084,N_610,N_21);
nor U1085 (N_1085,N_102,N_197);
and U1086 (N_1086,N_508,N_249);
nor U1087 (N_1087,N_651,N_289);
and U1088 (N_1088,N_594,N_478);
or U1089 (N_1089,N_399,N_128);
nand U1090 (N_1090,N_460,N_648);
nand U1091 (N_1091,N_18,N_71);
nor U1092 (N_1092,N_198,N_716);
and U1093 (N_1093,N_645,N_568);
or U1094 (N_1094,N_240,N_702);
nor U1095 (N_1095,N_634,N_266);
or U1096 (N_1096,N_451,N_259);
or U1097 (N_1097,N_576,N_729);
or U1098 (N_1098,N_182,N_41);
nand U1099 (N_1099,N_390,N_99);
nand U1100 (N_1100,N_589,N_108);
and U1101 (N_1101,N_643,N_565);
nand U1102 (N_1102,N_541,N_489);
or U1103 (N_1103,N_387,N_652);
and U1104 (N_1104,N_371,N_313);
and U1105 (N_1105,N_257,N_15);
nand U1106 (N_1106,N_633,N_667);
nand U1107 (N_1107,N_421,N_25);
nand U1108 (N_1108,N_517,N_34);
and U1109 (N_1109,N_389,N_416);
and U1110 (N_1110,N_563,N_467);
or U1111 (N_1111,N_691,N_139);
or U1112 (N_1112,N_19,N_138);
and U1113 (N_1113,N_143,N_606);
nand U1114 (N_1114,N_498,N_684);
nand U1115 (N_1115,N_516,N_192);
or U1116 (N_1116,N_721,N_486);
nand U1117 (N_1117,N_434,N_273);
or U1118 (N_1118,N_653,N_609);
nor U1119 (N_1119,N_575,N_655);
nand U1120 (N_1120,N_235,N_417);
and U1121 (N_1121,N_364,N_427);
nand U1122 (N_1122,N_483,N_686);
and U1123 (N_1123,N_685,N_422);
or U1124 (N_1124,N_343,N_136);
nor U1125 (N_1125,N_587,N_450);
nand U1126 (N_1126,N_124,N_511);
or U1127 (N_1127,N_205,N_85);
nor U1128 (N_1128,N_400,N_536);
nor U1129 (N_1129,N_120,N_123);
nor U1130 (N_1130,N_682,N_103);
xor U1131 (N_1131,N_740,N_733);
or U1132 (N_1132,N_105,N_23);
or U1133 (N_1133,N_149,N_141);
or U1134 (N_1134,N_307,N_521);
nor U1135 (N_1135,N_331,N_257);
or U1136 (N_1136,N_547,N_163);
nand U1137 (N_1137,N_692,N_238);
or U1138 (N_1138,N_657,N_64);
or U1139 (N_1139,N_173,N_635);
nand U1140 (N_1140,N_167,N_281);
or U1141 (N_1141,N_454,N_9);
or U1142 (N_1142,N_10,N_670);
nand U1143 (N_1143,N_513,N_667);
or U1144 (N_1144,N_735,N_657);
nor U1145 (N_1145,N_556,N_148);
or U1146 (N_1146,N_224,N_654);
or U1147 (N_1147,N_168,N_505);
and U1148 (N_1148,N_747,N_156);
and U1149 (N_1149,N_425,N_746);
and U1150 (N_1150,N_376,N_496);
nor U1151 (N_1151,N_271,N_526);
and U1152 (N_1152,N_353,N_179);
or U1153 (N_1153,N_385,N_678);
nor U1154 (N_1154,N_177,N_381);
and U1155 (N_1155,N_555,N_598);
nor U1156 (N_1156,N_240,N_523);
or U1157 (N_1157,N_79,N_95);
and U1158 (N_1158,N_387,N_235);
nand U1159 (N_1159,N_584,N_568);
nor U1160 (N_1160,N_328,N_690);
and U1161 (N_1161,N_194,N_240);
or U1162 (N_1162,N_198,N_356);
nand U1163 (N_1163,N_225,N_159);
nand U1164 (N_1164,N_596,N_694);
nor U1165 (N_1165,N_227,N_502);
nand U1166 (N_1166,N_110,N_419);
nand U1167 (N_1167,N_250,N_137);
nor U1168 (N_1168,N_583,N_579);
nor U1169 (N_1169,N_436,N_465);
nand U1170 (N_1170,N_472,N_498);
nor U1171 (N_1171,N_95,N_450);
nor U1172 (N_1172,N_290,N_286);
and U1173 (N_1173,N_736,N_160);
nor U1174 (N_1174,N_661,N_383);
nor U1175 (N_1175,N_155,N_284);
nand U1176 (N_1176,N_413,N_185);
and U1177 (N_1177,N_675,N_449);
nor U1178 (N_1178,N_263,N_540);
nand U1179 (N_1179,N_537,N_605);
and U1180 (N_1180,N_504,N_60);
and U1181 (N_1181,N_582,N_536);
and U1182 (N_1182,N_708,N_287);
nand U1183 (N_1183,N_503,N_182);
nor U1184 (N_1184,N_288,N_150);
or U1185 (N_1185,N_11,N_99);
or U1186 (N_1186,N_138,N_588);
nor U1187 (N_1187,N_496,N_116);
nand U1188 (N_1188,N_419,N_632);
and U1189 (N_1189,N_338,N_73);
or U1190 (N_1190,N_313,N_546);
nor U1191 (N_1191,N_327,N_165);
or U1192 (N_1192,N_430,N_115);
or U1193 (N_1193,N_582,N_721);
or U1194 (N_1194,N_312,N_472);
or U1195 (N_1195,N_170,N_320);
or U1196 (N_1196,N_471,N_312);
nand U1197 (N_1197,N_521,N_679);
and U1198 (N_1198,N_631,N_382);
nor U1199 (N_1199,N_443,N_606);
or U1200 (N_1200,N_203,N_300);
or U1201 (N_1201,N_306,N_496);
and U1202 (N_1202,N_53,N_44);
nor U1203 (N_1203,N_487,N_525);
nand U1204 (N_1204,N_171,N_147);
nand U1205 (N_1205,N_737,N_459);
nor U1206 (N_1206,N_80,N_366);
or U1207 (N_1207,N_410,N_547);
nand U1208 (N_1208,N_497,N_701);
or U1209 (N_1209,N_523,N_704);
nor U1210 (N_1210,N_107,N_412);
and U1211 (N_1211,N_409,N_26);
nand U1212 (N_1212,N_240,N_147);
nor U1213 (N_1213,N_748,N_187);
nand U1214 (N_1214,N_408,N_97);
nor U1215 (N_1215,N_749,N_528);
or U1216 (N_1216,N_559,N_29);
nor U1217 (N_1217,N_345,N_235);
and U1218 (N_1218,N_147,N_717);
or U1219 (N_1219,N_331,N_212);
or U1220 (N_1220,N_663,N_592);
or U1221 (N_1221,N_661,N_165);
or U1222 (N_1222,N_200,N_504);
nand U1223 (N_1223,N_346,N_471);
nor U1224 (N_1224,N_193,N_515);
or U1225 (N_1225,N_411,N_365);
nor U1226 (N_1226,N_190,N_378);
nor U1227 (N_1227,N_337,N_1);
and U1228 (N_1228,N_340,N_599);
or U1229 (N_1229,N_585,N_55);
and U1230 (N_1230,N_560,N_339);
nor U1231 (N_1231,N_107,N_249);
nand U1232 (N_1232,N_501,N_256);
nor U1233 (N_1233,N_559,N_331);
or U1234 (N_1234,N_492,N_294);
nand U1235 (N_1235,N_593,N_740);
nand U1236 (N_1236,N_305,N_534);
or U1237 (N_1237,N_214,N_77);
nor U1238 (N_1238,N_223,N_617);
nor U1239 (N_1239,N_54,N_173);
nor U1240 (N_1240,N_251,N_6);
and U1241 (N_1241,N_267,N_447);
and U1242 (N_1242,N_326,N_250);
nor U1243 (N_1243,N_101,N_745);
or U1244 (N_1244,N_2,N_219);
and U1245 (N_1245,N_361,N_663);
or U1246 (N_1246,N_686,N_744);
nand U1247 (N_1247,N_674,N_463);
or U1248 (N_1248,N_397,N_160);
or U1249 (N_1249,N_326,N_219);
and U1250 (N_1250,N_415,N_476);
and U1251 (N_1251,N_569,N_637);
nand U1252 (N_1252,N_133,N_630);
and U1253 (N_1253,N_153,N_702);
nand U1254 (N_1254,N_112,N_349);
or U1255 (N_1255,N_396,N_124);
nand U1256 (N_1256,N_454,N_188);
nand U1257 (N_1257,N_331,N_58);
nor U1258 (N_1258,N_272,N_281);
nor U1259 (N_1259,N_518,N_585);
nand U1260 (N_1260,N_31,N_395);
nand U1261 (N_1261,N_673,N_400);
nand U1262 (N_1262,N_618,N_685);
and U1263 (N_1263,N_319,N_347);
and U1264 (N_1264,N_63,N_385);
or U1265 (N_1265,N_380,N_206);
nand U1266 (N_1266,N_612,N_568);
nor U1267 (N_1267,N_512,N_72);
or U1268 (N_1268,N_579,N_611);
or U1269 (N_1269,N_604,N_649);
nand U1270 (N_1270,N_342,N_314);
and U1271 (N_1271,N_226,N_520);
and U1272 (N_1272,N_471,N_216);
nand U1273 (N_1273,N_108,N_12);
nor U1274 (N_1274,N_10,N_726);
nand U1275 (N_1275,N_485,N_212);
or U1276 (N_1276,N_737,N_348);
nor U1277 (N_1277,N_738,N_696);
and U1278 (N_1278,N_438,N_182);
and U1279 (N_1279,N_500,N_565);
and U1280 (N_1280,N_643,N_488);
nor U1281 (N_1281,N_299,N_632);
or U1282 (N_1282,N_6,N_694);
and U1283 (N_1283,N_117,N_555);
nor U1284 (N_1284,N_679,N_119);
or U1285 (N_1285,N_560,N_507);
nand U1286 (N_1286,N_267,N_732);
or U1287 (N_1287,N_113,N_371);
and U1288 (N_1288,N_211,N_615);
and U1289 (N_1289,N_577,N_325);
nor U1290 (N_1290,N_171,N_564);
or U1291 (N_1291,N_217,N_36);
and U1292 (N_1292,N_201,N_676);
and U1293 (N_1293,N_529,N_192);
or U1294 (N_1294,N_490,N_382);
or U1295 (N_1295,N_552,N_374);
nand U1296 (N_1296,N_673,N_393);
nand U1297 (N_1297,N_715,N_717);
nor U1298 (N_1298,N_185,N_444);
nor U1299 (N_1299,N_464,N_281);
and U1300 (N_1300,N_94,N_674);
or U1301 (N_1301,N_206,N_739);
and U1302 (N_1302,N_745,N_409);
and U1303 (N_1303,N_377,N_522);
nor U1304 (N_1304,N_39,N_375);
or U1305 (N_1305,N_154,N_446);
nand U1306 (N_1306,N_541,N_198);
and U1307 (N_1307,N_2,N_163);
nor U1308 (N_1308,N_486,N_633);
xnor U1309 (N_1309,N_339,N_17);
and U1310 (N_1310,N_267,N_130);
nand U1311 (N_1311,N_522,N_299);
nand U1312 (N_1312,N_219,N_407);
nand U1313 (N_1313,N_478,N_391);
nor U1314 (N_1314,N_82,N_533);
or U1315 (N_1315,N_599,N_196);
nor U1316 (N_1316,N_197,N_552);
and U1317 (N_1317,N_554,N_186);
or U1318 (N_1318,N_566,N_314);
or U1319 (N_1319,N_444,N_740);
nand U1320 (N_1320,N_328,N_273);
and U1321 (N_1321,N_637,N_428);
and U1322 (N_1322,N_497,N_379);
nor U1323 (N_1323,N_240,N_579);
nor U1324 (N_1324,N_98,N_548);
and U1325 (N_1325,N_65,N_122);
nand U1326 (N_1326,N_270,N_379);
nor U1327 (N_1327,N_80,N_482);
and U1328 (N_1328,N_83,N_125);
nor U1329 (N_1329,N_47,N_116);
and U1330 (N_1330,N_299,N_531);
nor U1331 (N_1331,N_708,N_294);
nor U1332 (N_1332,N_556,N_672);
or U1333 (N_1333,N_666,N_242);
nand U1334 (N_1334,N_679,N_401);
and U1335 (N_1335,N_183,N_110);
nor U1336 (N_1336,N_743,N_354);
and U1337 (N_1337,N_679,N_716);
and U1338 (N_1338,N_370,N_445);
and U1339 (N_1339,N_115,N_432);
nor U1340 (N_1340,N_526,N_683);
and U1341 (N_1341,N_118,N_318);
nand U1342 (N_1342,N_181,N_493);
and U1343 (N_1343,N_114,N_274);
or U1344 (N_1344,N_574,N_652);
nor U1345 (N_1345,N_212,N_168);
nand U1346 (N_1346,N_669,N_219);
nor U1347 (N_1347,N_654,N_720);
nand U1348 (N_1348,N_149,N_551);
xor U1349 (N_1349,N_443,N_235);
and U1350 (N_1350,N_657,N_326);
nor U1351 (N_1351,N_538,N_617);
nand U1352 (N_1352,N_678,N_17);
and U1353 (N_1353,N_29,N_60);
and U1354 (N_1354,N_350,N_266);
nor U1355 (N_1355,N_101,N_329);
nand U1356 (N_1356,N_576,N_20);
and U1357 (N_1357,N_722,N_66);
nand U1358 (N_1358,N_272,N_412);
nor U1359 (N_1359,N_86,N_359);
nand U1360 (N_1360,N_459,N_242);
nand U1361 (N_1361,N_83,N_436);
or U1362 (N_1362,N_501,N_7);
and U1363 (N_1363,N_0,N_274);
or U1364 (N_1364,N_589,N_220);
or U1365 (N_1365,N_33,N_149);
or U1366 (N_1366,N_452,N_396);
nand U1367 (N_1367,N_90,N_33);
nand U1368 (N_1368,N_28,N_31);
and U1369 (N_1369,N_404,N_427);
or U1370 (N_1370,N_500,N_18);
or U1371 (N_1371,N_440,N_373);
nand U1372 (N_1372,N_671,N_122);
or U1373 (N_1373,N_719,N_541);
or U1374 (N_1374,N_715,N_151);
nor U1375 (N_1375,N_590,N_252);
or U1376 (N_1376,N_26,N_290);
nand U1377 (N_1377,N_361,N_257);
nor U1378 (N_1378,N_443,N_121);
nor U1379 (N_1379,N_287,N_572);
nand U1380 (N_1380,N_376,N_147);
or U1381 (N_1381,N_589,N_97);
nor U1382 (N_1382,N_187,N_473);
nand U1383 (N_1383,N_690,N_559);
nand U1384 (N_1384,N_330,N_577);
and U1385 (N_1385,N_123,N_446);
or U1386 (N_1386,N_61,N_631);
nor U1387 (N_1387,N_149,N_525);
nor U1388 (N_1388,N_584,N_686);
and U1389 (N_1389,N_495,N_29);
nor U1390 (N_1390,N_146,N_570);
nand U1391 (N_1391,N_223,N_485);
nand U1392 (N_1392,N_94,N_327);
nand U1393 (N_1393,N_747,N_403);
nand U1394 (N_1394,N_107,N_277);
nor U1395 (N_1395,N_110,N_451);
nor U1396 (N_1396,N_472,N_553);
and U1397 (N_1397,N_430,N_597);
and U1398 (N_1398,N_120,N_204);
and U1399 (N_1399,N_493,N_145);
or U1400 (N_1400,N_95,N_218);
nand U1401 (N_1401,N_383,N_624);
or U1402 (N_1402,N_92,N_496);
nor U1403 (N_1403,N_138,N_366);
nand U1404 (N_1404,N_92,N_342);
and U1405 (N_1405,N_574,N_531);
or U1406 (N_1406,N_91,N_316);
nand U1407 (N_1407,N_327,N_204);
nor U1408 (N_1408,N_124,N_459);
or U1409 (N_1409,N_243,N_317);
or U1410 (N_1410,N_95,N_688);
and U1411 (N_1411,N_177,N_487);
nand U1412 (N_1412,N_65,N_4);
nor U1413 (N_1413,N_122,N_276);
nor U1414 (N_1414,N_399,N_50);
or U1415 (N_1415,N_93,N_23);
and U1416 (N_1416,N_436,N_641);
and U1417 (N_1417,N_620,N_339);
or U1418 (N_1418,N_574,N_82);
nand U1419 (N_1419,N_335,N_714);
and U1420 (N_1420,N_647,N_217);
xor U1421 (N_1421,N_442,N_90);
and U1422 (N_1422,N_12,N_456);
nor U1423 (N_1423,N_631,N_245);
or U1424 (N_1424,N_485,N_748);
and U1425 (N_1425,N_537,N_528);
or U1426 (N_1426,N_269,N_40);
xor U1427 (N_1427,N_307,N_331);
nand U1428 (N_1428,N_48,N_357);
and U1429 (N_1429,N_555,N_645);
nor U1430 (N_1430,N_163,N_715);
and U1431 (N_1431,N_584,N_720);
or U1432 (N_1432,N_586,N_20);
nor U1433 (N_1433,N_59,N_507);
nor U1434 (N_1434,N_616,N_39);
nand U1435 (N_1435,N_9,N_284);
nand U1436 (N_1436,N_33,N_612);
xnor U1437 (N_1437,N_129,N_147);
or U1438 (N_1438,N_388,N_632);
nor U1439 (N_1439,N_720,N_180);
nor U1440 (N_1440,N_127,N_266);
and U1441 (N_1441,N_643,N_8);
nor U1442 (N_1442,N_624,N_50);
nor U1443 (N_1443,N_189,N_327);
and U1444 (N_1444,N_634,N_521);
or U1445 (N_1445,N_656,N_493);
and U1446 (N_1446,N_404,N_718);
or U1447 (N_1447,N_191,N_55);
and U1448 (N_1448,N_188,N_442);
and U1449 (N_1449,N_740,N_641);
nor U1450 (N_1450,N_430,N_498);
and U1451 (N_1451,N_384,N_75);
nand U1452 (N_1452,N_228,N_720);
nand U1453 (N_1453,N_712,N_242);
nand U1454 (N_1454,N_445,N_694);
or U1455 (N_1455,N_377,N_97);
nor U1456 (N_1456,N_334,N_128);
or U1457 (N_1457,N_7,N_516);
nand U1458 (N_1458,N_401,N_374);
or U1459 (N_1459,N_401,N_392);
nand U1460 (N_1460,N_339,N_192);
xnor U1461 (N_1461,N_357,N_563);
nor U1462 (N_1462,N_167,N_435);
nor U1463 (N_1463,N_603,N_211);
nor U1464 (N_1464,N_727,N_254);
nor U1465 (N_1465,N_60,N_744);
or U1466 (N_1466,N_300,N_473);
or U1467 (N_1467,N_324,N_317);
and U1468 (N_1468,N_128,N_148);
nand U1469 (N_1469,N_185,N_36);
nor U1470 (N_1470,N_277,N_713);
nand U1471 (N_1471,N_538,N_129);
or U1472 (N_1472,N_264,N_688);
or U1473 (N_1473,N_299,N_87);
and U1474 (N_1474,N_37,N_568);
nand U1475 (N_1475,N_530,N_439);
and U1476 (N_1476,N_99,N_48);
and U1477 (N_1477,N_587,N_204);
nor U1478 (N_1478,N_691,N_1);
and U1479 (N_1479,N_603,N_126);
and U1480 (N_1480,N_507,N_153);
nor U1481 (N_1481,N_106,N_86);
nand U1482 (N_1482,N_297,N_707);
and U1483 (N_1483,N_75,N_624);
nand U1484 (N_1484,N_107,N_475);
or U1485 (N_1485,N_161,N_151);
and U1486 (N_1486,N_293,N_300);
nor U1487 (N_1487,N_602,N_12);
nor U1488 (N_1488,N_401,N_434);
nand U1489 (N_1489,N_500,N_364);
nand U1490 (N_1490,N_441,N_359);
and U1491 (N_1491,N_515,N_89);
or U1492 (N_1492,N_315,N_90);
nor U1493 (N_1493,N_15,N_74);
or U1494 (N_1494,N_749,N_122);
nand U1495 (N_1495,N_368,N_495);
or U1496 (N_1496,N_71,N_465);
nand U1497 (N_1497,N_539,N_58);
or U1498 (N_1498,N_571,N_418);
or U1499 (N_1499,N_191,N_731);
nor U1500 (N_1500,N_1345,N_935);
nor U1501 (N_1501,N_1052,N_817);
nand U1502 (N_1502,N_836,N_909);
nand U1503 (N_1503,N_756,N_1471);
or U1504 (N_1504,N_1374,N_1140);
or U1505 (N_1505,N_1199,N_785);
and U1506 (N_1506,N_1108,N_1128);
or U1507 (N_1507,N_1184,N_758);
and U1508 (N_1508,N_1430,N_1318);
nor U1509 (N_1509,N_1103,N_1284);
or U1510 (N_1510,N_779,N_846);
and U1511 (N_1511,N_1141,N_1458);
nor U1512 (N_1512,N_1372,N_907);
and U1513 (N_1513,N_1170,N_1124);
and U1514 (N_1514,N_976,N_1083);
nand U1515 (N_1515,N_1319,N_1278);
nor U1516 (N_1516,N_787,N_1195);
and U1517 (N_1517,N_1036,N_816);
nor U1518 (N_1518,N_1415,N_904);
nor U1519 (N_1519,N_1177,N_1260);
and U1520 (N_1520,N_1325,N_1234);
or U1521 (N_1521,N_1071,N_1077);
or U1522 (N_1522,N_1256,N_1365);
and U1523 (N_1523,N_1157,N_979);
nand U1524 (N_1524,N_793,N_1439);
nand U1525 (N_1525,N_1009,N_1338);
nor U1526 (N_1526,N_1019,N_1204);
and U1527 (N_1527,N_1292,N_1249);
nand U1528 (N_1528,N_1223,N_1159);
nor U1529 (N_1529,N_1344,N_1106);
or U1530 (N_1530,N_1064,N_1237);
nand U1531 (N_1531,N_777,N_1239);
or U1532 (N_1532,N_1253,N_802);
or U1533 (N_1533,N_853,N_900);
nand U1534 (N_1534,N_1307,N_1397);
nor U1535 (N_1535,N_1030,N_1333);
and U1536 (N_1536,N_1401,N_1163);
and U1537 (N_1537,N_1025,N_989);
nand U1538 (N_1538,N_828,N_1169);
nand U1539 (N_1539,N_1181,N_1480);
or U1540 (N_1540,N_1355,N_1228);
nand U1541 (N_1541,N_1472,N_1102);
or U1542 (N_1542,N_1012,N_1148);
nand U1543 (N_1543,N_1015,N_1217);
nand U1544 (N_1544,N_962,N_1363);
nor U1545 (N_1545,N_1109,N_869);
or U1546 (N_1546,N_780,N_937);
nand U1547 (N_1547,N_1155,N_1214);
nand U1548 (N_1548,N_1351,N_1436);
and U1549 (N_1549,N_913,N_1481);
or U1550 (N_1550,N_1117,N_1118);
nor U1551 (N_1551,N_1194,N_774);
and U1552 (N_1552,N_1297,N_1346);
and U1553 (N_1553,N_923,N_1306);
nor U1554 (N_1554,N_868,N_1000);
nor U1555 (N_1555,N_1440,N_1242);
nand U1556 (N_1556,N_1287,N_951);
nor U1557 (N_1557,N_812,N_903);
nor U1558 (N_1558,N_1488,N_1271);
and U1559 (N_1559,N_1200,N_965);
or U1560 (N_1560,N_983,N_1267);
or U1561 (N_1561,N_1315,N_1136);
and U1562 (N_1562,N_1396,N_1087);
nor U1563 (N_1563,N_1298,N_1266);
nor U1564 (N_1564,N_1100,N_1144);
and U1565 (N_1565,N_805,N_1011);
nand U1566 (N_1566,N_838,N_1206);
nor U1567 (N_1567,N_1469,N_1347);
nor U1568 (N_1568,N_1336,N_1384);
nand U1569 (N_1569,N_1288,N_768);
nor U1570 (N_1570,N_1153,N_1165);
or U1571 (N_1571,N_1069,N_752);
and U1572 (N_1572,N_1388,N_1129);
nor U1573 (N_1573,N_1489,N_1038);
nor U1574 (N_1574,N_860,N_1186);
or U1575 (N_1575,N_1008,N_1014);
or U1576 (N_1576,N_924,N_1245);
nand U1577 (N_1577,N_1201,N_1020);
or U1578 (N_1578,N_1092,N_1142);
nand U1579 (N_1579,N_893,N_1276);
nor U1580 (N_1580,N_1322,N_792);
and U1581 (N_1581,N_1189,N_1460);
and U1582 (N_1582,N_769,N_1431);
nand U1583 (N_1583,N_1273,N_1004);
and U1584 (N_1584,N_1235,N_1107);
or U1585 (N_1585,N_1205,N_1497);
nor U1586 (N_1586,N_1252,N_906);
and U1587 (N_1587,N_920,N_798);
nand U1588 (N_1588,N_1167,N_799);
and U1589 (N_1589,N_931,N_1045);
nand U1590 (N_1590,N_1173,N_1392);
and U1591 (N_1591,N_1358,N_784);
or U1592 (N_1592,N_1050,N_1437);
and U1593 (N_1593,N_808,N_1243);
nand U1594 (N_1594,N_1134,N_761);
nor U1595 (N_1595,N_1127,N_1393);
nand U1596 (N_1596,N_936,N_1022);
nand U1597 (N_1597,N_1147,N_1326);
or U1598 (N_1598,N_940,N_1323);
nand U1599 (N_1599,N_1085,N_1058);
nor U1600 (N_1600,N_1139,N_964);
nand U1601 (N_1601,N_1312,N_946);
and U1602 (N_1602,N_1411,N_804);
nor U1603 (N_1603,N_1099,N_894);
nand U1604 (N_1604,N_1031,N_783);
nand U1605 (N_1605,N_1265,N_1233);
nand U1606 (N_1606,N_1041,N_1224);
nor U1607 (N_1607,N_1465,N_885);
nand U1608 (N_1608,N_824,N_1427);
and U1609 (N_1609,N_794,N_810);
or U1610 (N_1610,N_1185,N_1027);
nor U1611 (N_1611,N_944,N_1227);
and U1612 (N_1612,N_835,N_760);
or U1613 (N_1613,N_974,N_1407);
nor U1614 (N_1614,N_973,N_1080);
or U1615 (N_1615,N_1434,N_1280);
or U1616 (N_1616,N_753,N_1176);
or U1617 (N_1617,N_864,N_1274);
nor U1618 (N_1618,N_1482,N_1309);
and U1619 (N_1619,N_1328,N_1037);
or U1620 (N_1620,N_925,N_895);
or U1621 (N_1621,N_1091,N_1360);
nor U1622 (N_1622,N_1275,N_1335);
nand U1623 (N_1623,N_1453,N_1414);
nand U1624 (N_1624,N_1054,N_1123);
nor U1625 (N_1625,N_1409,N_1003);
nand U1626 (N_1626,N_1111,N_1382);
nand U1627 (N_1627,N_1316,N_754);
or U1628 (N_1628,N_1295,N_1076);
nand U1629 (N_1629,N_1244,N_781);
nor U1630 (N_1630,N_873,N_1192);
or U1631 (N_1631,N_1479,N_1188);
and U1632 (N_1632,N_1162,N_899);
nand U1633 (N_1633,N_1493,N_987);
nor U1634 (N_1634,N_806,N_1420);
xnor U1635 (N_1635,N_1332,N_1090);
and U1636 (N_1636,N_999,N_902);
nand U1637 (N_1637,N_1405,N_1166);
and U1638 (N_1638,N_1079,N_1476);
nand U1639 (N_1639,N_1208,N_1095);
nand U1640 (N_1640,N_992,N_1241);
and U1641 (N_1641,N_1313,N_1218);
nand U1642 (N_1642,N_763,N_1135);
or U1643 (N_1643,N_1101,N_874);
nand U1644 (N_1644,N_1018,N_782);
and U1645 (N_1645,N_1310,N_1051);
nand U1646 (N_1646,N_850,N_826);
nand U1647 (N_1647,N_1468,N_1408);
or U1648 (N_1648,N_1435,N_1272);
nor U1649 (N_1649,N_1448,N_872);
xor U1650 (N_1650,N_1057,N_1289);
nor U1651 (N_1651,N_1219,N_911);
nand U1652 (N_1652,N_773,N_790);
nand U1653 (N_1653,N_856,N_1403);
nand U1654 (N_1654,N_1340,N_910);
nor U1655 (N_1655,N_1178,N_1417);
and U1656 (N_1656,N_1475,N_1362);
nand U1657 (N_1657,N_1389,N_1290);
nor U1658 (N_1658,N_982,N_859);
nand U1659 (N_1659,N_1246,N_916);
and U1660 (N_1660,N_1121,N_1105);
xor U1661 (N_1661,N_1073,N_1391);
and U1662 (N_1662,N_1492,N_1232);
and U1663 (N_1663,N_1158,N_1028);
and U1664 (N_1664,N_1423,N_852);
xor U1665 (N_1665,N_1098,N_1291);
nand U1666 (N_1666,N_918,N_994);
nand U1667 (N_1667,N_919,N_829);
nor U1668 (N_1668,N_1317,N_933);
or U1669 (N_1669,N_1477,N_975);
and U1670 (N_1670,N_847,N_1151);
nor U1671 (N_1671,N_905,N_1089);
nor U1672 (N_1672,N_786,N_1305);
or U1673 (N_1673,N_1063,N_1464);
nand U1674 (N_1674,N_797,N_915);
nor U1675 (N_1675,N_938,N_1293);
and U1676 (N_1676,N_834,N_827);
or U1677 (N_1677,N_966,N_1207);
nor U1678 (N_1678,N_821,N_1226);
nand U1679 (N_1679,N_803,N_1327);
nor U1680 (N_1680,N_917,N_1251);
nand U1681 (N_1681,N_1418,N_1255);
nor U1682 (N_1682,N_1161,N_922);
and U1683 (N_1683,N_1324,N_1197);
nor U1684 (N_1684,N_1211,N_1075);
and U1685 (N_1685,N_1386,N_875);
or U1686 (N_1686,N_952,N_985);
or U1687 (N_1687,N_1277,N_1074);
or U1688 (N_1688,N_1442,N_912);
nor U1689 (N_1689,N_1032,N_1441);
nand U1690 (N_1690,N_1138,N_958);
nor U1691 (N_1691,N_823,N_1164);
and U1692 (N_1692,N_908,N_1122);
and U1693 (N_1693,N_948,N_809);
nor U1694 (N_1694,N_1149,N_1380);
and U1695 (N_1695,N_1196,N_957);
nor U1696 (N_1696,N_1329,N_815);
or U1697 (N_1697,N_1096,N_800);
and U1698 (N_1698,N_883,N_825);
nand U1699 (N_1699,N_884,N_879);
or U1700 (N_1700,N_861,N_819);
and U1701 (N_1701,N_1115,N_1330);
nor U1702 (N_1702,N_1250,N_1056);
nor U1703 (N_1703,N_1299,N_766);
and U1704 (N_1704,N_841,N_791);
and U1705 (N_1705,N_1466,N_1433);
nor U1706 (N_1706,N_1131,N_1044);
or U1707 (N_1707,N_1404,N_1093);
and U1708 (N_1708,N_1387,N_870);
or U1709 (N_1709,N_1203,N_1042);
or U1710 (N_1710,N_1390,N_1007);
and U1711 (N_1711,N_914,N_1210);
nor U1712 (N_1712,N_1168,N_887);
and U1713 (N_1713,N_1449,N_1160);
nand U1714 (N_1714,N_789,N_1446);
and U1715 (N_1715,N_881,N_839);
or U1716 (N_1716,N_959,N_1094);
nand U1717 (N_1717,N_1416,N_1156);
and U1718 (N_1718,N_943,N_1447);
nor U1719 (N_1719,N_837,N_941);
or U1720 (N_1720,N_770,N_1356);
or U1721 (N_1721,N_954,N_1248);
nand U1722 (N_1722,N_1321,N_1478);
and U1723 (N_1723,N_1212,N_993);
and U1724 (N_1724,N_942,N_1375);
nor U1725 (N_1725,N_1357,N_1238);
nor U1726 (N_1726,N_857,N_765);
nand U1727 (N_1727,N_1183,N_1498);
or U1728 (N_1728,N_1078,N_1331);
nor U1729 (N_1729,N_1279,N_1342);
or U1730 (N_1730,N_1114,N_1254);
nand U1731 (N_1731,N_1450,N_848);
and U1732 (N_1732,N_1366,N_1146);
and U1733 (N_1733,N_1231,N_788);
or U1734 (N_1734,N_795,N_778);
and U1735 (N_1735,N_833,N_1270);
nor U1736 (N_1736,N_867,N_1132);
nand U1737 (N_1737,N_929,N_851);
or U1738 (N_1738,N_1373,N_1432);
or U1739 (N_1739,N_1002,N_1283);
and U1740 (N_1740,N_1145,N_1048);
nand U1741 (N_1741,N_1303,N_997);
or U1742 (N_1742,N_984,N_926);
and U1743 (N_1743,N_1024,N_876);
or U1744 (N_1744,N_772,N_1359);
or U1745 (N_1745,N_1062,N_1443);
or U1746 (N_1746,N_1496,N_969);
nand U1747 (N_1747,N_1171,N_1172);
and U1748 (N_1748,N_1339,N_1486);
nor U1749 (N_1749,N_1422,N_1154);
and U1750 (N_1750,N_1017,N_820);
nor U1751 (N_1751,N_1296,N_968);
or U1752 (N_1752,N_934,N_1059);
or U1753 (N_1753,N_807,N_1463);
nand U1754 (N_1754,N_1383,N_759);
nand U1755 (N_1755,N_840,N_1459);
nand U1756 (N_1756,N_1053,N_1072);
nand U1757 (N_1757,N_1484,N_1070);
and U1758 (N_1758,N_1229,N_1143);
or U1759 (N_1759,N_1398,N_1308);
nand U1760 (N_1760,N_1371,N_1110);
nand U1761 (N_1761,N_855,N_1180);
nor U1762 (N_1762,N_1043,N_882);
and U1763 (N_1763,N_1126,N_1381);
nor U1764 (N_1764,N_1467,N_1055);
and U1765 (N_1765,N_921,N_956);
or U1766 (N_1766,N_1113,N_1282);
or U1767 (N_1767,N_822,N_1258);
and U1768 (N_1768,N_928,N_1301);
nand U1769 (N_1769,N_1474,N_1419);
and U1770 (N_1770,N_1485,N_1368);
and U1771 (N_1771,N_751,N_1361);
or U1772 (N_1772,N_949,N_1320);
nand U1773 (N_1773,N_967,N_1262);
nor U1774 (N_1774,N_1236,N_1084);
nand U1775 (N_1775,N_1202,N_898);
nand U1776 (N_1776,N_901,N_1395);
nor U1777 (N_1777,N_1425,N_814);
nand U1778 (N_1778,N_1349,N_897);
and U1779 (N_1779,N_1445,N_1152);
nand U1780 (N_1780,N_862,N_1081);
nor U1781 (N_1781,N_877,N_1193);
nor U1782 (N_1782,N_932,N_991);
and U1783 (N_1783,N_947,N_1334);
nor U1784 (N_1784,N_1379,N_1175);
and U1785 (N_1785,N_977,N_1259);
and U1786 (N_1786,N_1046,N_1005);
nor U1787 (N_1787,N_1263,N_1473);
nand U1788 (N_1788,N_762,N_1490);
nor U1789 (N_1789,N_831,N_1350);
nor U1790 (N_1790,N_1230,N_1499);
and U1791 (N_1791,N_1487,N_1029);
and U1792 (N_1792,N_1120,N_801);
or U1793 (N_1793,N_1494,N_1086);
or U1794 (N_1794,N_1285,N_1454);
nand U1795 (N_1795,N_1268,N_1444);
or U1796 (N_1796,N_1191,N_886);
nand U1797 (N_1797,N_1426,N_978);
or U1798 (N_1798,N_1049,N_981);
and U1799 (N_1799,N_843,N_1377);
or U1800 (N_1800,N_858,N_980);
and U1801 (N_1801,N_950,N_1209);
nor U1802 (N_1802,N_890,N_960);
nand U1803 (N_1803,N_871,N_889);
nor U1804 (N_1804,N_1341,N_1410);
and U1805 (N_1805,N_1491,N_1026);
nor U1806 (N_1806,N_1040,N_1001);
and U1807 (N_1807,N_1137,N_1213);
nor U1808 (N_1808,N_955,N_757);
or U1809 (N_1809,N_1179,N_1006);
nor U1810 (N_1810,N_1424,N_1104);
nor U1811 (N_1811,N_1457,N_945);
and U1812 (N_1812,N_1462,N_1065);
and U1813 (N_1813,N_1399,N_1337);
nand U1814 (N_1814,N_1378,N_927);
or U1815 (N_1815,N_995,N_1311);
or U1816 (N_1816,N_1385,N_1455);
and U1817 (N_1817,N_880,N_1034);
and U1818 (N_1818,N_1016,N_1281);
or U1819 (N_1819,N_842,N_1352);
nor U1820 (N_1820,N_1215,N_1394);
nor U1821 (N_1821,N_1033,N_845);
nand U1822 (N_1822,N_1456,N_1364);
and U1823 (N_1823,N_1343,N_1294);
and U1824 (N_1824,N_832,N_811);
nor U1825 (N_1825,N_775,N_771);
and U1826 (N_1826,N_1221,N_866);
nor U1827 (N_1827,N_888,N_1369);
and U1828 (N_1828,N_764,N_1021);
or U1829 (N_1829,N_1483,N_939);
nand U1830 (N_1830,N_1216,N_1068);
and U1831 (N_1831,N_1082,N_878);
or U1832 (N_1832,N_1348,N_1300);
or U1833 (N_1833,N_1067,N_891);
or U1834 (N_1834,N_755,N_1406);
or U1835 (N_1835,N_972,N_1367);
nand U1836 (N_1836,N_1412,N_1198);
nand U1837 (N_1837,N_1257,N_849);
and U1838 (N_1838,N_1428,N_988);
nand U1839 (N_1839,N_1269,N_1222);
nor U1840 (N_1840,N_1190,N_963);
or U1841 (N_1841,N_1039,N_970);
nor U1842 (N_1842,N_1066,N_1220);
and U1843 (N_1843,N_1354,N_1182);
nor U1844 (N_1844,N_896,N_961);
and U1845 (N_1845,N_1130,N_1495);
nand U1846 (N_1846,N_1023,N_1088);
or U1847 (N_1847,N_990,N_796);
or U1848 (N_1848,N_1451,N_1060);
or U1849 (N_1849,N_1187,N_750);
nand U1850 (N_1850,N_1302,N_1314);
nor U1851 (N_1851,N_1116,N_1264);
and U1852 (N_1852,N_863,N_1240);
and U1853 (N_1853,N_1370,N_1452);
or U1854 (N_1854,N_1247,N_854);
and U1855 (N_1855,N_1286,N_971);
and U1856 (N_1856,N_1150,N_830);
and U1857 (N_1857,N_1353,N_1470);
nand U1858 (N_1858,N_953,N_1010);
or U1859 (N_1859,N_1304,N_998);
nand U1860 (N_1860,N_1376,N_776);
nor U1861 (N_1861,N_1119,N_892);
nor U1862 (N_1862,N_1225,N_813);
nor U1863 (N_1863,N_1097,N_1013);
or U1864 (N_1864,N_1438,N_1174);
or U1865 (N_1865,N_767,N_1061);
nand U1866 (N_1866,N_1261,N_1429);
or U1867 (N_1867,N_1035,N_1112);
nor U1868 (N_1868,N_1133,N_1461);
nor U1869 (N_1869,N_1413,N_986);
nor U1870 (N_1870,N_1125,N_844);
nor U1871 (N_1871,N_996,N_818);
or U1872 (N_1872,N_930,N_1421);
nor U1873 (N_1873,N_1047,N_1402);
and U1874 (N_1874,N_865,N_1400);
or U1875 (N_1875,N_997,N_1302);
and U1876 (N_1876,N_1187,N_877);
or U1877 (N_1877,N_1464,N_851);
nor U1878 (N_1878,N_791,N_819);
or U1879 (N_1879,N_1303,N_849);
and U1880 (N_1880,N_941,N_1137);
nor U1881 (N_1881,N_1044,N_1059);
nor U1882 (N_1882,N_1053,N_1482);
nor U1883 (N_1883,N_828,N_872);
nor U1884 (N_1884,N_796,N_1413);
nand U1885 (N_1885,N_1372,N_1327);
nand U1886 (N_1886,N_790,N_937);
and U1887 (N_1887,N_882,N_916);
nor U1888 (N_1888,N_1027,N_1485);
and U1889 (N_1889,N_1200,N_1430);
nand U1890 (N_1890,N_1334,N_1036);
or U1891 (N_1891,N_750,N_866);
nor U1892 (N_1892,N_1077,N_1452);
nand U1893 (N_1893,N_795,N_1486);
and U1894 (N_1894,N_1227,N_1096);
and U1895 (N_1895,N_944,N_1011);
and U1896 (N_1896,N_1020,N_1066);
nand U1897 (N_1897,N_886,N_894);
nand U1898 (N_1898,N_1026,N_1382);
or U1899 (N_1899,N_982,N_966);
or U1900 (N_1900,N_1098,N_882);
nand U1901 (N_1901,N_993,N_1351);
nor U1902 (N_1902,N_1327,N_1411);
nand U1903 (N_1903,N_1046,N_1284);
nand U1904 (N_1904,N_960,N_843);
and U1905 (N_1905,N_1269,N_1413);
nand U1906 (N_1906,N_1405,N_921);
nand U1907 (N_1907,N_804,N_900);
nor U1908 (N_1908,N_769,N_1343);
nand U1909 (N_1909,N_1385,N_1267);
xor U1910 (N_1910,N_948,N_984);
and U1911 (N_1911,N_1152,N_910);
nor U1912 (N_1912,N_1262,N_1296);
or U1913 (N_1913,N_1445,N_1056);
nand U1914 (N_1914,N_810,N_1237);
nand U1915 (N_1915,N_1186,N_1330);
or U1916 (N_1916,N_1438,N_1473);
nand U1917 (N_1917,N_766,N_1135);
nor U1918 (N_1918,N_1166,N_1101);
nor U1919 (N_1919,N_1472,N_848);
and U1920 (N_1920,N_799,N_1286);
nor U1921 (N_1921,N_1248,N_1151);
nor U1922 (N_1922,N_1484,N_971);
nor U1923 (N_1923,N_1176,N_1455);
and U1924 (N_1924,N_1185,N_878);
and U1925 (N_1925,N_1335,N_1201);
and U1926 (N_1926,N_1173,N_911);
nand U1927 (N_1927,N_820,N_1061);
nor U1928 (N_1928,N_1447,N_951);
and U1929 (N_1929,N_1419,N_961);
nand U1930 (N_1930,N_772,N_803);
or U1931 (N_1931,N_995,N_1364);
and U1932 (N_1932,N_1217,N_815);
and U1933 (N_1933,N_772,N_1143);
and U1934 (N_1934,N_1294,N_1323);
nor U1935 (N_1935,N_1048,N_856);
nor U1936 (N_1936,N_1186,N_1109);
and U1937 (N_1937,N_1151,N_919);
nand U1938 (N_1938,N_1149,N_1294);
or U1939 (N_1939,N_1476,N_774);
nor U1940 (N_1940,N_982,N_1002);
or U1941 (N_1941,N_1345,N_1402);
nor U1942 (N_1942,N_865,N_761);
and U1943 (N_1943,N_1379,N_1265);
and U1944 (N_1944,N_1069,N_804);
nor U1945 (N_1945,N_1374,N_1380);
nor U1946 (N_1946,N_983,N_1195);
nand U1947 (N_1947,N_1242,N_1227);
or U1948 (N_1948,N_1020,N_887);
nand U1949 (N_1949,N_1332,N_796);
or U1950 (N_1950,N_883,N_1180);
and U1951 (N_1951,N_1454,N_923);
nor U1952 (N_1952,N_998,N_1038);
or U1953 (N_1953,N_1020,N_1251);
nand U1954 (N_1954,N_1324,N_1174);
or U1955 (N_1955,N_1057,N_1047);
nor U1956 (N_1956,N_1291,N_981);
nand U1957 (N_1957,N_1092,N_968);
nand U1958 (N_1958,N_1261,N_1263);
and U1959 (N_1959,N_1446,N_1496);
nand U1960 (N_1960,N_763,N_1154);
nor U1961 (N_1961,N_1194,N_775);
nand U1962 (N_1962,N_1245,N_1301);
or U1963 (N_1963,N_1246,N_1189);
and U1964 (N_1964,N_980,N_1387);
xnor U1965 (N_1965,N_962,N_813);
nand U1966 (N_1966,N_1484,N_840);
nand U1967 (N_1967,N_1458,N_1435);
and U1968 (N_1968,N_778,N_971);
or U1969 (N_1969,N_1478,N_1333);
or U1970 (N_1970,N_1153,N_1190);
or U1971 (N_1971,N_1452,N_1096);
nand U1972 (N_1972,N_1025,N_1291);
nor U1973 (N_1973,N_1155,N_1356);
and U1974 (N_1974,N_803,N_794);
nand U1975 (N_1975,N_761,N_1425);
or U1976 (N_1976,N_888,N_1296);
and U1977 (N_1977,N_1468,N_1287);
or U1978 (N_1978,N_1363,N_1328);
nand U1979 (N_1979,N_886,N_1312);
or U1980 (N_1980,N_1442,N_1039);
nand U1981 (N_1981,N_853,N_1420);
nor U1982 (N_1982,N_960,N_1259);
nand U1983 (N_1983,N_888,N_1071);
nor U1984 (N_1984,N_1468,N_1284);
and U1985 (N_1985,N_1114,N_1264);
nand U1986 (N_1986,N_1420,N_1267);
nand U1987 (N_1987,N_1238,N_1272);
or U1988 (N_1988,N_913,N_1151);
nand U1989 (N_1989,N_1335,N_993);
and U1990 (N_1990,N_1483,N_966);
nand U1991 (N_1991,N_1109,N_834);
nand U1992 (N_1992,N_1266,N_1433);
nand U1993 (N_1993,N_1438,N_1104);
and U1994 (N_1994,N_1288,N_1386);
nor U1995 (N_1995,N_1337,N_994);
or U1996 (N_1996,N_1139,N_1413);
nor U1997 (N_1997,N_1008,N_1325);
and U1998 (N_1998,N_956,N_1309);
nor U1999 (N_1999,N_1325,N_1230);
nand U2000 (N_2000,N_1163,N_1260);
nand U2001 (N_2001,N_913,N_1190);
nand U2002 (N_2002,N_924,N_1199);
nor U2003 (N_2003,N_979,N_1319);
nand U2004 (N_2004,N_1307,N_777);
and U2005 (N_2005,N_1036,N_919);
and U2006 (N_2006,N_1442,N_1191);
nand U2007 (N_2007,N_1482,N_924);
and U2008 (N_2008,N_852,N_898);
nand U2009 (N_2009,N_970,N_1474);
or U2010 (N_2010,N_1363,N_987);
nand U2011 (N_2011,N_1454,N_1080);
nor U2012 (N_2012,N_923,N_1455);
and U2013 (N_2013,N_1012,N_1131);
and U2014 (N_2014,N_1447,N_1478);
and U2015 (N_2015,N_1215,N_1301);
nor U2016 (N_2016,N_1296,N_1099);
nor U2017 (N_2017,N_851,N_1417);
or U2018 (N_2018,N_942,N_834);
nor U2019 (N_2019,N_833,N_1287);
and U2020 (N_2020,N_819,N_1308);
and U2021 (N_2021,N_1019,N_1109);
and U2022 (N_2022,N_984,N_1350);
xnor U2023 (N_2023,N_1349,N_1437);
nand U2024 (N_2024,N_844,N_781);
nand U2025 (N_2025,N_1436,N_1070);
nor U2026 (N_2026,N_961,N_1246);
nand U2027 (N_2027,N_1325,N_1422);
nand U2028 (N_2028,N_1177,N_1110);
and U2029 (N_2029,N_1279,N_965);
nor U2030 (N_2030,N_1181,N_773);
nor U2031 (N_2031,N_1494,N_769);
and U2032 (N_2032,N_938,N_1220);
or U2033 (N_2033,N_1263,N_1428);
or U2034 (N_2034,N_1480,N_1046);
nor U2035 (N_2035,N_777,N_792);
nor U2036 (N_2036,N_995,N_1080);
xor U2037 (N_2037,N_1022,N_1190);
nand U2038 (N_2038,N_1257,N_1207);
and U2039 (N_2039,N_1011,N_929);
nor U2040 (N_2040,N_899,N_1487);
or U2041 (N_2041,N_870,N_971);
or U2042 (N_2042,N_858,N_1387);
or U2043 (N_2043,N_1083,N_1233);
nand U2044 (N_2044,N_1226,N_1187);
or U2045 (N_2045,N_1358,N_1024);
nor U2046 (N_2046,N_937,N_1185);
nor U2047 (N_2047,N_939,N_902);
nand U2048 (N_2048,N_1449,N_945);
nor U2049 (N_2049,N_815,N_804);
or U2050 (N_2050,N_1021,N_996);
nand U2051 (N_2051,N_1444,N_1308);
nand U2052 (N_2052,N_1222,N_845);
or U2053 (N_2053,N_1040,N_1118);
nand U2054 (N_2054,N_1378,N_1463);
and U2055 (N_2055,N_1236,N_1109);
nor U2056 (N_2056,N_1313,N_1217);
and U2057 (N_2057,N_1357,N_1032);
and U2058 (N_2058,N_1442,N_1411);
nor U2059 (N_2059,N_886,N_1347);
and U2060 (N_2060,N_1401,N_962);
and U2061 (N_2061,N_1025,N_1336);
or U2062 (N_2062,N_1234,N_1097);
nand U2063 (N_2063,N_1187,N_782);
or U2064 (N_2064,N_951,N_1155);
nand U2065 (N_2065,N_1389,N_1303);
nor U2066 (N_2066,N_1251,N_1318);
xnor U2067 (N_2067,N_980,N_1180);
and U2068 (N_2068,N_773,N_1027);
or U2069 (N_2069,N_1220,N_1231);
nand U2070 (N_2070,N_1211,N_1187);
nand U2071 (N_2071,N_1192,N_1041);
nand U2072 (N_2072,N_849,N_1404);
nor U2073 (N_2073,N_918,N_791);
or U2074 (N_2074,N_924,N_1462);
nor U2075 (N_2075,N_770,N_1190);
and U2076 (N_2076,N_1182,N_924);
nor U2077 (N_2077,N_812,N_1368);
nand U2078 (N_2078,N_798,N_1480);
nand U2079 (N_2079,N_1330,N_1400);
or U2080 (N_2080,N_1267,N_1376);
or U2081 (N_2081,N_1310,N_983);
nand U2082 (N_2082,N_1222,N_1493);
and U2083 (N_2083,N_905,N_994);
nor U2084 (N_2084,N_1376,N_788);
nand U2085 (N_2085,N_1342,N_1383);
and U2086 (N_2086,N_799,N_1115);
or U2087 (N_2087,N_1490,N_909);
nor U2088 (N_2088,N_1207,N_1080);
or U2089 (N_2089,N_1018,N_1146);
nand U2090 (N_2090,N_806,N_1048);
nand U2091 (N_2091,N_1011,N_1423);
and U2092 (N_2092,N_1020,N_1182);
or U2093 (N_2093,N_1244,N_1067);
and U2094 (N_2094,N_769,N_914);
or U2095 (N_2095,N_758,N_811);
nand U2096 (N_2096,N_828,N_990);
or U2097 (N_2097,N_1138,N_1288);
and U2098 (N_2098,N_1438,N_1305);
and U2099 (N_2099,N_1064,N_772);
nor U2100 (N_2100,N_822,N_1254);
or U2101 (N_2101,N_1231,N_924);
and U2102 (N_2102,N_1163,N_830);
or U2103 (N_2103,N_1135,N_814);
xor U2104 (N_2104,N_1434,N_1452);
or U2105 (N_2105,N_1080,N_1000);
nand U2106 (N_2106,N_1039,N_1363);
and U2107 (N_2107,N_858,N_1119);
nor U2108 (N_2108,N_909,N_1378);
nand U2109 (N_2109,N_912,N_1015);
and U2110 (N_2110,N_1347,N_1350);
or U2111 (N_2111,N_1370,N_1124);
and U2112 (N_2112,N_1086,N_1327);
or U2113 (N_2113,N_1057,N_1305);
or U2114 (N_2114,N_1234,N_1117);
nand U2115 (N_2115,N_1106,N_1359);
nand U2116 (N_2116,N_1357,N_1242);
or U2117 (N_2117,N_1010,N_866);
or U2118 (N_2118,N_1092,N_891);
nor U2119 (N_2119,N_1414,N_859);
or U2120 (N_2120,N_1315,N_1376);
or U2121 (N_2121,N_960,N_788);
nand U2122 (N_2122,N_773,N_854);
or U2123 (N_2123,N_1167,N_1190);
or U2124 (N_2124,N_940,N_1478);
nor U2125 (N_2125,N_1379,N_1151);
or U2126 (N_2126,N_1131,N_1073);
nor U2127 (N_2127,N_826,N_1311);
nor U2128 (N_2128,N_924,N_766);
or U2129 (N_2129,N_1379,N_1072);
or U2130 (N_2130,N_1219,N_1312);
nor U2131 (N_2131,N_789,N_1308);
nor U2132 (N_2132,N_1440,N_1386);
and U2133 (N_2133,N_862,N_1487);
or U2134 (N_2134,N_1290,N_1352);
and U2135 (N_2135,N_1007,N_925);
nand U2136 (N_2136,N_765,N_1050);
nor U2137 (N_2137,N_766,N_1372);
nand U2138 (N_2138,N_842,N_961);
and U2139 (N_2139,N_1461,N_1329);
nand U2140 (N_2140,N_1352,N_1158);
and U2141 (N_2141,N_1280,N_1150);
or U2142 (N_2142,N_1138,N_1279);
or U2143 (N_2143,N_814,N_1248);
nand U2144 (N_2144,N_950,N_884);
or U2145 (N_2145,N_754,N_1195);
or U2146 (N_2146,N_941,N_859);
and U2147 (N_2147,N_800,N_1372);
nand U2148 (N_2148,N_947,N_1048);
nor U2149 (N_2149,N_790,N_1011);
nor U2150 (N_2150,N_1045,N_860);
nand U2151 (N_2151,N_793,N_1441);
nor U2152 (N_2152,N_1086,N_904);
nor U2153 (N_2153,N_763,N_1171);
nor U2154 (N_2154,N_1442,N_845);
and U2155 (N_2155,N_757,N_1055);
or U2156 (N_2156,N_1169,N_1388);
nand U2157 (N_2157,N_1449,N_1067);
or U2158 (N_2158,N_1355,N_1479);
nand U2159 (N_2159,N_1117,N_921);
nand U2160 (N_2160,N_998,N_871);
nand U2161 (N_2161,N_785,N_916);
nand U2162 (N_2162,N_1341,N_949);
nand U2163 (N_2163,N_1256,N_786);
nor U2164 (N_2164,N_941,N_1370);
and U2165 (N_2165,N_1295,N_1162);
and U2166 (N_2166,N_1467,N_912);
and U2167 (N_2167,N_1070,N_1081);
and U2168 (N_2168,N_1286,N_882);
nand U2169 (N_2169,N_1470,N_1437);
and U2170 (N_2170,N_1383,N_1023);
and U2171 (N_2171,N_825,N_998);
nor U2172 (N_2172,N_1300,N_1131);
or U2173 (N_2173,N_925,N_1437);
or U2174 (N_2174,N_1321,N_1225);
or U2175 (N_2175,N_1281,N_836);
or U2176 (N_2176,N_1437,N_812);
and U2177 (N_2177,N_1020,N_889);
or U2178 (N_2178,N_1307,N_913);
nor U2179 (N_2179,N_1468,N_903);
or U2180 (N_2180,N_1041,N_1147);
nor U2181 (N_2181,N_979,N_1423);
nor U2182 (N_2182,N_1460,N_1181);
or U2183 (N_2183,N_973,N_821);
or U2184 (N_2184,N_1316,N_1344);
nand U2185 (N_2185,N_1125,N_1296);
nand U2186 (N_2186,N_1289,N_1482);
nand U2187 (N_2187,N_781,N_1237);
and U2188 (N_2188,N_1409,N_1353);
or U2189 (N_2189,N_1278,N_818);
or U2190 (N_2190,N_1325,N_981);
and U2191 (N_2191,N_979,N_1357);
nand U2192 (N_2192,N_1162,N_1255);
nand U2193 (N_2193,N_1439,N_806);
nand U2194 (N_2194,N_970,N_1184);
nand U2195 (N_2195,N_864,N_1029);
nand U2196 (N_2196,N_1256,N_792);
or U2197 (N_2197,N_761,N_1135);
nand U2198 (N_2198,N_1259,N_1345);
nand U2199 (N_2199,N_1034,N_804);
nor U2200 (N_2200,N_1093,N_1056);
or U2201 (N_2201,N_1327,N_1408);
nor U2202 (N_2202,N_1048,N_1261);
and U2203 (N_2203,N_1457,N_1034);
nand U2204 (N_2204,N_1431,N_931);
nor U2205 (N_2205,N_1300,N_963);
nor U2206 (N_2206,N_1224,N_1430);
and U2207 (N_2207,N_823,N_915);
nor U2208 (N_2208,N_1323,N_1092);
nor U2209 (N_2209,N_1460,N_1286);
and U2210 (N_2210,N_1356,N_1406);
nand U2211 (N_2211,N_1324,N_1032);
and U2212 (N_2212,N_982,N_1324);
or U2213 (N_2213,N_1088,N_1137);
and U2214 (N_2214,N_1289,N_1101);
and U2215 (N_2215,N_1313,N_1281);
nand U2216 (N_2216,N_1199,N_1417);
nor U2217 (N_2217,N_1456,N_1352);
or U2218 (N_2218,N_1357,N_1340);
or U2219 (N_2219,N_1416,N_1377);
and U2220 (N_2220,N_995,N_881);
or U2221 (N_2221,N_1243,N_1045);
and U2222 (N_2222,N_962,N_1064);
or U2223 (N_2223,N_965,N_1203);
nor U2224 (N_2224,N_1441,N_1240);
nor U2225 (N_2225,N_938,N_1155);
nor U2226 (N_2226,N_1146,N_1029);
or U2227 (N_2227,N_1434,N_1241);
nand U2228 (N_2228,N_1009,N_857);
or U2229 (N_2229,N_1407,N_1263);
or U2230 (N_2230,N_955,N_904);
or U2231 (N_2231,N_976,N_1086);
nand U2232 (N_2232,N_1205,N_859);
nand U2233 (N_2233,N_1392,N_1110);
nor U2234 (N_2234,N_1163,N_1249);
nor U2235 (N_2235,N_1030,N_1472);
nand U2236 (N_2236,N_1210,N_953);
nor U2237 (N_2237,N_1051,N_774);
nand U2238 (N_2238,N_1200,N_1161);
nand U2239 (N_2239,N_1070,N_752);
nand U2240 (N_2240,N_1104,N_1453);
nor U2241 (N_2241,N_1116,N_1369);
nand U2242 (N_2242,N_1353,N_1369);
nand U2243 (N_2243,N_949,N_965);
nand U2244 (N_2244,N_935,N_863);
or U2245 (N_2245,N_762,N_820);
nor U2246 (N_2246,N_781,N_1224);
and U2247 (N_2247,N_1110,N_1260);
and U2248 (N_2248,N_1275,N_1082);
nor U2249 (N_2249,N_1188,N_985);
nand U2250 (N_2250,N_1818,N_1800);
and U2251 (N_2251,N_1558,N_2247);
or U2252 (N_2252,N_1516,N_1847);
xor U2253 (N_2253,N_1965,N_2241);
and U2254 (N_2254,N_1568,N_1628);
nand U2255 (N_2255,N_1890,N_2114);
nor U2256 (N_2256,N_1569,N_1626);
nand U2257 (N_2257,N_2035,N_1987);
or U2258 (N_2258,N_2151,N_1605);
nor U2259 (N_2259,N_2193,N_2033);
or U2260 (N_2260,N_1678,N_1868);
and U2261 (N_2261,N_1713,N_1662);
nor U2262 (N_2262,N_1637,N_2233);
or U2263 (N_2263,N_1921,N_1724);
or U2264 (N_2264,N_2089,N_1880);
nor U2265 (N_2265,N_1769,N_1993);
nor U2266 (N_2266,N_1524,N_1795);
nand U2267 (N_2267,N_1961,N_2084);
or U2268 (N_2268,N_1913,N_2112);
or U2269 (N_2269,N_1956,N_1946);
or U2270 (N_2270,N_1525,N_2166);
nor U2271 (N_2271,N_1739,N_2020);
nor U2272 (N_2272,N_1758,N_1634);
nand U2273 (N_2273,N_1792,N_2230);
or U2274 (N_2274,N_2107,N_2021);
or U2275 (N_2275,N_2153,N_1819);
xor U2276 (N_2276,N_1911,N_2212);
nand U2277 (N_2277,N_1740,N_1589);
and U2278 (N_2278,N_2170,N_2177);
and U2279 (N_2279,N_1580,N_2126);
xnor U2280 (N_2280,N_2064,N_2055);
or U2281 (N_2281,N_2186,N_1508);
nand U2282 (N_2282,N_2156,N_1572);
and U2283 (N_2283,N_1518,N_1991);
and U2284 (N_2284,N_1728,N_1875);
nor U2285 (N_2285,N_2174,N_1658);
nor U2286 (N_2286,N_2147,N_1561);
or U2287 (N_2287,N_2092,N_1839);
or U2288 (N_2288,N_1682,N_1867);
nand U2289 (N_2289,N_1900,N_1559);
nor U2290 (N_2290,N_2205,N_1884);
or U2291 (N_2291,N_1846,N_2108);
or U2292 (N_2292,N_1644,N_1708);
nor U2293 (N_2293,N_1711,N_1777);
or U2294 (N_2294,N_1738,N_1659);
nand U2295 (N_2295,N_1726,N_2217);
nor U2296 (N_2296,N_1958,N_1891);
nor U2297 (N_2297,N_1825,N_1601);
nand U2298 (N_2298,N_1530,N_2145);
and U2299 (N_2299,N_1754,N_2219);
and U2300 (N_2300,N_1920,N_1521);
and U2301 (N_2301,N_1977,N_1794);
xnor U2302 (N_2302,N_1994,N_1814);
and U2303 (N_2303,N_1618,N_1630);
and U2304 (N_2304,N_1934,N_2066);
and U2305 (N_2305,N_1592,N_2201);
and U2306 (N_2306,N_1995,N_2133);
and U2307 (N_2307,N_1859,N_2125);
or U2308 (N_2308,N_1865,N_1504);
nand U2309 (N_2309,N_1509,N_1849);
and U2310 (N_2310,N_2063,N_2218);
or U2311 (N_2311,N_1517,N_1645);
and U2312 (N_2312,N_2185,N_1749);
xor U2313 (N_2313,N_1663,N_2142);
and U2314 (N_2314,N_2175,N_2083);
nand U2315 (N_2315,N_1673,N_2011);
or U2316 (N_2316,N_1586,N_1863);
nor U2317 (N_2317,N_2208,N_1801);
nor U2318 (N_2318,N_1514,N_2103);
nor U2319 (N_2319,N_1510,N_1979);
nand U2320 (N_2320,N_1941,N_1939);
nor U2321 (N_2321,N_2051,N_2008);
and U2322 (N_2322,N_1883,N_2235);
nor U2323 (N_2323,N_1808,N_2221);
or U2324 (N_2324,N_1803,N_1692);
nor U2325 (N_2325,N_1748,N_1523);
nand U2326 (N_2326,N_1700,N_2067);
nand U2327 (N_2327,N_1540,N_1789);
nor U2328 (N_2328,N_1973,N_2072);
nand U2329 (N_2329,N_1940,N_1538);
or U2330 (N_2330,N_1683,N_1963);
nor U2331 (N_2331,N_2016,N_2117);
nand U2332 (N_2332,N_1886,N_1674);
or U2333 (N_2333,N_1797,N_1985);
nand U2334 (N_2334,N_2206,N_1791);
nand U2335 (N_2335,N_1968,N_1858);
xor U2336 (N_2336,N_1710,N_2227);
nand U2337 (N_2337,N_2118,N_1672);
and U2338 (N_2338,N_1997,N_1768);
nor U2339 (N_2339,N_2044,N_1652);
nand U2340 (N_2340,N_2123,N_1746);
and U2341 (N_2341,N_1571,N_1869);
nor U2342 (N_2342,N_1501,N_1786);
nand U2343 (N_2343,N_2018,N_1541);
nand U2344 (N_2344,N_2113,N_1547);
and U2345 (N_2345,N_1766,N_2138);
and U2346 (N_2346,N_1996,N_2000);
or U2347 (N_2347,N_1930,N_2246);
or U2348 (N_2348,N_2229,N_1604);
nand U2349 (N_2349,N_1550,N_1902);
nor U2350 (N_2350,N_1924,N_1776);
nand U2351 (N_2351,N_2155,N_2100);
nor U2352 (N_2352,N_2028,N_1815);
nand U2353 (N_2353,N_1585,N_2149);
nor U2354 (N_2354,N_1506,N_2095);
or U2355 (N_2355,N_2025,N_1704);
and U2356 (N_2356,N_1533,N_2101);
or U2357 (N_2357,N_2176,N_2096);
nor U2358 (N_2358,N_2098,N_1870);
or U2359 (N_2359,N_1836,N_1755);
nand U2360 (N_2360,N_1646,N_1929);
nor U2361 (N_2361,N_2168,N_1966);
nand U2362 (N_2362,N_1842,N_1602);
and U2363 (N_2363,N_1519,N_1608);
and U2364 (N_2364,N_1744,N_1681);
nor U2365 (N_2365,N_2165,N_2194);
or U2366 (N_2366,N_1730,N_2191);
xnor U2367 (N_2367,N_1885,N_1654);
nand U2368 (N_2368,N_1838,N_2248);
nand U2369 (N_2369,N_2071,N_1935);
or U2370 (N_2370,N_2013,N_2074);
or U2371 (N_2371,N_1596,N_2130);
nor U2372 (N_2372,N_2243,N_1898);
and U2373 (N_2373,N_1822,N_1906);
nor U2374 (N_2374,N_2187,N_1856);
nor U2375 (N_2375,N_2214,N_1931);
nor U2376 (N_2376,N_1600,N_1549);
or U2377 (N_2377,N_2245,N_1553);
nor U2378 (N_2378,N_1745,N_1761);
nor U2379 (N_2379,N_2228,N_1736);
nand U2380 (N_2380,N_1999,N_1820);
or U2381 (N_2381,N_1715,N_1503);
nor U2382 (N_2382,N_1986,N_2036);
and U2383 (N_2383,N_1593,N_1942);
nor U2384 (N_2384,N_1679,N_1691);
xor U2385 (N_2385,N_1882,N_1537);
nand U2386 (N_2386,N_2158,N_2057);
or U2387 (N_2387,N_2132,N_1978);
or U2388 (N_2388,N_1741,N_2034);
or U2389 (N_2389,N_1775,N_1716);
or U2390 (N_2390,N_2124,N_1639);
nor U2391 (N_2391,N_2070,N_1778);
or U2392 (N_2392,N_1823,N_2102);
or U2393 (N_2393,N_1937,N_1955);
or U2394 (N_2394,N_2090,N_1765);
nand U2395 (N_2395,N_2062,N_1845);
and U2396 (N_2396,N_1718,N_2082);
or U2397 (N_2397,N_1699,N_1922);
or U2398 (N_2398,N_1657,N_1927);
nor U2399 (N_2399,N_1742,N_1636);
and U2400 (N_2400,N_2146,N_1841);
or U2401 (N_2401,N_2068,N_1623);
or U2402 (N_2402,N_2189,N_1960);
nand U2403 (N_2403,N_1954,N_1528);
nand U2404 (N_2404,N_2197,N_2047);
or U2405 (N_2405,N_1899,N_1563);
and U2406 (N_2406,N_1896,N_2224);
nand U2407 (N_2407,N_2129,N_1835);
or U2408 (N_2408,N_1722,N_2131);
nor U2409 (N_2409,N_1629,N_1735);
nand U2410 (N_2410,N_2003,N_1560);
nor U2411 (N_2411,N_2210,N_2216);
and U2412 (N_2412,N_2014,N_1953);
nor U2413 (N_2413,N_1638,N_1879);
nor U2414 (N_2414,N_1535,N_1829);
nand U2415 (N_2415,N_2106,N_1779);
and U2416 (N_2416,N_1774,N_1689);
or U2417 (N_2417,N_2198,N_2204);
nand U2418 (N_2418,N_1967,N_1980);
or U2419 (N_2419,N_1969,N_1762);
and U2420 (N_2420,N_2086,N_2046);
nand U2421 (N_2421,N_2136,N_2094);
nand U2422 (N_2422,N_1680,N_2069);
nor U2423 (N_2423,N_1983,N_2183);
nand U2424 (N_2424,N_2009,N_1947);
nand U2425 (N_2425,N_1964,N_1976);
or U2426 (N_2426,N_1734,N_1824);
nand U2427 (N_2427,N_1709,N_1731);
and U2428 (N_2428,N_1587,N_1564);
nand U2429 (N_2429,N_1633,N_2052);
nand U2430 (N_2430,N_1944,N_1671);
nor U2431 (N_2431,N_1893,N_2211);
or U2432 (N_2432,N_1767,N_1871);
or U2433 (N_2433,N_1613,N_1799);
or U2434 (N_2434,N_2060,N_1698);
nor U2435 (N_2435,N_2111,N_1543);
or U2436 (N_2436,N_1677,N_1915);
nand U2437 (N_2437,N_1990,N_1759);
and U2438 (N_2438,N_2099,N_1594);
or U2439 (N_2439,N_1932,N_1912);
nor U2440 (N_2440,N_2030,N_2029);
and U2441 (N_2441,N_1850,N_1567);
and U2442 (N_2442,N_2043,N_1751);
or U2443 (N_2443,N_1579,N_1661);
nor U2444 (N_2444,N_1784,N_2244);
nor U2445 (N_2445,N_1702,N_2157);
or U2446 (N_2446,N_1536,N_2154);
xor U2447 (N_2447,N_1620,N_1574);
nor U2448 (N_2448,N_1840,N_1526);
or U2449 (N_2449,N_2007,N_1720);
or U2450 (N_2450,N_1887,N_1612);
nor U2451 (N_2451,N_2061,N_1916);
and U2452 (N_2452,N_1998,N_2002);
nor U2453 (N_2453,N_1705,N_1752);
nor U2454 (N_2454,N_1539,N_1649);
and U2455 (N_2455,N_2143,N_1575);
nor U2456 (N_2456,N_2249,N_1812);
or U2457 (N_2457,N_1643,N_1675);
or U2458 (N_2458,N_1546,N_1610);
nor U2459 (N_2459,N_1562,N_1527);
nand U2460 (N_2460,N_2160,N_1952);
or U2461 (N_2461,N_1771,N_2027);
nand U2462 (N_2462,N_1693,N_1895);
or U2463 (N_2463,N_1544,N_1642);
nand U2464 (N_2464,N_2164,N_2182);
and U2465 (N_2465,N_1810,N_1548);
or U2466 (N_2466,N_2234,N_1584);
nand U2467 (N_2467,N_1876,N_1905);
nor U2468 (N_2468,N_1670,N_1936);
nand U2469 (N_2469,N_2159,N_1591);
nor U2470 (N_2470,N_1798,N_1772);
xor U2471 (N_2471,N_1655,N_1512);
nand U2472 (N_2472,N_1757,N_1793);
nand U2473 (N_2473,N_2137,N_1889);
or U2474 (N_2474,N_1933,N_1703);
and U2475 (N_2475,N_1597,N_1743);
and U2476 (N_2476,N_1534,N_2163);
nand U2477 (N_2477,N_1872,N_1653);
or U2478 (N_2478,N_2073,N_2161);
nor U2479 (N_2479,N_1529,N_2110);
or U2480 (N_2480,N_2032,N_2215);
nor U2481 (N_2481,N_1668,N_2041);
and U2482 (N_2482,N_2237,N_1500);
and U2483 (N_2483,N_2076,N_1764);
xnor U2484 (N_2484,N_1938,N_2022);
and U2485 (N_2485,N_1783,N_1656);
or U2486 (N_2486,N_1611,N_2152);
or U2487 (N_2487,N_1619,N_1844);
and U2488 (N_2488,N_1923,N_1949);
nor U2489 (N_2489,N_2162,N_1982);
or U2490 (N_2490,N_2012,N_2209);
nor U2491 (N_2491,N_1917,N_1542);
nor U2492 (N_2492,N_2037,N_1837);
and U2493 (N_2493,N_1894,N_1651);
nor U2494 (N_2494,N_2220,N_2150);
nor U2495 (N_2495,N_1972,N_2202);
nor U2496 (N_2496,N_1522,N_1888);
nor U2497 (N_2497,N_2223,N_1635);
or U2498 (N_2498,N_1854,N_2139);
nand U2499 (N_2499,N_2226,N_2038);
and U2500 (N_2500,N_1588,N_1945);
and U2501 (N_2501,N_1811,N_1622);
and U2502 (N_2502,N_1816,N_1780);
nor U2503 (N_2503,N_1796,N_1957);
nor U2504 (N_2504,N_1545,N_1781);
or U2505 (N_2505,N_1782,N_1690);
or U2506 (N_2506,N_1821,N_2054);
or U2507 (N_2507,N_2023,N_1763);
nor U2508 (N_2508,N_1950,N_1919);
or U2509 (N_2509,N_2105,N_1790);
or U2510 (N_2510,N_2173,N_2109);
or U2511 (N_2511,N_1531,N_1832);
nand U2512 (N_2512,N_2196,N_2119);
nor U2513 (N_2513,N_1632,N_2207);
nand U2514 (N_2514,N_2039,N_1862);
nor U2515 (N_2515,N_1992,N_1852);
nor U2516 (N_2516,N_1903,N_1570);
nor U2517 (N_2517,N_1648,N_1551);
or U2518 (N_2518,N_1590,N_2134);
or U2519 (N_2519,N_1855,N_1687);
nor U2520 (N_2520,N_1750,N_1732);
nor U2521 (N_2521,N_1647,N_1603);
nand U2522 (N_2522,N_1676,N_1640);
and U2523 (N_2523,N_2144,N_2075);
or U2524 (N_2524,N_2141,N_1599);
or U2525 (N_2525,N_2093,N_1621);
nand U2526 (N_2526,N_1686,N_2081);
nand U2527 (N_2527,N_1918,N_1688);
xnor U2528 (N_2528,N_1773,N_1970);
nand U2529 (N_2529,N_1520,N_1909);
and U2530 (N_2530,N_2120,N_1733);
and U2531 (N_2531,N_2050,N_1714);
nor U2532 (N_2532,N_1834,N_2087);
nand U2533 (N_2533,N_1723,N_1555);
or U2534 (N_2534,N_1747,N_1928);
and U2535 (N_2535,N_2225,N_1507);
nor U2536 (N_2536,N_1907,N_1984);
nor U2537 (N_2537,N_1566,N_1582);
nor U2538 (N_2538,N_1873,N_2040);
and U2539 (N_2539,N_2042,N_1664);
nor U2540 (N_2540,N_1717,N_1513);
nand U2541 (N_2541,N_1625,N_1515);
and U2542 (N_2542,N_1827,N_2015);
or U2543 (N_2543,N_1813,N_1577);
or U2544 (N_2544,N_1866,N_2053);
nor U2545 (N_2545,N_1556,N_1696);
nand U2546 (N_2546,N_1805,N_1573);
or U2547 (N_2547,N_1989,N_1951);
nor U2548 (N_2548,N_1877,N_1914);
or U2549 (N_2549,N_1861,N_1830);
nor U2550 (N_2550,N_2167,N_1685);
nand U2551 (N_2551,N_1697,N_2058);
and U2552 (N_2552,N_1615,N_1616);
nor U2553 (N_2553,N_2078,N_2188);
and U2554 (N_2554,N_1910,N_1727);
nand U2555 (N_2555,N_1806,N_1753);
or U2556 (N_2556,N_1502,N_2080);
or U2557 (N_2557,N_1650,N_2178);
or U2558 (N_2558,N_2238,N_2240);
and U2559 (N_2559,N_2059,N_2077);
and U2560 (N_2560,N_2065,N_2231);
nand U2561 (N_2561,N_1843,N_2031);
and U2562 (N_2562,N_1881,N_2199);
or U2563 (N_2563,N_1729,N_1988);
nor U2564 (N_2564,N_2184,N_1864);
or U2565 (N_2565,N_2171,N_1943);
nand U2566 (N_2566,N_2200,N_2181);
and U2567 (N_2567,N_2091,N_1807);
or U2568 (N_2568,N_1557,N_2079);
nor U2569 (N_2569,N_2104,N_1667);
nor U2570 (N_2570,N_2148,N_1878);
or U2571 (N_2571,N_1857,N_2135);
or U2572 (N_2572,N_2085,N_1701);
or U2573 (N_2573,N_2190,N_1897);
nor U2574 (N_2574,N_2140,N_1770);
nor U2575 (N_2575,N_1552,N_2017);
nand U2576 (N_2576,N_1860,N_2088);
nand U2577 (N_2577,N_2010,N_1848);
nand U2578 (N_2578,N_2222,N_1631);
and U2579 (N_2579,N_2172,N_2122);
and U2580 (N_2580,N_1641,N_1607);
and U2581 (N_2581,N_1712,N_2006);
and U2582 (N_2582,N_1706,N_1511);
or U2583 (N_2583,N_1609,N_2056);
or U2584 (N_2584,N_1926,N_1554);
or U2585 (N_2585,N_2242,N_1725);
and U2586 (N_2586,N_1660,N_1581);
nor U2587 (N_2587,N_2239,N_1892);
and U2588 (N_2588,N_1853,N_1802);
nand U2589 (N_2589,N_2121,N_1974);
nor U2590 (N_2590,N_1756,N_2097);
nand U2591 (N_2591,N_1606,N_1975);
and U2592 (N_2592,N_2213,N_2127);
nand U2593 (N_2593,N_1669,N_1707);
and U2594 (N_2594,N_2179,N_1981);
nor U2595 (N_2595,N_1826,N_2048);
or U2596 (N_2596,N_1532,N_1833);
and U2597 (N_2597,N_2180,N_1908);
nand U2598 (N_2598,N_2195,N_1694);
nor U2599 (N_2599,N_1719,N_1851);
nor U2600 (N_2600,N_2192,N_1948);
and U2601 (N_2601,N_1578,N_2001);
or U2602 (N_2602,N_2128,N_1831);
nor U2603 (N_2603,N_1576,N_1925);
nand U2604 (N_2604,N_1901,N_1760);
and U2605 (N_2605,N_1788,N_1624);
or U2606 (N_2606,N_2169,N_2045);
nand U2607 (N_2607,N_1565,N_1959);
xor U2608 (N_2608,N_1665,N_1962);
nor U2609 (N_2609,N_1695,N_1684);
nor U2610 (N_2610,N_1666,N_1737);
and U2611 (N_2611,N_2049,N_2232);
nor U2612 (N_2612,N_1785,N_2115);
or U2613 (N_2613,N_1505,N_2019);
nor U2614 (N_2614,N_1787,N_1721);
nand U2615 (N_2615,N_2203,N_1583);
nand U2616 (N_2616,N_1828,N_2116);
or U2617 (N_2617,N_2004,N_1598);
nor U2618 (N_2618,N_1595,N_1809);
or U2619 (N_2619,N_1804,N_1904);
and U2620 (N_2620,N_1874,N_1614);
and U2621 (N_2621,N_1617,N_1971);
nor U2622 (N_2622,N_1817,N_1627);
nor U2623 (N_2623,N_2024,N_2026);
or U2624 (N_2624,N_2005,N_2236);
nand U2625 (N_2625,N_1946,N_1724);
and U2626 (N_2626,N_1998,N_1986);
or U2627 (N_2627,N_1888,N_1997);
or U2628 (N_2628,N_1790,N_1549);
and U2629 (N_2629,N_1666,N_1539);
nor U2630 (N_2630,N_2014,N_2218);
nor U2631 (N_2631,N_1841,N_1932);
nor U2632 (N_2632,N_1590,N_1909);
and U2633 (N_2633,N_1652,N_1799);
xnor U2634 (N_2634,N_1869,N_1975);
nor U2635 (N_2635,N_1894,N_1620);
and U2636 (N_2636,N_1500,N_1726);
or U2637 (N_2637,N_2012,N_1621);
nor U2638 (N_2638,N_1931,N_1680);
nor U2639 (N_2639,N_1752,N_1680);
and U2640 (N_2640,N_1705,N_1789);
nor U2641 (N_2641,N_2200,N_2092);
nand U2642 (N_2642,N_1833,N_2172);
and U2643 (N_2643,N_1658,N_1768);
nand U2644 (N_2644,N_1870,N_1810);
nor U2645 (N_2645,N_1554,N_1580);
and U2646 (N_2646,N_1974,N_1567);
or U2647 (N_2647,N_1780,N_2171);
and U2648 (N_2648,N_1835,N_1596);
and U2649 (N_2649,N_1563,N_2168);
nor U2650 (N_2650,N_2152,N_1977);
or U2651 (N_2651,N_1612,N_2132);
nand U2652 (N_2652,N_1605,N_1922);
nor U2653 (N_2653,N_1710,N_1784);
or U2654 (N_2654,N_2184,N_1872);
or U2655 (N_2655,N_1660,N_1821);
and U2656 (N_2656,N_2098,N_1609);
nor U2657 (N_2657,N_1967,N_1580);
or U2658 (N_2658,N_1715,N_2081);
nand U2659 (N_2659,N_2219,N_1816);
or U2660 (N_2660,N_2210,N_1768);
and U2661 (N_2661,N_2226,N_1879);
or U2662 (N_2662,N_2096,N_1635);
and U2663 (N_2663,N_1903,N_1677);
and U2664 (N_2664,N_1990,N_2156);
or U2665 (N_2665,N_1760,N_1629);
and U2666 (N_2666,N_1724,N_1694);
or U2667 (N_2667,N_1938,N_2144);
nor U2668 (N_2668,N_1924,N_2083);
and U2669 (N_2669,N_1746,N_1903);
nor U2670 (N_2670,N_2196,N_2192);
and U2671 (N_2671,N_2069,N_2126);
nand U2672 (N_2672,N_1755,N_2120);
nor U2673 (N_2673,N_2207,N_2072);
nand U2674 (N_2674,N_1694,N_1616);
nor U2675 (N_2675,N_1727,N_1710);
nand U2676 (N_2676,N_1658,N_1906);
nor U2677 (N_2677,N_1893,N_2053);
nor U2678 (N_2678,N_1747,N_1688);
xor U2679 (N_2679,N_1547,N_1510);
and U2680 (N_2680,N_1904,N_2119);
or U2681 (N_2681,N_1856,N_2018);
nand U2682 (N_2682,N_2124,N_1689);
or U2683 (N_2683,N_1959,N_1582);
or U2684 (N_2684,N_1870,N_1909);
nand U2685 (N_2685,N_1963,N_1639);
and U2686 (N_2686,N_2111,N_1629);
or U2687 (N_2687,N_1865,N_1982);
xor U2688 (N_2688,N_1785,N_1765);
nand U2689 (N_2689,N_2142,N_1598);
nand U2690 (N_2690,N_1956,N_1897);
nand U2691 (N_2691,N_1757,N_1709);
nor U2692 (N_2692,N_1833,N_1741);
nor U2693 (N_2693,N_1840,N_1579);
and U2694 (N_2694,N_1592,N_1582);
and U2695 (N_2695,N_1913,N_1934);
nand U2696 (N_2696,N_2224,N_1598);
nand U2697 (N_2697,N_1974,N_1661);
and U2698 (N_2698,N_2155,N_1945);
nand U2699 (N_2699,N_1798,N_1648);
nor U2700 (N_2700,N_2004,N_1618);
or U2701 (N_2701,N_1609,N_2173);
nor U2702 (N_2702,N_1863,N_1898);
and U2703 (N_2703,N_2106,N_1621);
and U2704 (N_2704,N_1992,N_1600);
and U2705 (N_2705,N_2150,N_1829);
xor U2706 (N_2706,N_1943,N_1559);
nand U2707 (N_2707,N_1730,N_1663);
nand U2708 (N_2708,N_2229,N_2090);
and U2709 (N_2709,N_1833,N_1795);
and U2710 (N_2710,N_2239,N_2098);
or U2711 (N_2711,N_1901,N_1538);
nor U2712 (N_2712,N_1805,N_1501);
nor U2713 (N_2713,N_1926,N_2242);
nand U2714 (N_2714,N_1551,N_2232);
or U2715 (N_2715,N_1634,N_1694);
nor U2716 (N_2716,N_2174,N_2210);
and U2717 (N_2717,N_1976,N_2204);
or U2718 (N_2718,N_1902,N_1672);
nand U2719 (N_2719,N_1565,N_1507);
nor U2720 (N_2720,N_1991,N_1876);
nor U2721 (N_2721,N_2243,N_1798);
nor U2722 (N_2722,N_2017,N_1761);
nand U2723 (N_2723,N_1817,N_1870);
and U2724 (N_2724,N_2023,N_1564);
or U2725 (N_2725,N_2025,N_1674);
nor U2726 (N_2726,N_1793,N_1929);
nor U2727 (N_2727,N_1576,N_1851);
or U2728 (N_2728,N_1951,N_2006);
and U2729 (N_2729,N_1825,N_1705);
nor U2730 (N_2730,N_2141,N_1503);
nand U2731 (N_2731,N_1561,N_1617);
nor U2732 (N_2732,N_1623,N_2072);
or U2733 (N_2733,N_1973,N_1765);
nand U2734 (N_2734,N_1613,N_1596);
or U2735 (N_2735,N_1630,N_1553);
and U2736 (N_2736,N_1570,N_2091);
nor U2737 (N_2737,N_1662,N_2083);
nor U2738 (N_2738,N_2034,N_2025);
and U2739 (N_2739,N_2215,N_1785);
and U2740 (N_2740,N_1997,N_1783);
and U2741 (N_2741,N_2109,N_1553);
or U2742 (N_2742,N_1829,N_1930);
or U2743 (N_2743,N_1546,N_1612);
or U2744 (N_2744,N_1722,N_1592);
nand U2745 (N_2745,N_1758,N_1533);
nor U2746 (N_2746,N_2087,N_1629);
nor U2747 (N_2747,N_2041,N_1505);
and U2748 (N_2748,N_1655,N_1680);
xor U2749 (N_2749,N_1812,N_1510);
nand U2750 (N_2750,N_1673,N_1695);
nor U2751 (N_2751,N_1536,N_1895);
nor U2752 (N_2752,N_1793,N_1962);
nor U2753 (N_2753,N_1920,N_1539);
and U2754 (N_2754,N_2083,N_1622);
nand U2755 (N_2755,N_1672,N_2197);
and U2756 (N_2756,N_2005,N_1860);
or U2757 (N_2757,N_1815,N_2130);
nor U2758 (N_2758,N_2237,N_1762);
nand U2759 (N_2759,N_1912,N_1998);
nand U2760 (N_2760,N_1529,N_1520);
nor U2761 (N_2761,N_1506,N_2205);
nor U2762 (N_2762,N_1945,N_1649);
nand U2763 (N_2763,N_2100,N_2064);
or U2764 (N_2764,N_1992,N_2053);
nand U2765 (N_2765,N_1775,N_1852);
nor U2766 (N_2766,N_2143,N_1951);
or U2767 (N_2767,N_2148,N_1831);
or U2768 (N_2768,N_2016,N_1678);
and U2769 (N_2769,N_1811,N_1807);
and U2770 (N_2770,N_1872,N_1556);
or U2771 (N_2771,N_2066,N_1724);
nand U2772 (N_2772,N_2079,N_1643);
and U2773 (N_2773,N_1919,N_1536);
nand U2774 (N_2774,N_2124,N_2088);
or U2775 (N_2775,N_2145,N_1522);
nor U2776 (N_2776,N_1978,N_2068);
or U2777 (N_2777,N_1519,N_2191);
nor U2778 (N_2778,N_2204,N_1955);
nand U2779 (N_2779,N_1549,N_2011);
nor U2780 (N_2780,N_2114,N_2003);
and U2781 (N_2781,N_2133,N_2039);
and U2782 (N_2782,N_1956,N_1539);
nand U2783 (N_2783,N_2056,N_1986);
nor U2784 (N_2784,N_2008,N_1841);
nand U2785 (N_2785,N_1853,N_1805);
nor U2786 (N_2786,N_1525,N_2177);
nand U2787 (N_2787,N_1632,N_1798);
or U2788 (N_2788,N_1872,N_2224);
or U2789 (N_2789,N_1810,N_1652);
or U2790 (N_2790,N_1947,N_1796);
nand U2791 (N_2791,N_1930,N_1954);
nand U2792 (N_2792,N_1640,N_1894);
nor U2793 (N_2793,N_1884,N_1881);
and U2794 (N_2794,N_2102,N_2248);
and U2795 (N_2795,N_2092,N_1615);
nor U2796 (N_2796,N_1951,N_1712);
nand U2797 (N_2797,N_1912,N_2129);
nand U2798 (N_2798,N_1608,N_1656);
nor U2799 (N_2799,N_1949,N_1970);
and U2800 (N_2800,N_2076,N_1808);
or U2801 (N_2801,N_1719,N_1612);
or U2802 (N_2802,N_2097,N_1930);
and U2803 (N_2803,N_1720,N_1739);
or U2804 (N_2804,N_1929,N_1529);
or U2805 (N_2805,N_1922,N_1642);
nand U2806 (N_2806,N_1700,N_2017);
or U2807 (N_2807,N_1675,N_2200);
nor U2808 (N_2808,N_1539,N_1841);
nand U2809 (N_2809,N_1852,N_1773);
or U2810 (N_2810,N_2051,N_1931);
or U2811 (N_2811,N_1598,N_1515);
nand U2812 (N_2812,N_1507,N_1533);
nand U2813 (N_2813,N_1554,N_1894);
and U2814 (N_2814,N_2246,N_1978);
and U2815 (N_2815,N_1690,N_1544);
xnor U2816 (N_2816,N_2141,N_2182);
nor U2817 (N_2817,N_2154,N_1579);
nand U2818 (N_2818,N_1622,N_2152);
and U2819 (N_2819,N_1821,N_2203);
nand U2820 (N_2820,N_1752,N_2054);
or U2821 (N_2821,N_1868,N_1898);
or U2822 (N_2822,N_1909,N_1626);
or U2823 (N_2823,N_1708,N_2239);
nor U2824 (N_2824,N_2019,N_1567);
and U2825 (N_2825,N_1798,N_1640);
and U2826 (N_2826,N_2218,N_2083);
nor U2827 (N_2827,N_1530,N_1967);
nand U2828 (N_2828,N_2126,N_1911);
nand U2829 (N_2829,N_1897,N_1508);
nand U2830 (N_2830,N_1547,N_1565);
nand U2831 (N_2831,N_2013,N_2216);
and U2832 (N_2832,N_2100,N_1523);
nor U2833 (N_2833,N_1948,N_2007);
and U2834 (N_2834,N_2171,N_1670);
nand U2835 (N_2835,N_1944,N_2185);
nand U2836 (N_2836,N_1775,N_1739);
or U2837 (N_2837,N_2099,N_1616);
nor U2838 (N_2838,N_1732,N_1951);
or U2839 (N_2839,N_2032,N_1900);
nor U2840 (N_2840,N_1649,N_2087);
and U2841 (N_2841,N_1680,N_1922);
nor U2842 (N_2842,N_1888,N_1699);
nand U2843 (N_2843,N_1906,N_1639);
or U2844 (N_2844,N_1680,N_1587);
nand U2845 (N_2845,N_1859,N_2109);
nand U2846 (N_2846,N_1988,N_2009);
nor U2847 (N_2847,N_2204,N_1767);
and U2848 (N_2848,N_2048,N_1746);
nand U2849 (N_2849,N_2104,N_1802);
and U2850 (N_2850,N_2204,N_1918);
and U2851 (N_2851,N_1635,N_1557);
nand U2852 (N_2852,N_1787,N_2163);
or U2853 (N_2853,N_1677,N_2066);
and U2854 (N_2854,N_1996,N_1945);
nor U2855 (N_2855,N_2233,N_1593);
or U2856 (N_2856,N_2042,N_1780);
nand U2857 (N_2857,N_2189,N_1695);
or U2858 (N_2858,N_1681,N_1853);
or U2859 (N_2859,N_1575,N_1548);
nor U2860 (N_2860,N_1877,N_1948);
nor U2861 (N_2861,N_1550,N_2113);
nand U2862 (N_2862,N_1951,N_1888);
and U2863 (N_2863,N_2112,N_2227);
nor U2864 (N_2864,N_1555,N_1909);
nor U2865 (N_2865,N_1654,N_2029);
or U2866 (N_2866,N_1991,N_1578);
nand U2867 (N_2867,N_1978,N_1833);
or U2868 (N_2868,N_2124,N_2015);
nand U2869 (N_2869,N_1891,N_2238);
and U2870 (N_2870,N_2067,N_1560);
nor U2871 (N_2871,N_2159,N_1752);
and U2872 (N_2872,N_2159,N_2126);
nor U2873 (N_2873,N_1764,N_1830);
and U2874 (N_2874,N_1760,N_1989);
or U2875 (N_2875,N_2016,N_2168);
or U2876 (N_2876,N_1987,N_1530);
or U2877 (N_2877,N_1533,N_1916);
xnor U2878 (N_2878,N_2047,N_1564);
nor U2879 (N_2879,N_1609,N_2169);
or U2880 (N_2880,N_2090,N_1882);
or U2881 (N_2881,N_1952,N_2194);
nand U2882 (N_2882,N_1858,N_2070);
nand U2883 (N_2883,N_2094,N_1514);
nor U2884 (N_2884,N_2170,N_1539);
nor U2885 (N_2885,N_2237,N_2157);
nand U2886 (N_2886,N_2248,N_2021);
nor U2887 (N_2887,N_1822,N_1548);
nor U2888 (N_2888,N_1686,N_2112);
and U2889 (N_2889,N_2130,N_1779);
and U2890 (N_2890,N_2238,N_2004);
nor U2891 (N_2891,N_1579,N_2157);
nor U2892 (N_2892,N_2080,N_2207);
and U2893 (N_2893,N_1639,N_2057);
and U2894 (N_2894,N_2113,N_1957);
or U2895 (N_2895,N_2051,N_1851);
nand U2896 (N_2896,N_1540,N_1506);
nor U2897 (N_2897,N_1514,N_1504);
nor U2898 (N_2898,N_1901,N_1947);
and U2899 (N_2899,N_1832,N_1907);
or U2900 (N_2900,N_2209,N_1757);
and U2901 (N_2901,N_1580,N_1716);
nand U2902 (N_2902,N_1504,N_1713);
nand U2903 (N_2903,N_2220,N_1866);
or U2904 (N_2904,N_1861,N_1995);
or U2905 (N_2905,N_1912,N_1893);
nand U2906 (N_2906,N_2005,N_1704);
nor U2907 (N_2907,N_1592,N_2149);
nor U2908 (N_2908,N_1506,N_2184);
nand U2909 (N_2909,N_1867,N_2041);
nor U2910 (N_2910,N_2136,N_1766);
nor U2911 (N_2911,N_1998,N_1966);
nor U2912 (N_2912,N_2083,N_1572);
and U2913 (N_2913,N_1686,N_1691);
nor U2914 (N_2914,N_1587,N_1500);
or U2915 (N_2915,N_1775,N_2220);
nand U2916 (N_2916,N_1784,N_1956);
or U2917 (N_2917,N_2002,N_2107);
nor U2918 (N_2918,N_1887,N_1741);
nor U2919 (N_2919,N_1797,N_2201);
nor U2920 (N_2920,N_1787,N_1901);
and U2921 (N_2921,N_1916,N_1997);
nor U2922 (N_2922,N_1890,N_1960);
nand U2923 (N_2923,N_1954,N_2111);
nor U2924 (N_2924,N_2173,N_2248);
and U2925 (N_2925,N_1704,N_1754);
nand U2926 (N_2926,N_1522,N_1577);
or U2927 (N_2927,N_1782,N_1928);
or U2928 (N_2928,N_1779,N_1817);
nor U2929 (N_2929,N_1541,N_2128);
nor U2930 (N_2930,N_1801,N_1704);
nor U2931 (N_2931,N_2215,N_1546);
nand U2932 (N_2932,N_1737,N_2091);
nor U2933 (N_2933,N_1739,N_1520);
nand U2934 (N_2934,N_1810,N_1520);
nor U2935 (N_2935,N_1708,N_2154);
nand U2936 (N_2936,N_1638,N_1534);
nor U2937 (N_2937,N_1768,N_1995);
nor U2938 (N_2938,N_1584,N_1670);
nor U2939 (N_2939,N_2242,N_2169);
nand U2940 (N_2940,N_1679,N_2025);
and U2941 (N_2941,N_1861,N_2065);
and U2942 (N_2942,N_1590,N_2065);
or U2943 (N_2943,N_1532,N_1842);
or U2944 (N_2944,N_1744,N_1835);
or U2945 (N_2945,N_1872,N_1691);
nand U2946 (N_2946,N_1686,N_1871);
nand U2947 (N_2947,N_1929,N_2084);
nand U2948 (N_2948,N_2202,N_2063);
nand U2949 (N_2949,N_2215,N_1588);
or U2950 (N_2950,N_1932,N_1622);
or U2951 (N_2951,N_1752,N_2122);
nor U2952 (N_2952,N_2097,N_1902);
nand U2953 (N_2953,N_1853,N_2243);
nand U2954 (N_2954,N_1660,N_2245);
nor U2955 (N_2955,N_1502,N_1968);
and U2956 (N_2956,N_1919,N_1650);
nor U2957 (N_2957,N_1878,N_1731);
and U2958 (N_2958,N_1867,N_2186);
nor U2959 (N_2959,N_1660,N_1869);
nor U2960 (N_2960,N_1663,N_2214);
nor U2961 (N_2961,N_2174,N_1737);
or U2962 (N_2962,N_1647,N_1769);
and U2963 (N_2963,N_1552,N_1811);
and U2964 (N_2964,N_1751,N_1931);
or U2965 (N_2965,N_1890,N_2034);
or U2966 (N_2966,N_2242,N_2072);
or U2967 (N_2967,N_1534,N_1881);
or U2968 (N_2968,N_1838,N_1504);
xor U2969 (N_2969,N_1806,N_2020);
nand U2970 (N_2970,N_1909,N_1817);
and U2971 (N_2971,N_1505,N_1654);
and U2972 (N_2972,N_1902,N_1626);
or U2973 (N_2973,N_2030,N_1805);
and U2974 (N_2974,N_1876,N_2069);
and U2975 (N_2975,N_1743,N_2117);
and U2976 (N_2976,N_2235,N_1541);
or U2977 (N_2977,N_1969,N_2079);
nand U2978 (N_2978,N_1658,N_1551);
nand U2979 (N_2979,N_1765,N_1536);
nor U2980 (N_2980,N_1854,N_2098);
xor U2981 (N_2981,N_1555,N_1958);
or U2982 (N_2982,N_2210,N_1615);
nor U2983 (N_2983,N_2150,N_1571);
and U2984 (N_2984,N_1633,N_1727);
nor U2985 (N_2985,N_2124,N_1658);
nor U2986 (N_2986,N_1870,N_1959);
nor U2987 (N_2987,N_1535,N_2051);
and U2988 (N_2988,N_1659,N_2039);
or U2989 (N_2989,N_1769,N_2215);
nand U2990 (N_2990,N_2052,N_1855);
and U2991 (N_2991,N_2178,N_2170);
nand U2992 (N_2992,N_2236,N_1674);
or U2993 (N_2993,N_1751,N_2186);
and U2994 (N_2994,N_1721,N_2240);
nand U2995 (N_2995,N_1882,N_1654);
or U2996 (N_2996,N_1950,N_1861);
and U2997 (N_2997,N_1968,N_1642);
or U2998 (N_2998,N_1582,N_2088);
nand U2999 (N_2999,N_2139,N_1793);
nand UO_0 (O_0,N_2398,N_2691);
nand UO_1 (O_1,N_2445,N_2976);
nor UO_2 (O_2,N_2596,N_2916);
or UO_3 (O_3,N_2870,N_2426);
and UO_4 (O_4,N_2685,N_2969);
and UO_5 (O_5,N_2577,N_2931);
nor UO_6 (O_6,N_2489,N_2463);
and UO_7 (O_7,N_2462,N_2318);
and UO_8 (O_8,N_2741,N_2303);
and UO_9 (O_9,N_2374,N_2472);
nand UO_10 (O_10,N_2401,N_2560);
and UO_11 (O_11,N_2536,N_2387);
and UO_12 (O_12,N_2295,N_2833);
or UO_13 (O_13,N_2350,N_2688);
and UO_14 (O_14,N_2863,N_2565);
and UO_15 (O_15,N_2461,N_2359);
or UO_16 (O_16,N_2621,N_2780);
nor UO_17 (O_17,N_2868,N_2497);
and UO_18 (O_18,N_2332,N_2537);
nand UO_19 (O_19,N_2875,N_2951);
or UO_20 (O_20,N_2635,N_2906);
or UO_21 (O_21,N_2665,N_2442);
and UO_22 (O_22,N_2479,N_2737);
nor UO_23 (O_23,N_2603,N_2519);
or UO_24 (O_24,N_2348,N_2764);
or UO_25 (O_25,N_2858,N_2954);
nor UO_26 (O_26,N_2490,N_2409);
nand UO_27 (O_27,N_2312,N_2844);
or UO_28 (O_28,N_2842,N_2689);
and UO_29 (O_29,N_2559,N_2797);
xnor UO_30 (O_30,N_2676,N_2440);
or UO_31 (O_31,N_2437,N_2404);
and UO_32 (O_32,N_2758,N_2376);
and UO_33 (O_33,N_2418,N_2922);
nor UO_34 (O_34,N_2653,N_2423);
nand UO_35 (O_35,N_2871,N_2602);
and UO_36 (O_36,N_2747,N_2540);
and UO_37 (O_37,N_2711,N_2402);
and UO_38 (O_38,N_2932,N_2852);
and UO_39 (O_39,N_2710,N_2992);
nand UO_40 (O_40,N_2848,N_2471);
xor UO_41 (O_41,N_2891,N_2674);
nor UO_42 (O_42,N_2314,N_2995);
or UO_43 (O_43,N_2802,N_2309);
or UO_44 (O_44,N_2860,N_2601);
and UO_45 (O_45,N_2448,N_2508);
nor UO_46 (O_46,N_2935,N_2584);
or UO_47 (O_47,N_2953,N_2999);
nand UO_48 (O_48,N_2420,N_2680);
nand UO_49 (O_49,N_2591,N_2518);
nand UO_50 (O_50,N_2260,N_2512);
nor UO_51 (O_51,N_2966,N_2517);
nor UO_52 (O_52,N_2934,N_2622);
or UO_53 (O_53,N_2368,N_2849);
or UO_54 (O_54,N_2444,N_2499);
nand UO_55 (O_55,N_2980,N_2470);
or UO_56 (O_56,N_2640,N_2532);
nor UO_57 (O_57,N_2452,N_2269);
nand UO_58 (O_58,N_2322,N_2386);
or UO_59 (O_59,N_2294,N_2415);
nand UO_60 (O_60,N_2738,N_2381);
or UO_61 (O_61,N_2446,N_2832);
and UO_62 (O_62,N_2717,N_2564);
nand UO_63 (O_63,N_2755,N_2553);
and UO_64 (O_64,N_2772,N_2405);
and UO_65 (O_65,N_2261,N_2855);
and UO_66 (O_66,N_2750,N_2830);
and UO_67 (O_67,N_2587,N_2407);
nor UO_68 (O_68,N_2769,N_2439);
nor UO_69 (O_69,N_2687,N_2905);
nor UO_70 (O_70,N_2297,N_2422);
nor UO_71 (O_71,N_2654,N_2250);
or UO_72 (O_72,N_2306,N_2956);
xor UO_73 (O_73,N_2866,N_2826);
nand UO_74 (O_74,N_2666,N_2585);
or UO_75 (O_75,N_2996,N_2697);
and UO_76 (O_76,N_2973,N_2283);
nand UO_77 (O_77,N_2647,N_2997);
or UO_78 (O_78,N_2854,N_2946);
nor UO_79 (O_79,N_2690,N_2828);
nand UO_80 (O_80,N_2695,N_2329);
nand UO_81 (O_81,N_2330,N_2880);
nand UO_82 (O_82,N_2798,N_2626);
and UO_83 (O_83,N_2903,N_2307);
nor UO_84 (O_84,N_2829,N_2790);
and UO_85 (O_85,N_2593,N_2686);
nor UO_86 (O_86,N_2867,N_2841);
nand UO_87 (O_87,N_2943,N_2476);
and UO_88 (O_88,N_2961,N_2554);
nand UO_89 (O_89,N_2364,N_2892);
nor UO_90 (O_90,N_2617,N_2449);
and UO_91 (O_91,N_2313,N_2488);
nand UO_92 (O_92,N_2558,N_2563);
nor UO_93 (O_93,N_2334,N_2734);
or UO_94 (O_94,N_2733,N_2965);
or UO_95 (O_95,N_2949,N_2473);
nand UO_96 (O_96,N_2254,N_2395);
nor UO_97 (O_97,N_2618,N_2958);
nand UO_98 (O_98,N_2457,N_2884);
and UO_99 (O_99,N_2947,N_2881);
nand UO_100 (O_100,N_2373,N_2466);
nand UO_101 (O_101,N_2761,N_2274);
and UO_102 (O_102,N_2713,N_2352);
nand UO_103 (O_103,N_2255,N_2925);
nor UO_104 (O_104,N_2722,N_2664);
or UO_105 (O_105,N_2464,N_2339);
nor UO_106 (O_106,N_2384,N_2263);
and UO_107 (O_107,N_2580,N_2443);
and UO_108 (O_108,N_2456,N_2270);
xor UO_109 (O_109,N_2672,N_2974);
or UO_110 (O_110,N_2824,N_2336);
or UO_111 (O_111,N_2719,N_2290);
and UO_112 (O_112,N_2728,N_2777);
nand UO_113 (O_113,N_2575,N_2643);
and UO_114 (O_114,N_2425,N_2696);
nand UO_115 (O_115,N_2562,N_2576);
or UO_116 (O_116,N_2919,N_2763);
or UO_117 (O_117,N_2438,N_2785);
nor UO_118 (O_118,N_2704,N_2351);
nand UO_119 (O_119,N_2412,N_2474);
and UO_120 (O_120,N_2998,N_2390);
nor UO_121 (O_121,N_2876,N_2740);
and UO_122 (O_122,N_2288,N_2428);
nor UO_123 (O_123,N_2392,N_2963);
nor UO_124 (O_124,N_2441,N_2586);
or UO_125 (O_125,N_2378,N_2421);
nand UO_126 (O_126,N_2846,N_2788);
nand UO_127 (O_127,N_2890,N_2652);
and UO_128 (O_128,N_2569,N_2727);
or UO_129 (O_129,N_2803,N_2492);
or UO_130 (O_130,N_2725,N_2619);
nand UO_131 (O_131,N_2258,N_2262);
and UO_132 (O_132,N_2605,N_2280);
nand UO_133 (O_133,N_2491,N_2944);
and UO_134 (O_134,N_2606,N_2816);
and UO_135 (O_135,N_2272,N_2572);
nand UO_136 (O_136,N_2515,N_2743);
nand UO_137 (O_137,N_2897,N_2343);
nor UO_138 (O_138,N_2311,N_2320);
or UO_139 (O_139,N_2960,N_2305);
or UO_140 (O_140,N_2266,N_2774);
or UO_141 (O_141,N_2450,N_2543);
nor UO_142 (O_142,N_2607,N_2615);
and UO_143 (O_143,N_2534,N_2411);
nor UO_144 (O_144,N_2520,N_2886);
nand UO_145 (O_145,N_2791,N_2549);
nand UO_146 (O_146,N_2732,N_2817);
nand UO_147 (O_147,N_2941,N_2362);
or UO_148 (O_148,N_2358,N_2410);
and UO_149 (O_149,N_2921,N_2708);
or UO_150 (O_150,N_2256,N_2677);
and UO_151 (O_151,N_2590,N_2289);
and UO_152 (O_152,N_2278,N_2639);
or UO_153 (O_153,N_2784,N_2433);
nand UO_154 (O_154,N_2901,N_2762);
nand UO_155 (O_155,N_2918,N_2432);
nor UO_156 (O_156,N_2651,N_2545);
nor UO_157 (O_157,N_2872,N_2909);
nand UO_158 (O_158,N_2782,N_2573);
nand UO_159 (O_159,N_2355,N_2889);
nand UO_160 (O_160,N_2337,N_2693);
or UO_161 (O_161,N_2714,N_2970);
nor UO_162 (O_162,N_2326,N_2478);
and UO_163 (O_163,N_2669,N_2597);
or UO_164 (O_164,N_2513,N_2773);
nor UO_165 (O_165,N_2865,N_2353);
or UO_166 (O_166,N_2363,N_2649);
or UO_167 (O_167,N_2729,N_2557);
and UO_168 (O_168,N_2360,N_2469);
or UO_169 (O_169,N_2942,N_2783);
nand UO_170 (O_170,N_2521,N_2787);
or UO_171 (O_171,N_2838,N_2776);
nor UO_172 (O_172,N_2502,N_2589);
nand UO_173 (O_173,N_2767,N_2582);
and UO_174 (O_174,N_2781,N_2331);
nor UO_175 (O_175,N_2546,N_2988);
nor UO_176 (O_176,N_2718,N_2625);
or UO_177 (O_177,N_2673,N_2367);
nand UO_178 (O_178,N_2709,N_2896);
or UO_179 (O_179,N_2393,N_2668);
nor UO_180 (O_180,N_2806,N_2375);
and UO_181 (O_181,N_2869,N_2372);
and UO_182 (O_182,N_2419,N_2483);
or UO_183 (O_183,N_2952,N_2716);
or UO_184 (O_184,N_2933,N_2955);
and UO_185 (O_185,N_2539,N_2937);
and UO_186 (O_186,N_2583,N_2435);
or UO_187 (O_187,N_2631,N_2335);
or UO_188 (O_188,N_2388,N_2757);
or UO_189 (O_189,N_2771,N_2819);
nand UO_190 (O_190,N_2851,N_2770);
nor UO_191 (O_191,N_2950,N_2568);
and UO_192 (O_192,N_2252,N_2962);
or UO_193 (O_193,N_2913,N_2671);
xor UO_194 (O_194,N_2301,N_2879);
or UO_195 (O_195,N_2611,N_2794);
or UO_196 (O_196,N_2396,N_2659);
nand UO_197 (O_197,N_2389,N_2588);
nor UO_198 (O_198,N_2968,N_2477);
and UO_199 (O_199,N_2427,N_2538);
and UO_200 (O_200,N_2574,N_2636);
and UO_201 (O_201,N_2873,N_2800);
nor UO_202 (O_202,N_2749,N_2501);
and UO_203 (O_203,N_2883,N_2675);
or UO_204 (O_204,N_2662,N_2795);
or UO_205 (O_205,N_2333,N_2315);
or UO_206 (O_206,N_2533,N_2730);
or UO_207 (O_207,N_2936,N_2799);
and UO_208 (O_208,N_2264,N_2825);
nor UO_209 (O_209,N_2623,N_2682);
nand UO_210 (O_210,N_2746,N_2940);
or UO_211 (O_211,N_2592,N_2304);
and UO_212 (O_212,N_2756,N_2712);
nand UO_213 (O_213,N_2612,N_2509);
nand UO_214 (O_214,N_2914,N_2856);
nand UO_215 (O_215,N_2805,N_2661);
nand UO_216 (O_216,N_2551,N_2751);
nand UO_217 (O_217,N_2945,N_2644);
nor UO_218 (O_218,N_2453,N_2406);
nand UO_219 (O_219,N_2399,N_2645);
nand UO_220 (O_220,N_2820,N_2804);
nor UO_221 (O_221,N_2357,N_2391);
or UO_222 (O_222,N_2813,N_2505);
nand UO_223 (O_223,N_2324,N_2342);
nor UO_224 (O_224,N_2801,N_2417);
nor UO_225 (O_225,N_2810,N_2259);
or UO_226 (O_226,N_2616,N_2609);
nor UO_227 (O_227,N_2277,N_2630);
and UO_228 (O_228,N_2681,N_2978);
and UO_229 (O_229,N_2982,N_2993);
nand UO_230 (O_230,N_2356,N_2516);
or UO_231 (O_231,N_2507,N_2524);
nor UO_232 (O_232,N_2361,N_2796);
and UO_233 (O_233,N_2341,N_2494);
nor UO_234 (O_234,N_2434,N_2300);
and UO_235 (O_235,N_2862,N_2977);
nand UO_236 (O_236,N_2990,N_2887);
or UO_237 (O_237,N_2344,N_2291);
and UO_238 (O_238,N_2850,N_2811);
or UO_239 (O_239,N_2745,N_2809);
nor UO_240 (O_240,N_2299,N_2877);
or UO_241 (O_241,N_2808,N_2964);
nor UO_242 (O_242,N_2271,N_2698);
nand UO_243 (O_243,N_2459,N_2510);
or UO_244 (O_244,N_2836,N_2768);
and UO_245 (O_245,N_2285,N_2663);
or UO_246 (O_246,N_2323,N_2566);
and UO_247 (O_247,N_2571,N_2416);
nor UO_248 (O_248,N_2904,N_2959);
and UO_249 (O_249,N_2986,N_2920);
and UO_250 (O_250,N_2279,N_2646);
nor UO_251 (O_251,N_2338,N_2613);
xnor UO_252 (O_252,N_2281,N_2641);
xnor UO_253 (O_253,N_2678,N_2910);
or UO_254 (O_254,N_2482,N_2431);
nor UO_255 (O_255,N_2971,N_2684);
and UO_256 (O_256,N_2400,N_2522);
and UO_257 (O_257,N_2328,N_2276);
and UO_258 (O_258,N_2506,N_2514);
nand UO_259 (O_259,N_2789,N_2983);
or UO_260 (O_260,N_2475,N_2792);
and UO_261 (O_261,N_2778,N_2346);
or UO_262 (O_262,N_2610,N_2900);
or UO_263 (O_263,N_2284,N_2818);
nor UO_264 (O_264,N_2455,N_2503);
nor UO_265 (O_265,N_2912,N_2317);
and UO_266 (O_266,N_2321,N_2628);
and UO_267 (O_267,N_2275,N_2253);
nor UO_268 (O_268,N_2298,N_2765);
or UO_269 (O_269,N_2600,N_2926);
nor UO_270 (O_270,N_2377,N_2552);
nor UO_271 (O_271,N_2547,N_2927);
or UO_272 (O_272,N_2430,N_2907);
and UO_273 (O_273,N_2939,N_2578);
or UO_274 (O_274,N_2929,N_2251);
nand UO_275 (O_275,N_2424,N_2975);
nand UO_276 (O_276,N_2380,N_2465);
or UO_277 (O_277,N_2484,N_2561);
or UO_278 (O_278,N_2604,N_2370);
and UO_279 (O_279,N_2454,N_2325);
or UO_280 (O_280,N_2327,N_2408);
nor UO_281 (O_281,N_2928,N_2468);
and UO_282 (O_282,N_2638,N_2366);
nor UO_283 (O_283,N_2382,N_2930);
and UO_284 (O_284,N_2911,N_2938);
nor UO_285 (O_285,N_2985,N_2882);
and UO_286 (O_286,N_2570,N_2831);
or UO_287 (O_287,N_2614,N_2793);
nor UO_288 (O_288,N_2827,N_2394);
or UO_289 (O_289,N_2385,N_2286);
or UO_290 (O_290,N_2753,N_2267);
nor UO_291 (O_291,N_2308,N_2656);
nor UO_292 (O_292,N_2744,N_2504);
or UO_293 (O_293,N_2548,N_2840);
xor UO_294 (O_294,N_2581,N_2957);
nand UO_295 (O_295,N_2650,N_2667);
and UO_296 (O_296,N_2349,N_2541);
nand UO_297 (O_297,N_2861,N_2726);
nor UO_298 (O_298,N_2525,N_2486);
nand UO_299 (O_299,N_2397,N_2723);
and UO_300 (O_300,N_2268,N_2705);
nor UO_301 (O_301,N_2979,N_2864);
or UO_302 (O_302,N_2915,N_2821);
nor UO_303 (O_303,N_2496,N_2748);
nor UO_304 (O_304,N_2908,N_2347);
and UO_305 (O_305,N_2436,N_2627);
nand UO_306 (O_306,N_2735,N_2495);
and UO_307 (O_307,N_2371,N_2528);
xnor UO_308 (O_308,N_2815,N_2991);
nor UO_309 (O_309,N_2620,N_2660);
and UO_310 (O_310,N_2633,N_2500);
nand UO_311 (O_311,N_2823,N_2634);
nor UO_312 (O_312,N_2293,N_2493);
nor UO_313 (O_313,N_2487,N_2888);
nand UO_314 (O_314,N_2701,N_2429);
nand UO_315 (O_315,N_2670,N_2853);
nand UO_316 (O_316,N_2981,N_2812);
and UO_317 (O_317,N_2715,N_2724);
nor UO_318 (O_318,N_2595,N_2987);
nand UO_319 (O_319,N_2754,N_2902);
or UO_320 (O_320,N_2531,N_2739);
or UO_321 (O_321,N_2414,N_2608);
or UO_322 (O_322,N_2527,N_2599);
or UO_323 (O_323,N_2451,N_2874);
and UO_324 (O_324,N_2498,N_2403);
and UO_325 (O_325,N_2535,N_2657);
or UO_326 (O_326,N_2948,N_2837);
nor UO_327 (O_327,N_2316,N_2721);
nor UO_328 (O_328,N_2885,N_2658);
nor UO_329 (O_329,N_2699,N_2485);
nor UO_330 (O_330,N_2292,N_2766);
nor UO_331 (O_331,N_2296,N_2759);
and UO_332 (O_332,N_2655,N_2624);
and UO_333 (O_333,N_2354,N_2265);
or UO_334 (O_334,N_2523,N_2567);
nor UO_335 (O_335,N_2822,N_2835);
and UO_336 (O_336,N_2731,N_2526);
nor UO_337 (O_337,N_2859,N_2847);
or UO_338 (O_338,N_2839,N_2544);
or UO_339 (O_339,N_2834,N_2700);
and UO_340 (O_340,N_2447,N_2542);
or UO_341 (O_341,N_2287,N_2458);
nand UO_342 (O_342,N_2579,N_2530);
nand UO_343 (O_343,N_2917,N_2893);
and UO_344 (O_344,N_2703,N_2302);
or UO_345 (O_345,N_2779,N_2924);
nand UO_346 (O_346,N_2511,N_2720);
and UO_347 (O_347,N_2786,N_2598);
nor UO_348 (O_348,N_2807,N_2878);
or UO_349 (O_349,N_2899,N_2972);
or UO_350 (O_350,N_2895,N_2845);
or UO_351 (O_351,N_2257,N_2679);
nor UO_352 (O_352,N_2345,N_2629);
nor UO_353 (O_353,N_2683,N_2967);
and UO_354 (O_354,N_2319,N_2556);
and UO_355 (O_355,N_2273,N_2369);
or UO_356 (O_356,N_2632,N_2594);
and UO_357 (O_357,N_2481,N_2379);
nor UO_358 (O_358,N_2340,N_2984);
or UO_359 (O_359,N_2642,N_2383);
or UO_360 (O_360,N_2843,N_2760);
or UO_361 (O_361,N_2555,N_2707);
nor UO_362 (O_362,N_2989,N_2648);
xnor UO_363 (O_363,N_2706,N_2742);
nor UO_364 (O_364,N_2310,N_2814);
nand UO_365 (O_365,N_2775,N_2694);
nand UO_366 (O_366,N_2923,N_2480);
or UO_367 (O_367,N_2550,N_2736);
nand UO_368 (O_368,N_2702,N_2894);
nand UO_369 (O_369,N_2898,N_2994);
nand UO_370 (O_370,N_2692,N_2282);
nand UO_371 (O_371,N_2857,N_2460);
nor UO_372 (O_372,N_2467,N_2365);
nand UO_373 (O_373,N_2529,N_2637);
nand UO_374 (O_374,N_2413,N_2752);
nor UO_375 (O_375,N_2314,N_2733);
nand UO_376 (O_376,N_2657,N_2485);
nor UO_377 (O_377,N_2782,N_2489);
nand UO_378 (O_378,N_2398,N_2871);
or UO_379 (O_379,N_2785,N_2539);
nor UO_380 (O_380,N_2623,N_2362);
nand UO_381 (O_381,N_2602,N_2771);
nor UO_382 (O_382,N_2312,N_2887);
nand UO_383 (O_383,N_2614,N_2319);
nor UO_384 (O_384,N_2463,N_2412);
and UO_385 (O_385,N_2929,N_2687);
nor UO_386 (O_386,N_2494,N_2726);
nor UO_387 (O_387,N_2368,N_2817);
and UO_388 (O_388,N_2747,N_2513);
or UO_389 (O_389,N_2555,N_2824);
nand UO_390 (O_390,N_2559,N_2991);
nor UO_391 (O_391,N_2465,N_2403);
or UO_392 (O_392,N_2784,N_2760);
nand UO_393 (O_393,N_2456,N_2251);
nand UO_394 (O_394,N_2702,N_2626);
nor UO_395 (O_395,N_2792,N_2819);
and UO_396 (O_396,N_2809,N_2617);
nor UO_397 (O_397,N_2348,N_2394);
or UO_398 (O_398,N_2998,N_2638);
nor UO_399 (O_399,N_2963,N_2780);
nor UO_400 (O_400,N_2302,N_2832);
or UO_401 (O_401,N_2796,N_2273);
nand UO_402 (O_402,N_2386,N_2924);
nand UO_403 (O_403,N_2796,N_2397);
or UO_404 (O_404,N_2309,N_2433);
or UO_405 (O_405,N_2373,N_2312);
or UO_406 (O_406,N_2815,N_2287);
nand UO_407 (O_407,N_2781,N_2913);
nand UO_408 (O_408,N_2666,N_2556);
nor UO_409 (O_409,N_2566,N_2337);
nor UO_410 (O_410,N_2792,N_2590);
or UO_411 (O_411,N_2931,N_2623);
nand UO_412 (O_412,N_2726,N_2625);
or UO_413 (O_413,N_2783,N_2994);
and UO_414 (O_414,N_2807,N_2829);
nor UO_415 (O_415,N_2653,N_2817);
or UO_416 (O_416,N_2345,N_2599);
nor UO_417 (O_417,N_2536,N_2648);
or UO_418 (O_418,N_2285,N_2771);
nand UO_419 (O_419,N_2417,N_2348);
and UO_420 (O_420,N_2984,N_2495);
nand UO_421 (O_421,N_2555,N_2499);
or UO_422 (O_422,N_2748,N_2376);
or UO_423 (O_423,N_2276,N_2648);
nand UO_424 (O_424,N_2352,N_2919);
or UO_425 (O_425,N_2791,N_2534);
and UO_426 (O_426,N_2453,N_2938);
nand UO_427 (O_427,N_2743,N_2527);
nand UO_428 (O_428,N_2479,N_2582);
nor UO_429 (O_429,N_2291,N_2447);
nor UO_430 (O_430,N_2382,N_2973);
or UO_431 (O_431,N_2321,N_2749);
xor UO_432 (O_432,N_2918,N_2749);
and UO_433 (O_433,N_2724,N_2458);
nor UO_434 (O_434,N_2924,N_2780);
nand UO_435 (O_435,N_2743,N_2687);
and UO_436 (O_436,N_2828,N_2540);
nand UO_437 (O_437,N_2713,N_2520);
nor UO_438 (O_438,N_2538,N_2835);
and UO_439 (O_439,N_2584,N_2509);
nor UO_440 (O_440,N_2655,N_2916);
nor UO_441 (O_441,N_2330,N_2545);
nor UO_442 (O_442,N_2947,N_2708);
nor UO_443 (O_443,N_2851,N_2306);
and UO_444 (O_444,N_2805,N_2601);
or UO_445 (O_445,N_2960,N_2752);
nor UO_446 (O_446,N_2593,N_2858);
and UO_447 (O_447,N_2510,N_2533);
or UO_448 (O_448,N_2774,N_2691);
or UO_449 (O_449,N_2441,N_2706);
or UO_450 (O_450,N_2938,N_2653);
nand UO_451 (O_451,N_2851,N_2748);
and UO_452 (O_452,N_2374,N_2922);
nor UO_453 (O_453,N_2842,N_2637);
nand UO_454 (O_454,N_2339,N_2687);
nor UO_455 (O_455,N_2520,N_2538);
nand UO_456 (O_456,N_2842,N_2697);
nand UO_457 (O_457,N_2285,N_2506);
nand UO_458 (O_458,N_2983,N_2777);
nand UO_459 (O_459,N_2315,N_2493);
or UO_460 (O_460,N_2456,N_2919);
nor UO_461 (O_461,N_2449,N_2859);
and UO_462 (O_462,N_2944,N_2916);
and UO_463 (O_463,N_2983,N_2521);
nor UO_464 (O_464,N_2265,N_2356);
or UO_465 (O_465,N_2533,N_2841);
nor UO_466 (O_466,N_2726,N_2964);
nand UO_467 (O_467,N_2504,N_2734);
and UO_468 (O_468,N_2252,N_2989);
nor UO_469 (O_469,N_2639,N_2559);
and UO_470 (O_470,N_2553,N_2901);
and UO_471 (O_471,N_2690,N_2758);
or UO_472 (O_472,N_2848,N_2874);
and UO_473 (O_473,N_2270,N_2381);
nor UO_474 (O_474,N_2811,N_2986);
nand UO_475 (O_475,N_2528,N_2327);
nor UO_476 (O_476,N_2570,N_2753);
or UO_477 (O_477,N_2537,N_2662);
and UO_478 (O_478,N_2808,N_2862);
nand UO_479 (O_479,N_2942,N_2301);
nand UO_480 (O_480,N_2580,N_2801);
nor UO_481 (O_481,N_2606,N_2359);
nor UO_482 (O_482,N_2618,N_2933);
nand UO_483 (O_483,N_2923,N_2973);
nand UO_484 (O_484,N_2503,N_2308);
or UO_485 (O_485,N_2691,N_2280);
or UO_486 (O_486,N_2681,N_2353);
and UO_487 (O_487,N_2507,N_2775);
nor UO_488 (O_488,N_2410,N_2576);
or UO_489 (O_489,N_2432,N_2746);
nor UO_490 (O_490,N_2696,N_2734);
and UO_491 (O_491,N_2983,N_2751);
nand UO_492 (O_492,N_2454,N_2315);
nand UO_493 (O_493,N_2532,N_2950);
nand UO_494 (O_494,N_2392,N_2696);
or UO_495 (O_495,N_2479,N_2258);
nor UO_496 (O_496,N_2546,N_2663);
and UO_497 (O_497,N_2772,N_2655);
nand UO_498 (O_498,N_2675,N_2831);
and UO_499 (O_499,N_2379,N_2354);
endmodule