module basic_2500_25000_3000_4_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18762,N_18763,N_18764,N_18765,N_18766,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18792,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18880,N_18881,N_18882,N_18883,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18900,N_18901,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18912,N_18913,N_18914,N_18915,N_18916,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19305,N_19306,N_19307,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20291,N_20292,N_20294,N_20295,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20372,N_20373,N_20374,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20622,N_20624,N_20625,N_20626,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20652,N_20653,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20906,N_20907,N_20908,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20925,N_20926,N_20927,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20983,N_20984,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21081,N_21082,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21119,N_21120,N_21121,N_21122,N_21123,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21429,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21465,N_21466,N_21467,N_21469,N_21470,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21514,N_21515,N_21516,N_21517,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21599,N_21600,N_21601,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21767,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21903,N_21904,N_21905,N_21907,N_21908,N_21910,N_21911,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22031,N_22032,N_22033,N_22034,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22058,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22287,N_22288,N_22289,N_22290,N_22291,N_22293,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22358,N_22359,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22507,N_22508,N_22509,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22741,N_22742,N_22743,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22941,N_22942,N_22943,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23010,N_23011,N_23012,N_23013,N_23014,N_23016,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23028,N_23029,N_23030,N_23031,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23331,N_23332,N_23333,N_23334,N_23335,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23717,N_23718,N_23719,N_23720,N_23721,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24046,N_24047,N_24049,N_24050,N_24051,N_24052,N_24053,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24081,N_24082,N_24083,N_24084,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24141,N_24142,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24201,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24247,N_24248,N_24249,N_24250,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24478,N_24479,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24497,N_24498,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24607,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24680,N_24681,N_24682,N_24683,N_24684,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xor U0 (N_0,In_2207,In_323);
nor U1 (N_1,In_1485,In_1959);
or U2 (N_2,In_256,In_1208);
nand U3 (N_3,In_2063,In_1417);
and U4 (N_4,In_22,In_129);
nand U5 (N_5,In_1712,In_602);
nor U6 (N_6,In_1669,In_1963);
nor U7 (N_7,In_2342,In_50);
nor U8 (N_8,In_1345,In_2005);
nand U9 (N_9,In_1369,In_725);
and U10 (N_10,In_993,In_1135);
nor U11 (N_11,In_2286,In_18);
nor U12 (N_12,In_1326,In_879);
nor U13 (N_13,In_983,In_1764);
or U14 (N_14,In_20,In_1153);
and U15 (N_15,In_1616,In_2493);
and U16 (N_16,In_2235,In_223);
and U17 (N_17,In_2231,In_330);
nand U18 (N_18,In_1930,In_2153);
or U19 (N_19,In_787,In_529);
and U20 (N_20,In_101,In_2211);
or U21 (N_21,In_2155,In_2440);
and U22 (N_22,In_1978,In_468);
and U23 (N_23,In_41,In_754);
or U24 (N_24,In_2484,In_1638);
or U25 (N_25,In_2255,In_564);
nor U26 (N_26,In_1387,In_2393);
or U27 (N_27,In_1565,In_1335);
and U28 (N_28,In_945,In_583);
or U29 (N_29,In_1294,In_181);
and U30 (N_30,In_1200,In_1632);
nor U31 (N_31,In_453,In_131);
and U32 (N_32,In_203,In_2452);
nor U33 (N_33,In_2001,In_2379);
and U34 (N_34,In_506,In_627);
nand U35 (N_35,In_385,In_883);
xnor U36 (N_36,In_1261,In_1242);
nand U37 (N_37,In_1173,In_773);
and U38 (N_38,In_1272,In_804);
nor U39 (N_39,In_1503,In_1745);
nor U40 (N_40,In_2449,In_1831);
or U41 (N_41,In_1996,In_1218);
nand U42 (N_42,In_167,In_1196);
nor U43 (N_43,In_2076,In_1702);
and U44 (N_44,In_1327,In_1923);
and U45 (N_45,In_705,In_116);
nand U46 (N_46,In_169,In_1970);
nand U47 (N_47,In_941,In_2218);
or U48 (N_48,In_1328,In_2145);
or U49 (N_49,In_278,In_1176);
nand U50 (N_50,In_1062,In_1673);
or U51 (N_51,In_26,In_1846);
and U52 (N_52,In_596,In_793);
xor U53 (N_53,In_340,In_629);
and U54 (N_54,In_2366,In_2085);
or U55 (N_55,In_1756,In_1136);
and U56 (N_56,In_368,In_2309);
nand U57 (N_57,In_2217,In_914);
xor U58 (N_58,In_1641,In_1661);
or U59 (N_59,In_1587,In_837);
nand U60 (N_60,In_708,In_1410);
or U61 (N_61,In_523,In_626);
or U62 (N_62,In_461,In_2400);
or U63 (N_63,In_652,In_1432);
and U64 (N_64,In_333,In_1812);
nand U65 (N_65,In_933,In_1896);
or U66 (N_66,In_1672,In_2428);
and U67 (N_67,In_2310,In_1227);
nand U68 (N_68,In_864,In_1446);
nor U69 (N_69,In_1469,In_1161);
nand U70 (N_70,In_1449,In_2474);
nand U71 (N_71,In_2131,In_1620);
xnor U72 (N_72,In_1310,In_1518);
or U73 (N_73,In_1308,In_1311);
and U74 (N_74,In_519,In_528);
nor U75 (N_75,In_2156,In_1053);
nand U76 (N_76,In_1857,In_1194);
nand U77 (N_77,In_294,In_1826);
and U78 (N_78,In_2159,In_613);
or U79 (N_79,In_2042,In_70);
or U80 (N_80,In_2105,In_625);
or U81 (N_81,In_1928,In_406);
nor U82 (N_82,In_2160,In_778);
and U83 (N_83,In_2234,In_1052);
nand U84 (N_84,In_1341,In_1849);
and U85 (N_85,In_2083,In_1146);
nand U86 (N_86,In_2441,In_25);
and U87 (N_87,In_1119,In_263);
nand U88 (N_88,In_462,In_232);
xnor U89 (N_89,In_1521,In_1213);
or U90 (N_90,In_207,In_1944);
nand U91 (N_91,In_320,In_541);
and U92 (N_92,In_222,In_634);
xor U93 (N_93,In_89,In_721);
and U94 (N_94,In_1393,In_2210);
nor U95 (N_95,In_2346,In_766);
and U96 (N_96,In_1258,In_433);
and U97 (N_97,In_936,In_130);
xor U98 (N_98,In_2205,In_1398);
nor U99 (N_99,In_316,In_862);
nand U100 (N_100,In_2271,In_2321);
and U101 (N_101,In_473,In_439);
nor U102 (N_102,In_1350,In_2443);
nor U103 (N_103,In_1654,In_1734);
nor U104 (N_104,In_1291,In_1151);
and U105 (N_105,In_1754,In_71);
xor U106 (N_106,In_146,In_2254);
or U107 (N_107,In_1753,In_1142);
nor U108 (N_108,In_145,In_1428);
or U109 (N_109,In_1694,In_2361);
or U110 (N_110,In_1732,In_2);
and U111 (N_111,In_1199,In_2143);
and U112 (N_112,In_1799,In_405);
xor U113 (N_113,In_1837,In_1663);
or U114 (N_114,In_180,In_758);
nand U115 (N_115,In_2092,In_859);
nor U116 (N_116,In_243,In_603);
nand U117 (N_117,In_952,In_2483);
nor U118 (N_118,In_2311,In_1969);
nor U119 (N_119,In_731,In_1402);
and U120 (N_120,In_2209,In_1080);
and U121 (N_121,In_2223,In_1739);
and U122 (N_122,In_1539,In_698);
nand U123 (N_123,In_2436,In_975);
nor U124 (N_124,In_2185,In_2038);
nor U125 (N_125,In_867,In_2340);
and U126 (N_126,In_709,In_2370);
xnor U127 (N_127,In_561,In_678);
or U128 (N_128,In_1459,In_2178);
or U129 (N_129,In_356,In_2448);
nand U130 (N_130,In_1643,In_769);
nand U131 (N_131,In_514,In_2335);
and U132 (N_132,In_925,In_2396);
nand U133 (N_133,In_1595,In_503);
nor U134 (N_134,In_639,In_821);
or U135 (N_135,In_444,In_432);
nor U136 (N_136,In_1755,In_296);
nor U137 (N_137,In_1475,In_13);
nor U138 (N_138,In_46,In_1263);
and U139 (N_139,In_1675,In_1365);
or U140 (N_140,In_1180,In_408);
nor U141 (N_141,In_1337,In_969);
nand U142 (N_142,In_204,In_1735);
and U143 (N_143,In_1909,In_1319);
or U144 (N_144,In_1808,In_1660);
or U145 (N_145,In_2055,In_252);
nor U146 (N_146,In_502,In_2064);
or U147 (N_147,In_1132,In_112);
nor U148 (N_148,In_72,In_2377);
and U149 (N_149,In_85,In_1137);
and U150 (N_150,In_2058,In_746);
nor U151 (N_151,In_2432,In_1901);
nor U152 (N_152,In_2051,In_1193);
nand U153 (N_153,In_1113,In_1079);
or U154 (N_154,In_2439,In_803);
xnor U155 (N_155,In_2142,In_446);
nand U156 (N_156,In_1279,In_2166);
or U157 (N_157,In_1942,In_2025);
nand U158 (N_158,In_664,In_637);
or U159 (N_159,In_137,In_1768);
nor U160 (N_160,In_1803,In_249);
xnor U161 (N_161,In_2380,In_756);
or U162 (N_162,In_1219,In_2315);
xor U163 (N_163,In_687,In_1339);
nand U164 (N_164,In_404,In_1430);
or U165 (N_165,In_2481,In_1298);
xnor U166 (N_166,In_796,In_812);
and U167 (N_167,In_2442,In_1315);
nor U168 (N_168,In_753,In_866);
and U169 (N_169,In_1815,In_479);
xnor U170 (N_170,In_858,In_834);
nor U171 (N_171,In_1234,In_1711);
or U172 (N_172,In_92,In_31);
nor U173 (N_173,In_82,In_492);
and U174 (N_174,In_1461,In_1236);
nor U175 (N_175,In_464,In_122);
nor U176 (N_176,In_710,In_621);
nand U177 (N_177,In_1886,In_411);
nand U178 (N_178,In_811,In_465);
and U179 (N_179,In_559,In_2308);
nand U180 (N_180,In_1718,In_1635);
nand U181 (N_181,In_818,In_782);
or U182 (N_182,In_1491,In_1481);
nor U183 (N_183,In_305,In_279);
nor U184 (N_184,In_2415,In_1256);
nor U185 (N_185,In_655,In_1650);
or U186 (N_186,In_1851,In_1697);
and U187 (N_187,In_1127,In_2041);
nor U188 (N_188,In_1588,In_1374);
nor U189 (N_189,In_152,In_1828);
nand U190 (N_190,In_805,In_427);
nand U191 (N_191,In_2067,In_1577);
xor U192 (N_192,In_727,In_186);
and U193 (N_193,In_1947,In_2093);
or U194 (N_194,In_1434,In_23);
or U195 (N_195,In_2086,In_807);
nand U196 (N_196,In_121,In_438);
nand U197 (N_197,In_1332,In_2435);
nor U198 (N_198,In_1555,In_1174);
nand U199 (N_199,In_174,In_1708);
or U200 (N_200,In_2123,In_600);
nor U201 (N_201,In_2100,In_1715);
or U202 (N_202,In_2456,In_2398);
or U203 (N_203,In_1414,In_929);
or U204 (N_204,In_358,In_269);
nand U205 (N_205,In_170,In_2296);
or U206 (N_206,In_1,In_1346);
or U207 (N_207,In_1513,In_1203);
nor U208 (N_208,In_2192,In_164);
or U209 (N_209,In_212,In_1128);
nand U210 (N_210,In_1592,In_934);
or U211 (N_211,In_965,In_845);
nand U212 (N_212,In_2183,In_836);
nor U213 (N_213,In_1101,In_744);
and U214 (N_214,In_497,In_1703);
and U215 (N_215,In_1019,In_1184);
nor U216 (N_216,In_672,In_1950);
and U217 (N_217,In_605,In_1625);
nand U218 (N_218,In_1240,In_620);
nand U219 (N_219,In_706,In_293);
or U220 (N_220,In_329,In_2478);
nand U221 (N_221,In_1017,In_2165);
nor U222 (N_222,In_1925,In_877);
or U223 (N_223,In_2035,In_403);
xnor U224 (N_224,In_2097,In_2490);
or U225 (N_225,In_317,In_1902);
or U226 (N_226,In_17,In_3);
xor U227 (N_227,In_2181,In_1992);
and U228 (N_228,In_258,In_915);
nand U229 (N_229,In_2230,In_2292);
nor U230 (N_230,In_1811,In_874);
nand U231 (N_231,In_703,In_48);
and U232 (N_232,In_2199,In_846);
nor U233 (N_233,In_1500,In_1465);
nand U234 (N_234,In_91,In_376);
or U235 (N_235,In_1576,In_885);
or U236 (N_236,In_1380,In_1510);
nand U237 (N_237,In_2251,In_65);
xor U238 (N_238,In_1309,In_1351);
or U239 (N_239,In_1771,In_2162);
nand U240 (N_240,In_233,In_1425);
and U241 (N_241,In_1550,In_802);
and U242 (N_242,In_1162,In_2233);
or U243 (N_243,In_1467,In_1452);
nor U244 (N_244,In_1788,In_873);
or U245 (N_245,In_1888,In_570);
xnor U246 (N_246,In_36,In_1334);
and U247 (N_247,In_496,In_1704);
and U248 (N_248,In_1069,In_113);
and U249 (N_249,In_2082,In_300);
nor U250 (N_250,In_1571,In_2019);
nor U251 (N_251,In_1323,In_2045);
nor U252 (N_252,In_280,In_264);
and U253 (N_253,In_2206,In_1878);
nand U254 (N_254,In_1418,In_1295);
nor U255 (N_255,In_2349,In_2334);
nand U256 (N_256,In_225,In_370);
and U257 (N_257,In_1235,In_2161);
and U258 (N_258,In_1482,In_978);
and U259 (N_259,In_262,In_474);
and U260 (N_260,In_282,In_824);
nand U261 (N_261,In_610,In_1889);
and U262 (N_262,In_1985,In_374);
or U263 (N_263,In_536,In_1233);
nor U264 (N_264,In_1847,In_2194);
nand U265 (N_265,In_2466,In_1264);
xor U266 (N_266,In_799,In_1383);
nor U267 (N_267,In_1986,In_110);
or U268 (N_268,In_53,In_500);
and U269 (N_269,In_253,In_2017);
nand U270 (N_270,In_2354,In_882);
xor U271 (N_271,In_1361,In_1832);
and U272 (N_272,In_7,In_1931);
or U273 (N_273,In_960,In_2214);
and U274 (N_274,In_2262,In_1834);
or U275 (N_275,In_545,In_775);
nor U276 (N_276,In_304,In_261);
nor U277 (N_277,In_2227,In_1867);
nand U278 (N_278,In_1445,In_2498);
xor U279 (N_279,In_861,In_44);
and U280 (N_280,In_1552,In_448);
nor U281 (N_281,In_1584,In_688);
nand U282 (N_282,In_2355,In_127);
nand U283 (N_283,In_2167,In_1605);
nor U284 (N_284,In_825,In_2429);
or U285 (N_285,In_118,In_547);
xor U286 (N_286,In_1125,In_1746);
and U287 (N_287,In_1979,In_902);
nand U288 (N_288,In_173,In_1906);
xor U289 (N_289,In_1809,In_1188);
nor U290 (N_290,In_1793,In_1453);
nand U291 (N_291,In_1050,In_913);
or U292 (N_292,In_1827,In_40);
nand U293 (N_293,In_641,In_1864);
xor U294 (N_294,In_1581,In_1438);
nor U295 (N_295,In_257,In_2208);
and U296 (N_296,In_2290,In_1435);
or U297 (N_297,In_593,In_2002);
xnor U298 (N_298,In_1223,In_328);
or U299 (N_299,In_1594,In_714);
xnor U300 (N_300,In_900,In_2070);
nand U301 (N_301,In_1010,In_1046);
and U302 (N_302,In_1385,In_585);
or U303 (N_303,In_996,In_2032);
and U304 (N_304,In_842,In_1564);
or U305 (N_305,In_2148,In_2327);
nor U306 (N_306,In_1658,In_379);
nand U307 (N_307,In_322,In_240);
nand U308 (N_308,In_1706,In_2284);
nor U309 (N_309,In_831,In_1621);
nor U310 (N_310,In_504,In_1843);
nor U311 (N_311,In_2147,In_2226);
and U312 (N_312,In_601,In_1879);
or U313 (N_313,In_926,In_211);
nand U314 (N_314,In_2149,In_277);
or U315 (N_315,In_1110,In_2399);
and U316 (N_316,In_1772,In_2191);
or U317 (N_317,In_604,In_387);
nand U318 (N_318,In_633,In_309);
nor U319 (N_319,In_1532,In_380);
or U320 (N_320,In_1089,In_1454);
nor U321 (N_321,In_162,In_2491);
or U322 (N_322,In_676,In_924);
or U323 (N_323,In_467,In_1767);
nand U324 (N_324,In_303,In_909);
nor U325 (N_325,In_381,In_1529);
nand U326 (N_326,In_1579,In_2353);
nor U327 (N_327,In_1519,In_2128);
nor U328 (N_328,In_197,In_631);
or U329 (N_329,In_1290,In_2004);
nor U330 (N_330,In_580,In_1059);
xnor U331 (N_331,In_265,In_1591);
or U332 (N_332,In_970,In_1817);
or U333 (N_333,In_813,In_510);
or U334 (N_334,In_1104,In_2479);
xnor U335 (N_335,In_1822,In_1456);
nor U336 (N_336,In_2472,In_171);
xor U337 (N_337,In_193,In_729);
nor U338 (N_338,In_1025,In_1829);
nand U339 (N_339,In_533,In_2305);
or U340 (N_340,In_1224,In_2318);
nor U341 (N_341,In_1656,In_2107);
and U342 (N_342,In_1984,In_937);
nor U343 (N_343,In_635,In_272);
nand U344 (N_344,In_154,In_1171);
and U345 (N_345,In_1064,In_1504);
nor U346 (N_346,In_235,In_2467);
and U347 (N_347,In_1841,In_1823);
or U348 (N_348,In_283,In_1685);
nand U349 (N_349,In_2261,In_314);
or U350 (N_350,In_1399,In_431);
or U351 (N_351,In_2278,In_1450);
and U352 (N_352,In_1508,In_2280);
or U353 (N_353,In_1566,In_981);
or U354 (N_354,In_77,In_1042);
nor U355 (N_355,In_1018,In_1876);
nand U356 (N_356,In_125,In_1389);
or U357 (N_357,In_1786,In_1700);
nor U358 (N_358,In_1277,In_511);
nor U359 (N_359,In_597,In_1789);
nor U360 (N_360,In_117,In_1964);
nand U361 (N_361,In_1617,In_979);
nor U362 (N_362,In_142,In_2302);
or U363 (N_363,In_1557,In_1805);
or U364 (N_364,In_572,In_2499);
or U365 (N_365,In_1282,In_1614);
nand U366 (N_366,In_1593,In_1763);
or U367 (N_367,In_66,In_2259);
and U368 (N_368,In_1000,In_1514);
and U369 (N_369,In_2324,In_365);
and U370 (N_370,In_1994,In_1253);
and U371 (N_371,In_415,In_1918);
nor U372 (N_372,In_1216,In_976);
and U373 (N_373,In_538,In_1693);
or U374 (N_374,In_228,In_1894);
or U375 (N_375,In_1861,In_704);
nand U376 (N_376,In_96,In_400);
nand U377 (N_377,In_904,In_1349);
nor U378 (N_378,In_720,In_1589);
nor U379 (N_379,In_241,In_1709);
and U380 (N_380,In_977,In_220);
nand U381 (N_381,In_1765,In_16);
xor U382 (N_382,In_1273,In_1073);
or U383 (N_383,In_1109,In_2113);
nand U384 (N_384,In_617,In_2071);
nand U385 (N_385,In_1076,In_1117);
or U386 (N_386,In_743,In_1897);
and U387 (N_387,In_1416,In_1687);
xor U388 (N_388,In_916,In_2464);
nand U389 (N_389,In_987,In_692);
and U390 (N_390,In_206,In_1980);
or U391 (N_391,In_668,In_336);
nor U392 (N_392,In_417,In_890);
and U393 (N_393,In_2426,In_1221);
nor U394 (N_394,In_569,In_2133);
nor U395 (N_395,In_1848,In_1628);
and U396 (N_396,In_2222,In_1280);
and U397 (N_397,In_875,In_0);
xor U398 (N_398,In_1382,In_1795);
and U399 (N_399,In_2312,In_147);
nor U400 (N_400,In_394,In_1478);
and U401 (N_401,In_1265,In_1773);
or U402 (N_402,In_281,In_2084);
or U403 (N_403,In_650,In_1856);
and U404 (N_404,In_449,In_1197);
or U405 (N_405,In_2108,In_42);
xor U406 (N_406,In_2263,In_224);
and U407 (N_407,In_1744,In_2291);
or U408 (N_408,In_2368,In_966);
nand U409 (N_409,In_350,In_1705);
or U410 (N_410,In_591,In_190);
nand U411 (N_411,In_521,In_565);
or U412 (N_412,In_184,In_34);
and U413 (N_413,In_99,In_435);
nand U414 (N_414,In_1204,In_414);
or U415 (N_415,In_1781,In_499);
nand U416 (N_416,In_1926,In_209);
or U417 (N_417,In_2369,In_1289);
nor U418 (N_418,In_838,In_1126);
or U419 (N_419,In_1943,In_2492);
nor U420 (N_420,In_486,In_798);
and U421 (N_421,In_1743,In_1412);
nor U422 (N_422,In_516,In_760);
and U423 (N_423,In_313,In_1209);
and U424 (N_424,In_2106,In_1304);
nor U425 (N_425,In_741,In_2250);
nand U426 (N_426,In_1120,In_1483);
and U427 (N_427,In_2332,In_670);
nand U428 (N_428,In_1630,In_55);
nand U429 (N_429,In_1875,In_2134);
and U430 (N_430,In_1528,In_245);
nor U431 (N_431,In_1479,In_512);
nand U432 (N_432,In_1626,In_1186);
nor U433 (N_433,In_378,In_1007);
or U434 (N_434,In_1338,In_615);
nor U435 (N_435,In_1612,In_307);
xor U436 (N_436,In_986,In_391);
nand U437 (N_437,In_1946,In_1406);
xor U438 (N_438,In_643,In_1413);
nand U439 (N_439,In_1437,In_2197);
nand U440 (N_440,In_2257,In_1336);
or U441 (N_441,In_815,In_1839);
nand U442 (N_442,In_1190,In_1244);
and U443 (N_443,In_1511,In_1178);
nand U444 (N_444,In_701,In_105);
nand U445 (N_445,In_1222,In_56);
nand U446 (N_446,In_2482,In_1071);
or U447 (N_447,In_43,In_1056);
xor U448 (N_448,In_540,In_120);
nand U449 (N_449,In_2360,In_470);
and U450 (N_450,In_872,In_2187);
nor U451 (N_451,In_1855,In_1535);
and U452 (N_452,In_992,In_244);
and U453 (N_453,In_800,In_166);
xnor U454 (N_454,In_1472,In_592);
nand U455 (N_455,In_1362,In_1138);
nor U456 (N_456,In_2325,In_1377);
or U457 (N_457,In_2023,In_632);
and U458 (N_458,In_677,In_2179);
nand U459 (N_459,In_587,In_1573);
and U460 (N_460,In_1559,In_1257);
nand U461 (N_461,In_2014,In_2487);
nor U462 (N_462,In_892,In_2496);
nand U463 (N_463,In_371,In_1872);
nor U464 (N_464,In_662,In_1606);
nand U465 (N_465,In_1574,In_1551);
or U466 (N_466,In_1610,In_37);
or U467 (N_467,In_1087,In_2073);
and U468 (N_468,In_2044,In_157);
nor U469 (N_469,In_1881,In_518);
nand U470 (N_470,In_1759,In_384);
or U471 (N_471,In_1515,In_893);
xnor U472 (N_472,In_689,In_2356);
nand U473 (N_473,In_809,In_2357);
nor U474 (N_474,In_2135,In_527);
nor U475 (N_475,In_472,In_421);
or U476 (N_476,In_271,In_2411);
and U477 (N_477,In_2089,In_990);
nor U478 (N_478,In_155,In_829);
nor U479 (N_479,In_1363,In_611);
and U480 (N_480,In_1262,In_1601);
nor U481 (N_481,In_58,In_2300);
nor U482 (N_482,In_11,In_1243);
and U483 (N_483,In_624,In_686);
nand U484 (N_484,In_942,In_711);
nor U485 (N_485,In_1749,In_2126);
nor U486 (N_486,In_2028,In_1299);
nand U487 (N_487,In_2130,In_2281);
and U488 (N_488,In_172,In_2331);
xor U489 (N_489,In_2422,In_946);
and U490 (N_490,In_1466,In_483);
nand U491 (N_491,In_1534,In_188);
and U492 (N_492,In_1501,In_1664);
or U493 (N_493,In_2326,In_2406);
nand U494 (N_494,In_691,In_716);
and U495 (N_495,In_1710,In_2328);
xor U496 (N_496,In_372,In_2256);
or U497 (N_497,In_2477,In_143);
nand U498 (N_498,In_239,In_1198);
or U499 (N_499,In_2236,In_1887);
or U500 (N_500,In_1024,In_104);
or U501 (N_501,In_1157,In_2219);
nand U502 (N_502,In_2090,In_2447);
nand U503 (N_503,In_1585,In_1480);
or U504 (N_504,In_1791,In_1192);
nand U505 (N_505,In_822,In_413);
nor U506 (N_506,In_651,In_2080);
or U507 (N_507,In_780,In_988);
and U508 (N_508,In_1476,In_1689);
nor U509 (N_509,In_1536,In_1586);
nand U510 (N_510,In_828,In_1777);
nor U511 (N_511,In_679,In_869);
nand U512 (N_512,In_2260,In_1288);
nor U513 (N_513,In_1782,In_103);
nand U514 (N_514,In_562,In_2329);
nor U515 (N_515,In_2072,In_2339);
nor U516 (N_516,In_908,In_745);
and U517 (N_517,In_1624,In_1870);
or U518 (N_518,In_1520,In_1636);
nand U519 (N_519,In_1955,In_1347);
nor U520 (N_520,In_383,In_683);
xor U521 (N_521,In_1441,In_2322);
and U522 (N_522,In_680,In_1099);
xnor U523 (N_523,In_2111,In_2200);
and U524 (N_524,In_1844,In_2431);
nor U525 (N_525,In_2387,In_2094);
nand U526 (N_526,In_1956,In_826);
nor U527 (N_527,In_2104,In_2407);
xor U528 (N_528,In_2198,In_2465);
xnor U529 (N_529,In_2221,In_614);
nand U530 (N_530,In_390,In_1030);
nand U531 (N_531,In_288,In_2272);
nand U532 (N_532,In_324,In_1517);
xnor U533 (N_533,In_522,In_2119);
nand U534 (N_534,In_2253,In_1150);
xnor U535 (N_535,In_175,In_1250);
nand U536 (N_536,In_2297,In_1232);
nor U537 (N_537,In_2371,In_1684);
and U538 (N_538,In_1613,In_566);
xor U539 (N_539,In_1394,In_98);
and U540 (N_540,In_1995,In_1306);
or U541 (N_541,In_1952,In_2164);
and U542 (N_542,In_1830,In_2195);
nand U543 (N_543,In_94,In_1022);
nand U544 (N_544,In_201,In_1400);
nor U545 (N_545,In_2362,In_1381);
and U546 (N_546,In_1411,In_268);
nand U547 (N_547,In_764,In_88);
and U548 (N_548,In_1877,In_1390);
or U549 (N_549,In_424,In_254);
nand U550 (N_550,In_755,In_1471);
nand U551 (N_551,In_475,In_1769);
and U552 (N_552,In_2497,In_1143);
nand U553 (N_553,In_1760,In_546);
nand U554 (N_554,In_2203,In_568);
nor U555 (N_555,In_1429,In_1836);
nand U556 (N_556,In_2409,In_1998);
and U557 (N_557,In_1597,In_360);
and U558 (N_558,In_638,In_2184);
or U559 (N_559,In_1860,In_1558);
or U560 (N_560,In_797,In_2402);
xnor U561 (N_561,In_2129,In_1360);
nor U562 (N_562,In_237,In_1063);
nor U563 (N_563,In_2101,In_1609);
xor U564 (N_564,In_1741,In_236);
and U565 (N_565,In_747,In_1164);
and U566 (N_566,In_548,In_2015);
and U567 (N_567,In_742,In_816);
xnor U568 (N_568,In_1993,In_2420);
nor U569 (N_569,In_2390,In_375);
nand U570 (N_570,In_786,In_1238);
nor U571 (N_571,In_1049,In_1727);
or U572 (N_572,In_1252,In_1463);
and U573 (N_573,In_1737,In_1634);
or U574 (N_574,In_354,In_823);
nand U575 (N_575,In_923,In_2295);
xor U576 (N_576,In_2283,In_732);
and U577 (N_577,In_2489,In_1248);
nand U578 (N_578,In_1618,In_1651);
nor U579 (N_579,In_1800,In_337);
and U580 (N_580,In_761,In_1778);
nor U581 (N_581,In_959,In_581);
or U582 (N_582,In_1976,In_1627);
xor U583 (N_583,In_1239,In_1214);
and U584 (N_584,In_49,In_139);
nor U585 (N_585,In_1880,In_401);
nor U586 (N_586,In_1116,In_250);
nor U587 (N_587,In_2463,In_153);
or U588 (N_588,In_1733,In_2372);
nand U589 (N_589,In_1431,In_555);
nand U590 (N_590,In_1070,In_791);
nand U591 (N_591,In_69,In_2405);
nand U592 (N_592,In_801,In_2121);
and U593 (N_593,In_1991,In_1895);
nand U594 (N_594,In_1082,In_918);
nand U595 (N_595,In_1724,In_1433);
or U596 (N_596,In_213,In_1247);
or U597 (N_597,In_349,In_1134);
xnor U598 (N_598,In_215,In_657);
and U599 (N_599,In_1293,In_1270);
nand U600 (N_600,In_1013,In_341);
nand U601 (N_601,In_2049,In_943);
and U602 (N_602,In_534,In_550);
or U603 (N_603,In_1835,In_1284);
or U604 (N_604,In_2301,In_1182);
and U605 (N_605,In_2122,In_1936);
or U606 (N_606,In_1077,In_62);
nor U607 (N_607,In_1181,In_2303);
nand U608 (N_608,In_544,In_618);
and U609 (N_609,In_1312,In_1569);
xor U610 (N_610,In_1563,In_1231);
nand U611 (N_611,In_1405,In_513);
xor U612 (N_612,In_1078,In_2098);
nand U613 (N_613,In_1874,In_410);
nor U614 (N_614,In_2109,In_2480);
nor U615 (N_615,In_273,In_735);
nand U616 (N_616,In_367,In_395);
xor U617 (N_617,In_2468,In_2418);
xnor U618 (N_618,In_1899,In_1572);
nor U619 (N_619,In_1691,In_1619);
xor U620 (N_620,In_814,In_1716);
nand U621 (N_621,In_2266,In_717);
nand U622 (N_622,In_412,In_1269);
nor U623 (N_623,In_1611,In_884);
nand U624 (N_624,In_346,In_1736);
or U625 (N_625,In_2423,In_357);
nand U626 (N_626,In_2413,In_1961);
nor U627 (N_627,In_2375,In_290);
and U628 (N_628,In_697,In_1907);
xnor U629 (N_629,In_1348,In_949);
nand U630 (N_630,In_1353,In_648);
and U631 (N_631,In_1882,In_1945);
nor U632 (N_632,In_442,In_78);
and U633 (N_633,In_217,In_1873);
or U634 (N_634,In_1160,In_2351);
nor U635 (N_635,In_1916,In_1230);
nor U636 (N_636,In_230,In_674);
and U637 (N_637,In_27,In_1506);
nor U638 (N_638,In_857,In_1578);
and U639 (N_639,In_2282,In_2476);
nand U640 (N_640,In_1012,In_2434);
and U641 (N_641,In_1156,In_1858);
nand U642 (N_642,In_724,In_889);
nand U643 (N_643,In_1268,In_1783);
or U644 (N_644,In_1102,In_2246);
or U645 (N_645,In_1029,In_286);
or U646 (N_646,In_246,In_702);
and U647 (N_647,In_179,In_348);
nand U648 (N_648,In_1245,In_917);
nand U649 (N_649,In_319,In_2053);
xor U650 (N_650,In_176,In_1957);
nor U651 (N_651,In_2358,In_2232);
nor U652 (N_652,In_1468,In_334);
nor U653 (N_653,In_669,In_2039);
xnor U654 (N_654,In_830,In_2008);
or U655 (N_655,In_1570,In_443);
or U656 (N_656,In_1093,In_2124);
xor U657 (N_657,In_622,In_178);
or U658 (N_658,In_1451,In_447);
and U659 (N_659,In_740,In_1443);
nand U660 (N_660,In_870,In_2220);
nor U661 (N_661,In_997,In_312);
nor U662 (N_662,In_2374,In_905);
and U663 (N_663,In_531,In_609);
nor U664 (N_664,In_1175,In_1530);
or U665 (N_665,In_2445,In_1427);
nor U666 (N_666,In_1133,In_2173);
nor U667 (N_667,In_920,In_2127);
xnor U668 (N_668,In_1891,In_854);
xnor U669 (N_669,In_1026,In_1386);
nand U670 (N_670,In_418,In_1766);
or U671 (N_671,In_1933,In_1397);
xnor U672 (N_672,In_355,In_436);
and U673 (N_673,In_2457,In_364);
and U674 (N_674,In_1321,In_1055);
nand U675 (N_675,In_1266,In_1538);
xor U676 (N_676,In_776,In_808);
and U677 (N_677,In_267,In_2401);
or U678 (N_678,In_1921,In_1662);
and U679 (N_679,In_849,In_430);
nor U680 (N_680,In_1962,In_2430);
or U681 (N_681,In_2455,In_999);
nor U682 (N_682,In_1048,In_191);
or U683 (N_683,In_198,In_1462);
and U684 (N_684,In_598,In_456);
or U685 (N_685,In_189,In_73);
xnor U686 (N_686,In_1547,In_373);
nand U687 (N_687,In_1105,In_1287);
and U688 (N_688,In_2114,In_928);
nor U689 (N_689,In_2470,In_2269);
nor U690 (N_690,In_35,In_1499);
xnor U691 (N_691,In_848,In_1436);
nand U692 (N_692,In_1647,In_2424);
nand U693 (N_693,In_767,In_2391);
or U694 (N_694,In_1356,In_2425);
and U695 (N_695,In_359,In_111);
or U696 (N_696,In_287,In_1982);
or U697 (N_697,In_452,In_573);
nand U698 (N_698,In_1929,In_2437);
or U699 (N_699,In_1490,In_501);
nand U700 (N_700,In_477,In_623);
nand U701 (N_701,In_795,In_2247);
nand U702 (N_702,In_2433,In_1922);
and U703 (N_703,In_1031,In_1898);
and U704 (N_704,In_1645,In_948);
nor U705 (N_705,In_84,In_2469);
xor U706 (N_706,In_75,In_964);
nand U707 (N_707,In_1935,In_361);
or U708 (N_708,In_777,In_1545);
or U709 (N_709,In_1655,In_83);
or U710 (N_710,In_1671,In_226);
and U711 (N_711,In_144,In_2313);
and U712 (N_712,In_2471,In_1187);
and U713 (N_713,In_2252,In_827);
and U714 (N_714,In_1494,In_255);
nand U715 (N_715,In_1790,In_783);
xor U716 (N_716,In_2056,In_221);
nand U717 (N_717,In_843,In_1255);
and U718 (N_718,In_1354,In_440);
or U719 (N_719,In_1977,In_183);
or U720 (N_720,In_1833,In_1201);
or U721 (N_721,In_1670,In_2016);
nor U722 (N_722,In_2386,In_86);
nor U723 (N_723,In_2125,In_1542);
nand U724 (N_724,In_2137,In_1302);
or U725 (N_725,In_1183,In_2196);
or U726 (N_726,In_119,In_1086);
nand U727 (N_727,In_1968,In_1488);
or U728 (N_728,In_728,In_114);
or U729 (N_729,In_10,In_1202);
or U730 (N_730,In_2363,In_1316);
nand U731 (N_731,In_784,In_2068);
nand U732 (N_732,In_1560,In_1568);
and U733 (N_733,In_2066,In_1644);
nor U734 (N_734,In_1862,In_1544);
nand U735 (N_735,In_1842,In_1553);
xor U736 (N_736,In_524,In_1170);
or U737 (N_737,In_1748,In_260);
xnor U738 (N_738,In_886,In_2307);
and U739 (N_739,In_30,In_1719);
and U740 (N_740,In_1129,In_1179);
nor U741 (N_741,In_1533,In_1810);
or U742 (N_742,In_1083,In_2204);
xor U743 (N_743,In_1068,In_1512);
and U744 (N_744,In_315,In_1123);
or U745 (N_745,In_1040,In_985);
nand U746 (N_746,In_2154,In_897);
nor U747 (N_747,In_1172,In_458);
and U748 (N_748,In_2010,In_730);
nand U749 (N_749,In_1954,In_1067);
or U750 (N_750,In_1541,In_2240);
and U751 (N_751,In_1726,In_1364);
or U752 (N_752,In_2169,In_1088);
or U753 (N_753,In_2060,In_1686);
nand U754 (N_754,In_1604,In_1787);
nor U755 (N_755,In_2454,In_2151);
and U756 (N_756,In_106,In_989);
nor U757 (N_757,In_899,In_126);
or U758 (N_758,In_542,In_749);
nand U759 (N_759,In_739,In_318);
or U760 (N_760,In_2228,In_1690);
or U761 (N_761,In_2388,In_819);
nor U762 (N_762,In_1368,In_699);
and U763 (N_763,In_158,In_947);
nor U764 (N_764,In_1797,In_661);
nand U765 (N_765,In_939,In_1779);
xnor U766 (N_766,In_1714,In_177);
and U767 (N_767,In_369,In_712);
xor U768 (N_768,In_971,In_1296);
nor U769 (N_769,In_185,In_128);
or U770 (N_770,In_1983,In_654);
nand U771 (N_771,In_2193,In_2000);
nand U772 (N_772,In_1098,In_87);
nand U773 (N_773,In_2029,In_1131);
xor U774 (N_774,In_1927,In_1044);
nor U775 (N_775,In_1917,In_1111);
nand U776 (N_776,In_1470,In_2027);
and U777 (N_777,In_695,In_2412);
nand U778 (N_778,In_90,In_463);
and U779 (N_779,In_1608,In_1775);
nor U780 (N_780,In_1990,In_820);
and U781 (N_781,In_832,In_853);
xnor U782 (N_782,In_80,In_1531);
nand U783 (N_783,In_61,In_835);
and U784 (N_784,In_789,In_1575);
nor U785 (N_785,In_557,In_247);
or U786 (N_786,In_388,In_1859);
nand U787 (N_787,In_1527,In_1292);
or U788 (N_788,In_1124,In_1988);
and U789 (N_789,In_441,In_719);
xor U790 (N_790,In_1752,In_100);
and U791 (N_791,In_21,In_2382);
or U792 (N_792,In_1801,In_723);
or U793 (N_793,In_1717,In_289);
nand U794 (N_794,In_1599,In_47);
or U795 (N_795,In_1725,In_1212);
nor U796 (N_796,In_972,In_563);
nor U797 (N_797,In_202,In_161);
nand U798 (N_798,In_1653,In_2348);
nand U799 (N_799,In_33,In_2343);
or U800 (N_800,In_1496,In_967);
nor U801 (N_801,In_471,In_2410);
or U802 (N_802,In_1320,In_1331);
or U803 (N_803,In_54,In_1051);
and U804 (N_804,In_426,In_628);
or U805 (N_805,In_1657,In_1602);
nor U806 (N_806,In_2264,In_2249);
nor U807 (N_807,In_28,In_1967);
nor U808 (N_808,In_2012,In_489);
and U809 (N_809,In_1722,In_1516);
nor U810 (N_810,In_1818,In_231);
xor U811 (N_811,In_2115,In_998);
xnor U812 (N_812,In_445,In_93);
nand U813 (N_813,In_1281,In_751);
and U814 (N_814,In_109,In_2189);
nand U815 (N_815,In_107,In_1314);
and U816 (N_816,In_2385,In_840);
nand U817 (N_817,In_658,In_944);
xor U818 (N_818,In_1751,In_956);
and U819 (N_819,In_1036,In_1408);
or U820 (N_820,In_1158,In_1495);
nand U821 (N_821,In_507,In_1761);
or U822 (N_822,In_1852,In_1149);
nor U823 (N_823,In_2414,In_1646);
and U824 (N_824,In_586,In_1667);
nand U825 (N_825,In_1330,In_1999);
and U826 (N_826,In_1251,In_1561);
xnor U827 (N_827,In_306,In_229);
nand U828 (N_828,In_509,In_1384);
and U829 (N_829,In_1953,In_363);
or U830 (N_830,In_1804,In_526);
nand U831 (N_831,In_399,In_781);
or U832 (N_832,In_1884,In_1629);
xor U833 (N_833,In_881,In_757);
nor U834 (N_834,In_132,In_1502);
xor U835 (N_835,In_590,In_1404);
and U836 (N_836,In_1274,In_833);
or U837 (N_837,In_327,In_2037);
nand U838 (N_838,In_1642,In_335);
nor U839 (N_839,In_2298,In_1596);
nor U840 (N_840,In_640,In_1409);
and U841 (N_841,In_571,In_339);
nor U842 (N_842,In_1057,In_505);
nor U843 (N_843,In_1526,In_1939);
and U844 (N_844,In_2417,In_1072);
xor U845 (N_845,In_1373,In_1455);
nand U846 (N_846,In_1001,In_1041);
nand U847 (N_847,In_1537,In_2359);
or U848 (N_848,In_2333,In_1546);
or U849 (N_849,In_429,In_59);
or U850 (N_850,In_491,In_259);
and U851 (N_851,In_1300,In_266);
nor U852 (N_852,In_311,In_841);
nor U853 (N_853,In_806,In_2163);
nand U854 (N_854,In_1285,In_397);
and U855 (N_855,In_1912,In_480);
and U856 (N_856,In_961,In_2273);
and U857 (N_857,In_481,In_1014);
or U858 (N_858,In_1668,In_2047);
nor U859 (N_859,In_2168,In_79);
and U860 (N_860,In_1492,In_165);
xor U861 (N_861,In_1011,In_32);
xnor U862 (N_862,In_1148,In_1020);
or U863 (N_863,In_579,In_2043);
and U864 (N_864,In_352,In_14);
or U865 (N_865,In_894,In_2061);
nand U866 (N_866,In_576,In_2172);
or U867 (N_867,In_67,In_792);
nor U868 (N_868,In_1523,In_2215);
xor U869 (N_869,In_589,In_2040);
xnor U870 (N_870,In_150,In_478);
and U871 (N_871,In_2404,In_938);
and U872 (N_872,In_2381,In_1780);
nand U873 (N_873,In_2033,In_2397);
or U874 (N_874,In_1210,In_645);
nor U875 (N_875,In_930,In_588);
nor U876 (N_876,In_2136,In_1448);
and U877 (N_877,In_251,In_484);
nand U878 (N_878,In_663,In_2146);
and U879 (N_879,In_1824,In_1220);
nor U880 (N_880,In_1958,In_1600);
or U881 (N_881,In_763,In_931);
or U882 (N_882,In_2336,In_1960);
nand U883 (N_883,In_737,In_876);
nor U884 (N_884,In_734,In_1910);
xor U885 (N_885,In_160,In_1740);
or U886 (N_886,In_301,In_1421);
nand U887 (N_887,In_700,In_2229);
nand U888 (N_888,In_205,In_1278);
or U889 (N_889,In_2081,In_1924);
nand U890 (N_890,In_1505,In_968);
nand U891 (N_891,In_1965,In_1185);
nand U892 (N_892,In_97,In_1474);
nand U893 (N_893,In_353,In_1447);
and U894 (N_894,In_1191,In_962);
and U895 (N_895,In_1820,In_1165);
nand U896 (N_896,In_1297,In_1301);
xor U897 (N_897,In_298,In_1407);
nand U898 (N_898,In_490,In_2112);
xor U899 (N_899,In_630,In_362);
and U900 (N_900,In_2050,In_1118);
or U901 (N_901,In_922,In_29);
and U902 (N_902,In_2057,In_1392);
xnor U903 (N_903,In_216,In_927);
nor U904 (N_904,In_2186,In_1893);
nand U905 (N_905,In_1009,In_1792);
nor U906 (N_906,In_762,In_2319);
nor U907 (N_907,In_326,In_2248);
or U908 (N_908,In_1419,In_2444);
nand U909 (N_909,In_1155,In_2174);
or U910 (N_910,In_2077,In_2316);
or U911 (N_911,In_2344,In_578);
nand U912 (N_912,In_1167,In_1106);
nand U913 (N_913,In_338,In_901);
nor U914 (N_914,In_1358,In_1549);
nand U915 (N_915,In_310,In_847);
nand U916 (N_916,In_187,In_919);
and U917 (N_917,In_149,In_1913);
nor U918 (N_918,In_227,In_1034);
and U919 (N_919,In_957,In_64);
and U920 (N_920,In_342,In_567);
or U921 (N_921,In_136,In_451);
nor U922 (N_922,In_584,In_1762);
and U923 (N_923,In_718,In_1283);
nand U924 (N_924,In_2314,In_1060);
or U925 (N_925,In_38,In_1908);
or U926 (N_926,In_577,In_1457);
nand U927 (N_927,In_666,In_1871);
nand U928 (N_928,In_1177,In_647);
or U929 (N_929,In_2345,In_554);
nand U930 (N_930,In_1498,In_344);
or U931 (N_931,In_2451,In_284);
or U932 (N_932,In_1603,In_1215);
and U933 (N_933,In_2473,In_1701);
nand U934 (N_934,In_608,In_1325);
and U935 (N_935,In_1206,In_1688);
nand U936 (N_936,In_1987,In_1806);
or U937 (N_937,In_1840,In_2394);
nor U938 (N_938,In_995,In_1444);
nand U939 (N_939,In_733,In_2294);
nor U940 (N_940,In_2150,In_487);
nor U941 (N_941,In_2450,In_2054);
and U942 (N_942,In_785,In_954);
xor U943 (N_943,In_45,In_2201);
nand U944 (N_944,In_1682,In_63);
nor U945 (N_945,In_1489,In_285);
nor U946 (N_946,In_182,In_1738);
and U947 (N_947,In_1259,In_1005);
nor U948 (N_948,In_159,In_520);
or U949 (N_949,In_1477,In_1322);
or U950 (N_950,In_1066,In_2239);
or U951 (N_951,In_2238,In_1313);
or U952 (N_952,In_1938,In_1821);
nand U953 (N_953,In_398,In_416);
nand U954 (N_954,In_1914,In_2341);
xor U955 (N_955,In_2003,In_2267);
xor U956 (N_956,In_1195,In_1698);
nand U957 (N_957,In_863,In_560);
or U958 (N_958,In_1023,In_1058);
nand U959 (N_959,In_2376,In_1796);
nor U960 (N_960,In_910,In_907);
nand U961 (N_961,In_2188,In_1091);
nand U962 (N_962,In_2389,In_123);
or U963 (N_963,In_839,In_1037);
nand U964 (N_964,In_2285,In_1439);
nor U965 (N_965,In_331,In_1554);
nor U966 (N_966,In_1205,In_537);
nor U967 (N_967,In_1464,In_525);
nand U968 (N_968,In_810,In_2132);
or U969 (N_969,In_2453,In_1027);
nand U970 (N_970,In_984,In_865);
or U971 (N_971,In_1141,In_1275);
nand U972 (N_972,In_2171,In_2485);
and U973 (N_973,In_1731,In_51);
or U974 (N_974,In_1169,In_1352);
xnor U975 (N_975,In_1865,In_2013);
nor U976 (N_976,In_1045,In_1900);
and U977 (N_977,In_1802,In_1548);
and U978 (N_978,In_1850,In_1260);
nand U979 (N_979,In_888,In_2157);
nand U980 (N_980,In_1246,In_493);
nand U981 (N_981,In_195,In_1975);
or U982 (N_982,In_1130,In_1100);
and U983 (N_983,In_208,In_1237);
nor U984 (N_984,In_1674,In_457);
and U985 (N_985,In_2026,In_1695);
and U986 (N_986,In_1486,In_2320);
or U987 (N_987,In_1974,In_636);
xor U988 (N_988,In_248,In_1084);
nor U989 (N_989,In_2103,In_2416);
nand U990 (N_990,In_1039,In_1103);
or U991 (N_991,In_1757,In_321);
or U992 (N_992,In_2110,In_1989);
nor U993 (N_993,In_1396,In_1640);
and U994 (N_994,In_2277,In_1035);
nor U995 (N_995,In_1065,In_134);
nor U996 (N_996,In_133,In_1680);
or U997 (N_997,In_425,In_1038);
and U998 (N_998,In_715,In_1507);
nand U999 (N_999,In_1487,In_1728);
and U1000 (N_1000,In_308,In_2034);
nand U1001 (N_1001,In_1622,In_1699);
nand U1002 (N_1002,In_594,In_469);
and U1003 (N_1003,In_1152,In_1692);
nand U1004 (N_1004,In_1318,In_2352);
or U1005 (N_1005,In_325,In_771);
nand U1006 (N_1006,In_2177,In_2158);
nand U1007 (N_1007,In_880,In_2304);
xnor U1008 (N_1008,In_752,In_2212);
or U1009 (N_1009,In_2144,In_9);
nand U1010 (N_1010,In_218,In_1816);
nor U1011 (N_1011,In_1598,In_2116);
and U1012 (N_1012,In_2462,In_690);
and U1013 (N_1013,In_2059,In_2287);
and U1014 (N_1014,In_2403,In_768);
nor U1015 (N_1015,In_1951,In_402);
nor U1016 (N_1016,In_955,In_2102);
xnor U1017 (N_1017,In_667,In_515);
nor U1018 (N_1018,In_12,In_2289);
and U1019 (N_1019,In_275,In_1590);
xor U1020 (N_1020,In_1422,In_1567);
or U1021 (N_1021,In_1940,In_2350);
or U1022 (N_1022,In_466,In_1615);
nor U1023 (N_1023,In_575,In_2216);
nand U1024 (N_1024,In_1730,In_5);
and U1025 (N_1025,In_1509,In_1370);
xnor U1026 (N_1026,In_552,In_722);
and U1027 (N_1027,In_2446,In_1681);
nand U1028 (N_1028,In_906,In_1371);
nand U1029 (N_1029,In_1905,In_685);
or U1030 (N_1030,In_1484,In_345);
nand U1031 (N_1031,In_115,In_2152);
nor U1032 (N_1032,In_1228,In_297);
nand U1033 (N_1033,In_1147,In_494);
xor U1034 (N_1034,In_878,In_1678);
xnor U1035 (N_1035,In_991,In_2048);
and U1036 (N_1036,In_1966,In_386);
and U1037 (N_1037,In_903,In_1344);
nor U1038 (N_1038,In_1276,In_1372);
nand U1039 (N_1039,In_377,In_437);
or U1040 (N_1040,In_1785,In_2384);
nor U1041 (N_1041,In_1707,In_612);
and U1042 (N_1042,In_1813,In_982);
nand U1043 (N_1043,In_1649,In_2006);
or U1044 (N_1044,In_1807,In_4);
or U1045 (N_1045,In_707,In_736);
and U1046 (N_1046,In_2190,In_574);
xor U1047 (N_1047,In_2224,In_1207);
nand U1048 (N_1048,In_2270,In_2096);
or U1049 (N_1049,In_2213,In_1121);
and U1050 (N_1050,In_774,In_665);
xnor U1051 (N_1051,In_455,In_291);
and U1052 (N_1052,In_2031,In_2141);
or U1053 (N_1053,In_932,In_619);
nand U1054 (N_1054,In_15,In_1096);
or U1055 (N_1055,In_1869,In_844);
nand U1056 (N_1056,In_656,In_1623);
and U1057 (N_1057,In_1742,In_1305);
nor U1058 (N_1058,In_2117,In_2427);
nor U1059 (N_1059,In_2176,In_1004);
nand U1060 (N_1060,In_646,In_1047);
xnor U1061 (N_1061,In_1652,In_817);
or U1062 (N_1062,In_887,In_2079);
xnor U1063 (N_1063,In_1140,In_135);
or U1064 (N_1064,In_738,In_2099);
nand U1065 (N_1065,In_1145,In_482);
nor U1066 (N_1066,In_1114,In_681);
xor U1067 (N_1067,In_420,In_2306);
and U1068 (N_1068,In_765,In_1340);
nor U1069 (N_1069,In_1648,In_2138);
and U1070 (N_1070,In_682,In_911);
or U1071 (N_1071,In_1225,In_1903);
nand U1072 (N_1072,In_1580,In_1329);
or U1073 (N_1073,In_963,In_1081);
xnor U1074 (N_1074,In_748,In_2120);
nor U1075 (N_1075,In_1919,In_1075);
xor U1076 (N_1076,In_539,In_459);
or U1077 (N_1077,In_649,In_1442);
or U1078 (N_1078,In_1395,In_2009);
nor U1079 (N_1079,In_2170,In_1420);
nand U1080 (N_1080,In_1750,In_2337);
and U1081 (N_1081,In_1426,In_192);
and U1082 (N_1082,In_2408,In_1853);
nor U1083 (N_1083,In_2074,In_694);
xor U1084 (N_1084,In_1424,In_1679);
nand U1085 (N_1085,In_299,In_790);
xnor U1086 (N_1086,In_1758,In_1189);
and U1087 (N_1087,In_1583,In_351);
or U1088 (N_1088,In_794,In_1562);
nand U1089 (N_1089,In_1217,In_2052);
and U1090 (N_1090,In_19,In_1949);
or U1091 (N_1091,In_1854,In_1920);
and U1092 (N_1092,In_1043,In_200);
and U1093 (N_1093,In_2364,In_1211);
nand U1094 (N_1094,In_508,In_1074);
or U1095 (N_1095,In_156,In_1163);
xnor U1096 (N_1096,In_6,In_407);
nor U1097 (N_1097,In_582,In_52);
nor U1098 (N_1098,In_1403,In_1659);
and U1099 (N_1099,In_891,In_2046);
or U1100 (N_1100,In_2175,In_343);
nand U1101 (N_1101,In_898,In_2242);
or U1102 (N_1102,In_108,In_2378);
or U1103 (N_1103,In_1144,In_896);
nor U1104 (N_1104,In_543,In_302);
nor U1105 (N_1105,In_2091,In_1637);
or U1106 (N_1106,In_1981,In_1342);
or U1107 (N_1107,In_1440,In_141);
nand U1108 (N_1108,In_495,In_1825);
nor U1109 (N_1109,In_1973,In_1607);
nand U1110 (N_1110,In_1972,In_868);
nor U1111 (N_1111,In_850,In_2243);
nand U1112 (N_1112,In_1525,In_1097);
nand U1113 (N_1113,In_1378,In_2395);
xnor U1114 (N_1114,In_779,In_951);
and U1115 (N_1115,In_2140,In_274);
nand U1116 (N_1116,In_1317,In_2279);
or U1117 (N_1117,In_1415,In_856);
and U1118 (N_1118,In_2419,In_8);
nor U1119 (N_1119,In_1166,In_1493);
nand U1120 (N_1120,In_1366,In_1122);
nor U1121 (N_1121,In_1683,In_770);
and U1122 (N_1122,In_1948,In_1633);
nor U1123 (N_1123,In_76,In_1355);
and U1124 (N_1124,In_595,In_95);
or U1125 (N_1125,In_1911,In_750);
nand U1126 (N_1126,In_292,In_1159);
or U1127 (N_1127,In_1112,In_1303);
nand U1128 (N_1128,In_558,In_102);
and U1129 (N_1129,In_2494,In_1241);
nand U1130 (N_1130,In_1002,In_2276);
xnor U1131 (N_1131,In_644,In_2330);
nand U1132 (N_1132,In_476,In_210);
and U1133 (N_1133,In_851,In_772);
nor U1134 (N_1134,In_1543,In_1729);
nor U1135 (N_1135,In_974,In_1357);
nand U1136 (N_1136,In_671,In_2338);
nand U1137 (N_1137,In_419,In_1115);
nor U1138 (N_1138,In_1904,In_2030);
nor U1139 (N_1139,In_980,In_366);
and U1140 (N_1140,In_422,In_1021);
or U1141 (N_1141,In_2495,In_2458);
nor U1142 (N_1142,In_659,In_148);
nand U1143 (N_1143,In_234,In_1866);
or U1144 (N_1144,In_392,In_1028);
or U1145 (N_1145,In_196,In_1497);
xor U1146 (N_1146,In_1892,In_1391);
nor U1147 (N_1147,In_696,In_460);
nor U1148 (N_1148,In_382,In_270);
nand U1149 (N_1149,In_498,In_1388);
or U1150 (N_1150,In_2018,In_2078);
or U1151 (N_1151,In_2036,In_194);
nor U1152 (N_1152,In_1819,In_2065);
nand U1153 (N_1153,In_1379,In_1061);
or U1154 (N_1154,In_2475,In_953);
xor U1155 (N_1155,In_1032,In_1890);
xnor U1156 (N_1156,In_713,In_1883);
and U1157 (N_1157,In_1794,In_2022);
or U1158 (N_1158,In_684,In_530);
nor U1159 (N_1159,In_2139,In_642);
and U1160 (N_1160,In_1838,In_1915);
and U1161 (N_1161,In_1229,In_1784);
nor U1162 (N_1162,In_517,In_163);
xnor U1163 (N_1163,In_1460,In_488);
nor U1164 (N_1164,In_1359,In_616);
or U1165 (N_1165,In_1271,In_1307);
or U1166 (N_1166,In_124,In_693);
nand U1167 (N_1167,In_788,In_2317);
and U1168 (N_1168,In_2021,In_2258);
and U1169 (N_1169,In_673,In_1582);
and U1170 (N_1170,In_2323,In_1375);
nor U1171 (N_1171,In_2274,In_1770);
and U1172 (N_1172,In_1774,In_242);
or U1173 (N_1173,In_2275,In_1798);
or U1174 (N_1174,In_2288,In_2062);
nor U1175 (N_1175,In_2075,In_1333);
and U1176 (N_1176,In_332,In_1934);
nand U1177 (N_1177,In_1863,In_2373);
nor U1178 (N_1178,In_409,In_935);
nor U1179 (N_1179,In_454,In_81);
nand U1180 (N_1180,In_1631,In_549);
and U1181 (N_1181,In_1094,In_1747);
and U1182 (N_1182,In_57,In_1006);
or U1183 (N_1183,In_852,In_1254);
xor U1184 (N_1184,In_1423,In_2095);
or U1185 (N_1185,In_2488,In_1107);
nand U1186 (N_1186,In_2293,In_1095);
nor U1187 (N_1187,In_1090,In_396);
or U1188 (N_1188,In_151,In_1054);
and U1189 (N_1189,In_606,In_1401);
nor U1190 (N_1190,In_1814,In_2265);
nand U1191 (N_1191,In_1941,In_994);
nand U1192 (N_1192,In_1139,In_1556);
xnor U1193 (N_1193,In_2421,In_2237);
xor U1194 (N_1194,In_2245,In_973);
or U1195 (N_1195,In_2367,In_1033);
or U1196 (N_1196,In_434,In_389);
nor U1197 (N_1197,In_276,In_532);
nor U1198 (N_1198,In_556,In_1720);
and U1199 (N_1199,In_2268,In_912);
xnor U1200 (N_1200,In_1721,In_219);
nor U1201 (N_1201,In_1524,In_1868);
nand U1202 (N_1202,In_1085,In_2241);
nor U1203 (N_1203,In_60,In_2182);
nor U1204 (N_1204,In_2461,In_2007);
nor U1205 (N_1205,In_2486,In_1249);
and U1206 (N_1206,In_1723,In_1522);
and U1207 (N_1207,In_450,In_1639);
nand U1208 (N_1208,In_2020,In_1286);
nor U1209 (N_1209,In_2225,In_1696);
nor U1210 (N_1210,In_1665,In_1008);
nand U1211 (N_1211,In_1092,In_1937);
or U1212 (N_1212,In_1713,In_950);
nor U1213 (N_1213,In_607,In_1226);
nor U1214 (N_1214,In_855,In_1885);
xnor U1215 (N_1215,In_675,In_140);
or U1216 (N_1216,In_138,In_1458);
or U1217 (N_1217,In_2024,In_68);
nand U1218 (N_1218,In_1154,In_2088);
or U1219 (N_1219,In_921,In_895);
or U1220 (N_1220,In_39,In_1677);
xnor U1221 (N_1221,In_2438,In_1540);
nand U1222 (N_1222,In_1997,In_214);
or U1223 (N_1223,In_347,In_485);
and U1224 (N_1224,In_2459,In_2011);
nor U1225 (N_1225,In_1015,In_295);
and U1226 (N_1226,In_238,In_2383);
nor U1227 (N_1227,In_1376,In_2180);
nor U1228 (N_1228,In_1324,In_2347);
nand U1229 (N_1229,In_2202,In_1666);
and U1230 (N_1230,In_535,In_1932);
and U1231 (N_1231,In_1776,In_2069);
nor U1232 (N_1232,In_2118,In_599);
and U1233 (N_1233,In_653,In_2365);
nor U1234 (N_1234,In_2087,In_660);
nor U1235 (N_1235,In_759,In_1343);
nand U1236 (N_1236,In_1473,In_726);
nand U1237 (N_1237,In_871,In_2392);
xnor U1238 (N_1238,In_958,In_551);
nand U1239 (N_1239,In_1367,In_940);
and U1240 (N_1240,In_24,In_74);
nor U1241 (N_1241,In_2460,In_168);
xnor U1242 (N_1242,In_1016,In_423);
nand U1243 (N_1243,In_1003,In_428);
or U1244 (N_1244,In_553,In_2244);
and U1245 (N_1245,In_1267,In_2299);
nor U1246 (N_1246,In_1676,In_393);
or U1247 (N_1247,In_1971,In_860);
or U1248 (N_1248,In_199,In_1108);
nor U1249 (N_1249,In_1845,In_1168);
nor U1250 (N_1250,In_1326,In_1444);
nand U1251 (N_1251,In_790,In_1157);
and U1252 (N_1252,In_1065,In_2293);
and U1253 (N_1253,In_882,In_1141);
nand U1254 (N_1254,In_2338,In_1758);
nand U1255 (N_1255,In_127,In_910);
nand U1256 (N_1256,In_1385,In_230);
xnor U1257 (N_1257,In_2435,In_1222);
or U1258 (N_1258,In_2337,In_214);
or U1259 (N_1259,In_591,In_1949);
nand U1260 (N_1260,In_2157,In_2496);
and U1261 (N_1261,In_230,In_1340);
and U1262 (N_1262,In_895,In_501);
nor U1263 (N_1263,In_2487,In_1048);
or U1264 (N_1264,In_57,In_1905);
or U1265 (N_1265,In_2354,In_1179);
xor U1266 (N_1266,In_2292,In_1710);
and U1267 (N_1267,In_1482,In_361);
xor U1268 (N_1268,In_382,In_1613);
nor U1269 (N_1269,In_819,In_126);
or U1270 (N_1270,In_723,In_1071);
and U1271 (N_1271,In_2474,In_34);
and U1272 (N_1272,In_718,In_3);
and U1273 (N_1273,In_1706,In_970);
xnor U1274 (N_1274,In_1016,In_512);
and U1275 (N_1275,In_439,In_711);
and U1276 (N_1276,In_792,In_664);
nand U1277 (N_1277,In_437,In_973);
or U1278 (N_1278,In_132,In_745);
xnor U1279 (N_1279,In_1607,In_2240);
nand U1280 (N_1280,In_2317,In_1902);
xnor U1281 (N_1281,In_233,In_2028);
or U1282 (N_1282,In_1996,In_473);
or U1283 (N_1283,In_819,In_25);
and U1284 (N_1284,In_1324,In_1197);
nor U1285 (N_1285,In_148,In_379);
or U1286 (N_1286,In_2394,In_2120);
xor U1287 (N_1287,In_2,In_342);
and U1288 (N_1288,In_1187,In_1243);
and U1289 (N_1289,In_2274,In_1037);
or U1290 (N_1290,In_626,In_236);
xor U1291 (N_1291,In_1387,In_1920);
or U1292 (N_1292,In_66,In_304);
xor U1293 (N_1293,In_553,In_1599);
or U1294 (N_1294,In_1535,In_1136);
nor U1295 (N_1295,In_2339,In_1460);
and U1296 (N_1296,In_2134,In_801);
nor U1297 (N_1297,In_578,In_435);
nand U1298 (N_1298,In_2045,In_810);
or U1299 (N_1299,In_431,In_1607);
nor U1300 (N_1300,In_2293,In_2105);
or U1301 (N_1301,In_667,In_63);
or U1302 (N_1302,In_1747,In_1982);
nand U1303 (N_1303,In_1798,In_741);
nor U1304 (N_1304,In_1106,In_1565);
or U1305 (N_1305,In_1061,In_2259);
xnor U1306 (N_1306,In_1863,In_2404);
nand U1307 (N_1307,In_157,In_617);
or U1308 (N_1308,In_559,In_421);
or U1309 (N_1309,In_2414,In_1524);
or U1310 (N_1310,In_779,In_1426);
and U1311 (N_1311,In_1704,In_373);
xnor U1312 (N_1312,In_1526,In_985);
nand U1313 (N_1313,In_749,In_1797);
nand U1314 (N_1314,In_408,In_2118);
nor U1315 (N_1315,In_2044,In_1337);
nor U1316 (N_1316,In_1766,In_513);
and U1317 (N_1317,In_2191,In_822);
and U1318 (N_1318,In_1666,In_453);
nand U1319 (N_1319,In_1696,In_1526);
nor U1320 (N_1320,In_493,In_2377);
and U1321 (N_1321,In_1033,In_2392);
xor U1322 (N_1322,In_1599,In_108);
nand U1323 (N_1323,In_1187,In_1710);
nor U1324 (N_1324,In_1212,In_863);
nand U1325 (N_1325,In_574,In_1479);
nand U1326 (N_1326,In_1007,In_1062);
xor U1327 (N_1327,In_2344,In_1367);
or U1328 (N_1328,In_38,In_1123);
or U1329 (N_1329,In_1172,In_2419);
nor U1330 (N_1330,In_2434,In_2452);
xnor U1331 (N_1331,In_1219,In_1894);
or U1332 (N_1332,In_85,In_1652);
or U1333 (N_1333,In_917,In_893);
or U1334 (N_1334,In_1397,In_1280);
nand U1335 (N_1335,In_1815,In_1635);
nand U1336 (N_1336,In_614,In_2018);
nor U1337 (N_1337,In_230,In_1419);
xor U1338 (N_1338,In_1982,In_1799);
nor U1339 (N_1339,In_1693,In_1920);
nand U1340 (N_1340,In_308,In_108);
nand U1341 (N_1341,In_1209,In_423);
and U1342 (N_1342,In_2454,In_1832);
nand U1343 (N_1343,In_1199,In_118);
nand U1344 (N_1344,In_1236,In_242);
or U1345 (N_1345,In_1730,In_399);
or U1346 (N_1346,In_190,In_1128);
nand U1347 (N_1347,In_1001,In_447);
and U1348 (N_1348,In_252,In_955);
nor U1349 (N_1349,In_2302,In_1309);
and U1350 (N_1350,In_1683,In_112);
nor U1351 (N_1351,In_1199,In_1806);
or U1352 (N_1352,In_952,In_216);
and U1353 (N_1353,In_1710,In_1290);
nor U1354 (N_1354,In_2341,In_863);
or U1355 (N_1355,In_2161,In_1850);
or U1356 (N_1356,In_624,In_2031);
xor U1357 (N_1357,In_1169,In_335);
nand U1358 (N_1358,In_1121,In_723);
nor U1359 (N_1359,In_768,In_708);
nor U1360 (N_1360,In_2311,In_423);
xor U1361 (N_1361,In_569,In_314);
nand U1362 (N_1362,In_1692,In_1920);
or U1363 (N_1363,In_2293,In_422);
and U1364 (N_1364,In_1075,In_499);
nand U1365 (N_1365,In_474,In_1748);
nor U1366 (N_1366,In_2312,In_1527);
and U1367 (N_1367,In_173,In_1878);
and U1368 (N_1368,In_1529,In_1185);
or U1369 (N_1369,In_1691,In_537);
nand U1370 (N_1370,In_1667,In_194);
nand U1371 (N_1371,In_1285,In_1363);
or U1372 (N_1372,In_1924,In_832);
xnor U1373 (N_1373,In_2414,In_90);
xor U1374 (N_1374,In_902,In_1270);
nor U1375 (N_1375,In_794,In_799);
and U1376 (N_1376,In_1837,In_504);
nor U1377 (N_1377,In_1231,In_104);
nor U1378 (N_1378,In_1487,In_20);
nor U1379 (N_1379,In_4,In_354);
and U1380 (N_1380,In_675,In_1033);
nand U1381 (N_1381,In_1778,In_299);
or U1382 (N_1382,In_2434,In_22);
and U1383 (N_1383,In_291,In_597);
nand U1384 (N_1384,In_2492,In_322);
and U1385 (N_1385,In_727,In_446);
and U1386 (N_1386,In_512,In_2115);
and U1387 (N_1387,In_843,In_693);
or U1388 (N_1388,In_1769,In_132);
nand U1389 (N_1389,In_1884,In_1551);
nand U1390 (N_1390,In_592,In_2140);
nand U1391 (N_1391,In_214,In_703);
or U1392 (N_1392,In_764,In_2124);
nor U1393 (N_1393,In_2418,In_1543);
nand U1394 (N_1394,In_204,In_915);
nand U1395 (N_1395,In_2360,In_451);
or U1396 (N_1396,In_94,In_47);
nor U1397 (N_1397,In_1725,In_2262);
nor U1398 (N_1398,In_1487,In_740);
or U1399 (N_1399,In_506,In_1310);
or U1400 (N_1400,In_329,In_355);
and U1401 (N_1401,In_1986,In_2433);
nand U1402 (N_1402,In_1168,In_1609);
or U1403 (N_1403,In_178,In_2300);
xor U1404 (N_1404,In_1255,In_2230);
nor U1405 (N_1405,In_1637,In_522);
nor U1406 (N_1406,In_60,In_384);
xor U1407 (N_1407,In_1464,In_1343);
nor U1408 (N_1408,In_715,In_531);
nor U1409 (N_1409,In_636,In_2127);
nand U1410 (N_1410,In_1300,In_383);
or U1411 (N_1411,In_1312,In_738);
or U1412 (N_1412,In_2074,In_2329);
nor U1413 (N_1413,In_2337,In_920);
xnor U1414 (N_1414,In_2146,In_1904);
nor U1415 (N_1415,In_509,In_908);
nand U1416 (N_1416,In_2473,In_1355);
nand U1417 (N_1417,In_2029,In_638);
or U1418 (N_1418,In_517,In_2466);
nand U1419 (N_1419,In_578,In_1570);
nand U1420 (N_1420,In_790,In_1246);
nand U1421 (N_1421,In_212,In_2419);
or U1422 (N_1422,In_1615,In_1253);
or U1423 (N_1423,In_732,In_165);
and U1424 (N_1424,In_2189,In_1472);
or U1425 (N_1425,In_1145,In_1574);
and U1426 (N_1426,In_2433,In_2219);
nand U1427 (N_1427,In_2178,In_870);
nand U1428 (N_1428,In_1869,In_529);
or U1429 (N_1429,In_2039,In_594);
and U1430 (N_1430,In_104,In_734);
nand U1431 (N_1431,In_2382,In_1630);
xnor U1432 (N_1432,In_2328,In_1647);
and U1433 (N_1433,In_151,In_2417);
and U1434 (N_1434,In_1764,In_2161);
nor U1435 (N_1435,In_1243,In_596);
and U1436 (N_1436,In_2210,In_519);
xor U1437 (N_1437,In_436,In_505);
or U1438 (N_1438,In_1518,In_481);
nor U1439 (N_1439,In_2362,In_2031);
and U1440 (N_1440,In_884,In_2231);
or U1441 (N_1441,In_266,In_1466);
nand U1442 (N_1442,In_1550,In_1009);
xor U1443 (N_1443,In_486,In_300);
and U1444 (N_1444,In_1710,In_2430);
xor U1445 (N_1445,In_212,In_1699);
xnor U1446 (N_1446,In_442,In_177);
nor U1447 (N_1447,In_2275,In_7);
xor U1448 (N_1448,In_2263,In_908);
nor U1449 (N_1449,In_1333,In_1441);
nor U1450 (N_1450,In_1647,In_1035);
nand U1451 (N_1451,In_1454,In_2004);
nor U1452 (N_1452,In_1320,In_2356);
and U1453 (N_1453,In_2493,In_528);
or U1454 (N_1454,In_803,In_2319);
nand U1455 (N_1455,In_1806,In_908);
and U1456 (N_1456,In_1795,In_808);
or U1457 (N_1457,In_72,In_1019);
or U1458 (N_1458,In_92,In_1024);
or U1459 (N_1459,In_1764,In_1339);
nor U1460 (N_1460,In_893,In_2105);
xnor U1461 (N_1461,In_2373,In_443);
and U1462 (N_1462,In_589,In_1006);
and U1463 (N_1463,In_423,In_1688);
nand U1464 (N_1464,In_463,In_1005);
and U1465 (N_1465,In_1752,In_725);
nor U1466 (N_1466,In_621,In_1273);
nor U1467 (N_1467,In_96,In_1349);
nor U1468 (N_1468,In_1547,In_337);
and U1469 (N_1469,In_2117,In_315);
nand U1470 (N_1470,In_1328,In_1551);
or U1471 (N_1471,In_227,In_438);
or U1472 (N_1472,In_2459,In_1109);
and U1473 (N_1473,In_1317,In_1997);
nor U1474 (N_1474,In_2470,In_603);
nor U1475 (N_1475,In_516,In_2392);
and U1476 (N_1476,In_1748,In_917);
nor U1477 (N_1477,In_1227,In_1044);
nor U1478 (N_1478,In_957,In_515);
or U1479 (N_1479,In_1782,In_2038);
and U1480 (N_1480,In_1296,In_1677);
nand U1481 (N_1481,In_2301,In_2223);
or U1482 (N_1482,In_2380,In_383);
xnor U1483 (N_1483,In_2078,In_78);
and U1484 (N_1484,In_457,In_849);
and U1485 (N_1485,In_1543,In_2013);
or U1486 (N_1486,In_1840,In_1959);
xnor U1487 (N_1487,In_1213,In_54);
and U1488 (N_1488,In_1127,In_953);
xnor U1489 (N_1489,In_2240,In_2198);
and U1490 (N_1490,In_1603,In_1668);
nor U1491 (N_1491,In_2094,In_2269);
xor U1492 (N_1492,In_559,In_663);
or U1493 (N_1493,In_1048,In_1451);
and U1494 (N_1494,In_2372,In_2376);
and U1495 (N_1495,In_2034,In_282);
or U1496 (N_1496,In_560,In_188);
nand U1497 (N_1497,In_891,In_614);
or U1498 (N_1498,In_2313,In_1810);
and U1499 (N_1499,In_1756,In_653);
or U1500 (N_1500,In_1299,In_1136);
and U1501 (N_1501,In_103,In_2467);
nor U1502 (N_1502,In_1313,In_2406);
nor U1503 (N_1503,In_108,In_2402);
nand U1504 (N_1504,In_735,In_2436);
and U1505 (N_1505,In_396,In_553);
or U1506 (N_1506,In_1850,In_2030);
and U1507 (N_1507,In_366,In_314);
nor U1508 (N_1508,In_1129,In_1052);
nor U1509 (N_1509,In_1178,In_1228);
nand U1510 (N_1510,In_451,In_1734);
or U1511 (N_1511,In_1723,In_2290);
and U1512 (N_1512,In_1400,In_1734);
nor U1513 (N_1513,In_483,In_42);
nand U1514 (N_1514,In_2171,In_44);
nand U1515 (N_1515,In_152,In_425);
nor U1516 (N_1516,In_1098,In_620);
nor U1517 (N_1517,In_2191,In_1029);
or U1518 (N_1518,In_85,In_2015);
and U1519 (N_1519,In_448,In_852);
or U1520 (N_1520,In_1554,In_865);
xnor U1521 (N_1521,In_1307,In_2075);
nor U1522 (N_1522,In_1706,In_2188);
xor U1523 (N_1523,In_2460,In_372);
nor U1524 (N_1524,In_2206,In_2273);
nor U1525 (N_1525,In_15,In_1380);
and U1526 (N_1526,In_1512,In_486);
or U1527 (N_1527,In_1507,In_1311);
nand U1528 (N_1528,In_301,In_2076);
or U1529 (N_1529,In_856,In_1276);
xor U1530 (N_1530,In_255,In_212);
nand U1531 (N_1531,In_1472,In_708);
and U1532 (N_1532,In_1453,In_664);
nand U1533 (N_1533,In_1489,In_715);
or U1534 (N_1534,In_1432,In_1506);
or U1535 (N_1535,In_21,In_1630);
and U1536 (N_1536,In_2008,In_1355);
and U1537 (N_1537,In_942,In_120);
nor U1538 (N_1538,In_523,In_413);
or U1539 (N_1539,In_1587,In_1585);
nor U1540 (N_1540,In_1905,In_2357);
xnor U1541 (N_1541,In_1238,In_285);
nand U1542 (N_1542,In_944,In_1710);
nor U1543 (N_1543,In_1339,In_972);
and U1544 (N_1544,In_68,In_1030);
nor U1545 (N_1545,In_1660,In_686);
and U1546 (N_1546,In_2229,In_2366);
and U1547 (N_1547,In_1566,In_576);
nand U1548 (N_1548,In_1277,In_2362);
or U1549 (N_1549,In_1144,In_2180);
and U1550 (N_1550,In_1945,In_1128);
nor U1551 (N_1551,In_101,In_835);
nor U1552 (N_1552,In_428,In_1516);
nor U1553 (N_1553,In_278,In_996);
nand U1554 (N_1554,In_309,In_2179);
nand U1555 (N_1555,In_1695,In_2168);
and U1556 (N_1556,In_500,In_1807);
and U1557 (N_1557,In_1914,In_591);
or U1558 (N_1558,In_1057,In_193);
nand U1559 (N_1559,In_1758,In_1656);
and U1560 (N_1560,In_1429,In_354);
nor U1561 (N_1561,In_337,In_549);
and U1562 (N_1562,In_2335,In_917);
nor U1563 (N_1563,In_414,In_1290);
and U1564 (N_1564,In_59,In_2123);
nor U1565 (N_1565,In_2491,In_1548);
nand U1566 (N_1566,In_1913,In_1151);
nand U1567 (N_1567,In_2175,In_2168);
nor U1568 (N_1568,In_297,In_1964);
or U1569 (N_1569,In_2006,In_2285);
and U1570 (N_1570,In_1549,In_107);
nand U1571 (N_1571,In_867,In_2091);
nand U1572 (N_1572,In_1811,In_1036);
and U1573 (N_1573,In_1535,In_2314);
nand U1574 (N_1574,In_691,In_671);
or U1575 (N_1575,In_132,In_1971);
nor U1576 (N_1576,In_1396,In_966);
and U1577 (N_1577,In_2007,In_2427);
and U1578 (N_1578,In_2090,In_4);
nand U1579 (N_1579,In_55,In_1339);
nor U1580 (N_1580,In_3,In_934);
nor U1581 (N_1581,In_2011,In_726);
and U1582 (N_1582,In_2211,In_1504);
and U1583 (N_1583,In_1939,In_448);
nand U1584 (N_1584,In_2135,In_1458);
nor U1585 (N_1585,In_354,In_2437);
and U1586 (N_1586,In_1410,In_1567);
and U1587 (N_1587,In_1348,In_731);
nor U1588 (N_1588,In_359,In_1007);
nand U1589 (N_1589,In_1167,In_1416);
nand U1590 (N_1590,In_1641,In_1170);
or U1591 (N_1591,In_2396,In_32);
and U1592 (N_1592,In_1855,In_269);
nor U1593 (N_1593,In_880,In_295);
or U1594 (N_1594,In_1887,In_2447);
or U1595 (N_1595,In_1151,In_1773);
nand U1596 (N_1596,In_956,In_416);
xnor U1597 (N_1597,In_765,In_1917);
xnor U1598 (N_1598,In_1332,In_560);
or U1599 (N_1599,In_447,In_1742);
or U1600 (N_1600,In_1741,In_499);
or U1601 (N_1601,In_2208,In_94);
nor U1602 (N_1602,In_653,In_197);
and U1603 (N_1603,In_1109,In_1561);
and U1604 (N_1604,In_742,In_1703);
nand U1605 (N_1605,In_273,In_2380);
and U1606 (N_1606,In_1450,In_2491);
nand U1607 (N_1607,In_691,In_2195);
or U1608 (N_1608,In_2481,In_1962);
and U1609 (N_1609,In_1999,In_1732);
and U1610 (N_1610,In_339,In_2054);
nor U1611 (N_1611,In_2415,In_6);
nand U1612 (N_1612,In_1151,In_2198);
nand U1613 (N_1613,In_406,In_1357);
and U1614 (N_1614,In_845,In_1362);
and U1615 (N_1615,In_2422,In_1534);
or U1616 (N_1616,In_131,In_530);
nand U1617 (N_1617,In_1940,In_1814);
or U1618 (N_1618,In_343,In_1036);
and U1619 (N_1619,In_1838,In_1675);
xnor U1620 (N_1620,In_966,In_54);
and U1621 (N_1621,In_1511,In_507);
or U1622 (N_1622,In_2106,In_1506);
and U1623 (N_1623,In_1635,In_1069);
nand U1624 (N_1624,In_1875,In_619);
nand U1625 (N_1625,In_1091,In_414);
and U1626 (N_1626,In_1713,In_1077);
and U1627 (N_1627,In_2393,In_1204);
and U1628 (N_1628,In_1799,In_2129);
nand U1629 (N_1629,In_1709,In_1597);
or U1630 (N_1630,In_1494,In_699);
xnor U1631 (N_1631,In_1348,In_2112);
xnor U1632 (N_1632,In_1612,In_1069);
nand U1633 (N_1633,In_445,In_1173);
nor U1634 (N_1634,In_448,In_579);
nor U1635 (N_1635,In_1111,In_150);
nor U1636 (N_1636,In_1465,In_2396);
xnor U1637 (N_1637,In_480,In_2078);
and U1638 (N_1638,In_153,In_785);
and U1639 (N_1639,In_227,In_1994);
nand U1640 (N_1640,In_822,In_870);
nor U1641 (N_1641,In_1693,In_465);
and U1642 (N_1642,In_1639,In_1641);
xnor U1643 (N_1643,In_1093,In_660);
nand U1644 (N_1644,In_1405,In_972);
nand U1645 (N_1645,In_2114,In_1262);
nand U1646 (N_1646,In_1944,In_1676);
or U1647 (N_1647,In_82,In_1165);
xor U1648 (N_1648,In_842,In_1056);
nand U1649 (N_1649,In_1247,In_2156);
and U1650 (N_1650,In_1462,In_1806);
nor U1651 (N_1651,In_2366,In_301);
and U1652 (N_1652,In_492,In_1130);
and U1653 (N_1653,In_125,In_298);
or U1654 (N_1654,In_1895,In_155);
nand U1655 (N_1655,In_1304,In_1758);
nor U1656 (N_1656,In_707,In_2030);
nor U1657 (N_1657,In_856,In_1705);
and U1658 (N_1658,In_1866,In_1591);
xor U1659 (N_1659,In_1662,In_217);
nand U1660 (N_1660,In_2358,In_1104);
nor U1661 (N_1661,In_657,In_263);
nand U1662 (N_1662,In_99,In_328);
or U1663 (N_1663,In_72,In_1821);
and U1664 (N_1664,In_2181,In_1737);
or U1665 (N_1665,In_653,In_1380);
nor U1666 (N_1666,In_1065,In_740);
or U1667 (N_1667,In_1040,In_569);
nor U1668 (N_1668,In_850,In_1263);
nor U1669 (N_1669,In_1212,In_1271);
nand U1670 (N_1670,In_1851,In_573);
nor U1671 (N_1671,In_2276,In_1440);
and U1672 (N_1672,In_1485,In_1347);
nand U1673 (N_1673,In_1052,In_1689);
nand U1674 (N_1674,In_398,In_1340);
and U1675 (N_1675,In_113,In_2434);
or U1676 (N_1676,In_1119,In_1730);
xnor U1677 (N_1677,In_634,In_2230);
nand U1678 (N_1678,In_363,In_1132);
or U1679 (N_1679,In_2360,In_1253);
or U1680 (N_1680,In_1821,In_2482);
and U1681 (N_1681,In_592,In_1408);
and U1682 (N_1682,In_1500,In_568);
nor U1683 (N_1683,In_2349,In_1723);
or U1684 (N_1684,In_454,In_2394);
or U1685 (N_1685,In_1237,In_1660);
nand U1686 (N_1686,In_1347,In_294);
and U1687 (N_1687,In_1755,In_1275);
nor U1688 (N_1688,In_2125,In_473);
or U1689 (N_1689,In_2148,In_1559);
or U1690 (N_1690,In_1187,In_466);
nand U1691 (N_1691,In_1558,In_2126);
nand U1692 (N_1692,In_282,In_2023);
or U1693 (N_1693,In_1914,In_1274);
nor U1694 (N_1694,In_1922,In_232);
or U1695 (N_1695,In_2319,In_1241);
nand U1696 (N_1696,In_1283,In_1910);
or U1697 (N_1697,In_2009,In_332);
nor U1698 (N_1698,In_2290,In_2369);
nor U1699 (N_1699,In_1609,In_2001);
or U1700 (N_1700,In_0,In_524);
nor U1701 (N_1701,In_453,In_1774);
or U1702 (N_1702,In_1349,In_940);
xor U1703 (N_1703,In_1091,In_70);
or U1704 (N_1704,In_1452,In_795);
nand U1705 (N_1705,In_2422,In_732);
or U1706 (N_1706,In_1048,In_1066);
xor U1707 (N_1707,In_615,In_6);
or U1708 (N_1708,In_828,In_678);
xnor U1709 (N_1709,In_1309,In_1095);
nand U1710 (N_1710,In_77,In_2226);
nor U1711 (N_1711,In_1580,In_587);
nand U1712 (N_1712,In_1451,In_1507);
or U1713 (N_1713,In_1496,In_2088);
nand U1714 (N_1714,In_1058,In_1559);
xor U1715 (N_1715,In_1620,In_793);
nor U1716 (N_1716,In_1987,In_2314);
nand U1717 (N_1717,In_2428,In_2175);
and U1718 (N_1718,In_2438,In_2068);
or U1719 (N_1719,In_610,In_1599);
nor U1720 (N_1720,In_1031,In_1436);
nor U1721 (N_1721,In_1990,In_1543);
nor U1722 (N_1722,In_1781,In_1281);
nor U1723 (N_1723,In_2200,In_1978);
or U1724 (N_1724,In_1954,In_2112);
nor U1725 (N_1725,In_1501,In_681);
or U1726 (N_1726,In_1603,In_2406);
xor U1727 (N_1727,In_1237,In_1762);
xnor U1728 (N_1728,In_1091,In_1856);
and U1729 (N_1729,In_760,In_386);
xor U1730 (N_1730,In_2069,In_152);
nor U1731 (N_1731,In_1675,In_196);
nor U1732 (N_1732,In_1098,In_2099);
nor U1733 (N_1733,In_710,In_666);
nor U1734 (N_1734,In_2111,In_961);
nand U1735 (N_1735,In_1773,In_1024);
or U1736 (N_1736,In_295,In_602);
and U1737 (N_1737,In_2297,In_1538);
or U1738 (N_1738,In_1440,In_1108);
nand U1739 (N_1739,In_1753,In_657);
xnor U1740 (N_1740,In_2292,In_1115);
nand U1741 (N_1741,In_1155,In_1562);
and U1742 (N_1742,In_621,In_2212);
and U1743 (N_1743,In_711,In_411);
and U1744 (N_1744,In_533,In_1815);
nor U1745 (N_1745,In_1138,In_1335);
nand U1746 (N_1746,In_1356,In_2353);
nand U1747 (N_1747,In_1514,In_673);
xor U1748 (N_1748,In_1724,In_1785);
or U1749 (N_1749,In_1210,In_392);
or U1750 (N_1750,In_2268,In_2134);
and U1751 (N_1751,In_1537,In_484);
nor U1752 (N_1752,In_2406,In_281);
and U1753 (N_1753,In_1809,In_2129);
nand U1754 (N_1754,In_2493,In_36);
or U1755 (N_1755,In_553,In_1953);
and U1756 (N_1756,In_916,In_1482);
or U1757 (N_1757,In_1510,In_1043);
nand U1758 (N_1758,In_1344,In_517);
xnor U1759 (N_1759,In_554,In_384);
nand U1760 (N_1760,In_2029,In_504);
nor U1761 (N_1761,In_85,In_727);
nor U1762 (N_1762,In_101,In_2189);
and U1763 (N_1763,In_468,In_1913);
or U1764 (N_1764,In_644,In_1839);
nor U1765 (N_1765,In_2446,In_2381);
and U1766 (N_1766,In_2178,In_2354);
xnor U1767 (N_1767,In_1571,In_2143);
and U1768 (N_1768,In_954,In_847);
or U1769 (N_1769,In_870,In_1267);
or U1770 (N_1770,In_994,In_1209);
or U1771 (N_1771,In_51,In_2079);
and U1772 (N_1772,In_1200,In_894);
nand U1773 (N_1773,In_554,In_447);
nor U1774 (N_1774,In_530,In_910);
and U1775 (N_1775,In_1409,In_2063);
nand U1776 (N_1776,In_709,In_439);
nor U1777 (N_1777,In_1125,In_948);
nand U1778 (N_1778,In_2412,In_1086);
nor U1779 (N_1779,In_953,In_666);
xnor U1780 (N_1780,In_1442,In_675);
and U1781 (N_1781,In_1317,In_2238);
xor U1782 (N_1782,In_1879,In_1304);
nor U1783 (N_1783,In_554,In_1064);
or U1784 (N_1784,In_1241,In_724);
nor U1785 (N_1785,In_1641,In_457);
or U1786 (N_1786,In_91,In_1053);
nor U1787 (N_1787,In_1193,In_1868);
or U1788 (N_1788,In_353,In_256);
nand U1789 (N_1789,In_1140,In_2398);
nor U1790 (N_1790,In_605,In_528);
or U1791 (N_1791,In_702,In_2488);
nand U1792 (N_1792,In_2393,In_2007);
nand U1793 (N_1793,In_222,In_1926);
nand U1794 (N_1794,In_246,In_2378);
nand U1795 (N_1795,In_341,In_635);
or U1796 (N_1796,In_1991,In_517);
or U1797 (N_1797,In_32,In_1398);
nand U1798 (N_1798,In_2265,In_1594);
xor U1799 (N_1799,In_1156,In_2234);
and U1800 (N_1800,In_2090,In_1640);
nor U1801 (N_1801,In_1823,In_451);
nor U1802 (N_1802,In_352,In_726);
nor U1803 (N_1803,In_2077,In_1873);
or U1804 (N_1804,In_388,In_577);
and U1805 (N_1805,In_1771,In_1529);
or U1806 (N_1806,In_1047,In_1577);
nand U1807 (N_1807,In_1548,In_1900);
nand U1808 (N_1808,In_2290,In_1735);
or U1809 (N_1809,In_362,In_103);
nor U1810 (N_1810,In_765,In_372);
xnor U1811 (N_1811,In_2260,In_1819);
nor U1812 (N_1812,In_1926,In_432);
nor U1813 (N_1813,In_652,In_1072);
or U1814 (N_1814,In_164,In_342);
nand U1815 (N_1815,In_308,In_2326);
or U1816 (N_1816,In_1018,In_891);
and U1817 (N_1817,In_890,In_1638);
nor U1818 (N_1818,In_1495,In_225);
and U1819 (N_1819,In_64,In_856);
nor U1820 (N_1820,In_2306,In_1426);
or U1821 (N_1821,In_1082,In_259);
and U1822 (N_1822,In_2318,In_718);
nor U1823 (N_1823,In_1706,In_491);
and U1824 (N_1824,In_222,In_1590);
and U1825 (N_1825,In_1428,In_1882);
or U1826 (N_1826,In_1764,In_1373);
nand U1827 (N_1827,In_370,In_542);
and U1828 (N_1828,In_344,In_1933);
nor U1829 (N_1829,In_1379,In_829);
or U1830 (N_1830,In_1855,In_2379);
and U1831 (N_1831,In_297,In_88);
xnor U1832 (N_1832,In_409,In_612);
or U1833 (N_1833,In_542,In_1191);
nand U1834 (N_1834,In_2343,In_1371);
or U1835 (N_1835,In_2210,In_2066);
xnor U1836 (N_1836,In_341,In_2298);
or U1837 (N_1837,In_1297,In_939);
nand U1838 (N_1838,In_1580,In_167);
and U1839 (N_1839,In_116,In_1790);
and U1840 (N_1840,In_2229,In_1695);
nor U1841 (N_1841,In_1207,In_1261);
and U1842 (N_1842,In_2399,In_1923);
or U1843 (N_1843,In_2330,In_651);
nor U1844 (N_1844,In_1539,In_571);
and U1845 (N_1845,In_1988,In_2254);
or U1846 (N_1846,In_495,In_2137);
nor U1847 (N_1847,In_769,In_1208);
nand U1848 (N_1848,In_2007,In_688);
or U1849 (N_1849,In_419,In_2026);
nor U1850 (N_1850,In_1663,In_1130);
or U1851 (N_1851,In_2063,In_173);
nand U1852 (N_1852,In_1843,In_1491);
and U1853 (N_1853,In_2394,In_970);
or U1854 (N_1854,In_406,In_1474);
nor U1855 (N_1855,In_1965,In_2152);
and U1856 (N_1856,In_472,In_1764);
nor U1857 (N_1857,In_724,In_1364);
or U1858 (N_1858,In_2056,In_1354);
or U1859 (N_1859,In_2387,In_1700);
and U1860 (N_1860,In_1568,In_828);
xor U1861 (N_1861,In_716,In_1772);
nor U1862 (N_1862,In_729,In_746);
or U1863 (N_1863,In_1454,In_1046);
or U1864 (N_1864,In_1903,In_2158);
nand U1865 (N_1865,In_1732,In_1917);
nor U1866 (N_1866,In_458,In_1311);
nor U1867 (N_1867,In_1223,In_2254);
and U1868 (N_1868,In_408,In_2062);
nor U1869 (N_1869,In_2083,In_2134);
nor U1870 (N_1870,In_191,In_917);
nor U1871 (N_1871,In_305,In_1477);
or U1872 (N_1872,In_954,In_1103);
nand U1873 (N_1873,In_1707,In_114);
or U1874 (N_1874,In_622,In_2030);
or U1875 (N_1875,In_1662,In_275);
xor U1876 (N_1876,In_918,In_2257);
nand U1877 (N_1877,In_2124,In_704);
nand U1878 (N_1878,In_45,In_623);
and U1879 (N_1879,In_2319,In_1386);
nor U1880 (N_1880,In_764,In_2402);
xor U1881 (N_1881,In_2089,In_678);
and U1882 (N_1882,In_1007,In_850);
nand U1883 (N_1883,In_1767,In_669);
or U1884 (N_1884,In_1164,In_2082);
and U1885 (N_1885,In_2111,In_2156);
nor U1886 (N_1886,In_228,In_2055);
or U1887 (N_1887,In_22,In_1580);
xnor U1888 (N_1888,In_1395,In_2473);
and U1889 (N_1889,In_695,In_409);
or U1890 (N_1890,In_321,In_953);
or U1891 (N_1891,In_1823,In_1279);
nor U1892 (N_1892,In_842,In_210);
nand U1893 (N_1893,In_624,In_996);
nor U1894 (N_1894,In_1840,In_1723);
or U1895 (N_1895,In_1127,In_363);
and U1896 (N_1896,In_327,In_2474);
and U1897 (N_1897,In_33,In_524);
nor U1898 (N_1898,In_881,In_2037);
nand U1899 (N_1899,In_1883,In_316);
and U1900 (N_1900,In_889,In_1526);
or U1901 (N_1901,In_559,In_2370);
nand U1902 (N_1902,In_297,In_13);
nor U1903 (N_1903,In_1802,In_790);
or U1904 (N_1904,In_22,In_1671);
or U1905 (N_1905,In_1726,In_1993);
nand U1906 (N_1906,In_1253,In_2218);
nor U1907 (N_1907,In_1011,In_2047);
xor U1908 (N_1908,In_1216,In_1936);
nor U1909 (N_1909,In_1442,In_644);
or U1910 (N_1910,In_655,In_562);
nor U1911 (N_1911,In_112,In_396);
nor U1912 (N_1912,In_2448,In_2309);
nand U1913 (N_1913,In_2284,In_2486);
nand U1914 (N_1914,In_1269,In_747);
nor U1915 (N_1915,In_1294,In_1710);
and U1916 (N_1916,In_147,In_1040);
nand U1917 (N_1917,In_1753,In_624);
nor U1918 (N_1918,In_1459,In_2228);
nand U1919 (N_1919,In_2002,In_2058);
nor U1920 (N_1920,In_1407,In_2047);
nor U1921 (N_1921,In_1718,In_317);
nor U1922 (N_1922,In_815,In_1684);
nand U1923 (N_1923,In_1946,In_84);
and U1924 (N_1924,In_819,In_1102);
or U1925 (N_1925,In_1696,In_912);
and U1926 (N_1926,In_129,In_2468);
nand U1927 (N_1927,In_688,In_1632);
and U1928 (N_1928,In_489,In_1283);
nor U1929 (N_1929,In_869,In_717);
nand U1930 (N_1930,In_2174,In_2292);
nor U1931 (N_1931,In_568,In_1600);
nand U1932 (N_1932,In_98,In_1490);
nand U1933 (N_1933,In_1381,In_2127);
nor U1934 (N_1934,In_2170,In_86);
or U1935 (N_1935,In_2359,In_927);
or U1936 (N_1936,In_456,In_1681);
or U1937 (N_1937,In_2006,In_479);
nor U1938 (N_1938,In_10,In_2010);
nor U1939 (N_1939,In_1901,In_2451);
nand U1940 (N_1940,In_1644,In_1601);
xnor U1941 (N_1941,In_944,In_1813);
xnor U1942 (N_1942,In_905,In_1639);
nand U1943 (N_1943,In_1126,In_1018);
nand U1944 (N_1944,In_520,In_1346);
nand U1945 (N_1945,In_893,In_2349);
nor U1946 (N_1946,In_2061,In_1809);
or U1947 (N_1947,In_1476,In_1824);
or U1948 (N_1948,In_1414,In_222);
nand U1949 (N_1949,In_350,In_2151);
nand U1950 (N_1950,In_551,In_1670);
or U1951 (N_1951,In_127,In_1394);
xor U1952 (N_1952,In_1276,In_1006);
or U1953 (N_1953,In_2401,In_1196);
or U1954 (N_1954,In_2417,In_811);
xor U1955 (N_1955,In_885,In_2017);
nand U1956 (N_1956,In_792,In_688);
or U1957 (N_1957,In_2164,In_1765);
or U1958 (N_1958,In_408,In_228);
and U1959 (N_1959,In_1163,In_2200);
or U1960 (N_1960,In_1545,In_1883);
nand U1961 (N_1961,In_645,In_2264);
nor U1962 (N_1962,In_1091,In_2238);
and U1963 (N_1963,In_2222,In_1354);
nand U1964 (N_1964,In_691,In_2272);
and U1965 (N_1965,In_1839,In_461);
xor U1966 (N_1966,In_867,In_957);
and U1967 (N_1967,In_128,In_69);
and U1968 (N_1968,In_2177,In_456);
or U1969 (N_1969,In_1462,In_332);
and U1970 (N_1970,In_1495,In_303);
or U1971 (N_1971,In_689,In_2087);
and U1972 (N_1972,In_1682,In_1818);
nor U1973 (N_1973,In_1761,In_578);
or U1974 (N_1974,In_2080,In_2075);
nand U1975 (N_1975,In_1936,In_2024);
or U1976 (N_1976,In_104,In_784);
and U1977 (N_1977,In_1518,In_548);
nor U1978 (N_1978,In_1289,In_127);
and U1979 (N_1979,In_548,In_1693);
or U1980 (N_1980,In_1373,In_1040);
nand U1981 (N_1981,In_1403,In_1885);
nand U1982 (N_1982,In_676,In_45);
xor U1983 (N_1983,In_1990,In_1447);
and U1984 (N_1984,In_1930,In_1049);
nor U1985 (N_1985,In_2347,In_819);
xor U1986 (N_1986,In_2235,In_1811);
and U1987 (N_1987,In_890,In_1968);
nor U1988 (N_1988,In_1723,In_1075);
or U1989 (N_1989,In_2306,In_803);
or U1990 (N_1990,In_1273,In_2240);
nor U1991 (N_1991,In_493,In_830);
xor U1992 (N_1992,In_2090,In_1746);
nor U1993 (N_1993,In_107,In_2006);
nand U1994 (N_1994,In_875,In_1755);
nor U1995 (N_1995,In_1827,In_488);
nor U1996 (N_1996,In_1387,In_1659);
and U1997 (N_1997,In_1312,In_1145);
or U1998 (N_1998,In_531,In_117);
nand U1999 (N_1999,In_733,In_488);
nor U2000 (N_2000,In_53,In_1866);
and U2001 (N_2001,In_1360,In_1276);
nor U2002 (N_2002,In_2074,In_1515);
and U2003 (N_2003,In_1437,In_860);
nand U2004 (N_2004,In_1476,In_1955);
xnor U2005 (N_2005,In_711,In_925);
nand U2006 (N_2006,In_918,In_908);
or U2007 (N_2007,In_1629,In_1357);
and U2008 (N_2008,In_1207,In_1966);
or U2009 (N_2009,In_282,In_2494);
nand U2010 (N_2010,In_1369,In_1665);
xor U2011 (N_2011,In_238,In_2011);
xnor U2012 (N_2012,In_958,In_1985);
and U2013 (N_2013,In_1245,In_2406);
and U2014 (N_2014,In_800,In_2340);
or U2015 (N_2015,In_546,In_250);
xor U2016 (N_2016,In_2302,In_1578);
or U2017 (N_2017,In_1566,In_834);
and U2018 (N_2018,In_742,In_752);
nand U2019 (N_2019,In_512,In_1824);
nor U2020 (N_2020,In_913,In_1603);
nand U2021 (N_2021,In_746,In_1938);
and U2022 (N_2022,In_29,In_1982);
or U2023 (N_2023,In_1010,In_1356);
xnor U2024 (N_2024,In_1252,In_989);
nor U2025 (N_2025,In_2352,In_1214);
or U2026 (N_2026,In_357,In_1287);
nand U2027 (N_2027,In_384,In_1726);
and U2028 (N_2028,In_1764,In_1074);
and U2029 (N_2029,In_1916,In_497);
and U2030 (N_2030,In_1673,In_981);
or U2031 (N_2031,In_12,In_99);
nor U2032 (N_2032,In_2373,In_164);
or U2033 (N_2033,In_1302,In_213);
or U2034 (N_2034,In_874,In_801);
or U2035 (N_2035,In_840,In_383);
nand U2036 (N_2036,In_1984,In_1084);
and U2037 (N_2037,In_348,In_214);
xnor U2038 (N_2038,In_837,In_1422);
or U2039 (N_2039,In_475,In_632);
nand U2040 (N_2040,In_2190,In_1204);
or U2041 (N_2041,In_2136,In_1232);
xor U2042 (N_2042,In_1534,In_1885);
nor U2043 (N_2043,In_1460,In_955);
or U2044 (N_2044,In_1019,In_219);
nor U2045 (N_2045,In_1108,In_2483);
nor U2046 (N_2046,In_530,In_2068);
nor U2047 (N_2047,In_494,In_240);
or U2048 (N_2048,In_1347,In_2262);
or U2049 (N_2049,In_2267,In_885);
nor U2050 (N_2050,In_1992,In_2396);
and U2051 (N_2051,In_169,In_1559);
or U2052 (N_2052,In_1623,In_1392);
nor U2053 (N_2053,In_1674,In_1404);
nand U2054 (N_2054,In_712,In_1568);
or U2055 (N_2055,In_852,In_542);
nor U2056 (N_2056,In_856,In_2173);
nand U2057 (N_2057,In_1058,In_173);
and U2058 (N_2058,In_1507,In_138);
or U2059 (N_2059,In_1681,In_407);
or U2060 (N_2060,In_2470,In_2133);
nor U2061 (N_2061,In_1217,In_103);
nand U2062 (N_2062,In_2389,In_2243);
nand U2063 (N_2063,In_1696,In_176);
nor U2064 (N_2064,In_1420,In_1367);
or U2065 (N_2065,In_824,In_1259);
or U2066 (N_2066,In_185,In_1981);
and U2067 (N_2067,In_1402,In_547);
and U2068 (N_2068,In_1516,In_2348);
nand U2069 (N_2069,In_1882,In_1441);
nand U2070 (N_2070,In_366,In_1552);
nand U2071 (N_2071,In_1528,In_903);
nand U2072 (N_2072,In_1012,In_1113);
nand U2073 (N_2073,In_1247,In_2022);
nor U2074 (N_2074,In_1677,In_1759);
nor U2075 (N_2075,In_1908,In_1618);
or U2076 (N_2076,In_1024,In_1523);
nand U2077 (N_2077,In_886,In_872);
nor U2078 (N_2078,In_1325,In_103);
nor U2079 (N_2079,In_2344,In_1178);
nand U2080 (N_2080,In_1264,In_631);
or U2081 (N_2081,In_1945,In_342);
or U2082 (N_2082,In_1761,In_962);
and U2083 (N_2083,In_2067,In_335);
xnor U2084 (N_2084,In_1255,In_2226);
nor U2085 (N_2085,In_2007,In_2373);
xnor U2086 (N_2086,In_1026,In_698);
nand U2087 (N_2087,In_2195,In_2068);
nand U2088 (N_2088,In_60,In_1471);
or U2089 (N_2089,In_2334,In_1524);
and U2090 (N_2090,In_686,In_65);
nor U2091 (N_2091,In_1724,In_1583);
or U2092 (N_2092,In_443,In_926);
or U2093 (N_2093,In_828,In_1365);
or U2094 (N_2094,In_836,In_172);
and U2095 (N_2095,In_576,In_1432);
nor U2096 (N_2096,In_2003,In_133);
and U2097 (N_2097,In_889,In_68);
nor U2098 (N_2098,In_1599,In_961);
xor U2099 (N_2099,In_920,In_2027);
and U2100 (N_2100,In_276,In_1839);
and U2101 (N_2101,In_2056,In_1493);
nor U2102 (N_2102,In_1940,In_2409);
and U2103 (N_2103,In_2476,In_174);
xnor U2104 (N_2104,In_1386,In_1250);
nor U2105 (N_2105,In_1007,In_1911);
nor U2106 (N_2106,In_1364,In_1455);
nor U2107 (N_2107,In_2231,In_779);
and U2108 (N_2108,In_1699,In_539);
nor U2109 (N_2109,In_2469,In_1773);
nor U2110 (N_2110,In_1253,In_880);
xor U2111 (N_2111,In_2115,In_2026);
nand U2112 (N_2112,In_2277,In_1959);
or U2113 (N_2113,In_298,In_1816);
and U2114 (N_2114,In_744,In_974);
nor U2115 (N_2115,In_1885,In_2366);
and U2116 (N_2116,In_1266,In_669);
xor U2117 (N_2117,In_507,In_787);
nand U2118 (N_2118,In_39,In_2426);
or U2119 (N_2119,In_2169,In_1987);
and U2120 (N_2120,In_192,In_152);
nor U2121 (N_2121,In_1312,In_674);
and U2122 (N_2122,In_2097,In_1795);
and U2123 (N_2123,In_2428,In_1709);
and U2124 (N_2124,In_245,In_1015);
or U2125 (N_2125,In_722,In_277);
or U2126 (N_2126,In_718,In_669);
or U2127 (N_2127,In_1234,In_599);
nor U2128 (N_2128,In_1531,In_1976);
nor U2129 (N_2129,In_1645,In_875);
nand U2130 (N_2130,In_51,In_1167);
nand U2131 (N_2131,In_1677,In_1792);
and U2132 (N_2132,In_521,In_1253);
or U2133 (N_2133,In_1742,In_663);
nand U2134 (N_2134,In_1101,In_920);
nor U2135 (N_2135,In_1625,In_1908);
nand U2136 (N_2136,In_856,In_1534);
and U2137 (N_2137,In_1659,In_1763);
nor U2138 (N_2138,In_326,In_2062);
nor U2139 (N_2139,In_2147,In_1219);
or U2140 (N_2140,In_1227,In_1140);
and U2141 (N_2141,In_2028,In_794);
nor U2142 (N_2142,In_72,In_1580);
nor U2143 (N_2143,In_263,In_1281);
or U2144 (N_2144,In_1617,In_880);
nor U2145 (N_2145,In_65,In_1362);
nand U2146 (N_2146,In_1346,In_380);
nor U2147 (N_2147,In_104,In_1982);
and U2148 (N_2148,In_1914,In_1849);
or U2149 (N_2149,In_1789,In_1308);
and U2150 (N_2150,In_2467,In_232);
nor U2151 (N_2151,In_471,In_2072);
nor U2152 (N_2152,In_2293,In_626);
xor U2153 (N_2153,In_2213,In_462);
nand U2154 (N_2154,In_1923,In_1357);
or U2155 (N_2155,In_1459,In_76);
nor U2156 (N_2156,In_1639,In_1140);
nor U2157 (N_2157,In_309,In_1007);
nand U2158 (N_2158,In_889,In_108);
nor U2159 (N_2159,In_1647,In_100);
nor U2160 (N_2160,In_229,In_1419);
or U2161 (N_2161,In_1347,In_6);
or U2162 (N_2162,In_763,In_431);
nand U2163 (N_2163,In_1455,In_1493);
and U2164 (N_2164,In_2098,In_333);
nand U2165 (N_2165,In_1029,In_486);
and U2166 (N_2166,In_1570,In_2000);
xnor U2167 (N_2167,In_1440,In_1228);
xor U2168 (N_2168,In_260,In_1863);
nand U2169 (N_2169,In_752,In_2028);
xnor U2170 (N_2170,In_511,In_2389);
nand U2171 (N_2171,In_420,In_1719);
and U2172 (N_2172,In_2381,In_2335);
or U2173 (N_2173,In_898,In_305);
or U2174 (N_2174,In_68,In_724);
or U2175 (N_2175,In_591,In_209);
or U2176 (N_2176,In_982,In_28);
nand U2177 (N_2177,In_2241,In_677);
nor U2178 (N_2178,In_1166,In_2310);
nand U2179 (N_2179,In_781,In_306);
and U2180 (N_2180,In_1984,In_1699);
or U2181 (N_2181,In_2283,In_20);
nor U2182 (N_2182,In_634,In_2112);
nand U2183 (N_2183,In_1576,In_2105);
nor U2184 (N_2184,In_1270,In_2400);
and U2185 (N_2185,In_871,In_2330);
nand U2186 (N_2186,In_2442,In_866);
nand U2187 (N_2187,In_1996,In_2280);
or U2188 (N_2188,In_17,In_1209);
and U2189 (N_2189,In_1644,In_1836);
or U2190 (N_2190,In_467,In_1255);
and U2191 (N_2191,In_284,In_1312);
nand U2192 (N_2192,In_188,In_1543);
nand U2193 (N_2193,In_680,In_921);
nor U2194 (N_2194,In_704,In_415);
nand U2195 (N_2195,In_2130,In_61);
and U2196 (N_2196,In_185,In_149);
and U2197 (N_2197,In_2264,In_2419);
nor U2198 (N_2198,In_77,In_1340);
nand U2199 (N_2199,In_2253,In_1854);
xnor U2200 (N_2200,In_375,In_1005);
nand U2201 (N_2201,In_6,In_41);
and U2202 (N_2202,In_414,In_2395);
and U2203 (N_2203,In_2038,In_1203);
nand U2204 (N_2204,In_2248,In_2458);
nand U2205 (N_2205,In_1269,In_782);
and U2206 (N_2206,In_800,In_873);
nand U2207 (N_2207,In_665,In_1328);
nor U2208 (N_2208,In_850,In_2450);
nor U2209 (N_2209,In_886,In_2002);
nor U2210 (N_2210,In_1457,In_1402);
and U2211 (N_2211,In_2125,In_1829);
nand U2212 (N_2212,In_485,In_1399);
xnor U2213 (N_2213,In_2224,In_1148);
nand U2214 (N_2214,In_1181,In_2028);
xnor U2215 (N_2215,In_696,In_2399);
xor U2216 (N_2216,In_2049,In_898);
nor U2217 (N_2217,In_1005,In_2020);
or U2218 (N_2218,In_1501,In_627);
and U2219 (N_2219,In_1155,In_1591);
nand U2220 (N_2220,In_218,In_872);
nand U2221 (N_2221,In_984,In_1654);
and U2222 (N_2222,In_1004,In_2120);
or U2223 (N_2223,In_1263,In_1074);
and U2224 (N_2224,In_2269,In_809);
and U2225 (N_2225,In_884,In_2138);
nand U2226 (N_2226,In_294,In_1211);
or U2227 (N_2227,In_1499,In_1449);
nand U2228 (N_2228,In_2147,In_311);
and U2229 (N_2229,In_1146,In_1882);
xnor U2230 (N_2230,In_1788,In_2217);
or U2231 (N_2231,In_1373,In_1514);
and U2232 (N_2232,In_1764,In_805);
or U2233 (N_2233,In_1256,In_1900);
or U2234 (N_2234,In_1380,In_2181);
nor U2235 (N_2235,In_816,In_2181);
xor U2236 (N_2236,In_424,In_1246);
nor U2237 (N_2237,In_2365,In_193);
and U2238 (N_2238,In_937,In_101);
or U2239 (N_2239,In_2363,In_682);
nor U2240 (N_2240,In_155,In_950);
or U2241 (N_2241,In_1857,In_1649);
or U2242 (N_2242,In_99,In_1025);
nor U2243 (N_2243,In_1710,In_2321);
or U2244 (N_2244,In_1596,In_1886);
nor U2245 (N_2245,In_1323,In_1025);
nand U2246 (N_2246,In_2087,In_973);
and U2247 (N_2247,In_2403,In_2103);
and U2248 (N_2248,In_681,In_719);
or U2249 (N_2249,In_1282,In_634);
or U2250 (N_2250,In_2163,In_521);
nor U2251 (N_2251,In_1740,In_2090);
nand U2252 (N_2252,In_2162,In_680);
or U2253 (N_2253,In_44,In_297);
nand U2254 (N_2254,In_2382,In_2423);
or U2255 (N_2255,In_2237,In_611);
nor U2256 (N_2256,In_2280,In_1804);
nand U2257 (N_2257,In_402,In_1706);
xor U2258 (N_2258,In_2447,In_795);
nand U2259 (N_2259,In_1082,In_2443);
or U2260 (N_2260,In_611,In_1181);
nand U2261 (N_2261,In_1975,In_873);
and U2262 (N_2262,In_863,In_1807);
or U2263 (N_2263,In_1066,In_1649);
nor U2264 (N_2264,In_2445,In_1708);
nor U2265 (N_2265,In_1761,In_2368);
or U2266 (N_2266,In_1069,In_659);
nand U2267 (N_2267,In_2318,In_437);
xor U2268 (N_2268,In_855,In_1956);
nor U2269 (N_2269,In_865,In_1111);
or U2270 (N_2270,In_1086,In_582);
nand U2271 (N_2271,In_1818,In_852);
nand U2272 (N_2272,In_827,In_1040);
or U2273 (N_2273,In_1023,In_1019);
nand U2274 (N_2274,In_1912,In_958);
or U2275 (N_2275,In_441,In_1860);
xor U2276 (N_2276,In_1809,In_29);
nor U2277 (N_2277,In_1658,In_626);
nor U2278 (N_2278,In_1232,In_861);
and U2279 (N_2279,In_1792,In_1616);
or U2280 (N_2280,In_653,In_651);
nand U2281 (N_2281,In_1636,In_526);
nor U2282 (N_2282,In_1812,In_772);
or U2283 (N_2283,In_676,In_1454);
nor U2284 (N_2284,In_50,In_337);
nor U2285 (N_2285,In_144,In_350);
nor U2286 (N_2286,In_1745,In_38);
nor U2287 (N_2287,In_815,In_1662);
and U2288 (N_2288,In_735,In_1954);
and U2289 (N_2289,In_2197,In_1501);
nand U2290 (N_2290,In_1611,In_875);
nand U2291 (N_2291,In_1845,In_499);
and U2292 (N_2292,In_633,In_599);
nor U2293 (N_2293,In_1884,In_2153);
or U2294 (N_2294,In_751,In_2308);
or U2295 (N_2295,In_301,In_1796);
nor U2296 (N_2296,In_1858,In_736);
or U2297 (N_2297,In_2062,In_364);
or U2298 (N_2298,In_988,In_2019);
nor U2299 (N_2299,In_969,In_1060);
and U2300 (N_2300,In_502,In_1021);
and U2301 (N_2301,In_1483,In_1720);
or U2302 (N_2302,In_495,In_1476);
nand U2303 (N_2303,In_1760,In_2107);
nor U2304 (N_2304,In_2260,In_164);
nand U2305 (N_2305,In_395,In_332);
nand U2306 (N_2306,In_504,In_1249);
nor U2307 (N_2307,In_513,In_688);
nor U2308 (N_2308,In_1209,In_1842);
nand U2309 (N_2309,In_2070,In_2365);
nor U2310 (N_2310,In_2057,In_9);
and U2311 (N_2311,In_518,In_1446);
xor U2312 (N_2312,In_905,In_540);
or U2313 (N_2313,In_1231,In_1194);
or U2314 (N_2314,In_2342,In_1136);
or U2315 (N_2315,In_26,In_1522);
and U2316 (N_2316,In_2398,In_2347);
and U2317 (N_2317,In_2025,In_678);
xnor U2318 (N_2318,In_814,In_318);
or U2319 (N_2319,In_414,In_2393);
nor U2320 (N_2320,In_582,In_2471);
xnor U2321 (N_2321,In_229,In_1240);
and U2322 (N_2322,In_537,In_146);
nand U2323 (N_2323,In_1109,In_793);
nor U2324 (N_2324,In_2453,In_1716);
or U2325 (N_2325,In_2218,In_823);
nor U2326 (N_2326,In_564,In_139);
or U2327 (N_2327,In_1371,In_251);
nand U2328 (N_2328,In_1176,In_1908);
nor U2329 (N_2329,In_2196,In_1218);
and U2330 (N_2330,In_150,In_702);
nand U2331 (N_2331,In_1486,In_600);
and U2332 (N_2332,In_2218,In_1748);
or U2333 (N_2333,In_1287,In_366);
and U2334 (N_2334,In_2080,In_722);
nand U2335 (N_2335,In_1847,In_1984);
and U2336 (N_2336,In_2408,In_714);
nor U2337 (N_2337,In_2072,In_1952);
and U2338 (N_2338,In_372,In_985);
nand U2339 (N_2339,In_2429,In_89);
nand U2340 (N_2340,In_75,In_728);
and U2341 (N_2341,In_56,In_1180);
nor U2342 (N_2342,In_335,In_1738);
xnor U2343 (N_2343,In_2259,In_2146);
nor U2344 (N_2344,In_1529,In_2359);
and U2345 (N_2345,In_604,In_383);
nor U2346 (N_2346,In_2211,In_940);
and U2347 (N_2347,In_1183,In_1441);
xnor U2348 (N_2348,In_1724,In_500);
or U2349 (N_2349,In_390,In_375);
nand U2350 (N_2350,In_335,In_232);
or U2351 (N_2351,In_612,In_184);
and U2352 (N_2352,In_1540,In_315);
or U2353 (N_2353,In_1532,In_43);
xnor U2354 (N_2354,In_700,In_2292);
nand U2355 (N_2355,In_2448,In_2473);
nor U2356 (N_2356,In_122,In_2245);
xnor U2357 (N_2357,In_753,In_241);
nand U2358 (N_2358,In_2375,In_1719);
and U2359 (N_2359,In_1717,In_2139);
and U2360 (N_2360,In_1736,In_890);
nor U2361 (N_2361,In_1767,In_1762);
and U2362 (N_2362,In_723,In_2079);
and U2363 (N_2363,In_2291,In_1000);
and U2364 (N_2364,In_1365,In_465);
nand U2365 (N_2365,In_267,In_1377);
and U2366 (N_2366,In_2425,In_305);
or U2367 (N_2367,In_1696,In_1908);
nor U2368 (N_2368,In_2493,In_1021);
xor U2369 (N_2369,In_672,In_785);
nor U2370 (N_2370,In_2110,In_1939);
nor U2371 (N_2371,In_1774,In_1708);
nand U2372 (N_2372,In_277,In_877);
xor U2373 (N_2373,In_1340,In_205);
and U2374 (N_2374,In_2081,In_488);
nand U2375 (N_2375,In_1579,In_1172);
or U2376 (N_2376,In_1307,In_2467);
and U2377 (N_2377,In_1656,In_658);
or U2378 (N_2378,In_93,In_296);
nand U2379 (N_2379,In_1146,In_2016);
and U2380 (N_2380,In_2331,In_200);
or U2381 (N_2381,In_54,In_78);
nand U2382 (N_2382,In_673,In_595);
and U2383 (N_2383,In_438,In_708);
nor U2384 (N_2384,In_336,In_331);
nand U2385 (N_2385,In_152,In_2016);
nand U2386 (N_2386,In_1619,In_802);
or U2387 (N_2387,In_525,In_1150);
or U2388 (N_2388,In_2112,In_928);
nor U2389 (N_2389,In_1667,In_2156);
or U2390 (N_2390,In_1396,In_736);
and U2391 (N_2391,In_56,In_811);
or U2392 (N_2392,In_244,In_2048);
or U2393 (N_2393,In_1504,In_1060);
or U2394 (N_2394,In_1857,In_553);
and U2395 (N_2395,In_732,In_1529);
or U2396 (N_2396,In_198,In_2146);
and U2397 (N_2397,In_801,In_935);
nor U2398 (N_2398,In_1197,In_1605);
and U2399 (N_2399,In_1992,In_249);
nor U2400 (N_2400,In_1291,In_2283);
nor U2401 (N_2401,In_798,In_2448);
nor U2402 (N_2402,In_52,In_2379);
and U2403 (N_2403,In_2401,In_1869);
and U2404 (N_2404,In_1142,In_2315);
and U2405 (N_2405,In_1279,In_1745);
or U2406 (N_2406,In_958,In_2126);
or U2407 (N_2407,In_172,In_1075);
and U2408 (N_2408,In_2256,In_511);
nor U2409 (N_2409,In_379,In_809);
or U2410 (N_2410,In_387,In_298);
nor U2411 (N_2411,In_683,In_1269);
or U2412 (N_2412,In_2178,In_2016);
nor U2413 (N_2413,In_924,In_2274);
and U2414 (N_2414,In_112,In_172);
and U2415 (N_2415,In_1219,In_427);
nand U2416 (N_2416,In_2305,In_9);
or U2417 (N_2417,In_1468,In_537);
nor U2418 (N_2418,In_319,In_2092);
nor U2419 (N_2419,In_2157,In_31);
or U2420 (N_2420,In_1659,In_1590);
and U2421 (N_2421,In_1072,In_188);
and U2422 (N_2422,In_1408,In_646);
xnor U2423 (N_2423,In_1350,In_1586);
and U2424 (N_2424,In_1242,In_1636);
or U2425 (N_2425,In_2211,In_207);
or U2426 (N_2426,In_1041,In_2292);
nand U2427 (N_2427,In_787,In_626);
nor U2428 (N_2428,In_511,In_1110);
or U2429 (N_2429,In_828,In_1000);
nand U2430 (N_2430,In_1999,In_1667);
nand U2431 (N_2431,In_1162,In_2086);
nor U2432 (N_2432,In_913,In_911);
nand U2433 (N_2433,In_1232,In_1205);
and U2434 (N_2434,In_1803,In_1749);
or U2435 (N_2435,In_1126,In_202);
and U2436 (N_2436,In_1769,In_2417);
nor U2437 (N_2437,In_51,In_1229);
or U2438 (N_2438,In_2011,In_1490);
nor U2439 (N_2439,In_749,In_2043);
nand U2440 (N_2440,In_1196,In_2008);
nor U2441 (N_2441,In_34,In_324);
nand U2442 (N_2442,In_12,In_364);
nand U2443 (N_2443,In_1787,In_2195);
and U2444 (N_2444,In_1204,In_1917);
nand U2445 (N_2445,In_255,In_2190);
nand U2446 (N_2446,In_1306,In_2347);
nand U2447 (N_2447,In_2062,In_2392);
xnor U2448 (N_2448,In_72,In_1006);
nand U2449 (N_2449,In_1761,In_806);
and U2450 (N_2450,In_83,In_175);
nand U2451 (N_2451,In_1259,In_2204);
nor U2452 (N_2452,In_1450,In_993);
nor U2453 (N_2453,In_208,In_1255);
or U2454 (N_2454,In_616,In_974);
nor U2455 (N_2455,In_2385,In_1302);
nand U2456 (N_2456,In_1343,In_1328);
nor U2457 (N_2457,In_437,In_2240);
nand U2458 (N_2458,In_796,In_1995);
nand U2459 (N_2459,In_258,In_576);
nor U2460 (N_2460,In_1927,In_1108);
xnor U2461 (N_2461,In_1384,In_765);
nand U2462 (N_2462,In_1909,In_1132);
or U2463 (N_2463,In_2186,In_1930);
nor U2464 (N_2464,In_1067,In_28);
nand U2465 (N_2465,In_158,In_1457);
nor U2466 (N_2466,In_2091,In_1458);
or U2467 (N_2467,In_803,In_1183);
and U2468 (N_2468,In_561,In_209);
or U2469 (N_2469,In_680,In_1581);
and U2470 (N_2470,In_1674,In_2279);
and U2471 (N_2471,In_1183,In_334);
xnor U2472 (N_2472,In_1318,In_500);
nor U2473 (N_2473,In_942,In_1451);
nor U2474 (N_2474,In_1532,In_1061);
or U2475 (N_2475,In_468,In_87);
nor U2476 (N_2476,In_403,In_850);
or U2477 (N_2477,In_347,In_1282);
xnor U2478 (N_2478,In_851,In_1166);
nand U2479 (N_2479,In_2460,In_1108);
and U2480 (N_2480,In_915,In_1593);
nand U2481 (N_2481,In_768,In_2484);
or U2482 (N_2482,In_456,In_1298);
xor U2483 (N_2483,In_2197,In_1115);
nor U2484 (N_2484,In_1407,In_1044);
nand U2485 (N_2485,In_2260,In_715);
nor U2486 (N_2486,In_856,In_383);
or U2487 (N_2487,In_1207,In_1385);
nand U2488 (N_2488,In_1002,In_2203);
or U2489 (N_2489,In_2482,In_1594);
nand U2490 (N_2490,In_442,In_904);
and U2491 (N_2491,In_615,In_1814);
or U2492 (N_2492,In_150,In_195);
nand U2493 (N_2493,In_373,In_207);
nor U2494 (N_2494,In_70,In_2239);
xor U2495 (N_2495,In_1338,In_824);
and U2496 (N_2496,In_654,In_2467);
and U2497 (N_2497,In_1108,In_154);
or U2498 (N_2498,In_1291,In_1664);
nand U2499 (N_2499,In_1687,In_2200);
or U2500 (N_2500,In_94,In_1834);
nand U2501 (N_2501,In_526,In_299);
or U2502 (N_2502,In_1183,In_1424);
nor U2503 (N_2503,In_1006,In_1727);
or U2504 (N_2504,In_577,In_1779);
or U2505 (N_2505,In_845,In_644);
nand U2506 (N_2506,In_713,In_1400);
or U2507 (N_2507,In_287,In_2319);
or U2508 (N_2508,In_2262,In_1539);
nor U2509 (N_2509,In_1597,In_461);
and U2510 (N_2510,In_2012,In_47);
xnor U2511 (N_2511,In_1012,In_1432);
nand U2512 (N_2512,In_435,In_1955);
nand U2513 (N_2513,In_1512,In_1467);
nor U2514 (N_2514,In_226,In_659);
nand U2515 (N_2515,In_731,In_2345);
nand U2516 (N_2516,In_1967,In_2034);
or U2517 (N_2517,In_222,In_2433);
nand U2518 (N_2518,In_2119,In_2497);
and U2519 (N_2519,In_1246,In_82);
or U2520 (N_2520,In_1957,In_1400);
nand U2521 (N_2521,In_1280,In_371);
nor U2522 (N_2522,In_42,In_1345);
nor U2523 (N_2523,In_1924,In_603);
or U2524 (N_2524,In_57,In_1943);
nor U2525 (N_2525,In_186,In_519);
and U2526 (N_2526,In_2398,In_762);
nand U2527 (N_2527,In_235,In_1306);
or U2528 (N_2528,In_1708,In_817);
nor U2529 (N_2529,In_283,In_2067);
xnor U2530 (N_2530,In_1508,In_1886);
and U2531 (N_2531,In_1172,In_289);
xor U2532 (N_2532,In_1598,In_769);
nor U2533 (N_2533,In_2367,In_733);
nor U2534 (N_2534,In_510,In_351);
and U2535 (N_2535,In_1688,In_2137);
nor U2536 (N_2536,In_1454,In_256);
and U2537 (N_2537,In_867,In_1104);
nor U2538 (N_2538,In_755,In_1138);
and U2539 (N_2539,In_783,In_1296);
and U2540 (N_2540,In_1989,In_965);
and U2541 (N_2541,In_97,In_797);
nor U2542 (N_2542,In_1297,In_222);
xnor U2543 (N_2543,In_1482,In_1079);
nor U2544 (N_2544,In_742,In_2400);
nor U2545 (N_2545,In_1263,In_1891);
and U2546 (N_2546,In_2329,In_1845);
or U2547 (N_2547,In_2056,In_2047);
nor U2548 (N_2548,In_1221,In_333);
and U2549 (N_2549,In_1357,In_2430);
or U2550 (N_2550,In_1736,In_2083);
nor U2551 (N_2551,In_2051,In_1315);
xor U2552 (N_2552,In_882,In_942);
or U2553 (N_2553,In_1381,In_2331);
and U2554 (N_2554,In_607,In_883);
and U2555 (N_2555,In_1550,In_200);
and U2556 (N_2556,In_279,In_151);
nor U2557 (N_2557,In_532,In_348);
or U2558 (N_2558,In_2376,In_2402);
xor U2559 (N_2559,In_1371,In_1907);
and U2560 (N_2560,In_196,In_1515);
xnor U2561 (N_2561,In_2237,In_1175);
xor U2562 (N_2562,In_2486,In_219);
and U2563 (N_2563,In_2136,In_2203);
nor U2564 (N_2564,In_159,In_1432);
nand U2565 (N_2565,In_2085,In_1880);
or U2566 (N_2566,In_1732,In_1178);
nand U2567 (N_2567,In_215,In_2243);
or U2568 (N_2568,In_331,In_2388);
and U2569 (N_2569,In_846,In_1413);
or U2570 (N_2570,In_2338,In_7);
nand U2571 (N_2571,In_2276,In_2421);
nand U2572 (N_2572,In_459,In_538);
and U2573 (N_2573,In_1660,In_558);
or U2574 (N_2574,In_1059,In_1583);
and U2575 (N_2575,In_1090,In_1795);
nor U2576 (N_2576,In_1441,In_2076);
nand U2577 (N_2577,In_1764,In_1044);
and U2578 (N_2578,In_2446,In_280);
nand U2579 (N_2579,In_1592,In_597);
nand U2580 (N_2580,In_1582,In_919);
and U2581 (N_2581,In_713,In_1983);
or U2582 (N_2582,In_1052,In_1092);
xnor U2583 (N_2583,In_1981,In_2225);
or U2584 (N_2584,In_1511,In_1781);
nor U2585 (N_2585,In_436,In_1116);
or U2586 (N_2586,In_489,In_2326);
nand U2587 (N_2587,In_418,In_504);
nor U2588 (N_2588,In_762,In_737);
or U2589 (N_2589,In_172,In_1924);
or U2590 (N_2590,In_974,In_1003);
and U2591 (N_2591,In_1093,In_1046);
and U2592 (N_2592,In_1198,In_1995);
nor U2593 (N_2593,In_2369,In_351);
nor U2594 (N_2594,In_509,In_1201);
and U2595 (N_2595,In_2244,In_959);
nand U2596 (N_2596,In_2083,In_1418);
nor U2597 (N_2597,In_2344,In_1999);
nor U2598 (N_2598,In_836,In_1084);
or U2599 (N_2599,In_1327,In_1722);
xor U2600 (N_2600,In_490,In_1695);
nand U2601 (N_2601,In_1279,In_1636);
and U2602 (N_2602,In_22,In_2207);
or U2603 (N_2603,In_1633,In_115);
and U2604 (N_2604,In_1718,In_2452);
nor U2605 (N_2605,In_1126,In_117);
nor U2606 (N_2606,In_110,In_545);
and U2607 (N_2607,In_880,In_1974);
xnor U2608 (N_2608,In_203,In_2026);
nor U2609 (N_2609,In_2177,In_2381);
xnor U2610 (N_2610,In_157,In_2158);
nor U2611 (N_2611,In_1392,In_583);
nand U2612 (N_2612,In_814,In_1362);
nor U2613 (N_2613,In_566,In_1055);
nor U2614 (N_2614,In_710,In_2420);
nor U2615 (N_2615,In_1353,In_1599);
nand U2616 (N_2616,In_1518,In_1685);
nand U2617 (N_2617,In_2238,In_1157);
nand U2618 (N_2618,In_760,In_2215);
nand U2619 (N_2619,In_369,In_972);
or U2620 (N_2620,In_2166,In_546);
xnor U2621 (N_2621,In_1189,In_2364);
and U2622 (N_2622,In_651,In_2137);
xnor U2623 (N_2623,In_2414,In_1928);
nor U2624 (N_2624,In_543,In_2394);
and U2625 (N_2625,In_2144,In_1130);
or U2626 (N_2626,In_1129,In_696);
or U2627 (N_2627,In_1251,In_2126);
and U2628 (N_2628,In_336,In_28);
nand U2629 (N_2629,In_1783,In_329);
nand U2630 (N_2630,In_642,In_1370);
and U2631 (N_2631,In_906,In_615);
and U2632 (N_2632,In_170,In_2432);
nand U2633 (N_2633,In_1985,In_271);
and U2634 (N_2634,In_2074,In_487);
nor U2635 (N_2635,In_1683,In_2451);
nor U2636 (N_2636,In_1594,In_1237);
and U2637 (N_2637,In_855,In_305);
nor U2638 (N_2638,In_1819,In_616);
and U2639 (N_2639,In_620,In_242);
xor U2640 (N_2640,In_511,In_126);
or U2641 (N_2641,In_1273,In_520);
nand U2642 (N_2642,In_2112,In_1039);
or U2643 (N_2643,In_255,In_157);
nand U2644 (N_2644,In_610,In_1893);
or U2645 (N_2645,In_2482,In_1542);
nor U2646 (N_2646,In_2070,In_927);
nand U2647 (N_2647,In_1419,In_1686);
nand U2648 (N_2648,In_26,In_2359);
nor U2649 (N_2649,In_1107,In_93);
or U2650 (N_2650,In_833,In_48);
or U2651 (N_2651,In_1853,In_1279);
and U2652 (N_2652,In_1405,In_489);
and U2653 (N_2653,In_631,In_1090);
nor U2654 (N_2654,In_2419,In_934);
and U2655 (N_2655,In_2038,In_958);
and U2656 (N_2656,In_1505,In_316);
nand U2657 (N_2657,In_1768,In_1990);
nor U2658 (N_2658,In_873,In_2333);
and U2659 (N_2659,In_1683,In_2420);
nor U2660 (N_2660,In_2225,In_2435);
nand U2661 (N_2661,In_841,In_529);
and U2662 (N_2662,In_1998,In_353);
nor U2663 (N_2663,In_346,In_2227);
nor U2664 (N_2664,In_1488,In_2099);
nand U2665 (N_2665,In_942,In_1850);
nand U2666 (N_2666,In_2332,In_1300);
and U2667 (N_2667,In_1847,In_468);
nand U2668 (N_2668,In_317,In_1844);
nor U2669 (N_2669,In_313,In_2264);
or U2670 (N_2670,In_1507,In_1562);
nand U2671 (N_2671,In_763,In_1705);
and U2672 (N_2672,In_1898,In_1435);
xnor U2673 (N_2673,In_534,In_2279);
nand U2674 (N_2674,In_1629,In_406);
nor U2675 (N_2675,In_2499,In_865);
or U2676 (N_2676,In_451,In_335);
nand U2677 (N_2677,In_1681,In_2218);
and U2678 (N_2678,In_662,In_886);
or U2679 (N_2679,In_1784,In_821);
nor U2680 (N_2680,In_2134,In_418);
nor U2681 (N_2681,In_596,In_2358);
or U2682 (N_2682,In_2495,In_552);
nor U2683 (N_2683,In_2210,In_1946);
nand U2684 (N_2684,In_324,In_2161);
or U2685 (N_2685,In_155,In_167);
nor U2686 (N_2686,In_1360,In_1780);
nor U2687 (N_2687,In_1726,In_976);
nor U2688 (N_2688,In_1765,In_14);
nand U2689 (N_2689,In_337,In_1853);
and U2690 (N_2690,In_1322,In_137);
xnor U2691 (N_2691,In_1959,In_1386);
and U2692 (N_2692,In_1855,In_141);
and U2693 (N_2693,In_2074,In_995);
nand U2694 (N_2694,In_30,In_1006);
and U2695 (N_2695,In_976,In_1070);
or U2696 (N_2696,In_195,In_1962);
or U2697 (N_2697,In_2341,In_1762);
nor U2698 (N_2698,In_565,In_2471);
and U2699 (N_2699,In_110,In_1101);
and U2700 (N_2700,In_2370,In_473);
or U2701 (N_2701,In_1870,In_935);
nand U2702 (N_2702,In_1278,In_1418);
and U2703 (N_2703,In_1317,In_670);
or U2704 (N_2704,In_1648,In_193);
or U2705 (N_2705,In_237,In_2207);
or U2706 (N_2706,In_1098,In_2112);
nand U2707 (N_2707,In_1138,In_790);
nand U2708 (N_2708,In_634,In_931);
nand U2709 (N_2709,In_1156,In_2384);
xor U2710 (N_2710,In_872,In_146);
nor U2711 (N_2711,In_2080,In_1720);
nor U2712 (N_2712,In_433,In_1996);
nand U2713 (N_2713,In_1133,In_2449);
and U2714 (N_2714,In_1508,In_1072);
and U2715 (N_2715,In_189,In_1215);
nor U2716 (N_2716,In_1860,In_1099);
and U2717 (N_2717,In_541,In_1709);
and U2718 (N_2718,In_1472,In_2013);
and U2719 (N_2719,In_1644,In_2118);
nor U2720 (N_2720,In_399,In_1661);
or U2721 (N_2721,In_722,In_1538);
nor U2722 (N_2722,In_406,In_803);
nand U2723 (N_2723,In_1530,In_100);
or U2724 (N_2724,In_1644,In_1722);
nor U2725 (N_2725,In_1406,In_1787);
xor U2726 (N_2726,In_1465,In_512);
nor U2727 (N_2727,In_96,In_1235);
nand U2728 (N_2728,In_185,In_2065);
or U2729 (N_2729,In_2396,In_1342);
nor U2730 (N_2730,In_2225,In_50);
nor U2731 (N_2731,In_1080,In_2183);
nand U2732 (N_2732,In_885,In_99);
nand U2733 (N_2733,In_1111,In_1116);
nor U2734 (N_2734,In_2456,In_405);
or U2735 (N_2735,In_1717,In_1819);
nand U2736 (N_2736,In_1719,In_757);
xnor U2737 (N_2737,In_550,In_1837);
nand U2738 (N_2738,In_1049,In_991);
and U2739 (N_2739,In_472,In_192);
nand U2740 (N_2740,In_348,In_553);
nand U2741 (N_2741,In_864,In_1773);
or U2742 (N_2742,In_1109,In_828);
xor U2743 (N_2743,In_2111,In_246);
or U2744 (N_2744,In_1614,In_2252);
nand U2745 (N_2745,In_2211,In_789);
nand U2746 (N_2746,In_1311,In_1877);
or U2747 (N_2747,In_1587,In_589);
and U2748 (N_2748,In_2457,In_20);
or U2749 (N_2749,In_587,In_649);
nand U2750 (N_2750,In_975,In_1698);
and U2751 (N_2751,In_563,In_1030);
and U2752 (N_2752,In_695,In_1931);
nand U2753 (N_2753,In_364,In_1683);
nor U2754 (N_2754,In_474,In_1162);
xnor U2755 (N_2755,In_2173,In_601);
or U2756 (N_2756,In_2396,In_1053);
nor U2757 (N_2757,In_437,In_1732);
xor U2758 (N_2758,In_169,In_1238);
nor U2759 (N_2759,In_1394,In_1698);
nor U2760 (N_2760,In_1417,In_2214);
nor U2761 (N_2761,In_1480,In_299);
xor U2762 (N_2762,In_2156,In_1669);
and U2763 (N_2763,In_1372,In_2116);
and U2764 (N_2764,In_424,In_880);
nand U2765 (N_2765,In_292,In_1844);
nand U2766 (N_2766,In_442,In_1717);
nand U2767 (N_2767,In_739,In_1279);
or U2768 (N_2768,In_1636,In_2204);
or U2769 (N_2769,In_191,In_2499);
xnor U2770 (N_2770,In_1793,In_2472);
nand U2771 (N_2771,In_68,In_1504);
nor U2772 (N_2772,In_2091,In_735);
and U2773 (N_2773,In_182,In_280);
nand U2774 (N_2774,In_914,In_1611);
xnor U2775 (N_2775,In_2108,In_1022);
nand U2776 (N_2776,In_1796,In_1398);
nor U2777 (N_2777,In_775,In_1964);
xor U2778 (N_2778,In_1189,In_2352);
xor U2779 (N_2779,In_1393,In_1589);
nand U2780 (N_2780,In_1757,In_2238);
or U2781 (N_2781,In_336,In_2472);
xor U2782 (N_2782,In_47,In_1768);
nor U2783 (N_2783,In_1461,In_955);
nor U2784 (N_2784,In_198,In_546);
xor U2785 (N_2785,In_1123,In_1332);
nor U2786 (N_2786,In_168,In_1861);
nor U2787 (N_2787,In_2390,In_509);
nor U2788 (N_2788,In_1521,In_325);
or U2789 (N_2789,In_1425,In_1852);
nor U2790 (N_2790,In_30,In_1028);
or U2791 (N_2791,In_1697,In_2448);
nand U2792 (N_2792,In_118,In_729);
xor U2793 (N_2793,In_1455,In_1785);
or U2794 (N_2794,In_1593,In_2124);
and U2795 (N_2795,In_343,In_1150);
or U2796 (N_2796,In_1853,In_1650);
and U2797 (N_2797,In_1126,In_790);
xnor U2798 (N_2798,In_246,In_354);
and U2799 (N_2799,In_934,In_297);
nor U2800 (N_2800,In_1578,In_486);
and U2801 (N_2801,In_1197,In_525);
nand U2802 (N_2802,In_277,In_1609);
xnor U2803 (N_2803,In_300,In_391);
nand U2804 (N_2804,In_1444,In_2452);
nand U2805 (N_2805,In_978,In_194);
nor U2806 (N_2806,In_341,In_1872);
and U2807 (N_2807,In_506,In_1933);
xor U2808 (N_2808,In_1737,In_555);
xor U2809 (N_2809,In_2012,In_424);
or U2810 (N_2810,In_2114,In_300);
or U2811 (N_2811,In_1681,In_306);
and U2812 (N_2812,In_2046,In_1683);
nand U2813 (N_2813,In_1082,In_631);
nor U2814 (N_2814,In_269,In_1976);
nand U2815 (N_2815,In_710,In_2445);
and U2816 (N_2816,In_1554,In_325);
nand U2817 (N_2817,In_572,In_1508);
and U2818 (N_2818,In_1008,In_1001);
or U2819 (N_2819,In_1872,In_1030);
nor U2820 (N_2820,In_1970,In_2091);
nand U2821 (N_2821,In_2435,In_1678);
nand U2822 (N_2822,In_1566,In_415);
and U2823 (N_2823,In_1127,In_2442);
or U2824 (N_2824,In_697,In_468);
nand U2825 (N_2825,In_2222,In_2483);
or U2826 (N_2826,In_1425,In_2066);
and U2827 (N_2827,In_645,In_1673);
and U2828 (N_2828,In_2279,In_2499);
or U2829 (N_2829,In_1556,In_2321);
nor U2830 (N_2830,In_1101,In_2168);
and U2831 (N_2831,In_543,In_1972);
nand U2832 (N_2832,In_829,In_2196);
and U2833 (N_2833,In_1851,In_2234);
nor U2834 (N_2834,In_793,In_2425);
nand U2835 (N_2835,In_1018,In_955);
or U2836 (N_2836,In_725,In_1798);
xnor U2837 (N_2837,In_867,In_1739);
or U2838 (N_2838,In_707,In_2455);
nand U2839 (N_2839,In_1391,In_568);
xnor U2840 (N_2840,In_1220,In_971);
nor U2841 (N_2841,In_229,In_1618);
and U2842 (N_2842,In_1140,In_1878);
nand U2843 (N_2843,In_797,In_625);
or U2844 (N_2844,In_2484,In_762);
or U2845 (N_2845,In_330,In_190);
nor U2846 (N_2846,In_449,In_753);
nor U2847 (N_2847,In_637,In_1096);
and U2848 (N_2848,In_1647,In_1909);
and U2849 (N_2849,In_779,In_11);
nand U2850 (N_2850,In_793,In_1030);
nand U2851 (N_2851,In_1025,In_1086);
or U2852 (N_2852,In_1234,In_782);
xnor U2853 (N_2853,In_1612,In_387);
or U2854 (N_2854,In_457,In_78);
nand U2855 (N_2855,In_2017,In_1711);
or U2856 (N_2856,In_95,In_473);
nand U2857 (N_2857,In_1717,In_83);
or U2858 (N_2858,In_413,In_1683);
nand U2859 (N_2859,In_2094,In_1646);
nor U2860 (N_2860,In_2031,In_339);
or U2861 (N_2861,In_716,In_938);
or U2862 (N_2862,In_1338,In_2004);
nor U2863 (N_2863,In_1489,In_1957);
nor U2864 (N_2864,In_2397,In_2488);
nor U2865 (N_2865,In_1775,In_598);
nand U2866 (N_2866,In_572,In_1498);
nand U2867 (N_2867,In_2442,In_755);
nand U2868 (N_2868,In_1867,In_1492);
nand U2869 (N_2869,In_1002,In_906);
and U2870 (N_2870,In_1256,In_2340);
and U2871 (N_2871,In_490,In_1291);
nor U2872 (N_2872,In_1262,In_280);
nand U2873 (N_2873,In_753,In_704);
nand U2874 (N_2874,In_2437,In_1416);
or U2875 (N_2875,In_390,In_519);
or U2876 (N_2876,In_1874,In_1794);
and U2877 (N_2877,In_451,In_1144);
and U2878 (N_2878,In_2140,In_1565);
or U2879 (N_2879,In_2140,In_418);
nand U2880 (N_2880,In_1992,In_450);
nand U2881 (N_2881,In_884,In_1477);
nand U2882 (N_2882,In_1942,In_464);
and U2883 (N_2883,In_103,In_767);
nor U2884 (N_2884,In_1533,In_1193);
xor U2885 (N_2885,In_1452,In_1015);
nor U2886 (N_2886,In_1648,In_1614);
nand U2887 (N_2887,In_321,In_2042);
and U2888 (N_2888,In_1248,In_433);
nor U2889 (N_2889,In_180,In_2253);
nand U2890 (N_2890,In_869,In_2077);
nand U2891 (N_2891,In_1120,In_652);
and U2892 (N_2892,In_1867,In_747);
xnor U2893 (N_2893,In_1604,In_1228);
and U2894 (N_2894,In_376,In_1744);
or U2895 (N_2895,In_970,In_992);
and U2896 (N_2896,In_1254,In_405);
or U2897 (N_2897,In_2323,In_457);
xnor U2898 (N_2898,In_2227,In_13);
and U2899 (N_2899,In_241,In_1974);
nand U2900 (N_2900,In_754,In_16);
or U2901 (N_2901,In_1154,In_940);
or U2902 (N_2902,In_1207,In_1433);
xnor U2903 (N_2903,In_2458,In_25);
nor U2904 (N_2904,In_1116,In_330);
or U2905 (N_2905,In_2004,In_1817);
nand U2906 (N_2906,In_1635,In_748);
xor U2907 (N_2907,In_125,In_65);
and U2908 (N_2908,In_1820,In_1657);
nor U2909 (N_2909,In_564,In_1720);
nor U2910 (N_2910,In_1057,In_1861);
or U2911 (N_2911,In_1829,In_773);
nand U2912 (N_2912,In_1186,In_2127);
nor U2913 (N_2913,In_1067,In_1989);
nor U2914 (N_2914,In_1738,In_343);
nor U2915 (N_2915,In_867,In_774);
and U2916 (N_2916,In_760,In_586);
and U2917 (N_2917,In_236,In_487);
xor U2918 (N_2918,In_115,In_2490);
xnor U2919 (N_2919,In_1545,In_2198);
xor U2920 (N_2920,In_1604,In_551);
or U2921 (N_2921,In_859,In_1724);
nor U2922 (N_2922,In_702,In_1412);
xor U2923 (N_2923,In_845,In_84);
nand U2924 (N_2924,In_2430,In_992);
nor U2925 (N_2925,In_1606,In_332);
and U2926 (N_2926,In_1283,In_2214);
nand U2927 (N_2927,In_2217,In_326);
nor U2928 (N_2928,In_2048,In_2025);
and U2929 (N_2929,In_476,In_2328);
nor U2930 (N_2930,In_1746,In_2030);
nor U2931 (N_2931,In_1168,In_785);
xor U2932 (N_2932,In_804,In_1024);
nor U2933 (N_2933,In_1331,In_695);
nand U2934 (N_2934,In_2458,In_2344);
and U2935 (N_2935,In_364,In_217);
xor U2936 (N_2936,In_2453,In_61);
xnor U2937 (N_2937,In_99,In_2394);
and U2938 (N_2938,In_1057,In_1664);
or U2939 (N_2939,In_2072,In_449);
and U2940 (N_2940,In_2304,In_1773);
nand U2941 (N_2941,In_2316,In_130);
or U2942 (N_2942,In_733,In_1487);
and U2943 (N_2943,In_266,In_2033);
or U2944 (N_2944,In_890,In_1934);
or U2945 (N_2945,In_2048,In_2155);
nor U2946 (N_2946,In_116,In_1076);
nor U2947 (N_2947,In_1977,In_2391);
or U2948 (N_2948,In_1258,In_2496);
or U2949 (N_2949,In_1002,In_286);
or U2950 (N_2950,In_794,In_789);
or U2951 (N_2951,In_2089,In_53);
and U2952 (N_2952,In_2102,In_2466);
nor U2953 (N_2953,In_1335,In_2127);
and U2954 (N_2954,In_710,In_2183);
nor U2955 (N_2955,In_1767,In_2328);
and U2956 (N_2956,In_146,In_1079);
or U2957 (N_2957,In_1832,In_1990);
and U2958 (N_2958,In_2204,In_1893);
or U2959 (N_2959,In_827,In_279);
nand U2960 (N_2960,In_1921,In_876);
nand U2961 (N_2961,In_2441,In_616);
and U2962 (N_2962,In_594,In_83);
nor U2963 (N_2963,In_1797,In_832);
and U2964 (N_2964,In_1965,In_752);
and U2965 (N_2965,In_1691,In_1865);
and U2966 (N_2966,In_1287,In_2376);
and U2967 (N_2967,In_1275,In_1486);
and U2968 (N_2968,In_2215,In_303);
nor U2969 (N_2969,In_1858,In_2494);
xor U2970 (N_2970,In_1322,In_1308);
nand U2971 (N_2971,In_287,In_1146);
or U2972 (N_2972,In_308,In_301);
nand U2973 (N_2973,In_2012,In_1048);
and U2974 (N_2974,In_748,In_1736);
or U2975 (N_2975,In_644,In_353);
xnor U2976 (N_2976,In_709,In_1504);
and U2977 (N_2977,In_912,In_1212);
nand U2978 (N_2978,In_270,In_287);
xnor U2979 (N_2979,In_1655,In_2227);
nor U2980 (N_2980,In_626,In_335);
nor U2981 (N_2981,In_906,In_1168);
and U2982 (N_2982,In_833,In_908);
and U2983 (N_2983,In_1738,In_320);
and U2984 (N_2984,In_935,In_2103);
or U2985 (N_2985,In_1856,In_1733);
and U2986 (N_2986,In_1663,In_2361);
nor U2987 (N_2987,In_2498,In_2373);
nand U2988 (N_2988,In_232,In_445);
or U2989 (N_2989,In_2165,In_2235);
or U2990 (N_2990,In_730,In_190);
or U2991 (N_2991,In_1923,In_2276);
and U2992 (N_2992,In_1527,In_1244);
xor U2993 (N_2993,In_1217,In_77);
nand U2994 (N_2994,In_873,In_679);
or U2995 (N_2995,In_2269,In_2341);
nor U2996 (N_2996,In_546,In_2096);
and U2997 (N_2997,In_1033,In_2088);
and U2998 (N_2998,In_867,In_62);
or U2999 (N_2999,In_83,In_2231);
nor U3000 (N_3000,In_500,In_1644);
xnor U3001 (N_3001,In_1938,In_1432);
nor U3002 (N_3002,In_2138,In_1635);
nor U3003 (N_3003,In_1354,In_1728);
and U3004 (N_3004,In_570,In_1491);
nor U3005 (N_3005,In_1054,In_488);
or U3006 (N_3006,In_2125,In_271);
or U3007 (N_3007,In_1732,In_1575);
or U3008 (N_3008,In_1186,In_1992);
or U3009 (N_3009,In_620,In_1392);
nand U3010 (N_3010,In_867,In_1532);
nor U3011 (N_3011,In_1777,In_920);
nand U3012 (N_3012,In_2355,In_2075);
and U3013 (N_3013,In_1239,In_690);
nand U3014 (N_3014,In_641,In_405);
nand U3015 (N_3015,In_409,In_225);
nand U3016 (N_3016,In_1273,In_132);
nand U3017 (N_3017,In_2047,In_388);
nor U3018 (N_3018,In_663,In_1996);
nand U3019 (N_3019,In_281,In_1644);
and U3020 (N_3020,In_811,In_1219);
nand U3021 (N_3021,In_2169,In_2198);
nor U3022 (N_3022,In_1462,In_1017);
and U3023 (N_3023,In_992,In_687);
nand U3024 (N_3024,In_807,In_681);
nor U3025 (N_3025,In_2436,In_2084);
nor U3026 (N_3026,In_267,In_2185);
or U3027 (N_3027,In_212,In_929);
or U3028 (N_3028,In_377,In_935);
nor U3029 (N_3029,In_1822,In_1064);
or U3030 (N_3030,In_1118,In_496);
xnor U3031 (N_3031,In_371,In_541);
or U3032 (N_3032,In_1297,In_636);
and U3033 (N_3033,In_1107,In_1707);
nand U3034 (N_3034,In_444,In_6);
or U3035 (N_3035,In_1141,In_75);
nor U3036 (N_3036,In_116,In_1877);
and U3037 (N_3037,In_1378,In_2112);
nor U3038 (N_3038,In_1144,In_5);
xor U3039 (N_3039,In_2453,In_2105);
nand U3040 (N_3040,In_2414,In_220);
and U3041 (N_3041,In_53,In_898);
nor U3042 (N_3042,In_821,In_1017);
xnor U3043 (N_3043,In_2195,In_1036);
or U3044 (N_3044,In_994,In_1245);
and U3045 (N_3045,In_1808,In_1867);
and U3046 (N_3046,In_1943,In_1673);
nor U3047 (N_3047,In_460,In_119);
nand U3048 (N_3048,In_1422,In_830);
nand U3049 (N_3049,In_2336,In_1940);
and U3050 (N_3050,In_539,In_829);
nand U3051 (N_3051,In_1560,In_14);
nand U3052 (N_3052,In_2042,In_2122);
nor U3053 (N_3053,In_2074,In_2413);
nand U3054 (N_3054,In_1692,In_2116);
nand U3055 (N_3055,In_2289,In_1986);
or U3056 (N_3056,In_1961,In_120);
nand U3057 (N_3057,In_1323,In_1230);
nor U3058 (N_3058,In_999,In_2192);
xor U3059 (N_3059,In_945,In_2087);
or U3060 (N_3060,In_272,In_1133);
xnor U3061 (N_3061,In_304,In_354);
xnor U3062 (N_3062,In_2320,In_1466);
nand U3063 (N_3063,In_2285,In_2278);
and U3064 (N_3064,In_2010,In_519);
or U3065 (N_3065,In_335,In_1344);
xnor U3066 (N_3066,In_237,In_1646);
and U3067 (N_3067,In_2326,In_1831);
and U3068 (N_3068,In_1134,In_1718);
nor U3069 (N_3069,In_611,In_1446);
and U3070 (N_3070,In_415,In_1395);
xor U3071 (N_3071,In_1593,In_662);
and U3072 (N_3072,In_257,In_1052);
nand U3073 (N_3073,In_2360,In_2143);
or U3074 (N_3074,In_2289,In_654);
or U3075 (N_3075,In_689,In_209);
and U3076 (N_3076,In_1934,In_931);
nand U3077 (N_3077,In_2006,In_2226);
nand U3078 (N_3078,In_2450,In_1371);
nand U3079 (N_3079,In_233,In_2383);
nor U3080 (N_3080,In_168,In_629);
nor U3081 (N_3081,In_1998,In_1352);
and U3082 (N_3082,In_1303,In_1344);
nand U3083 (N_3083,In_2210,In_763);
nand U3084 (N_3084,In_291,In_292);
xor U3085 (N_3085,In_2266,In_2065);
and U3086 (N_3086,In_1757,In_1774);
nand U3087 (N_3087,In_1763,In_2216);
nor U3088 (N_3088,In_1544,In_1805);
nor U3089 (N_3089,In_1437,In_1332);
nor U3090 (N_3090,In_2269,In_463);
xor U3091 (N_3091,In_601,In_1998);
nor U3092 (N_3092,In_1919,In_2317);
or U3093 (N_3093,In_1655,In_1473);
nor U3094 (N_3094,In_374,In_967);
or U3095 (N_3095,In_2051,In_190);
nor U3096 (N_3096,In_985,In_1626);
and U3097 (N_3097,In_365,In_2318);
or U3098 (N_3098,In_1922,In_2367);
nor U3099 (N_3099,In_530,In_1779);
nor U3100 (N_3100,In_1734,In_901);
nand U3101 (N_3101,In_169,In_2087);
xor U3102 (N_3102,In_1678,In_661);
nand U3103 (N_3103,In_2325,In_1445);
or U3104 (N_3104,In_1950,In_203);
or U3105 (N_3105,In_331,In_772);
nand U3106 (N_3106,In_2492,In_37);
nor U3107 (N_3107,In_2075,In_251);
nand U3108 (N_3108,In_407,In_1137);
nand U3109 (N_3109,In_623,In_2305);
or U3110 (N_3110,In_1056,In_538);
xnor U3111 (N_3111,In_2000,In_2063);
nand U3112 (N_3112,In_387,In_1379);
and U3113 (N_3113,In_1138,In_1966);
xor U3114 (N_3114,In_892,In_579);
and U3115 (N_3115,In_790,In_501);
and U3116 (N_3116,In_303,In_1009);
and U3117 (N_3117,In_44,In_312);
and U3118 (N_3118,In_1203,In_552);
or U3119 (N_3119,In_59,In_622);
nand U3120 (N_3120,In_856,In_816);
and U3121 (N_3121,In_1131,In_1673);
nand U3122 (N_3122,In_803,In_1558);
xnor U3123 (N_3123,In_740,In_263);
nor U3124 (N_3124,In_1,In_2032);
and U3125 (N_3125,In_2090,In_1394);
nor U3126 (N_3126,In_1090,In_1768);
and U3127 (N_3127,In_1736,In_1266);
nor U3128 (N_3128,In_2228,In_1016);
nand U3129 (N_3129,In_2484,In_1522);
xnor U3130 (N_3130,In_2364,In_1401);
nor U3131 (N_3131,In_1637,In_742);
nand U3132 (N_3132,In_1050,In_56);
or U3133 (N_3133,In_1118,In_2187);
xnor U3134 (N_3134,In_1350,In_829);
or U3135 (N_3135,In_1458,In_1575);
or U3136 (N_3136,In_2033,In_1729);
nand U3137 (N_3137,In_642,In_2304);
nand U3138 (N_3138,In_1090,In_1502);
nor U3139 (N_3139,In_1055,In_1889);
nor U3140 (N_3140,In_1241,In_2004);
nor U3141 (N_3141,In_814,In_1175);
nor U3142 (N_3142,In_1042,In_2343);
nand U3143 (N_3143,In_2230,In_213);
nand U3144 (N_3144,In_951,In_1812);
nand U3145 (N_3145,In_1077,In_647);
nand U3146 (N_3146,In_1010,In_199);
or U3147 (N_3147,In_2130,In_482);
nor U3148 (N_3148,In_2288,In_1671);
nor U3149 (N_3149,In_534,In_2364);
and U3150 (N_3150,In_2073,In_323);
nor U3151 (N_3151,In_2497,In_1316);
or U3152 (N_3152,In_1510,In_1752);
nand U3153 (N_3153,In_1940,In_1981);
or U3154 (N_3154,In_456,In_1617);
nand U3155 (N_3155,In_42,In_1492);
nand U3156 (N_3156,In_126,In_746);
or U3157 (N_3157,In_2313,In_1439);
or U3158 (N_3158,In_1983,In_53);
nand U3159 (N_3159,In_1602,In_127);
nor U3160 (N_3160,In_49,In_689);
nor U3161 (N_3161,In_500,In_2131);
nand U3162 (N_3162,In_853,In_1347);
nor U3163 (N_3163,In_1707,In_2240);
nand U3164 (N_3164,In_950,In_1376);
and U3165 (N_3165,In_1858,In_2209);
nor U3166 (N_3166,In_2361,In_1875);
or U3167 (N_3167,In_1312,In_64);
and U3168 (N_3168,In_764,In_1962);
nor U3169 (N_3169,In_896,In_489);
and U3170 (N_3170,In_1559,In_2367);
and U3171 (N_3171,In_988,In_306);
nor U3172 (N_3172,In_2192,In_458);
nor U3173 (N_3173,In_1405,In_916);
nor U3174 (N_3174,In_276,In_2132);
nand U3175 (N_3175,In_305,In_1412);
xnor U3176 (N_3176,In_2094,In_1706);
and U3177 (N_3177,In_1201,In_346);
xnor U3178 (N_3178,In_1270,In_109);
and U3179 (N_3179,In_998,In_1681);
nor U3180 (N_3180,In_1386,In_98);
xor U3181 (N_3181,In_1357,In_754);
and U3182 (N_3182,In_1772,In_2037);
or U3183 (N_3183,In_1040,In_1191);
or U3184 (N_3184,In_2286,In_221);
or U3185 (N_3185,In_2176,In_111);
nand U3186 (N_3186,In_331,In_1721);
nand U3187 (N_3187,In_315,In_935);
or U3188 (N_3188,In_1987,In_444);
nand U3189 (N_3189,In_370,In_774);
or U3190 (N_3190,In_205,In_2481);
or U3191 (N_3191,In_1585,In_752);
nand U3192 (N_3192,In_987,In_2325);
and U3193 (N_3193,In_605,In_692);
nor U3194 (N_3194,In_1087,In_713);
and U3195 (N_3195,In_1417,In_1081);
nor U3196 (N_3196,In_1740,In_2322);
or U3197 (N_3197,In_1572,In_1444);
and U3198 (N_3198,In_1672,In_1761);
or U3199 (N_3199,In_2298,In_1832);
and U3200 (N_3200,In_1111,In_1905);
xnor U3201 (N_3201,In_2130,In_55);
nand U3202 (N_3202,In_1250,In_2382);
nor U3203 (N_3203,In_2328,In_1639);
or U3204 (N_3204,In_2058,In_136);
nand U3205 (N_3205,In_2292,In_2355);
xor U3206 (N_3206,In_2188,In_319);
xor U3207 (N_3207,In_419,In_1606);
nor U3208 (N_3208,In_586,In_311);
or U3209 (N_3209,In_1558,In_438);
nand U3210 (N_3210,In_1822,In_883);
or U3211 (N_3211,In_56,In_2392);
and U3212 (N_3212,In_98,In_89);
nor U3213 (N_3213,In_374,In_211);
or U3214 (N_3214,In_1332,In_1312);
and U3215 (N_3215,In_1532,In_2348);
nand U3216 (N_3216,In_1820,In_1708);
or U3217 (N_3217,In_2142,In_1400);
and U3218 (N_3218,In_291,In_2199);
or U3219 (N_3219,In_2438,In_1294);
nand U3220 (N_3220,In_637,In_2185);
or U3221 (N_3221,In_2004,In_1951);
nand U3222 (N_3222,In_381,In_1410);
nand U3223 (N_3223,In_1568,In_244);
and U3224 (N_3224,In_2270,In_226);
nand U3225 (N_3225,In_1133,In_2406);
or U3226 (N_3226,In_439,In_565);
nand U3227 (N_3227,In_1686,In_1220);
nor U3228 (N_3228,In_1902,In_865);
nor U3229 (N_3229,In_1066,In_2026);
or U3230 (N_3230,In_1988,In_2094);
or U3231 (N_3231,In_1925,In_2023);
nand U3232 (N_3232,In_1840,In_1577);
nor U3233 (N_3233,In_120,In_4);
or U3234 (N_3234,In_2246,In_1327);
nor U3235 (N_3235,In_730,In_991);
nor U3236 (N_3236,In_1339,In_202);
or U3237 (N_3237,In_52,In_1867);
or U3238 (N_3238,In_1031,In_1657);
nor U3239 (N_3239,In_1375,In_184);
or U3240 (N_3240,In_318,In_2377);
or U3241 (N_3241,In_1283,In_1042);
xnor U3242 (N_3242,In_2426,In_625);
nand U3243 (N_3243,In_1383,In_576);
xnor U3244 (N_3244,In_1309,In_62);
xnor U3245 (N_3245,In_1932,In_214);
nand U3246 (N_3246,In_1642,In_924);
and U3247 (N_3247,In_188,In_333);
nand U3248 (N_3248,In_187,In_805);
nor U3249 (N_3249,In_2301,In_1444);
nor U3250 (N_3250,In_1710,In_1909);
nor U3251 (N_3251,In_678,In_373);
or U3252 (N_3252,In_2261,In_372);
nand U3253 (N_3253,In_134,In_1509);
nor U3254 (N_3254,In_2495,In_1576);
or U3255 (N_3255,In_1896,In_846);
nand U3256 (N_3256,In_1265,In_242);
nor U3257 (N_3257,In_1176,In_675);
nand U3258 (N_3258,In_1793,In_454);
nand U3259 (N_3259,In_165,In_1638);
nand U3260 (N_3260,In_1659,In_26);
nand U3261 (N_3261,In_1103,In_2069);
nor U3262 (N_3262,In_1757,In_460);
and U3263 (N_3263,In_1413,In_2189);
and U3264 (N_3264,In_1656,In_1081);
or U3265 (N_3265,In_1905,In_904);
nor U3266 (N_3266,In_1339,In_836);
and U3267 (N_3267,In_430,In_1327);
or U3268 (N_3268,In_631,In_430);
nand U3269 (N_3269,In_1017,In_123);
nand U3270 (N_3270,In_2424,In_2020);
nor U3271 (N_3271,In_124,In_126);
or U3272 (N_3272,In_674,In_2226);
or U3273 (N_3273,In_751,In_548);
xor U3274 (N_3274,In_1404,In_1872);
nand U3275 (N_3275,In_2051,In_2053);
or U3276 (N_3276,In_1312,In_2163);
and U3277 (N_3277,In_748,In_2061);
nand U3278 (N_3278,In_1753,In_454);
and U3279 (N_3279,In_1878,In_119);
or U3280 (N_3280,In_1252,In_2155);
xor U3281 (N_3281,In_2266,In_293);
nor U3282 (N_3282,In_859,In_1548);
nor U3283 (N_3283,In_193,In_241);
nor U3284 (N_3284,In_88,In_139);
xor U3285 (N_3285,In_1468,In_2151);
nor U3286 (N_3286,In_374,In_538);
xor U3287 (N_3287,In_1992,In_2492);
and U3288 (N_3288,In_2031,In_1619);
xor U3289 (N_3289,In_132,In_468);
and U3290 (N_3290,In_2101,In_2008);
nor U3291 (N_3291,In_793,In_1116);
or U3292 (N_3292,In_1863,In_2063);
and U3293 (N_3293,In_1390,In_1408);
and U3294 (N_3294,In_2494,In_1836);
and U3295 (N_3295,In_1671,In_1245);
or U3296 (N_3296,In_1142,In_203);
or U3297 (N_3297,In_653,In_1703);
nand U3298 (N_3298,In_246,In_1874);
nor U3299 (N_3299,In_2289,In_2114);
or U3300 (N_3300,In_1486,In_1264);
or U3301 (N_3301,In_676,In_194);
nand U3302 (N_3302,In_2469,In_1344);
nand U3303 (N_3303,In_1586,In_2032);
or U3304 (N_3304,In_1706,In_427);
nor U3305 (N_3305,In_2342,In_257);
nand U3306 (N_3306,In_591,In_2337);
nand U3307 (N_3307,In_1500,In_2361);
nor U3308 (N_3308,In_101,In_597);
nand U3309 (N_3309,In_2031,In_765);
nand U3310 (N_3310,In_1644,In_1273);
or U3311 (N_3311,In_426,In_200);
nor U3312 (N_3312,In_1791,In_2392);
and U3313 (N_3313,In_1057,In_2137);
nand U3314 (N_3314,In_2043,In_1553);
nand U3315 (N_3315,In_568,In_1369);
xnor U3316 (N_3316,In_588,In_670);
nand U3317 (N_3317,In_1015,In_1788);
nand U3318 (N_3318,In_1028,In_155);
and U3319 (N_3319,In_2430,In_1046);
nand U3320 (N_3320,In_1998,In_1345);
and U3321 (N_3321,In_1372,In_981);
nand U3322 (N_3322,In_1986,In_1229);
nor U3323 (N_3323,In_213,In_1832);
xor U3324 (N_3324,In_511,In_2079);
nand U3325 (N_3325,In_208,In_2029);
and U3326 (N_3326,In_54,In_1901);
nor U3327 (N_3327,In_1031,In_339);
and U3328 (N_3328,In_1030,In_807);
or U3329 (N_3329,In_1261,In_2010);
or U3330 (N_3330,In_1814,In_2225);
xor U3331 (N_3331,In_1380,In_823);
nor U3332 (N_3332,In_2216,In_681);
nand U3333 (N_3333,In_1946,In_393);
nand U3334 (N_3334,In_1333,In_478);
nand U3335 (N_3335,In_1720,In_1337);
or U3336 (N_3336,In_1080,In_1037);
xor U3337 (N_3337,In_442,In_308);
nor U3338 (N_3338,In_2424,In_2052);
nand U3339 (N_3339,In_617,In_474);
and U3340 (N_3340,In_921,In_2368);
or U3341 (N_3341,In_1365,In_1795);
or U3342 (N_3342,In_927,In_1473);
and U3343 (N_3343,In_1596,In_2441);
nand U3344 (N_3344,In_939,In_1016);
nand U3345 (N_3345,In_2286,In_1501);
nor U3346 (N_3346,In_2366,In_650);
and U3347 (N_3347,In_2440,In_330);
nor U3348 (N_3348,In_1387,In_154);
nand U3349 (N_3349,In_1277,In_821);
or U3350 (N_3350,In_682,In_664);
nand U3351 (N_3351,In_521,In_1284);
nand U3352 (N_3352,In_1710,In_1371);
and U3353 (N_3353,In_183,In_1399);
nor U3354 (N_3354,In_1930,In_226);
nor U3355 (N_3355,In_2026,In_153);
or U3356 (N_3356,In_1683,In_2163);
nand U3357 (N_3357,In_331,In_2371);
xnor U3358 (N_3358,In_2343,In_2290);
or U3359 (N_3359,In_1269,In_704);
and U3360 (N_3360,In_78,In_317);
nand U3361 (N_3361,In_1124,In_1357);
nand U3362 (N_3362,In_547,In_843);
or U3363 (N_3363,In_1430,In_539);
or U3364 (N_3364,In_1175,In_92);
or U3365 (N_3365,In_823,In_179);
or U3366 (N_3366,In_1010,In_439);
or U3367 (N_3367,In_1299,In_571);
or U3368 (N_3368,In_1595,In_551);
and U3369 (N_3369,In_846,In_900);
nor U3370 (N_3370,In_1104,In_716);
xor U3371 (N_3371,In_473,In_2465);
nand U3372 (N_3372,In_1643,In_37);
or U3373 (N_3373,In_2352,In_1383);
or U3374 (N_3374,In_634,In_813);
nand U3375 (N_3375,In_354,In_1663);
and U3376 (N_3376,In_740,In_464);
or U3377 (N_3377,In_378,In_292);
xor U3378 (N_3378,In_1022,In_1659);
nor U3379 (N_3379,In_1584,In_702);
or U3380 (N_3380,In_1205,In_1167);
and U3381 (N_3381,In_913,In_88);
and U3382 (N_3382,In_1363,In_1661);
and U3383 (N_3383,In_501,In_1070);
nor U3384 (N_3384,In_2316,In_2472);
and U3385 (N_3385,In_1046,In_2008);
and U3386 (N_3386,In_2149,In_1969);
nand U3387 (N_3387,In_1601,In_250);
and U3388 (N_3388,In_1904,In_100);
nand U3389 (N_3389,In_556,In_1732);
xnor U3390 (N_3390,In_957,In_1989);
and U3391 (N_3391,In_1967,In_249);
nor U3392 (N_3392,In_971,In_287);
and U3393 (N_3393,In_1678,In_1016);
nor U3394 (N_3394,In_2243,In_291);
and U3395 (N_3395,In_148,In_1737);
and U3396 (N_3396,In_414,In_1836);
nand U3397 (N_3397,In_69,In_1483);
xnor U3398 (N_3398,In_1388,In_1629);
and U3399 (N_3399,In_1565,In_1158);
nor U3400 (N_3400,In_1406,In_2354);
xor U3401 (N_3401,In_810,In_1639);
and U3402 (N_3402,In_1789,In_1617);
or U3403 (N_3403,In_573,In_973);
nand U3404 (N_3404,In_758,In_526);
and U3405 (N_3405,In_157,In_1620);
or U3406 (N_3406,In_1273,In_1552);
and U3407 (N_3407,In_1429,In_573);
nand U3408 (N_3408,In_434,In_227);
nor U3409 (N_3409,In_862,In_406);
and U3410 (N_3410,In_940,In_903);
nor U3411 (N_3411,In_2171,In_1913);
nand U3412 (N_3412,In_1150,In_988);
or U3413 (N_3413,In_2472,In_725);
or U3414 (N_3414,In_515,In_1283);
xnor U3415 (N_3415,In_1884,In_2105);
nor U3416 (N_3416,In_1972,In_401);
or U3417 (N_3417,In_534,In_1114);
and U3418 (N_3418,In_500,In_2499);
and U3419 (N_3419,In_581,In_596);
nor U3420 (N_3420,In_2040,In_2049);
and U3421 (N_3421,In_1505,In_1176);
and U3422 (N_3422,In_1773,In_2052);
xnor U3423 (N_3423,In_825,In_1326);
or U3424 (N_3424,In_1138,In_577);
nor U3425 (N_3425,In_837,In_2372);
xnor U3426 (N_3426,In_654,In_2446);
nor U3427 (N_3427,In_1104,In_2023);
and U3428 (N_3428,In_746,In_588);
nor U3429 (N_3429,In_112,In_1976);
or U3430 (N_3430,In_74,In_2137);
and U3431 (N_3431,In_993,In_1947);
nand U3432 (N_3432,In_1789,In_299);
nand U3433 (N_3433,In_849,In_699);
nor U3434 (N_3434,In_2408,In_1070);
xor U3435 (N_3435,In_1937,In_2421);
nor U3436 (N_3436,In_295,In_1001);
xor U3437 (N_3437,In_1322,In_2046);
nor U3438 (N_3438,In_2360,In_2414);
and U3439 (N_3439,In_2045,In_235);
or U3440 (N_3440,In_2422,In_1131);
nand U3441 (N_3441,In_1291,In_301);
nor U3442 (N_3442,In_163,In_2308);
xnor U3443 (N_3443,In_1292,In_2050);
or U3444 (N_3444,In_212,In_1121);
and U3445 (N_3445,In_1838,In_2425);
or U3446 (N_3446,In_2416,In_1295);
nand U3447 (N_3447,In_472,In_1822);
or U3448 (N_3448,In_709,In_1788);
nor U3449 (N_3449,In_617,In_2201);
or U3450 (N_3450,In_1921,In_1674);
and U3451 (N_3451,In_1100,In_1355);
and U3452 (N_3452,In_238,In_1794);
nand U3453 (N_3453,In_1948,In_2386);
nand U3454 (N_3454,In_1011,In_78);
nor U3455 (N_3455,In_938,In_2259);
nand U3456 (N_3456,In_1867,In_1973);
xnor U3457 (N_3457,In_943,In_723);
or U3458 (N_3458,In_1239,In_1855);
or U3459 (N_3459,In_1460,In_264);
nand U3460 (N_3460,In_835,In_543);
nand U3461 (N_3461,In_2347,In_2146);
and U3462 (N_3462,In_743,In_1471);
and U3463 (N_3463,In_1447,In_2069);
nand U3464 (N_3464,In_2169,In_1672);
or U3465 (N_3465,In_1641,In_1693);
nand U3466 (N_3466,In_1686,In_1242);
xnor U3467 (N_3467,In_1450,In_867);
or U3468 (N_3468,In_2089,In_2165);
or U3469 (N_3469,In_1134,In_541);
nand U3470 (N_3470,In_2305,In_441);
and U3471 (N_3471,In_2478,In_2226);
xnor U3472 (N_3472,In_1131,In_1182);
or U3473 (N_3473,In_1723,In_788);
or U3474 (N_3474,In_28,In_582);
nand U3475 (N_3475,In_1316,In_1165);
nor U3476 (N_3476,In_174,In_878);
nor U3477 (N_3477,In_1374,In_793);
and U3478 (N_3478,In_1649,In_1866);
or U3479 (N_3479,In_83,In_242);
nor U3480 (N_3480,In_2436,In_102);
nor U3481 (N_3481,In_1091,In_1351);
nor U3482 (N_3482,In_688,In_234);
nand U3483 (N_3483,In_136,In_1091);
nand U3484 (N_3484,In_2300,In_2165);
nand U3485 (N_3485,In_1524,In_2018);
and U3486 (N_3486,In_784,In_1933);
or U3487 (N_3487,In_1563,In_1575);
nor U3488 (N_3488,In_1421,In_385);
xnor U3489 (N_3489,In_263,In_160);
nand U3490 (N_3490,In_379,In_2112);
and U3491 (N_3491,In_1261,In_2230);
or U3492 (N_3492,In_1212,In_980);
nor U3493 (N_3493,In_2303,In_1389);
or U3494 (N_3494,In_1895,In_1440);
or U3495 (N_3495,In_1577,In_2286);
and U3496 (N_3496,In_1762,In_1827);
or U3497 (N_3497,In_901,In_2345);
nor U3498 (N_3498,In_1304,In_597);
or U3499 (N_3499,In_2151,In_1934);
or U3500 (N_3500,In_1677,In_1472);
nor U3501 (N_3501,In_1749,In_2005);
and U3502 (N_3502,In_674,In_2080);
xor U3503 (N_3503,In_1014,In_2223);
and U3504 (N_3504,In_258,In_999);
or U3505 (N_3505,In_1857,In_472);
nand U3506 (N_3506,In_1555,In_158);
nand U3507 (N_3507,In_1324,In_146);
or U3508 (N_3508,In_783,In_2130);
or U3509 (N_3509,In_2436,In_508);
nor U3510 (N_3510,In_1379,In_558);
or U3511 (N_3511,In_2100,In_964);
nand U3512 (N_3512,In_2365,In_2004);
or U3513 (N_3513,In_2472,In_475);
and U3514 (N_3514,In_2413,In_1425);
xor U3515 (N_3515,In_945,In_2025);
nand U3516 (N_3516,In_621,In_2232);
nand U3517 (N_3517,In_41,In_2379);
xnor U3518 (N_3518,In_428,In_1454);
or U3519 (N_3519,In_1959,In_2147);
nor U3520 (N_3520,In_2149,In_1094);
or U3521 (N_3521,In_1377,In_371);
nor U3522 (N_3522,In_1051,In_1174);
nor U3523 (N_3523,In_1247,In_907);
and U3524 (N_3524,In_1309,In_2227);
xor U3525 (N_3525,In_1111,In_324);
or U3526 (N_3526,In_1054,In_228);
or U3527 (N_3527,In_1044,In_1672);
or U3528 (N_3528,In_1913,In_2436);
or U3529 (N_3529,In_823,In_2191);
or U3530 (N_3530,In_1463,In_922);
or U3531 (N_3531,In_601,In_946);
and U3532 (N_3532,In_833,In_1924);
nor U3533 (N_3533,In_904,In_865);
nand U3534 (N_3534,In_1349,In_1769);
nor U3535 (N_3535,In_2083,In_1686);
nand U3536 (N_3536,In_869,In_1938);
nor U3537 (N_3537,In_1866,In_2423);
and U3538 (N_3538,In_1061,In_1886);
or U3539 (N_3539,In_755,In_2431);
nor U3540 (N_3540,In_2263,In_962);
nor U3541 (N_3541,In_583,In_1739);
or U3542 (N_3542,In_1829,In_647);
or U3543 (N_3543,In_639,In_32);
or U3544 (N_3544,In_2395,In_1760);
xor U3545 (N_3545,In_821,In_2327);
or U3546 (N_3546,In_1518,In_1556);
xnor U3547 (N_3547,In_796,In_1386);
xor U3548 (N_3548,In_108,In_973);
nor U3549 (N_3549,In_1947,In_2492);
nand U3550 (N_3550,In_1171,In_158);
nand U3551 (N_3551,In_440,In_1964);
nor U3552 (N_3552,In_838,In_2381);
or U3553 (N_3553,In_251,In_1938);
xor U3554 (N_3554,In_1909,In_502);
nor U3555 (N_3555,In_252,In_2065);
nor U3556 (N_3556,In_345,In_117);
and U3557 (N_3557,In_2029,In_2489);
and U3558 (N_3558,In_1292,In_429);
and U3559 (N_3559,In_2381,In_1781);
nor U3560 (N_3560,In_754,In_2492);
xor U3561 (N_3561,In_644,In_1903);
xnor U3562 (N_3562,In_1836,In_802);
nand U3563 (N_3563,In_405,In_840);
nor U3564 (N_3564,In_2453,In_2462);
and U3565 (N_3565,In_1685,In_628);
nor U3566 (N_3566,In_2344,In_732);
nor U3567 (N_3567,In_1703,In_1884);
nand U3568 (N_3568,In_1922,In_717);
or U3569 (N_3569,In_1969,In_307);
nor U3570 (N_3570,In_864,In_1140);
nand U3571 (N_3571,In_1257,In_1757);
and U3572 (N_3572,In_2145,In_970);
and U3573 (N_3573,In_418,In_213);
nor U3574 (N_3574,In_10,In_551);
and U3575 (N_3575,In_115,In_1833);
nor U3576 (N_3576,In_832,In_854);
nor U3577 (N_3577,In_1229,In_944);
and U3578 (N_3578,In_1978,In_465);
and U3579 (N_3579,In_963,In_1403);
xor U3580 (N_3580,In_1403,In_134);
or U3581 (N_3581,In_48,In_1337);
and U3582 (N_3582,In_1737,In_1427);
nor U3583 (N_3583,In_272,In_1248);
nand U3584 (N_3584,In_1699,In_1147);
and U3585 (N_3585,In_672,In_885);
or U3586 (N_3586,In_1699,In_455);
or U3587 (N_3587,In_744,In_689);
nor U3588 (N_3588,In_2339,In_599);
nand U3589 (N_3589,In_2033,In_1052);
and U3590 (N_3590,In_591,In_909);
and U3591 (N_3591,In_601,In_837);
xor U3592 (N_3592,In_673,In_177);
and U3593 (N_3593,In_1668,In_1429);
or U3594 (N_3594,In_1843,In_463);
nand U3595 (N_3595,In_1426,In_2134);
and U3596 (N_3596,In_230,In_1531);
or U3597 (N_3597,In_503,In_2186);
xor U3598 (N_3598,In_1256,In_301);
nand U3599 (N_3599,In_2407,In_574);
nand U3600 (N_3600,In_642,In_2396);
and U3601 (N_3601,In_533,In_446);
and U3602 (N_3602,In_1349,In_1027);
and U3603 (N_3603,In_348,In_1641);
nor U3604 (N_3604,In_49,In_1705);
nand U3605 (N_3605,In_1450,In_2231);
xnor U3606 (N_3606,In_953,In_242);
or U3607 (N_3607,In_2345,In_334);
xor U3608 (N_3608,In_406,In_37);
or U3609 (N_3609,In_1888,In_2396);
or U3610 (N_3610,In_1260,In_1082);
or U3611 (N_3611,In_978,In_750);
nand U3612 (N_3612,In_1891,In_2410);
nand U3613 (N_3613,In_1786,In_2322);
nor U3614 (N_3614,In_536,In_2300);
and U3615 (N_3615,In_1823,In_241);
nor U3616 (N_3616,In_1418,In_1335);
nand U3617 (N_3617,In_1266,In_1404);
and U3618 (N_3618,In_222,In_379);
nor U3619 (N_3619,In_630,In_821);
nand U3620 (N_3620,In_461,In_852);
nand U3621 (N_3621,In_298,In_42);
or U3622 (N_3622,In_2496,In_149);
nand U3623 (N_3623,In_328,In_626);
xor U3624 (N_3624,In_749,In_2065);
and U3625 (N_3625,In_2404,In_20);
and U3626 (N_3626,In_273,In_1765);
nor U3627 (N_3627,In_397,In_273);
xnor U3628 (N_3628,In_1283,In_993);
and U3629 (N_3629,In_999,In_1);
nor U3630 (N_3630,In_1541,In_1109);
nor U3631 (N_3631,In_1159,In_1121);
nand U3632 (N_3632,In_1592,In_2406);
xnor U3633 (N_3633,In_2347,In_1343);
nor U3634 (N_3634,In_1513,In_1338);
nand U3635 (N_3635,In_2009,In_958);
nor U3636 (N_3636,In_1244,In_1751);
and U3637 (N_3637,In_2332,In_2007);
xnor U3638 (N_3638,In_1644,In_1075);
or U3639 (N_3639,In_1782,In_1081);
nand U3640 (N_3640,In_1928,In_1773);
nor U3641 (N_3641,In_869,In_2223);
and U3642 (N_3642,In_1758,In_2413);
nor U3643 (N_3643,In_1995,In_2216);
or U3644 (N_3644,In_1808,In_1077);
or U3645 (N_3645,In_442,In_1888);
and U3646 (N_3646,In_1255,In_936);
or U3647 (N_3647,In_2096,In_1974);
nand U3648 (N_3648,In_1791,In_2104);
and U3649 (N_3649,In_2401,In_123);
nand U3650 (N_3650,In_2181,In_1517);
nand U3651 (N_3651,In_2409,In_711);
nand U3652 (N_3652,In_2459,In_1350);
or U3653 (N_3653,In_913,In_1517);
or U3654 (N_3654,In_259,In_2122);
and U3655 (N_3655,In_1526,In_1534);
nor U3656 (N_3656,In_64,In_610);
nand U3657 (N_3657,In_1728,In_1586);
nor U3658 (N_3658,In_178,In_614);
xor U3659 (N_3659,In_905,In_1136);
nand U3660 (N_3660,In_1267,In_485);
xor U3661 (N_3661,In_1339,In_2062);
and U3662 (N_3662,In_84,In_515);
and U3663 (N_3663,In_1439,In_63);
and U3664 (N_3664,In_1719,In_1170);
nand U3665 (N_3665,In_1165,In_488);
nand U3666 (N_3666,In_241,In_198);
nor U3667 (N_3667,In_1507,In_918);
and U3668 (N_3668,In_2228,In_1970);
or U3669 (N_3669,In_344,In_811);
nor U3670 (N_3670,In_765,In_2478);
and U3671 (N_3671,In_493,In_1518);
and U3672 (N_3672,In_1642,In_701);
nand U3673 (N_3673,In_724,In_994);
and U3674 (N_3674,In_788,In_192);
nand U3675 (N_3675,In_2062,In_236);
nor U3676 (N_3676,In_8,In_882);
xor U3677 (N_3677,In_1846,In_388);
nand U3678 (N_3678,In_2197,In_1284);
nand U3679 (N_3679,In_30,In_1846);
nor U3680 (N_3680,In_963,In_1342);
and U3681 (N_3681,In_754,In_1816);
and U3682 (N_3682,In_2233,In_590);
or U3683 (N_3683,In_714,In_613);
nand U3684 (N_3684,In_1796,In_1143);
xor U3685 (N_3685,In_1923,In_489);
nand U3686 (N_3686,In_2262,In_1870);
nand U3687 (N_3687,In_2281,In_1547);
and U3688 (N_3688,In_827,In_1486);
or U3689 (N_3689,In_1183,In_1559);
and U3690 (N_3690,In_1452,In_59);
nand U3691 (N_3691,In_1287,In_2064);
nand U3692 (N_3692,In_1876,In_2179);
nor U3693 (N_3693,In_247,In_160);
xor U3694 (N_3694,In_600,In_392);
and U3695 (N_3695,In_1691,In_190);
or U3696 (N_3696,In_1001,In_2257);
nor U3697 (N_3697,In_2180,In_744);
nand U3698 (N_3698,In_1998,In_1441);
and U3699 (N_3699,In_54,In_1742);
and U3700 (N_3700,In_723,In_1027);
nor U3701 (N_3701,In_2460,In_1262);
nor U3702 (N_3702,In_465,In_1777);
nand U3703 (N_3703,In_1217,In_662);
and U3704 (N_3704,In_557,In_769);
and U3705 (N_3705,In_1573,In_2478);
nand U3706 (N_3706,In_1221,In_61);
or U3707 (N_3707,In_1601,In_1058);
and U3708 (N_3708,In_1913,In_539);
nor U3709 (N_3709,In_1148,In_808);
nor U3710 (N_3710,In_849,In_1132);
xor U3711 (N_3711,In_90,In_1504);
nor U3712 (N_3712,In_1274,In_383);
or U3713 (N_3713,In_471,In_286);
or U3714 (N_3714,In_1173,In_261);
xor U3715 (N_3715,In_585,In_425);
and U3716 (N_3716,In_958,In_393);
nor U3717 (N_3717,In_108,In_1648);
or U3718 (N_3718,In_2475,In_216);
nand U3719 (N_3719,In_1676,In_1316);
nor U3720 (N_3720,In_1271,In_760);
nor U3721 (N_3721,In_1667,In_1485);
or U3722 (N_3722,In_996,In_258);
or U3723 (N_3723,In_808,In_461);
and U3724 (N_3724,In_436,In_248);
and U3725 (N_3725,In_2388,In_105);
nand U3726 (N_3726,In_120,In_165);
and U3727 (N_3727,In_2141,In_1080);
or U3728 (N_3728,In_212,In_217);
nor U3729 (N_3729,In_1771,In_1033);
nand U3730 (N_3730,In_2360,In_2011);
and U3731 (N_3731,In_1329,In_2245);
xnor U3732 (N_3732,In_18,In_2000);
nor U3733 (N_3733,In_624,In_1350);
nand U3734 (N_3734,In_1477,In_1336);
or U3735 (N_3735,In_1061,In_751);
and U3736 (N_3736,In_2027,In_1917);
or U3737 (N_3737,In_1423,In_1270);
nand U3738 (N_3738,In_1426,In_518);
nor U3739 (N_3739,In_964,In_2481);
nor U3740 (N_3740,In_1267,In_1006);
nand U3741 (N_3741,In_1916,In_2126);
nand U3742 (N_3742,In_1310,In_773);
nand U3743 (N_3743,In_2127,In_1984);
nor U3744 (N_3744,In_2258,In_1797);
or U3745 (N_3745,In_1534,In_87);
nand U3746 (N_3746,In_602,In_481);
or U3747 (N_3747,In_461,In_2077);
nand U3748 (N_3748,In_124,In_1207);
nand U3749 (N_3749,In_1754,In_913);
nand U3750 (N_3750,In_525,In_430);
and U3751 (N_3751,In_483,In_1743);
nor U3752 (N_3752,In_425,In_351);
nor U3753 (N_3753,In_1241,In_253);
nand U3754 (N_3754,In_1854,In_348);
nor U3755 (N_3755,In_697,In_1672);
or U3756 (N_3756,In_318,In_1302);
or U3757 (N_3757,In_1118,In_1187);
and U3758 (N_3758,In_602,In_695);
or U3759 (N_3759,In_941,In_2260);
or U3760 (N_3760,In_1222,In_1152);
xnor U3761 (N_3761,In_1674,In_945);
or U3762 (N_3762,In_663,In_424);
nand U3763 (N_3763,In_977,In_1027);
or U3764 (N_3764,In_1061,In_2454);
or U3765 (N_3765,In_562,In_1449);
or U3766 (N_3766,In_553,In_112);
nor U3767 (N_3767,In_1421,In_1225);
or U3768 (N_3768,In_16,In_1340);
and U3769 (N_3769,In_2394,In_1913);
nand U3770 (N_3770,In_616,In_286);
or U3771 (N_3771,In_752,In_568);
xnor U3772 (N_3772,In_1418,In_251);
and U3773 (N_3773,In_31,In_1423);
nand U3774 (N_3774,In_2072,In_2082);
nor U3775 (N_3775,In_532,In_1181);
and U3776 (N_3776,In_1579,In_1177);
nand U3777 (N_3777,In_368,In_2038);
or U3778 (N_3778,In_886,In_120);
nand U3779 (N_3779,In_2493,In_701);
or U3780 (N_3780,In_501,In_1774);
nor U3781 (N_3781,In_800,In_351);
nand U3782 (N_3782,In_1618,In_166);
nor U3783 (N_3783,In_151,In_758);
or U3784 (N_3784,In_815,In_1168);
nand U3785 (N_3785,In_638,In_2375);
or U3786 (N_3786,In_2070,In_691);
and U3787 (N_3787,In_151,In_1477);
or U3788 (N_3788,In_2047,In_1725);
and U3789 (N_3789,In_1162,In_2315);
or U3790 (N_3790,In_1312,In_1659);
nor U3791 (N_3791,In_2250,In_1089);
and U3792 (N_3792,In_2418,In_1519);
nor U3793 (N_3793,In_353,In_511);
and U3794 (N_3794,In_1645,In_2125);
and U3795 (N_3795,In_401,In_1806);
nand U3796 (N_3796,In_1325,In_2237);
and U3797 (N_3797,In_154,In_1708);
nand U3798 (N_3798,In_1619,In_432);
or U3799 (N_3799,In_178,In_539);
or U3800 (N_3800,In_890,In_548);
nand U3801 (N_3801,In_546,In_1992);
nor U3802 (N_3802,In_1204,In_2279);
xnor U3803 (N_3803,In_1926,In_527);
nor U3804 (N_3804,In_343,In_1622);
or U3805 (N_3805,In_2354,In_2080);
xor U3806 (N_3806,In_1202,In_2374);
nor U3807 (N_3807,In_1638,In_1704);
and U3808 (N_3808,In_2131,In_94);
and U3809 (N_3809,In_899,In_774);
xnor U3810 (N_3810,In_274,In_321);
and U3811 (N_3811,In_761,In_2470);
or U3812 (N_3812,In_830,In_2146);
nor U3813 (N_3813,In_838,In_85);
and U3814 (N_3814,In_2150,In_1276);
and U3815 (N_3815,In_1219,In_420);
nor U3816 (N_3816,In_737,In_914);
and U3817 (N_3817,In_1317,In_1705);
xnor U3818 (N_3818,In_887,In_1265);
or U3819 (N_3819,In_105,In_726);
or U3820 (N_3820,In_155,In_1933);
or U3821 (N_3821,In_2460,In_1851);
nor U3822 (N_3822,In_448,In_875);
nor U3823 (N_3823,In_171,In_1329);
and U3824 (N_3824,In_215,In_1062);
xor U3825 (N_3825,In_2380,In_1976);
nand U3826 (N_3826,In_697,In_674);
or U3827 (N_3827,In_627,In_437);
nand U3828 (N_3828,In_2258,In_2191);
nor U3829 (N_3829,In_1603,In_1057);
nand U3830 (N_3830,In_1714,In_1686);
nand U3831 (N_3831,In_1480,In_1712);
nor U3832 (N_3832,In_1801,In_1878);
or U3833 (N_3833,In_182,In_972);
and U3834 (N_3834,In_2259,In_600);
or U3835 (N_3835,In_2423,In_2354);
nand U3836 (N_3836,In_1622,In_588);
and U3837 (N_3837,In_600,In_1667);
and U3838 (N_3838,In_2081,In_2080);
or U3839 (N_3839,In_1319,In_1283);
nand U3840 (N_3840,In_1896,In_1755);
and U3841 (N_3841,In_1360,In_128);
nor U3842 (N_3842,In_518,In_2176);
and U3843 (N_3843,In_536,In_1892);
nor U3844 (N_3844,In_192,In_14);
nand U3845 (N_3845,In_87,In_1808);
nand U3846 (N_3846,In_1110,In_874);
nor U3847 (N_3847,In_145,In_940);
nor U3848 (N_3848,In_246,In_2223);
or U3849 (N_3849,In_120,In_818);
nand U3850 (N_3850,In_957,In_1338);
or U3851 (N_3851,In_266,In_610);
nand U3852 (N_3852,In_1646,In_27);
and U3853 (N_3853,In_1829,In_116);
and U3854 (N_3854,In_246,In_1613);
or U3855 (N_3855,In_1681,In_1257);
and U3856 (N_3856,In_1035,In_78);
nand U3857 (N_3857,In_1889,In_2484);
or U3858 (N_3858,In_1196,In_1577);
nand U3859 (N_3859,In_1032,In_2449);
nand U3860 (N_3860,In_1922,In_1050);
nand U3861 (N_3861,In_2122,In_657);
nand U3862 (N_3862,In_2095,In_800);
or U3863 (N_3863,In_1694,In_348);
nor U3864 (N_3864,In_1071,In_2471);
nand U3865 (N_3865,In_1180,In_1768);
and U3866 (N_3866,In_2067,In_1928);
or U3867 (N_3867,In_2197,In_59);
or U3868 (N_3868,In_634,In_18);
xnor U3869 (N_3869,In_1045,In_2428);
and U3870 (N_3870,In_2038,In_645);
nor U3871 (N_3871,In_1750,In_2262);
and U3872 (N_3872,In_1810,In_1123);
or U3873 (N_3873,In_819,In_1072);
nand U3874 (N_3874,In_254,In_2235);
and U3875 (N_3875,In_1302,In_585);
and U3876 (N_3876,In_1666,In_894);
nand U3877 (N_3877,In_1172,In_1323);
and U3878 (N_3878,In_1151,In_2061);
nand U3879 (N_3879,In_1560,In_1565);
nor U3880 (N_3880,In_2033,In_2328);
or U3881 (N_3881,In_2029,In_1395);
nor U3882 (N_3882,In_307,In_533);
nand U3883 (N_3883,In_1514,In_935);
nand U3884 (N_3884,In_167,In_2190);
or U3885 (N_3885,In_1161,In_143);
or U3886 (N_3886,In_2228,In_238);
or U3887 (N_3887,In_1802,In_317);
or U3888 (N_3888,In_1788,In_1849);
nor U3889 (N_3889,In_432,In_1873);
xnor U3890 (N_3890,In_954,In_488);
nand U3891 (N_3891,In_992,In_1435);
xor U3892 (N_3892,In_437,In_1208);
or U3893 (N_3893,In_1346,In_1426);
nand U3894 (N_3894,In_1787,In_2352);
or U3895 (N_3895,In_989,In_874);
nand U3896 (N_3896,In_832,In_71);
nor U3897 (N_3897,In_437,In_2448);
nor U3898 (N_3898,In_2363,In_2400);
or U3899 (N_3899,In_2293,In_601);
nor U3900 (N_3900,In_434,In_2017);
or U3901 (N_3901,In_295,In_2458);
or U3902 (N_3902,In_463,In_1556);
nand U3903 (N_3903,In_2465,In_21);
xor U3904 (N_3904,In_2355,In_571);
xnor U3905 (N_3905,In_892,In_1912);
and U3906 (N_3906,In_122,In_554);
nand U3907 (N_3907,In_1869,In_376);
xnor U3908 (N_3908,In_2033,In_1809);
nand U3909 (N_3909,In_2082,In_1191);
nand U3910 (N_3910,In_2301,In_1397);
or U3911 (N_3911,In_502,In_1367);
nand U3912 (N_3912,In_407,In_2299);
nor U3913 (N_3913,In_2201,In_2332);
xor U3914 (N_3914,In_1865,In_471);
nor U3915 (N_3915,In_1433,In_378);
and U3916 (N_3916,In_1924,In_834);
or U3917 (N_3917,In_629,In_374);
and U3918 (N_3918,In_1592,In_2065);
or U3919 (N_3919,In_866,In_594);
nor U3920 (N_3920,In_2424,In_1426);
or U3921 (N_3921,In_1422,In_820);
nand U3922 (N_3922,In_2423,In_2068);
and U3923 (N_3923,In_818,In_917);
nor U3924 (N_3924,In_1047,In_425);
nor U3925 (N_3925,In_982,In_1090);
nor U3926 (N_3926,In_425,In_2337);
nor U3927 (N_3927,In_1737,In_403);
and U3928 (N_3928,In_955,In_17);
nand U3929 (N_3929,In_904,In_966);
nor U3930 (N_3930,In_388,In_2486);
nor U3931 (N_3931,In_1305,In_270);
nand U3932 (N_3932,In_591,In_912);
xor U3933 (N_3933,In_841,In_368);
xor U3934 (N_3934,In_147,In_467);
nor U3935 (N_3935,In_2324,In_260);
xnor U3936 (N_3936,In_264,In_1732);
nand U3937 (N_3937,In_1991,In_2369);
or U3938 (N_3938,In_2115,In_1845);
and U3939 (N_3939,In_506,In_1160);
nor U3940 (N_3940,In_2267,In_187);
nand U3941 (N_3941,In_1271,In_1360);
nor U3942 (N_3942,In_911,In_165);
nor U3943 (N_3943,In_679,In_2306);
xor U3944 (N_3944,In_1051,In_227);
and U3945 (N_3945,In_1650,In_313);
or U3946 (N_3946,In_1854,In_2465);
xor U3947 (N_3947,In_2447,In_1447);
nand U3948 (N_3948,In_803,In_602);
or U3949 (N_3949,In_696,In_2299);
xor U3950 (N_3950,In_1733,In_1954);
or U3951 (N_3951,In_769,In_1889);
xnor U3952 (N_3952,In_2468,In_1214);
nor U3953 (N_3953,In_711,In_1029);
or U3954 (N_3954,In_1619,In_1841);
nor U3955 (N_3955,In_1803,In_102);
or U3956 (N_3956,In_1735,In_1241);
nand U3957 (N_3957,In_1563,In_214);
and U3958 (N_3958,In_1381,In_1100);
xor U3959 (N_3959,In_2403,In_1763);
nand U3960 (N_3960,In_2331,In_609);
nand U3961 (N_3961,In_111,In_2363);
nor U3962 (N_3962,In_156,In_2066);
or U3963 (N_3963,In_1814,In_192);
nand U3964 (N_3964,In_1410,In_313);
nor U3965 (N_3965,In_359,In_1130);
nand U3966 (N_3966,In_2293,In_1530);
or U3967 (N_3967,In_644,In_2226);
or U3968 (N_3968,In_338,In_1451);
and U3969 (N_3969,In_1136,In_1906);
nor U3970 (N_3970,In_766,In_1887);
and U3971 (N_3971,In_1608,In_2488);
nor U3972 (N_3972,In_1226,In_116);
and U3973 (N_3973,In_1054,In_1284);
or U3974 (N_3974,In_181,In_1627);
or U3975 (N_3975,In_2437,In_499);
nand U3976 (N_3976,In_938,In_2163);
nand U3977 (N_3977,In_2426,In_1849);
nand U3978 (N_3978,In_485,In_1599);
or U3979 (N_3979,In_918,In_1002);
nand U3980 (N_3980,In_1171,In_2204);
or U3981 (N_3981,In_746,In_1579);
xnor U3982 (N_3982,In_215,In_2294);
nand U3983 (N_3983,In_604,In_1972);
nor U3984 (N_3984,In_1866,In_1186);
nand U3985 (N_3985,In_1948,In_1815);
nor U3986 (N_3986,In_366,In_1938);
nand U3987 (N_3987,In_1988,In_760);
and U3988 (N_3988,In_244,In_1227);
nor U3989 (N_3989,In_205,In_985);
and U3990 (N_3990,In_886,In_1116);
xnor U3991 (N_3991,In_2095,In_1131);
nor U3992 (N_3992,In_209,In_1293);
and U3993 (N_3993,In_2343,In_1724);
xnor U3994 (N_3994,In_2108,In_1451);
nand U3995 (N_3995,In_430,In_906);
and U3996 (N_3996,In_377,In_1514);
nor U3997 (N_3997,In_1273,In_754);
or U3998 (N_3998,In_1827,In_390);
or U3999 (N_3999,In_5,In_1818);
nor U4000 (N_4000,In_1776,In_932);
xnor U4001 (N_4001,In_355,In_1676);
and U4002 (N_4002,In_1545,In_1990);
or U4003 (N_4003,In_1877,In_1168);
and U4004 (N_4004,In_862,In_1729);
and U4005 (N_4005,In_1405,In_1515);
nand U4006 (N_4006,In_2249,In_1147);
or U4007 (N_4007,In_1682,In_1913);
nor U4008 (N_4008,In_1376,In_2001);
nand U4009 (N_4009,In_636,In_535);
nand U4010 (N_4010,In_2419,In_1443);
nand U4011 (N_4011,In_758,In_1968);
nand U4012 (N_4012,In_2097,In_2450);
and U4013 (N_4013,In_1244,In_302);
nand U4014 (N_4014,In_504,In_479);
and U4015 (N_4015,In_1143,In_712);
or U4016 (N_4016,In_793,In_1605);
and U4017 (N_4017,In_2122,In_2351);
nand U4018 (N_4018,In_792,In_1942);
nor U4019 (N_4019,In_1599,In_1837);
nand U4020 (N_4020,In_846,In_907);
nor U4021 (N_4021,In_1570,In_711);
xor U4022 (N_4022,In_2438,In_2493);
and U4023 (N_4023,In_411,In_330);
and U4024 (N_4024,In_1574,In_633);
and U4025 (N_4025,In_897,In_2498);
and U4026 (N_4026,In_2258,In_362);
nor U4027 (N_4027,In_708,In_1008);
nand U4028 (N_4028,In_1829,In_1941);
and U4029 (N_4029,In_1767,In_300);
nand U4030 (N_4030,In_224,In_141);
nand U4031 (N_4031,In_835,In_2185);
and U4032 (N_4032,In_1185,In_857);
xnor U4033 (N_4033,In_404,In_99);
and U4034 (N_4034,In_1624,In_2449);
xnor U4035 (N_4035,In_802,In_1293);
or U4036 (N_4036,In_258,In_1703);
xor U4037 (N_4037,In_606,In_1606);
xor U4038 (N_4038,In_1285,In_1491);
and U4039 (N_4039,In_215,In_1274);
nor U4040 (N_4040,In_332,In_70);
xor U4041 (N_4041,In_132,In_2260);
and U4042 (N_4042,In_1563,In_619);
nor U4043 (N_4043,In_1702,In_1902);
nor U4044 (N_4044,In_1993,In_1644);
nand U4045 (N_4045,In_1994,In_42);
or U4046 (N_4046,In_570,In_2038);
nand U4047 (N_4047,In_1530,In_862);
or U4048 (N_4048,In_711,In_905);
or U4049 (N_4049,In_591,In_1518);
nor U4050 (N_4050,In_1096,In_1256);
or U4051 (N_4051,In_648,In_2276);
nand U4052 (N_4052,In_1432,In_1064);
nand U4053 (N_4053,In_236,In_1922);
nor U4054 (N_4054,In_7,In_776);
nand U4055 (N_4055,In_2,In_25);
or U4056 (N_4056,In_453,In_1967);
and U4057 (N_4057,In_309,In_180);
and U4058 (N_4058,In_1054,In_1324);
nand U4059 (N_4059,In_1778,In_116);
and U4060 (N_4060,In_1187,In_1563);
and U4061 (N_4061,In_2349,In_1983);
or U4062 (N_4062,In_439,In_354);
nor U4063 (N_4063,In_441,In_1880);
or U4064 (N_4064,In_1722,In_2015);
and U4065 (N_4065,In_1978,In_2075);
nor U4066 (N_4066,In_923,In_1790);
and U4067 (N_4067,In_2163,In_2470);
and U4068 (N_4068,In_916,In_2407);
nor U4069 (N_4069,In_1982,In_1635);
xnor U4070 (N_4070,In_1238,In_454);
nand U4071 (N_4071,In_1169,In_1744);
and U4072 (N_4072,In_2445,In_2466);
or U4073 (N_4073,In_2204,In_172);
xnor U4074 (N_4074,In_669,In_2336);
nand U4075 (N_4075,In_1912,In_2331);
nand U4076 (N_4076,In_442,In_500);
and U4077 (N_4077,In_975,In_1776);
xor U4078 (N_4078,In_2079,In_169);
nand U4079 (N_4079,In_840,In_888);
nor U4080 (N_4080,In_834,In_2467);
nor U4081 (N_4081,In_294,In_134);
xnor U4082 (N_4082,In_1557,In_1581);
xnor U4083 (N_4083,In_94,In_590);
or U4084 (N_4084,In_2007,In_1928);
nor U4085 (N_4085,In_1974,In_67);
or U4086 (N_4086,In_346,In_1530);
nor U4087 (N_4087,In_980,In_631);
nand U4088 (N_4088,In_42,In_1186);
nor U4089 (N_4089,In_359,In_304);
nand U4090 (N_4090,In_2286,In_1506);
and U4091 (N_4091,In_919,In_563);
or U4092 (N_4092,In_2310,In_1434);
nor U4093 (N_4093,In_506,In_732);
and U4094 (N_4094,In_299,In_941);
nor U4095 (N_4095,In_799,In_1488);
and U4096 (N_4096,In_1794,In_1586);
or U4097 (N_4097,In_682,In_2304);
and U4098 (N_4098,In_1017,In_75);
or U4099 (N_4099,In_1148,In_425);
nor U4100 (N_4100,In_2113,In_131);
nor U4101 (N_4101,In_1543,In_1179);
nor U4102 (N_4102,In_146,In_1775);
and U4103 (N_4103,In_310,In_260);
nand U4104 (N_4104,In_335,In_1898);
and U4105 (N_4105,In_471,In_823);
nand U4106 (N_4106,In_1099,In_997);
or U4107 (N_4107,In_2280,In_1717);
nand U4108 (N_4108,In_1378,In_348);
nor U4109 (N_4109,In_65,In_1040);
and U4110 (N_4110,In_1169,In_393);
nand U4111 (N_4111,In_964,In_750);
or U4112 (N_4112,In_194,In_2452);
and U4113 (N_4113,In_868,In_600);
or U4114 (N_4114,In_2443,In_1655);
nand U4115 (N_4115,In_401,In_2021);
or U4116 (N_4116,In_521,In_1181);
nand U4117 (N_4117,In_1960,In_1251);
nor U4118 (N_4118,In_962,In_1302);
nand U4119 (N_4119,In_419,In_158);
nand U4120 (N_4120,In_662,In_1033);
and U4121 (N_4121,In_2196,In_2444);
xor U4122 (N_4122,In_1773,In_2487);
and U4123 (N_4123,In_445,In_1930);
nand U4124 (N_4124,In_338,In_1369);
and U4125 (N_4125,In_1505,In_522);
nor U4126 (N_4126,In_845,In_809);
or U4127 (N_4127,In_954,In_385);
xnor U4128 (N_4128,In_889,In_1035);
and U4129 (N_4129,In_1997,In_2495);
or U4130 (N_4130,In_913,In_872);
nor U4131 (N_4131,In_2115,In_1919);
or U4132 (N_4132,In_2460,In_1436);
or U4133 (N_4133,In_2097,In_1637);
or U4134 (N_4134,In_1827,In_1491);
nand U4135 (N_4135,In_2107,In_2372);
or U4136 (N_4136,In_1104,In_1071);
or U4137 (N_4137,In_260,In_781);
and U4138 (N_4138,In_551,In_1637);
and U4139 (N_4139,In_2445,In_1241);
or U4140 (N_4140,In_2391,In_2454);
or U4141 (N_4141,In_1331,In_2328);
nand U4142 (N_4142,In_131,In_1199);
nor U4143 (N_4143,In_930,In_1250);
xnor U4144 (N_4144,In_407,In_1828);
and U4145 (N_4145,In_2492,In_2393);
or U4146 (N_4146,In_2494,In_383);
nand U4147 (N_4147,In_1607,In_160);
or U4148 (N_4148,In_268,In_267);
nand U4149 (N_4149,In_1199,In_514);
nand U4150 (N_4150,In_1796,In_519);
and U4151 (N_4151,In_1608,In_1197);
nor U4152 (N_4152,In_2080,In_2133);
nand U4153 (N_4153,In_2037,In_1410);
or U4154 (N_4154,In_1541,In_107);
and U4155 (N_4155,In_1914,In_844);
nor U4156 (N_4156,In_1953,In_2440);
and U4157 (N_4157,In_2043,In_2004);
or U4158 (N_4158,In_2486,In_887);
and U4159 (N_4159,In_217,In_1053);
nand U4160 (N_4160,In_1061,In_2175);
nor U4161 (N_4161,In_1898,In_1135);
nand U4162 (N_4162,In_2186,In_763);
nor U4163 (N_4163,In_1885,In_364);
or U4164 (N_4164,In_604,In_1575);
nand U4165 (N_4165,In_706,In_2246);
or U4166 (N_4166,In_285,In_923);
nand U4167 (N_4167,In_1219,In_1358);
nand U4168 (N_4168,In_1982,In_2018);
and U4169 (N_4169,In_245,In_2413);
and U4170 (N_4170,In_914,In_2445);
nor U4171 (N_4171,In_1713,In_654);
or U4172 (N_4172,In_673,In_111);
nand U4173 (N_4173,In_1339,In_1362);
and U4174 (N_4174,In_13,In_609);
nor U4175 (N_4175,In_1984,In_2034);
nor U4176 (N_4176,In_130,In_1493);
nand U4177 (N_4177,In_1947,In_1972);
xor U4178 (N_4178,In_915,In_1924);
and U4179 (N_4179,In_314,In_1165);
and U4180 (N_4180,In_1496,In_2331);
or U4181 (N_4181,In_1396,In_637);
nor U4182 (N_4182,In_900,In_1780);
nand U4183 (N_4183,In_2070,In_1696);
and U4184 (N_4184,In_2427,In_2486);
and U4185 (N_4185,In_1737,In_2299);
or U4186 (N_4186,In_1972,In_2097);
nand U4187 (N_4187,In_1458,In_738);
and U4188 (N_4188,In_1193,In_748);
or U4189 (N_4189,In_778,In_113);
or U4190 (N_4190,In_333,In_2458);
or U4191 (N_4191,In_778,In_1971);
and U4192 (N_4192,In_540,In_2000);
and U4193 (N_4193,In_548,In_1528);
nand U4194 (N_4194,In_1211,In_251);
and U4195 (N_4195,In_1757,In_613);
nand U4196 (N_4196,In_825,In_586);
or U4197 (N_4197,In_2089,In_2191);
or U4198 (N_4198,In_765,In_1247);
and U4199 (N_4199,In_799,In_2434);
nand U4200 (N_4200,In_1327,In_2438);
nor U4201 (N_4201,In_1115,In_2460);
nand U4202 (N_4202,In_1871,In_2002);
nand U4203 (N_4203,In_1907,In_2400);
nand U4204 (N_4204,In_1988,In_1557);
nor U4205 (N_4205,In_919,In_310);
or U4206 (N_4206,In_2303,In_536);
or U4207 (N_4207,In_1956,In_313);
nand U4208 (N_4208,In_907,In_1699);
nor U4209 (N_4209,In_359,In_1316);
or U4210 (N_4210,In_135,In_1202);
or U4211 (N_4211,In_635,In_736);
nor U4212 (N_4212,In_1478,In_1374);
or U4213 (N_4213,In_32,In_322);
or U4214 (N_4214,In_1607,In_2067);
and U4215 (N_4215,In_1353,In_2443);
and U4216 (N_4216,In_1583,In_265);
and U4217 (N_4217,In_2471,In_442);
or U4218 (N_4218,In_2136,In_2482);
or U4219 (N_4219,In_2187,In_591);
nor U4220 (N_4220,In_938,In_1688);
nor U4221 (N_4221,In_2130,In_2220);
or U4222 (N_4222,In_1075,In_1988);
and U4223 (N_4223,In_1732,In_75);
and U4224 (N_4224,In_1986,In_1601);
nand U4225 (N_4225,In_2301,In_1691);
nand U4226 (N_4226,In_1992,In_167);
nand U4227 (N_4227,In_1285,In_1556);
or U4228 (N_4228,In_1475,In_796);
and U4229 (N_4229,In_1915,In_227);
and U4230 (N_4230,In_2447,In_91);
and U4231 (N_4231,In_2186,In_1388);
xnor U4232 (N_4232,In_1040,In_1674);
nand U4233 (N_4233,In_692,In_36);
and U4234 (N_4234,In_1808,In_2133);
xnor U4235 (N_4235,In_1710,In_337);
or U4236 (N_4236,In_1425,In_1749);
or U4237 (N_4237,In_337,In_1501);
nor U4238 (N_4238,In_1011,In_311);
nor U4239 (N_4239,In_1420,In_934);
and U4240 (N_4240,In_20,In_2328);
nand U4241 (N_4241,In_1896,In_2212);
nand U4242 (N_4242,In_2331,In_1862);
nor U4243 (N_4243,In_2000,In_655);
nand U4244 (N_4244,In_254,In_36);
and U4245 (N_4245,In_1487,In_1332);
nand U4246 (N_4246,In_510,In_1491);
xor U4247 (N_4247,In_1161,In_1619);
or U4248 (N_4248,In_2302,In_515);
nor U4249 (N_4249,In_2051,In_942);
and U4250 (N_4250,In_1657,In_2165);
nor U4251 (N_4251,In_234,In_1277);
nand U4252 (N_4252,In_1531,In_337);
and U4253 (N_4253,In_2087,In_2370);
nor U4254 (N_4254,In_73,In_2139);
or U4255 (N_4255,In_2021,In_745);
and U4256 (N_4256,In_130,In_2049);
nor U4257 (N_4257,In_336,In_366);
and U4258 (N_4258,In_2062,In_1456);
xnor U4259 (N_4259,In_636,In_844);
nor U4260 (N_4260,In_2349,In_1619);
xnor U4261 (N_4261,In_1042,In_486);
nor U4262 (N_4262,In_1526,In_1162);
and U4263 (N_4263,In_324,In_2227);
or U4264 (N_4264,In_1437,In_1915);
nor U4265 (N_4265,In_2409,In_903);
and U4266 (N_4266,In_1106,In_2403);
xor U4267 (N_4267,In_765,In_1150);
nand U4268 (N_4268,In_1633,In_2329);
and U4269 (N_4269,In_614,In_1061);
nor U4270 (N_4270,In_647,In_1502);
nor U4271 (N_4271,In_531,In_230);
or U4272 (N_4272,In_1306,In_1830);
nor U4273 (N_4273,In_36,In_530);
and U4274 (N_4274,In_858,In_807);
nor U4275 (N_4275,In_262,In_2008);
xnor U4276 (N_4276,In_779,In_1416);
nor U4277 (N_4277,In_1602,In_2056);
and U4278 (N_4278,In_701,In_351);
or U4279 (N_4279,In_1341,In_2171);
and U4280 (N_4280,In_161,In_1247);
nor U4281 (N_4281,In_1452,In_1951);
and U4282 (N_4282,In_1666,In_2493);
or U4283 (N_4283,In_1643,In_1336);
nand U4284 (N_4284,In_1192,In_1760);
or U4285 (N_4285,In_1667,In_1844);
and U4286 (N_4286,In_946,In_1144);
nand U4287 (N_4287,In_2368,In_1016);
or U4288 (N_4288,In_123,In_143);
nor U4289 (N_4289,In_1957,In_283);
and U4290 (N_4290,In_2272,In_1161);
and U4291 (N_4291,In_1942,In_1374);
nor U4292 (N_4292,In_502,In_2421);
or U4293 (N_4293,In_1266,In_1320);
nand U4294 (N_4294,In_467,In_1884);
and U4295 (N_4295,In_1361,In_1739);
nand U4296 (N_4296,In_2383,In_467);
nand U4297 (N_4297,In_2018,In_2231);
and U4298 (N_4298,In_1342,In_2215);
or U4299 (N_4299,In_1429,In_101);
and U4300 (N_4300,In_1808,In_2135);
nand U4301 (N_4301,In_161,In_2369);
nor U4302 (N_4302,In_273,In_2116);
or U4303 (N_4303,In_534,In_2077);
or U4304 (N_4304,In_1063,In_2174);
nor U4305 (N_4305,In_2321,In_1693);
nand U4306 (N_4306,In_1276,In_638);
and U4307 (N_4307,In_1045,In_1460);
nand U4308 (N_4308,In_110,In_916);
or U4309 (N_4309,In_1771,In_1594);
nor U4310 (N_4310,In_564,In_1714);
nand U4311 (N_4311,In_2311,In_1466);
or U4312 (N_4312,In_1920,In_2443);
nor U4313 (N_4313,In_117,In_1531);
nand U4314 (N_4314,In_882,In_289);
xor U4315 (N_4315,In_2017,In_1415);
nor U4316 (N_4316,In_692,In_182);
and U4317 (N_4317,In_512,In_1414);
nand U4318 (N_4318,In_1851,In_1042);
and U4319 (N_4319,In_937,In_1724);
or U4320 (N_4320,In_520,In_2128);
nor U4321 (N_4321,In_797,In_62);
and U4322 (N_4322,In_1373,In_1555);
xnor U4323 (N_4323,In_1212,In_1966);
nand U4324 (N_4324,In_295,In_308);
or U4325 (N_4325,In_992,In_1268);
nor U4326 (N_4326,In_2490,In_2085);
or U4327 (N_4327,In_1724,In_972);
and U4328 (N_4328,In_111,In_713);
nor U4329 (N_4329,In_731,In_1270);
xor U4330 (N_4330,In_1455,In_1476);
nand U4331 (N_4331,In_1795,In_2103);
and U4332 (N_4332,In_251,In_1639);
nor U4333 (N_4333,In_602,In_1924);
xnor U4334 (N_4334,In_734,In_918);
nor U4335 (N_4335,In_1561,In_2040);
or U4336 (N_4336,In_1247,In_1851);
and U4337 (N_4337,In_2278,In_1262);
xnor U4338 (N_4338,In_254,In_663);
or U4339 (N_4339,In_115,In_2036);
or U4340 (N_4340,In_1382,In_398);
xnor U4341 (N_4341,In_624,In_1659);
or U4342 (N_4342,In_2107,In_1356);
and U4343 (N_4343,In_2103,In_237);
nor U4344 (N_4344,In_460,In_1110);
xnor U4345 (N_4345,In_683,In_2050);
nor U4346 (N_4346,In_1512,In_1491);
xnor U4347 (N_4347,In_1700,In_374);
nor U4348 (N_4348,In_1556,In_333);
xnor U4349 (N_4349,In_249,In_141);
nand U4350 (N_4350,In_1912,In_998);
nor U4351 (N_4351,In_709,In_2283);
nand U4352 (N_4352,In_429,In_1730);
and U4353 (N_4353,In_2037,In_2167);
xor U4354 (N_4354,In_370,In_1287);
and U4355 (N_4355,In_1193,In_119);
or U4356 (N_4356,In_351,In_1132);
nand U4357 (N_4357,In_107,In_2307);
and U4358 (N_4358,In_40,In_1997);
nor U4359 (N_4359,In_1678,In_989);
and U4360 (N_4360,In_2459,In_79);
nand U4361 (N_4361,In_1359,In_1836);
and U4362 (N_4362,In_939,In_1269);
nand U4363 (N_4363,In_966,In_478);
nand U4364 (N_4364,In_37,In_1277);
nor U4365 (N_4365,In_1419,In_139);
or U4366 (N_4366,In_551,In_545);
nand U4367 (N_4367,In_1159,In_1320);
or U4368 (N_4368,In_262,In_1876);
xnor U4369 (N_4369,In_1437,In_1037);
or U4370 (N_4370,In_1548,In_1144);
nor U4371 (N_4371,In_987,In_1790);
or U4372 (N_4372,In_1026,In_74);
nand U4373 (N_4373,In_1567,In_1705);
nor U4374 (N_4374,In_2015,In_693);
and U4375 (N_4375,In_2251,In_425);
nor U4376 (N_4376,In_2288,In_683);
nand U4377 (N_4377,In_96,In_8);
and U4378 (N_4378,In_450,In_1373);
nor U4379 (N_4379,In_1522,In_2272);
and U4380 (N_4380,In_113,In_375);
and U4381 (N_4381,In_2265,In_1957);
nor U4382 (N_4382,In_1647,In_576);
nor U4383 (N_4383,In_2424,In_635);
nand U4384 (N_4384,In_1334,In_2249);
nand U4385 (N_4385,In_1491,In_251);
or U4386 (N_4386,In_1337,In_1117);
and U4387 (N_4387,In_793,In_1847);
or U4388 (N_4388,In_1800,In_26);
nand U4389 (N_4389,In_2017,In_2034);
and U4390 (N_4390,In_325,In_1881);
xor U4391 (N_4391,In_12,In_1582);
and U4392 (N_4392,In_2274,In_1264);
or U4393 (N_4393,In_871,In_2066);
nand U4394 (N_4394,In_722,In_2377);
nor U4395 (N_4395,In_1146,In_2005);
nand U4396 (N_4396,In_461,In_1098);
nor U4397 (N_4397,In_2166,In_2244);
or U4398 (N_4398,In_1551,In_533);
nand U4399 (N_4399,In_629,In_1468);
and U4400 (N_4400,In_216,In_1816);
and U4401 (N_4401,In_2473,In_1580);
nor U4402 (N_4402,In_66,In_1652);
or U4403 (N_4403,In_93,In_8);
nor U4404 (N_4404,In_684,In_1421);
or U4405 (N_4405,In_1917,In_1696);
and U4406 (N_4406,In_2250,In_2246);
nor U4407 (N_4407,In_1003,In_1592);
xor U4408 (N_4408,In_1921,In_200);
and U4409 (N_4409,In_1877,In_1044);
nor U4410 (N_4410,In_615,In_404);
or U4411 (N_4411,In_1444,In_1479);
and U4412 (N_4412,In_1373,In_750);
or U4413 (N_4413,In_2447,In_1542);
or U4414 (N_4414,In_428,In_32);
nand U4415 (N_4415,In_1268,In_134);
and U4416 (N_4416,In_697,In_1071);
and U4417 (N_4417,In_769,In_1340);
xnor U4418 (N_4418,In_1386,In_1762);
or U4419 (N_4419,In_1430,In_1140);
or U4420 (N_4420,In_2100,In_638);
and U4421 (N_4421,In_1572,In_1916);
nand U4422 (N_4422,In_172,In_1143);
nor U4423 (N_4423,In_2412,In_1972);
and U4424 (N_4424,In_2106,In_1450);
and U4425 (N_4425,In_949,In_371);
or U4426 (N_4426,In_799,In_27);
or U4427 (N_4427,In_2128,In_117);
nor U4428 (N_4428,In_2494,In_1028);
nor U4429 (N_4429,In_392,In_730);
nand U4430 (N_4430,In_2440,In_2419);
xor U4431 (N_4431,In_54,In_1074);
nand U4432 (N_4432,In_10,In_588);
nand U4433 (N_4433,In_469,In_2243);
and U4434 (N_4434,In_1027,In_2415);
and U4435 (N_4435,In_2165,In_1214);
nand U4436 (N_4436,In_1698,In_949);
nand U4437 (N_4437,In_1506,In_1507);
nor U4438 (N_4438,In_728,In_1756);
nand U4439 (N_4439,In_1991,In_842);
nand U4440 (N_4440,In_2379,In_1364);
xnor U4441 (N_4441,In_814,In_833);
or U4442 (N_4442,In_2076,In_1065);
nor U4443 (N_4443,In_1280,In_1639);
xor U4444 (N_4444,In_1492,In_1199);
or U4445 (N_4445,In_1552,In_1826);
nor U4446 (N_4446,In_103,In_1147);
and U4447 (N_4447,In_2313,In_1873);
or U4448 (N_4448,In_1381,In_2012);
nand U4449 (N_4449,In_1321,In_640);
nor U4450 (N_4450,In_236,In_2069);
or U4451 (N_4451,In_2346,In_1219);
or U4452 (N_4452,In_135,In_1089);
nor U4453 (N_4453,In_1200,In_1690);
and U4454 (N_4454,In_1826,In_1072);
xnor U4455 (N_4455,In_2147,In_122);
and U4456 (N_4456,In_1658,In_922);
and U4457 (N_4457,In_1053,In_55);
and U4458 (N_4458,In_881,In_125);
nand U4459 (N_4459,In_90,In_920);
nand U4460 (N_4460,In_436,In_1239);
or U4461 (N_4461,In_2009,In_909);
nor U4462 (N_4462,In_1943,In_476);
nor U4463 (N_4463,In_490,In_1135);
or U4464 (N_4464,In_1523,In_1184);
and U4465 (N_4465,In_60,In_2356);
or U4466 (N_4466,In_696,In_862);
nand U4467 (N_4467,In_637,In_1558);
and U4468 (N_4468,In_1229,In_696);
nand U4469 (N_4469,In_2122,In_388);
and U4470 (N_4470,In_2160,In_1397);
nor U4471 (N_4471,In_2478,In_145);
and U4472 (N_4472,In_1232,In_2383);
nor U4473 (N_4473,In_1066,In_599);
or U4474 (N_4474,In_1255,In_755);
xor U4475 (N_4475,In_1274,In_326);
nand U4476 (N_4476,In_1956,In_729);
nand U4477 (N_4477,In_1575,In_628);
nand U4478 (N_4478,In_1018,In_1240);
and U4479 (N_4479,In_1175,In_238);
and U4480 (N_4480,In_27,In_854);
nand U4481 (N_4481,In_850,In_1108);
or U4482 (N_4482,In_177,In_444);
nand U4483 (N_4483,In_1657,In_876);
and U4484 (N_4484,In_24,In_540);
and U4485 (N_4485,In_339,In_670);
nor U4486 (N_4486,In_1985,In_1522);
nand U4487 (N_4487,In_1531,In_2146);
nor U4488 (N_4488,In_23,In_10);
nor U4489 (N_4489,In_1241,In_1992);
nand U4490 (N_4490,In_749,In_3);
nor U4491 (N_4491,In_1051,In_983);
xor U4492 (N_4492,In_454,In_624);
xor U4493 (N_4493,In_2082,In_365);
or U4494 (N_4494,In_177,In_1762);
nand U4495 (N_4495,In_2325,In_2285);
nor U4496 (N_4496,In_496,In_3);
nor U4497 (N_4497,In_1423,In_95);
nand U4498 (N_4498,In_1842,In_210);
xnor U4499 (N_4499,In_2274,In_1105);
and U4500 (N_4500,In_2262,In_2338);
or U4501 (N_4501,In_1705,In_467);
nand U4502 (N_4502,In_301,In_1325);
nor U4503 (N_4503,In_1783,In_1537);
or U4504 (N_4504,In_1500,In_1497);
or U4505 (N_4505,In_1804,In_1037);
nor U4506 (N_4506,In_2176,In_1301);
xnor U4507 (N_4507,In_801,In_2140);
or U4508 (N_4508,In_1428,In_591);
nor U4509 (N_4509,In_479,In_2073);
xor U4510 (N_4510,In_1205,In_1062);
or U4511 (N_4511,In_821,In_1391);
nor U4512 (N_4512,In_1951,In_2166);
xor U4513 (N_4513,In_2090,In_2207);
nor U4514 (N_4514,In_316,In_1249);
or U4515 (N_4515,In_767,In_354);
nor U4516 (N_4516,In_1847,In_836);
and U4517 (N_4517,In_2473,In_58);
nor U4518 (N_4518,In_2084,In_740);
or U4519 (N_4519,In_1942,In_2257);
or U4520 (N_4520,In_2427,In_202);
and U4521 (N_4521,In_514,In_2021);
xor U4522 (N_4522,In_392,In_1457);
nor U4523 (N_4523,In_1204,In_627);
and U4524 (N_4524,In_2096,In_1936);
xor U4525 (N_4525,In_144,In_2494);
or U4526 (N_4526,In_1887,In_1705);
and U4527 (N_4527,In_783,In_1336);
or U4528 (N_4528,In_82,In_2484);
nor U4529 (N_4529,In_835,In_703);
and U4530 (N_4530,In_1367,In_2289);
or U4531 (N_4531,In_1489,In_1620);
nor U4532 (N_4532,In_1290,In_749);
nand U4533 (N_4533,In_226,In_1836);
or U4534 (N_4534,In_1556,In_418);
and U4535 (N_4535,In_195,In_1645);
nor U4536 (N_4536,In_344,In_2179);
nand U4537 (N_4537,In_467,In_2258);
xnor U4538 (N_4538,In_1879,In_2163);
nor U4539 (N_4539,In_229,In_1289);
or U4540 (N_4540,In_1476,In_1220);
or U4541 (N_4541,In_433,In_1411);
or U4542 (N_4542,In_1218,In_295);
and U4543 (N_4543,In_1096,In_2193);
and U4544 (N_4544,In_1624,In_1784);
or U4545 (N_4545,In_1430,In_1103);
or U4546 (N_4546,In_2153,In_836);
nor U4547 (N_4547,In_2160,In_1390);
nor U4548 (N_4548,In_1783,In_271);
xor U4549 (N_4549,In_1200,In_668);
xnor U4550 (N_4550,In_2467,In_198);
or U4551 (N_4551,In_1580,In_1675);
and U4552 (N_4552,In_777,In_424);
nand U4553 (N_4553,In_2286,In_2251);
or U4554 (N_4554,In_805,In_611);
or U4555 (N_4555,In_999,In_2207);
or U4556 (N_4556,In_1743,In_1021);
and U4557 (N_4557,In_2167,In_198);
or U4558 (N_4558,In_2024,In_999);
and U4559 (N_4559,In_1968,In_1049);
and U4560 (N_4560,In_123,In_678);
or U4561 (N_4561,In_89,In_1518);
or U4562 (N_4562,In_1756,In_1733);
nor U4563 (N_4563,In_950,In_1196);
or U4564 (N_4564,In_524,In_1341);
or U4565 (N_4565,In_2034,In_214);
and U4566 (N_4566,In_2305,In_1627);
nand U4567 (N_4567,In_97,In_169);
and U4568 (N_4568,In_886,In_2280);
nor U4569 (N_4569,In_2027,In_949);
nand U4570 (N_4570,In_456,In_903);
xnor U4571 (N_4571,In_2025,In_671);
nor U4572 (N_4572,In_124,In_2388);
or U4573 (N_4573,In_327,In_1554);
and U4574 (N_4574,In_106,In_723);
xnor U4575 (N_4575,In_1134,In_1017);
or U4576 (N_4576,In_296,In_1336);
and U4577 (N_4577,In_1327,In_812);
or U4578 (N_4578,In_470,In_569);
nand U4579 (N_4579,In_369,In_876);
xnor U4580 (N_4580,In_952,In_1309);
nand U4581 (N_4581,In_1396,In_2474);
nor U4582 (N_4582,In_547,In_1044);
and U4583 (N_4583,In_1516,In_729);
xor U4584 (N_4584,In_236,In_972);
and U4585 (N_4585,In_1215,In_1369);
or U4586 (N_4586,In_1821,In_2033);
or U4587 (N_4587,In_1849,In_58);
nor U4588 (N_4588,In_1424,In_1547);
nor U4589 (N_4589,In_1824,In_1010);
or U4590 (N_4590,In_1961,In_2151);
xor U4591 (N_4591,In_2455,In_476);
nand U4592 (N_4592,In_2167,In_724);
and U4593 (N_4593,In_1235,In_1727);
nor U4594 (N_4594,In_2235,In_1915);
nor U4595 (N_4595,In_1964,In_787);
or U4596 (N_4596,In_768,In_2066);
nor U4597 (N_4597,In_1599,In_88);
xor U4598 (N_4598,In_1118,In_756);
and U4599 (N_4599,In_134,In_1398);
and U4600 (N_4600,In_845,In_660);
nor U4601 (N_4601,In_364,In_681);
nor U4602 (N_4602,In_2451,In_2490);
nor U4603 (N_4603,In_1739,In_2276);
or U4604 (N_4604,In_309,In_1567);
or U4605 (N_4605,In_1050,In_2030);
nor U4606 (N_4606,In_1338,In_281);
nor U4607 (N_4607,In_1001,In_1605);
and U4608 (N_4608,In_1090,In_1504);
nor U4609 (N_4609,In_1769,In_2328);
nor U4610 (N_4610,In_2004,In_377);
and U4611 (N_4611,In_2252,In_2467);
nand U4612 (N_4612,In_1097,In_1982);
and U4613 (N_4613,In_1776,In_615);
or U4614 (N_4614,In_1189,In_2335);
nor U4615 (N_4615,In_2421,In_475);
nand U4616 (N_4616,In_1045,In_2099);
or U4617 (N_4617,In_548,In_2414);
nor U4618 (N_4618,In_1160,In_270);
and U4619 (N_4619,In_157,In_2314);
xnor U4620 (N_4620,In_1352,In_2102);
nor U4621 (N_4621,In_1122,In_2348);
or U4622 (N_4622,In_1353,In_52);
xnor U4623 (N_4623,In_734,In_2150);
xnor U4624 (N_4624,In_909,In_1231);
nor U4625 (N_4625,In_1231,In_579);
nand U4626 (N_4626,In_323,In_254);
and U4627 (N_4627,In_1120,In_1214);
or U4628 (N_4628,In_1057,In_2239);
nand U4629 (N_4629,In_898,In_1754);
xnor U4630 (N_4630,In_1794,In_936);
nand U4631 (N_4631,In_762,In_2430);
or U4632 (N_4632,In_1315,In_2407);
nor U4633 (N_4633,In_545,In_401);
xor U4634 (N_4634,In_1330,In_779);
nand U4635 (N_4635,In_866,In_2196);
or U4636 (N_4636,In_439,In_643);
nor U4637 (N_4637,In_1556,In_1286);
and U4638 (N_4638,In_644,In_1176);
nor U4639 (N_4639,In_2301,In_50);
or U4640 (N_4640,In_855,In_1307);
or U4641 (N_4641,In_1499,In_422);
nor U4642 (N_4642,In_1946,In_1645);
nand U4643 (N_4643,In_2086,In_141);
and U4644 (N_4644,In_1259,In_1777);
nand U4645 (N_4645,In_2005,In_1243);
or U4646 (N_4646,In_2103,In_987);
or U4647 (N_4647,In_117,In_2110);
nor U4648 (N_4648,In_992,In_916);
nor U4649 (N_4649,In_2379,In_1695);
nor U4650 (N_4650,In_879,In_1873);
nor U4651 (N_4651,In_2171,In_2117);
and U4652 (N_4652,In_296,In_485);
and U4653 (N_4653,In_785,In_310);
or U4654 (N_4654,In_1076,In_261);
or U4655 (N_4655,In_2020,In_1862);
or U4656 (N_4656,In_2385,In_204);
nor U4657 (N_4657,In_1457,In_1848);
nor U4658 (N_4658,In_2068,In_764);
or U4659 (N_4659,In_1959,In_367);
nand U4660 (N_4660,In_2453,In_2119);
or U4661 (N_4661,In_574,In_1462);
xnor U4662 (N_4662,In_1666,In_2471);
nand U4663 (N_4663,In_2288,In_2097);
nor U4664 (N_4664,In_2001,In_1790);
xor U4665 (N_4665,In_1507,In_1306);
nand U4666 (N_4666,In_1932,In_1709);
and U4667 (N_4667,In_1589,In_1670);
nand U4668 (N_4668,In_2247,In_963);
or U4669 (N_4669,In_1750,In_1030);
nand U4670 (N_4670,In_745,In_497);
or U4671 (N_4671,In_2479,In_317);
or U4672 (N_4672,In_2190,In_1368);
or U4673 (N_4673,In_1335,In_1733);
nor U4674 (N_4674,In_625,In_1965);
nor U4675 (N_4675,In_606,In_1852);
or U4676 (N_4676,In_1860,In_42);
or U4677 (N_4677,In_589,In_697);
nor U4678 (N_4678,In_7,In_1714);
or U4679 (N_4679,In_1773,In_937);
nand U4680 (N_4680,In_625,In_1819);
and U4681 (N_4681,In_1665,In_1819);
nor U4682 (N_4682,In_1679,In_1593);
xnor U4683 (N_4683,In_2273,In_1220);
xnor U4684 (N_4684,In_2436,In_1459);
and U4685 (N_4685,In_266,In_2048);
and U4686 (N_4686,In_2382,In_1165);
nor U4687 (N_4687,In_1132,In_1247);
xor U4688 (N_4688,In_1239,In_516);
and U4689 (N_4689,In_351,In_1977);
and U4690 (N_4690,In_1586,In_1471);
and U4691 (N_4691,In_2220,In_637);
and U4692 (N_4692,In_1424,In_532);
nand U4693 (N_4693,In_1891,In_1813);
nand U4694 (N_4694,In_879,In_1155);
and U4695 (N_4695,In_1170,In_752);
xnor U4696 (N_4696,In_1822,In_2010);
and U4697 (N_4697,In_235,In_1467);
xor U4698 (N_4698,In_1399,In_92);
nand U4699 (N_4699,In_349,In_2029);
nand U4700 (N_4700,In_351,In_525);
or U4701 (N_4701,In_1567,In_949);
nor U4702 (N_4702,In_748,In_640);
nor U4703 (N_4703,In_2067,In_834);
nand U4704 (N_4704,In_219,In_2431);
and U4705 (N_4705,In_724,In_913);
or U4706 (N_4706,In_663,In_694);
nand U4707 (N_4707,In_627,In_455);
or U4708 (N_4708,In_294,In_755);
nor U4709 (N_4709,In_304,In_1593);
nand U4710 (N_4710,In_742,In_1948);
nor U4711 (N_4711,In_1236,In_877);
and U4712 (N_4712,In_448,In_651);
and U4713 (N_4713,In_875,In_2163);
and U4714 (N_4714,In_1265,In_2071);
or U4715 (N_4715,In_921,In_1577);
or U4716 (N_4716,In_484,In_2296);
and U4717 (N_4717,In_507,In_1883);
or U4718 (N_4718,In_914,In_2386);
nor U4719 (N_4719,In_1199,In_898);
nor U4720 (N_4720,In_944,In_318);
and U4721 (N_4721,In_946,In_2397);
nor U4722 (N_4722,In_392,In_2179);
nor U4723 (N_4723,In_1634,In_1496);
xor U4724 (N_4724,In_1502,In_1919);
and U4725 (N_4725,In_1975,In_924);
or U4726 (N_4726,In_2320,In_563);
or U4727 (N_4727,In_222,In_1022);
nor U4728 (N_4728,In_1653,In_118);
and U4729 (N_4729,In_2379,In_659);
or U4730 (N_4730,In_595,In_2267);
or U4731 (N_4731,In_863,In_844);
nand U4732 (N_4732,In_1923,In_1253);
nor U4733 (N_4733,In_1215,In_728);
nand U4734 (N_4734,In_1763,In_1293);
nand U4735 (N_4735,In_2145,In_1485);
or U4736 (N_4736,In_1746,In_467);
and U4737 (N_4737,In_1678,In_1250);
xnor U4738 (N_4738,In_257,In_1695);
nor U4739 (N_4739,In_612,In_2252);
and U4740 (N_4740,In_883,In_204);
nand U4741 (N_4741,In_56,In_1690);
nor U4742 (N_4742,In_555,In_153);
and U4743 (N_4743,In_1117,In_1012);
nor U4744 (N_4744,In_9,In_1864);
nand U4745 (N_4745,In_1876,In_556);
xor U4746 (N_4746,In_92,In_1389);
nand U4747 (N_4747,In_1610,In_2472);
nand U4748 (N_4748,In_2411,In_2051);
or U4749 (N_4749,In_2368,In_360);
nand U4750 (N_4750,In_1277,In_2010);
nand U4751 (N_4751,In_1980,In_1862);
nand U4752 (N_4752,In_614,In_337);
nor U4753 (N_4753,In_1445,In_276);
nor U4754 (N_4754,In_1171,In_1554);
nor U4755 (N_4755,In_842,In_100);
or U4756 (N_4756,In_1878,In_560);
and U4757 (N_4757,In_2318,In_2405);
nand U4758 (N_4758,In_528,In_339);
or U4759 (N_4759,In_1466,In_1033);
nor U4760 (N_4760,In_333,In_641);
nand U4761 (N_4761,In_1974,In_97);
nor U4762 (N_4762,In_1852,In_1134);
or U4763 (N_4763,In_509,In_188);
nand U4764 (N_4764,In_1548,In_113);
and U4765 (N_4765,In_1499,In_386);
nor U4766 (N_4766,In_366,In_599);
nand U4767 (N_4767,In_1955,In_1906);
or U4768 (N_4768,In_128,In_161);
or U4769 (N_4769,In_603,In_60);
and U4770 (N_4770,In_868,In_1052);
xnor U4771 (N_4771,In_2258,In_1946);
nor U4772 (N_4772,In_109,In_572);
and U4773 (N_4773,In_733,In_2173);
or U4774 (N_4774,In_1735,In_640);
nand U4775 (N_4775,In_465,In_2274);
nand U4776 (N_4776,In_2257,In_2019);
or U4777 (N_4777,In_122,In_518);
nand U4778 (N_4778,In_1508,In_1865);
nand U4779 (N_4779,In_1653,In_1084);
and U4780 (N_4780,In_1408,In_1777);
and U4781 (N_4781,In_2078,In_860);
and U4782 (N_4782,In_1831,In_2453);
nor U4783 (N_4783,In_1889,In_2011);
and U4784 (N_4784,In_2294,In_1359);
or U4785 (N_4785,In_551,In_2020);
nor U4786 (N_4786,In_436,In_1359);
nand U4787 (N_4787,In_1772,In_1202);
nor U4788 (N_4788,In_1427,In_623);
and U4789 (N_4789,In_1315,In_2440);
or U4790 (N_4790,In_821,In_1724);
or U4791 (N_4791,In_1183,In_65);
nand U4792 (N_4792,In_1784,In_1815);
and U4793 (N_4793,In_1601,In_1491);
xor U4794 (N_4794,In_1977,In_235);
nor U4795 (N_4795,In_1113,In_391);
nand U4796 (N_4796,In_336,In_1556);
nand U4797 (N_4797,In_2401,In_935);
or U4798 (N_4798,In_593,In_2401);
or U4799 (N_4799,In_969,In_1680);
nor U4800 (N_4800,In_615,In_532);
nand U4801 (N_4801,In_1593,In_2369);
or U4802 (N_4802,In_1858,In_916);
nand U4803 (N_4803,In_1021,In_476);
xor U4804 (N_4804,In_2145,In_348);
or U4805 (N_4805,In_1285,In_25);
nor U4806 (N_4806,In_2067,In_2229);
nor U4807 (N_4807,In_2254,In_2499);
and U4808 (N_4808,In_66,In_1367);
nand U4809 (N_4809,In_2414,In_1902);
and U4810 (N_4810,In_1672,In_2258);
and U4811 (N_4811,In_838,In_432);
or U4812 (N_4812,In_1014,In_1428);
nand U4813 (N_4813,In_1378,In_2080);
or U4814 (N_4814,In_613,In_1232);
nand U4815 (N_4815,In_2152,In_2352);
nand U4816 (N_4816,In_847,In_1187);
and U4817 (N_4817,In_426,In_1588);
xor U4818 (N_4818,In_1898,In_1470);
or U4819 (N_4819,In_31,In_1107);
or U4820 (N_4820,In_2264,In_1691);
xor U4821 (N_4821,In_1294,In_1188);
and U4822 (N_4822,In_505,In_1746);
or U4823 (N_4823,In_503,In_368);
and U4824 (N_4824,In_1152,In_1730);
nand U4825 (N_4825,In_187,In_1934);
nor U4826 (N_4826,In_968,In_325);
and U4827 (N_4827,In_268,In_120);
nand U4828 (N_4828,In_836,In_1532);
and U4829 (N_4829,In_2006,In_558);
nor U4830 (N_4830,In_1112,In_2372);
nor U4831 (N_4831,In_2218,In_325);
xnor U4832 (N_4832,In_1928,In_699);
and U4833 (N_4833,In_2300,In_1132);
and U4834 (N_4834,In_587,In_1388);
or U4835 (N_4835,In_220,In_286);
nand U4836 (N_4836,In_364,In_647);
nand U4837 (N_4837,In_671,In_1596);
or U4838 (N_4838,In_1780,In_175);
or U4839 (N_4839,In_2480,In_74);
or U4840 (N_4840,In_1605,In_1716);
and U4841 (N_4841,In_333,In_555);
or U4842 (N_4842,In_2436,In_136);
or U4843 (N_4843,In_92,In_1888);
or U4844 (N_4844,In_839,In_176);
and U4845 (N_4845,In_159,In_1679);
xor U4846 (N_4846,In_2058,In_1264);
nor U4847 (N_4847,In_722,In_1091);
or U4848 (N_4848,In_62,In_1764);
and U4849 (N_4849,In_1886,In_1144);
or U4850 (N_4850,In_711,In_844);
and U4851 (N_4851,In_2149,In_2442);
and U4852 (N_4852,In_86,In_2044);
nand U4853 (N_4853,In_2083,In_1503);
nor U4854 (N_4854,In_1222,In_817);
nor U4855 (N_4855,In_2136,In_2444);
or U4856 (N_4856,In_1026,In_1352);
nor U4857 (N_4857,In_206,In_2092);
nand U4858 (N_4858,In_418,In_2290);
xor U4859 (N_4859,In_2016,In_378);
xor U4860 (N_4860,In_1193,In_2071);
or U4861 (N_4861,In_2261,In_2373);
and U4862 (N_4862,In_2145,In_461);
and U4863 (N_4863,In_1255,In_2405);
or U4864 (N_4864,In_594,In_2186);
xor U4865 (N_4865,In_352,In_2426);
and U4866 (N_4866,In_1046,In_163);
nor U4867 (N_4867,In_2009,In_1285);
nand U4868 (N_4868,In_1051,In_1525);
and U4869 (N_4869,In_1906,In_1248);
nor U4870 (N_4870,In_340,In_726);
nand U4871 (N_4871,In_1867,In_150);
xnor U4872 (N_4872,In_1772,In_74);
nand U4873 (N_4873,In_425,In_1838);
nor U4874 (N_4874,In_1555,In_1768);
and U4875 (N_4875,In_1057,In_1862);
xor U4876 (N_4876,In_572,In_2479);
or U4877 (N_4877,In_1824,In_429);
nand U4878 (N_4878,In_579,In_2232);
nor U4879 (N_4879,In_913,In_2416);
nor U4880 (N_4880,In_1852,In_929);
and U4881 (N_4881,In_684,In_112);
and U4882 (N_4882,In_69,In_1784);
nand U4883 (N_4883,In_1849,In_2189);
nor U4884 (N_4884,In_1485,In_526);
xor U4885 (N_4885,In_445,In_1439);
and U4886 (N_4886,In_997,In_1755);
and U4887 (N_4887,In_815,In_1898);
or U4888 (N_4888,In_2393,In_1755);
and U4889 (N_4889,In_781,In_1632);
nor U4890 (N_4890,In_301,In_124);
and U4891 (N_4891,In_2384,In_1223);
nand U4892 (N_4892,In_1846,In_1396);
nor U4893 (N_4893,In_1722,In_1074);
nand U4894 (N_4894,In_824,In_1325);
or U4895 (N_4895,In_2128,In_1155);
and U4896 (N_4896,In_1000,In_494);
and U4897 (N_4897,In_1326,In_71);
nor U4898 (N_4898,In_954,In_1381);
and U4899 (N_4899,In_1246,In_2031);
and U4900 (N_4900,In_644,In_48);
nor U4901 (N_4901,In_1892,In_1438);
xor U4902 (N_4902,In_1507,In_2314);
or U4903 (N_4903,In_21,In_1232);
nand U4904 (N_4904,In_234,In_327);
or U4905 (N_4905,In_523,In_1554);
nor U4906 (N_4906,In_1061,In_990);
nor U4907 (N_4907,In_411,In_2164);
nor U4908 (N_4908,In_582,In_1661);
nor U4909 (N_4909,In_2072,In_1144);
or U4910 (N_4910,In_875,In_1618);
and U4911 (N_4911,In_1857,In_427);
or U4912 (N_4912,In_48,In_2038);
nor U4913 (N_4913,In_1665,In_1682);
nand U4914 (N_4914,In_219,In_913);
and U4915 (N_4915,In_1304,In_2240);
and U4916 (N_4916,In_1347,In_365);
nand U4917 (N_4917,In_572,In_1452);
nand U4918 (N_4918,In_1562,In_1067);
or U4919 (N_4919,In_12,In_1556);
nand U4920 (N_4920,In_1877,In_2315);
nand U4921 (N_4921,In_1321,In_775);
and U4922 (N_4922,In_45,In_561);
or U4923 (N_4923,In_1861,In_989);
and U4924 (N_4924,In_1836,In_390);
and U4925 (N_4925,In_1805,In_1234);
and U4926 (N_4926,In_709,In_2187);
nor U4927 (N_4927,In_2474,In_1468);
nand U4928 (N_4928,In_1007,In_974);
xnor U4929 (N_4929,In_1446,In_1036);
and U4930 (N_4930,In_1576,In_1742);
nor U4931 (N_4931,In_1229,In_873);
nand U4932 (N_4932,In_780,In_1506);
or U4933 (N_4933,In_2489,In_372);
and U4934 (N_4934,In_1086,In_310);
nor U4935 (N_4935,In_2349,In_1232);
nand U4936 (N_4936,In_905,In_486);
or U4937 (N_4937,In_1934,In_2141);
or U4938 (N_4938,In_1951,In_1857);
xnor U4939 (N_4939,In_1396,In_686);
nor U4940 (N_4940,In_1128,In_938);
nor U4941 (N_4941,In_2091,In_162);
and U4942 (N_4942,In_480,In_1077);
nand U4943 (N_4943,In_1268,In_2434);
nand U4944 (N_4944,In_1312,In_2405);
nor U4945 (N_4945,In_2023,In_1089);
and U4946 (N_4946,In_657,In_614);
nor U4947 (N_4947,In_2180,In_2436);
nor U4948 (N_4948,In_2059,In_28);
nor U4949 (N_4949,In_1281,In_632);
xor U4950 (N_4950,In_587,In_21);
xnor U4951 (N_4951,In_1007,In_2335);
nor U4952 (N_4952,In_1179,In_591);
or U4953 (N_4953,In_1232,In_1180);
nor U4954 (N_4954,In_2182,In_163);
and U4955 (N_4955,In_1957,In_1007);
nor U4956 (N_4956,In_2406,In_2480);
or U4957 (N_4957,In_858,In_1901);
xnor U4958 (N_4958,In_356,In_2386);
nand U4959 (N_4959,In_855,In_798);
nor U4960 (N_4960,In_156,In_1655);
nand U4961 (N_4961,In_1920,In_604);
xor U4962 (N_4962,In_645,In_1804);
nand U4963 (N_4963,In_2308,In_2469);
or U4964 (N_4964,In_273,In_1541);
or U4965 (N_4965,In_1491,In_1065);
nor U4966 (N_4966,In_233,In_2058);
or U4967 (N_4967,In_672,In_1521);
nand U4968 (N_4968,In_238,In_1303);
xnor U4969 (N_4969,In_1504,In_606);
nor U4970 (N_4970,In_46,In_434);
nand U4971 (N_4971,In_1724,In_2164);
or U4972 (N_4972,In_1222,In_37);
nor U4973 (N_4973,In_1818,In_134);
or U4974 (N_4974,In_1630,In_1434);
nor U4975 (N_4975,In_1489,In_275);
xor U4976 (N_4976,In_2319,In_2308);
and U4977 (N_4977,In_521,In_653);
nand U4978 (N_4978,In_38,In_1519);
nand U4979 (N_4979,In_129,In_1632);
nor U4980 (N_4980,In_201,In_1362);
or U4981 (N_4981,In_794,In_2165);
nand U4982 (N_4982,In_306,In_1288);
or U4983 (N_4983,In_1105,In_1075);
nand U4984 (N_4984,In_364,In_1193);
or U4985 (N_4985,In_525,In_45);
and U4986 (N_4986,In_1572,In_380);
xnor U4987 (N_4987,In_1931,In_326);
xnor U4988 (N_4988,In_308,In_562);
nand U4989 (N_4989,In_1409,In_1179);
and U4990 (N_4990,In_1445,In_2166);
nor U4991 (N_4991,In_927,In_2117);
or U4992 (N_4992,In_1296,In_2422);
nor U4993 (N_4993,In_905,In_304);
or U4994 (N_4994,In_148,In_175);
nor U4995 (N_4995,In_2024,In_160);
nand U4996 (N_4996,In_250,In_1048);
nor U4997 (N_4997,In_2248,In_33);
nand U4998 (N_4998,In_634,In_994);
nor U4999 (N_4999,In_1235,In_1908);
or U5000 (N_5000,In_2494,In_2152);
or U5001 (N_5001,In_63,In_1943);
nor U5002 (N_5002,In_2406,In_1366);
and U5003 (N_5003,In_1506,In_2294);
or U5004 (N_5004,In_331,In_1480);
and U5005 (N_5005,In_871,In_57);
and U5006 (N_5006,In_1275,In_1898);
nand U5007 (N_5007,In_1163,In_3);
and U5008 (N_5008,In_1005,In_1901);
or U5009 (N_5009,In_1651,In_636);
nor U5010 (N_5010,In_843,In_847);
nor U5011 (N_5011,In_209,In_815);
and U5012 (N_5012,In_978,In_2404);
or U5013 (N_5013,In_1205,In_2025);
nor U5014 (N_5014,In_405,In_1444);
or U5015 (N_5015,In_1504,In_1990);
nor U5016 (N_5016,In_1451,In_2070);
nor U5017 (N_5017,In_1093,In_2191);
xnor U5018 (N_5018,In_261,In_2424);
nor U5019 (N_5019,In_1442,In_1361);
and U5020 (N_5020,In_1585,In_1929);
nand U5021 (N_5021,In_131,In_287);
or U5022 (N_5022,In_1457,In_253);
nand U5023 (N_5023,In_676,In_1469);
or U5024 (N_5024,In_1278,In_371);
nor U5025 (N_5025,In_247,In_296);
nor U5026 (N_5026,In_171,In_2367);
nand U5027 (N_5027,In_803,In_12);
nand U5028 (N_5028,In_2038,In_41);
or U5029 (N_5029,In_2147,In_2463);
and U5030 (N_5030,In_503,In_1358);
nor U5031 (N_5031,In_135,In_2085);
nand U5032 (N_5032,In_1883,In_1062);
and U5033 (N_5033,In_1374,In_2211);
nor U5034 (N_5034,In_831,In_2299);
nand U5035 (N_5035,In_1971,In_1232);
nand U5036 (N_5036,In_1133,In_73);
nor U5037 (N_5037,In_303,In_1080);
or U5038 (N_5038,In_963,In_649);
and U5039 (N_5039,In_468,In_1070);
nand U5040 (N_5040,In_1188,In_491);
xor U5041 (N_5041,In_2414,In_1110);
or U5042 (N_5042,In_692,In_726);
nor U5043 (N_5043,In_1224,In_713);
or U5044 (N_5044,In_921,In_502);
and U5045 (N_5045,In_2452,In_1805);
nand U5046 (N_5046,In_1662,In_509);
or U5047 (N_5047,In_381,In_484);
or U5048 (N_5048,In_2273,In_1363);
nor U5049 (N_5049,In_986,In_964);
and U5050 (N_5050,In_2251,In_34);
nand U5051 (N_5051,In_545,In_2135);
nor U5052 (N_5052,In_910,In_2053);
and U5053 (N_5053,In_490,In_1930);
nand U5054 (N_5054,In_460,In_856);
nor U5055 (N_5055,In_1129,In_749);
xnor U5056 (N_5056,In_1217,In_1386);
xor U5057 (N_5057,In_1893,In_1609);
nand U5058 (N_5058,In_1208,In_1980);
and U5059 (N_5059,In_1859,In_308);
and U5060 (N_5060,In_276,In_421);
nand U5061 (N_5061,In_901,In_818);
and U5062 (N_5062,In_1119,In_132);
nand U5063 (N_5063,In_603,In_980);
xor U5064 (N_5064,In_1633,In_943);
and U5065 (N_5065,In_566,In_557);
or U5066 (N_5066,In_2195,In_925);
or U5067 (N_5067,In_1421,In_1076);
or U5068 (N_5068,In_2371,In_1772);
or U5069 (N_5069,In_1162,In_2495);
nor U5070 (N_5070,In_2363,In_1956);
and U5071 (N_5071,In_209,In_1451);
and U5072 (N_5072,In_640,In_33);
and U5073 (N_5073,In_316,In_48);
or U5074 (N_5074,In_1408,In_1095);
or U5075 (N_5075,In_1430,In_585);
xor U5076 (N_5076,In_508,In_1941);
nor U5077 (N_5077,In_2106,In_823);
and U5078 (N_5078,In_2181,In_1931);
and U5079 (N_5079,In_503,In_2065);
nor U5080 (N_5080,In_1636,In_1790);
or U5081 (N_5081,In_1177,In_328);
or U5082 (N_5082,In_2478,In_2375);
xor U5083 (N_5083,In_831,In_1353);
nand U5084 (N_5084,In_4,In_2389);
and U5085 (N_5085,In_1109,In_400);
nand U5086 (N_5086,In_147,In_1972);
or U5087 (N_5087,In_1701,In_90);
nand U5088 (N_5088,In_1960,In_2124);
or U5089 (N_5089,In_679,In_1557);
nor U5090 (N_5090,In_583,In_1733);
and U5091 (N_5091,In_558,In_2318);
nor U5092 (N_5092,In_2429,In_673);
and U5093 (N_5093,In_960,In_1708);
and U5094 (N_5094,In_1537,In_835);
nor U5095 (N_5095,In_1813,In_500);
and U5096 (N_5096,In_1702,In_1120);
and U5097 (N_5097,In_508,In_1957);
nand U5098 (N_5098,In_2012,In_80);
or U5099 (N_5099,In_148,In_1151);
xor U5100 (N_5100,In_614,In_1921);
xor U5101 (N_5101,In_2162,In_384);
nand U5102 (N_5102,In_1438,In_455);
nand U5103 (N_5103,In_123,In_1690);
nor U5104 (N_5104,In_722,In_2156);
xor U5105 (N_5105,In_1758,In_1726);
or U5106 (N_5106,In_1571,In_1222);
and U5107 (N_5107,In_1965,In_1332);
nand U5108 (N_5108,In_1218,In_211);
nand U5109 (N_5109,In_74,In_2054);
or U5110 (N_5110,In_1010,In_1295);
nor U5111 (N_5111,In_698,In_2200);
or U5112 (N_5112,In_815,In_1633);
or U5113 (N_5113,In_2142,In_2151);
xor U5114 (N_5114,In_717,In_2499);
nand U5115 (N_5115,In_892,In_1936);
nand U5116 (N_5116,In_379,In_2140);
nor U5117 (N_5117,In_630,In_1739);
nand U5118 (N_5118,In_591,In_1073);
nand U5119 (N_5119,In_837,In_1429);
and U5120 (N_5120,In_2394,In_1594);
or U5121 (N_5121,In_817,In_2238);
nand U5122 (N_5122,In_1061,In_1744);
xnor U5123 (N_5123,In_1936,In_782);
or U5124 (N_5124,In_52,In_2388);
and U5125 (N_5125,In_1239,In_724);
and U5126 (N_5126,In_1854,In_2075);
and U5127 (N_5127,In_2248,In_2246);
nand U5128 (N_5128,In_369,In_231);
and U5129 (N_5129,In_1024,In_1480);
or U5130 (N_5130,In_131,In_1906);
and U5131 (N_5131,In_1789,In_1190);
nand U5132 (N_5132,In_68,In_636);
nand U5133 (N_5133,In_1871,In_23);
or U5134 (N_5134,In_127,In_978);
and U5135 (N_5135,In_1142,In_588);
xnor U5136 (N_5136,In_189,In_204);
and U5137 (N_5137,In_1260,In_1306);
or U5138 (N_5138,In_420,In_2200);
xor U5139 (N_5139,In_2246,In_1886);
nor U5140 (N_5140,In_1152,In_506);
and U5141 (N_5141,In_1173,In_689);
nor U5142 (N_5142,In_1237,In_448);
nand U5143 (N_5143,In_1128,In_1707);
and U5144 (N_5144,In_934,In_2308);
or U5145 (N_5145,In_1700,In_2314);
and U5146 (N_5146,In_1133,In_2046);
xor U5147 (N_5147,In_40,In_816);
and U5148 (N_5148,In_606,In_1656);
and U5149 (N_5149,In_2,In_218);
or U5150 (N_5150,In_1026,In_200);
and U5151 (N_5151,In_1741,In_437);
and U5152 (N_5152,In_480,In_855);
nand U5153 (N_5153,In_2317,In_2355);
or U5154 (N_5154,In_229,In_1494);
nor U5155 (N_5155,In_2314,In_1740);
and U5156 (N_5156,In_678,In_1162);
xnor U5157 (N_5157,In_1331,In_1697);
nand U5158 (N_5158,In_160,In_758);
and U5159 (N_5159,In_1837,In_1916);
or U5160 (N_5160,In_2122,In_2385);
nand U5161 (N_5161,In_241,In_1922);
and U5162 (N_5162,In_873,In_1301);
nor U5163 (N_5163,In_414,In_996);
nor U5164 (N_5164,In_1270,In_2439);
nand U5165 (N_5165,In_2011,In_510);
nand U5166 (N_5166,In_1411,In_221);
and U5167 (N_5167,In_1958,In_1898);
nand U5168 (N_5168,In_1757,In_1701);
nor U5169 (N_5169,In_132,In_1817);
nor U5170 (N_5170,In_100,In_577);
and U5171 (N_5171,In_1075,In_2032);
nand U5172 (N_5172,In_2107,In_1307);
and U5173 (N_5173,In_1996,In_1671);
and U5174 (N_5174,In_1321,In_99);
nand U5175 (N_5175,In_1842,In_2069);
nor U5176 (N_5176,In_206,In_1268);
or U5177 (N_5177,In_916,In_1999);
or U5178 (N_5178,In_1571,In_265);
or U5179 (N_5179,In_724,In_309);
nand U5180 (N_5180,In_1988,In_1715);
or U5181 (N_5181,In_2335,In_2065);
nor U5182 (N_5182,In_815,In_1721);
nor U5183 (N_5183,In_854,In_1955);
nand U5184 (N_5184,In_122,In_1136);
xnor U5185 (N_5185,In_1993,In_2014);
or U5186 (N_5186,In_2380,In_1213);
nand U5187 (N_5187,In_841,In_360);
or U5188 (N_5188,In_748,In_454);
xor U5189 (N_5189,In_2391,In_2156);
and U5190 (N_5190,In_722,In_236);
nor U5191 (N_5191,In_1360,In_192);
and U5192 (N_5192,In_1899,In_915);
or U5193 (N_5193,In_2316,In_2134);
and U5194 (N_5194,In_2290,In_755);
and U5195 (N_5195,In_1342,In_142);
xnor U5196 (N_5196,In_2338,In_1663);
and U5197 (N_5197,In_107,In_853);
xor U5198 (N_5198,In_2075,In_358);
or U5199 (N_5199,In_1790,In_469);
xor U5200 (N_5200,In_332,In_1621);
nand U5201 (N_5201,In_1040,In_1307);
or U5202 (N_5202,In_2462,In_1617);
or U5203 (N_5203,In_558,In_1553);
xor U5204 (N_5204,In_2137,In_1758);
and U5205 (N_5205,In_437,In_846);
xnor U5206 (N_5206,In_793,In_1762);
nand U5207 (N_5207,In_258,In_1688);
xnor U5208 (N_5208,In_1181,In_414);
and U5209 (N_5209,In_565,In_1045);
nor U5210 (N_5210,In_1454,In_806);
nand U5211 (N_5211,In_191,In_384);
or U5212 (N_5212,In_1518,In_1436);
and U5213 (N_5213,In_484,In_1707);
xor U5214 (N_5214,In_1398,In_1446);
nand U5215 (N_5215,In_710,In_540);
nor U5216 (N_5216,In_1345,In_28);
and U5217 (N_5217,In_23,In_1412);
nand U5218 (N_5218,In_1961,In_1401);
nor U5219 (N_5219,In_329,In_2280);
nand U5220 (N_5220,In_2251,In_2137);
nor U5221 (N_5221,In_977,In_2494);
nor U5222 (N_5222,In_765,In_294);
or U5223 (N_5223,In_463,In_1959);
and U5224 (N_5224,In_1697,In_307);
nor U5225 (N_5225,In_685,In_2008);
nand U5226 (N_5226,In_1485,In_450);
or U5227 (N_5227,In_260,In_160);
or U5228 (N_5228,In_108,In_2477);
nor U5229 (N_5229,In_681,In_217);
nor U5230 (N_5230,In_1832,In_162);
nor U5231 (N_5231,In_1719,In_1460);
or U5232 (N_5232,In_561,In_833);
nand U5233 (N_5233,In_499,In_2107);
or U5234 (N_5234,In_447,In_600);
and U5235 (N_5235,In_1352,In_577);
nand U5236 (N_5236,In_2219,In_761);
nor U5237 (N_5237,In_1217,In_1448);
xor U5238 (N_5238,In_2087,In_949);
xnor U5239 (N_5239,In_583,In_2325);
xor U5240 (N_5240,In_1695,In_1270);
nand U5241 (N_5241,In_1379,In_1305);
nor U5242 (N_5242,In_1080,In_60);
nor U5243 (N_5243,In_249,In_94);
nand U5244 (N_5244,In_2367,In_760);
nor U5245 (N_5245,In_1974,In_1209);
or U5246 (N_5246,In_1652,In_54);
and U5247 (N_5247,In_2274,In_1989);
nor U5248 (N_5248,In_354,In_1665);
and U5249 (N_5249,In_150,In_2484);
nand U5250 (N_5250,In_913,In_1041);
nor U5251 (N_5251,In_2395,In_1093);
nand U5252 (N_5252,In_2281,In_770);
nor U5253 (N_5253,In_2209,In_2144);
and U5254 (N_5254,In_1627,In_2179);
xnor U5255 (N_5255,In_622,In_466);
and U5256 (N_5256,In_211,In_1443);
nand U5257 (N_5257,In_1817,In_436);
nor U5258 (N_5258,In_890,In_2368);
nor U5259 (N_5259,In_1790,In_1454);
nor U5260 (N_5260,In_1772,In_534);
or U5261 (N_5261,In_515,In_2469);
nor U5262 (N_5262,In_1491,In_156);
nor U5263 (N_5263,In_2182,In_2186);
nand U5264 (N_5264,In_639,In_491);
or U5265 (N_5265,In_1206,In_847);
or U5266 (N_5266,In_1657,In_996);
and U5267 (N_5267,In_1467,In_1811);
and U5268 (N_5268,In_615,In_1135);
nor U5269 (N_5269,In_1842,In_1043);
nor U5270 (N_5270,In_320,In_1827);
nand U5271 (N_5271,In_106,In_2288);
or U5272 (N_5272,In_1827,In_930);
and U5273 (N_5273,In_2361,In_413);
or U5274 (N_5274,In_209,In_1457);
nand U5275 (N_5275,In_2071,In_717);
nor U5276 (N_5276,In_1268,In_1591);
or U5277 (N_5277,In_748,In_785);
nand U5278 (N_5278,In_2489,In_1103);
nor U5279 (N_5279,In_992,In_1622);
or U5280 (N_5280,In_1606,In_776);
nand U5281 (N_5281,In_461,In_545);
and U5282 (N_5282,In_1297,In_188);
or U5283 (N_5283,In_1196,In_1295);
and U5284 (N_5284,In_1805,In_661);
nand U5285 (N_5285,In_1157,In_136);
nor U5286 (N_5286,In_770,In_2363);
and U5287 (N_5287,In_1022,In_2282);
and U5288 (N_5288,In_1743,In_1539);
or U5289 (N_5289,In_1147,In_1108);
nand U5290 (N_5290,In_569,In_1758);
or U5291 (N_5291,In_310,In_1764);
or U5292 (N_5292,In_1712,In_15);
nand U5293 (N_5293,In_1328,In_216);
or U5294 (N_5294,In_314,In_867);
nand U5295 (N_5295,In_2071,In_1256);
and U5296 (N_5296,In_393,In_410);
and U5297 (N_5297,In_1431,In_2240);
or U5298 (N_5298,In_1198,In_746);
nor U5299 (N_5299,In_1226,In_947);
and U5300 (N_5300,In_1476,In_983);
and U5301 (N_5301,In_2419,In_1847);
nand U5302 (N_5302,In_182,In_2272);
and U5303 (N_5303,In_412,In_1998);
nor U5304 (N_5304,In_641,In_356);
nand U5305 (N_5305,In_2224,In_371);
nand U5306 (N_5306,In_1811,In_1132);
and U5307 (N_5307,In_1408,In_1309);
nand U5308 (N_5308,In_56,In_2179);
nor U5309 (N_5309,In_298,In_2109);
or U5310 (N_5310,In_1146,In_1222);
nand U5311 (N_5311,In_397,In_1915);
nand U5312 (N_5312,In_248,In_872);
or U5313 (N_5313,In_689,In_2230);
and U5314 (N_5314,In_1692,In_2499);
xnor U5315 (N_5315,In_2341,In_722);
or U5316 (N_5316,In_262,In_2135);
nand U5317 (N_5317,In_2141,In_774);
nand U5318 (N_5318,In_2325,In_1489);
and U5319 (N_5319,In_1702,In_234);
nand U5320 (N_5320,In_426,In_1399);
and U5321 (N_5321,In_1675,In_2090);
nor U5322 (N_5322,In_285,In_1694);
nand U5323 (N_5323,In_880,In_722);
and U5324 (N_5324,In_39,In_1877);
nor U5325 (N_5325,In_191,In_1870);
nand U5326 (N_5326,In_820,In_29);
nor U5327 (N_5327,In_508,In_2483);
xor U5328 (N_5328,In_1570,In_1788);
or U5329 (N_5329,In_2042,In_2283);
xor U5330 (N_5330,In_1591,In_2143);
nand U5331 (N_5331,In_939,In_578);
nor U5332 (N_5332,In_2195,In_1860);
and U5333 (N_5333,In_1308,In_1330);
and U5334 (N_5334,In_1780,In_1409);
and U5335 (N_5335,In_1309,In_2292);
or U5336 (N_5336,In_1822,In_2451);
nand U5337 (N_5337,In_1553,In_908);
nand U5338 (N_5338,In_2117,In_1236);
and U5339 (N_5339,In_1758,In_1419);
nand U5340 (N_5340,In_850,In_1262);
nand U5341 (N_5341,In_626,In_330);
nand U5342 (N_5342,In_147,In_1038);
and U5343 (N_5343,In_2471,In_1826);
and U5344 (N_5344,In_315,In_1860);
and U5345 (N_5345,In_1033,In_557);
or U5346 (N_5346,In_1099,In_1943);
nand U5347 (N_5347,In_1279,In_561);
nand U5348 (N_5348,In_1717,In_929);
or U5349 (N_5349,In_438,In_911);
or U5350 (N_5350,In_2336,In_873);
nand U5351 (N_5351,In_196,In_2214);
nor U5352 (N_5352,In_936,In_127);
nor U5353 (N_5353,In_1664,In_2042);
and U5354 (N_5354,In_1656,In_391);
and U5355 (N_5355,In_921,In_555);
nand U5356 (N_5356,In_553,In_2269);
and U5357 (N_5357,In_1261,In_1548);
nor U5358 (N_5358,In_2332,In_2475);
or U5359 (N_5359,In_1957,In_2047);
and U5360 (N_5360,In_2334,In_796);
xor U5361 (N_5361,In_521,In_2045);
xnor U5362 (N_5362,In_1201,In_38);
xor U5363 (N_5363,In_1872,In_38);
and U5364 (N_5364,In_2387,In_3);
or U5365 (N_5365,In_1122,In_1836);
nor U5366 (N_5366,In_537,In_212);
xor U5367 (N_5367,In_331,In_1035);
nor U5368 (N_5368,In_1106,In_1631);
nor U5369 (N_5369,In_2323,In_1766);
or U5370 (N_5370,In_121,In_1881);
nand U5371 (N_5371,In_1658,In_301);
nand U5372 (N_5372,In_1350,In_207);
or U5373 (N_5373,In_2020,In_768);
nor U5374 (N_5374,In_431,In_653);
or U5375 (N_5375,In_1803,In_97);
and U5376 (N_5376,In_2472,In_1743);
nor U5377 (N_5377,In_1661,In_1557);
nand U5378 (N_5378,In_1234,In_2199);
nor U5379 (N_5379,In_1631,In_2225);
and U5380 (N_5380,In_778,In_463);
xnor U5381 (N_5381,In_1872,In_752);
nand U5382 (N_5382,In_783,In_512);
and U5383 (N_5383,In_1864,In_327);
and U5384 (N_5384,In_206,In_745);
nor U5385 (N_5385,In_615,In_2228);
xor U5386 (N_5386,In_46,In_2172);
xor U5387 (N_5387,In_1463,In_938);
nor U5388 (N_5388,In_2109,In_1713);
nor U5389 (N_5389,In_2029,In_1359);
or U5390 (N_5390,In_2170,In_1393);
xnor U5391 (N_5391,In_710,In_1734);
and U5392 (N_5392,In_1648,In_712);
nand U5393 (N_5393,In_522,In_448);
nand U5394 (N_5394,In_969,In_1844);
nor U5395 (N_5395,In_2384,In_1934);
and U5396 (N_5396,In_800,In_1890);
nor U5397 (N_5397,In_1194,In_1607);
nor U5398 (N_5398,In_2407,In_1548);
and U5399 (N_5399,In_526,In_1148);
and U5400 (N_5400,In_1025,In_217);
nand U5401 (N_5401,In_27,In_2475);
nor U5402 (N_5402,In_2302,In_1446);
nand U5403 (N_5403,In_1586,In_1187);
xor U5404 (N_5404,In_125,In_88);
and U5405 (N_5405,In_1695,In_774);
and U5406 (N_5406,In_1935,In_504);
or U5407 (N_5407,In_926,In_292);
nor U5408 (N_5408,In_1212,In_33);
nor U5409 (N_5409,In_1010,In_1335);
nand U5410 (N_5410,In_1283,In_113);
xnor U5411 (N_5411,In_893,In_2167);
nor U5412 (N_5412,In_2432,In_1267);
nor U5413 (N_5413,In_528,In_452);
or U5414 (N_5414,In_1235,In_2255);
and U5415 (N_5415,In_2316,In_1131);
nor U5416 (N_5416,In_1224,In_711);
nor U5417 (N_5417,In_2386,In_2376);
and U5418 (N_5418,In_1043,In_35);
nor U5419 (N_5419,In_1128,In_2465);
nand U5420 (N_5420,In_1278,In_146);
nor U5421 (N_5421,In_2359,In_1407);
and U5422 (N_5422,In_527,In_729);
nor U5423 (N_5423,In_1947,In_1336);
xor U5424 (N_5424,In_1010,In_1022);
and U5425 (N_5425,In_1798,In_379);
xnor U5426 (N_5426,In_1181,In_1118);
nor U5427 (N_5427,In_2264,In_126);
or U5428 (N_5428,In_1195,In_712);
and U5429 (N_5429,In_2130,In_451);
and U5430 (N_5430,In_69,In_2498);
and U5431 (N_5431,In_22,In_244);
or U5432 (N_5432,In_2148,In_338);
and U5433 (N_5433,In_2343,In_1435);
and U5434 (N_5434,In_1015,In_657);
and U5435 (N_5435,In_188,In_1043);
or U5436 (N_5436,In_1781,In_66);
xnor U5437 (N_5437,In_52,In_1586);
and U5438 (N_5438,In_952,In_1740);
and U5439 (N_5439,In_581,In_1041);
nor U5440 (N_5440,In_878,In_1384);
nand U5441 (N_5441,In_2084,In_353);
nor U5442 (N_5442,In_711,In_1178);
nand U5443 (N_5443,In_1957,In_820);
and U5444 (N_5444,In_2349,In_593);
nor U5445 (N_5445,In_136,In_2001);
nor U5446 (N_5446,In_2008,In_1733);
or U5447 (N_5447,In_574,In_93);
nand U5448 (N_5448,In_1529,In_2415);
xor U5449 (N_5449,In_1033,In_1641);
nor U5450 (N_5450,In_1787,In_1720);
nand U5451 (N_5451,In_1491,In_859);
nand U5452 (N_5452,In_382,In_367);
nand U5453 (N_5453,In_1995,In_528);
nand U5454 (N_5454,In_1583,In_1890);
and U5455 (N_5455,In_733,In_1274);
and U5456 (N_5456,In_2485,In_1840);
or U5457 (N_5457,In_740,In_543);
xnor U5458 (N_5458,In_1056,In_271);
and U5459 (N_5459,In_1792,In_712);
nor U5460 (N_5460,In_1957,In_1450);
nor U5461 (N_5461,In_1970,In_2215);
nand U5462 (N_5462,In_2283,In_450);
nor U5463 (N_5463,In_1842,In_581);
or U5464 (N_5464,In_1929,In_249);
nand U5465 (N_5465,In_194,In_1222);
or U5466 (N_5466,In_510,In_2486);
and U5467 (N_5467,In_80,In_182);
nor U5468 (N_5468,In_1052,In_1055);
and U5469 (N_5469,In_1241,In_1995);
xnor U5470 (N_5470,In_887,In_2253);
and U5471 (N_5471,In_1229,In_1802);
and U5472 (N_5472,In_2497,In_1285);
and U5473 (N_5473,In_525,In_1766);
nand U5474 (N_5474,In_98,In_418);
nand U5475 (N_5475,In_1223,In_2241);
nand U5476 (N_5476,In_877,In_1096);
and U5477 (N_5477,In_1582,In_579);
xnor U5478 (N_5478,In_877,In_1501);
nand U5479 (N_5479,In_1655,In_1383);
and U5480 (N_5480,In_1943,In_1873);
and U5481 (N_5481,In_808,In_6);
nand U5482 (N_5482,In_508,In_1602);
nand U5483 (N_5483,In_560,In_1735);
xnor U5484 (N_5484,In_2227,In_2466);
nand U5485 (N_5485,In_1225,In_1987);
and U5486 (N_5486,In_779,In_1811);
and U5487 (N_5487,In_154,In_1605);
nand U5488 (N_5488,In_678,In_746);
nor U5489 (N_5489,In_1791,In_2034);
nand U5490 (N_5490,In_2251,In_785);
nor U5491 (N_5491,In_1554,In_135);
or U5492 (N_5492,In_277,In_2271);
nand U5493 (N_5493,In_2222,In_2329);
nor U5494 (N_5494,In_2402,In_794);
nor U5495 (N_5495,In_2495,In_595);
or U5496 (N_5496,In_1219,In_1264);
nand U5497 (N_5497,In_1572,In_1317);
and U5498 (N_5498,In_1868,In_271);
nand U5499 (N_5499,In_2084,In_1473);
nor U5500 (N_5500,In_2152,In_116);
or U5501 (N_5501,In_1989,In_2393);
nand U5502 (N_5502,In_2260,In_1958);
and U5503 (N_5503,In_1065,In_362);
and U5504 (N_5504,In_231,In_1082);
and U5505 (N_5505,In_1333,In_2024);
nand U5506 (N_5506,In_1413,In_751);
and U5507 (N_5507,In_674,In_1691);
nor U5508 (N_5508,In_436,In_153);
or U5509 (N_5509,In_1954,In_991);
and U5510 (N_5510,In_379,In_141);
or U5511 (N_5511,In_2326,In_1503);
and U5512 (N_5512,In_788,In_507);
xnor U5513 (N_5513,In_79,In_66);
and U5514 (N_5514,In_2346,In_791);
and U5515 (N_5515,In_2383,In_2442);
or U5516 (N_5516,In_1061,In_2048);
or U5517 (N_5517,In_929,In_1606);
xnor U5518 (N_5518,In_2161,In_409);
and U5519 (N_5519,In_7,In_1612);
nand U5520 (N_5520,In_1577,In_99);
xor U5521 (N_5521,In_1579,In_848);
xnor U5522 (N_5522,In_2114,In_961);
nor U5523 (N_5523,In_1063,In_1943);
or U5524 (N_5524,In_643,In_1495);
nand U5525 (N_5525,In_665,In_447);
and U5526 (N_5526,In_28,In_53);
nor U5527 (N_5527,In_117,In_988);
xor U5528 (N_5528,In_1318,In_40);
or U5529 (N_5529,In_2498,In_40);
nand U5530 (N_5530,In_1352,In_1664);
and U5531 (N_5531,In_858,In_2275);
or U5532 (N_5532,In_235,In_2432);
or U5533 (N_5533,In_1508,In_1437);
nand U5534 (N_5534,In_1494,In_4);
nand U5535 (N_5535,In_362,In_1722);
xor U5536 (N_5536,In_1837,In_953);
nand U5537 (N_5537,In_825,In_2171);
nor U5538 (N_5538,In_962,In_450);
nor U5539 (N_5539,In_18,In_2053);
nor U5540 (N_5540,In_1873,In_570);
nand U5541 (N_5541,In_522,In_768);
and U5542 (N_5542,In_848,In_714);
nand U5543 (N_5543,In_1330,In_2365);
or U5544 (N_5544,In_1225,In_1283);
nand U5545 (N_5545,In_1444,In_2302);
nor U5546 (N_5546,In_1104,In_718);
and U5547 (N_5547,In_1856,In_1283);
or U5548 (N_5548,In_2391,In_1102);
and U5549 (N_5549,In_1367,In_194);
nand U5550 (N_5550,In_1635,In_1145);
or U5551 (N_5551,In_1438,In_919);
or U5552 (N_5552,In_2136,In_2350);
xor U5553 (N_5553,In_508,In_779);
and U5554 (N_5554,In_1404,In_916);
or U5555 (N_5555,In_621,In_811);
and U5556 (N_5556,In_2438,In_40);
nand U5557 (N_5557,In_941,In_1707);
or U5558 (N_5558,In_995,In_48);
nor U5559 (N_5559,In_2244,In_2387);
or U5560 (N_5560,In_316,In_1177);
nand U5561 (N_5561,In_1580,In_473);
nor U5562 (N_5562,In_2076,In_2345);
nor U5563 (N_5563,In_925,In_2095);
or U5564 (N_5564,In_1431,In_1935);
and U5565 (N_5565,In_1653,In_1237);
nand U5566 (N_5566,In_380,In_2232);
nand U5567 (N_5567,In_911,In_125);
nand U5568 (N_5568,In_139,In_1600);
and U5569 (N_5569,In_673,In_1382);
nor U5570 (N_5570,In_1965,In_785);
or U5571 (N_5571,In_2034,In_614);
or U5572 (N_5572,In_23,In_1340);
nand U5573 (N_5573,In_2441,In_623);
nand U5574 (N_5574,In_2132,In_208);
and U5575 (N_5575,In_1616,In_1352);
and U5576 (N_5576,In_1894,In_1915);
xor U5577 (N_5577,In_148,In_739);
nor U5578 (N_5578,In_1105,In_164);
and U5579 (N_5579,In_1355,In_54);
or U5580 (N_5580,In_1813,In_1213);
or U5581 (N_5581,In_978,In_1467);
nand U5582 (N_5582,In_1989,In_2310);
and U5583 (N_5583,In_237,In_1780);
nor U5584 (N_5584,In_1832,In_2165);
and U5585 (N_5585,In_1971,In_2107);
xnor U5586 (N_5586,In_263,In_1408);
nor U5587 (N_5587,In_730,In_538);
nand U5588 (N_5588,In_2313,In_6);
and U5589 (N_5589,In_478,In_2257);
xor U5590 (N_5590,In_97,In_1798);
nand U5591 (N_5591,In_325,In_2143);
nand U5592 (N_5592,In_1614,In_802);
nand U5593 (N_5593,In_427,In_2027);
or U5594 (N_5594,In_1881,In_461);
xnor U5595 (N_5595,In_1523,In_275);
nor U5596 (N_5596,In_2247,In_1051);
nor U5597 (N_5597,In_1056,In_2258);
nand U5598 (N_5598,In_413,In_144);
and U5599 (N_5599,In_1440,In_1626);
xnor U5600 (N_5600,In_1957,In_994);
nor U5601 (N_5601,In_491,In_2315);
nand U5602 (N_5602,In_42,In_525);
nor U5603 (N_5603,In_1001,In_199);
nor U5604 (N_5604,In_1484,In_1298);
and U5605 (N_5605,In_1470,In_476);
nor U5606 (N_5606,In_2105,In_688);
nor U5607 (N_5607,In_247,In_1191);
nor U5608 (N_5608,In_1323,In_459);
xor U5609 (N_5609,In_2213,In_25);
and U5610 (N_5610,In_448,In_319);
nand U5611 (N_5611,In_797,In_64);
or U5612 (N_5612,In_2483,In_761);
and U5613 (N_5613,In_44,In_309);
xnor U5614 (N_5614,In_2006,In_1678);
or U5615 (N_5615,In_1114,In_284);
nand U5616 (N_5616,In_1520,In_1577);
nor U5617 (N_5617,In_2345,In_1894);
nor U5618 (N_5618,In_1537,In_973);
nand U5619 (N_5619,In_1057,In_2364);
nor U5620 (N_5620,In_1493,In_628);
nor U5621 (N_5621,In_1470,In_2035);
or U5622 (N_5622,In_1900,In_2022);
nor U5623 (N_5623,In_1966,In_1179);
nand U5624 (N_5624,In_1415,In_211);
xor U5625 (N_5625,In_1005,In_2479);
or U5626 (N_5626,In_2031,In_2069);
nor U5627 (N_5627,In_1439,In_539);
or U5628 (N_5628,In_2153,In_2158);
nor U5629 (N_5629,In_1684,In_1552);
or U5630 (N_5630,In_433,In_1609);
nor U5631 (N_5631,In_1665,In_653);
nand U5632 (N_5632,In_46,In_1459);
nor U5633 (N_5633,In_860,In_2034);
nor U5634 (N_5634,In_782,In_1826);
and U5635 (N_5635,In_1532,In_764);
or U5636 (N_5636,In_1177,In_1033);
nand U5637 (N_5637,In_413,In_1527);
nand U5638 (N_5638,In_1147,In_1415);
nand U5639 (N_5639,In_1049,In_15);
xnor U5640 (N_5640,In_532,In_1861);
or U5641 (N_5641,In_2437,In_1667);
nand U5642 (N_5642,In_2127,In_1898);
or U5643 (N_5643,In_1918,In_558);
or U5644 (N_5644,In_2243,In_1001);
and U5645 (N_5645,In_1373,In_283);
or U5646 (N_5646,In_1057,In_1351);
nor U5647 (N_5647,In_1966,In_2333);
and U5648 (N_5648,In_2393,In_2275);
nand U5649 (N_5649,In_1481,In_2255);
and U5650 (N_5650,In_621,In_1593);
nor U5651 (N_5651,In_765,In_839);
nor U5652 (N_5652,In_1082,In_636);
nor U5653 (N_5653,In_1433,In_2472);
or U5654 (N_5654,In_576,In_1702);
and U5655 (N_5655,In_403,In_1411);
nor U5656 (N_5656,In_1488,In_2108);
or U5657 (N_5657,In_1434,In_689);
or U5658 (N_5658,In_2325,In_369);
and U5659 (N_5659,In_516,In_1595);
nand U5660 (N_5660,In_2378,In_248);
nor U5661 (N_5661,In_97,In_2396);
and U5662 (N_5662,In_1348,In_562);
or U5663 (N_5663,In_2129,In_1405);
nor U5664 (N_5664,In_1716,In_1899);
nand U5665 (N_5665,In_188,In_1644);
or U5666 (N_5666,In_341,In_1261);
and U5667 (N_5667,In_956,In_293);
nand U5668 (N_5668,In_1441,In_1648);
nor U5669 (N_5669,In_1488,In_2359);
and U5670 (N_5670,In_1700,In_1826);
nand U5671 (N_5671,In_575,In_1307);
and U5672 (N_5672,In_714,In_1105);
nor U5673 (N_5673,In_1952,In_2256);
or U5674 (N_5674,In_433,In_2061);
xnor U5675 (N_5675,In_2135,In_158);
and U5676 (N_5676,In_2097,In_1800);
nor U5677 (N_5677,In_352,In_77);
nand U5678 (N_5678,In_130,In_2112);
or U5679 (N_5679,In_1207,In_1232);
nand U5680 (N_5680,In_2451,In_1278);
xnor U5681 (N_5681,In_1034,In_2156);
nor U5682 (N_5682,In_2075,In_1344);
nor U5683 (N_5683,In_1229,In_1797);
and U5684 (N_5684,In_1951,In_1778);
nor U5685 (N_5685,In_648,In_918);
nand U5686 (N_5686,In_758,In_72);
or U5687 (N_5687,In_1561,In_2186);
nor U5688 (N_5688,In_1954,In_96);
or U5689 (N_5689,In_1064,In_1975);
or U5690 (N_5690,In_1991,In_1132);
nand U5691 (N_5691,In_1772,In_1252);
or U5692 (N_5692,In_1131,In_2101);
xnor U5693 (N_5693,In_108,In_2327);
nand U5694 (N_5694,In_726,In_804);
or U5695 (N_5695,In_459,In_2467);
or U5696 (N_5696,In_406,In_2151);
or U5697 (N_5697,In_1095,In_611);
and U5698 (N_5698,In_950,In_1806);
xor U5699 (N_5699,In_932,In_1877);
or U5700 (N_5700,In_1954,In_1098);
nand U5701 (N_5701,In_2385,In_1933);
nor U5702 (N_5702,In_161,In_1190);
nand U5703 (N_5703,In_2081,In_1402);
and U5704 (N_5704,In_617,In_1633);
and U5705 (N_5705,In_1523,In_969);
nand U5706 (N_5706,In_1445,In_2233);
or U5707 (N_5707,In_2128,In_1809);
or U5708 (N_5708,In_983,In_2457);
nor U5709 (N_5709,In_1088,In_131);
or U5710 (N_5710,In_452,In_2273);
nor U5711 (N_5711,In_1851,In_1766);
or U5712 (N_5712,In_632,In_811);
nand U5713 (N_5713,In_1664,In_2119);
or U5714 (N_5714,In_57,In_119);
and U5715 (N_5715,In_127,In_1825);
nand U5716 (N_5716,In_2216,In_47);
or U5717 (N_5717,In_483,In_267);
nor U5718 (N_5718,In_1069,In_1931);
and U5719 (N_5719,In_2161,In_112);
or U5720 (N_5720,In_2172,In_541);
or U5721 (N_5721,In_1663,In_233);
xor U5722 (N_5722,In_74,In_2040);
nor U5723 (N_5723,In_1343,In_2121);
or U5724 (N_5724,In_715,In_2324);
nor U5725 (N_5725,In_416,In_908);
or U5726 (N_5726,In_2090,In_1768);
and U5727 (N_5727,In_2333,In_1011);
nand U5728 (N_5728,In_10,In_91);
and U5729 (N_5729,In_803,In_1871);
or U5730 (N_5730,In_1272,In_1670);
nand U5731 (N_5731,In_481,In_153);
nand U5732 (N_5732,In_1225,In_2127);
nor U5733 (N_5733,In_1589,In_27);
or U5734 (N_5734,In_683,In_278);
or U5735 (N_5735,In_999,In_974);
nand U5736 (N_5736,In_2249,In_367);
nor U5737 (N_5737,In_699,In_108);
and U5738 (N_5738,In_1958,In_1968);
and U5739 (N_5739,In_493,In_2368);
and U5740 (N_5740,In_1167,In_202);
and U5741 (N_5741,In_2370,In_1266);
xnor U5742 (N_5742,In_505,In_1589);
nor U5743 (N_5743,In_321,In_1067);
nand U5744 (N_5744,In_1566,In_224);
or U5745 (N_5745,In_641,In_1286);
xnor U5746 (N_5746,In_695,In_965);
nand U5747 (N_5747,In_436,In_790);
and U5748 (N_5748,In_1142,In_1268);
nor U5749 (N_5749,In_1689,In_314);
nor U5750 (N_5750,In_1087,In_921);
or U5751 (N_5751,In_990,In_787);
and U5752 (N_5752,In_398,In_1854);
and U5753 (N_5753,In_521,In_2387);
or U5754 (N_5754,In_1766,In_1826);
nand U5755 (N_5755,In_2406,In_664);
xnor U5756 (N_5756,In_2473,In_508);
and U5757 (N_5757,In_863,In_705);
nand U5758 (N_5758,In_157,In_2137);
or U5759 (N_5759,In_1431,In_1658);
nor U5760 (N_5760,In_234,In_900);
and U5761 (N_5761,In_941,In_881);
nand U5762 (N_5762,In_1824,In_1606);
xor U5763 (N_5763,In_536,In_1136);
xnor U5764 (N_5764,In_20,In_1333);
nor U5765 (N_5765,In_1515,In_829);
nand U5766 (N_5766,In_3,In_1787);
xor U5767 (N_5767,In_755,In_1549);
xnor U5768 (N_5768,In_294,In_1237);
nor U5769 (N_5769,In_2467,In_1748);
and U5770 (N_5770,In_2047,In_1424);
or U5771 (N_5771,In_465,In_388);
xnor U5772 (N_5772,In_2324,In_1945);
and U5773 (N_5773,In_2464,In_1697);
and U5774 (N_5774,In_1821,In_2112);
xor U5775 (N_5775,In_1731,In_163);
xor U5776 (N_5776,In_71,In_1446);
nor U5777 (N_5777,In_1598,In_710);
nand U5778 (N_5778,In_720,In_1735);
or U5779 (N_5779,In_2119,In_1294);
or U5780 (N_5780,In_2075,In_1079);
nor U5781 (N_5781,In_118,In_2041);
and U5782 (N_5782,In_1587,In_819);
xor U5783 (N_5783,In_213,In_1246);
nand U5784 (N_5784,In_1300,In_1448);
or U5785 (N_5785,In_2413,In_2263);
nand U5786 (N_5786,In_361,In_2485);
and U5787 (N_5787,In_1594,In_1633);
xnor U5788 (N_5788,In_1728,In_673);
or U5789 (N_5789,In_2128,In_246);
nand U5790 (N_5790,In_2287,In_2450);
nor U5791 (N_5791,In_1259,In_96);
nand U5792 (N_5792,In_998,In_629);
nand U5793 (N_5793,In_1997,In_1643);
and U5794 (N_5794,In_721,In_1588);
or U5795 (N_5795,In_542,In_2485);
and U5796 (N_5796,In_825,In_2052);
nor U5797 (N_5797,In_1699,In_2392);
and U5798 (N_5798,In_133,In_1855);
or U5799 (N_5799,In_94,In_1928);
nand U5800 (N_5800,In_585,In_2344);
nand U5801 (N_5801,In_1378,In_1985);
nand U5802 (N_5802,In_2015,In_1307);
and U5803 (N_5803,In_1078,In_290);
nor U5804 (N_5804,In_1336,In_1262);
nand U5805 (N_5805,In_1930,In_245);
nand U5806 (N_5806,In_558,In_2394);
or U5807 (N_5807,In_1673,In_988);
and U5808 (N_5808,In_669,In_11);
nand U5809 (N_5809,In_2216,In_1420);
and U5810 (N_5810,In_652,In_1380);
nand U5811 (N_5811,In_885,In_286);
nor U5812 (N_5812,In_2422,In_1120);
nand U5813 (N_5813,In_1049,In_1466);
and U5814 (N_5814,In_845,In_638);
nor U5815 (N_5815,In_453,In_1400);
nor U5816 (N_5816,In_1013,In_259);
nor U5817 (N_5817,In_669,In_168);
or U5818 (N_5818,In_2358,In_1210);
nand U5819 (N_5819,In_443,In_1693);
and U5820 (N_5820,In_1939,In_1805);
nor U5821 (N_5821,In_753,In_624);
or U5822 (N_5822,In_1391,In_851);
nor U5823 (N_5823,In_942,In_1116);
or U5824 (N_5824,In_1600,In_2491);
or U5825 (N_5825,In_625,In_1405);
or U5826 (N_5826,In_2248,In_1039);
or U5827 (N_5827,In_1982,In_1135);
or U5828 (N_5828,In_359,In_1923);
and U5829 (N_5829,In_894,In_328);
nand U5830 (N_5830,In_242,In_2288);
or U5831 (N_5831,In_190,In_473);
or U5832 (N_5832,In_849,In_1387);
and U5833 (N_5833,In_1850,In_2040);
xnor U5834 (N_5834,In_365,In_398);
nand U5835 (N_5835,In_241,In_97);
nand U5836 (N_5836,In_2357,In_1291);
nor U5837 (N_5837,In_2384,In_1037);
nor U5838 (N_5838,In_2448,In_285);
or U5839 (N_5839,In_513,In_1386);
nand U5840 (N_5840,In_1727,In_2490);
nor U5841 (N_5841,In_1993,In_1970);
xor U5842 (N_5842,In_674,In_2047);
and U5843 (N_5843,In_2154,In_2283);
xnor U5844 (N_5844,In_877,In_85);
xor U5845 (N_5845,In_1062,In_935);
and U5846 (N_5846,In_361,In_1639);
nor U5847 (N_5847,In_448,In_1953);
nand U5848 (N_5848,In_904,In_431);
and U5849 (N_5849,In_2337,In_931);
nor U5850 (N_5850,In_1117,In_2276);
or U5851 (N_5851,In_1297,In_2298);
or U5852 (N_5852,In_2080,In_830);
nand U5853 (N_5853,In_2214,In_1978);
nand U5854 (N_5854,In_879,In_1611);
xnor U5855 (N_5855,In_151,In_2010);
nand U5856 (N_5856,In_949,In_445);
nand U5857 (N_5857,In_1096,In_365);
nor U5858 (N_5858,In_1851,In_1449);
nor U5859 (N_5859,In_840,In_2067);
nor U5860 (N_5860,In_1758,In_870);
and U5861 (N_5861,In_2380,In_584);
or U5862 (N_5862,In_2250,In_399);
nor U5863 (N_5863,In_2107,In_1298);
and U5864 (N_5864,In_1080,In_705);
and U5865 (N_5865,In_1883,In_1607);
and U5866 (N_5866,In_1989,In_1279);
nand U5867 (N_5867,In_2267,In_464);
and U5868 (N_5868,In_1703,In_1182);
nand U5869 (N_5869,In_2247,In_1064);
nor U5870 (N_5870,In_1751,In_254);
xnor U5871 (N_5871,In_149,In_1405);
or U5872 (N_5872,In_1454,In_1735);
nor U5873 (N_5873,In_308,In_2315);
nor U5874 (N_5874,In_1920,In_2386);
nand U5875 (N_5875,In_543,In_1093);
nand U5876 (N_5876,In_884,In_576);
nor U5877 (N_5877,In_1058,In_1492);
or U5878 (N_5878,In_610,In_113);
nand U5879 (N_5879,In_861,In_2207);
xor U5880 (N_5880,In_75,In_431);
and U5881 (N_5881,In_248,In_274);
or U5882 (N_5882,In_1293,In_342);
nor U5883 (N_5883,In_2142,In_1608);
nor U5884 (N_5884,In_2274,In_2130);
nand U5885 (N_5885,In_613,In_1526);
nand U5886 (N_5886,In_1323,In_1165);
nor U5887 (N_5887,In_1239,In_788);
xor U5888 (N_5888,In_2235,In_359);
nand U5889 (N_5889,In_171,In_2275);
and U5890 (N_5890,In_1905,In_899);
nor U5891 (N_5891,In_357,In_1186);
nor U5892 (N_5892,In_1330,In_402);
or U5893 (N_5893,In_1304,In_1777);
nor U5894 (N_5894,In_2062,In_2113);
or U5895 (N_5895,In_1064,In_536);
nand U5896 (N_5896,In_956,In_2409);
nand U5897 (N_5897,In_2016,In_1700);
nor U5898 (N_5898,In_2439,In_2226);
nand U5899 (N_5899,In_1134,In_2150);
nor U5900 (N_5900,In_864,In_1967);
nor U5901 (N_5901,In_2432,In_431);
nand U5902 (N_5902,In_557,In_2010);
nand U5903 (N_5903,In_797,In_837);
and U5904 (N_5904,In_2470,In_1182);
and U5905 (N_5905,In_778,In_2440);
and U5906 (N_5906,In_1799,In_2298);
nor U5907 (N_5907,In_1935,In_1363);
or U5908 (N_5908,In_409,In_1123);
xor U5909 (N_5909,In_1931,In_2016);
or U5910 (N_5910,In_2148,In_278);
nor U5911 (N_5911,In_2083,In_1694);
or U5912 (N_5912,In_1452,In_1556);
or U5913 (N_5913,In_989,In_336);
nand U5914 (N_5914,In_1359,In_2389);
or U5915 (N_5915,In_2090,In_392);
xnor U5916 (N_5916,In_1381,In_947);
or U5917 (N_5917,In_2185,In_1964);
and U5918 (N_5918,In_623,In_2168);
nor U5919 (N_5919,In_144,In_2090);
and U5920 (N_5920,In_100,In_1867);
or U5921 (N_5921,In_688,In_207);
nand U5922 (N_5922,In_1092,In_855);
nor U5923 (N_5923,In_53,In_2109);
and U5924 (N_5924,In_1967,In_2358);
nor U5925 (N_5925,In_2476,In_2432);
and U5926 (N_5926,In_2342,In_1336);
nor U5927 (N_5927,In_1798,In_2019);
nor U5928 (N_5928,In_2198,In_2397);
or U5929 (N_5929,In_2383,In_2425);
or U5930 (N_5930,In_198,In_1775);
or U5931 (N_5931,In_1934,In_1109);
and U5932 (N_5932,In_219,In_1495);
nand U5933 (N_5933,In_575,In_1034);
nor U5934 (N_5934,In_1722,In_1234);
nand U5935 (N_5935,In_2303,In_1541);
or U5936 (N_5936,In_2119,In_1478);
xnor U5937 (N_5937,In_546,In_2293);
and U5938 (N_5938,In_1546,In_2136);
and U5939 (N_5939,In_1509,In_2207);
nand U5940 (N_5940,In_2392,In_605);
nand U5941 (N_5941,In_1789,In_2266);
nor U5942 (N_5942,In_273,In_521);
or U5943 (N_5943,In_2068,In_1730);
or U5944 (N_5944,In_776,In_2141);
nor U5945 (N_5945,In_145,In_397);
nand U5946 (N_5946,In_1909,In_855);
nor U5947 (N_5947,In_1425,In_271);
xor U5948 (N_5948,In_2055,In_2409);
or U5949 (N_5949,In_1182,In_458);
nand U5950 (N_5950,In_2321,In_1664);
nor U5951 (N_5951,In_1902,In_399);
or U5952 (N_5952,In_690,In_1798);
and U5953 (N_5953,In_201,In_2285);
or U5954 (N_5954,In_1640,In_2143);
nor U5955 (N_5955,In_2354,In_1175);
or U5956 (N_5956,In_1357,In_385);
and U5957 (N_5957,In_475,In_1491);
or U5958 (N_5958,In_2410,In_1529);
or U5959 (N_5959,In_2046,In_1251);
and U5960 (N_5960,In_1337,In_477);
nor U5961 (N_5961,In_155,In_1017);
xor U5962 (N_5962,In_322,In_2135);
nor U5963 (N_5963,In_322,In_557);
or U5964 (N_5964,In_164,In_2292);
nor U5965 (N_5965,In_2399,In_341);
or U5966 (N_5966,In_305,In_547);
or U5967 (N_5967,In_1753,In_190);
or U5968 (N_5968,In_1756,In_2486);
nor U5969 (N_5969,In_234,In_910);
nor U5970 (N_5970,In_2329,In_2333);
nor U5971 (N_5971,In_2476,In_1694);
nor U5972 (N_5972,In_431,In_2456);
xor U5973 (N_5973,In_1343,In_635);
nand U5974 (N_5974,In_282,In_575);
or U5975 (N_5975,In_435,In_2309);
and U5976 (N_5976,In_1436,In_324);
and U5977 (N_5977,In_1322,In_366);
xnor U5978 (N_5978,In_2329,In_2315);
or U5979 (N_5979,In_1138,In_96);
nor U5980 (N_5980,In_2245,In_474);
or U5981 (N_5981,In_1582,In_1060);
nand U5982 (N_5982,In_336,In_1272);
and U5983 (N_5983,In_1957,In_1325);
nor U5984 (N_5984,In_1163,In_582);
nand U5985 (N_5985,In_2438,In_1618);
nor U5986 (N_5986,In_935,In_1476);
nand U5987 (N_5987,In_2471,In_1531);
and U5988 (N_5988,In_2411,In_2147);
and U5989 (N_5989,In_1478,In_1515);
or U5990 (N_5990,In_856,In_322);
nor U5991 (N_5991,In_970,In_1270);
or U5992 (N_5992,In_2223,In_416);
nand U5993 (N_5993,In_146,In_2419);
and U5994 (N_5994,In_1183,In_1343);
nand U5995 (N_5995,In_720,In_294);
nor U5996 (N_5996,In_2091,In_1858);
nor U5997 (N_5997,In_2287,In_296);
nor U5998 (N_5998,In_1307,In_1708);
or U5999 (N_5999,In_2042,In_505);
nand U6000 (N_6000,In_1581,In_1800);
nand U6001 (N_6001,In_1591,In_236);
or U6002 (N_6002,In_8,In_2326);
or U6003 (N_6003,In_768,In_611);
and U6004 (N_6004,In_2479,In_2176);
nand U6005 (N_6005,In_1931,In_908);
or U6006 (N_6006,In_1341,In_1427);
nand U6007 (N_6007,In_2084,In_2381);
xor U6008 (N_6008,In_1534,In_2112);
and U6009 (N_6009,In_1419,In_1577);
or U6010 (N_6010,In_1191,In_2039);
or U6011 (N_6011,In_1915,In_1822);
nand U6012 (N_6012,In_1606,In_1058);
and U6013 (N_6013,In_1202,In_631);
nor U6014 (N_6014,In_1502,In_2126);
and U6015 (N_6015,In_2247,In_2361);
and U6016 (N_6016,In_2328,In_2390);
and U6017 (N_6017,In_871,In_2177);
xnor U6018 (N_6018,In_2085,In_707);
and U6019 (N_6019,In_1910,In_1152);
nand U6020 (N_6020,In_890,In_1553);
nand U6021 (N_6021,In_232,In_1649);
nand U6022 (N_6022,In_404,In_1470);
nor U6023 (N_6023,In_1569,In_1620);
nor U6024 (N_6024,In_1994,In_301);
or U6025 (N_6025,In_2154,In_1119);
xnor U6026 (N_6026,In_1246,In_1170);
and U6027 (N_6027,In_379,In_134);
nor U6028 (N_6028,In_2254,In_1385);
nor U6029 (N_6029,In_342,In_1967);
xor U6030 (N_6030,In_1544,In_987);
and U6031 (N_6031,In_2039,In_2416);
xor U6032 (N_6032,In_575,In_499);
and U6033 (N_6033,In_1108,In_2100);
nor U6034 (N_6034,In_2369,In_1994);
and U6035 (N_6035,In_1462,In_2053);
and U6036 (N_6036,In_734,In_902);
and U6037 (N_6037,In_973,In_1405);
xor U6038 (N_6038,In_1753,In_1722);
and U6039 (N_6039,In_2326,In_1588);
or U6040 (N_6040,In_1638,In_1127);
or U6041 (N_6041,In_1585,In_1904);
nand U6042 (N_6042,In_773,In_549);
nand U6043 (N_6043,In_1123,In_1969);
nor U6044 (N_6044,In_1017,In_503);
nand U6045 (N_6045,In_1830,In_2238);
nor U6046 (N_6046,In_113,In_1659);
and U6047 (N_6047,In_847,In_72);
or U6048 (N_6048,In_837,In_1384);
nand U6049 (N_6049,In_1723,In_2050);
nand U6050 (N_6050,In_1881,In_281);
and U6051 (N_6051,In_2388,In_1754);
xor U6052 (N_6052,In_2421,In_2019);
nand U6053 (N_6053,In_2412,In_831);
and U6054 (N_6054,In_1381,In_1929);
nand U6055 (N_6055,In_1853,In_304);
nand U6056 (N_6056,In_1397,In_739);
nand U6057 (N_6057,In_859,In_1017);
xnor U6058 (N_6058,In_934,In_2195);
nor U6059 (N_6059,In_1395,In_2285);
or U6060 (N_6060,In_1941,In_540);
xnor U6061 (N_6061,In_635,In_183);
nand U6062 (N_6062,In_2469,In_2445);
nor U6063 (N_6063,In_595,In_794);
or U6064 (N_6064,In_773,In_579);
or U6065 (N_6065,In_1572,In_165);
and U6066 (N_6066,In_1451,In_1001);
or U6067 (N_6067,In_2009,In_1230);
or U6068 (N_6068,In_1896,In_2240);
or U6069 (N_6069,In_218,In_1611);
xor U6070 (N_6070,In_255,In_1122);
nor U6071 (N_6071,In_1423,In_523);
xnor U6072 (N_6072,In_632,In_1510);
and U6073 (N_6073,In_978,In_132);
nand U6074 (N_6074,In_116,In_1238);
nor U6075 (N_6075,In_2052,In_1209);
xnor U6076 (N_6076,In_1885,In_238);
nor U6077 (N_6077,In_1450,In_2134);
nor U6078 (N_6078,In_401,In_2417);
or U6079 (N_6079,In_1237,In_1018);
or U6080 (N_6080,In_1774,In_2309);
and U6081 (N_6081,In_906,In_10);
and U6082 (N_6082,In_478,In_2325);
xnor U6083 (N_6083,In_1399,In_663);
or U6084 (N_6084,In_910,In_1138);
xor U6085 (N_6085,In_733,In_840);
and U6086 (N_6086,In_522,In_1117);
xor U6087 (N_6087,In_533,In_1934);
nand U6088 (N_6088,In_2238,In_2167);
and U6089 (N_6089,In_129,In_2132);
or U6090 (N_6090,In_1049,In_1215);
nor U6091 (N_6091,In_537,In_315);
xor U6092 (N_6092,In_897,In_1430);
nand U6093 (N_6093,In_303,In_390);
nand U6094 (N_6094,In_215,In_738);
and U6095 (N_6095,In_542,In_725);
or U6096 (N_6096,In_1815,In_1012);
xnor U6097 (N_6097,In_1051,In_1680);
nand U6098 (N_6098,In_421,In_2054);
or U6099 (N_6099,In_1374,In_816);
nor U6100 (N_6100,In_696,In_1270);
nor U6101 (N_6101,In_1451,In_1412);
and U6102 (N_6102,In_2412,In_1542);
and U6103 (N_6103,In_228,In_1818);
nand U6104 (N_6104,In_1480,In_2202);
nor U6105 (N_6105,In_1741,In_997);
or U6106 (N_6106,In_2177,In_923);
and U6107 (N_6107,In_683,In_1111);
nand U6108 (N_6108,In_532,In_2039);
and U6109 (N_6109,In_2090,In_1824);
nand U6110 (N_6110,In_816,In_300);
and U6111 (N_6111,In_2086,In_2304);
nor U6112 (N_6112,In_1646,In_2454);
nand U6113 (N_6113,In_1593,In_586);
and U6114 (N_6114,In_2076,In_2348);
nand U6115 (N_6115,In_1078,In_1205);
xor U6116 (N_6116,In_1334,In_1901);
nor U6117 (N_6117,In_712,In_2302);
and U6118 (N_6118,In_81,In_1745);
and U6119 (N_6119,In_83,In_960);
or U6120 (N_6120,In_1876,In_1453);
nand U6121 (N_6121,In_1675,In_530);
xor U6122 (N_6122,In_514,In_348);
nand U6123 (N_6123,In_1805,In_50);
or U6124 (N_6124,In_1800,In_2038);
nor U6125 (N_6125,In_1593,In_253);
nor U6126 (N_6126,In_860,In_794);
and U6127 (N_6127,In_768,In_614);
nor U6128 (N_6128,In_1424,In_2151);
xor U6129 (N_6129,In_1508,In_205);
nand U6130 (N_6130,In_694,In_1481);
nand U6131 (N_6131,In_520,In_2025);
and U6132 (N_6132,In_414,In_296);
nor U6133 (N_6133,In_2442,In_896);
and U6134 (N_6134,In_1877,In_1153);
nand U6135 (N_6135,In_1053,In_1457);
or U6136 (N_6136,In_265,In_2404);
xor U6137 (N_6137,In_1304,In_1202);
and U6138 (N_6138,In_928,In_398);
nand U6139 (N_6139,In_2435,In_1395);
and U6140 (N_6140,In_2211,In_2189);
nor U6141 (N_6141,In_202,In_1059);
nor U6142 (N_6142,In_1324,In_582);
and U6143 (N_6143,In_1357,In_391);
and U6144 (N_6144,In_474,In_942);
or U6145 (N_6145,In_1727,In_1091);
nor U6146 (N_6146,In_368,In_616);
nor U6147 (N_6147,In_349,In_54);
xor U6148 (N_6148,In_1842,In_2156);
nand U6149 (N_6149,In_2340,In_218);
and U6150 (N_6150,In_838,In_2016);
nand U6151 (N_6151,In_2263,In_25);
nor U6152 (N_6152,In_386,In_747);
or U6153 (N_6153,In_817,In_2048);
nand U6154 (N_6154,In_889,In_1053);
and U6155 (N_6155,In_2125,In_199);
and U6156 (N_6156,In_1288,In_2429);
or U6157 (N_6157,In_355,In_1146);
or U6158 (N_6158,In_1768,In_2029);
nor U6159 (N_6159,In_1694,In_1776);
nor U6160 (N_6160,In_584,In_1725);
or U6161 (N_6161,In_635,In_2255);
nor U6162 (N_6162,In_638,In_584);
and U6163 (N_6163,In_2460,In_1000);
nor U6164 (N_6164,In_1053,In_479);
and U6165 (N_6165,In_1383,In_999);
nor U6166 (N_6166,In_2290,In_1346);
nor U6167 (N_6167,In_2310,In_245);
nand U6168 (N_6168,In_1872,In_1228);
and U6169 (N_6169,In_1521,In_1691);
or U6170 (N_6170,In_2200,In_860);
and U6171 (N_6171,In_978,In_1008);
or U6172 (N_6172,In_2443,In_2050);
and U6173 (N_6173,In_409,In_2019);
xnor U6174 (N_6174,In_2374,In_1064);
and U6175 (N_6175,In_835,In_1784);
nand U6176 (N_6176,In_1360,In_429);
and U6177 (N_6177,In_2294,In_1251);
and U6178 (N_6178,In_2046,In_665);
or U6179 (N_6179,In_1556,In_375);
or U6180 (N_6180,In_970,In_697);
and U6181 (N_6181,In_1564,In_2091);
and U6182 (N_6182,In_2330,In_2440);
nand U6183 (N_6183,In_1848,In_910);
or U6184 (N_6184,In_252,In_948);
or U6185 (N_6185,In_1398,In_7);
xor U6186 (N_6186,In_1595,In_1888);
xor U6187 (N_6187,In_2073,In_1741);
nor U6188 (N_6188,In_2009,In_978);
nor U6189 (N_6189,In_471,In_2119);
nand U6190 (N_6190,In_1595,In_1305);
nor U6191 (N_6191,In_2458,In_1659);
and U6192 (N_6192,In_1856,In_130);
nand U6193 (N_6193,In_1896,In_382);
and U6194 (N_6194,In_1515,In_1721);
nand U6195 (N_6195,In_291,In_910);
nand U6196 (N_6196,In_221,In_584);
or U6197 (N_6197,In_270,In_1217);
or U6198 (N_6198,In_1957,In_882);
xnor U6199 (N_6199,In_2055,In_2402);
or U6200 (N_6200,In_583,In_1671);
nor U6201 (N_6201,In_870,In_2005);
and U6202 (N_6202,In_978,In_536);
and U6203 (N_6203,In_2202,In_1080);
and U6204 (N_6204,In_1414,In_1223);
nor U6205 (N_6205,In_1873,In_212);
and U6206 (N_6206,In_2421,In_506);
nor U6207 (N_6207,In_848,In_297);
or U6208 (N_6208,In_1155,In_58);
or U6209 (N_6209,In_111,In_84);
or U6210 (N_6210,In_2181,In_390);
and U6211 (N_6211,In_855,In_2205);
nor U6212 (N_6212,In_1608,In_2303);
nor U6213 (N_6213,In_389,In_2414);
nor U6214 (N_6214,In_12,In_2171);
or U6215 (N_6215,In_2017,In_621);
or U6216 (N_6216,In_563,In_205);
nor U6217 (N_6217,In_426,In_970);
and U6218 (N_6218,In_2288,In_692);
nor U6219 (N_6219,In_1743,In_403);
nor U6220 (N_6220,In_961,In_1318);
and U6221 (N_6221,In_1393,In_882);
nor U6222 (N_6222,In_2482,In_1010);
nand U6223 (N_6223,In_702,In_900);
nor U6224 (N_6224,In_935,In_1152);
and U6225 (N_6225,In_1398,In_2209);
and U6226 (N_6226,In_80,In_2456);
or U6227 (N_6227,In_500,In_1238);
xor U6228 (N_6228,In_2445,In_156);
nor U6229 (N_6229,In_1443,In_1732);
xor U6230 (N_6230,In_2409,In_235);
nand U6231 (N_6231,In_2315,In_1916);
nand U6232 (N_6232,In_27,In_1031);
and U6233 (N_6233,In_2292,In_1472);
nand U6234 (N_6234,In_126,In_1870);
xnor U6235 (N_6235,In_2332,In_9);
and U6236 (N_6236,In_77,In_1390);
nor U6237 (N_6237,In_2146,In_1501);
or U6238 (N_6238,In_1287,In_640);
or U6239 (N_6239,In_1251,In_1613);
nor U6240 (N_6240,In_17,In_1444);
xor U6241 (N_6241,In_641,In_2263);
xor U6242 (N_6242,In_1332,In_57);
nor U6243 (N_6243,In_688,In_2312);
and U6244 (N_6244,In_1410,In_2489);
xnor U6245 (N_6245,In_584,In_1243);
xor U6246 (N_6246,In_1733,In_1683);
or U6247 (N_6247,In_1072,In_110);
nand U6248 (N_6248,In_197,In_733);
or U6249 (N_6249,In_1359,In_1677);
xnor U6250 (N_6250,N_1491,N_1421);
nor U6251 (N_6251,N_3173,N_1053);
nor U6252 (N_6252,N_5516,N_4365);
or U6253 (N_6253,N_4484,N_2825);
and U6254 (N_6254,N_3980,N_4379);
nand U6255 (N_6255,N_4296,N_2004);
nand U6256 (N_6256,N_965,N_5183);
xnor U6257 (N_6257,N_6103,N_1969);
nor U6258 (N_6258,N_848,N_450);
xnor U6259 (N_6259,N_1681,N_804);
nor U6260 (N_6260,N_751,N_1467);
or U6261 (N_6261,N_5170,N_6073);
nand U6262 (N_6262,N_1692,N_1536);
nand U6263 (N_6263,N_3888,N_5883);
and U6264 (N_6264,N_4571,N_4579);
or U6265 (N_6265,N_2776,N_2333);
and U6266 (N_6266,N_5642,N_3991);
nor U6267 (N_6267,N_2048,N_1135);
or U6268 (N_6268,N_4052,N_1941);
nor U6269 (N_6269,N_2810,N_1189);
or U6270 (N_6270,N_858,N_5607);
and U6271 (N_6271,N_3975,N_6204);
or U6272 (N_6272,N_924,N_1523);
or U6273 (N_6273,N_5485,N_4454);
nand U6274 (N_6274,N_4605,N_516);
nor U6275 (N_6275,N_877,N_2457);
or U6276 (N_6276,N_3263,N_4587);
xor U6277 (N_6277,N_897,N_4528);
xnor U6278 (N_6278,N_4827,N_2889);
and U6279 (N_6279,N_546,N_5254);
nor U6280 (N_6280,N_888,N_4374);
nand U6281 (N_6281,N_2199,N_605);
or U6282 (N_6282,N_5052,N_1717);
nor U6283 (N_6283,N_5178,N_2947);
nor U6284 (N_6284,N_4930,N_2781);
and U6285 (N_6285,N_526,N_383);
nand U6286 (N_6286,N_1530,N_1817);
nand U6287 (N_6287,N_14,N_4487);
nor U6288 (N_6288,N_3670,N_2753);
and U6289 (N_6289,N_5159,N_4691);
nand U6290 (N_6290,N_5173,N_4072);
and U6291 (N_6291,N_2713,N_4339);
or U6292 (N_6292,N_3167,N_5697);
xor U6293 (N_6293,N_3508,N_6243);
xnor U6294 (N_6294,N_3278,N_2643);
nor U6295 (N_6295,N_312,N_3480);
nand U6296 (N_6296,N_1628,N_1201);
or U6297 (N_6297,N_927,N_5741);
or U6298 (N_6298,N_5804,N_3731);
nor U6299 (N_6299,N_5821,N_1736);
nor U6300 (N_6300,N_2299,N_5181);
nor U6301 (N_6301,N_5470,N_955);
and U6302 (N_6302,N_1193,N_4896);
nor U6303 (N_6303,N_2324,N_2394);
and U6304 (N_6304,N_345,N_892);
and U6305 (N_6305,N_4117,N_1771);
or U6306 (N_6306,N_4793,N_3634);
or U6307 (N_6307,N_486,N_1379);
and U6308 (N_6308,N_3621,N_5836);
nor U6309 (N_6309,N_640,N_1587);
nand U6310 (N_6310,N_4898,N_214);
or U6311 (N_6311,N_4888,N_2057);
nor U6312 (N_6312,N_5288,N_678);
nor U6313 (N_6313,N_1440,N_505);
or U6314 (N_6314,N_2763,N_1990);
nand U6315 (N_6315,N_386,N_3482);
or U6316 (N_6316,N_4126,N_223);
xnor U6317 (N_6317,N_2282,N_932);
nor U6318 (N_6318,N_15,N_232);
nor U6319 (N_6319,N_2801,N_6116);
or U6320 (N_6320,N_811,N_3632);
or U6321 (N_6321,N_373,N_5500);
and U6322 (N_6322,N_2498,N_33);
nand U6323 (N_6323,N_202,N_6011);
or U6324 (N_6324,N_534,N_2647);
and U6325 (N_6325,N_3882,N_613);
nor U6326 (N_6326,N_2486,N_2599);
nor U6327 (N_6327,N_3082,N_2002);
nand U6328 (N_6328,N_5997,N_4711);
xnor U6329 (N_6329,N_3658,N_6217);
nor U6330 (N_6330,N_2441,N_339);
nand U6331 (N_6331,N_3815,N_5626);
and U6332 (N_6332,N_3635,N_3387);
and U6333 (N_6333,N_4224,N_2704);
nand U6334 (N_6334,N_4663,N_191);
or U6335 (N_6335,N_3148,N_1217);
nand U6336 (N_6336,N_3998,N_6238);
nand U6337 (N_6337,N_4724,N_77);
nand U6338 (N_6338,N_822,N_102);
and U6339 (N_6339,N_2092,N_2641);
nand U6340 (N_6340,N_4275,N_5056);
and U6341 (N_6341,N_6086,N_1585);
and U6342 (N_6342,N_3329,N_2232);
and U6343 (N_6343,N_750,N_5542);
xor U6344 (N_6344,N_352,N_6182);
nand U6345 (N_6345,N_592,N_5157);
nand U6346 (N_6346,N_2165,N_1539);
nand U6347 (N_6347,N_5623,N_524);
or U6348 (N_6348,N_2860,N_4722);
and U6349 (N_6349,N_610,N_2315);
xor U6350 (N_6350,N_830,N_3341);
or U6351 (N_6351,N_1701,N_3025);
nor U6352 (N_6352,N_5737,N_1586);
or U6353 (N_6353,N_3091,N_919);
or U6354 (N_6354,N_2521,N_948);
or U6355 (N_6355,N_1289,N_3138);
xor U6356 (N_6356,N_3129,N_2135);
and U6357 (N_6357,N_1735,N_4078);
nand U6358 (N_6358,N_2190,N_2533);
and U6359 (N_6359,N_6236,N_2522);
and U6360 (N_6360,N_704,N_2462);
or U6361 (N_6361,N_2212,N_4601);
xnor U6362 (N_6362,N_3610,N_5942);
nor U6363 (N_6363,N_5368,N_3075);
nand U6364 (N_6364,N_1420,N_5127);
xor U6365 (N_6365,N_2818,N_2407);
nor U6366 (N_6366,N_4734,N_6222);
nand U6367 (N_6367,N_1091,N_4560);
nor U6368 (N_6368,N_1690,N_4730);
xor U6369 (N_6369,N_4949,N_4166);
or U6370 (N_6370,N_2539,N_4141);
xnor U6371 (N_6371,N_797,N_5193);
nand U6372 (N_6372,N_4941,N_4806);
or U6373 (N_6373,N_5184,N_3517);
nand U6374 (N_6374,N_2391,N_187);
or U6375 (N_6375,N_6199,N_3017);
and U6376 (N_6376,N_418,N_831);
nand U6377 (N_6377,N_5442,N_2025);
nand U6378 (N_6378,N_4869,N_233);
xor U6379 (N_6379,N_4829,N_2708);
nor U6380 (N_6380,N_23,N_773);
nand U6381 (N_6381,N_1557,N_2714);
nor U6382 (N_6382,N_3713,N_2274);
nand U6383 (N_6383,N_2369,N_6050);
nand U6384 (N_6384,N_3344,N_2344);
and U6385 (N_6385,N_3532,N_2275);
nor U6386 (N_6386,N_5010,N_2728);
or U6387 (N_6387,N_2466,N_1742);
and U6388 (N_6388,N_817,N_5436);
nor U6389 (N_6389,N_3143,N_3768);
nand U6390 (N_6390,N_4727,N_2623);
nor U6391 (N_6391,N_819,N_4522);
or U6392 (N_6392,N_2502,N_4045);
nor U6393 (N_6393,N_2663,N_4708);
or U6394 (N_6394,N_2311,N_4776);
nor U6395 (N_6395,N_40,N_5208);
or U6396 (N_6396,N_4502,N_2388);
nand U6397 (N_6397,N_3649,N_5329);
nor U6398 (N_6398,N_5247,N_5979);
and U6399 (N_6399,N_2666,N_5083);
and U6400 (N_6400,N_4813,N_2906);
or U6401 (N_6401,N_2565,N_1351);
nand U6402 (N_6402,N_1583,N_5335);
and U6403 (N_6403,N_2305,N_4124);
nor U6404 (N_6404,N_5411,N_3229);
or U6405 (N_6405,N_2553,N_2444);
nor U6406 (N_6406,N_3030,N_2604);
xor U6407 (N_6407,N_902,N_5396);
and U6408 (N_6408,N_4410,N_6022);
nand U6409 (N_6409,N_3363,N_2103);
nor U6410 (N_6410,N_913,N_4069);
nor U6411 (N_6411,N_5926,N_2674);
nor U6412 (N_6412,N_248,N_2187);
nor U6413 (N_6413,N_4448,N_2106);
or U6414 (N_6414,N_5226,N_1609);
or U6415 (N_6415,N_256,N_3972);
or U6416 (N_6416,N_5005,N_1873);
nand U6417 (N_6417,N_3429,N_3059);
nor U6418 (N_6418,N_3425,N_497);
xnor U6419 (N_6419,N_1079,N_189);
nand U6420 (N_6420,N_6017,N_1521);
xor U6421 (N_6421,N_1296,N_3166);
nand U6422 (N_6422,N_3958,N_5662);
xor U6423 (N_6423,N_3806,N_3664);
xnor U6424 (N_6424,N_2816,N_2181);
nor U6425 (N_6425,N_2570,N_4616);
or U6426 (N_6426,N_4998,N_5412);
or U6427 (N_6427,N_5070,N_6147);
or U6428 (N_6428,N_3995,N_6087);
or U6429 (N_6429,N_4515,N_4274);
nand U6430 (N_6430,N_2918,N_3733);
nor U6431 (N_6431,N_3916,N_6145);
nand U6432 (N_6432,N_3944,N_5944);
nor U6433 (N_6433,N_4043,N_1021);
xor U6434 (N_6434,N_2630,N_28);
xor U6435 (N_6435,N_2850,N_3356);
or U6436 (N_6436,N_3624,N_1556);
and U6437 (N_6437,N_960,N_2900);
nand U6438 (N_6438,N_1697,N_375);
nor U6439 (N_6439,N_4160,N_1473);
and U6440 (N_6440,N_1288,N_4324);
and U6441 (N_6441,N_4053,N_2872);
and U6442 (N_6442,N_1429,N_2428);
and U6443 (N_6443,N_4264,N_3230);
nand U6444 (N_6444,N_3495,N_4889);
or U6445 (N_6445,N_4683,N_5624);
and U6446 (N_6446,N_707,N_3040);
nor U6447 (N_6447,N_488,N_2073);
and U6448 (N_6448,N_1611,N_1202);
xnor U6449 (N_6449,N_1286,N_3557);
nor U6450 (N_6450,N_1368,N_108);
and U6451 (N_6451,N_5104,N_304);
xor U6452 (N_6452,N_4899,N_4646);
nand U6453 (N_6453,N_2691,N_2151);
xor U6454 (N_6454,N_514,N_4830);
nand U6455 (N_6455,N_5976,N_4636);
nor U6456 (N_6456,N_3103,N_1909);
nor U6457 (N_6457,N_5816,N_5456);
and U6458 (N_6458,N_1487,N_4895);
nor U6459 (N_6459,N_5866,N_1834);
and U6460 (N_6460,N_2617,N_1457);
and U6461 (N_6461,N_4157,N_4098);
xnor U6462 (N_6462,N_5295,N_4282);
and U6463 (N_6463,N_3638,N_936);
and U6464 (N_6464,N_676,N_4721);
nand U6465 (N_6465,N_2509,N_1950);
nor U6466 (N_6466,N_5192,N_3812);
nor U6467 (N_6467,N_2950,N_1031);
nand U6468 (N_6468,N_966,N_4915);
and U6469 (N_6469,N_2110,N_6149);
xnor U6470 (N_6470,N_5538,N_1542);
nor U6471 (N_6471,N_466,N_0);
and U6472 (N_6472,N_4247,N_1112);
or U6473 (N_6473,N_1117,N_2952);
nor U6474 (N_6474,N_5510,N_4064);
nor U6475 (N_6475,N_1037,N_481);
nand U6476 (N_6476,N_5079,N_4285);
or U6477 (N_6477,N_1694,N_1165);
nor U6478 (N_6478,N_1669,N_5068);
or U6479 (N_6479,N_367,N_4625);
nor U6480 (N_6480,N_3603,N_4990);
nand U6481 (N_6481,N_4859,N_4745);
and U6482 (N_6482,N_4731,N_462);
nor U6483 (N_6483,N_1656,N_1745);
xor U6484 (N_6484,N_4598,N_53);
or U6485 (N_6485,N_3493,N_299);
nor U6486 (N_6486,N_834,N_2141);
or U6487 (N_6487,N_1899,N_1084);
or U6488 (N_6488,N_195,N_1216);
nand U6489 (N_6489,N_1349,N_2686);
nand U6490 (N_6490,N_6053,N_2717);
nor U6491 (N_6491,N_1398,N_2839);
and U6492 (N_6492,N_3097,N_452);
xor U6493 (N_6493,N_1748,N_301);
nand U6494 (N_6494,N_4197,N_5695);
nand U6495 (N_6495,N_5131,N_5932);
and U6496 (N_6496,N_4828,N_547);
and U6497 (N_6497,N_1125,N_1744);
and U6498 (N_6498,N_1483,N_5887);
nand U6499 (N_6499,N_3487,N_2870);
nand U6500 (N_6500,N_1926,N_2490);
or U6501 (N_6501,N_2297,N_6152);
nor U6502 (N_6502,N_3988,N_3565);
nand U6503 (N_6503,N_636,N_3012);
or U6504 (N_6504,N_766,N_4362);
or U6505 (N_6505,N_3739,N_2113);
and U6506 (N_6506,N_4497,N_2939);
nand U6507 (N_6507,N_2400,N_5433);
xor U6508 (N_6508,N_595,N_1034);
nand U6509 (N_6509,N_5930,N_2018);
nand U6510 (N_6510,N_4378,N_4087);
nand U6511 (N_6511,N_2052,N_1672);
or U6512 (N_6512,N_2660,N_5647);
and U6513 (N_6513,N_110,N_624);
and U6514 (N_6514,N_4303,N_4879);
xnor U6515 (N_6515,N_1612,N_1321);
nor U6516 (N_6516,N_1277,N_5479);
nor U6517 (N_6517,N_2312,N_5385);
and U6518 (N_6518,N_4059,N_1755);
nor U6519 (N_6519,N_2302,N_5894);
nand U6520 (N_6520,N_438,N_2208);
or U6521 (N_6521,N_1997,N_4682);
nand U6522 (N_6522,N_3709,N_2795);
nor U6523 (N_6523,N_4753,N_3013);
xnor U6524 (N_6524,N_2329,N_6008);
nand U6525 (N_6525,N_3695,N_5467);
and U6526 (N_6526,N_4989,N_2045);
and U6527 (N_6527,N_1638,N_1984);
nor U6528 (N_6528,N_3918,N_2615);
and U6529 (N_6529,N_2347,N_4027);
nand U6530 (N_6530,N_5840,N_147);
nor U6531 (N_6531,N_6220,N_1213);
or U6532 (N_6532,N_4143,N_3513);
nor U6533 (N_6533,N_5016,N_5994);
xor U6534 (N_6534,N_6009,N_3711);
or U6535 (N_6535,N_3239,N_779);
or U6536 (N_6536,N_1702,N_527);
nand U6537 (N_6537,N_3016,N_3725);
nor U6538 (N_6538,N_5921,N_2955);
xor U6539 (N_6539,N_2170,N_5488);
nor U6540 (N_6540,N_2916,N_6100);
nor U6541 (N_6541,N_1826,N_5570);
and U6542 (N_6542,N_3024,N_2272);
or U6543 (N_6543,N_403,N_4486);
nand U6544 (N_6544,N_4581,N_1438);
or U6545 (N_6545,N_3585,N_3851);
nor U6546 (N_6546,N_3022,N_4890);
xnor U6547 (N_6547,N_5933,N_1258);
or U6548 (N_6548,N_4337,N_1495);
or U6549 (N_6549,N_3477,N_41);
and U6550 (N_6550,N_5886,N_545);
nor U6551 (N_6551,N_4505,N_2039);
and U6552 (N_6552,N_2238,N_5936);
or U6553 (N_6553,N_2065,N_1914);
xnor U6554 (N_6554,N_4133,N_5354);
and U6555 (N_6555,N_1892,N_5080);
or U6556 (N_6556,N_1283,N_371);
nor U6557 (N_6557,N_5913,N_6025);
or U6558 (N_6558,N_5120,N_2633);
and U6559 (N_6559,N_5164,N_5273);
or U6560 (N_6560,N_3858,N_641);
or U6561 (N_6561,N_1360,N_400);
or U6562 (N_6562,N_2276,N_1036);
and U6563 (N_6563,N_4749,N_1600);
nand U6564 (N_6564,N_899,N_5029);
nor U6565 (N_6565,N_1679,N_5058);
and U6566 (N_6566,N_3755,N_5478);
or U6567 (N_6567,N_1174,N_3920);
nor U6568 (N_6568,N_747,N_1953);
and U6569 (N_6569,N_5884,N_3784);
nand U6570 (N_6570,N_324,N_922);
or U6571 (N_6571,N_1439,N_5549);
nand U6572 (N_6572,N_2224,N_4084);
and U6573 (N_6573,N_2259,N_5338);
nor U6574 (N_6574,N_4739,N_4519);
xnor U6575 (N_6575,N_3843,N_6055);
or U6576 (N_6576,N_3941,N_5537);
nor U6577 (N_6577,N_4152,N_1668);
nand U6578 (N_6578,N_4777,N_4139);
and U6579 (N_6579,N_4544,N_2695);
or U6580 (N_6580,N_4447,N_2062);
nand U6581 (N_6581,N_3574,N_4032);
and U6582 (N_6582,N_2371,N_59);
nor U6583 (N_6583,N_5434,N_4402);
nor U6584 (N_6584,N_1376,N_939);
and U6585 (N_6585,N_231,N_5204);
nor U6586 (N_6586,N_3298,N_5163);
xnor U6587 (N_6587,N_1069,N_240);
and U6588 (N_6588,N_1102,N_6034);
nor U6589 (N_6589,N_4313,N_2013);
xor U6590 (N_6590,N_2067,N_4760);
or U6591 (N_6591,N_1943,N_5767);
or U6592 (N_6592,N_1478,N_4451);
or U6593 (N_6593,N_6172,N_5613);
or U6594 (N_6594,N_1490,N_381);
nand U6595 (N_6595,N_94,N_3209);
and U6596 (N_6596,N_886,N_946);
and U6597 (N_6597,N_3449,N_1263);
or U6598 (N_6598,N_5091,N_4476);
xor U6599 (N_6599,N_1657,N_3824);
or U6600 (N_6600,N_1610,N_5961);
and U6601 (N_6601,N_4535,N_5671);
or U6602 (N_6602,N_5285,N_3475);
nor U6603 (N_6603,N_4853,N_1548);
nand U6604 (N_6604,N_5620,N_2390);
nand U6605 (N_6605,N_3161,N_379);
xor U6606 (N_6606,N_4426,N_1226);
or U6607 (N_6607,N_5829,N_3836);
or U6608 (N_6608,N_2940,N_5879);
nor U6609 (N_6609,N_84,N_4135);
nand U6610 (N_6610,N_3290,N_323);
or U6611 (N_6611,N_630,N_3932);
and U6612 (N_6612,N_4526,N_5701);
and U6613 (N_6613,N_517,N_765);
nor U6614 (N_6614,N_5097,N_1965);
nand U6615 (N_6615,N_3677,N_5723);
nor U6616 (N_6616,N_2771,N_4199);
xnor U6617 (N_6617,N_5319,N_5677);
or U6618 (N_6618,N_3394,N_4129);
nand U6619 (N_6619,N_1847,N_4875);
nor U6620 (N_6620,N_4283,N_2150);
or U6621 (N_6621,N_5771,N_4332);
or U6622 (N_6622,N_3646,N_1024);
nor U6623 (N_6623,N_3301,N_267);
nor U6624 (N_6624,N_2454,N_3072);
and U6625 (N_6625,N_4765,N_3068);
and U6626 (N_6626,N_5574,N_4784);
nor U6627 (N_6627,N_1866,N_4832);
or U6628 (N_6628,N_2746,N_5006);
nor U6629 (N_6629,N_5062,N_4521);
and U6630 (N_6630,N_1956,N_5202);
and U6631 (N_6631,N_5528,N_5931);
or U6632 (N_6632,N_6134,N_2205);
nand U6633 (N_6633,N_5639,N_758);
or U6634 (N_6634,N_5,N_5293);
xor U6635 (N_6635,N_1636,N_5205);
nand U6636 (N_6636,N_612,N_6097);
nand U6637 (N_6637,N_484,N_5235);
or U6638 (N_6638,N_717,N_5506);
nor U6639 (N_6639,N_4311,N_35);
and U6640 (N_6640,N_3339,N_681);
nor U6641 (N_6641,N_995,N_224);
and U6642 (N_6642,N_5043,N_1381);
nor U6643 (N_6643,N_4433,N_1940);
nor U6644 (N_6644,N_4621,N_4886);
or U6645 (N_6645,N_5735,N_1815);
or U6646 (N_6646,N_2374,N_4872);
and U6647 (N_6647,N_4300,N_3903);
and U6648 (N_6648,N_111,N_4914);
nor U6649 (N_6649,N_1804,N_60);
or U6650 (N_6650,N_5860,N_5362);
nor U6651 (N_6651,N_3939,N_364);
or U6652 (N_6652,N_4801,N_4111);
xnor U6653 (N_6653,N_331,N_5521);
xnor U6654 (N_6654,N_3316,N_4661);
nor U6655 (N_6655,N_5310,N_5325);
nor U6656 (N_6656,N_5561,N_5614);
or U6657 (N_6657,N_1671,N_332);
xnor U6658 (N_6658,N_2377,N_2654);
or U6659 (N_6659,N_3297,N_1330);
nor U6660 (N_6660,N_2336,N_170);
nand U6661 (N_6661,N_1642,N_2147);
and U6662 (N_6662,N_3866,N_5633);
nand U6663 (N_6663,N_4343,N_5901);
or U6664 (N_6664,N_4929,N_1220);
or U6665 (N_6665,N_368,N_3362);
nor U6666 (N_6666,N_1785,N_4954);
and U6667 (N_6667,N_1477,N_3149);
nand U6668 (N_6668,N_1803,N_687);
or U6669 (N_6669,N_602,N_4863);
or U6670 (N_6670,N_2267,N_5489);
and U6671 (N_6671,N_30,N_5405);
and U6672 (N_6672,N_4916,N_2619);
nand U6673 (N_6673,N_4017,N_5182);
xnor U6674 (N_6674,N_327,N_5761);
nand U6675 (N_6675,N_5458,N_5371);
xor U6676 (N_6676,N_787,N_6130);
nor U6677 (N_6677,N_937,N_2343);
or U6678 (N_6678,N_1905,N_3561);
xnor U6679 (N_6679,N_1828,N_4965);
or U6680 (N_6680,N_4979,N_5365);
and U6681 (N_6681,N_2523,N_5684);
nor U6682 (N_6682,N_2136,N_2264);
or U6683 (N_6683,N_2153,N_4472);
and U6684 (N_6684,N_4694,N_917);
nand U6685 (N_6685,N_5679,N_3431);
nor U6686 (N_6686,N_4079,N_495);
nor U6687 (N_6687,N_4946,N_4719);
nor U6688 (N_6688,N_3950,N_1047);
or U6689 (N_6689,N_4715,N_2707);
xnor U6690 (N_6690,N_4018,N_1666);
or U6691 (N_6691,N_623,N_1391);
nor U6692 (N_6692,N_2295,N_1088);
nand U6693 (N_6693,N_3539,N_3355);
nand U6694 (N_6694,N_5999,N_4452);
xnor U6695 (N_6695,N_1018,N_695);
xnor U6696 (N_6696,N_2219,N_1540);
nor U6697 (N_6697,N_1684,N_5355);
or U6698 (N_6698,N_4993,N_3586);
and U6699 (N_6699,N_3497,N_4307);
or U6700 (N_6700,N_4630,N_5520);
or U6701 (N_6701,N_5518,N_3524);
nor U6702 (N_6702,N_2887,N_1331);
nand U6703 (N_6703,N_5832,N_565);
and U6704 (N_6704,N_4980,N_166);
or U6705 (N_6705,N_3124,N_5591);
nand U6706 (N_6706,N_3809,N_1759);
and U6707 (N_6707,N_791,N_4594);
and U6708 (N_6708,N_2693,N_34);
xor U6709 (N_6709,N_3974,N_445);
xor U6710 (N_6710,N_1718,N_2882);
nand U6711 (N_6711,N_3118,N_1741);
nand U6712 (N_6712,N_3422,N_2005);
nand U6713 (N_6713,N_2284,N_1040);
nand U6714 (N_6714,N_2855,N_3896);
nand U6715 (N_6715,N_1810,N_3247);
or U6716 (N_6716,N_5323,N_5661);
or U6717 (N_6717,N_5511,N_3369);
xnor U6718 (N_6718,N_151,N_645);
nor U6719 (N_6719,N_5486,N_3570);
and U6720 (N_6720,N_346,N_4858);
nor U6721 (N_6721,N_5611,N_4241);
or U6722 (N_6722,N_728,N_5417);
nor U6723 (N_6723,N_3427,N_4913);
or U6724 (N_6724,N_49,N_5158);
nor U6725 (N_6725,N_4650,N_3292);
and U6726 (N_6726,N_1375,N_4210);
xor U6727 (N_6727,N_2114,N_1145);
or U6728 (N_6728,N_2662,N_1013);
nand U6729 (N_6729,N_665,N_3364);
nor U6730 (N_6730,N_6098,N_4261);
nor U6731 (N_6731,N_3259,N_3569);
and U6732 (N_6732,N_3101,N_4216);
and U6733 (N_6733,N_3264,N_2246);
nand U6734 (N_6734,N_1845,N_1299);
or U6735 (N_6735,N_5953,N_82);
or U6736 (N_6736,N_5215,N_2167);
or U6737 (N_6737,N_4912,N_273);
nor U6738 (N_6738,N_5265,N_5014);
nand U6739 (N_6739,N_3073,N_5406);
or U6740 (N_6740,N_1566,N_3488);
nor U6741 (N_6741,N_956,N_4825);
nand U6742 (N_6742,N_2881,N_3067);
nor U6743 (N_6743,N_912,N_1562);
or U6744 (N_6744,N_5220,N_1703);
or U6745 (N_6745,N_1868,N_3639);
and U6746 (N_6746,N_1942,N_2574);
nand U6747 (N_6747,N_5099,N_2531);
or U6748 (N_6748,N_4237,N_1249);
and U6749 (N_6749,N_2721,N_1081);
or U6750 (N_6750,N_1348,N_5276);
nor U6751 (N_6751,N_2108,N_3358);
or U6752 (N_6752,N_5952,N_6155);
nor U6753 (N_6753,N_3845,N_5216);
nor U6754 (N_6754,N_6188,N_4769);
or U6755 (N_6755,N_3692,N_2375);
and U6756 (N_6756,N_6240,N_1293);
and U6757 (N_6757,N_3965,N_5197);
or U6758 (N_6758,N_576,N_3010);
nor U6759 (N_6759,N_3198,N_1639);
nor U6760 (N_6760,N_574,N_4773);
nor U6761 (N_6761,N_1132,N_5221);
xor U6762 (N_6762,N_4764,N_353);
nand U6763 (N_6763,N_266,N_2249);
and U6764 (N_6764,N_2239,N_6225);
and U6765 (N_6765,N_4942,N_3752);
or U6766 (N_6766,N_3246,N_4293);
xor U6767 (N_6767,N_4702,N_2321);
nand U6768 (N_6768,N_4738,N_1714);
or U6769 (N_6769,N_206,N_951);
nand U6770 (N_6770,N_3107,N_1016);
xnor U6771 (N_6771,N_5289,N_1461);
and U6772 (N_6772,N_5369,N_540);
nand U6773 (N_6773,N_2427,N_98);
nand U6774 (N_6774,N_378,N_1635);
nor U6775 (N_6775,N_667,N_5589);
nor U6776 (N_6776,N_2893,N_358);
nand U6777 (N_6777,N_617,N_5364);
nor U6778 (N_6778,N_2075,N_5859);
nand U6779 (N_6779,N_2145,N_3114);
nand U6780 (N_6780,N_2518,N_977);
and U6781 (N_6781,N_3009,N_4208);
xnor U6782 (N_6782,N_5249,N_5222);
or U6783 (N_6783,N_5604,N_2492);
or U6784 (N_6784,N_548,N_3415);
nor U6785 (N_6785,N_5051,N_4235);
nor U6786 (N_6786,N_4910,N_2084);
nand U6787 (N_6787,N_118,N_1696);
nand U6788 (N_6788,N_1187,N_2448);
or U6789 (N_6789,N_4228,N_2750);
or U6790 (N_6790,N_6239,N_2440);
and U6791 (N_6791,N_6226,N_2086);
and U6792 (N_6792,N_1778,N_5213);
and U6793 (N_6793,N_123,N_3318);
or U6794 (N_6794,N_6164,N_5752);
xnor U6795 (N_6795,N_6038,N_3281);
nor U6796 (N_6796,N_3174,N_300);
nand U6797 (N_6797,N_3277,N_2536);
and U6798 (N_6798,N_5945,N_5664);
nor U6799 (N_6799,N_105,N_3630);
nor U6800 (N_6800,N_4156,N_2868);
and U6801 (N_6801,N_5706,N_598);
nand U6802 (N_6802,N_3535,N_3669);
nor U6803 (N_6803,N_1342,N_2439);
or U6804 (N_6804,N_5794,N_710);
nand U6805 (N_6805,N_1114,N_247);
or U6806 (N_6806,N_2864,N_2354);
nand U6807 (N_6807,N_2649,N_5269);
xnor U6808 (N_6808,N_1253,N_768);
nand U6809 (N_6809,N_572,N_6141);
xnor U6810 (N_6810,N_496,N_1652);
and U6811 (N_6811,N_148,N_544);
or U6812 (N_6812,N_5210,N_2851);
and U6813 (N_6813,N_4155,N_2467);
nand U6814 (N_6814,N_2520,N_1463);
nand U6815 (N_6815,N_5237,N_3598);
and U6816 (N_6816,N_1798,N_3228);
nor U6817 (N_6817,N_823,N_1169);
nor U6818 (N_6818,N_5747,N_1469);
nand U6819 (N_6819,N_3973,N_5758);
nor U6820 (N_6820,N_2719,N_2938);
and U6821 (N_6821,N_5093,N_3642);
nor U6822 (N_6822,N_5617,N_1241);
or U6823 (N_6823,N_5851,N_2410);
nand U6824 (N_6824,N_2813,N_164);
nor U6825 (N_6825,N_5874,N_3345);
nor U6826 (N_6826,N_19,N_3056);
nand U6827 (N_6827,N_2821,N_3325);
nand U6828 (N_6828,N_2992,N_1030);
nor U6829 (N_6829,N_5721,N_3880);
and U6830 (N_6830,N_1854,N_3807);
xor U6831 (N_6831,N_1544,N_910);
xnor U6832 (N_6832,N_5141,N_609);
nand U6833 (N_6833,N_1148,N_5464);
nor U6834 (N_6834,N_5318,N_4288);
xnor U6835 (N_6835,N_5796,N_1517);
or U6836 (N_6836,N_5227,N_529);
nor U6837 (N_6837,N_4845,N_2314);
or U6838 (N_6838,N_5982,N_3979);
or U6839 (N_6839,N_5410,N_4567);
nand U6840 (N_6840,N_4978,N_2665);
or U6841 (N_6841,N_4613,N_5086);
or U6842 (N_6842,N_2642,N_2703);
nor U6843 (N_6843,N_4444,N_447);
nand U6844 (N_6844,N_746,N_3179);
or U6845 (N_6845,N_4504,N_1149);
or U6846 (N_6846,N_5900,N_1916);
or U6847 (N_6847,N_3581,N_3864);
nand U6848 (N_6848,N_458,N_1840);
and U6849 (N_6849,N_3032,N_4563);
nand U6850 (N_6850,N_325,N_1917);
nor U6851 (N_6851,N_5648,N_1369);
and U6852 (N_6852,N_2863,N_4540);
and U6853 (N_6853,N_3000,N_2985);
nand U6854 (N_6854,N_4269,N_938);
and U6855 (N_6855,N_283,N_3351);
nand U6856 (N_6856,N_2689,N_5004);
nand U6857 (N_6857,N_5943,N_1301);
nor U6858 (N_6858,N_3104,N_374);
and U6859 (N_6859,N_5581,N_5228);
nand U6860 (N_6860,N_5654,N_1912);
nor U6861 (N_6861,N_844,N_1294);
xnor U6862 (N_6862,N_1897,N_5791);
or U6863 (N_6863,N_2352,N_5367);
or U6864 (N_6864,N_4258,N_5251);
nor U6865 (N_6865,N_183,N_3510);
or U6866 (N_6866,N_427,N_3145);
and U6867 (N_6867,N_3934,N_286);
or U6868 (N_6868,N_1768,N_6231);
and U6869 (N_6869,N_1648,N_4783);
or U6870 (N_6870,N_1911,N_1830);
nand U6871 (N_6871,N_5774,N_4592);
and U6872 (N_6872,N_4437,N_738);
or U6873 (N_6873,N_2929,N_1096);
xor U6874 (N_6874,N_1448,N_465);
and U6875 (N_6875,N_3360,N_1514);
nor U6876 (N_6876,N_2234,N_5077);
nand U6877 (N_6877,N_4539,N_589);
or U6878 (N_6878,N_5359,N_1528);
or U6879 (N_6879,N_4918,N_5722);
nor U6880 (N_6880,N_3719,N_756);
and U6881 (N_6881,N_853,N_1560);
nand U6882 (N_6882,N_5792,N_2716);
nand U6883 (N_6883,N_2221,N_333);
or U6884 (N_6884,N_2460,N_833);
nor U6885 (N_6885,N_5496,N_3884);
nand U6886 (N_6886,N_5813,N_4024);
or U6887 (N_6887,N_215,N_6107);
xor U6888 (N_6888,N_1849,N_5420);
xnor U6889 (N_6889,N_5003,N_3550);
nor U6890 (N_6890,N_764,N_1971);
and U6891 (N_6891,N_476,N_3391);
and U6892 (N_6892,N_2386,N_506);
nor U6893 (N_6893,N_4710,N_1285);
and U6894 (N_6894,N_4415,N_3566);
and U6895 (N_6895,N_4971,N_29);
xnor U6896 (N_6896,N_2620,N_2121);
nor U6897 (N_6897,N_2139,N_3879);
nand U6898 (N_6898,N_3204,N_4195);
nand U6899 (N_6899,N_3559,N_2572);
and U6900 (N_6900,N_895,N_1152);
or U6901 (N_6901,N_5906,N_4676);
nor U6902 (N_6902,N_5324,N_601);
or U6903 (N_6903,N_3343,N_437);
nor U6904 (N_6904,N_1163,N_5888);
or U6905 (N_6905,N_639,N_671);
xor U6906 (N_6906,N_4717,N_199);
xor U6907 (N_6907,N_4047,N_4549);
or U6908 (N_6908,N_4038,N_593);
nor U6909 (N_6909,N_3892,N_889);
and U6910 (N_6910,N_4004,N_3074);
and U6911 (N_6911,N_5196,N_5008);
nor U6912 (N_6912,N_4525,N_2035);
or U6913 (N_6913,N_1056,N_3165);
xnor U6914 (N_6914,N_998,N_5152);
or U6915 (N_6915,N_4639,N_3891);
nor U6916 (N_6916,N_1670,N_3342);
nand U6917 (N_6917,N_1746,N_2398);
and U6918 (N_6918,N_3152,N_2326);
and U6919 (N_6919,N_5240,N_244);
xnor U6920 (N_6920,N_860,N_237);
or U6921 (N_6921,N_3,N_753);
nor U6922 (N_6922,N_91,N_5799);
nand U6923 (N_6923,N_1352,N_5150);
nor U6924 (N_6924,N_329,N_5059);
and U6925 (N_6925,N_211,N_5555);
or U6926 (N_6926,N_5407,N_3746);
nor U6927 (N_6927,N_2587,N_3863);
or U6928 (N_6928,N_5194,N_6066);
nor U6929 (N_6929,N_2550,N_4364);
and U6930 (N_6930,N_4273,N_2317);
or U6931 (N_6931,N_2203,N_20);
and U6932 (N_6932,N_6060,N_4386);
nand U6933 (N_6933,N_4060,N_197);
nand U6934 (N_6934,N_2724,N_2547);
nor U6935 (N_6935,N_1927,N_3685);
or U6936 (N_6936,N_167,N_4624);
and U6937 (N_6937,N_5560,N_1214);
nor U6938 (N_6938,N_2843,N_4552);
or U6939 (N_6939,N_2242,N_631);
nand U6940 (N_6940,N_1654,N_2318);
or U6941 (N_6941,N_2527,N_4012);
nand U6942 (N_6942,N_2884,N_396);
xnor U6943 (N_6943,N_2698,N_3823);
and U6944 (N_6944,N_2741,N_4039);
nand U6945 (N_6945,N_4503,N_3584);
nand U6946 (N_6946,N_5377,N_1058);
or U6947 (N_6947,N_4514,N_42);
and U6948 (N_6948,N_2791,N_3266);
nor U6949 (N_6949,N_2257,N_4115);
or U6950 (N_6950,N_4441,N_4358);
nand U6951 (N_6951,N_2726,N_1818);
nor U6952 (N_6952,N_4943,N_3041);
nor U6953 (N_6953,N_5267,N_5439);
or U6954 (N_6954,N_430,N_5529);
xor U6955 (N_6955,N_2867,N_3412);
and U6956 (N_6956,N_1252,N_6163);
nand U6957 (N_6957,N_478,N_3168);
and U6958 (N_6958,N_1064,N_5258);
and U6959 (N_6959,N_4583,N_5606);
and U6960 (N_6960,N_1430,N_5209);
nor U6961 (N_6961,N_568,N_2255);
or U6962 (N_6962,N_2975,N_5937);
and U6963 (N_6963,N_2001,N_5383);
and U6964 (N_6964,N_3255,N_2207);
and U6965 (N_6965,N_1945,N_1191);
and U6966 (N_6966,N_4394,N_4499);
or U6967 (N_6967,N_1077,N_2452);
or U6968 (N_6968,N_5343,N_2034);
xor U6969 (N_6969,N_3956,N_6035);
xnor U6970 (N_6970,N_606,N_4036);
and U6971 (N_6971,N_2577,N_3096);
or U6972 (N_6972,N_3441,N_3180);
xor U6973 (N_6973,N_6132,N_4336);
or U6974 (N_6974,N_1831,N_933);
nand U6975 (N_6975,N_5954,N_5873);
nand U6976 (N_6976,N_3968,N_350);
and U6977 (N_6977,N_1498,N_3390);
nand U6978 (N_6978,N_2193,N_2331);
nor U6979 (N_6979,N_2530,N_3287);
nand U6980 (N_6980,N_451,N_5195);
and U6981 (N_6981,N_1176,N_3151);
and U6982 (N_6982,N_4659,N_5892);
or U6983 (N_6983,N_5880,N_2098);
or U6984 (N_6984,N_5833,N_6013);
or U6985 (N_6985,N_2571,N_5539);
and U6986 (N_6986,N_5531,N_2700);
and U6987 (N_6987,N_615,N_4042);
xor U6988 (N_6988,N_1472,N_4229);
or U6989 (N_6989,N_2974,N_5023);
nand U6990 (N_6990,N_1505,N_5045);
or U6991 (N_6991,N_1625,N_561);
or U6992 (N_6992,N_4533,N_3789);
nor U6993 (N_6993,N_1300,N_228);
or U6994 (N_6994,N_5871,N_4440);
or U6995 (N_6995,N_2127,N_62);
or U6996 (N_6996,N_2059,N_3035);
xor U6997 (N_6997,N_3842,N_2729);
and U6998 (N_6998,N_3523,N_4000);
nor U6999 (N_6999,N_4871,N_355);
or U7000 (N_7000,N_3045,N_690);
nor U7001 (N_7001,N_3270,N_4754);
and U7002 (N_7002,N_4076,N_1599);
xnor U7003 (N_7003,N_3811,N_1454);
xnor U7004 (N_7004,N_5315,N_5790);
and U7005 (N_7005,N_1178,N_4360);
or U7006 (N_7006,N_1052,N_3788);
nand U7007 (N_7007,N_3350,N_1417);
or U7008 (N_7008,N_5212,N_1182);
nand U7009 (N_7009,N_3401,N_1343);
xnor U7010 (N_7010,N_3682,N_200);
and U7011 (N_7011,N_4822,N_4326);
xor U7012 (N_7012,N_1157,N_5380);
nor U7013 (N_7013,N_1537,N_4510);
nand U7014 (N_7014,N_5756,N_4788);
or U7015 (N_7015,N_410,N_1266);
nand U7016 (N_7016,N_5474,N_5490);
nor U7017 (N_7017,N_1022,N_4354);
and U7018 (N_7018,N_4668,N_359);
and U7019 (N_7019,N_348,N_2945);
nor U7020 (N_7020,N_727,N_2058);
and U7021 (N_7021,N_4384,N_262);
xor U7022 (N_7022,N_3691,N_2485);
xnor U7023 (N_7023,N_4527,N_492);
and U7024 (N_7024,N_4002,N_3066);
or U7025 (N_7025,N_3541,N_2847);
xor U7026 (N_7026,N_1488,N_1295);
and U7027 (N_7027,N_6030,N_796);
xnor U7028 (N_7028,N_5793,N_5919);
nor U7029 (N_7029,N_4094,N_6084);
or U7030 (N_7030,N_4193,N_967);
nor U7031 (N_7031,N_2206,N_1709);
or U7032 (N_7032,N_5350,N_2891);
nand U7033 (N_7033,N_2636,N_2337);
xor U7034 (N_7034,N_3648,N_4220);
or U7035 (N_7035,N_5509,N_3127);
nor U7036 (N_7036,N_1468,N_6083);
xor U7037 (N_7037,N_771,N_3481);
nor U7038 (N_7038,N_6169,N_1185);
nor U7039 (N_7039,N_1629,N_726);
nor U7040 (N_7040,N_1933,N_795);
nor U7041 (N_7041,N_5000,N_2890);
nor U7042 (N_7042,N_2672,N_3782);
nor U7043 (N_7043,N_2325,N_487);
and U7044 (N_7044,N_4921,N_4368);
nand U7045 (N_7045,N_6216,N_5652);
or U7046 (N_7046,N_173,N_3197);
nor U7047 (N_7047,N_5713,N_4101);
and U7048 (N_7048,N_6058,N_2965);
nand U7049 (N_7049,N_4885,N_3023);
or U7050 (N_7050,N_5956,N_5641);
nor U7051 (N_7051,N_5631,N_4606);
nor U7052 (N_7052,N_757,N_5780);
and U7053 (N_7053,N_3485,N_1355);
or U7054 (N_7054,N_180,N_1946);
nor U7055 (N_7055,N_2681,N_4736);
nor U7056 (N_7056,N_2775,N_969);
xor U7057 (N_7057,N_900,N_4140);
nand U7058 (N_7058,N_774,N_3234);
nand U7059 (N_7059,N_2613,N_5036);
nor U7060 (N_7060,N_5545,N_3943);
or U7061 (N_7061,N_4917,N_5063);
nand U7062 (N_7062,N_3872,N_1316);
and U7063 (N_7063,N_723,N_3420);
and U7064 (N_7064,N_2777,N_3219);
nor U7065 (N_7065,N_3969,N_5111);
nand U7066 (N_7066,N_3680,N_177);
or U7067 (N_7067,N_2180,N_6190);
and U7068 (N_7068,N_3338,N_983);
and U7069 (N_7069,N_1113,N_3336);
or U7070 (N_7070,N_4392,N_4417);
and U7071 (N_7071,N_3568,N_557);
nand U7072 (N_7072,N_3984,N_5585);
and U7073 (N_7073,N_2125,N_444);
and U7074 (N_7074,N_1829,N_3810);
or U7075 (N_7075,N_3505,N_1939);
or U7076 (N_7076,N_1995,N_5934);
nor U7077 (N_7077,N_3141,N_4243);
nand U7078 (N_7078,N_1446,N_4870);
nand U7079 (N_7079,N_4741,N_3744);
or U7080 (N_7080,N_3820,N_1032);
nor U7081 (N_7081,N_3900,N_5657);
xnor U7082 (N_7082,N_1497,N_3933);
and U7083 (N_7083,N_4695,N_4611);
xor U7084 (N_7084,N_2051,N_1141);
nor U7085 (N_7085,N_4289,N_4459);
or U7086 (N_7086,N_990,N_508);
or U7087 (N_7087,N_4095,N_3468);
nand U7088 (N_7088,N_4048,N_3047);
or U7089 (N_7089,N_2365,N_3499);
and U7090 (N_7090,N_4812,N_742);
nand U7091 (N_7091,N_1967,N_5908);
nand U7092 (N_7092,N_1172,N_2711);
or U7093 (N_7093,N_563,N_1383);
and U7094 (N_7094,N_3454,N_522);
and U7095 (N_7095,N_3078,N_2463);
nor U7096 (N_7096,N_2266,N_3754);
nand U7097 (N_7097,N_2007,N_2037);
and U7098 (N_7098,N_93,N_5484);
and U7099 (N_7099,N_3006,N_5007);
and U7100 (N_7100,N_1859,N_2877);
nor U7101 (N_7101,N_5174,N_404);
nor U7102 (N_7102,N_5122,N_6002);
or U7103 (N_7103,N_5135,N_3829);
nand U7104 (N_7104,N_4810,N_632);
nor U7105 (N_7105,N_1371,N_3442);
nor U7106 (N_7106,N_3280,N_3289);
and U7107 (N_7107,N_4108,N_4726);
and U7108 (N_7108,N_2376,N_4277);
nor U7109 (N_7109,N_1820,N_408);
or U7110 (N_7110,N_1115,N_2552);
nor U7111 (N_7111,N_6143,N_3119);
and U7112 (N_7112,N_828,N_556);
or U7113 (N_7113,N_4276,N_5853);
nand U7114 (N_7114,N_3827,N_6113);
or U7115 (N_7115,N_5342,N_2935);
nand U7116 (N_7116,N_1124,N_3899);
and U7117 (N_7117,N_2822,N_5186);
nand U7118 (N_7118,N_453,N_682);
nor U7119 (N_7119,N_1327,N_5480);
nor U7120 (N_7120,N_4328,N_4508);
and U7121 (N_7121,N_2733,N_1850);
nand U7122 (N_7122,N_6115,N_5250);
and U7123 (N_7123,N_2735,N_669);
and U7124 (N_7124,N_55,N_281);
nor U7125 (N_7125,N_1569,N_5435);
nor U7126 (N_7126,N_3170,N_5782);
and U7127 (N_7127,N_3286,N_5123);
nand U7128 (N_7128,N_1761,N_1593);
nor U7129 (N_7129,N_309,N_4172);
or U7130 (N_7130,N_1234,N_1257);
xor U7131 (N_7131,N_961,N_1179);
nor U7132 (N_7132,N_1747,N_4816);
or U7133 (N_7133,N_2417,N_3512);
xnor U7134 (N_7134,N_1751,N_162);
or U7135 (N_7135,N_3506,N_1297);
or U7136 (N_7136,N_1307,N_3712);
and U7137 (N_7137,N_4774,N_1168);
nor U7138 (N_7138,N_964,N_2805);
nor U7139 (N_7139,N_6049,N_1384);
or U7140 (N_7140,N_3130,N_5386);
or U7141 (N_7141,N_1459,N_1627);
and U7142 (N_7142,N_314,N_5586);
nand U7143 (N_7143,N_5602,N_2316);
nand U7144 (N_7144,N_3440,N_4353);
nand U7145 (N_7145,N_821,N_2254);
or U7146 (N_7146,N_2999,N_798);
or U7147 (N_7147,N_908,N_2461);
nor U7148 (N_7148,N_4623,N_685);
or U7149 (N_7149,N_464,N_1923);
nor U7150 (N_7150,N_4566,N_3542);
or U7151 (N_7151,N_2338,N_5712);
nand U7152 (N_7152,N_65,N_4092);
and U7153 (N_7153,N_2800,N_5409);
xor U7154 (N_7154,N_5605,N_3178);
or U7155 (N_7155,N_5850,N_274);
or U7156 (N_7156,N_2853,N_5450);
or U7157 (N_7157,N_2408,N_5637);
and U7158 (N_7158,N_2280,N_2290);
and U7159 (N_7159,N_5330,N_1688);
nor U7160 (N_7160,N_2684,N_594);
and U7161 (N_7161,N_957,N_4615);
nand U7162 (N_7162,N_4488,N_1235);
nand U7163 (N_7163,N_3452,N_1492);
or U7164 (N_7164,N_5408,N_2426);
nor U7165 (N_7165,N_2178,N_3833);
xnor U7166 (N_7166,N_5776,N_1649);
and U7167 (N_7167,N_3905,N_2414);
and U7168 (N_7168,N_5568,N_4420);
and U7169 (N_7169,N_4995,N_463);
nand U7170 (N_7170,N_5065,N_691);
nand U7171 (N_7171,N_5878,N_2911);
nand U7172 (N_7172,N_3710,N_1130);
or U7173 (N_7173,N_1199,N_1553);
or U7174 (N_7174,N_3268,N_5578);
nor U7175 (N_7175,N_5453,N_2857);
and U7176 (N_7176,N_4620,N_6158);
or U7177 (N_7177,N_4669,N_1046);
and U7178 (N_7178,N_4170,N_2173);
nand U7179 (N_7179,N_2567,N_5425);
xnor U7180 (N_7180,N_4455,N_3413);
nor U7181 (N_7181,N_3530,N_6148);
nor U7182 (N_7182,N_2404,N_4286);
nor U7183 (N_7183,N_6138,N_5646);
xnor U7184 (N_7184,N_134,N_3126);
and U7185 (N_7185,N_4590,N_4882);
nor U7186 (N_7186,N_6082,N_5798);
xnor U7187 (N_7187,N_5615,N_5468);
or U7188 (N_7188,N_4926,N_5978);
nand U7189 (N_7189,N_3199,N_3935);
or U7190 (N_7190,N_2237,N_4955);
xnor U7191 (N_7191,N_3773,N_2420);
nand U7192 (N_7192,N_5965,N_1450);
and U7193 (N_7193,N_1043,N_5416);
and U7194 (N_7194,N_4633,N_5818);
nor U7195 (N_7195,N_1190,N_6012);
or U7196 (N_7196,N_2409,N_5278);
and U7197 (N_7197,N_3397,N_5986);
nand U7198 (N_7198,N_5465,N_4013);
and U7199 (N_7199,N_4707,N_4545);
or U7200 (N_7200,N_1140,N_5852);
nor U7201 (N_7201,N_1337,N_4902);
and U7202 (N_7202,N_3236,N_4856);
or U7203 (N_7203,N_1377,N_5770);
xor U7204 (N_7204,N_6154,N_313);
and U7205 (N_7205,N_5136,N_1930);
or U7206 (N_7206,N_2556,N_5274);
and U7207 (N_7207,N_5789,N_1486);
nor U7208 (N_7208,N_2809,N_4665);
xnor U7209 (N_7209,N_4213,N_2768);
nor U7210 (N_7210,N_1613,N_4740);
nand U7211 (N_7211,N_981,N_5563);
nand U7212 (N_7212,N_3217,N_2525);
nor U7213 (N_7213,N_1807,N_1315);
nand U7214 (N_7214,N_6026,N_4512);
nor U7215 (N_7215,N_2089,N_5048);
or U7216 (N_7216,N_4729,N_6094);
and U7217 (N_7217,N_5115,N_1362);
xor U7218 (N_7218,N_5146,N_1650);
xor U7219 (N_7219,N_365,N_1605);
xnor U7220 (N_7220,N_3388,N_1044);
xnor U7221 (N_7221,N_1992,N_952);
nor U7222 (N_7222,N_4609,N_261);
nand U7223 (N_7223,N_4185,N_3718);
and U7224 (N_7224,N_2088,N_265);
nand U7225 (N_7225,N_6032,N_1471);
or U7226 (N_7226,N_5786,N_2364);
nor U7227 (N_7227,N_3430,N_2973);
and U7228 (N_7228,N_5460,N_3729);
or U7229 (N_7229,N_5717,N_4612);
xor U7230 (N_7230,N_3323,N_2840);
nand U7231 (N_7231,N_1886,N_2984);
nor U7232 (N_7232,N_4489,N_5784);
nor U7233 (N_7233,N_1836,N_5650);
nor U7234 (N_7234,N_3990,N_5011);
or U7235 (N_7235,N_3835,N_1325);
or U7236 (N_7236,N_5809,N_5317);
and U7237 (N_7237,N_3953,N_1239);
and U7238 (N_7238,N_3893,N_4785);
nand U7239 (N_7239,N_10,N_4778);
nand U7240 (N_7240,N_1456,N_5950);
nor U7241 (N_7241,N_2080,N_3679);
and U7242 (N_7242,N_3549,N_5777);
xor U7243 (N_7243,N_3402,N_4132);
xor U7244 (N_7244,N_5972,N_3043);
nand U7245 (N_7245,N_3765,N_3393);
and U7246 (N_7246,N_1323,N_2323);
and U7247 (N_7247,N_1273,N_4215);
and U7248 (N_7248,N_1094,N_5935);
or U7249 (N_7249,N_6117,N_874);
or U7250 (N_7250,N_6044,N_3376);
nand U7251 (N_7251,N_1480,N_648);
and U7252 (N_7252,N_2370,N_3225);
or U7253 (N_7253,N_3724,N_3408);
or U7254 (N_7254,N_5885,N_3697);
and U7255 (N_7255,N_4696,N_3955);
nor U7256 (N_7256,N_2885,N_4557);
nor U7257 (N_7257,N_5842,N_2696);
nand U7258 (N_7258,N_1903,N_3966);
nand U7259 (N_7259,N_2197,N_4465);
xor U7260 (N_7260,N_5138,N_2871);
and U7261 (N_7261,N_1111,N_5601);
xor U7262 (N_7262,N_5428,N_5636);
or U7263 (N_7263,N_1183,N_3348);
nand U7264 (N_7264,N_566,N_2626);
and U7265 (N_7265,N_5621,N_2050);
or U7266 (N_7266,N_1092,N_4257);
xor U7267 (N_7267,N_389,N_5101);
nor U7268 (N_7268,N_2015,N_4654);
nand U7269 (N_7269,N_3206,N_2677);
and U7270 (N_7270,N_3817,N_4619);
and U7271 (N_7271,N_6247,N_2071);
nand U7272 (N_7272,N_2568,N_5590);
and U7273 (N_7273,N_5920,N_2506);
and U7274 (N_7274,N_1874,N_1065);
and U7275 (N_7275,N_1565,N_3919);
nor U7276 (N_7276,N_2873,N_4507);
nor U7277 (N_7277,N_6237,N_554);
nand U7278 (N_7278,N_3357,N_3291);
and U7279 (N_7279,N_2727,N_2436);
nor U7280 (N_7280,N_1789,N_1568);
or U7281 (N_7281,N_3705,N_5082);
nand U7282 (N_7282,N_1589,N_461);
nand U7283 (N_7283,N_4191,N_1180);
or U7284 (N_7284,N_2772,N_4050);
nand U7285 (N_7285,N_1003,N_4381);
nor U7286 (N_7286,N_5959,N_5754);
nor U7287 (N_7287,N_406,N_5666);
nand U7288 (N_7288,N_3821,N_3655);
nand U7289 (N_7289,N_5245,N_1822);
and U7290 (N_7290,N_1691,N_730);
nand U7291 (N_7291,N_3582,N_3556);
or U7292 (N_7292,N_3001,N_3947);
and U7293 (N_7293,N_5137,N_2828);
xor U7294 (N_7294,N_5983,N_5739);
xor U7295 (N_7295,N_2910,N_4589);
nand U7296 (N_7296,N_2803,N_3489);
xor U7297 (N_7297,N_2557,N_3354);
and U7298 (N_7298,N_1123,N_6118);
or U7299 (N_7299,N_5476,N_3317);
xor U7300 (N_7300,N_4770,N_349);
nand U7301 (N_7301,N_455,N_2159);
nor U7302 (N_7302,N_625,N_5211);
nor U7303 (N_7303,N_2152,N_1192);
xnor U7304 (N_7304,N_4400,N_642);
or U7305 (N_7305,N_1618,N_2830);
nand U7306 (N_7306,N_2683,N_5113);
or U7307 (N_7307,N_3511,N_3020);
and U7308 (N_7308,N_2148,N_4648);
and U7309 (N_7309,N_11,N_3128);
nand U7310 (N_7310,N_1653,N_2747);
nand U7311 (N_7311,N_2117,N_2730);
nor U7312 (N_7312,N_4292,N_5255);
nor U7313 (N_7313,N_1054,N_3518);
nor U7314 (N_7314,N_581,N_4748);
nand U7315 (N_7315,N_4836,N_3456);
nor U7316 (N_7316,N_1978,N_457);
and U7317 (N_7317,N_1952,N_4766);
nor U7318 (N_7318,N_3095,N_3099);
and U7319 (N_7319,N_4934,N_36);
nor U7320 (N_7320,N_2752,N_5728);
nand U7321 (N_7321,N_1061,N_6124);
nor U7322 (N_7322,N_1764,N_4985);
and U7323 (N_7323,N_393,N_5760);
nand U7324 (N_7324,N_1008,N_2497);
and U7325 (N_7325,N_6007,N_4349);
xor U7326 (N_7326,N_86,N_1643);
nor U7327 (N_7327,N_5116,N_3240);
or U7328 (N_7328,N_4120,N_1212);
nand U7329 (N_7329,N_1267,N_6015);
nand U7330 (N_7330,N_761,N_1921);
nor U7331 (N_7331,N_3085,N_3769);
nor U7332 (N_7332,N_179,N_1466);
or U7333 (N_7333,N_611,N_2260);
nand U7334 (N_7334,N_57,N_5841);
nor U7335 (N_7335,N_6139,N_950);
and U7336 (N_7336,N_2953,N_1980);
nand U7337 (N_7337,N_4316,N_483);
xnor U7338 (N_7338,N_4699,N_4920);
and U7339 (N_7339,N_2158,N_5577);
nand U7340 (N_7340,N_1103,N_288);
xnor U7341 (N_7341,N_654,N_3192);
nor U7342 (N_7342,N_174,N_5971);
xor U7343 (N_7343,N_5955,N_5763);
nand U7344 (N_7344,N_3785,N_2096);
and U7345 (N_7345,N_471,N_5795);
or U7346 (N_7346,N_3982,N_1503);
nand U7347 (N_7347,N_4602,N_5663);
or U7348 (N_7348,N_3190,N_1104);
xor U7349 (N_7349,N_5402,N_6187);
and U7350 (N_7350,N_635,N_3602);
xor U7351 (N_7351,N_3708,N_5702);
xnor U7352 (N_7352,N_2968,N_1350);
or U7353 (N_7353,N_3181,N_3134);
and U7354 (N_7354,N_3862,N_5190);
or U7355 (N_7355,N_3741,N_512);
nand U7356 (N_7356,N_748,N_4158);
nor U7357 (N_7357,N_4466,N_3678);
and U7358 (N_7358,N_4456,N_1211);
and U7359 (N_7359,N_4644,N_1105);
nand U7360 (N_7360,N_5580,N_6234);
nand U7361 (N_7361,N_3463,N_109);
nor U7362 (N_7362,N_2047,N_4338);
and U7363 (N_7363,N_2078,N_3650);
nor U7364 (N_7364,N_1272,N_5838);
and U7365 (N_7365,N_347,N_1074);
and U7366 (N_7366,N_1647,N_6181);
nor U7367 (N_7367,N_3033,N_4561);
nor U7368 (N_7368,N_2812,N_782);
nand U7369 (N_7369,N_3707,N_3282);
and U7370 (N_7370,N_5525,N_6198);
and U7371 (N_7371,N_5185,N_1665);
nand U7372 (N_7372,N_4607,N_1961);
nor U7373 (N_7373,N_4007,N_5144);
xnor U7374 (N_7374,N_4938,N_4628);
nand U7375 (N_7375,N_3155,N_712);
xor U7376 (N_7376,N_100,N_871);
xnor U7377 (N_7377,N_2072,N_2582);
nand U7378 (N_7378,N_2003,N_5028);
and U7379 (N_7379,N_138,N_2921);
or U7380 (N_7380,N_958,N_1722);
and U7381 (N_7381,N_805,N_133);
and U7382 (N_7382,N_3992,N_2964);
nor U7383 (N_7383,N_596,N_1378);
or U7384 (N_7384,N_788,N_5426);
nor U7385 (N_7385,N_4231,N_569);
nor U7386 (N_7386,N_3552,N_3675);
xnor U7387 (N_7387,N_3313,N_2608);
nand U7388 (N_7388,N_2966,N_577);
or U7389 (N_7389,N_6146,N_5839);
xor U7390 (N_7390,N_692,N_1861);
nand U7391 (N_7391,N_2687,N_4805);
and U7392 (N_7392,N_4742,N_5075);
nor U7393 (N_7393,N_1314,N_1262);
and U7394 (N_7394,N_4003,N_1441);
and U7395 (N_7395,N_4884,N_4880);
nand U7396 (N_7396,N_54,N_3976);
or U7397 (N_7397,N_268,N_22);
nand U7398 (N_7398,N_5638,N_5980);
nand U7399 (N_7399,N_1039,N_1870);
and U7400 (N_7400,N_3686,N_838);
nor U7401 (N_7401,N_3337,N_3218);
and U7402 (N_7402,N_2176,N_2102);
nor U7403 (N_7403,N_4911,N_4772);
xor U7404 (N_7404,N_5046,N_2258);
or U7405 (N_7405,N_3871,N_1740);
xor U7406 (N_7406,N_1298,N_71);
nor U7407 (N_7407,N_3637,N_155);
or U7408 (N_7408,N_509,N_1760);
or U7409 (N_7409,N_3367,N_4799);
and U7410 (N_7410,N_423,N_3799);
nor U7411 (N_7411,N_5593,N_745);
xnor U7412 (N_7412,N_2754,N_5483);
and U7413 (N_7413,N_3433,N_2179);
or U7414 (N_7414,N_818,N_5775);
and U7415 (N_7415,N_2806,N_5559);
nor U7416 (N_7416,N_3372,N_5875);
and U7417 (N_7417,N_4850,N_1455);
nor U7418 (N_7418,N_6242,N_962);
and U7419 (N_7419,N_3653,N_1200);
nand U7420 (N_7420,N_4306,N_2824);
nand U7421 (N_7421,N_4200,N_1857);
nor U7422 (N_7422,N_3320,N_2859);
xnor U7423 (N_7423,N_3647,N_3153);
nor U7424 (N_7424,N_2363,N_1631);
nor U7425 (N_7425,N_4222,N_4553);
or U7426 (N_7426,N_3262,N_5105);
nor U7427 (N_7427,N_1236,N_5332);
and U7428 (N_7428,N_693,N_4977);
xor U7429 (N_7429,N_963,N_794);
or U7430 (N_7430,N_1324,N_320);
nor U7431 (N_7431,N_3273,N_3776);
nand U7432 (N_7432,N_4887,N_1915);
nor U7433 (N_7433,N_5692,N_6168);
nand U7434 (N_7434,N_5562,N_1531);
nor U7435 (N_7435,N_4671,N_984);
nand U7436 (N_7436,N_1025,N_5688);
nand U7437 (N_7437,N_1432,N_6);
or U7438 (N_7438,N_251,N_356);
or U7439 (N_7439,N_2948,N_3526);
or U7440 (N_7440,N_5340,N_1475);
nor U7441 (N_7441,N_3396,N_5177);
xnor U7442 (N_7442,N_559,N_3312);
or U7443 (N_7443,N_4187,N_4299);
or U7444 (N_7444,N_5253,N_1772);
or U7445 (N_7445,N_989,N_5805);
or U7446 (N_7446,N_6040,N_5297);
nand U7447 (N_7447,N_2495,N_1501);
and U7448 (N_7448,N_1076,N_1138);
and U7449 (N_7449,N_3560,N_3215);
and U7450 (N_7450,N_4333,N_1621);
and U7451 (N_7451,N_2581,N_4116);
nand U7452 (N_7452,N_4281,N_2192);
or U7453 (N_7453,N_591,N_3404);
and U7454 (N_7454,N_394,N_5609);
nand U7455 (N_7455,N_4122,N_4967);
nand U7456 (N_7456,N_1678,N_5314);
and U7457 (N_7457,N_1985,N_405);
xor U7458 (N_7458,N_4473,N_158);
and U7459 (N_7459,N_5498,N_1413);
xnor U7460 (N_7460,N_4188,N_2470);
and U7461 (N_7461,N_3296,N_3295);
nor U7462 (N_7462,N_1805,N_1936);
and U7463 (N_7463,N_6197,N_5985);
and U7464 (N_7464,N_4457,N_2262);
and U7465 (N_7465,N_2956,N_2236);
xnor U7466 (N_7466,N_1924,N_1767);
nor U7467 (N_7467,N_3531,N_2798);
or U7468 (N_7468,N_3443,N_473);
or U7469 (N_7469,N_5918,N_5924);
or U7470 (N_7470,N_6218,N_4388);
nand U7471 (N_7471,N_194,N_3333);
nand U7472 (N_7472,N_5627,N_3898);
and U7473 (N_7473,N_5431,N_1524);
nand U7474 (N_7474,N_2590,N_160);
nand U7475 (N_7475,N_530,N_2980);
xnor U7476 (N_7476,N_5320,N_2405);
and U7477 (N_7477,N_1494,N_5998);
nand U7478 (N_7478,N_4056,N_4492);
and U7479 (N_7479,N_1525,N_5305);
xor U7480 (N_7480,N_4100,N_2279);
xor U7481 (N_7481,N_4250,N_5703);
nand U7482 (N_7482,N_5964,N_6006);
or U7483 (N_7483,N_4548,N_699);
and U7484 (N_7484,N_3426,N_2972);
nand U7485 (N_7485,N_5925,N_786);
nand U7486 (N_7486,N_3948,N_2748);
nor U7487 (N_7487,N_5941,N_3235);
or U7488 (N_7488,N_5519,N_1982);
and U7489 (N_7489,N_849,N_6031);
xnor U7490 (N_7490,N_1230,N_655);
and U7491 (N_7491,N_3260,N_3855);
nor U7492 (N_7492,N_4431,N_1393);
and U7493 (N_7493,N_3036,N_5088);
nand U7494 (N_7494,N_813,N_1938);
nor U7495 (N_7495,N_4065,N_4330);
nor U7496 (N_7496,N_6106,N_2659);
nand U7497 (N_7497,N_2228,N_2740);
and U7498 (N_7498,N_2421,N_4657);
nand U7499 (N_7499,N_3750,N_926);
and U7500 (N_7500,N_3242,N_564);
or U7501 (N_7501,N_5272,N_2738);
and U7502 (N_7502,N_4511,N_4960);
and U7503 (N_7503,N_715,N_5501);
xor U7504 (N_7504,N_4532,N_904);
and U7505 (N_7505,N_3790,N_2892);
nand U7506 (N_7506,N_5072,N_510);
or U7507 (N_7507,N_597,N_258);
or U7508 (N_7508,N_1630,N_1987);
nand U7509 (N_7509,N_4348,N_4647);
or U7510 (N_7510,N_4932,N_647);
nand U7511 (N_7511,N_5001,N_1790);
and U7512 (N_7512,N_4263,N_5106);
and U7513 (N_7513,N_4370,N_2012);
xnor U7514 (N_7514,N_4746,N_4037);
or U7515 (N_7515,N_3231,N_4090);
and U7516 (N_7516,N_1160,N_276);
xor U7517 (N_7517,N_729,N_2780);
nor U7518 (N_7518,N_5573,N_1608);
and U7519 (N_7519,N_1581,N_1991);
and U7520 (N_7520,N_754,N_4067);
or U7521 (N_7521,N_3389,N_3694);
nand U7522 (N_7522,N_5547,N_3185);
and U7523 (N_7523,N_1758,N_4881);
nand U7524 (N_7524,N_2555,N_4093);
nor U7525 (N_7525,N_2990,N_4780);
nor U7526 (N_7526,N_3158,N_3672);
and U7527 (N_7527,N_599,N_4421);
nand U7528 (N_7528,N_5108,N_5471);
nor U7529 (N_7529,N_5882,N_5430);
and U7530 (N_7530,N_1518,N_5189);
or U7531 (N_7531,N_5389,N_909);
or U7532 (N_7532,N_1108,N_542);
xor U7533 (N_7533,N_3840,N_4113);
xnor U7534 (N_7534,N_4207,N_644);
and U7535 (N_7535,N_1651,N_2895);
or U7536 (N_7536,N_181,N_3859);
nand U7537 (N_7537,N_4725,N_1727);
nor U7538 (N_7538,N_921,N_2356);
nand U7539 (N_7539,N_4262,N_4653);
nand U7540 (N_7540,N_6125,N_2517);
or U7541 (N_7541,N_3676,N_5455);
nand U7542 (N_7542,N_3248,N_3626);
and U7543 (N_7543,N_5304,N_3805);
or U7544 (N_7544,N_3361,N_2432);
or U7545 (N_7545,N_4586,N_6184);
or U7546 (N_7546,N_1019,N_3850);
or U7547 (N_7547,N_6114,N_5939);
nor U7548 (N_7548,N_6079,N_1957);
and U7549 (N_7549,N_3105,N_1476);
nor U7550 (N_7550,N_2845,N_5507);
nand U7551 (N_7551,N_2742,N_1920);
or U7552 (N_7552,N_2396,N_5988);
and U7553 (N_7553,N_1506,N_4309);
and U7554 (N_7554,N_1133,N_254);
nand U7555 (N_7555,N_2223,N_5899);
nand U7556 (N_7556,N_1825,N_700);
nand U7557 (N_7557,N_1775,N_3241);
xnor U7558 (N_7558,N_5341,N_3405);
or U7559 (N_7559,N_743,N_3946);
nor U7560 (N_7560,N_3324,N_1910);
nand U7561 (N_7561,N_3439,N_4287);
and U7562 (N_7562,N_2739,N_5811);
nor U7563 (N_7563,N_4382,N_4427);
or U7564 (N_7564,N_1246,N_5870);
nor U7565 (N_7565,N_1661,N_5268);
or U7566 (N_7566,N_3303,N_4767);
nand U7567 (N_7567,N_3803,N_1880);
nor U7568 (N_7568,N_2029,N_5889);
nor U7569 (N_7569,N_1687,N_4425);
nand U7570 (N_7570,N_6142,N_5785);
and U7571 (N_7571,N_2751,N_2450);
or U7572 (N_7572,N_3283,N_334);
nor U7573 (N_7573,N_4490,N_2701);
or U7574 (N_7574,N_2989,N_306);
nor U7575 (N_7575,N_3516,N_934);
and U7576 (N_7576,N_3202,N_2163);
or U7577 (N_7577,N_6233,N_3832);
nand U7578 (N_7578,N_257,N_5658);
nand U7579 (N_7579,N_2725,N_4291);
or U7580 (N_7580,N_422,N_2635);
nor U7581 (N_7581,N_3870,N_3418);
and U7582 (N_7582,N_806,N_2534);
and U7583 (N_7583,N_5345,N_39);
and U7584 (N_7584,N_3385,N_2898);
nand U7585 (N_7585,N_4127,N_2922);
or U7586 (N_7586,N_1814,N_578);
nand U7587 (N_7587,N_5085,N_942);
xnor U7588 (N_7588,N_5653,N_4265);
or U7589 (N_7589,N_4040,N_662);
nor U7590 (N_7590,N_3088,N_4629);
nor U7591 (N_7591,N_5130,N_1049);
nand U7592 (N_7592,N_882,N_490);
nor U7593 (N_7593,N_2603,N_3034);
nand U7594 (N_7594,N_3279,N_3734);
nand U7595 (N_7595,N_5967,N_1063);
or U7596 (N_7596,N_5280,N_2634);
xnor U7597 (N_7597,N_1385,N_277);
and U7598 (N_7598,N_5153,N_1394);
and U7599 (N_7599,N_3054,N_832);
and U7600 (N_7600,N_1255,N_4670);
nand U7601 (N_7601,N_2473,N_3267);
or U7602 (N_7602,N_1000,N_5803);
nand U7603 (N_7603,N_5025,N_3706);
xnor U7604 (N_7604,N_2348,N_16);
nor U7605 (N_7605,N_5729,N_6064);
xor U7606 (N_7606,N_2535,N_3996);
nand U7607 (N_7607,N_92,N_6246);
and U7608 (N_7608,N_5201,N_219);
nor U7609 (N_7609,N_6089,N_4110);
nand U7610 (N_7610,N_1728,N_2804);
or U7611 (N_7611,N_6201,N_336);
or U7612 (N_7612,N_814,N_1280);
or U7613 (N_7613,N_2598,N_2449);
nor U7614 (N_7614,N_1493,N_1667);
xor U7615 (N_7615,N_2489,N_2920);
nand U7616 (N_7616,N_4146,N_5907);
or U7617 (N_7617,N_2064,N_976);
or U7618 (N_7618,N_2993,N_5753);
or U7619 (N_7619,N_4582,N_4436);
or U7620 (N_7620,N_3157,N_2757);
nor U7621 (N_7621,N_1607,N_5814);
or U7622 (N_7622,N_878,N_3288);
nor U7623 (N_7623,N_5418,N_5143);
nor U7624 (N_7624,N_3501,N_4428);
nor U7625 (N_7625,N_491,N_3874);
nor U7626 (N_7626,N_4789,N_978);
nand U7627 (N_7627,N_2866,N_4407);
nor U7628 (N_7628,N_864,N_4148);
nand U7629 (N_7629,N_6235,N_5566);
nor U7630 (N_7630,N_3432,N_4171);
nor U7631 (N_7631,N_238,N_5419);
or U7632 (N_7632,N_2043,N_6157);
or U7633 (N_7633,N_1842,N_3083);
nand U7634 (N_7634,N_4617,N_3136);
and U7635 (N_7635,N_959,N_1934);
nand U7636 (N_7636,N_3520,N_533);
or U7637 (N_7637,N_4543,N_3778);
xor U7638 (N_7638,N_1547,N_1436);
and U7639 (N_7639,N_1641,N_4574);
nor U7640 (N_7640,N_3514,N_3058);
nand U7641 (N_7641,N_2958,N_3667);
and U7642 (N_7642,N_296,N_1322);
nor U7643 (N_7643,N_3671,N_1749);
or U7644 (N_7644,N_3090,N_4814);
nor U7645 (N_7645,N_5234,N_980);
nor U7646 (N_7646,N_3657,N_503);
nor U7647 (N_7647,N_735,N_1552);
nor U7648 (N_7648,N_4854,N_2624);
and U7649 (N_7649,N_3476,N_144);
nand U7650 (N_7650,N_5864,N_734);
nor U7651 (N_7651,N_4900,N_5669);
or U7652 (N_7652,N_5759,N_70);
nor U7653 (N_7653,N_4403,N_5672);
or U7654 (N_7654,N_2869,N_6200);
or U7655 (N_7655,N_1006,N_4575);
and U7656 (N_7656,N_2359,N_6020);
nor U7657 (N_7657,N_2524,N_4600);
and U7658 (N_7658,N_5708,N_1507);
nand U7659 (N_7659,N_1072,N_3309);
nor U7660 (N_7660,N_2360,N_2465);
nor U7661 (N_7661,N_6048,N_2313);
and U7662 (N_7662,N_5180,N_385);
nor U7663 (N_7663,N_1574,N_203);
nor U7664 (N_7664,N_1906,N_5634);
nor U7665 (N_7665,N_1882,N_3826);
and U7666 (N_7666,N_38,N_3092);
or U7667 (N_7667,N_1304,N_1919);
nand U7668 (N_7668,N_4178,N_696);
nor U7669 (N_7669,N_1313,N_2794);
nor U7670 (N_7670,N_3949,N_1823);
nand U7671 (N_7671,N_1068,N_4284);
nor U7672 (N_7672,N_3046,N_4538);
or U7673 (N_7673,N_4838,N_4562);
and U7674 (N_7674,N_824,N_3749);
nor U7675 (N_7675,N_3923,N_3160);
nand U7676 (N_7676,N_5264,N_3759);
and U7677 (N_7677,N_1059,N_135);
and U7678 (N_7678,N_5166,N_5347);
nor U7679 (N_7679,N_4556,N_4112);
nor U7680 (N_7680,N_4248,N_1887);
and U7681 (N_7681,N_2694,N_701);
nand U7682 (N_7682,N_2591,N_836);
or U7683 (N_7683,N_5806,N_1089);
xor U7684 (N_7684,N_469,N_3214);
nand U7685 (N_7685,N_1791,N_1474);
xor U7686 (N_7686,N_2493,N_8);
nor U7687 (N_7687,N_2621,N_4570);
xor U7688 (N_7688,N_702,N_156);
nor U7689 (N_7689,N_1800,N_2549);
xnor U7690 (N_7690,N_3365,N_2998);
nand U7691 (N_7691,N_3986,N_2184);
or U7692 (N_7692,N_511,N_4406);
nor U7693 (N_7693,N_363,N_901);
xor U7694 (N_7694,N_5241,N_4689);
or U7695 (N_7695,N_2115,N_3193);
or U7696 (N_7696,N_4009,N_724);
and U7697 (N_7697,N_384,N_1066);
nand U7698 (N_7698,N_493,N_785);
nor U7699 (N_7699,N_3486,N_2971);
or U7700 (N_7700,N_697,N_3703);
and U7701 (N_7701,N_6215,N_3258);
nand U7702 (N_7702,N_207,N_2601);
and U7703 (N_7703,N_4096,N_975);
xnor U7704 (N_7704,N_1110,N_7);
or U7705 (N_7705,N_4996,N_2353);
nor U7706 (N_7706,N_3373,N_1545);
nor U7707 (N_7707,N_5026,N_3618);
nor U7708 (N_7708,N_1774,N_1415);
and U7709 (N_7709,N_4970,N_2629);
or U7710 (N_7710,N_1129,N_2160);
and U7711 (N_7711,N_5822,N_4974);
nor U7712 (N_7712,N_1534,N_4347);
nor U7713 (N_7713,N_972,N_4021);
nor U7714 (N_7714,N_1012,N_2222);
or U7715 (N_7715,N_4876,N_1271);
and U7716 (N_7716,N_243,N_2300);
xnor U7717 (N_7717,N_4154,N_3693);
nand U7718 (N_7718,N_1595,N_308);
and U7719 (N_7719,N_2032,N_3910);
nand U7720 (N_7720,N_1403,N_1334);
xor U7721 (N_7721,N_1588,N_5401);
nand U7722 (N_7722,N_2216,N_1673);
nor U7723 (N_7723,N_3875,N_5291);
nand U7724 (N_7724,N_4786,N_5300);
nand U7725 (N_7725,N_3469,N_2960);
or U7726 (N_7726,N_6081,N_5504);
and U7727 (N_7727,N_5682,N_6059);
and U7728 (N_7728,N_141,N_4981);
xnor U7729 (N_7729,N_5248,N_5243);
or U7730 (N_7730,N_2053,N_3533);
nor U7731 (N_7731,N_1634,N_459);
nand U7732 (N_7732,N_550,N_1232);
or U7733 (N_7733,N_4596,N_5041);
or U7734 (N_7734,N_3881,N_4412);
and U7735 (N_7735,N_3319,N_3395);
xor U7736 (N_7736,N_5990,N_5246);
and U7737 (N_7737,N_2099,N_1354);
xor U7738 (N_7738,N_338,N_945);
nor U7739 (N_7739,N_3599,N_2773);
nor U7740 (N_7740,N_987,N_3492);
nand U7741 (N_7741,N_434,N_3937);
and U7742 (N_7742,N_5858,N_4305);
nand U7743 (N_7743,N_1028,N_5441);
xor U7744 (N_7744,N_6102,N_891);
or U7745 (N_7745,N_31,N_2903);
xor U7746 (N_7746,N_176,N_5353);
or U7747 (N_7747,N_4130,N_2406);
or U7748 (N_7748,N_1734,N_5393);
or U7749 (N_7749,N_1769,N_5665);
and U7750 (N_7750,N_2538,N_468);
nand U7751 (N_7751,N_1055,N_2215);
and U7752 (N_7752,N_4460,N_5893);
nor U7753 (N_7753,N_855,N_3265);
nand U7754 (N_7754,N_5629,N_3308);
nand U7755 (N_7755,N_1975,N_1626);
xor U7756 (N_7756,N_2055,N_1427);
or U7757 (N_7757,N_6093,N_4580);
nor U7758 (N_7758,N_5125,N_3930);
nand U7759 (N_7759,N_5279,N_3460);
nand U7760 (N_7760,N_6248,N_5308);
and U7761 (N_7761,N_185,N_3077);
nand U7762 (N_7762,N_6153,N_1878);
nand U7763 (N_7763,N_4246,N_4572);
xnor U7764 (N_7764,N_4958,N_2269);
nand U7765 (N_7765,N_2715,N_3666);
nor U7766 (N_7766,N_1259,N_3037);
nand U7767 (N_7767,N_2383,N_4462);
nor U7768 (N_7768,N_1406,N_5905);
or U7769 (N_7769,N_5454,N_303);
and U7770 (N_7770,N_943,N_3885);
nand U7771 (N_7771,N_428,N_2382);
and U7772 (N_7772,N_3226,N_847);
nand U7773 (N_7773,N_3057,N_6211);
xor U7774 (N_7774,N_3359,N_6224);
nand U7775 (N_7775,N_1318,N_1811);
nor U7776 (N_7776,N_2614,N_1279);
or U7777 (N_7777,N_4181,N_776);
and U7778 (N_7778,N_354,N_3674);
nor U7779 (N_7779,N_4461,N_4680);
or U7780 (N_7780,N_4280,N_6167);
nor U7781 (N_7781,N_6112,N_3857);
nor U7782 (N_7782,N_3366,N_2856);
xor U7783 (N_7783,N_5755,N_2679);
nor U7784 (N_7784,N_5415,N_3256);
and U7785 (N_7785,N_2357,N_5398);
xnor U7786 (N_7786,N_5394,N_5846);
nand U7787 (N_7787,N_2983,N_4831);
and U7788 (N_7788,N_2116,N_1620);
xor U7789 (N_7789,N_4893,N_4874);
nand U7790 (N_7790,N_5718,N_4371);
and U7791 (N_7791,N_2834,N_4205);
or U7792 (N_7792,N_3502,N_3251);
and U7793 (N_7793,N_3931,N_2675);
and U7794 (N_7794,N_5413,N_5444);
nor U7795 (N_7795,N_2411,N_439);
or U7796 (N_7796,N_4555,N_1577);
and U7797 (N_7797,N_5448,N_5200);
and U7798 (N_7798,N_1929,N_2610);
and U7799 (N_7799,N_903,N_1373);
nand U7800 (N_7800,N_2508,N_3659);
and U7801 (N_7801,N_3521,N_1312);
nand U7802 (N_7802,N_1276,N_1196);
xor U7803 (N_7803,N_502,N_1872);
xor U7804 (N_7804,N_2526,N_703);
xnor U7805 (N_7805,N_2074,N_5569);
nor U7806 (N_7806,N_409,N_5595);
nand U7807 (N_7807,N_3051,N_1511);
nor U7808 (N_7808,N_4972,N_1237);
and U7809 (N_7809,N_3346,N_3007);
nor U7810 (N_7810,N_5461,N_172);
nand U7811 (N_7811,N_2499,N_3704);
nor U7812 (N_7812,N_1513,N_2095);
nor U7813 (N_7813,N_504,N_5076);
or U7814 (N_7814,N_4118,N_2387);
or U7815 (N_7815,N_2585,N_6092);
and U7816 (N_7816,N_2090,N_4070);
or U7817 (N_7817,N_2899,N_854);
xnor U7818 (N_7818,N_5716,N_3188);
and U7819 (N_7819,N_5499,N_4662);
nor U7820 (N_7820,N_5133,N_2656);
nand U7821 (N_7821,N_3728,N_837);
nand U7822 (N_7822,N_5331,N_1248);
and U7823 (N_7823,N_4168,N_3232);
nor U7824 (N_7824,N_2494,N_3490);
or U7825 (N_7825,N_182,N_21);
nor U7826 (N_7826,N_2350,N_1146);
nor U7827 (N_7827,N_4033,N_856);
and U7828 (N_7828,N_101,N_3740);
and U7829 (N_7829,N_4848,N_5596);
nor U7830 (N_7830,N_290,N_2602);
and U7831 (N_7831,N_638,N_351);
nor U7832 (N_7832,N_5992,N_4520);
nor U7833 (N_7833,N_2609,N_1782);
or U7834 (N_7834,N_3108,N_5457);
xor U7835 (N_7835,N_2240,N_5463);
nand U7836 (N_7836,N_4692,N_2959);
and U7837 (N_7837,N_3742,N_3714);
and U7838 (N_7838,N_4703,N_4272);
nor U7839 (N_7839,N_2397,N_1287);
and U7840 (N_7840,N_5301,N_3407);
nor U7841 (N_7841,N_6131,N_1721);
and U7842 (N_7842,N_292,N_1210);
or U7843 (N_7843,N_3210,N_985);
nor U7844 (N_7844,N_4396,N_1328);
or U7845 (N_7845,N_1093,N_4823);
or U7846 (N_7846,N_6033,N_5742);
or U7847 (N_7847,N_1966,N_3132);
nor U7848 (N_7848,N_3353,N_1320);
nand U7849 (N_7849,N_1424,N_1864);
and U7850 (N_7850,N_988,N_4672);
nand U7851 (N_7851,N_4509,N_4470);
nor U7852 (N_7852,N_1244,N_1763);
and U7853 (N_7853,N_4408,N_230);
nor U7854 (N_7854,N_5421,N_2782);
and U7855 (N_7855,N_2451,N_3538);
or U7856 (N_7856,N_4173,N_869);
or U7857 (N_7857,N_5429,N_2334);
xnor U7858 (N_7858,N_204,N_5553);
nor U7859 (N_7859,N_1904,N_1719);
or U7860 (N_7860,N_421,N_3853);
or U7861 (N_7861,N_3238,N_3738);
nand U7862 (N_7862,N_342,N_4475);
or U7863 (N_7863,N_1783,N_5608);
or U7864 (N_7864,N_2472,N_3597);
xor U7865 (N_7865,N_2446,N_3249);
and U7866 (N_7866,N_1841,N_1622);
nor U7867 (N_7867,N_1576,N_6136);
nand U7868 (N_7868,N_4445,N_840);
xnor U7869 (N_7869,N_3049,N_5128);
or U7870 (N_7870,N_4196,N_2548);
nor U7871 (N_7871,N_5991,N_5118);
nand U7872 (N_7872,N_1445,N_193);
nand U7873 (N_7873,N_4294,N_4712);
nor U7874 (N_7874,N_5903,N_861);
nor U7875 (N_7875,N_4530,N_4182);
nand U7876 (N_7876,N_2010,N_4835);
and U7877 (N_7877,N_136,N_6203);
or U7878 (N_7878,N_420,N_143);
nor U7879 (N_7879,N_2627,N_5024);
or U7880 (N_7880,N_5018,N_3684);
or U7881 (N_7881,N_5673,N_58);
nand U7882 (N_7882,N_999,N_4819);
nor U7883 (N_7883,N_720,N_4020);
nor U7884 (N_7884,N_1852,N_2996);
nor U7885 (N_7885,N_436,N_528);
or U7886 (N_7886,N_1340,N_6209);
and U7887 (N_7887,N_5475,N_5912);
nor U7888 (N_7888,N_4851,N_482);
xnor U7889 (N_7889,N_2650,N_1776);
or U7890 (N_7890,N_2784,N_2285);
and U7891 (N_7891,N_2849,N_1254);
nand U7892 (N_7892,N_5855,N_2041);
and U7893 (N_7893,N_3633,N_479);
nand U7894 (N_7894,N_5299,N_4804);
nand U7895 (N_7895,N_5951,N_800);
nand U7896 (N_7896,N_1932,N_95);
and U7897 (N_7897,N_1680,N_5778);
nor U7898 (N_7898,N_6077,N_2393);
and U7899 (N_7899,N_4091,N_973);
and U7900 (N_7900,N_3802,N_1695);
and U7901 (N_7901,N_1171,N_5975);
nand U7902 (N_7902,N_3447,N_4546);
nand U7903 (N_7903,N_2419,N_5256);
nor U7904 (N_7904,N_2760,N_4498);
nand U7905 (N_7905,N_2837,N_643);
nor U7906 (N_7906,N_3592,N_3216);
nor U7907 (N_7907,N_5302,N_1848);
or U7908 (N_7908,N_1462,N_72);
and U7909 (N_7909,N_2688,N_3720);
or U7910 (N_7910,N_4125,N_4704);
nor U7911 (N_7911,N_2185,N_5738);
nand U7912 (N_7912,N_868,N_1366);
or U7913 (N_7913,N_6245,N_4071);
or U7914 (N_7914,N_3182,N_3656);
nand U7915 (N_7915,N_2384,N_4554);
xor U7916 (N_7916,N_1205,N_4242);
nor U7917 (N_7917,N_4950,N_5094);
nand U7918 (N_7918,N_5266,N_3562);
nand U7919 (N_7919,N_2434,N_4723);
nand U7920 (N_7920,N_4046,N_1443);
and U7921 (N_7921,N_5321,N_9);
and U7922 (N_7922,N_4103,N_6171);
or U7923 (N_7923,N_6105,N_5667);
nand U7924 (N_7924,N_5382,N_5449);
or U7925 (N_7925,N_4713,N_472);
xnor U7926 (N_7926,N_4558,N_2142);
nor U7927 (N_7927,N_810,N_431);
and U7928 (N_7928,N_5854,N_2734);
nand U7929 (N_7929,N_1326,N_996);
nor U7930 (N_7930,N_291,N_2858);
nor U7931 (N_7931,N_4922,N_319);
nand U7932 (N_7932,N_3424,N_918);
xor U7933 (N_7933,N_4252,N_5751);
nand U7934 (N_7934,N_6108,N_1290);
and U7935 (N_7935,N_1964,N_5424);
and U7936 (N_7936,N_3109,N_4818);
nand U7937 (N_7937,N_1243,N_227);
or U7938 (N_7938,N_501,N_5473);
and U7939 (N_7939,N_2438,N_225);
or U7940 (N_7940,N_2392,N_4969);
nand U7941 (N_7941,N_1029,N_4759);
or U7942 (N_7942,N_3617,N_25);
nor U7943 (N_7943,N_4413,N_4369);
and U7944 (N_7944,N_2301,N_2902);
nor U7945 (N_7945,N_190,N_3873);
nor U7946 (N_7946,N_5233,N_5257);
nor U7947 (N_7947,N_4588,N_6150);
nand U7948 (N_7948,N_5923,N_4375);
nor U7949 (N_7949,N_3453,N_4494);
nor U7950 (N_7950,N_2373,N_2690);
nand U7951 (N_7951,N_684,N_4937);
nor U7952 (N_7952,N_4775,N_749);
and U7953 (N_7953,N_1733,N_5388);
nor U7954 (N_7954,N_1571,N_4474);
or U7955 (N_7955,N_4430,N_4346);
or U7956 (N_7956,N_3640,N_130);
nor U7957 (N_7957,N_3660,N_2049);
and U7958 (N_7958,N_1188,N_4988);
nor U7959 (N_7959,N_1095,N_1405);
or U7960 (N_7960,N_6191,N_4404);
and U7961 (N_7961,N_152,N_150);
nor U7962 (N_7962,N_5598,N_2657);
or U7963 (N_7963,N_2154,N_5378);
nor U7964 (N_7964,N_125,N_5987);
nand U7965 (N_7965,N_6024,N_3978);
nand U7966 (N_7966,N_4260,N_4271);
and U7967 (N_7967,N_1624,N_6069);
or U7968 (N_7968,N_2759,N_4907);
nand U7969 (N_7969,N_2038,N_4595);
and U7970 (N_7970,N_494,N_582);
and U7971 (N_7971,N_6192,N_5030);
nand U7972 (N_7972,N_1564,N_562);
or U7973 (N_7973,N_1365,N_2063);
and U7974 (N_7974,N_1937,N_5387);
or U7975 (N_7975,N_3509,N_443);
nand U7976 (N_7976,N_1107,N_5719);
nand U7977 (N_7977,N_5783,N_4279);
xor U7978 (N_7978,N_4085,N_2195);
xor U7979 (N_7979,N_4779,N_3121);
or U7980 (N_7980,N_3772,N_621);
nor U7981 (N_7981,N_652,N_6170);
or U7982 (N_7982,N_3311,N_5698);
nand U7983 (N_7983,N_1433,N_5958);
or U7984 (N_7984,N_3474,N_3473);
or U7985 (N_7985,N_2402,N_4843);
or U7986 (N_7986,N_4952,N_6104);
xor U7987 (N_7987,N_4295,N_5027);
nor U7988 (N_7988,N_5270,N_1955);
and U7989 (N_7989,N_1871,N_3014);
and U7990 (N_7990,N_1414,N_3464);
and U7991 (N_7991,N_295,N_2021);
xor U7992 (N_7992,N_4114,N_6228);
xor U7993 (N_7993,N_2104,N_6001);
nand U7994 (N_7994,N_2351,N_711);
nor U7995 (N_7995,N_664,N_2330);
nor U7996 (N_7996,N_4304,N_3444);
xnor U7997 (N_7997,N_4501,N_90);
and U7998 (N_7998,N_4256,N_3914);
or U7999 (N_7999,N_4106,N_658);
xor U8000 (N_8000,N_1228,N_475);
or U8001 (N_8001,N_2355,N_2628);
and U8002 (N_8002,N_3027,N_725);
or U8003 (N_8003,N_3762,N_3071);
nor U8004 (N_8004,N_2380,N_1219);
nand U8005 (N_8005,N_3233,N_1522);
nand U8006 (N_8006,N_3466,N_6041);
nor U8007 (N_8007,N_5800,N_6123);
or U8008 (N_8008,N_1499,N_775);
nand U8009 (N_8009,N_2761,N_4782);
nand U8010 (N_8010,N_4675,N_5223);
and U8011 (N_8011,N_5670,N_5744);
xnor U8012 (N_8012,N_4137,N_115);
or U8013 (N_8013,N_3261,N_1363);
nor U8014 (N_8014,N_3465,N_2252);
nor U8015 (N_8015,N_3461,N_5740);
nand U8016 (N_8016,N_1963,N_2637);
nand U8017 (N_8017,N_127,N_931);
nand U8018 (N_8018,N_2044,N_263);
and U8019 (N_8019,N_5403,N_6137);
nand U8020 (N_8020,N_284,N_1543);
nand U8021 (N_8021,N_3019,N_5134);
or U8022 (N_8022,N_3722,N_6241);
or U8023 (N_8023,N_1801,N_5820);
and U8024 (N_8024,N_3623,N_4550);
and U8025 (N_8025,N_2957,N_2042);
and U8026 (N_8026,N_5031,N_1578);
nor U8027 (N_8027,N_4102,N_5497);
nor U8028 (N_8028,N_4398,N_783);
and U8029 (N_8029,N_1597,N_1529);
nor U8030 (N_8030,N_4569,N_2140);
or U8031 (N_8031,N_2934,N_2174);
or U8032 (N_8032,N_1526,N_5306);
nand U8033 (N_8033,N_4211,N_398);
and U8034 (N_8034,N_3400,N_4356);
nor U8035 (N_8035,N_5788,N_1308);
nor U8036 (N_8036,N_4867,N_4467);
xor U8037 (N_8037,N_1644,N_2692);
nor U8038 (N_8038,N_3382,N_543);
xnor U8039 (N_8039,N_513,N_2907);
nand U8040 (N_8040,N_925,N_250);
nor U8041 (N_8041,N_4802,N_1575);
nor U8042 (N_8042,N_4429,N_1245);
nand U8043 (N_8043,N_3060,N_3651);
or U8044 (N_8044,N_898,N_2962);
nor U8045 (N_8045,N_1305,N_5588);
and U8046 (N_8046,N_2202,N_993);
or U8047 (N_8047,N_1070,N_3123);
or U8048 (N_8048,N_5154,N_2268);
xnor U8049 (N_8049,N_2504,N_2671);
and U8050 (N_8050,N_6175,N_1153);
or U8051 (N_8051,N_3579,N_5375);
nor U8052 (N_8052,N_5823,N_4351);
and U8053 (N_8053,N_5651,N_1004);
nor U8054 (N_8054,N_4212,N_1080);
xnor U8055 (N_8055,N_5098,N_1592);
nand U8056 (N_8056,N_5524,N_5096);
nand U8057 (N_8057,N_1663,N_1693);
or U8058 (N_8058,N_5224,N_2123);
or U8059 (N_8059,N_1730,N_4631);
nor U8060 (N_8060,N_1835,N_75);
and U8061 (N_8061,N_1925,N_3753);
nand U8062 (N_8062,N_1233,N_1813);
xor U8063 (N_8063,N_3663,N_5660);
nand U8064 (N_8064,N_5779,N_2593);
nand U8065 (N_8065,N_390,N_3102);
and U8066 (N_8066,N_1041,N_518);
or U8067 (N_8067,N_5824,N_5922);
nand U8068 (N_8068,N_2981,N_2852);
xnor U8069 (N_8069,N_1195,N_1484);
nor U8070 (N_8070,N_6037,N_6047);
nor U8071 (N_8071,N_4442,N_376);
or U8072 (N_8072,N_5100,N_1979);
nor U8073 (N_8073,N_2040,N_3015);
xor U8074 (N_8074,N_4667,N_2416);
nor U8075 (N_8075,N_1167,N_4055);
nand U8076 (N_8076,N_1464,N_2573);
and U8077 (N_8077,N_2000,N_4706);
or U8078 (N_8078,N_5147,N_3625);
nor U8079 (N_8079,N_2009,N_5374);
nand U8080 (N_8080,N_2283,N_6021);
nand U8081 (N_8081,N_2942,N_2954);
and U8082 (N_8082,N_5039,N_1948);
nand U8083 (N_8083,N_2640,N_4705);
nor U8084 (N_8084,N_229,N_4134);
nand U8085 (N_8085,N_3758,N_2218);
and U8086 (N_8086,N_4164,N_3142);
nor U8087 (N_8087,N_968,N_1792);
nor U8088 (N_8088,N_3028,N_73);
nand U8089 (N_8089,N_2381,N_2769);
and U8090 (N_8090,N_5835,N_218);
nor U8091 (N_8091,N_4861,N_3177);
and U8092 (N_8092,N_5725,N_4167);
or U8093 (N_8093,N_3736,N_1890);
nor U8094 (N_8094,N_441,N_5252);
nand U8095 (N_8095,N_3608,N_5328);
or U8096 (N_8096,N_2501,N_2081);
xor U8097 (N_8097,N_433,N_2651);
nor U8098 (N_8098,N_3575,N_2513);
or U8099 (N_8099,N_2491,N_302);
or U8100 (N_8100,N_5124,N_5261);
nor U8101 (N_8101,N_1716,N_6110);
nand U8102 (N_8102,N_3590,N_474);
or U8103 (N_8103,N_192,N_3732);
nor U8104 (N_8104,N_1087,N_3945);
nor U8105 (N_8105,N_413,N_4693);
and U8106 (N_8106,N_4992,N_5768);
nand U8107 (N_8107,N_1799,N_744);
and U8108 (N_8108,N_2982,N_5491);
nor U8109 (N_8109,N_1884,N_1712);
nor U8110 (N_8110,N_1282,N_809);
or U8111 (N_8111,N_3117,N_2146);
nand U8112 (N_8112,N_1396,N_3496);
and U8113 (N_8113,N_4058,N_3748);
nor U8114 (N_8114,N_2247,N_689);
xnor U8115 (N_8115,N_5857,N_454);
or U8116 (N_8116,N_4933,N_5349);
nand U8117 (N_8117,N_816,N_6014);
nand U8118 (N_8118,N_651,N_4642);
nor U8119 (N_8119,N_740,N_2157);
xnor U8120 (N_8120,N_2149,N_3819);
nand U8121 (N_8121,N_3952,N_607);
or U8122 (N_8122,N_5522,N_2596);
and U8123 (N_8123,N_4150,N_1423);
or U8124 (N_8124,N_4720,N_5696);
or U8125 (N_8125,N_67,N_2335);
or U8126 (N_8126,N_5060,N_107);
nor U8127 (N_8127,N_3384,N_5707);
nand U8128 (N_8128,N_3867,N_1780);
nor U8129 (N_8129,N_3399,N_2027);
and U8130 (N_8130,N_4278,N_6052);
or U8131 (N_8131,N_2788,N_1960);
and U8132 (N_8132,N_3368,N_5260);
or U8133 (N_8133,N_1136,N_5727);
nand U8134 (N_8134,N_3005,N_5298);
or U8135 (N_8135,N_2256,N_264);
xor U8136 (N_8136,N_169,N_3304);
nand U8137 (N_8137,N_500,N_3347);
or U8138 (N_8138,N_4204,N_780);
or U8139 (N_8139,N_4153,N_2277);
nand U8140 (N_8140,N_2831,N_2453);
nor U8141 (N_8141,N_672,N_3580);
nor U8142 (N_8142,N_3629,N_3491);
or U8143 (N_8143,N_4144,N_5126);
nand U8144 (N_8144,N_3600,N_5239);
nand U8145 (N_8145,N_149,N_1614);
nor U8146 (N_8146,N_3002,N_4897);
nor U8147 (N_8147,N_5179,N_5508);
or U8148 (N_8148,N_5333,N_2298);
or U8149 (N_8149,N_4577,N_1535);
xor U8150 (N_8150,N_5038,N_1546);
xnor U8151 (N_8151,N_1485,N_1900);
nor U8152 (N_8152,N_3419,N_2362);
and U8153 (N_8153,N_2433,N_1465);
or U8154 (N_8154,N_2349,N_113);
nor U8155 (N_8155,N_6043,N_3911);
nand U8156 (N_8156,N_5527,N_1186);
nand U8157 (N_8157,N_4865,N_896);
or U8158 (N_8158,N_357,N_6065);
nor U8159 (N_8159,N_5155,N_4019);
or U8160 (N_8160,N_4491,N_2778);
nand U8161 (N_8161,N_571,N_4841);
or U8162 (N_8162,N_1306,N_2785);
nor U8163 (N_8163,N_5069,N_2412);
and U8164 (N_8164,N_694,N_2100);
nand U8165 (N_8165,N_3798,N_3912);
and U8166 (N_8166,N_1973,N_1128);
nor U8167 (N_8167,N_3841,N_2588);
or U8168 (N_8168,N_3478,N_3689);
and U8169 (N_8169,N_1265,N_3245);
nand U8170 (N_8170,N_953,N_4714);
nand U8171 (N_8171,N_1098,N_1275);
nor U8172 (N_8172,N_2829,N_5459);
and U8173 (N_8173,N_5017,N_3079);
xor U8174 (N_8174,N_2293,N_1907);
nand U8175 (N_8175,N_4495,N_1242);
and U8176 (N_8176,N_6202,N_5700);
and U8177 (N_8177,N_1408,N_4603);
or U8178 (N_8178,N_5334,N_3760);
or U8179 (N_8179,N_4251,N_4658);
nor U8180 (N_8180,N_1106,N_3987);
or U8181 (N_8181,N_2797,N_175);
xor U8182 (N_8182,N_344,N_1551);
nor U8183 (N_8183,N_5379,N_5711);
or U8184 (N_8184,N_3213,N_5064);
nand U8185 (N_8185,N_1017,N_4449);
xor U8186 (N_8186,N_6174,N_5339);
and U8187 (N_8187,N_5477,N_4159);
nand U8188 (N_8188,N_519,N_6057);
nor U8189 (N_8189,N_992,N_157);
nor U8190 (N_8190,N_5681,N_6195);
and U8191 (N_8191,N_3726,N_201);
nor U8192 (N_8192,N_1206,N_3098);
nor U8193 (N_8193,N_5649,N_5632);
and U8194 (N_8194,N_4022,N_3200);
nand U8195 (N_8195,N_6004,N_4846);
and U8196 (N_8196,N_361,N_1361);
and U8197 (N_8197,N_4482,N_3589);
or U8198 (N_8198,N_2697,N_5132);
nand U8199 (N_8199,N_769,N_432);
xnor U8200 (N_8200,N_2558,N_5686);
or U8201 (N_8201,N_4331,N_2210);
nand U8202 (N_8202,N_2033,N_2932);
or U8203 (N_8203,N_668,N_5312);
nor U8204 (N_8204,N_4147,N_6003);
xnor U8205 (N_8205,N_2022,N_1122);
xnor U8206 (N_8206,N_970,N_4797);
and U8207 (N_8207,N_3196,N_5110);
and U8208 (N_8208,N_1197,N_3928);
or U8209 (N_8209,N_841,N_3070);
or U8210 (N_8210,N_275,N_2967);
or U8211 (N_8211,N_2575,N_3917);
nand U8212 (N_8212,N_657,N_767);
and U8213 (N_8213,N_4743,N_1616);
nand U8214 (N_8214,N_3374,N_5848);
and U8215 (N_8215,N_4352,N_4994);
or U8216 (N_8216,N_507,N_5078);
xnor U8217 (N_8217,N_2069,N_2930);
or U8218 (N_8218,N_5865,N_2586);
nand U8219 (N_8219,N_5095,N_2120);
and U8220 (N_8220,N_3591,N_4458);
nand U8221 (N_8221,N_5810,N_3483);
nand U8222 (N_8222,N_1109,N_736);
nor U8223 (N_8223,N_1395,N_627);
nor U8224 (N_8224,N_4434,N_5807);
nor U8225 (N_8225,N_5390,N_1428);
and U8226 (N_8226,N_3307,N_1127);
and U8227 (N_8227,N_1706,N_3479);
and U8228 (N_8228,N_5172,N_2479);
or U8229 (N_8229,N_1256,N_4363);
nand U8230 (N_8230,N_1683,N_679);
nor U8231 (N_8231,N_1261,N_448);
xor U8232 (N_8232,N_2191,N_3321);
or U8233 (N_8233,N_4035,N_5290);
or U8234 (N_8234,N_3578,N_4438);
nand U8235 (N_8235,N_3252,N_770);
nand U8236 (N_8236,N_1623,N_3999);
nor U8237 (N_8237,N_675,N_3545);
nor U8238 (N_8238,N_51,N_2455);
nor U8239 (N_8239,N_5092,N_1410);
and U8240 (N_8240,N_3507,N_4389);
and U8241 (N_8241,N_322,N_3951);
or U8242 (N_8242,N_553,N_5736);
nand U8243 (N_8243,N_3814,N_4685);
nand U8244 (N_8244,N_2271,N_1994);
or U8245 (N_8245,N_587,N_5140);
nor U8246 (N_8246,N_4758,N_1527);
xnor U8247 (N_8247,N_4591,N_5705);
or U8248 (N_8248,N_835,N_573);
nor U8249 (N_8249,N_4314,N_890);
nor U8250 (N_8250,N_3494,N_894);
nand U8251 (N_8251,N_5316,N_3652);
nor U8252 (N_8252,N_280,N_2510);
and U8253 (N_8253,N_1793,N_1579);
nand U8254 (N_8254,N_5322,N_5962);
or U8255 (N_8255,N_1346,N_424);
nor U8256 (N_8256,N_5949,N_784);
nor U8257 (N_8257,N_2611,N_112);
nand U8258 (N_8258,N_5443,N_395);
or U8259 (N_8259,N_881,N_241);
nor U8260 (N_8260,N_3825,N_6095);
nor U8261 (N_8261,N_2767,N_1949);
nor U8262 (N_8262,N_616,N_762);
and U8263 (N_8263,N_3223,N_1533);
and U8264 (N_8264,N_5114,N_2886);
nand U8265 (N_8265,N_2923,N_1988);
nand U8266 (N_8266,N_3156,N_2068);
nand U8267 (N_8267,N_2031,N_3537);
and U8268 (N_8268,N_3737,N_1116);
nand U8269 (N_8269,N_3794,N_119);
and U8270 (N_8270,N_5544,N_2737);
nor U8271 (N_8271,N_4849,N_5370);
nor U8272 (N_8272,N_2288,N_1131);
nor U8273 (N_8273,N_4034,N_5787);
nor U8274 (N_8274,N_1005,N_446);
and U8275 (N_8275,N_1402,N_2796);
nor U8276 (N_8276,N_2944,N_5546);
nand U8277 (N_8277,N_4245,N_6068);
nor U8278 (N_8278,N_3434,N_4513);
nor U8279 (N_8279,N_2799,N_2808);
nand U8280 (N_8280,N_6179,N_4075);
or U8281 (N_8281,N_2991,N_3086);
or U8282 (N_8282,N_6229,N_3808);
or U8283 (N_8283,N_87,N_2020);
and U8284 (N_8284,N_2294,N_2807);
or U8285 (N_8285,N_914,N_3414);
nor U8286 (N_8286,N_3837,N_5517);
nand U8287 (N_8287,N_1332,N_6165);
and U8288 (N_8288,N_812,N_3274);
and U8289 (N_8289,N_1773,N_1787);
and U8290 (N_8290,N_5466,N_6189);
nand U8291 (N_8291,N_3961,N_4383);
xor U8292 (N_8292,N_5505,N_4183);
nor U8293 (N_8293,N_4678,N_552);
nand U8294 (N_8294,N_2977,N_3924);
nand U8295 (N_8295,N_2667,N_5242);
nor U8296 (N_8296,N_5363,N_3498);
and U8297 (N_8297,N_2093,N_3548);
or U8298 (N_8298,N_1082,N_2622);
and U8299 (N_8299,N_4656,N_5845);
or U8300 (N_8300,N_2676,N_5049);
nand U8301 (N_8301,N_2456,N_3201);
nor U8302 (N_8302,N_3380,N_3926);
and U8303 (N_8303,N_3967,N_5861);
and U8304 (N_8304,N_6140,N_5214);
nor U8305 (N_8305,N_2424,N_583);
nand U8306 (N_8306,N_3470,N_2132);
xor U8307 (N_8307,N_2483,N_2066);
and U8308 (N_8308,N_4270,N_272);
and U8309 (N_8309,N_3696,N_2600);
and U8310 (N_8310,N_1284,N_2310);
nor U8311 (N_8311,N_3631,N_4068);
and U8312 (N_8312,N_1222,N_104);
nand U8313 (N_8313,N_3379,N_253);
nand U8314 (N_8314,N_1532,N_6062);
or U8315 (N_8315,N_1725,N_4319);
nor U8316 (N_8316,N_5020,N_3113);
nor U8317 (N_8317,N_3403,N_5392);
nor U8318 (N_8318,N_3605,N_6054);
nor U8319 (N_8319,N_1770,N_1901);
nand U8320 (N_8320,N_401,N_2372);
nand U8321 (N_8321,N_3661,N_3052);
nor U8322 (N_8322,N_1033,N_5311);
xnor U8323 (N_8323,N_1794,N_2435);
and U8324 (N_8324,N_2814,N_2101);
and U8325 (N_8325,N_2091,N_106);
and U8326 (N_8326,N_4081,N_4864);
nand U8327 (N_8327,N_3062,N_4254);
and U8328 (N_8328,N_3889,N_5683);
and U8329 (N_8329,N_721,N_5984);
nand U8330 (N_8330,N_5053,N_1358);
and U8331 (N_8331,N_2286,N_3985);
and U8332 (N_8332,N_3250,N_4082);
or U8333 (N_8333,N_50,N_4800);
or U8334 (N_8334,N_4666,N_5019);
and U8335 (N_8335,N_4380,N_1802);
nor U8336 (N_8336,N_1144,N_4757);
nand U8337 (N_8337,N_2306,N_4792);
and U8338 (N_8338,N_4302,N_2291);
nand U8339 (N_8339,N_731,N_1561);
nor U8340 (N_8340,N_2625,N_5535);
nand U8341 (N_8341,N_5057,N_1118);
or U8342 (N_8342,N_1865,N_4325);
and U8343 (N_8343,N_4226,N_3065);
and U8344 (N_8344,N_2774,N_79);
or U8345 (N_8345,N_5229,N_1855);
nand U8346 (N_8346,N_1292,N_3416);
and U8347 (N_8347,N_188,N_3822);
or U8348 (N_8348,N_3207,N_5042);
xnor U8349 (N_8349,N_1177,N_4576);
or U8350 (N_8350,N_4744,N_5033);
nor U8351 (N_8351,N_5977,N_2917);
nand U8352 (N_8352,N_5357,N_722);
nor U8353 (N_8353,N_4755,N_3159);
or U8354 (N_8354,N_2346,N_5361);
and U8355 (N_8355,N_3504,N_2648);
nand U8356 (N_8356,N_6249,N_2415);
or U8357 (N_8357,N_3786,N_392);
and U8358 (N_8358,N_46,N_80);
xor U8359 (N_8359,N_2963,N_6071);
or U8360 (N_8360,N_575,N_4298);
nor U8361 (N_8361,N_733,N_4627);
nor U8362 (N_8362,N_5536,N_3601);
nor U8363 (N_8363,N_5558,N_2144);
nor U8364 (N_8364,N_4240,N_4128);
nor U8365 (N_8365,N_772,N_2919);
xnor U8366 (N_8366,N_1311,N_2111);
nor U8367 (N_8367,N_4878,N_3620);
or U8368 (N_8368,N_96,N_2109);
nor U8369 (N_8369,N_1151,N_3894);
nand U8370 (N_8370,N_1335,N_4905);
or U8371 (N_8371,N_1821,N_3622);
and U8372 (N_8372,N_1020,N_259);
and U8373 (N_8373,N_217,N_4318);
or U8374 (N_8374,N_2511,N_5044);
nand U8375 (N_8375,N_4411,N_2437);
and U8376 (N_8376,N_2014,N_1336);
nand U8377 (N_8377,N_5733,N_5526);
and U8378 (N_8378,N_604,N_4214);
nand U8379 (N_8379,N_4551,N_6096);
or U8380 (N_8380,N_1898,N_2987);
nand U8381 (N_8381,N_1270,N_634);
nor U8382 (N_8382,N_6070,N_4329);
and U8383 (N_8383,N_3887,N_2281);
xor U8384 (N_8384,N_5495,N_5514);
or U8385 (N_8385,N_196,N_5440);
nand U8386 (N_8386,N_6061,N_12);
or U8387 (N_8387,N_5616,N_537);
nor U8388 (N_8388,N_4634,N_2287);
or U8389 (N_8389,N_414,N_4453);
or U8390 (N_8390,N_3299,N_2186);
or U8391 (N_8391,N_4928,N_3438);
and U8392 (N_8392,N_4698,N_6206);
or U8393 (N_8393,N_1729,N_4088);
or U8394 (N_8394,N_2878,N_3902);
and U8395 (N_8395,N_5957,N_4026);
and U8396 (N_8396,N_3120,N_2211);
or U8397 (N_8397,N_6039,N_48);
xnor U8398 (N_8398,N_2475,N_6161);
or U8399 (N_8399,N_6063,N_1715);
and U8400 (N_8400,N_6223,N_4367);
or U8401 (N_8401,N_2669,N_2720);
or U8402 (N_8402,N_1339,N_1184);
nand U8403 (N_8403,N_880,N_402);
xor U8404 (N_8404,N_4439,N_2951);
nand U8405 (N_8405,N_1010,N_5898);
xnor U8406 (N_8406,N_3831,N_3771);
nor U8407 (N_8407,N_2924,N_5891);
nor U8408 (N_8408,N_4405,N_1877);
or U8409 (N_8409,N_2542,N_5826);
or U8410 (N_8410,N_1738,N_5966);
or U8411 (N_8411,N_1221,N_1541);
nand U8412 (N_8412,N_5352,N_4951);
nand U8413 (N_8413,N_2085,N_1386);
and U8414 (N_8414,N_705,N_417);
nand U8415 (N_8415,N_142,N_4232);
nand U8416 (N_8416,N_3890,N_935);
or U8417 (N_8417,N_5351,N_4687);
xnor U8418 (N_8418,N_2579,N_3699);
or U8419 (N_8419,N_4542,N_2540);
xnor U8420 (N_8420,N_2979,N_3922);
and U8421 (N_8421,N_5515,N_372);
nand U8422 (N_8422,N_6029,N_5640);
and U8423 (N_8423,N_2263,N_4424);
or U8424 (N_8424,N_656,N_4842);
nand U8425 (N_8425,N_3008,N_216);
nor U8426 (N_8426,N_1422,N_1632);
or U8427 (N_8427,N_1347,N_83);
nand U8428 (N_8428,N_3816,N_5548);
nand U8429 (N_8429,N_5970,N_1713);
or U8430 (N_8430,N_3331,N_388);
nor U8431 (N_8431,N_6042,N_2848);
and U8432 (N_8432,N_739,N_5685);
nand U8433 (N_8433,N_2030,N_3852);
nor U8434 (N_8434,N_2528,N_1382);
or U8435 (N_8435,N_2233,N_3269);
or U8436 (N_8436,N_5579,N_2476);
nand U8437 (N_8437,N_3421,N_4855);
nand U8438 (N_8438,N_3144,N_4677);
nor U8439 (N_8439,N_5346,N_2722);
or U8440 (N_8440,N_1662,N_4837);
nor U8441 (N_8441,N_649,N_4464);
nand U8442 (N_8442,N_2595,N_2054);
and U8443 (N_8443,N_1633,N_4866);
nand U8444 (N_8444,N_2464,N_4169);
nand U8445 (N_8445,N_3131,N_1570);
nor U8446 (N_8446,N_2189,N_2680);
nor U8447 (N_8447,N_5765,N_37);
or U8448 (N_8448,N_2896,N_2480);
and U8449 (N_8449,N_1143,N_2914);
and U8450 (N_8450,N_5432,N_4030);
nand U8451 (N_8451,N_1580,N_5445);
or U8452 (N_8452,N_2709,N_2702);
nand U8453 (N_8453,N_4927,N_4218);
nand U8454 (N_8454,N_3175,N_1894);
nand U8455 (N_8455,N_1931,N_2731);
or U8456 (N_8456,N_5469,N_5262);
nor U8457 (N_8457,N_3112,N_5904);
nand U8458 (N_8458,N_1009,N_139);
nand U8459 (N_8459,N_5513,N_1269);
nor U8460 (N_8460,N_271,N_6219);
nand U8461 (N_8461,N_5326,N_1390);
or U8462 (N_8462,N_5156,N_2399);
and U8463 (N_8463,N_1026,N_1302);
nand U8464 (N_8464,N_5231,N_1048);
xnor U8465 (N_8465,N_3683,N_467);
xnor U8466 (N_8466,N_4957,N_4357);
or U8467 (N_8467,N_1504,N_3723);
nor U8468 (N_8468,N_161,N_5437);
or U8469 (N_8469,N_2779,N_3865);
and U8470 (N_8470,N_1891,N_2762);
nand U8471 (N_8471,N_4062,N_4756);
nor U8472 (N_8472,N_4186,N_2551);
nand U8473 (N_8473,N_803,N_293);
and U8474 (N_8474,N_3048,N_2503);
and U8475 (N_8475,N_6016,N_5571);
and U8476 (N_8476,N_1809,N_6121);
nand U8477 (N_8477,N_52,N_3328);
nand U8478 (N_8478,N_3183,N_3055);
or U8479 (N_8479,N_4844,N_2578);
or U8480 (N_8480,N_3909,N_1142);
xor U8481 (N_8481,N_1516,N_2790);
or U8482 (N_8482,N_6085,N_2736);
nand U8483 (N_8483,N_1119,N_2632);
nor U8484 (N_8484,N_1602,N_2162);
xnor U8485 (N_8485,N_620,N_4397);
xnor U8486 (N_8486,N_3334,N_4862);
and U8487 (N_8487,N_4179,N_2678);
and U8488 (N_8488,N_994,N_317);
nand U8489 (N_8489,N_982,N_6046);
nor U8490 (N_8490,N_2129,N_846);
xnor U8491 (N_8491,N_3294,N_63);
nor U8492 (N_8492,N_1097,N_5199);
or U8493 (N_8493,N_4468,N_3063);
xnor U8494 (N_8494,N_5238,N_2342);
or U8495 (N_8495,N_1520,N_1863);
nor U8496 (N_8496,N_3244,N_4161);
nand U8497 (N_8497,N_4,N_1617);
or U8498 (N_8498,N_6128,N_2705);
or U8499 (N_8499,N_4500,N_5149);
nor U8500 (N_8500,N_2543,N_1598);
nand U8501 (N_8501,N_1090,N_4701);
xnor U8502 (N_8502,N_4074,N_1968);
nor U8503 (N_8503,N_1981,N_3962);
nand U8504 (N_8504,N_5451,N_3021);
and U8505 (N_8505,N_4463,N_6067);
xnor U8506 (N_8506,N_4798,N_907);
nor U8507 (N_8507,N_2477,N_3448);
nor U8508 (N_8508,N_1796,N_1399);
or U8509 (N_8509,N_4190,N_3253);
nor U8510 (N_8510,N_5674,N_3558);
xor U8511 (N_8511,N_4443,N_3997);
nand U8512 (N_8512,N_2541,N_1023);
nand U8513 (N_8513,N_4192,N_1685);
or U8514 (N_8514,N_3340,N_1392);
xor U8515 (N_8515,N_3467,N_5160);
and U8516 (N_8516,N_4142,N_5714);
xor U8517 (N_8517,N_3847,N_1085);
xor U8518 (N_8518,N_3081,N_4315);
nor U8519 (N_8519,N_2612,N_4104);
and U8520 (N_8520,N_5188,N_1051);
nand U8521 (N_8521,N_4664,N_4350);
and U8522 (N_8522,N_3567,N_5067);
or U8523 (N_8523,N_4637,N_5427);
or U8524 (N_8524,N_2912,N_5530);
nand U8525 (N_8525,N_1329,N_5107);
and U8526 (N_8526,N_2087,N_3774);
nand U8527 (N_8527,N_4565,N_2529);
nor U8528 (N_8528,N_3801,N_2913);
nor U8529 (N_8529,N_538,N_3662);
xor U8530 (N_8530,N_442,N_1816);
nand U8531 (N_8531,N_4826,N_5902);
or U8532 (N_8532,N_5286,N_3908);
nor U8533 (N_8533,N_477,N_5699);
xnor U8534 (N_8534,N_1038,N_5533);
and U8535 (N_8535,N_1689,N_633);
nor U8536 (N_8536,N_4145,N_5575);
nand U8537 (N_8537,N_3205,N_2723);
nor U8538 (N_8538,N_3110,N_2995);
nand U8539 (N_8539,N_5592,N_2289);
nand U8540 (N_8540,N_2006,N_460);
and U8541 (N_8541,N_4857,N_1159);
nand U8542 (N_8542,N_5271,N_4733);
and U8543 (N_8543,N_3423,N_686);
or U8544 (N_8544,N_4202,N_2243);
or U8545 (N_8545,N_714,N_1126);
nand U8546 (N_8546,N_799,N_1947);
and U8547 (N_8547,N_3293,N_4728);
xnor U8548 (N_8548,N_6074,N_661);
xor U8549 (N_8549,N_1519,N_4840);
or U8550 (N_8550,N_2645,N_2838);
or U8551 (N_8551,N_4771,N_1341);
nand U8552 (N_8552,N_1777,N_3064);
or U8553 (N_8553,N_3915,N_3844);
or U8554 (N_8554,N_4493,N_4175);
or U8555 (N_8555,N_1707,N_670);
or U8556 (N_8556,N_570,N_5710);
nand U8557 (N_8557,N_3411,N_1784);
nand U8558 (N_8558,N_5294,N_5012);
nand U8559 (N_8559,N_5348,N_4626);
or U8560 (N_8560,N_3529,N_1839);
xnor U8561 (N_8561,N_3747,N_6160);
xnor U8562 (N_8562,N_5073,N_719);
nor U8563 (N_8563,N_1596,N_2105);
nand U8564 (N_8564,N_3115,N_5423);
xnor U8565 (N_8565,N_27,N_4097);
nand U8566 (N_8566,N_4737,N_3315);
or U8567 (N_8567,N_307,N_3137);
xnor U8568 (N_8568,N_5584,N_4790);
and U8569 (N_8569,N_5618,N_872);
and U8570 (N_8570,N_3029,N_3042);
nand U8571 (N_8571,N_6244,N_1640);
and U8572 (N_8572,N_825,N_1594);
nor U8573 (N_8573,N_103,N_1739);
nand U8574 (N_8574,N_5996,N_2682);
and U8575 (N_8575,N_5828,N_4718);
and U8576 (N_8576,N_586,N_2592);
xor U8577 (N_8577,N_2783,N_3125);
or U8578 (N_8578,N_663,N_6005);
nor U8579 (N_8579,N_4762,N_4649);
xnor U8580 (N_8580,N_4355,N_3305);
nand U8581 (N_8581,N_32,N_4559);
and U8582 (N_8582,N_3417,N_3189);
nand U8583 (N_8583,N_1860,N_4948);
nand U8584 (N_8584,N_2471,N_1637);
nand U8585 (N_8585,N_3383,N_5769);
and U8586 (N_8586,N_5492,N_6221);
or U8587 (N_8587,N_1251,N_4107);
nand U8588 (N_8588,N_1397,N_5230);
and U8589 (N_8589,N_3227,N_369);
and U8590 (N_8590,N_3766,N_3472);
nand U8591 (N_8591,N_3254,N_2631);
and U8592 (N_8592,N_3701,N_3458);
and U8593 (N_8593,N_3839,N_1549);
nand U8594 (N_8594,N_5981,N_732);
xor U8595 (N_8595,N_4809,N_5691);
nand U8596 (N_8596,N_1922,N_5960);
nand U8597 (N_8597,N_5974,N_5927);
and U8598 (N_8598,N_979,N_3654);
nand U8599 (N_8599,N_114,N_4366);
or U8600 (N_8600,N_3619,N_4066);
nor U8601 (N_8601,N_3093,N_1158);
or U8602 (N_8602,N_212,N_3300);
or U8603 (N_8603,N_4253,N_2583);
nor U8604 (N_8604,N_5414,N_826);
and U8605 (N_8605,N_2875,N_4393);
and U8606 (N_8606,N_1844,N_4735);
nor U8607 (N_8607,N_1489,N_5995);
nand U8608 (N_8608,N_1700,N_391);
xnor U8609 (N_8609,N_1281,N_2036);
nand U8610 (N_8610,N_3551,N_6162);
nand U8611 (N_8611,N_1078,N_1060);
nor U8612 (N_8612,N_4344,N_429);
nand U8613 (N_8613,N_326,N_5757);
xnor U8614 (N_8614,N_1550,N_5750);
nand U8615 (N_8615,N_2094,N_2664);
and U8616 (N_8616,N_5103,N_3195);
nand U8617 (N_8617,N_763,N_5600);
nor U8618 (N_8618,N_5244,N_2413);
and U8619 (N_8619,N_5550,N_4230);
and U8620 (N_8620,N_2745,N_4847);
and U8621 (N_8621,N_4028,N_3163);
nand U8622 (N_8622,N_255,N_3983);
or U8623 (N_8623,N_5236,N_485);
and U8624 (N_8624,N_4524,N_3546);
nand U8625 (N_8625,N_5724,N_4925);
or U8626 (N_8626,N_1827,N_5797);
and U8627 (N_8627,N_2819,N_2879);
or U8628 (N_8628,N_3135,N_5567);
or U8629 (N_8629,N_1711,N_6036);
or U8630 (N_8630,N_2425,N_585);
xor U8631 (N_8631,N_1705,N_4953);
or U8632 (N_8632,N_1101,N_154);
or U8633 (N_8633,N_278,N_2563);
nand U8634 (N_8634,N_3921,N_3381);
nand U8635 (N_8635,N_5169,N_6122);
nor U8636 (N_8636,N_3793,N_4390);
nor U8637 (N_8637,N_4423,N_131);
nor U8638 (N_8638,N_2817,N_3332);
nand U8639 (N_8639,N_2755,N_5102);
nor U8640 (N_8640,N_1229,N_2303);
and U8641 (N_8641,N_3613,N_1057);
or U8642 (N_8642,N_2056,N_2296);
or U8643 (N_8643,N_1902,N_1139);
nor U8644 (N_8644,N_3779,N_5808);
and U8645 (N_8645,N_2201,N_3455);
nor U8646 (N_8646,N_2484,N_5540);
or U8647 (N_8647,N_1404,N_4016);
or U8648 (N_8648,N_4001,N_789);
nor U8649 (N_8649,N_5909,N_3050);
nand U8650 (N_8650,N_4372,N_3767);
nor U8651 (N_8651,N_1976,N_3122);
or U8652 (N_8652,N_3310,N_5773);
xnor U8653 (N_8653,N_4219,N_6019);
nor U8654 (N_8654,N_397,N_4883);
and U8655 (N_8655,N_4781,N_3398);
or U8656 (N_8656,N_2442,N_1309);
and U8657 (N_8657,N_5022,N_5032);
and U8658 (N_8658,N_523,N_4684);
xnor U8659 (N_8659,N_4651,N_3756);
and U8660 (N_8660,N_5066,N_535);
and U8661 (N_8661,N_4795,N_2569);
or U8662 (N_8662,N_1972,N_2046);
xnor U8663 (N_8663,N_209,N_44);
and U8664 (N_8664,N_5619,N_5917);
nor U8665 (N_8665,N_1962,N_2655);
xor U8666 (N_8666,N_3053,N_2097);
xnor U8667 (N_8667,N_3795,N_3925);
xor U8668 (N_8668,N_252,N_1367);
nand U8669 (N_8669,N_567,N_4121);
or U8670 (N_8670,N_2345,N_2304);
nand U8671 (N_8671,N_3764,N_2888);
nor U8672 (N_8672,N_2171,N_5948);
or U8673 (N_8673,N_4894,N_1161);
nand U8674 (N_8674,N_716,N_3459);
nor U8675 (N_8675,N_3989,N_1372);
nand U8676 (N_8676,N_5543,N_1431);
or U8677 (N_8677,N_1838,N_4976);
nand U8678 (N_8678,N_870,N_4341);
nor U8679 (N_8679,N_5877,N_1356);
nand U8680 (N_8680,N_4244,N_5869);
nor U8681 (N_8681,N_4049,N_4029);
nor U8682 (N_8682,N_708,N_2107);
or U8683 (N_8683,N_425,N_4051);
or U8684 (N_8684,N_416,N_4815);
nand U8685 (N_8685,N_3462,N_718);
nor U8686 (N_8686,N_5283,N_1812);
nand U8687 (N_8687,N_4578,N_2418);
nand U8688 (N_8688,N_1380,N_2265);
or U8689 (N_8689,N_126,N_5856);
nand U8690 (N_8690,N_646,N_1944);
nand U8691 (N_8691,N_121,N_4194);
nand U8692 (N_8692,N_5630,N_1510);
and U8693 (N_8693,N_3860,N_5557);
or U8694 (N_8694,N_3673,N_3929);
nand U8695 (N_8695,N_5802,N_2876);
nand U8696 (N_8696,N_3540,N_1209);
nand U8697 (N_8697,N_3960,N_4584);
nor U8698 (N_8698,N_2241,N_947);
or U8699 (N_8699,N_666,N_6180);
and U8700 (N_8700,N_3901,N_1218);
xor U8701 (N_8701,N_4903,N_3727);
nand U8702 (N_8702,N_5358,N_499);
or U8703 (N_8703,N_3615,N_4604);
nor U8704 (N_8704,N_997,N_6088);
and U8705 (N_8705,N_5655,N_4640);
and U8706 (N_8706,N_660,N_1062);
and U8707 (N_8707,N_2765,N_4593);
and U8708 (N_8708,N_2227,N_1698);
nand U8709 (N_8709,N_3314,N_5872);
nand U8710 (N_8710,N_6196,N_760);
and U8711 (N_8711,N_2937,N_3069);
or U8712 (N_8712,N_4599,N_2401);
and U8713 (N_8713,N_3904,N_5863);
xor U8714 (N_8714,N_3643,N_4015);
nor U8715 (N_8715,N_5089,N_5762);
or U8716 (N_8716,N_2883,N_873);
nand U8717 (N_8717,N_4506,N_2445);
nand U8718 (N_8718,N_3306,N_1333);
and U8719 (N_8719,N_5582,N_4290);
nor U8720 (N_8720,N_5356,N_3616);
and U8721 (N_8721,N_2764,N_5831);
or U8722 (N_8722,N_2231,N_2319);
and U8723 (N_8723,N_3094,N_1011);
nand U8724 (N_8724,N_412,N_1359);
or U8725 (N_8725,N_1819,N_3211);
nand U8726 (N_8726,N_887,N_4531);
xor U8727 (N_8727,N_116,N_3878);
or U8728 (N_8728,N_178,N_2341);
nor U8729 (N_8729,N_5749,N_2459);
and U8730 (N_8730,N_5203,N_673);
and U8731 (N_8731,N_5021,N_4301);
or U8732 (N_8732,N_2546,N_884);
or U8733 (N_8733,N_1247,N_2580);
nand U8734 (N_8734,N_6159,N_5512);
nand U8735 (N_8735,N_4414,N_1983);
nor U8736 (N_8736,N_1204,N_5914);
nor U8737 (N_8737,N_4334,N_6173);
and U8738 (N_8738,N_1100,N_387);
or U8739 (N_8739,N_184,N_1572);
nand U8740 (N_8740,N_435,N_2023);
nand U8741 (N_8741,N_4480,N_5129);
nand U8742 (N_8742,N_340,N_2482);
and U8743 (N_8743,N_3907,N_1225);
and U8744 (N_8744,N_2685,N_2505);
and U8745 (N_8745,N_6101,N_5890);
or U8746 (N_8746,N_3133,N_89);
or U8747 (N_8747,N_3536,N_213);
xor U8748 (N_8748,N_81,N_4852);
nand U8749 (N_8749,N_1908,N_3515);
nor U8750 (N_8750,N_4643,N_2225);
nor U8751 (N_8751,N_6018,N_4924);
or U8752 (N_8752,N_4416,N_4259);
or U8753 (N_8753,N_3854,N_1045);
and U8754 (N_8754,N_3606,N_4608);
nand U8755 (N_8755,N_1374,N_6076);
and U8756 (N_8756,N_4031,N_3609);
nand U8757 (N_8757,N_1645,N_5015);
or U8758 (N_8758,N_335,N_906);
and U8759 (N_8759,N_3031,N_2235);
or U8760 (N_8760,N_3076,N_2594);
and U8761 (N_8761,N_4180,N_3435);
and U8762 (N_8762,N_555,N_1134);
nand U8763 (N_8763,N_5764,N_2423);
nand U8764 (N_8764,N_366,N_2842);
and U8765 (N_8765,N_69,N_1317);
nand U8766 (N_8766,N_2077,N_128);
and U8767 (N_8767,N_2928,N_2997);
nor U8768 (N_8768,N_4523,N_2339);
nand U8769 (N_8769,N_4811,N_3147);
or U8770 (N_8770,N_618,N_2138);
xor U8771 (N_8771,N_3665,N_1658);
nor U8772 (N_8772,N_5327,N_3222);
nor U8773 (N_8773,N_1704,N_3471);
nor U8774 (N_8774,N_5054,N_949);
or U8775 (N_8775,N_3596,N_120);
nor U8776 (N_8776,N_4541,N_4688);
or U8777 (N_8777,N_2946,N_3846);
nand U8778 (N_8778,N_5109,N_1224);
or U8779 (N_8779,N_489,N_5709);
or U8780 (N_8780,N_677,N_1708);
and U8781 (N_8781,N_1893,N_4471);
and U8782 (N_8782,N_5161,N_4225);
xor U8783 (N_8783,N_1291,N_1425);
xnor U8784 (N_8784,N_2389,N_2070);
nand U8785 (N_8785,N_2646,N_5372);
nor U8786 (N_8786,N_4645,N_2616);
nand U8787 (N_8787,N_205,N_2011);
nor U8788 (N_8788,N_5009,N_6045);
or U8789 (N_8789,N_5344,N_4201);
and U8790 (N_8790,N_1750,N_4761);
nand U8791 (N_8791,N_377,N_3039);
and U8792 (N_8792,N_2566,N_4901);
xnor U8793 (N_8793,N_4808,N_1215);
nand U8794 (N_8794,N_1846,N_2137);
xor U8795 (N_8795,N_2008,N_5938);
or U8796 (N_8796,N_4632,N_4697);
and U8797 (N_8797,N_827,N_3534);
nand U8798 (N_8798,N_3743,N_1002);
nand U8799 (N_8799,N_45,N_1515);
nor U8800 (N_8800,N_2512,N_525);
and U8801 (N_8801,N_3272,N_3751);
nor U8802 (N_8802,N_3607,N_1310);
or U8803 (N_8803,N_4529,N_5087);
or U8804 (N_8804,N_2943,N_4534);
nor U8805 (N_8805,N_2422,N_3856);
nor U8806 (N_8806,N_3745,N_1027);
nand U8807 (N_8807,N_5819,N_2718);
and U8808 (N_8808,N_4939,N_426);
or U8809 (N_8809,N_5603,N_1918);
nand U8810 (N_8810,N_1788,N_1173);
nor U8811 (N_8811,N_842,N_674);
nand U8812 (N_8812,N_236,N_863);
nor U8813 (N_8813,N_737,N_61);
and U8814 (N_8814,N_4221,N_186);
nand U8815 (N_8815,N_2507,N_5534);
and U8816 (N_8816,N_5404,N_4873);
nor U8817 (N_8817,N_2488,N_2658);
xnor U8818 (N_8818,N_4892,N_3895);
nand U8819 (N_8819,N_5897,N_1954);
nor U8820 (N_8820,N_2194,N_5599);
xnor U8821 (N_8821,N_5050,N_2134);
and U8822 (N_8822,N_2823,N_4238);
nand U8823 (N_8823,N_343,N_4080);
or U8824 (N_8824,N_2758,N_3781);
and U8825 (N_8825,N_1646,N_5438);
xnor U8826 (N_8826,N_321,N_4909);
and U8827 (N_8827,N_3883,N_6193);
or U8828 (N_8828,N_876,N_2880);
nand U8829 (N_8829,N_2712,N_5452);
and U8830 (N_8830,N_3172,N_2118);
or U8831 (N_8831,N_4618,N_4391);
and U8832 (N_8832,N_807,N_1674);
or U8833 (N_8833,N_3877,N_1573);
and U8834 (N_8834,N_5165,N_3203);
or U8835 (N_8835,N_2183,N_3162);
and U8836 (N_8836,N_2961,N_498);
xor U8837 (N_8837,N_2787,N_4131);
or U8838 (N_8838,N_3594,N_88);
or U8839 (N_8839,N_1851,N_5576);
xnor U8840 (N_8840,N_4138,N_1731);
nor U8841 (N_8841,N_1824,N_3187);
and U8842 (N_8842,N_6208,N_6099);
and U8843 (N_8843,N_4517,N_5812);
xor U8844 (N_8844,N_3681,N_3576);
nand U8845 (N_8845,N_3849,N_1387);
nand U8846 (N_8846,N_5659,N_759);
and U8847 (N_8847,N_1099,N_650);
nor U8848 (N_8848,N_1797,N_2854);
and U8849 (N_8849,N_3004,N_449);
nor U8850 (N_8850,N_3044,N_1042);
and U8851 (N_8851,N_3525,N_4877);
nand U8852 (N_8852,N_1766,N_5565);
nor U8853 (N_8853,N_5675,N_249);
xor U8854 (N_8854,N_3716,N_2028);
and U8855 (N_8855,N_5482,N_2447);
xor U8856 (N_8856,N_2515,N_4345);
nand U8857 (N_8857,N_1240,N_2994);
nand U8858 (N_8858,N_2024,N_1986);
or U8859 (N_8859,N_4968,N_5376);
and U8860 (N_8860,N_4820,N_1303);
or U8861 (N_8861,N_2927,N_282);
or U8862 (N_8862,N_239,N_3061);
xnor U8863 (N_8863,N_140,N_2124);
and U8864 (N_8864,N_584,N_5263);
or U8865 (N_8865,N_5556,N_3543);
and U8866 (N_8866,N_3688,N_2841);
xor U8867 (N_8867,N_3208,N_4041);
xnor U8868 (N_8868,N_777,N_2743);
nand U8869 (N_8869,N_5061,N_5218);
xnor U8870 (N_8870,N_3818,N_208);
or U8871 (N_8871,N_4089,N_1808);
xor U8872 (N_8872,N_839,N_1198);
and U8873 (N_8873,N_3547,N_4652);
nor U8874 (N_8874,N_755,N_3994);
nand U8875 (N_8875,N_5781,N_4518);
or U8876 (N_8876,N_3668,N_2554);
nand U8877 (N_8877,N_5175,N_5643);
or U8878 (N_8878,N_5587,N_5847);
and U8879 (N_8879,N_3428,N_26);
and U8880 (N_8880,N_5090,N_3243);
and U8881 (N_8881,N_4310,N_4987);
xnor U8882 (N_8882,N_1434,N_5034);
xor U8883 (N_8883,N_2133,N_4983);
or U8884 (N_8884,N_1449,N_4961);
and U8885 (N_8885,N_2639,N_2706);
nand U8886 (N_8886,N_2789,N_1344);
nand U8887 (N_8887,N_521,N_341);
and U8888 (N_8888,N_3100,N_3770);
or U8889 (N_8889,N_1437,N_4997);
and U8890 (N_8890,N_3555,N_168);
and U8891 (N_8891,N_362,N_680);
and U8892 (N_8892,N_3111,N_3378);
or U8893 (N_8893,N_5391,N_5399);
nor U8894 (N_8894,N_1370,N_1853);
and U8895 (N_8895,N_1660,N_1559);
or U8896 (N_8896,N_1958,N_4217);
nand U8897 (N_8897,N_3386,N_580);
nor U8898 (N_8898,N_2978,N_171);
xnor U8899 (N_8899,N_2606,N_1604);
and U8900 (N_8900,N_1194,N_4077);
nor U8901 (N_8901,N_1538,N_4312);
or U8902 (N_8902,N_5731,N_608);
nand U8903 (N_8903,N_4340,N_3450);
or U8904 (N_8904,N_1502,N_1833);
or U8905 (N_8905,N_3604,N_3869);
xor U8906 (N_8906,N_4791,N_3377);
or U8907 (N_8907,N_3224,N_5693);
nor U8908 (N_8908,N_3437,N_2469);
and U8909 (N_8909,N_1726,N_5827);
or U8910 (N_8910,N_2514,N_5745);
nor U8911 (N_8911,N_5915,N_294);
and U8912 (N_8912,N_1453,N_5397);
nand U8913 (N_8913,N_4234,N_5541);
xnor U8914 (N_8914,N_619,N_653);
nor U8915 (N_8915,N_2544,N_1007);
nand U8916 (N_8916,N_1278,N_2175);
xor U8917 (N_8917,N_4044,N_2792);
nand U8918 (N_8918,N_3164,N_1762);
nor U8919 (N_8919,N_2532,N_2248);
and U8920 (N_8920,N_954,N_915);
xnor U8921 (N_8921,N_407,N_6129);
nand U8922 (N_8922,N_2970,N_2379);
or U8923 (N_8923,N_929,N_4940);
nand U8924 (N_8924,N_4063,N_5825);
nand U8925 (N_8925,N_590,N_4803);
and U8926 (N_8926,N_3284,N_6227);
nand U8927 (N_8927,N_337,N_5989);
or U8928 (N_8928,N_4189,N_2710);
xor U8929 (N_8929,N_382,N_5635);
or U8930 (N_8930,N_2168,N_2481);
nand U8931 (N_8931,N_3886,N_4975);
or U8932 (N_8932,N_4083,N_2122);
and U8933 (N_8933,N_6185,N_3611);
or U8934 (N_8934,N_3588,N_706);
nand U8935 (N_8935,N_2161,N_1075);
nand U8936 (N_8936,N_2941,N_560);
and U8937 (N_8937,N_137,N_5313);
nand U8938 (N_8938,N_2487,N_1998);
nor U8939 (N_8939,N_3011,N_1832);
nand U8940 (N_8940,N_5876,N_399);
and U8941 (N_8941,N_2082,N_1837);
and U8942 (N_8942,N_5868,N_4747);
and U8943 (N_8943,N_883,N_1407);
and U8944 (N_8944,N_5366,N_5704);
nor U8945 (N_8945,N_1806,N_3804);
xnor U8946 (N_8946,N_3457,N_1223);
or U8947 (N_8947,N_1856,N_1508);
or U8948 (N_8948,N_1989,N_2988);
or U8949 (N_8949,N_1364,N_5969);
or U8950 (N_8950,N_802,N_5748);
nand U8951 (N_8951,N_2644,N_2827);
or U8952 (N_8952,N_5746,N_4660);
nor U8953 (N_8953,N_5472,N_5171);
nor U8954 (N_8954,N_480,N_4700);
or U8955 (N_8955,N_3687,N_3796);
and U8956 (N_8956,N_56,N_2894);
or U8957 (N_8957,N_3335,N_1401);
nor U8958 (N_8958,N_6120,N_2198);
xor U8959 (N_8959,N_3636,N_1452);
nand U8960 (N_8960,N_3322,N_4833);
nand U8961 (N_8961,N_1447,N_3644);
nand U8962 (N_8962,N_2079,N_5047);
and U8963 (N_8963,N_4891,N_6051);
nor U8964 (N_8964,N_4255,N_5689);
nor U8965 (N_8965,N_1150,N_4947);
and U8966 (N_8966,N_3484,N_2169);
nor U8967 (N_8967,N_2560,N_875);
nor U8968 (N_8968,N_6177,N_2443);
nor U8969 (N_8969,N_6166,N_5644);
nand U8970 (N_8970,N_4163,N_3150);
nand U8971 (N_8971,N_6023,N_4690);
or U8972 (N_8972,N_3212,N_5564);
and U8973 (N_8973,N_3285,N_3146);
nor U8974 (N_8974,N_5690,N_911);
nor U8975 (N_8975,N_3564,N_4904);
xor U8976 (N_8976,N_1710,N_5625);
nand U8977 (N_8977,N_4573,N_4011);
xnor U8978 (N_8978,N_24,N_709);
nor U8979 (N_8979,N_3326,N_3106);
nor U8980 (N_8980,N_5373,N_1686);
and U8981 (N_8981,N_3349,N_5968);
xnor U8982 (N_8982,N_2017,N_1601);
nand U8983 (N_8983,N_285,N_1895);
nor U8984 (N_8984,N_4006,N_470);
nand U8985 (N_8985,N_4547,N_1319);
and U8986 (N_8986,N_3409,N_4931);
xnor U8987 (N_8987,N_3275,N_3577);
xnor U8988 (N_8988,N_3906,N_5119);
nor U8989 (N_8989,N_2229,N_5139);
nor U8990 (N_8990,N_2500,N_328);
nor U8991 (N_8991,N_2307,N_3276);
or U8992 (N_8992,N_1753,N_4236);
xnor U8993 (N_8993,N_1977,N_1999);
or U8994 (N_8994,N_843,N_2083);
and U8995 (N_8995,N_3593,N_2576);
or U8996 (N_8996,N_2395,N_4422);
or U8997 (N_8997,N_4268,N_4944);
nor U8998 (N_8998,N_5481,N_5494);
and U8999 (N_8999,N_6126,N_2251);
nand U9000 (N_9000,N_221,N_1951);
or U9001 (N_9001,N_380,N_3528);
nand U9002 (N_9002,N_1858,N_2332);
and U9003 (N_9003,N_2209,N_2833);
or U9004 (N_9004,N_287,N_1353);
nor U9005 (N_9005,N_5715,N_3938);
or U9006 (N_9006,N_305,N_310);
or U9007 (N_9007,N_4025,N_628);
and U9008 (N_9008,N_4794,N_5734);
and U9009 (N_9009,N_1913,N_4956);
nor U9010 (N_9010,N_2155,N_3392);
nand U9011 (N_9011,N_3446,N_4377);
nand U9012 (N_9012,N_3641,N_3503);
or U9013 (N_9013,N_1411,N_4073);
xnor U9014 (N_9014,N_5117,N_4399);
or U9015 (N_9015,N_1001,N_5911);
nand U9016 (N_9016,N_3271,N_2537);
nand U9017 (N_9017,N_5447,N_4373);
nand U9018 (N_9018,N_551,N_752);
nand U9019 (N_9019,N_781,N_1677);
or U9020 (N_9020,N_2270,N_5597);
xor U9021 (N_9021,N_579,N_5656);
nor U9022 (N_9022,N_3171,N_4982);
and U9023 (N_9023,N_5002,N_76);
or U9024 (N_9024,N_2474,N_2429);
or U9025 (N_9025,N_3698,N_2278);
or U9026 (N_9026,N_4177,N_370);
or U9027 (N_9027,N_3080,N_5037);
nor U9028 (N_9028,N_1732,N_246);
and U9029 (N_9029,N_4610,N_3519);
nand U9030 (N_9030,N_297,N_6214);
nor U9031 (N_9031,N_1756,N_2793);
or U9032 (N_9032,N_1724,N_5676);
or U9033 (N_9033,N_865,N_3595);
or U9034 (N_9034,N_5628,N_5207);
and U9035 (N_9035,N_1869,N_4796);
and U9036 (N_9036,N_2366,N_2589);
or U9037 (N_9037,N_5232,N_3614);
or U9038 (N_9038,N_1435,N_1400);
nand U9039 (N_9039,N_2815,N_3375);
and U9040 (N_9040,N_4321,N_1154);
and U9041 (N_9041,N_5817,N_1175);
or U9042 (N_9042,N_3830,N_5225);
nor U9043 (N_9043,N_850,N_456);
nor U9044 (N_9044,N_1121,N_2936);
nor U9045 (N_9045,N_132,N_97);
or U9046 (N_9046,N_741,N_4496);
nand U9047 (N_9047,N_145,N_2744);
nor U9048 (N_9048,N_4401,N_1147);
xor U9049 (N_9049,N_5583,N_5259);
and U9050 (N_9050,N_3194,N_5849);
or U9051 (N_9051,N_2770,N_1120);
or U9052 (N_9052,N_5815,N_4824);
or U9053 (N_9053,N_4963,N_4419);
xnor U9054 (N_9054,N_2164,N_122);
xnor U9055 (N_9055,N_1659,N_5801);
xor U9056 (N_9056,N_3761,N_3612);
and U9057 (N_9057,N_1862,N_4478);
nand U9058 (N_9058,N_3572,N_2976);
and U9059 (N_9059,N_2925,N_4014);
nand U9060 (N_9060,N_4485,N_1071);
nor U9061 (N_9061,N_5772,N_5277);
or U9062 (N_9062,N_5284,N_4206);
nand U9063 (N_9063,N_3927,N_5993);
xnor U9064 (N_9064,N_2926,N_298);
nor U9065 (N_9065,N_2,N_5503);
and U9066 (N_9066,N_2361,N_6183);
nand U9067 (N_9067,N_66,N_2516);
or U9068 (N_9068,N_845,N_1786);
nor U9069 (N_9069,N_3959,N_2378);
nor U9070 (N_9070,N_235,N_17);
xnor U9071 (N_9071,N_4223,N_2245);
nor U9072 (N_9072,N_4335,N_2874);
or U9073 (N_9073,N_4010,N_536);
nor U9074 (N_9074,N_2766,N_3327);
or U9075 (N_9075,N_2811,N_5303);
and U9076 (N_9076,N_3936,N_2196);
nand U9077 (N_9077,N_2430,N_4387);
xor U9078 (N_9078,N_549,N_4923);
or U9079 (N_9079,N_3717,N_2478);
or U9080 (N_9080,N_3876,N_1460);
or U9081 (N_9081,N_2668,N_419);
or U9082 (N_9082,N_4817,N_4716);
or U9083 (N_9083,N_2846,N_5622);
and U9084 (N_9084,N_3571,N_43);
and U9085 (N_9085,N_1993,N_3942);
nand U9086 (N_9086,N_2253,N_4787);
xnor U9087 (N_9087,N_2862,N_4327);
nand U9088 (N_9088,N_5035,N_1881);
or U9089 (N_9089,N_3700,N_3370);
nor U9090 (N_9090,N_5732,N_18);
or U9091 (N_9091,N_4308,N_4935);
xnor U9092 (N_9092,N_3800,N_269);
or U9093 (N_9093,N_2561,N_3940);
nand U9094 (N_9094,N_4054,N_1416);
and U9095 (N_9095,N_2261,N_3191);
nand U9096 (N_9096,N_4119,N_5381);
xor U9097 (N_9097,N_941,N_2320);
and U9098 (N_9098,N_4184,N_1867);
nor U9099 (N_9099,N_4973,N_3087);
nor U9100 (N_9100,N_1412,N_5071);
or U9101 (N_9101,N_790,N_5594);
or U9102 (N_9102,N_1067,N_4483);
nor U9103 (N_9103,N_5726,N_5896);
xor U9104 (N_9104,N_2519,N_1563);
or U9105 (N_9105,N_2749,N_866);
or U9106 (N_9106,N_1590,N_928);
xnor U9107 (N_9107,N_85,N_531);
nor U9108 (N_9108,N_3971,N_4209);
nand U9109 (N_9109,N_1451,N_944);
nand U9110 (N_9110,N_1603,N_2908);
and U9111 (N_9111,N_4008,N_1682);
and U9112 (N_9112,N_415,N_3184);
xor U9113 (N_9113,N_2564,N_1664);
xnor U9114 (N_9114,N_801,N_4359);
and U9115 (N_9115,N_64,N_1162);
nand U9116 (N_9116,N_2200,N_520);
or U9117 (N_9117,N_3220,N_3838);
and U9118 (N_9118,N_4936,N_4568);
nand U9119 (N_9119,N_198,N_1896);
xor U9120 (N_9120,N_1512,N_1500);
and U9121 (N_9121,N_4516,N_4320);
nor U9122 (N_9122,N_3169,N_5296);
nor U9123 (N_9123,N_2901,N_2226);
nand U9124 (N_9124,N_6144,N_1426);
nand U9125 (N_9125,N_1757,N_1419);
nor U9126 (N_9126,N_5947,N_2969);
nand U9127 (N_9127,N_2327,N_2182);
nand U9128 (N_9128,N_5730,N_1260);
and U9129 (N_9129,N_4057,N_1250);
nor U9130 (N_9130,N_4641,N_4005);
and U9131 (N_9131,N_4395,N_1737);
and U9132 (N_9132,N_4908,N_1470);
xor U9133 (N_9133,N_2618,N_1389);
or U9134 (N_9134,N_659,N_1889);
nand U9135 (N_9135,N_857,N_6213);
nand U9136 (N_9136,N_6212,N_5112);
nor U9137 (N_9137,N_1409,N_5281);
nand U9138 (N_9138,N_6135,N_3352);
nor U9139 (N_9139,N_1675,N_5148);
or U9140 (N_9140,N_1765,N_2188);
nor U9141 (N_9141,N_1227,N_4945);
xnor U9142 (N_9142,N_3702,N_129);
xor U9143 (N_9143,N_5400,N_1035);
nor U9144 (N_9144,N_3868,N_4342);
nand U9145 (N_9145,N_4964,N_2562);
nand U9146 (N_9146,N_991,N_4469);
nor U9147 (N_9147,N_5384,N_5862);
nor U9148 (N_9148,N_6010,N_4481);
nand U9149 (N_9149,N_1338,N_5395);
nand U9150 (N_9150,N_1509,N_4149);
xnor U9151 (N_9151,N_4638,N_2931);
nand U9152 (N_9152,N_2699,N_1444);
nand U9153 (N_9153,N_637,N_5198);
nand U9154 (N_9154,N_778,N_5668);
nor U9155 (N_9155,N_4109,N_2130);
xnor U9156 (N_9156,N_3792,N_2865);
nand U9157 (N_9157,N_4198,N_4227);
nand U9158 (N_9158,N_3913,N_1496);
nand U9159 (N_9159,N_3797,N_6178);
nand U9160 (N_9160,N_3154,N_318);
nand U9161 (N_9161,N_4322,N_4966);
and U9162 (N_9162,N_515,N_5743);
and U9163 (N_9163,N_859,N_163);
nor U9164 (N_9164,N_4409,N_4564);
xor U9165 (N_9165,N_4479,N_5446);
nor U9166 (N_9166,N_4839,N_600);
and U9167 (N_9167,N_1970,N_6028);
and U9168 (N_9168,N_5282,N_1554);
and U9169 (N_9169,N_698,N_4174);
nor U9170 (N_9170,N_3084,N_3977);
and U9171 (N_9171,N_279,N_5121);
nand U9172 (N_9172,N_226,N_1357);
nor U9173 (N_9173,N_99,N_867);
nand U9174 (N_9174,N_5275,N_1879);
and U9175 (N_9175,N_5867,N_4165);
or U9176 (N_9176,N_5678,N_3302);
nor U9177 (N_9177,N_2820,N_2172);
and U9178 (N_9178,N_4086,N_165);
or U9179 (N_9179,N_3690,N_1268);
nand U9180 (N_9180,N_6072,N_4991);
nor U9181 (N_9181,N_3410,N_2732);
nor U9182 (N_9182,N_532,N_629);
or U9183 (N_9183,N_6091,N_3026);
and U9184 (N_9184,N_1699,N_4323);
nor U9185 (N_9185,N_3787,N_603);
or U9186 (N_9186,N_4136,N_3897);
or U9187 (N_9187,N_683,N_3780);
nand U9188 (N_9188,N_234,N_1086);
or U9189 (N_9189,N_974,N_4655);
nor U9190 (N_9190,N_5523,N_2861);
nor U9191 (N_9191,N_5910,N_5645);
nand U9192 (N_9192,N_4752,N_78);
nand U9193 (N_9193,N_792,N_3573);
xor U9194 (N_9194,N_5219,N_2026);
nor U9195 (N_9195,N_4732,N_5881);
nand U9196 (N_9196,N_2458,N_1274);
nor U9197 (N_9197,N_1238,N_1558);
and U9198 (N_9198,N_4768,N_440);
nand U9199 (N_9199,N_2584,N_986);
or U9200 (N_9200,N_4686,N_1458);
nand U9201 (N_9201,N_893,N_4999);
nand U9202 (N_9202,N_6207,N_6000);
nand U9203 (N_9203,N_1050,N_3813);
or U9204 (N_9204,N_3775,N_4763);
nor U9205 (N_9205,N_1582,N_5287);
xnor U9206 (N_9206,N_4622,N_3018);
and U9207 (N_9207,N_3848,N_5612);
nand U9208 (N_9208,N_4297,N_2909);
or U9209 (N_9209,N_5963,N_3116);
xor U9210 (N_9210,N_4751,N_270);
nand U9211 (N_9211,N_3861,N_6194);
nand U9212 (N_9212,N_4317,N_6230);
nor U9213 (N_9213,N_5895,N_2756);
and U9214 (N_9214,N_2156,N_2016);
and U9215 (N_9215,N_2652,N_289);
or U9216 (N_9216,N_920,N_6080);
nand U9217 (N_9217,N_4537,N_1591);
and U9218 (N_9218,N_2496,N_4023);
or U9219 (N_9219,N_330,N_3777);
xnor U9220 (N_9220,N_3522,N_4105);
nor U9221 (N_9221,N_2292,N_3645);
nand U9222 (N_9222,N_1655,N_3721);
and U9223 (N_9223,N_4821,N_3954);
nor U9224 (N_9224,N_5837,N_3500);
and U9225 (N_9225,N_1885,N_6186);
nor U9226 (N_9226,N_4681,N_360);
nor U9227 (N_9227,N_5074,N_1156);
nand U9228 (N_9228,N_2786,N_74);
or U9229 (N_9229,N_1555,N_2076);
and U9230 (N_9230,N_5487,N_2340);
and U9231 (N_9231,N_5532,N_2905);
nor U9232 (N_9232,N_1876,N_851);
or U9233 (N_9233,N_5176,N_4536);
and U9234 (N_9234,N_2126,N_6205);
and U9235 (N_9235,N_2638,N_5081);
and U9236 (N_9236,N_539,N_5145);
nor U9237 (N_9237,N_47,N_2368);
xnor U9238 (N_9238,N_4750,N_5834);
and U9239 (N_9239,N_2673,N_1231);
nand U9240 (N_9240,N_3791,N_3735);
nor U9241 (N_9241,N_3237,N_315);
nand U9242 (N_9242,N_940,N_3436);
nand U9243 (N_9243,N_4176,N_242);
nor U9244 (N_9244,N_3957,N_2128);
and U9245 (N_9245,N_2244,N_5493);
nor U9246 (N_9246,N_5462,N_6056);
and U9247 (N_9247,N_4635,N_3583);
or U9248 (N_9248,N_5687,N_3828);
and U9249 (N_9249,N_13,N_4233);
nor U9250 (N_9250,N_5307,N_2308);
nand U9251 (N_9251,N_815,N_5309);
and U9252 (N_9252,N_3186,N_4061);
and U9253 (N_9253,N_2653,N_1164);
and U9254 (N_9254,N_5422,N_4376);
or U9255 (N_9255,N_2986,N_4807);
and U9256 (N_9256,N_3445,N_622);
nand U9257 (N_9257,N_2468,N_2358);
nand U9258 (N_9258,N_3970,N_6151);
and U9259 (N_9259,N_2217,N_3003);
or U9260 (N_9260,N_5502,N_4674);
xnor U9261 (N_9261,N_2802,N_4860);
and U9262 (N_9262,N_3981,N_5055);
nand U9263 (N_9263,N_1720,N_2385);
nand U9264 (N_9264,N_1442,N_2367);
nor U9265 (N_9265,N_4906,N_4435);
xor U9266 (N_9266,N_4203,N_1606);
or U9267 (N_9267,N_5946,N_5292);
and U9268 (N_9268,N_1203,N_2204);
and U9269 (N_9269,N_6232,N_2545);
nand U9270 (N_9270,N_1935,N_2915);
or U9271 (N_9271,N_411,N_2949);
or U9272 (N_9272,N_3628,N_6127);
nand U9273 (N_9273,N_5336,N_1181);
nand U9274 (N_9274,N_808,N_5916);
or U9275 (N_9275,N_2559,N_3783);
nor U9276 (N_9276,N_2897,N_2835);
and U9277 (N_9277,N_2844,N_5928);
xor U9278 (N_9278,N_6090,N_220);
nor U9279 (N_9279,N_614,N_2403);
or U9280 (N_9280,N_1567,N_688);
nor U9281 (N_9281,N_3757,N_210);
nor U9282 (N_9282,N_6027,N_6109);
or U9283 (N_9283,N_5084,N_3406);
xor U9284 (N_9284,N_541,N_2933);
xnor U9285 (N_9285,N_4834,N_2019);
nor U9286 (N_9286,N_1208,N_3140);
or U9287 (N_9287,N_5844,N_4959);
nor U9288 (N_9288,N_885,N_5168);
nor U9289 (N_9289,N_4585,N_1795);
and U9290 (N_9290,N_4249,N_5337);
or U9291 (N_9291,N_1207,N_5973);
nor U9292 (N_9292,N_5360,N_852);
nor U9293 (N_9293,N_879,N_2143);
nand U9294 (N_9294,N_1723,N_117);
and U9295 (N_9295,N_713,N_4151);
xnor U9296 (N_9296,N_222,N_4385);
and U9297 (N_9297,N_971,N_1959);
and U9298 (N_9298,N_3038,N_1779);
or U9299 (N_9299,N_2322,N_5217);
or U9300 (N_9300,N_3715,N_3964);
xnor U9301 (N_9301,N_2060,N_3963);
nand U9302 (N_9302,N_2112,N_5040);
and U9303 (N_9303,N_1,N_4679);
and U9304 (N_9304,N_5013,N_1974);
nor U9305 (N_9305,N_3730,N_3763);
and U9306 (N_9306,N_1754,N_5572);
nor U9307 (N_9307,N_1481,N_1137);
nand U9308 (N_9308,N_1418,N_4418);
and U9309 (N_9309,N_4450,N_2250);
nor U9310 (N_9310,N_2832,N_4962);
nand U9311 (N_9311,N_4099,N_4361);
nor U9312 (N_9312,N_6176,N_3451);
or U9313 (N_9313,N_6119,N_1619);
and U9314 (N_9314,N_1883,N_1170);
nor U9315 (N_9315,N_5940,N_3834);
or U9316 (N_9316,N_68,N_5610);
nor U9317 (N_9317,N_3089,N_2309);
nor U9318 (N_9318,N_3553,N_1014);
or U9319 (N_9319,N_3563,N_4239);
nand U9320 (N_9320,N_5929,N_4984);
nand U9321 (N_9321,N_5680,N_3527);
nand U9322 (N_9322,N_5552,N_2214);
nand U9323 (N_9323,N_6075,N_5694);
and U9324 (N_9324,N_1752,N_2607);
nor U9325 (N_9325,N_4123,N_558);
or U9326 (N_9326,N_2131,N_5551);
xor U9327 (N_9327,N_316,N_1015);
and U9328 (N_9328,N_2431,N_5167);
nor U9329 (N_9329,N_2119,N_4868);
or U9330 (N_9330,N_3330,N_1888);
nor U9331 (N_9331,N_5151,N_3544);
xor U9332 (N_9332,N_1875,N_3139);
nand U9333 (N_9333,N_311,N_2597);
nand U9334 (N_9334,N_3221,N_2273);
or U9335 (N_9335,N_260,N_2836);
or U9336 (N_9336,N_5830,N_2166);
nand U9337 (N_9337,N_5766,N_862);
nor U9338 (N_9338,N_2904,N_1743);
nor U9339 (N_9339,N_4477,N_3371);
nand U9340 (N_9340,N_1781,N_1345);
nand U9341 (N_9341,N_1083,N_2061);
nand U9342 (N_9342,N_3554,N_5720);
nand U9343 (N_9343,N_2230,N_4986);
nor U9344 (N_9344,N_930,N_916);
or U9345 (N_9345,N_1073,N_1615);
xnor U9346 (N_9346,N_4432,N_1155);
or U9347 (N_9347,N_5843,N_3627);
or U9348 (N_9348,N_153,N_2661);
nand U9349 (N_9349,N_6210,N_5187);
nor U9350 (N_9350,N_159,N_1264);
and U9351 (N_9351,N_4267,N_1676);
and U9352 (N_9352,N_245,N_3257);
and U9353 (N_9353,N_829,N_124);
nor U9354 (N_9354,N_2177,N_4446);
nand U9355 (N_9355,N_2328,N_2220);
nor U9356 (N_9356,N_5206,N_923);
nor U9357 (N_9357,N_146,N_2605);
or U9358 (N_9358,N_1928,N_2670);
nand U9359 (N_9359,N_2213,N_3587);
or U9360 (N_9360,N_3176,N_820);
or U9361 (N_9361,N_4673,N_793);
or U9362 (N_9362,N_4597,N_4266);
nor U9363 (N_9363,N_5162,N_6078);
nand U9364 (N_9364,N_5554,N_1479);
nand U9365 (N_9365,N_6111,N_1482);
or U9366 (N_9366,N_1584,N_1843);
nor U9367 (N_9367,N_6133,N_3993);
nand U9368 (N_9368,N_5191,N_1166);
and U9369 (N_9369,N_1996,N_626);
or U9370 (N_9370,N_4919,N_4614);
xor U9371 (N_9371,N_905,N_4162);
xor U9372 (N_9372,N_6156,N_5142);
or U9373 (N_9373,N_588,N_4709);
and U9374 (N_9374,N_2826,N_1388);
nand U9375 (N_9375,N_3899,N_5427);
or U9376 (N_9376,N_2135,N_948);
xor U9377 (N_9377,N_2780,N_2615);
and U9378 (N_9378,N_503,N_3090);
nor U9379 (N_9379,N_1123,N_3807);
nor U9380 (N_9380,N_5870,N_69);
nand U9381 (N_9381,N_2677,N_3246);
and U9382 (N_9382,N_1826,N_1917);
or U9383 (N_9383,N_2242,N_5367);
nor U9384 (N_9384,N_5998,N_3383);
nor U9385 (N_9385,N_385,N_4953);
nand U9386 (N_9386,N_4026,N_3526);
nand U9387 (N_9387,N_1811,N_4162);
nand U9388 (N_9388,N_5118,N_4173);
or U9389 (N_9389,N_6195,N_3845);
or U9390 (N_9390,N_2116,N_4219);
and U9391 (N_9391,N_4219,N_2453);
nor U9392 (N_9392,N_4416,N_3937);
and U9393 (N_9393,N_6079,N_610);
or U9394 (N_9394,N_32,N_1311);
nor U9395 (N_9395,N_1546,N_5315);
nor U9396 (N_9396,N_5040,N_3308);
or U9397 (N_9397,N_2840,N_6018);
or U9398 (N_9398,N_2997,N_5504);
nor U9399 (N_9399,N_2387,N_4570);
nand U9400 (N_9400,N_1388,N_2113);
or U9401 (N_9401,N_643,N_141);
and U9402 (N_9402,N_5125,N_1820);
or U9403 (N_9403,N_6086,N_1749);
and U9404 (N_9404,N_3312,N_5540);
and U9405 (N_9405,N_1127,N_4830);
nand U9406 (N_9406,N_1670,N_5003);
xor U9407 (N_9407,N_1295,N_5575);
nand U9408 (N_9408,N_1855,N_3684);
nand U9409 (N_9409,N_3609,N_1109);
nor U9410 (N_9410,N_3842,N_5958);
or U9411 (N_9411,N_4438,N_5059);
nor U9412 (N_9412,N_3549,N_3180);
xnor U9413 (N_9413,N_4365,N_4207);
and U9414 (N_9414,N_2931,N_6147);
nor U9415 (N_9415,N_6129,N_2853);
xor U9416 (N_9416,N_271,N_3444);
xnor U9417 (N_9417,N_5680,N_3725);
nand U9418 (N_9418,N_3734,N_2498);
or U9419 (N_9419,N_230,N_141);
and U9420 (N_9420,N_2254,N_585);
or U9421 (N_9421,N_85,N_581);
or U9422 (N_9422,N_2327,N_4435);
nor U9423 (N_9423,N_48,N_3921);
nand U9424 (N_9424,N_2058,N_5363);
nand U9425 (N_9425,N_2233,N_1171);
or U9426 (N_9426,N_5168,N_6121);
nor U9427 (N_9427,N_1262,N_1955);
nand U9428 (N_9428,N_344,N_4005);
nor U9429 (N_9429,N_511,N_3908);
nand U9430 (N_9430,N_5489,N_3210);
and U9431 (N_9431,N_1226,N_2092);
nand U9432 (N_9432,N_6082,N_5878);
or U9433 (N_9433,N_3470,N_4561);
and U9434 (N_9434,N_996,N_2638);
or U9435 (N_9435,N_5732,N_2569);
and U9436 (N_9436,N_209,N_2884);
nand U9437 (N_9437,N_1082,N_1890);
or U9438 (N_9438,N_5100,N_1577);
nand U9439 (N_9439,N_992,N_2171);
nor U9440 (N_9440,N_1021,N_5914);
nor U9441 (N_9441,N_5906,N_3356);
nand U9442 (N_9442,N_3681,N_2005);
nand U9443 (N_9443,N_1087,N_1000);
and U9444 (N_9444,N_2909,N_930);
nor U9445 (N_9445,N_866,N_1963);
or U9446 (N_9446,N_6247,N_2658);
or U9447 (N_9447,N_3640,N_4338);
and U9448 (N_9448,N_1379,N_4571);
xor U9449 (N_9449,N_1630,N_2055);
xnor U9450 (N_9450,N_2631,N_3347);
nor U9451 (N_9451,N_2759,N_2028);
nor U9452 (N_9452,N_29,N_2208);
and U9453 (N_9453,N_6057,N_4077);
nand U9454 (N_9454,N_5007,N_5214);
xor U9455 (N_9455,N_2842,N_5242);
nor U9456 (N_9456,N_3725,N_4895);
nor U9457 (N_9457,N_6217,N_5495);
nand U9458 (N_9458,N_3021,N_1310);
nor U9459 (N_9459,N_4327,N_383);
nand U9460 (N_9460,N_60,N_1713);
nand U9461 (N_9461,N_1546,N_5314);
or U9462 (N_9462,N_5734,N_3256);
xor U9463 (N_9463,N_3603,N_4127);
nand U9464 (N_9464,N_550,N_1186);
nand U9465 (N_9465,N_1577,N_1997);
nor U9466 (N_9466,N_1991,N_5984);
nand U9467 (N_9467,N_4340,N_1405);
or U9468 (N_9468,N_1348,N_4245);
or U9469 (N_9469,N_2387,N_2081);
nor U9470 (N_9470,N_2114,N_2184);
or U9471 (N_9471,N_4758,N_2500);
nand U9472 (N_9472,N_370,N_3940);
xor U9473 (N_9473,N_1474,N_2586);
or U9474 (N_9474,N_5945,N_4492);
nand U9475 (N_9475,N_4070,N_3032);
xor U9476 (N_9476,N_2250,N_2357);
and U9477 (N_9477,N_2251,N_1463);
xnor U9478 (N_9478,N_5695,N_6086);
nor U9479 (N_9479,N_2849,N_815);
xnor U9480 (N_9480,N_2478,N_2839);
or U9481 (N_9481,N_1532,N_36);
or U9482 (N_9482,N_1751,N_4348);
xor U9483 (N_9483,N_1345,N_2644);
and U9484 (N_9484,N_4013,N_5681);
nor U9485 (N_9485,N_708,N_5696);
and U9486 (N_9486,N_24,N_5437);
and U9487 (N_9487,N_4734,N_648);
nor U9488 (N_9488,N_3355,N_5115);
nor U9489 (N_9489,N_779,N_3775);
and U9490 (N_9490,N_726,N_4310);
or U9491 (N_9491,N_5944,N_1492);
nand U9492 (N_9492,N_5822,N_6167);
nand U9493 (N_9493,N_1924,N_3001);
nand U9494 (N_9494,N_5467,N_4647);
xor U9495 (N_9495,N_1540,N_133);
nand U9496 (N_9496,N_4757,N_6067);
nand U9497 (N_9497,N_1129,N_1211);
or U9498 (N_9498,N_5889,N_5969);
or U9499 (N_9499,N_1115,N_5371);
xnor U9500 (N_9500,N_2167,N_3862);
nand U9501 (N_9501,N_5328,N_2192);
and U9502 (N_9502,N_5474,N_5762);
nand U9503 (N_9503,N_5970,N_1483);
and U9504 (N_9504,N_3381,N_4597);
nor U9505 (N_9505,N_4408,N_2371);
nor U9506 (N_9506,N_3544,N_3792);
and U9507 (N_9507,N_1835,N_4839);
nor U9508 (N_9508,N_307,N_4670);
xnor U9509 (N_9509,N_5379,N_5209);
nor U9510 (N_9510,N_2627,N_2854);
nand U9511 (N_9511,N_448,N_5395);
nor U9512 (N_9512,N_2449,N_6196);
nor U9513 (N_9513,N_5745,N_4831);
xnor U9514 (N_9514,N_3938,N_5482);
or U9515 (N_9515,N_668,N_4584);
nand U9516 (N_9516,N_4326,N_4177);
nor U9517 (N_9517,N_806,N_2729);
or U9518 (N_9518,N_4610,N_5087);
or U9519 (N_9519,N_6240,N_5897);
xor U9520 (N_9520,N_1889,N_759);
nand U9521 (N_9521,N_4098,N_3248);
or U9522 (N_9522,N_4009,N_1040);
nand U9523 (N_9523,N_3949,N_4256);
nand U9524 (N_9524,N_4830,N_4134);
or U9525 (N_9525,N_4354,N_4552);
or U9526 (N_9526,N_4702,N_3028);
and U9527 (N_9527,N_2335,N_4919);
and U9528 (N_9528,N_2985,N_2040);
or U9529 (N_9529,N_1678,N_2055);
xnor U9530 (N_9530,N_5957,N_3233);
nand U9531 (N_9531,N_4356,N_348);
or U9532 (N_9532,N_2208,N_1487);
or U9533 (N_9533,N_527,N_3661);
nand U9534 (N_9534,N_5026,N_181);
xor U9535 (N_9535,N_1160,N_5573);
and U9536 (N_9536,N_5197,N_3763);
nor U9537 (N_9537,N_7,N_2936);
and U9538 (N_9538,N_1218,N_1477);
xor U9539 (N_9539,N_5501,N_2750);
nand U9540 (N_9540,N_322,N_685);
and U9541 (N_9541,N_6129,N_2508);
nor U9542 (N_9542,N_1959,N_3103);
nor U9543 (N_9543,N_890,N_4864);
and U9544 (N_9544,N_582,N_1313);
or U9545 (N_9545,N_5268,N_644);
xor U9546 (N_9546,N_1682,N_5210);
or U9547 (N_9547,N_1892,N_4651);
nand U9548 (N_9548,N_2801,N_2235);
xor U9549 (N_9549,N_929,N_5007);
xnor U9550 (N_9550,N_5203,N_219);
nand U9551 (N_9551,N_604,N_401);
nor U9552 (N_9552,N_1965,N_4776);
or U9553 (N_9553,N_629,N_2127);
or U9554 (N_9554,N_2130,N_2616);
or U9555 (N_9555,N_1266,N_4398);
or U9556 (N_9556,N_4253,N_4163);
nor U9557 (N_9557,N_3731,N_2782);
or U9558 (N_9558,N_4698,N_5303);
or U9559 (N_9559,N_5577,N_3837);
or U9560 (N_9560,N_5347,N_3929);
and U9561 (N_9561,N_59,N_3631);
and U9562 (N_9562,N_4062,N_2272);
nor U9563 (N_9563,N_1663,N_5898);
and U9564 (N_9564,N_3353,N_3617);
or U9565 (N_9565,N_1609,N_3002);
xor U9566 (N_9566,N_5419,N_5797);
nor U9567 (N_9567,N_5482,N_3251);
nand U9568 (N_9568,N_4435,N_27);
nor U9569 (N_9569,N_3754,N_1629);
and U9570 (N_9570,N_2868,N_3055);
and U9571 (N_9571,N_42,N_5671);
or U9572 (N_9572,N_193,N_70);
xor U9573 (N_9573,N_654,N_4098);
nor U9574 (N_9574,N_539,N_4708);
and U9575 (N_9575,N_2418,N_5893);
and U9576 (N_9576,N_2451,N_251);
nor U9577 (N_9577,N_2307,N_5366);
xnor U9578 (N_9578,N_603,N_2109);
xnor U9579 (N_9579,N_159,N_2532);
or U9580 (N_9580,N_3414,N_784);
nor U9581 (N_9581,N_3907,N_364);
nand U9582 (N_9582,N_372,N_749);
nand U9583 (N_9583,N_5864,N_4169);
nor U9584 (N_9584,N_5890,N_1441);
nor U9585 (N_9585,N_821,N_1724);
or U9586 (N_9586,N_4039,N_5995);
or U9587 (N_9587,N_1828,N_1417);
nand U9588 (N_9588,N_1046,N_1036);
nor U9589 (N_9589,N_1086,N_1364);
nand U9590 (N_9590,N_2516,N_4726);
nor U9591 (N_9591,N_1265,N_3035);
nor U9592 (N_9592,N_3506,N_418);
or U9593 (N_9593,N_4015,N_2229);
nor U9594 (N_9594,N_4359,N_4693);
nand U9595 (N_9595,N_5409,N_935);
and U9596 (N_9596,N_5458,N_5930);
or U9597 (N_9597,N_2869,N_2909);
or U9598 (N_9598,N_2870,N_307);
nand U9599 (N_9599,N_5876,N_2229);
and U9600 (N_9600,N_3177,N_5653);
xnor U9601 (N_9601,N_1344,N_6097);
nand U9602 (N_9602,N_38,N_910);
and U9603 (N_9603,N_827,N_354);
and U9604 (N_9604,N_5579,N_2901);
or U9605 (N_9605,N_621,N_1658);
and U9606 (N_9606,N_108,N_5159);
xnor U9607 (N_9607,N_1879,N_3075);
or U9608 (N_9608,N_590,N_3850);
nor U9609 (N_9609,N_350,N_4436);
xor U9610 (N_9610,N_3244,N_1687);
and U9611 (N_9611,N_5879,N_1773);
and U9612 (N_9612,N_2155,N_5145);
and U9613 (N_9613,N_1474,N_5884);
or U9614 (N_9614,N_5809,N_5638);
nand U9615 (N_9615,N_5601,N_1144);
and U9616 (N_9616,N_3809,N_3352);
or U9617 (N_9617,N_4585,N_836);
and U9618 (N_9618,N_2518,N_5816);
and U9619 (N_9619,N_1074,N_334);
nand U9620 (N_9620,N_2094,N_3093);
and U9621 (N_9621,N_1830,N_3371);
and U9622 (N_9622,N_4448,N_2194);
nor U9623 (N_9623,N_1651,N_6093);
nor U9624 (N_9624,N_2307,N_3208);
and U9625 (N_9625,N_1080,N_3401);
and U9626 (N_9626,N_3302,N_4687);
and U9627 (N_9627,N_277,N_2273);
or U9628 (N_9628,N_735,N_82);
nor U9629 (N_9629,N_2283,N_2963);
and U9630 (N_9630,N_2276,N_17);
and U9631 (N_9631,N_1108,N_3725);
nor U9632 (N_9632,N_4419,N_927);
nand U9633 (N_9633,N_368,N_5205);
and U9634 (N_9634,N_4509,N_3755);
nand U9635 (N_9635,N_2415,N_2191);
and U9636 (N_9636,N_6166,N_244);
or U9637 (N_9637,N_556,N_4370);
xor U9638 (N_9638,N_6201,N_258);
or U9639 (N_9639,N_58,N_4994);
and U9640 (N_9640,N_363,N_4920);
and U9641 (N_9641,N_4052,N_4920);
and U9642 (N_9642,N_5585,N_917);
or U9643 (N_9643,N_862,N_1496);
and U9644 (N_9644,N_5122,N_3251);
nor U9645 (N_9645,N_5962,N_2786);
nand U9646 (N_9646,N_3374,N_91);
and U9647 (N_9647,N_1786,N_4508);
and U9648 (N_9648,N_4932,N_1880);
and U9649 (N_9649,N_5893,N_3487);
and U9650 (N_9650,N_529,N_1764);
and U9651 (N_9651,N_568,N_567);
and U9652 (N_9652,N_5635,N_5744);
or U9653 (N_9653,N_2573,N_989);
nand U9654 (N_9654,N_2310,N_2895);
or U9655 (N_9655,N_2629,N_338);
or U9656 (N_9656,N_350,N_4075);
and U9657 (N_9657,N_5041,N_3042);
or U9658 (N_9658,N_2102,N_1881);
nor U9659 (N_9659,N_3885,N_1642);
and U9660 (N_9660,N_5633,N_600);
or U9661 (N_9661,N_4837,N_774);
or U9662 (N_9662,N_1668,N_4015);
nor U9663 (N_9663,N_1106,N_1543);
and U9664 (N_9664,N_2185,N_2285);
and U9665 (N_9665,N_5997,N_511);
or U9666 (N_9666,N_5163,N_5679);
xnor U9667 (N_9667,N_2816,N_5072);
nor U9668 (N_9668,N_4722,N_4551);
xnor U9669 (N_9669,N_1068,N_2383);
xnor U9670 (N_9670,N_2431,N_735);
and U9671 (N_9671,N_1783,N_2145);
and U9672 (N_9672,N_41,N_3165);
nand U9673 (N_9673,N_4782,N_2271);
nor U9674 (N_9674,N_2749,N_1829);
nand U9675 (N_9675,N_5747,N_2445);
xor U9676 (N_9676,N_2293,N_710);
or U9677 (N_9677,N_126,N_4092);
or U9678 (N_9678,N_4506,N_3390);
nand U9679 (N_9679,N_3225,N_3336);
nor U9680 (N_9680,N_408,N_3118);
or U9681 (N_9681,N_5530,N_5220);
or U9682 (N_9682,N_2595,N_1277);
nand U9683 (N_9683,N_4706,N_2280);
nand U9684 (N_9684,N_154,N_6064);
and U9685 (N_9685,N_2203,N_5840);
nor U9686 (N_9686,N_4753,N_3372);
nor U9687 (N_9687,N_1250,N_5559);
xnor U9688 (N_9688,N_4688,N_3119);
nor U9689 (N_9689,N_5971,N_5633);
nand U9690 (N_9690,N_5229,N_4864);
nor U9691 (N_9691,N_2461,N_5063);
nand U9692 (N_9692,N_4284,N_5004);
nand U9693 (N_9693,N_5181,N_365);
nand U9694 (N_9694,N_2712,N_748);
nand U9695 (N_9695,N_4982,N_3242);
or U9696 (N_9696,N_6027,N_1911);
and U9697 (N_9697,N_2147,N_3104);
or U9698 (N_9698,N_75,N_4955);
nand U9699 (N_9699,N_105,N_3009);
nand U9700 (N_9700,N_4756,N_2771);
or U9701 (N_9701,N_814,N_1795);
nor U9702 (N_9702,N_5227,N_1417);
xnor U9703 (N_9703,N_1043,N_1778);
nand U9704 (N_9704,N_2993,N_2024);
nand U9705 (N_9705,N_1984,N_4333);
or U9706 (N_9706,N_4784,N_400);
and U9707 (N_9707,N_1584,N_5610);
or U9708 (N_9708,N_2059,N_3594);
or U9709 (N_9709,N_3583,N_1087);
nand U9710 (N_9710,N_3058,N_247);
nand U9711 (N_9711,N_856,N_5016);
or U9712 (N_9712,N_325,N_4535);
nor U9713 (N_9713,N_5121,N_6140);
or U9714 (N_9714,N_999,N_1450);
or U9715 (N_9715,N_4916,N_2735);
nor U9716 (N_9716,N_2895,N_4942);
nor U9717 (N_9717,N_4438,N_5293);
and U9718 (N_9718,N_3397,N_290);
nand U9719 (N_9719,N_4069,N_174);
or U9720 (N_9720,N_6103,N_4355);
nand U9721 (N_9721,N_1844,N_1746);
and U9722 (N_9722,N_2664,N_2804);
nand U9723 (N_9723,N_3485,N_1860);
or U9724 (N_9724,N_2390,N_5198);
and U9725 (N_9725,N_1326,N_1107);
nand U9726 (N_9726,N_1220,N_3750);
and U9727 (N_9727,N_1982,N_876);
nor U9728 (N_9728,N_5417,N_2872);
and U9729 (N_9729,N_1919,N_221);
nand U9730 (N_9730,N_920,N_2847);
and U9731 (N_9731,N_2974,N_3553);
or U9732 (N_9732,N_3886,N_2947);
nand U9733 (N_9733,N_2199,N_3322);
and U9734 (N_9734,N_3231,N_498);
nor U9735 (N_9735,N_5851,N_4636);
xnor U9736 (N_9736,N_3864,N_5788);
and U9737 (N_9737,N_4535,N_5197);
nand U9738 (N_9738,N_6204,N_3001);
nor U9739 (N_9739,N_1834,N_5875);
nor U9740 (N_9740,N_3527,N_4502);
or U9741 (N_9741,N_1331,N_2727);
or U9742 (N_9742,N_4564,N_5366);
and U9743 (N_9743,N_4701,N_4742);
nor U9744 (N_9744,N_1276,N_1081);
nand U9745 (N_9745,N_1305,N_2416);
and U9746 (N_9746,N_5894,N_2403);
nand U9747 (N_9747,N_4877,N_2079);
nor U9748 (N_9748,N_5648,N_713);
nor U9749 (N_9749,N_5023,N_2281);
xor U9750 (N_9750,N_942,N_4003);
nand U9751 (N_9751,N_583,N_4056);
or U9752 (N_9752,N_1948,N_2634);
nor U9753 (N_9753,N_21,N_2070);
nand U9754 (N_9754,N_1323,N_5085);
nand U9755 (N_9755,N_2187,N_3049);
nand U9756 (N_9756,N_4835,N_3875);
nand U9757 (N_9757,N_1947,N_1941);
or U9758 (N_9758,N_4043,N_3421);
nand U9759 (N_9759,N_3801,N_478);
and U9760 (N_9760,N_916,N_1679);
or U9761 (N_9761,N_1714,N_1006);
nand U9762 (N_9762,N_5138,N_4974);
or U9763 (N_9763,N_5729,N_5022);
xor U9764 (N_9764,N_3004,N_3161);
or U9765 (N_9765,N_121,N_6053);
nand U9766 (N_9766,N_4058,N_2238);
nand U9767 (N_9767,N_6113,N_3087);
nor U9768 (N_9768,N_3397,N_1291);
and U9769 (N_9769,N_835,N_1007);
nor U9770 (N_9770,N_545,N_5214);
or U9771 (N_9771,N_515,N_1376);
nor U9772 (N_9772,N_1058,N_6191);
xor U9773 (N_9773,N_5413,N_6043);
xor U9774 (N_9774,N_671,N_2747);
nand U9775 (N_9775,N_1060,N_502);
and U9776 (N_9776,N_4768,N_1545);
or U9777 (N_9777,N_5406,N_5361);
or U9778 (N_9778,N_2907,N_3323);
nand U9779 (N_9779,N_2960,N_1430);
nor U9780 (N_9780,N_3033,N_5988);
xnor U9781 (N_9781,N_4492,N_5415);
and U9782 (N_9782,N_1192,N_3880);
nand U9783 (N_9783,N_673,N_1336);
or U9784 (N_9784,N_2965,N_3598);
xnor U9785 (N_9785,N_6244,N_2494);
and U9786 (N_9786,N_3376,N_4101);
and U9787 (N_9787,N_2104,N_412);
xnor U9788 (N_9788,N_901,N_1895);
and U9789 (N_9789,N_2031,N_1297);
nor U9790 (N_9790,N_3993,N_1832);
nor U9791 (N_9791,N_675,N_5535);
nor U9792 (N_9792,N_1648,N_2442);
xnor U9793 (N_9793,N_3332,N_4058);
nand U9794 (N_9794,N_4070,N_3697);
and U9795 (N_9795,N_3469,N_1606);
nand U9796 (N_9796,N_2460,N_4146);
and U9797 (N_9797,N_2253,N_910);
nand U9798 (N_9798,N_3645,N_2806);
or U9799 (N_9799,N_882,N_5289);
nand U9800 (N_9800,N_4769,N_1123);
nand U9801 (N_9801,N_2119,N_3653);
or U9802 (N_9802,N_2324,N_516);
nor U9803 (N_9803,N_2603,N_3488);
and U9804 (N_9804,N_2304,N_2814);
and U9805 (N_9805,N_2899,N_2844);
and U9806 (N_9806,N_3564,N_2359);
or U9807 (N_9807,N_2103,N_4489);
xnor U9808 (N_9808,N_3072,N_2409);
nand U9809 (N_9809,N_3654,N_4088);
and U9810 (N_9810,N_1249,N_4035);
and U9811 (N_9811,N_5574,N_5320);
xnor U9812 (N_9812,N_4919,N_5959);
nand U9813 (N_9813,N_4187,N_2314);
and U9814 (N_9814,N_1920,N_732);
xor U9815 (N_9815,N_4263,N_4298);
and U9816 (N_9816,N_3722,N_1618);
nor U9817 (N_9817,N_3498,N_5049);
nand U9818 (N_9818,N_5493,N_6085);
nor U9819 (N_9819,N_31,N_736);
and U9820 (N_9820,N_1979,N_1599);
nor U9821 (N_9821,N_5965,N_3004);
and U9822 (N_9822,N_538,N_2577);
nand U9823 (N_9823,N_1123,N_4668);
nor U9824 (N_9824,N_2471,N_153);
xnor U9825 (N_9825,N_4847,N_1380);
nand U9826 (N_9826,N_755,N_4116);
nand U9827 (N_9827,N_4935,N_4112);
xnor U9828 (N_9828,N_230,N_3198);
nand U9829 (N_9829,N_1147,N_5843);
nor U9830 (N_9830,N_3631,N_1233);
or U9831 (N_9831,N_592,N_1571);
or U9832 (N_9832,N_2791,N_761);
and U9833 (N_9833,N_2947,N_39);
and U9834 (N_9834,N_6104,N_1576);
or U9835 (N_9835,N_3006,N_2539);
or U9836 (N_9836,N_407,N_4552);
nor U9837 (N_9837,N_5050,N_3552);
or U9838 (N_9838,N_6129,N_5280);
nor U9839 (N_9839,N_5764,N_2778);
or U9840 (N_9840,N_4918,N_5868);
nor U9841 (N_9841,N_537,N_1181);
or U9842 (N_9842,N_5966,N_1990);
or U9843 (N_9843,N_2819,N_2673);
nor U9844 (N_9844,N_1913,N_4592);
nor U9845 (N_9845,N_5897,N_5214);
and U9846 (N_9846,N_3795,N_454);
or U9847 (N_9847,N_1192,N_5102);
and U9848 (N_9848,N_3713,N_1035);
or U9849 (N_9849,N_1181,N_3239);
nor U9850 (N_9850,N_5247,N_2030);
nor U9851 (N_9851,N_418,N_370);
nand U9852 (N_9852,N_6029,N_4907);
or U9853 (N_9853,N_1667,N_1968);
or U9854 (N_9854,N_4665,N_727);
nand U9855 (N_9855,N_1706,N_4712);
or U9856 (N_9856,N_2897,N_1391);
and U9857 (N_9857,N_2431,N_5775);
nand U9858 (N_9858,N_5713,N_4781);
nand U9859 (N_9859,N_4831,N_1689);
or U9860 (N_9860,N_5329,N_3443);
and U9861 (N_9861,N_4718,N_4532);
or U9862 (N_9862,N_4807,N_2277);
nor U9863 (N_9863,N_329,N_977);
xor U9864 (N_9864,N_5615,N_4716);
xnor U9865 (N_9865,N_4298,N_6232);
or U9866 (N_9866,N_5271,N_4467);
nor U9867 (N_9867,N_5710,N_6175);
or U9868 (N_9868,N_1350,N_2469);
nand U9869 (N_9869,N_5778,N_535);
xnor U9870 (N_9870,N_3290,N_2584);
or U9871 (N_9871,N_2567,N_1093);
and U9872 (N_9872,N_538,N_6078);
nor U9873 (N_9873,N_5328,N_2767);
and U9874 (N_9874,N_5386,N_459);
or U9875 (N_9875,N_6026,N_1877);
nand U9876 (N_9876,N_1983,N_5364);
or U9877 (N_9877,N_2976,N_2578);
xnor U9878 (N_9878,N_6087,N_1349);
or U9879 (N_9879,N_4806,N_4870);
nand U9880 (N_9880,N_4404,N_1429);
and U9881 (N_9881,N_2157,N_181);
or U9882 (N_9882,N_5507,N_5000);
nand U9883 (N_9883,N_80,N_254);
nand U9884 (N_9884,N_384,N_1964);
nor U9885 (N_9885,N_3352,N_5849);
and U9886 (N_9886,N_183,N_3787);
or U9887 (N_9887,N_1166,N_2077);
and U9888 (N_9888,N_3755,N_5838);
and U9889 (N_9889,N_3415,N_257);
or U9890 (N_9890,N_2753,N_297);
nand U9891 (N_9891,N_802,N_4530);
and U9892 (N_9892,N_1876,N_1157);
and U9893 (N_9893,N_1130,N_2257);
or U9894 (N_9894,N_3481,N_3161);
nor U9895 (N_9895,N_4564,N_806);
nor U9896 (N_9896,N_6228,N_739);
nand U9897 (N_9897,N_948,N_3355);
nand U9898 (N_9898,N_1472,N_5514);
nor U9899 (N_9899,N_1519,N_1236);
and U9900 (N_9900,N_4522,N_2410);
nand U9901 (N_9901,N_382,N_2834);
xnor U9902 (N_9902,N_532,N_2908);
nor U9903 (N_9903,N_266,N_2564);
xnor U9904 (N_9904,N_3477,N_131);
nor U9905 (N_9905,N_1196,N_1832);
nor U9906 (N_9906,N_4693,N_3085);
nor U9907 (N_9907,N_1457,N_4907);
nand U9908 (N_9908,N_2366,N_2105);
nand U9909 (N_9909,N_2695,N_2704);
nor U9910 (N_9910,N_961,N_962);
nand U9911 (N_9911,N_4234,N_269);
nand U9912 (N_9912,N_1008,N_2618);
nor U9913 (N_9913,N_2299,N_2758);
nor U9914 (N_9914,N_2139,N_1445);
nor U9915 (N_9915,N_3315,N_3058);
nor U9916 (N_9916,N_5420,N_4466);
nand U9917 (N_9917,N_2647,N_2885);
nor U9918 (N_9918,N_3644,N_4066);
nor U9919 (N_9919,N_5762,N_3931);
nor U9920 (N_9920,N_189,N_4918);
nor U9921 (N_9921,N_75,N_4934);
xnor U9922 (N_9922,N_1992,N_3093);
nand U9923 (N_9923,N_3990,N_3599);
nor U9924 (N_9924,N_5932,N_5490);
nand U9925 (N_9925,N_2424,N_4347);
xnor U9926 (N_9926,N_4456,N_918);
and U9927 (N_9927,N_5776,N_1244);
xnor U9928 (N_9928,N_5282,N_4630);
nor U9929 (N_9929,N_1015,N_29);
nand U9930 (N_9930,N_6088,N_2826);
nor U9931 (N_9931,N_854,N_5600);
nor U9932 (N_9932,N_4857,N_4425);
nand U9933 (N_9933,N_2335,N_6015);
or U9934 (N_9934,N_846,N_2658);
and U9935 (N_9935,N_841,N_1470);
or U9936 (N_9936,N_3265,N_55);
or U9937 (N_9937,N_689,N_1273);
and U9938 (N_9938,N_4514,N_3653);
nor U9939 (N_9939,N_376,N_4204);
nor U9940 (N_9940,N_3684,N_4843);
or U9941 (N_9941,N_847,N_1966);
or U9942 (N_9942,N_3761,N_5130);
or U9943 (N_9943,N_4014,N_621);
nor U9944 (N_9944,N_256,N_4845);
and U9945 (N_9945,N_2600,N_5105);
or U9946 (N_9946,N_1219,N_284);
and U9947 (N_9947,N_1319,N_5869);
or U9948 (N_9948,N_979,N_4434);
and U9949 (N_9949,N_4134,N_3355);
nand U9950 (N_9950,N_3949,N_407);
and U9951 (N_9951,N_1953,N_614);
or U9952 (N_9952,N_2159,N_5119);
xor U9953 (N_9953,N_4795,N_4797);
or U9954 (N_9954,N_6018,N_2299);
nor U9955 (N_9955,N_293,N_5891);
or U9956 (N_9956,N_3675,N_6030);
nand U9957 (N_9957,N_2005,N_1786);
nor U9958 (N_9958,N_2154,N_2411);
nor U9959 (N_9959,N_1876,N_3577);
nor U9960 (N_9960,N_3714,N_2130);
and U9961 (N_9961,N_108,N_3668);
nand U9962 (N_9962,N_2158,N_3500);
and U9963 (N_9963,N_5878,N_5961);
or U9964 (N_9964,N_1241,N_3941);
or U9965 (N_9965,N_4847,N_1446);
nor U9966 (N_9966,N_2802,N_1328);
nor U9967 (N_9967,N_3372,N_1330);
nand U9968 (N_9968,N_3611,N_117);
xor U9969 (N_9969,N_1643,N_954);
or U9970 (N_9970,N_5169,N_2468);
nand U9971 (N_9971,N_5394,N_4629);
nand U9972 (N_9972,N_3033,N_3528);
and U9973 (N_9973,N_405,N_5072);
nor U9974 (N_9974,N_6206,N_2661);
xnor U9975 (N_9975,N_1067,N_4635);
nor U9976 (N_9976,N_3332,N_5531);
or U9977 (N_9977,N_792,N_2028);
and U9978 (N_9978,N_6192,N_155);
or U9979 (N_9979,N_6180,N_1952);
xor U9980 (N_9980,N_1657,N_3035);
nor U9981 (N_9981,N_1311,N_5837);
nand U9982 (N_9982,N_688,N_5407);
xor U9983 (N_9983,N_4494,N_3150);
and U9984 (N_9984,N_3065,N_3750);
nand U9985 (N_9985,N_1650,N_1072);
nand U9986 (N_9986,N_964,N_1578);
xor U9987 (N_9987,N_1676,N_4349);
nand U9988 (N_9988,N_566,N_3560);
nor U9989 (N_9989,N_4777,N_4681);
and U9990 (N_9990,N_5379,N_2834);
nand U9991 (N_9991,N_3948,N_4016);
or U9992 (N_9992,N_1114,N_2620);
and U9993 (N_9993,N_1921,N_3796);
xnor U9994 (N_9994,N_770,N_3318);
nor U9995 (N_9995,N_2109,N_5054);
nand U9996 (N_9996,N_5450,N_2547);
nand U9997 (N_9997,N_76,N_1353);
xnor U9998 (N_9998,N_3395,N_1226);
and U9999 (N_9999,N_4052,N_5603);
nor U10000 (N_10000,N_1076,N_2057);
and U10001 (N_10001,N_4721,N_6132);
or U10002 (N_10002,N_1296,N_593);
nor U10003 (N_10003,N_2750,N_2920);
nand U10004 (N_10004,N_4611,N_5108);
nand U10005 (N_10005,N_736,N_4305);
nor U10006 (N_10006,N_1167,N_204);
and U10007 (N_10007,N_1364,N_484);
nand U10008 (N_10008,N_5372,N_4259);
or U10009 (N_10009,N_6065,N_1694);
or U10010 (N_10010,N_4574,N_1841);
nand U10011 (N_10011,N_4256,N_4913);
xor U10012 (N_10012,N_4591,N_5142);
nor U10013 (N_10013,N_1900,N_4656);
and U10014 (N_10014,N_1718,N_640);
or U10015 (N_10015,N_1068,N_2587);
nor U10016 (N_10016,N_4997,N_1389);
or U10017 (N_10017,N_5715,N_6095);
nand U10018 (N_10018,N_4358,N_5853);
nand U10019 (N_10019,N_3852,N_3859);
or U10020 (N_10020,N_4578,N_1190);
and U10021 (N_10021,N_5635,N_2497);
xnor U10022 (N_10022,N_4043,N_2072);
or U10023 (N_10023,N_4083,N_4348);
nand U10024 (N_10024,N_2891,N_6069);
and U10025 (N_10025,N_5812,N_352);
and U10026 (N_10026,N_1434,N_4005);
nor U10027 (N_10027,N_4408,N_3854);
or U10028 (N_10028,N_1515,N_6021);
nor U10029 (N_10029,N_5653,N_5673);
xor U10030 (N_10030,N_3270,N_64);
nor U10031 (N_10031,N_5005,N_4037);
nand U10032 (N_10032,N_8,N_342);
and U10033 (N_10033,N_3456,N_2280);
xor U10034 (N_10034,N_124,N_1401);
nand U10035 (N_10035,N_12,N_5806);
and U10036 (N_10036,N_4646,N_3847);
or U10037 (N_10037,N_3397,N_5814);
and U10038 (N_10038,N_2868,N_4700);
and U10039 (N_10039,N_5491,N_3126);
nand U10040 (N_10040,N_3336,N_2159);
nand U10041 (N_10041,N_4797,N_157);
or U10042 (N_10042,N_3708,N_4744);
or U10043 (N_10043,N_1773,N_276);
nand U10044 (N_10044,N_3083,N_870);
xor U10045 (N_10045,N_1028,N_1702);
nand U10046 (N_10046,N_3583,N_3257);
or U10047 (N_10047,N_5910,N_4059);
and U10048 (N_10048,N_243,N_1373);
nor U10049 (N_10049,N_2365,N_5092);
xnor U10050 (N_10050,N_2234,N_2254);
nor U10051 (N_10051,N_402,N_4732);
nand U10052 (N_10052,N_1410,N_4037);
nor U10053 (N_10053,N_4547,N_880);
and U10054 (N_10054,N_4043,N_6187);
or U10055 (N_10055,N_3053,N_969);
nor U10056 (N_10056,N_3870,N_3479);
and U10057 (N_10057,N_161,N_5997);
and U10058 (N_10058,N_4547,N_5445);
nand U10059 (N_10059,N_2700,N_1018);
nand U10060 (N_10060,N_4311,N_3441);
or U10061 (N_10061,N_6095,N_4676);
nor U10062 (N_10062,N_734,N_4686);
nor U10063 (N_10063,N_3115,N_5462);
nand U10064 (N_10064,N_4906,N_2565);
or U10065 (N_10065,N_2307,N_2145);
nand U10066 (N_10066,N_2117,N_5275);
and U10067 (N_10067,N_4825,N_2103);
and U10068 (N_10068,N_3480,N_5160);
nand U10069 (N_10069,N_1854,N_2831);
or U10070 (N_10070,N_5201,N_3451);
and U10071 (N_10071,N_4950,N_2767);
nand U10072 (N_10072,N_3161,N_3060);
nand U10073 (N_10073,N_321,N_300);
nor U10074 (N_10074,N_4180,N_2171);
nor U10075 (N_10075,N_4459,N_3964);
nand U10076 (N_10076,N_4718,N_2730);
nand U10077 (N_10077,N_1526,N_5299);
nand U10078 (N_10078,N_6155,N_4863);
nor U10079 (N_10079,N_6078,N_1452);
or U10080 (N_10080,N_6122,N_4989);
nor U10081 (N_10081,N_551,N_550);
and U10082 (N_10082,N_6172,N_4611);
and U10083 (N_10083,N_782,N_2393);
and U10084 (N_10084,N_5443,N_3511);
or U10085 (N_10085,N_1924,N_5095);
or U10086 (N_10086,N_4079,N_1439);
xnor U10087 (N_10087,N_3246,N_2457);
nor U10088 (N_10088,N_749,N_4979);
and U10089 (N_10089,N_5459,N_5382);
nor U10090 (N_10090,N_4393,N_4146);
nor U10091 (N_10091,N_233,N_676);
and U10092 (N_10092,N_344,N_1391);
or U10093 (N_10093,N_597,N_5203);
or U10094 (N_10094,N_5034,N_1867);
nand U10095 (N_10095,N_5072,N_1514);
and U10096 (N_10096,N_1903,N_3345);
or U10097 (N_10097,N_384,N_4407);
nand U10098 (N_10098,N_4958,N_1711);
and U10099 (N_10099,N_2043,N_3455);
or U10100 (N_10100,N_3271,N_1212);
or U10101 (N_10101,N_1656,N_3687);
nor U10102 (N_10102,N_4636,N_413);
nand U10103 (N_10103,N_3031,N_701);
or U10104 (N_10104,N_4849,N_4356);
or U10105 (N_10105,N_4164,N_3810);
xor U10106 (N_10106,N_940,N_4386);
and U10107 (N_10107,N_2838,N_752);
or U10108 (N_10108,N_1142,N_2860);
or U10109 (N_10109,N_1965,N_5438);
xnor U10110 (N_10110,N_3449,N_4539);
nand U10111 (N_10111,N_760,N_5577);
nand U10112 (N_10112,N_3468,N_2046);
nand U10113 (N_10113,N_353,N_2366);
xnor U10114 (N_10114,N_3632,N_6080);
xor U10115 (N_10115,N_4656,N_2843);
nor U10116 (N_10116,N_385,N_416);
and U10117 (N_10117,N_4398,N_2110);
nor U10118 (N_10118,N_3210,N_5692);
or U10119 (N_10119,N_443,N_5410);
or U10120 (N_10120,N_753,N_3350);
or U10121 (N_10121,N_5564,N_2843);
nand U10122 (N_10122,N_3572,N_473);
or U10123 (N_10123,N_5890,N_3427);
nor U10124 (N_10124,N_3672,N_957);
nor U10125 (N_10125,N_3806,N_2478);
xnor U10126 (N_10126,N_5902,N_599);
or U10127 (N_10127,N_1735,N_3790);
nor U10128 (N_10128,N_6111,N_3485);
or U10129 (N_10129,N_888,N_3863);
nand U10130 (N_10130,N_2521,N_5007);
nor U10131 (N_10131,N_4408,N_1909);
nor U10132 (N_10132,N_656,N_245);
nand U10133 (N_10133,N_1983,N_5366);
and U10134 (N_10134,N_840,N_188);
xnor U10135 (N_10135,N_3831,N_3216);
xnor U10136 (N_10136,N_5531,N_5660);
nand U10137 (N_10137,N_2025,N_594);
nor U10138 (N_10138,N_908,N_2815);
and U10139 (N_10139,N_3032,N_4146);
and U10140 (N_10140,N_2544,N_3578);
nor U10141 (N_10141,N_4352,N_1563);
nor U10142 (N_10142,N_5422,N_4878);
nand U10143 (N_10143,N_2979,N_673);
or U10144 (N_10144,N_4395,N_636);
nand U10145 (N_10145,N_2123,N_1324);
and U10146 (N_10146,N_1665,N_245);
nand U10147 (N_10147,N_1316,N_3406);
nor U10148 (N_10148,N_5487,N_5900);
or U10149 (N_10149,N_4204,N_1883);
and U10150 (N_10150,N_2833,N_2569);
xor U10151 (N_10151,N_4841,N_2035);
and U10152 (N_10152,N_5451,N_3370);
xor U10153 (N_10153,N_5325,N_2866);
or U10154 (N_10154,N_4782,N_386);
nand U10155 (N_10155,N_583,N_4594);
and U10156 (N_10156,N_5380,N_5736);
nand U10157 (N_10157,N_4169,N_3874);
nand U10158 (N_10158,N_5682,N_2806);
nand U10159 (N_10159,N_841,N_2199);
nand U10160 (N_10160,N_1311,N_3970);
or U10161 (N_10161,N_3752,N_4825);
xor U10162 (N_10162,N_1003,N_4474);
nor U10163 (N_10163,N_493,N_3835);
nor U10164 (N_10164,N_1897,N_5654);
xor U10165 (N_10165,N_496,N_522);
and U10166 (N_10166,N_849,N_3445);
and U10167 (N_10167,N_1410,N_4480);
nor U10168 (N_10168,N_4887,N_3523);
xnor U10169 (N_10169,N_2678,N_729);
nor U10170 (N_10170,N_5473,N_293);
nor U10171 (N_10171,N_3035,N_5302);
or U10172 (N_10172,N_4557,N_4804);
or U10173 (N_10173,N_5956,N_3988);
nor U10174 (N_10174,N_3038,N_3226);
nor U10175 (N_10175,N_5782,N_5559);
or U10176 (N_10176,N_286,N_188);
xnor U10177 (N_10177,N_4526,N_4280);
xor U10178 (N_10178,N_1870,N_2041);
nor U10179 (N_10179,N_2471,N_3478);
nand U10180 (N_10180,N_4169,N_5663);
xnor U10181 (N_10181,N_5009,N_1747);
xnor U10182 (N_10182,N_1931,N_2776);
or U10183 (N_10183,N_5397,N_2350);
or U10184 (N_10184,N_85,N_5089);
and U10185 (N_10185,N_2496,N_3147);
nor U10186 (N_10186,N_5182,N_2790);
xnor U10187 (N_10187,N_1118,N_4225);
and U10188 (N_10188,N_3555,N_6098);
and U10189 (N_10189,N_3839,N_3691);
xor U10190 (N_10190,N_899,N_442);
nor U10191 (N_10191,N_5091,N_800);
and U10192 (N_10192,N_4918,N_2648);
and U10193 (N_10193,N_3193,N_587);
nand U10194 (N_10194,N_4715,N_548);
nand U10195 (N_10195,N_1556,N_1945);
or U10196 (N_10196,N_170,N_5149);
nor U10197 (N_10197,N_4510,N_2223);
xor U10198 (N_10198,N_1885,N_5518);
nand U10199 (N_10199,N_4363,N_4836);
and U10200 (N_10200,N_4175,N_5043);
and U10201 (N_10201,N_4952,N_1856);
and U10202 (N_10202,N_1364,N_3554);
and U10203 (N_10203,N_2985,N_1410);
and U10204 (N_10204,N_3610,N_2189);
nor U10205 (N_10205,N_1289,N_3290);
and U10206 (N_10206,N_4524,N_3304);
nor U10207 (N_10207,N_5115,N_2016);
nor U10208 (N_10208,N_2701,N_1936);
xor U10209 (N_10209,N_5436,N_2812);
xor U10210 (N_10210,N_5046,N_2473);
and U10211 (N_10211,N_3172,N_3894);
xnor U10212 (N_10212,N_4998,N_2694);
nand U10213 (N_10213,N_392,N_6075);
xor U10214 (N_10214,N_127,N_1065);
or U10215 (N_10215,N_5559,N_2203);
xor U10216 (N_10216,N_4865,N_159);
or U10217 (N_10217,N_2330,N_3071);
and U10218 (N_10218,N_3408,N_3522);
or U10219 (N_10219,N_2221,N_278);
nand U10220 (N_10220,N_5118,N_3102);
nand U10221 (N_10221,N_120,N_843);
nand U10222 (N_10222,N_3012,N_3976);
nor U10223 (N_10223,N_5648,N_3841);
or U10224 (N_10224,N_2490,N_847);
and U10225 (N_10225,N_4880,N_3244);
or U10226 (N_10226,N_5924,N_22);
nor U10227 (N_10227,N_616,N_3478);
nor U10228 (N_10228,N_381,N_4682);
or U10229 (N_10229,N_61,N_5263);
or U10230 (N_10230,N_3952,N_4994);
nand U10231 (N_10231,N_4177,N_2836);
and U10232 (N_10232,N_3782,N_5490);
nor U10233 (N_10233,N_2276,N_332);
nand U10234 (N_10234,N_5089,N_2542);
xnor U10235 (N_10235,N_488,N_2733);
and U10236 (N_10236,N_5272,N_5411);
and U10237 (N_10237,N_1310,N_1656);
nand U10238 (N_10238,N_6237,N_471);
nor U10239 (N_10239,N_505,N_1481);
and U10240 (N_10240,N_3189,N_4364);
or U10241 (N_10241,N_680,N_5583);
and U10242 (N_10242,N_80,N_675);
nor U10243 (N_10243,N_1196,N_4118);
nand U10244 (N_10244,N_3869,N_5316);
nor U10245 (N_10245,N_278,N_3460);
nor U10246 (N_10246,N_5585,N_125);
nor U10247 (N_10247,N_3226,N_4027);
nor U10248 (N_10248,N_6202,N_1925);
and U10249 (N_10249,N_5765,N_2126);
nand U10250 (N_10250,N_4693,N_4123);
nand U10251 (N_10251,N_2622,N_3908);
nor U10252 (N_10252,N_3634,N_2809);
or U10253 (N_10253,N_4471,N_3132);
nor U10254 (N_10254,N_883,N_1631);
nor U10255 (N_10255,N_5640,N_6197);
nand U10256 (N_10256,N_3333,N_5865);
or U10257 (N_10257,N_3950,N_54);
xor U10258 (N_10258,N_1356,N_788);
nor U10259 (N_10259,N_1405,N_4930);
or U10260 (N_10260,N_1043,N_929);
and U10261 (N_10261,N_5864,N_1248);
xor U10262 (N_10262,N_1150,N_4386);
and U10263 (N_10263,N_2049,N_2583);
xnor U10264 (N_10264,N_5407,N_1193);
and U10265 (N_10265,N_5487,N_4093);
and U10266 (N_10266,N_883,N_3683);
nand U10267 (N_10267,N_2707,N_1627);
or U10268 (N_10268,N_523,N_2070);
or U10269 (N_10269,N_4398,N_949);
and U10270 (N_10270,N_442,N_69);
xnor U10271 (N_10271,N_4808,N_389);
and U10272 (N_10272,N_2516,N_2310);
nor U10273 (N_10273,N_5281,N_963);
nand U10274 (N_10274,N_5079,N_5874);
nand U10275 (N_10275,N_435,N_5316);
or U10276 (N_10276,N_2225,N_2612);
nor U10277 (N_10277,N_2468,N_1089);
xnor U10278 (N_10278,N_5966,N_4965);
or U10279 (N_10279,N_3179,N_865);
nor U10280 (N_10280,N_3316,N_4098);
nand U10281 (N_10281,N_4127,N_5127);
nand U10282 (N_10282,N_1759,N_1778);
or U10283 (N_10283,N_3016,N_2656);
nand U10284 (N_10284,N_3935,N_2309);
nor U10285 (N_10285,N_4346,N_3259);
and U10286 (N_10286,N_2425,N_1679);
nand U10287 (N_10287,N_4768,N_1273);
xnor U10288 (N_10288,N_1708,N_5926);
and U10289 (N_10289,N_3267,N_1617);
and U10290 (N_10290,N_555,N_4940);
nor U10291 (N_10291,N_4474,N_5489);
nand U10292 (N_10292,N_4784,N_6019);
nor U10293 (N_10293,N_4612,N_290);
and U10294 (N_10294,N_3342,N_3796);
and U10295 (N_10295,N_302,N_4737);
nand U10296 (N_10296,N_1789,N_5954);
or U10297 (N_10297,N_5171,N_3559);
and U10298 (N_10298,N_942,N_3389);
nor U10299 (N_10299,N_291,N_5161);
nor U10300 (N_10300,N_5003,N_1374);
and U10301 (N_10301,N_844,N_5772);
nor U10302 (N_10302,N_5062,N_1631);
nor U10303 (N_10303,N_3761,N_839);
xnor U10304 (N_10304,N_2314,N_5840);
xnor U10305 (N_10305,N_970,N_719);
or U10306 (N_10306,N_1197,N_413);
nand U10307 (N_10307,N_3638,N_2860);
and U10308 (N_10308,N_5431,N_2133);
nor U10309 (N_10309,N_1023,N_2982);
nand U10310 (N_10310,N_3221,N_5859);
or U10311 (N_10311,N_5474,N_5657);
and U10312 (N_10312,N_6141,N_3364);
nor U10313 (N_10313,N_2162,N_4979);
or U10314 (N_10314,N_5602,N_187);
or U10315 (N_10315,N_1547,N_2273);
nand U10316 (N_10316,N_1317,N_348);
or U10317 (N_10317,N_1654,N_4152);
nand U10318 (N_10318,N_5838,N_3539);
nand U10319 (N_10319,N_3,N_1537);
nand U10320 (N_10320,N_4843,N_3857);
xor U10321 (N_10321,N_4953,N_885);
nand U10322 (N_10322,N_3786,N_1350);
and U10323 (N_10323,N_284,N_2476);
and U10324 (N_10324,N_3014,N_769);
or U10325 (N_10325,N_2690,N_222);
and U10326 (N_10326,N_3079,N_229);
nor U10327 (N_10327,N_2052,N_4030);
nand U10328 (N_10328,N_799,N_6027);
xnor U10329 (N_10329,N_53,N_6208);
nand U10330 (N_10330,N_2288,N_2940);
nor U10331 (N_10331,N_200,N_3095);
or U10332 (N_10332,N_862,N_2443);
xor U10333 (N_10333,N_1679,N_1856);
nand U10334 (N_10334,N_6233,N_1564);
xnor U10335 (N_10335,N_4194,N_5321);
nor U10336 (N_10336,N_3693,N_4814);
nor U10337 (N_10337,N_2327,N_5378);
nand U10338 (N_10338,N_2451,N_4380);
or U10339 (N_10339,N_1427,N_1945);
and U10340 (N_10340,N_233,N_4483);
or U10341 (N_10341,N_4886,N_3840);
or U10342 (N_10342,N_1744,N_215);
nand U10343 (N_10343,N_1178,N_1397);
or U10344 (N_10344,N_4091,N_1109);
nand U10345 (N_10345,N_4162,N_323);
and U10346 (N_10346,N_5549,N_5303);
nand U10347 (N_10347,N_156,N_5749);
nor U10348 (N_10348,N_4289,N_957);
or U10349 (N_10349,N_1874,N_4604);
nand U10350 (N_10350,N_2588,N_2141);
xor U10351 (N_10351,N_5820,N_3377);
and U10352 (N_10352,N_5050,N_4266);
xor U10353 (N_10353,N_2066,N_4287);
and U10354 (N_10354,N_876,N_4847);
nand U10355 (N_10355,N_690,N_579);
nand U10356 (N_10356,N_780,N_3086);
nand U10357 (N_10357,N_5929,N_3122);
and U10358 (N_10358,N_5956,N_2403);
or U10359 (N_10359,N_3791,N_4516);
and U10360 (N_10360,N_309,N_3670);
and U10361 (N_10361,N_5854,N_911);
nand U10362 (N_10362,N_1165,N_2630);
and U10363 (N_10363,N_3082,N_5988);
nor U10364 (N_10364,N_4186,N_1037);
nor U10365 (N_10365,N_4168,N_3993);
or U10366 (N_10366,N_857,N_1920);
and U10367 (N_10367,N_5633,N_6050);
nand U10368 (N_10368,N_4854,N_2175);
nor U10369 (N_10369,N_2732,N_2684);
nor U10370 (N_10370,N_498,N_3086);
and U10371 (N_10371,N_5875,N_881);
and U10372 (N_10372,N_4179,N_1049);
or U10373 (N_10373,N_654,N_5875);
nor U10374 (N_10374,N_799,N_2205);
or U10375 (N_10375,N_293,N_5862);
and U10376 (N_10376,N_5260,N_3682);
nand U10377 (N_10377,N_5222,N_2623);
and U10378 (N_10378,N_6068,N_5681);
and U10379 (N_10379,N_3522,N_4256);
nor U10380 (N_10380,N_1564,N_2594);
or U10381 (N_10381,N_4644,N_4291);
nor U10382 (N_10382,N_4081,N_3344);
and U10383 (N_10383,N_217,N_1770);
nand U10384 (N_10384,N_5517,N_3363);
xor U10385 (N_10385,N_2944,N_5687);
nand U10386 (N_10386,N_4732,N_2215);
or U10387 (N_10387,N_1080,N_2306);
nor U10388 (N_10388,N_3268,N_4204);
nor U10389 (N_10389,N_1877,N_2926);
nand U10390 (N_10390,N_3818,N_218);
or U10391 (N_10391,N_817,N_776);
xnor U10392 (N_10392,N_216,N_3455);
and U10393 (N_10393,N_4985,N_812);
nor U10394 (N_10394,N_4536,N_1921);
xnor U10395 (N_10395,N_4330,N_4674);
and U10396 (N_10396,N_3562,N_5451);
xor U10397 (N_10397,N_2352,N_3810);
or U10398 (N_10398,N_1161,N_5210);
xor U10399 (N_10399,N_5746,N_2699);
or U10400 (N_10400,N_1431,N_2842);
and U10401 (N_10401,N_3192,N_3251);
nor U10402 (N_10402,N_2756,N_6245);
or U10403 (N_10403,N_2758,N_1056);
nor U10404 (N_10404,N_6036,N_2386);
nand U10405 (N_10405,N_4938,N_5565);
xor U10406 (N_10406,N_445,N_3962);
or U10407 (N_10407,N_1158,N_4191);
nor U10408 (N_10408,N_1431,N_6065);
or U10409 (N_10409,N_6242,N_1747);
nand U10410 (N_10410,N_4548,N_5702);
or U10411 (N_10411,N_5312,N_2231);
xor U10412 (N_10412,N_3001,N_5048);
and U10413 (N_10413,N_2777,N_515);
or U10414 (N_10414,N_3443,N_2873);
nor U10415 (N_10415,N_4186,N_2672);
and U10416 (N_10416,N_1329,N_675);
or U10417 (N_10417,N_1709,N_4717);
nor U10418 (N_10418,N_3172,N_2846);
nand U10419 (N_10419,N_1818,N_4463);
or U10420 (N_10420,N_2837,N_3607);
nand U10421 (N_10421,N_1615,N_4263);
nand U10422 (N_10422,N_5232,N_2705);
or U10423 (N_10423,N_3115,N_4351);
nor U10424 (N_10424,N_5084,N_5850);
nor U10425 (N_10425,N_4771,N_1473);
or U10426 (N_10426,N_4312,N_312);
and U10427 (N_10427,N_2044,N_4902);
nor U10428 (N_10428,N_1456,N_4951);
nand U10429 (N_10429,N_1928,N_4532);
nand U10430 (N_10430,N_1228,N_4130);
and U10431 (N_10431,N_3902,N_3179);
or U10432 (N_10432,N_399,N_3440);
and U10433 (N_10433,N_124,N_2343);
nor U10434 (N_10434,N_1702,N_2088);
nand U10435 (N_10435,N_4797,N_5569);
nor U10436 (N_10436,N_2641,N_1932);
and U10437 (N_10437,N_2476,N_1392);
nand U10438 (N_10438,N_288,N_1556);
and U10439 (N_10439,N_6228,N_2459);
and U10440 (N_10440,N_576,N_1267);
and U10441 (N_10441,N_951,N_3061);
or U10442 (N_10442,N_941,N_1989);
nor U10443 (N_10443,N_451,N_5889);
nand U10444 (N_10444,N_4555,N_3761);
or U10445 (N_10445,N_1659,N_2171);
nor U10446 (N_10446,N_3394,N_1639);
nand U10447 (N_10447,N_2277,N_6220);
nand U10448 (N_10448,N_4274,N_32);
nor U10449 (N_10449,N_4210,N_2955);
and U10450 (N_10450,N_291,N_4738);
nand U10451 (N_10451,N_2079,N_3500);
or U10452 (N_10452,N_4362,N_869);
or U10453 (N_10453,N_266,N_1053);
or U10454 (N_10454,N_2217,N_1611);
nand U10455 (N_10455,N_1393,N_785);
nand U10456 (N_10456,N_3328,N_3138);
and U10457 (N_10457,N_1189,N_1933);
nand U10458 (N_10458,N_5242,N_2240);
nor U10459 (N_10459,N_5075,N_4524);
nor U10460 (N_10460,N_2461,N_5759);
or U10461 (N_10461,N_1497,N_4591);
and U10462 (N_10462,N_4885,N_4488);
xnor U10463 (N_10463,N_2251,N_1669);
or U10464 (N_10464,N_1281,N_5965);
nand U10465 (N_10465,N_1108,N_2248);
and U10466 (N_10466,N_2999,N_5034);
and U10467 (N_10467,N_1335,N_553);
or U10468 (N_10468,N_4532,N_1906);
and U10469 (N_10469,N_3706,N_3249);
xnor U10470 (N_10470,N_3045,N_3897);
xor U10471 (N_10471,N_629,N_5204);
nor U10472 (N_10472,N_23,N_441);
nor U10473 (N_10473,N_6094,N_3451);
and U10474 (N_10474,N_3826,N_5934);
or U10475 (N_10475,N_4449,N_2733);
or U10476 (N_10476,N_3278,N_2147);
nand U10477 (N_10477,N_1780,N_2117);
nor U10478 (N_10478,N_759,N_6064);
and U10479 (N_10479,N_523,N_5825);
nand U10480 (N_10480,N_677,N_2808);
and U10481 (N_10481,N_1656,N_1150);
nand U10482 (N_10482,N_2309,N_4462);
or U10483 (N_10483,N_906,N_3001);
nor U10484 (N_10484,N_454,N_628);
or U10485 (N_10485,N_3874,N_2861);
xnor U10486 (N_10486,N_2838,N_4046);
nand U10487 (N_10487,N_4086,N_1278);
xor U10488 (N_10488,N_1491,N_5740);
and U10489 (N_10489,N_230,N_2186);
nor U10490 (N_10490,N_315,N_5259);
xor U10491 (N_10491,N_2273,N_447);
or U10492 (N_10492,N_1377,N_3571);
or U10493 (N_10493,N_6200,N_1411);
nor U10494 (N_10494,N_2829,N_678);
or U10495 (N_10495,N_676,N_780);
nor U10496 (N_10496,N_6170,N_374);
or U10497 (N_10497,N_4248,N_4359);
and U10498 (N_10498,N_5416,N_936);
and U10499 (N_10499,N_6092,N_6137);
nand U10500 (N_10500,N_3263,N_5245);
nand U10501 (N_10501,N_1858,N_6150);
xnor U10502 (N_10502,N_5043,N_585);
nand U10503 (N_10503,N_3648,N_1961);
or U10504 (N_10504,N_899,N_3408);
xnor U10505 (N_10505,N_5399,N_1380);
and U10506 (N_10506,N_202,N_3836);
or U10507 (N_10507,N_5398,N_5207);
or U10508 (N_10508,N_4948,N_1442);
nand U10509 (N_10509,N_4816,N_2968);
and U10510 (N_10510,N_4156,N_4418);
nor U10511 (N_10511,N_4752,N_2908);
nor U10512 (N_10512,N_756,N_5753);
nand U10513 (N_10513,N_5925,N_1589);
and U10514 (N_10514,N_4694,N_1327);
nor U10515 (N_10515,N_3555,N_2924);
nor U10516 (N_10516,N_1731,N_3558);
xnor U10517 (N_10517,N_2212,N_2881);
and U10518 (N_10518,N_6136,N_3049);
or U10519 (N_10519,N_387,N_6248);
and U10520 (N_10520,N_5895,N_2702);
nand U10521 (N_10521,N_505,N_2655);
nand U10522 (N_10522,N_4023,N_994);
and U10523 (N_10523,N_69,N_1365);
nor U10524 (N_10524,N_5360,N_5436);
and U10525 (N_10525,N_1294,N_3132);
nor U10526 (N_10526,N_3432,N_1495);
or U10527 (N_10527,N_2305,N_5992);
nor U10528 (N_10528,N_3140,N_2753);
nor U10529 (N_10529,N_1127,N_1099);
nor U10530 (N_10530,N_6030,N_2762);
nor U10531 (N_10531,N_460,N_2534);
and U10532 (N_10532,N_4586,N_2057);
and U10533 (N_10533,N_3756,N_4214);
and U10534 (N_10534,N_4414,N_3122);
nor U10535 (N_10535,N_4715,N_2661);
nand U10536 (N_10536,N_3109,N_1011);
or U10537 (N_10537,N_2785,N_2779);
nor U10538 (N_10538,N_259,N_1873);
nor U10539 (N_10539,N_6108,N_3686);
or U10540 (N_10540,N_3499,N_244);
nor U10541 (N_10541,N_1756,N_1975);
nor U10542 (N_10542,N_1241,N_5830);
xor U10543 (N_10543,N_5376,N_437);
xor U10544 (N_10544,N_4588,N_1701);
nor U10545 (N_10545,N_5940,N_4854);
nand U10546 (N_10546,N_743,N_4345);
or U10547 (N_10547,N_305,N_2219);
xnor U10548 (N_10548,N_4545,N_5647);
nand U10549 (N_10549,N_1283,N_5517);
nand U10550 (N_10550,N_1192,N_5047);
nor U10551 (N_10551,N_717,N_4221);
nor U10552 (N_10552,N_5292,N_389);
xor U10553 (N_10553,N_12,N_47);
nor U10554 (N_10554,N_3162,N_2780);
nor U10555 (N_10555,N_1079,N_1700);
nor U10556 (N_10556,N_1976,N_1623);
or U10557 (N_10557,N_4892,N_5123);
or U10558 (N_10558,N_3180,N_3106);
nand U10559 (N_10559,N_955,N_86);
or U10560 (N_10560,N_4816,N_3005);
nor U10561 (N_10561,N_160,N_3773);
or U10562 (N_10562,N_5361,N_4631);
nor U10563 (N_10563,N_6034,N_4770);
nor U10564 (N_10564,N_4834,N_1750);
or U10565 (N_10565,N_4301,N_3271);
nand U10566 (N_10566,N_890,N_1261);
and U10567 (N_10567,N_2099,N_4266);
or U10568 (N_10568,N_895,N_4866);
nor U10569 (N_10569,N_2481,N_1059);
xnor U10570 (N_10570,N_287,N_5185);
nand U10571 (N_10571,N_772,N_1396);
xnor U10572 (N_10572,N_5336,N_4494);
nand U10573 (N_10573,N_1483,N_6208);
and U10574 (N_10574,N_27,N_2403);
nand U10575 (N_10575,N_5204,N_3451);
nor U10576 (N_10576,N_4865,N_4129);
nand U10577 (N_10577,N_2461,N_849);
nor U10578 (N_10578,N_2310,N_1025);
and U10579 (N_10579,N_955,N_5886);
nor U10580 (N_10580,N_5824,N_2150);
or U10581 (N_10581,N_5199,N_4472);
nand U10582 (N_10582,N_3524,N_5314);
or U10583 (N_10583,N_5135,N_4838);
nand U10584 (N_10584,N_4618,N_3333);
and U10585 (N_10585,N_3569,N_2376);
and U10586 (N_10586,N_1878,N_1060);
nor U10587 (N_10587,N_2263,N_2235);
nor U10588 (N_10588,N_1587,N_1700);
and U10589 (N_10589,N_850,N_60);
or U10590 (N_10590,N_3867,N_3740);
and U10591 (N_10591,N_4640,N_5852);
nand U10592 (N_10592,N_2321,N_164);
nor U10593 (N_10593,N_5099,N_5165);
or U10594 (N_10594,N_2356,N_4853);
xnor U10595 (N_10595,N_4227,N_6067);
and U10596 (N_10596,N_6154,N_5613);
nand U10597 (N_10597,N_4818,N_5323);
nand U10598 (N_10598,N_3329,N_5112);
nor U10599 (N_10599,N_664,N_61);
or U10600 (N_10600,N_444,N_1179);
nor U10601 (N_10601,N_2708,N_2914);
nand U10602 (N_10602,N_4874,N_1399);
nand U10603 (N_10603,N_3022,N_4245);
and U10604 (N_10604,N_3907,N_557);
nor U10605 (N_10605,N_256,N_763);
xor U10606 (N_10606,N_6181,N_1561);
nor U10607 (N_10607,N_1495,N_822);
or U10608 (N_10608,N_3010,N_1481);
nand U10609 (N_10609,N_4486,N_4232);
nand U10610 (N_10610,N_120,N_875);
and U10611 (N_10611,N_2054,N_386);
or U10612 (N_10612,N_2429,N_5856);
and U10613 (N_10613,N_2365,N_3259);
nor U10614 (N_10614,N_710,N_4905);
nand U10615 (N_10615,N_4274,N_6249);
xnor U10616 (N_10616,N_3604,N_5339);
nand U10617 (N_10617,N_5750,N_2842);
or U10618 (N_10618,N_3315,N_366);
nand U10619 (N_10619,N_1082,N_2997);
or U10620 (N_10620,N_3857,N_2437);
and U10621 (N_10621,N_5947,N_2247);
xor U10622 (N_10622,N_2575,N_3345);
nand U10623 (N_10623,N_4750,N_3521);
or U10624 (N_10624,N_2366,N_479);
xor U10625 (N_10625,N_1272,N_4436);
nor U10626 (N_10626,N_1129,N_1518);
and U10627 (N_10627,N_1777,N_3327);
and U10628 (N_10628,N_5928,N_1620);
nor U10629 (N_10629,N_1394,N_5482);
or U10630 (N_10630,N_794,N_4270);
xor U10631 (N_10631,N_463,N_1467);
or U10632 (N_10632,N_4806,N_5295);
and U10633 (N_10633,N_1349,N_3205);
nand U10634 (N_10634,N_3422,N_3081);
or U10635 (N_10635,N_4629,N_508);
or U10636 (N_10636,N_5434,N_2531);
nor U10637 (N_10637,N_3137,N_5491);
and U10638 (N_10638,N_5172,N_5718);
or U10639 (N_10639,N_2756,N_1141);
nor U10640 (N_10640,N_1728,N_3613);
nand U10641 (N_10641,N_5395,N_4638);
or U10642 (N_10642,N_1362,N_2873);
nor U10643 (N_10643,N_5173,N_3202);
nor U10644 (N_10644,N_2104,N_2619);
or U10645 (N_10645,N_891,N_2567);
or U10646 (N_10646,N_495,N_2754);
and U10647 (N_10647,N_1946,N_3599);
and U10648 (N_10648,N_5737,N_6127);
or U10649 (N_10649,N_5443,N_2686);
nand U10650 (N_10650,N_6080,N_5134);
nor U10651 (N_10651,N_579,N_2149);
or U10652 (N_10652,N_5778,N_5029);
nor U10653 (N_10653,N_344,N_412);
nand U10654 (N_10654,N_4557,N_2133);
and U10655 (N_10655,N_1744,N_1418);
nor U10656 (N_10656,N_6126,N_5018);
nand U10657 (N_10657,N_5536,N_6148);
nand U10658 (N_10658,N_2109,N_1956);
xnor U10659 (N_10659,N_224,N_84);
and U10660 (N_10660,N_4821,N_585);
nor U10661 (N_10661,N_3114,N_6034);
nand U10662 (N_10662,N_715,N_5667);
xor U10663 (N_10663,N_4081,N_382);
xor U10664 (N_10664,N_3425,N_4062);
nand U10665 (N_10665,N_5306,N_5446);
nand U10666 (N_10666,N_1848,N_3470);
nor U10667 (N_10667,N_4879,N_6142);
nand U10668 (N_10668,N_5677,N_385);
nor U10669 (N_10669,N_4800,N_231);
xnor U10670 (N_10670,N_670,N_2452);
xor U10671 (N_10671,N_3128,N_1273);
xor U10672 (N_10672,N_3966,N_2786);
nand U10673 (N_10673,N_4838,N_3655);
nor U10674 (N_10674,N_5611,N_4328);
nor U10675 (N_10675,N_4911,N_5851);
and U10676 (N_10676,N_3583,N_3500);
nor U10677 (N_10677,N_3846,N_2538);
or U10678 (N_10678,N_5036,N_5041);
nand U10679 (N_10679,N_1095,N_741);
nor U10680 (N_10680,N_4370,N_468);
or U10681 (N_10681,N_2141,N_233);
and U10682 (N_10682,N_3932,N_4579);
or U10683 (N_10683,N_4835,N_4128);
or U10684 (N_10684,N_5790,N_2905);
and U10685 (N_10685,N_823,N_4984);
and U10686 (N_10686,N_3263,N_4342);
nor U10687 (N_10687,N_3618,N_5720);
and U10688 (N_10688,N_5665,N_3821);
nand U10689 (N_10689,N_942,N_563);
and U10690 (N_10690,N_2215,N_4322);
nor U10691 (N_10691,N_2410,N_1033);
and U10692 (N_10692,N_3938,N_5842);
nand U10693 (N_10693,N_445,N_4495);
nand U10694 (N_10694,N_3210,N_2677);
nor U10695 (N_10695,N_5857,N_74);
or U10696 (N_10696,N_6135,N_2066);
or U10697 (N_10697,N_4339,N_6069);
and U10698 (N_10698,N_4278,N_2266);
or U10699 (N_10699,N_5738,N_6175);
xnor U10700 (N_10700,N_760,N_3444);
nand U10701 (N_10701,N_5682,N_6030);
and U10702 (N_10702,N_3786,N_2070);
nand U10703 (N_10703,N_3428,N_3891);
and U10704 (N_10704,N_3695,N_1028);
and U10705 (N_10705,N_4711,N_2704);
nor U10706 (N_10706,N_4538,N_3467);
xnor U10707 (N_10707,N_4220,N_2368);
nor U10708 (N_10708,N_2912,N_5646);
and U10709 (N_10709,N_718,N_3058);
and U10710 (N_10710,N_188,N_3208);
and U10711 (N_10711,N_2815,N_4862);
xor U10712 (N_10712,N_3016,N_1236);
or U10713 (N_10713,N_513,N_2841);
and U10714 (N_10714,N_4231,N_1180);
or U10715 (N_10715,N_2,N_2850);
or U10716 (N_10716,N_6088,N_2017);
nand U10717 (N_10717,N_49,N_2645);
or U10718 (N_10718,N_3725,N_5312);
xor U10719 (N_10719,N_965,N_752);
nor U10720 (N_10720,N_4390,N_664);
nor U10721 (N_10721,N_135,N_2443);
xor U10722 (N_10722,N_2539,N_6130);
xor U10723 (N_10723,N_829,N_5408);
or U10724 (N_10724,N_5865,N_3030);
nand U10725 (N_10725,N_2153,N_4095);
nand U10726 (N_10726,N_745,N_2373);
or U10727 (N_10727,N_3637,N_721);
and U10728 (N_10728,N_4250,N_4450);
nor U10729 (N_10729,N_2509,N_347);
xor U10730 (N_10730,N_506,N_5023);
or U10731 (N_10731,N_5057,N_2032);
nor U10732 (N_10732,N_5645,N_3502);
or U10733 (N_10733,N_4850,N_4396);
and U10734 (N_10734,N_440,N_3074);
xnor U10735 (N_10735,N_3012,N_1145);
nand U10736 (N_10736,N_2512,N_2929);
and U10737 (N_10737,N_761,N_5249);
nor U10738 (N_10738,N_3062,N_3611);
nand U10739 (N_10739,N_1499,N_424);
nand U10740 (N_10740,N_1588,N_3379);
and U10741 (N_10741,N_3850,N_5604);
xnor U10742 (N_10742,N_1269,N_1545);
nor U10743 (N_10743,N_3675,N_1165);
and U10744 (N_10744,N_348,N_3230);
or U10745 (N_10745,N_227,N_4511);
and U10746 (N_10746,N_616,N_5446);
and U10747 (N_10747,N_5124,N_1612);
nand U10748 (N_10748,N_2478,N_3533);
nand U10749 (N_10749,N_1131,N_1205);
and U10750 (N_10750,N_145,N_2270);
nor U10751 (N_10751,N_2614,N_1082);
or U10752 (N_10752,N_4775,N_2891);
or U10753 (N_10753,N_2433,N_1662);
xor U10754 (N_10754,N_2502,N_3686);
nor U10755 (N_10755,N_3071,N_3862);
nand U10756 (N_10756,N_11,N_2232);
xor U10757 (N_10757,N_433,N_505);
nand U10758 (N_10758,N_1144,N_683);
xor U10759 (N_10759,N_3898,N_1469);
and U10760 (N_10760,N_4720,N_3908);
nor U10761 (N_10761,N_2611,N_265);
and U10762 (N_10762,N_947,N_165);
nor U10763 (N_10763,N_5021,N_2381);
nor U10764 (N_10764,N_4698,N_3022);
nor U10765 (N_10765,N_365,N_5877);
or U10766 (N_10766,N_1670,N_1868);
nand U10767 (N_10767,N_3981,N_4126);
and U10768 (N_10768,N_2113,N_1565);
nor U10769 (N_10769,N_2451,N_3840);
nand U10770 (N_10770,N_3201,N_1179);
or U10771 (N_10771,N_5184,N_5395);
and U10772 (N_10772,N_618,N_2613);
or U10773 (N_10773,N_4877,N_2681);
nand U10774 (N_10774,N_3608,N_3210);
and U10775 (N_10775,N_3978,N_6194);
or U10776 (N_10776,N_6096,N_5480);
or U10777 (N_10777,N_4435,N_3105);
nor U10778 (N_10778,N_4603,N_4379);
or U10779 (N_10779,N_2635,N_4442);
nor U10780 (N_10780,N_3953,N_1238);
nor U10781 (N_10781,N_4752,N_5951);
or U10782 (N_10782,N_1641,N_5380);
nand U10783 (N_10783,N_2166,N_3808);
and U10784 (N_10784,N_336,N_3067);
nor U10785 (N_10785,N_4881,N_3837);
and U10786 (N_10786,N_3428,N_2896);
nor U10787 (N_10787,N_5337,N_2046);
nand U10788 (N_10788,N_5951,N_201);
or U10789 (N_10789,N_3762,N_2399);
nand U10790 (N_10790,N_6033,N_2809);
nor U10791 (N_10791,N_5360,N_1690);
nor U10792 (N_10792,N_105,N_5166);
nand U10793 (N_10793,N_819,N_1161);
xnor U10794 (N_10794,N_5179,N_5067);
or U10795 (N_10795,N_3905,N_5343);
and U10796 (N_10796,N_4993,N_19);
nand U10797 (N_10797,N_4592,N_2980);
and U10798 (N_10798,N_1518,N_2145);
nor U10799 (N_10799,N_51,N_4805);
and U10800 (N_10800,N_5040,N_4538);
or U10801 (N_10801,N_4946,N_358);
nor U10802 (N_10802,N_3327,N_2647);
nand U10803 (N_10803,N_1451,N_4780);
nor U10804 (N_10804,N_2595,N_2300);
nand U10805 (N_10805,N_239,N_2921);
nand U10806 (N_10806,N_2658,N_4228);
nor U10807 (N_10807,N_1856,N_3360);
nor U10808 (N_10808,N_3437,N_1688);
xor U10809 (N_10809,N_3823,N_6146);
nor U10810 (N_10810,N_2852,N_3757);
nor U10811 (N_10811,N_4674,N_4320);
and U10812 (N_10812,N_3881,N_337);
and U10813 (N_10813,N_5662,N_194);
nor U10814 (N_10814,N_1417,N_4742);
xor U10815 (N_10815,N_3208,N_4953);
nand U10816 (N_10816,N_1544,N_3040);
nand U10817 (N_10817,N_3722,N_2641);
or U10818 (N_10818,N_5715,N_87);
nand U10819 (N_10819,N_1038,N_3407);
nand U10820 (N_10820,N_4524,N_2073);
nand U10821 (N_10821,N_2929,N_225);
nand U10822 (N_10822,N_4094,N_184);
and U10823 (N_10823,N_3329,N_275);
and U10824 (N_10824,N_4938,N_4293);
nand U10825 (N_10825,N_3986,N_3416);
nor U10826 (N_10826,N_139,N_628);
nor U10827 (N_10827,N_1672,N_1312);
nand U10828 (N_10828,N_2988,N_4445);
nor U10829 (N_10829,N_5557,N_3471);
nor U10830 (N_10830,N_5110,N_2605);
nor U10831 (N_10831,N_4511,N_2807);
nand U10832 (N_10832,N_3387,N_2233);
nand U10833 (N_10833,N_1110,N_1605);
nor U10834 (N_10834,N_5799,N_4057);
nand U10835 (N_10835,N_5739,N_4307);
and U10836 (N_10836,N_2450,N_268);
and U10837 (N_10837,N_5184,N_820);
nor U10838 (N_10838,N_5942,N_1091);
nor U10839 (N_10839,N_3113,N_4448);
and U10840 (N_10840,N_3684,N_2119);
xor U10841 (N_10841,N_5400,N_4363);
or U10842 (N_10842,N_4263,N_4352);
nor U10843 (N_10843,N_4264,N_3804);
nand U10844 (N_10844,N_5272,N_2680);
and U10845 (N_10845,N_2491,N_525);
and U10846 (N_10846,N_5574,N_981);
xnor U10847 (N_10847,N_3239,N_953);
or U10848 (N_10848,N_2123,N_4295);
nand U10849 (N_10849,N_4466,N_5607);
xnor U10850 (N_10850,N_2898,N_4966);
nand U10851 (N_10851,N_5637,N_5816);
nand U10852 (N_10852,N_3384,N_1490);
nor U10853 (N_10853,N_3779,N_4944);
nand U10854 (N_10854,N_2160,N_5465);
nand U10855 (N_10855,N_6160,N_6101);
or U10856 (N_10856,N_1689,N_1635);
and U10857 (N_10857,N_4063,N_857);
and U10858 (N_10858,N_2741,N_5963);
nor U10859 (N_10859,N_2473,N_2764);
nor U10860 (N_10860,N_4942,N_4492);
nand U10861 (N_10861,N_4359,N_96);
nand U10862 (N_10862,N_5181,N_1551);
or U10863 (N_10863,N_2985,N_751);
xor U10864 (N_10864,N_2942,N_4607);
nor U10865 (N_10865,N_816,N_4975);
or U10866 (N_10866,N_3631,N_263);
xor U10867 (N_10867,N_399,N_3802);
nor U10868 (N_10868,N_3850,N_3917);
nand U10869 (N_10869,N_2146,N_4514);
nand U10870 (N_10870,N_926,N_385);
xor U10871 (N_10871,N_1254,N_3837);
and U10872 (N_10872,N_85,N_249);
nand U10873 (N_10873,N_3424,N_792);
nor U10874 (N_10874,N_387,N_5486);
xor U10875 (N_10875,N_4854,N_1282);
nand U10876 (N_10876,N_273,N_384);
nor U10877 (N_10877,N_4849,N_4568);
or U10878 (N_10878,N_2663,N_1158);
nand U10879 (N_10879,N_5837,N_5761);
nor U10880 (N_10880,N_1441,N_855);
or U10881 (N_10881,N_2709,N_4589);
or U10882 (N_10882,N_1949,N_1685);
and U10883 (N_10883,N_5478,N_2025);
xor U10884 (N_10884,N_5080,N_4289);
and U10885 (N_10885,N_3010,N_1248);
or U10886 (N_10886,N_4198,N_1426);
nand U10887 (N_10887,N_5268,N_990);
or U10888 (N_10888,N_2688,N_5791);
and U10889 (N_10889,N_56,N_3150);
nand U10890 (N_10890,N_1375,N_2404);
xnor U10891 (N_10891,N_4925,N_4614);
nor U10892 (N_10892,N_136,N_1092);
nand U10893 (N_10893,N_3565,N_4574);
nor U10894 (N_10894,N_5645,N_3137);
or U10895 (N_10895,N_4370,N_2980);
or U10896 (N_10896,N_4618,N_53);
xor U10897 (N_10897,N_185,N_439);
or U10898 (N_10898,N_5727,N_5122);
nand U10899 (N_10899,N_1377,N_1708);
or U10900 (N_10900,N_3762,N_1893);
nor U10901 (N_10901,N_5768,N_5019);
or U10902 (N_10902,N_5931,N_3705);
and U10903 (N_10903,N_136,N_4702);
nand U10904 (N_10904,N_2586,N_3328);
nand U10905 (N_10905,N_5641,N_1197);
nor U10906 (N_10906,N_4742,N_1774);
and U10907 (N_10907,N_1583,N_2868);
xor U10908 (N_10908,N_1187,N_6021);
and U10909 (N_10909,N_131,N_5334);
nor U10910 (N_10910,N_473,N_5208);
and U10911 (N_10911,N_2571,N_3958);
or U10912 (N_10912,N_5980,N_3457);
nor U10913 (N_10913,N_3149,N_519);
and U10914 (N_10914,N_932,N_5555);
nor U10915 (N_10915,N_487,N_22);
nand U10916 (N_10916,N_2,N_4088);
or U10917 (N_10917,N_1269,N_4728);
nor U10918 (N_10918,N_769,N_5348);
nand U10919 (N_10919,N_373,N_753);
and U10920 (N_10920,N_6061,N_3690);
and U10921 (N_10921,N_1394,N_1501);
nor U10922 (N_10922,N_2415,N_3137);
nand U10923 (N_10923,N_4254,N_4188);
nor U10924 (N_10924,N_5465,N_5395);
xnor U10925 (N_10925,N_73,N_2633);
nor U10926 (N_10926,N_3924,N_5746);
nand U10927 (N_10927,N_2103,N_3350);
or U10928 (N_10928,N_4488,N_2513);
xor U10929 (N_10929,N_2661,N_5564);
or U10930 (N_10930,N_1622,N_41);
or U10931 (N_10931,N_2652,N_512);
and U10932 (N_10932,N_4635,N_5055);
nor U10933 (N_10933,N_2113,N_1825);
nor U10934 (N_10934,N_4318,N_1169);
nor U10935 (N_10935,N_4338,N_1027);
nand U10936 (N_10936,N_4972,N_1819);
or U10937 (N_10937,N_3124,N_796);
or U10938 (N_10938,N_2047,N_3723);
or U10939 (N_10939,N_348,N_5702);
nor U10940 (N_10940,N_2845,N_3383);
xor U10941 (N_10941,N_2155,N_649);
nor U10942 (N_10942,N_2508,N_1588);
nor U10943 (N_10943,N_5102,N_1863);
nor U10944 (N_10944,N_2070,N_6093);
nor U10945 (N_10945,N_269,N_4769);
or U10946 (N_10946,N_3185,N_2041);
or U10947 (N_10947,N_753,N_6122);
nand U10948 (N_10948,N_5596,N_2777);
nor U10949 (N_10949,N_1470,N_2684);
nand U10950 (N_10950,N_432,N_4422);
nand U10951 (N_10951,N_2174,N_2356);
or U10952 (N_10952,N_5013,N_1377);
xor U10953 (N_10953,N_1214,N_6201);
nor U10954 (N_10954,N_3304,N_4034);
nor U10955 (N_10955,N_4501,N_2551);
nand U10956 (N_10956,N_3942,N_4504);
nor U10957 (N_10957,N_5836,N_3551);
and U10958 (N_10958,N_4561,N_213);
nand U10959 (N_10959,N_2444,N_4400);
or U10960 (N_10960,N_214,N_2429);
nand U10961 (N_10961,N_2672,N_2694);
nand U10962 (N_10962,N_3144,N_1805);
nor U10963 (N_10963,N_2257,N_3340);
nor U10964 (N_10964,N_66,N_283);
and U10965 (N_10965,N_4325,N_2943);
and U10966 (N_10966,N_5986,N_4380);
xor U10967 (N_10967,N_3057,N_3661);
and U10968 (N_10968,N_3943,N_2732);
nand U10969 (N_10969,N_424,N_2212);
nand U10970 (N_10970,N_3501,N_1303);
nor U10971 (N_10971,N_5876,N_6078);
nand U10972 (N_10972,N_256,N_2682);
xnor U10973 (N_10973,N_408,N_4196);
and U10974 (N_10974,N_3239,N_1657);
or U10975 (N_10975,N_2450,N_2148);
and U10976 (N_10976,N_3709,N_1564);
nor U10977 (N_10977,N_5426,N_1441);
nor U10978 (N_10978,N_6184,N_6077);
nand U10979 (N_10979,N_3647,N_2580);
and U10980 (N_10980,N_2465,N_4472);
nor U10981 (N_10981,N_2935,N_3083);
or U10982 (N_10982,N_350,N_304);
and U10983 (N_10983,N_1584,N_2555);
nand U10984 (N_10984,N_2959,N_2551);
and U10985 (N_10985,N_696,N_6246);
nor U10986 (N_10986,N_1416,N_6007);
and U10987 (N_10987,N_4970,N_3318);
nor U10988 (N_10988,N_921,N_5695);
or U10989 (N_10989,N_524,N_855);
xor U10990 (N_10990,N_3150,N_1841);
and U10991 (N_10991,N_5936,N_5560);
nor U10992 (N_10992,N_2334,N_1206);
nand U10993 (N_10993,N_4775,N_3850);
or U10994 (N_10994,N_2147,N_5152);
and U10995 (N_10995,N_4762,N_6076);
nand U10996 (N_10996,N_4505,N_6116);
nor U10997 (N_10997,N_1637,N_1741);
nand U10998 (N_10998,N_939,N_4524);
or U10999 (N_10999,N_5498,N_2843);
or U11000 (N_11000,N_603,N_4836);
or U11001 (N_11001,N_2881,N_3671);
nand U11002 (N_11002,N_1489,N_2775);
and U11003 (N_11003,N_3547,N_2498);
or U11004 (N_11004,N_6226,N_1441);
nand U11005 (N_11005,N_4834,N_1201);
or U11006 (N_11006,N_5963,N_5069);
nand U11007 (N_11007,N_2494,N_6059);
nor U11008 (N_11008,N_5797,N_2967);
nor U11009 (N_11009,N_4989,N_177);
or U11010 (N_11010,N_2369,N_1202);
nor U11011 (N_11011,N_935,N_1600);
or U11012 (N_11012,N_3180,N_1171);
nand U11013 (N_11013,N_4893,N_1362);
xor U11014 (N_11014,N_3343,N_2299);
xor U11015 (N_11015,N_1040,N_2661);
nand U11016 (N_11016,N_5286,N_2855);
nor U11017 (N_11017,N_1353,N_5694);
nor U11018 (N_11018,N_3071,N_3807);
nand U11019 (N_11019,N_2135,N_4254);
xnor U11020 (N_11020,N_3774,N_5317);
nor U11021 (N_11021,N_5412,N_1970);
xnor U11022 (N_11022,N_1184,N_3911);
nor U11023 (N_11023,N_3454,N_5274);
and U11024 (N_11024,N_852,N_1636);
nand U11025 (N_11025,N_1044,N_1420);
nor U11026 (N_11026,N_4084,N_68);
nand U11027 (N_11027,N_1490,N_5977);
and U11028 (N_11028,N_2204,N_608);
nand U11029 (N_11029,N_382,N_5178);
xnor U11030 (N_11030,N_2630,N_5115);
nor U11031 (N_11031,N_3181,N_2033);
nand U11032 (N_11032,N_5095,N_1357);
or U11033 (N_11033,N_3390,N_1128);
nor U11034 (N_11034,N_2204,N_5752);
or U11035 (N_11035,N_1059,N_5878);
or U11036 (N_11036,N_3667,N_5952);
nor U11037 (N_11037,N_296,N_1094);
and U11038 (N_11038,N_4204,N_6002);
nor U11039 (N_11039,N_4422,N_1766);
xor U11040 (N_11040,N_2191,N_3327);
or U11041 (N_11041,N_4011,N_379);
or U11042 (N_11042,N_2806,N_2451);
xnor U11043 (N_11043,N_1563,N_700);
xor U11044 (N_11044,N_2689,N_3942);
or U11045 (N_11045,N_4502,N_5204);
nor U11046 (N_11046,N_727,N_2962);
nor U11047 (N_11047,N_67,N_1916);
and U11048 (N_11048,N_4991,N_2392);
nor U11049 (N_11049,N_4140,N_280);
or U11050 (N_11050,N_2537,N_5317);
or U11051 (N_11051,N_12,N_4648);
or U11052 (N_11052,N_2608,N_4478);
nor U11053 (N_11053,N_388,N_4950);
or U11054 (N_11054,N_1001,N_5708);
nand U11055 (N_11055,N_23,N_67);
and U11056 (N_11056,N_4063,N_6127);
nand U11057 (N_11057,N_209,N_3475);
nand U11058 (N_11058,N_1957,N_3679);
or U11059 (N_11059,N_312,N_5594);
and U11060 (N_11060,N_1758,N_3923);
xnor U11061 (N_11061,N_3305,N_6247);
nor U11062 (N_11062,N_3120,N_1726);
and U11063 (N_11063,N_2934,N_2670);
or U11064 (N_11064,N_4298,N_338);
and U11065 (N_11065,N_1890,N_2719);
nor U11066 (N_11066,N_5623,N_4194);
or U11067 (N_11067,N_1428,N_373);
and U11068 (N_11068,N_2351,N_3061);
xor U11069 (N_11069,N_1177,N_3254);
nor U11070 (N_11070,N_2762,N_3113);
and U11071 (N_11071,N_1095,N_5028);
nand U11072 (N_11072,N_745,N_1690);
or U11073 (N_11073,N_3153,N_2820);
and U11074 (N_11074,N_3109,N_3979);
and U11075 (N_11075,N_487,N_988);
nand U11076 (N_11076,N_6173,N_3075);
nand U11077 (N_11077,N_2425,N_1965);
and U11078 (N_11078,N_2451,N_5663);
nor U11079 (N_11079,N_4422,N_2659);
xnor U11080 (N_11080,N_5687,N_5892);
nor U11081 (N_11081,N_3333,N_1808);
and U11082 (N_11082,N_1408,N_5763);
nor U11083 (N_11083,N_1659,N_2852);
nor U11084 (N_11084,N_3929,N_3604);
xnor U11085 (N_11085,N_6232,N_5684);
nor U11086 (N_11086,N_4940,N_568);
nand U11087 (N_11087,N_2099,N_3948);
nand U11088 (N_11088,N_2498,N_5736);
and U11089 (N_11089,N_1734,N_5158);
or U11090 (N_11090,N_2124,N_962);
nand U11091 (N_11091,N_5127,N_5050);
nor U11092 (N_11092,N_3812,N_4730);
and U11093 (N_11093,N_2105,N_1622);
nand U11094 (N_11094,N_4501,N_2723);
nor U11095 (N_11095,N_4281,N_343);
and U11096 (N_11096,N_2585,N_55);
xor U11097 (N_11097,N_4890,N_5155);
and U11098 (N_11098,N_212,N_2388);
nor U11099 (N_11099,N_2219,N_1873);
and U11100 (N_11100,N_2542,N_3399);
nor U11101 (N_11101,N_2542,N_5172);
nor U11102 (N_11102,N_4494,N_2293);
nor U11103 (N_11103,N_103,N_4653);
xnor U11104 (N_11104,N_1153,N_1674);
nand U11105 (N_11105,N_326,N_5099);
and U11106 (N_11106,N_1774,N_887);
nor U11107 (N_11107,N_4106,N_3766);
nor U11108 (N_11108,N_338,N_606);
and U11109 (N_11109,N_2061,N_4803);
and U11110 (N_11110,N_5701,N_4457);
nor U11111 (N_11111,N_5058,N_3316);
or U11112 (N_11112,N_1570,N_3569);
nand U11113 (N_11113,N_2900,N_872);
xor U11114 (N_11114,N_2473,N_2668);
nand U11115 (N_11115,N_6120,N_3349);
nand U11116 (N_11116,N_4545,N_1803);
nor U11117 (N_11117,N_5991,N_5370);
and U11118 (N_11118,N_1067,N_126);
or U11119 (N_11119,N_3295,N_1564);
and U11120 (N_11120,N_4953,N_1001);
nand U11121 (N_11121,N_4988,N_5802);
or U11122 (N_11122,N_1832,N_150);
or U11123 (N_11123,N_1010,N_4894);
or U11124 (N_11124,N_3851,N_3268);
nand U11125 (N_11125,N_1884,N_2785);
nor U11126 (N_11126,N_5164,N_2445);
or U11127 (N_11127,N_4159,N_3953);
xnor U11128 (N_11128,N_5437,N_4312);
xnor U11129 (N_11129,N_4367,N_4974);
nand U11130 (N_11130,N_3139,N_4942);
nor U11131 (N_11131,N_5634,N_2462);
and U11132 (N_11132,N_4441,N_486);
xnor U11133 (N_11133,N_3783,N_4660);
nor U11134 (N_11134,N_986,N_1042);
nand U11135 (N_11135,N_4461,N_1279);
and U11136 (N_11136,N_824,N_2305);
nand U11137 (N_11137,N_29,N_759);
xor U11138 (N_11138,N_3728,N_798);
nand U11139 (N_11139,N_3391,N_4414);
or U11140 (N_11140,N_3316,N_5531);
nor U11141 (N_11141,N_512,N_5174);
or U11142 (N_11142,N_761,N_2162);
or U11143 (N_11143,N_19,N_4273);
xor U11144 (N_11144,N_4991,N_6132);
xnor U11145 (N_11145,N_1412,N_4628);
or U11146 (N_11146,N_1956,N_2145);
and U11147 (N_11147,N_5384,N_2872);
nand U11148 (N_11148,N_2195,N_5398);
nor U11149 (N_11149,N_3230,N_634);
or U11150 (N_11150,N_455,N_2303);
nand U11151 (N_11151,N_3933,N_3370);
nor U11152 (N_11152,N_1726,N_2403);
nand U11153 (N_11153,N_1586,N_3509);
and U11154 (N_11154,N_756,N_2259);
or U11155 (N_11155,N_3960,N_6126);
nand U11156 (N_11156,N_4550,N_4614);
nand U11157 (N_11157,N_1907,N_4238);
or U11158 (N_11158,N_27,N_983);
nor U11159 (N_11159,N_436,N_4351);
nand U11160 (N_11160,N_4799,N_2232);
and U11161 (N_11161,N_5487,N_2577);
nor U11162 (N_11162,N_5511,N_3098);
and U11163 (N_11163,N_1029,N_4517);
nor U11164 (N_11164,N_5481,N_3199);
nor U11165 (N_11165,N_3461,N_377);
or U11166 (N_11166,N_175,N_1805);
or U11167 (N_11167,N_2518,N_1877);
or U11168 (N_11168,N_1865,N_5182);
or U11169 (N_11169,N_2560,N_4563);
xor U11170 (N_11170,N_5585,N_5960);
nor U11171 (N_11171,N_1259,N_6148);
or U11172 (N_11172,N_3684,N_768);
and U11173 (N_11173,N_4103,N_2883);
and U11174 (N_11174,N_86,N_139);
and U11175 (N_11175,N_3333,N_3778);
nor U11176 (N_11176,N_5425,N_5584);
or U11177 (N_11177,N_2421,N_3031);
nand U11178 (N_11178,N_1093,N_5782);
or U11179 (N_11179,N_2801,N_3676);
or U11180 (N_11180,N_3805,N_936);
and U11181 (N_11181,N_1209,N_2108);
nand U11182 (N_11182,N_3006,N_2975);
xor U11183 (N_11183,N_1504,N_4041);
xnor U11184 (N_11184,N_4737,N_588);
nor U11185 (N_11185,N_865,N_3711);
or U11186 (N_11186,N_525,N_4983);
and U11187 (N_11187,N_1263,N_1115);
or U11188 (N_11188,N_1682,N_3179);
and U11189 (N_11189,N_2743,N_4050);
nand U11190 (N_11190,N_5586,N_5424);
nor U11191 (N_11191,N_1581,N_6058);
nand U11192 (N_11192,N_4613,N_2916);
or U11193 (N_11193,N_1522,N_4899);
nand U11194 (N_11194,N_989,N_2457);
and U11195 (N_11195,N_901,N_5488);
nor U11196 (N_11196,N_3796,N_3644);
nor U11197 (N_11197,N_1614,N_3293);
nand U11198 (N_11198,N_5136,N_408);
or U11199 (N_11199,N_572,N_5009);
and U11200 (N_11200,N_4012,N_4671);
nand U11201 (N_11201,N_4356,N_365);
and U11202 (N_11202,N_3553,N_2423);
xor U11203 (N_11203,N_3942,N_5542);
nor U11204 (N_11204,N_439,N_2442);
nand U11205 (N_11205,N_1110,N_1891);
and U11206 (N_11206,N_771,N_1741);
nand U11207 (N_11207,N_1778,N_353);
nor U11208 (N_11208,N_2028,N_4816);
nor U11209 (N_11209,N_175,N_368);
or U11210 (N_11210,N_3323,N_745);
and U11211 (N_11211,N_5093,N_1170);
nor U11212 (N_11212,N_6177,N_1972);
or U11213 (N_11213,N_6197,N_5967);
nand U11214 (N_11214,N_5788,N_5390);
nor U11215 (N_11215,N_1788,N_1883);
and U11216 (N_11216,N_2751,N_3707);
nor U11217 (N_11217,N_6028,N_2862);
nand U11218 (N_11218,N_4548,N_3866);
xnor U11219 (N_11219,N_2558,N_6010);
and U11220 (N_11220,N_4170,N_4364);
nor U11221 (N_11221,N_6161,N_5247);
nand U11222 (N_11222,N_2850,N_2207);
nor U11223 (N_11223,N_5938,N_3614);
and U11224 (N_11224,N_720,N_2031);
or U11225 (N_11225,N_3219,N_4512);
or U11226 (N_11226,N_5555,N_3375);
nand U11227 (N_11227,N_5752,N_2393);
nor U11228 (N_11228,N_3134,N_301);
nand U11229 (N_11229,N_1606,N_5957);
xnor U11230 (N_11230,N_1750,N_3662);
and U11231 (N_11231,N_4955,N_645);
or U11232 (N_11232,N_5914,N_3992);
nor U11233 (N_11233,N_5285,N_4579);
or U11234 (N_11234,N_1973,N_4537);
or U11235 (N_11235,N_5543,N_4630);
xor U11236 (N_11236,N_2820,N_5356);
and U11237 (N_11237,N_1195,N_5119);
and U11238 (N_11238,N_3786,N_4583);
and U11239 (N_11239,N_4037,N_2486);
or U11240 (N_11240,N_1702,N_2532);
and U11241 (N_11241,N_3123,N_306);
nand U11242 (N_11242,N_2328,N_1213);
or U11243 (N_11243,N_4825,N_2896);
nor U11244 (N_11244,N_1266,N_5434);
and U11245 (N_11245,N_5559,N_2779);
nand U11246 (N_11246,N_4345,N_5289);
or U11247 (N_11247,N_532,N_1350);
and U11248 (N_11248,N_1309,N_3422);
or U11249 (N_11249,N_3476,N_519);
nand U11250 (N_11250,N_2726,N_2026);
or U11251 (N_11251,N_1574,N_2840);
nor U11252 (N_11252,N_5838,N_4442);
nand U11253 (N_11253,N_5968,N_1249);
nor U11254 (N_11254,N_4431,N_862);
and U11255 (N_11255,N_4408,N_4322);
nand U11256 (N_11256,N_884,N_2408);
nand U11257 (N_11257,N_1314,N_1021);
and U11258 (N_11258,N_4388,N_3002);
and U11259 (N_11259,N_205,N_3158);
and U11260 (N_11260,N_1333,N_5972);
or U11261 (N_11261,N_5200,N_2781);
nand U11262 (N_11262,N_3162,N_5236);
xnor U11263 (N_11263,N_222,N_4671);
and U11264 (N_11264,N_5014,N_6209);
or U11265 (N_11265,N_4734,N_4332);
nand U11266 (N_11266,N_5532,N_1791);
or U11267 (N_11267,N_6110,N_2606);
nor U11268 (N_11268,N_2430,N_3947);
nor U11269 (N_11269,N_578,N_1599);
nand U11270 (N_11270,N_1608,N_2686);
xnor U11271 (N_11271,N_1714,N_416);
or U11272 (N_11272,N_749,N_107);
nand U11273 (N_11273,N_2956,N_4535);
nand U11274 (N_11274,N_763,N_5921);
or U11275 (N_11275,N_1231,N_5609);
nor U11276 (N_11276,N_2003,N_4644);
and U11277 (N_11277,N_5622,N_2459);
nand U11278 (N_11278,N_775,N_212);
nor U11279 (N_11279,N_2850,N_3593);
nand U11280 (N_11280,N_2458,N_186);
or U11281 (N_11281,N_3691,N_1846);
or U11282 (N_11282,N_3486,N_6025);
xor U11283 (N_11283,N_1028,N_3465);
nor U11284 (N_11284,N_4930,N_3561);
nand U11285 (N_11285,N_4142,N_2562);
and U11286 (N_11286,N_2383,N_429);
nor U11287 (N_11287,N_4956,N_399);
or U11288 (N_11288,N_3319,N_3698);
xnor U11289 (N_11289,N_1954,N_3898);
nand U11290 (N_11290,N_5832,N_2434);
or U11291 (N_11291,N_1539,N_3140);
nor U11292 (N_11292,N_379,N_2156);
nor U11293 (N_11293,N_5581,N_1879);
or U11294 (N_11294,N_589,N_5991);
nor U11295 (N_11295,N_3174,N_470);
or U11296 (N_11296,N_2573,N_2578);
nand U11297 (N_11297,N_14,N_239);
nor U11298 (N_11298,N_2842,N_3739);
nor U11299 (N_11299,N_4127,N_5966);
xnor U11300 (N_11300,N_3375,N_3969);
nor U11301 (N_11301,N_256,N_3998);
nand U11302 (N_11302,N_3203,N_1522);
and U11303 (N_11303,N_632,N_3950);
and U11304 (N_11304,N_2729,N_4200);
nor U11305 (N_11305,N_2982,N_3444);
or U11306 (N_11306,N_1659,N_1960);
nor U11307 (N_11307,N_536,N_1753);
nand U11308 (N_11308,N_629,N_6215);
xor U11309 (N_11309,N_4727,N_6000);
nand U11310 (N_11310,N_332,N_5738);
nor U11311 (N_11311,N_2271,N_5055);
or U11312 (N_11312,N_3367,N_2235);
xnor U11313 (N_11313,N_5764,N_280);
or U11314 (N_11314,N_1879,N_972);
nor U11315 (N_11315,N_2769,N_288);
nor U11316 (N_11316,N_342,N_2271);
nand U11317 (N_11317,N_1890,N_40);
and U11318 (N_11318,N_959,N_3339);
nor U11319 (N_11319,N_622,N_4669);
and U11320 (N_11320,N_4418,N_854);
nand U11321 (N_11321,N_1837,N_824);
nor U11322 (N_11322,N_6240,N_4454);
and U11323 (N_11323,N_2787,N_3005);
xnor U11324 (N_11324,N_283,N_825);
nor U11325 (N_11325,N_721,N_4624);
nand U11326 (N_11326,N_1611,N_5343);
or U11327 (N_11327,N_3563,N_6188);
or U11328 (N_11328,N_3256,N_167);
nor U11329 (N_11329,N_1951,N_1279);
and U11330 (N_11330,N_2240,N_1589);
nor U11331 (N_11331,N_4779,N_3143);
xor U11332 (N_11332,N_1624,N_465);
or U11333 (N_11333,N_677,N_1226);
or U11334 (N_11334,N_4433,N_5135);
nand U11335 (N_11335,N_3690,N_5343);
xor U11336 (N_11336,N_6222,N_4594);
nand U11337 (N_11337,N_2334,N_857);
nor U11338 (N_11338,N_3151,N_4206);
and U11339 (N_11339,N_2310,N_5103);
nor U11340 (N_11340,N_1144,N_5010);
nand U11341 (N_11341,N_5527,N_1114);
or U11342 (N_11342,N_1264,N_5951);
and U11343 (N_11343,N_988,N_1290);
and U11344 (N_11344,N_2372,N_1780);
nor U11345 (N_11345,N_5684,N_978);
nand U11346 (N_11346,N_4541,N_5021);
nand U11347 (N_11347,N_1075,N_3492);
nor U11348 (N_11348,N_1195,N_5018);
or U11349 (N_11349,N_3204,N_1756);
nor U11350 (N_11350,N_2691,N_1802);
nor U11351 (N_11351,N_5550,N_4346);
and U11352 (N_11352,N_1097,N_134);
and U11353 (N_11353,N_2776,N_5284);
and U11354 (N_11354,N_5616,N_1757);
or U11355 (N_11355,N_3362,N_5934);
nor U11356 (N_11356,N_5290,N_4286);
or U11357 (N_11357,N_1584,N_846);
or U11358 (N_11358,N_3606,N_3430);
or U11359 (N_11359,N_182,N_1875);
nand U11360 (N_11360,N_1996,N_388);
nand U11361 (N_11361,N_6010,N_2582);
nand U11362 (N_11362,N_6018,N_3106);
and U11363 (N_11363,N_4845,N_4966);
and U11364 (N_11364,N_1715,N_1226);
nor U11365 (N_11365,N_3158,N_3296);
nand U11366 (N_11366,N_1,N_4599);
and U11367 (N_11367,N_2841,N_4091);
nand U11368 (N_11368,N_4930,N_2970);
nor U11369 (N_11369,N_4216,N_5352);
nand U11370 (N_11370,N_3312,N_5532);
nor U11371 (N_11371,N_2255,N_3343);
xor U11372 (N_11372,N_242,N_3006);
nor U11373 (N_11373,N_3490,N_4864);
and U11374 (N_11374,N_2045,N_6004);
or U11375 (N_11375,N_4008,N_5701);
nor U11376 (N_11376,N_1186,N_1101);
nor U11377 (N_11377,N_5486,N_1287);
xnor U11378 (N_11378,N_3003,N_1872);
nor U11379 (N_11379,N_414,N_5524);
nor U11380 (N_11380,N_2476,N_3020);
nand U11381 (N_11381,N_3957,N_2988);
and U11382 (N_11382,N_3082,N_3823);
and U11383 (N_11383,N_4201,N_3476);
nand U11384 (N_11384,N_42,N_299);
or U11385 (N_11385,N_1779,N_5747);
and U11386 (N_11386,N_5383,N_5219);
or U11387 (N_11387,N_3687,N_5336);
or U11388 (N_11388,N_3578,N_6094);
or U11389 (N_11389,N_3564,N_3013);
nor U11390 (N_11390,N_3744,N_790);
xor U11391 (N_11391,N_3856,N_4835);
or U11392 (N_11392,N_4544,N_3462);
or U11393 (N_11393,N_743,N_2247);
and U11394 (N_11394,N_3366,N_2349);
and U11395 (N_11395,N_428,N_5619);
or U11396 (N_11396,N_4628,N_5156);
or U11397 (N_11397,N_115,N_2150);
or U11398 (N_11398,N_769,N_27);
nor U11399 (N_11399,N_3034,N_3360);
or U11400 (N_11400,N_4382,N_6172);
or U11401 (N_11401,N_5472,N_199);
xnor U11402 (N_11402,N_3740,N_1319);
xnor U11403 (N_11403,N_2404,N_1452);
or U11404 (N_11404,N_1147,N_643);
or U11405 (N_11405,N_1760,N_1580);
nor U11406 (N_11406,N_4273,N_6126);
nand U11407 (N_11407,N_5712,N_128);
and U11408 (N_11408,N_150,N_5527);
and U11409 (N_11409,N_2180,N_1272);
or U11410 (N_11410,N_2043,N_460);
nor U11411 (N_11411,N_4969,N_2321);
nor U11412 (N_11412,N_2311,N_4761);
and U11413 (N_11413,N_3498,N_676);
nand U11414 (N_11414,N_4640,N_2059);
and U11415 (N_11415,N_195,N_3890);
or U11416 (N_11416,N_1409,N_5386);
and U11417 (N_11417,N_2895,N_151);
or U11418 (N_11418,N_5848,N_6099);
and U11419 (N_11419,N_2070,N_3273);
and U11420 (N_11420,N_1782,N_5384);
nand U11421 (N_11421,N_6021,N_3022);
nand U11422 (N_11422,N_1643,N_4615);
xor U11423 (N_11423,N_5016,N_5033);
nand U11424 (N_11424,N_2044,N_2487);
nand U11425 (N_11425,N_425,N_5929);
nor U11426 (N_11426,N_807,N_6197);
or U11427 (N_11427,N_1000,N_1839);
and U11428 (N_11428,N_2806,N_3050);
and U11429 (N_11429,N_2066,N_5503);
nand U11430 (N_11430,N_4583,N_4375);
nand U11431 (N_11431,N_292,N_1787);
nand U11432 (N_11432,N_132,N_75);
or U11433 (N_11433,N_5071,N_2962);
nand U11434 (N_11434,N_1088,N_3149);
and U11435 (N_11435,N_331,N_5053);
nand U11436 (N_11436,N_2595,N_5375);
nor U11437 (N_11437,N_3673,N_2897);
and U11438 (N_11438,N_4073,N_1209);
nand U11439 (N_11439,N_5545,N_368);
nand U11440 (N_11440,N_3435,N_3090);
nand U11441 (N_11441,N_3980,N_4477);
nor U11442 (N_11442,N_4618,N_4556);
xnor U11443 (N_11443,N_2655,N_2515);
nand U11444 (N_11444,N_1764,N_3322);
nand U11445 (N_11445,N_2847,N_1741);
and U11446 (N_11446,N_1284,N_2810);
xor U11447 (N_11447,N_2150,N_4080);
nand U11448 (N_11448,N_4560,N_579);
xnor U11449 (N_11449,N_4491,N_2766);
nor U11450 (N_11450,N_5344,N_5366);
nand U11451 (N_11451,N_5229,N_2797);
or U11452 (N_11452,N_3695,N_3018);
nand U11453 (N_11453,N_3141,N_2831);
xnor U11454 (N_11454,N_5151,N_3490);
or U11455 (N_11455,N_4471,N_836);
nor U11456 (N_11456,N_293,N_2898);
and U11457 (N_11457,N_4146,N_5061);
or U11458 (N_11458,N_1848,N_1739);
nor U11459 (N_11459,N_564,N_2766);
or U11460 (N_11460,N_2760,N_1321);
nor U11461 (N_11461,N_4424,N_4366);
nand U11462 (N_11462,N_3106,N_1093);
nor U11463 (N_11463,N_3741,N_1891);
nand U11464 (N_11464,N_5698,N_3250);
nor U11465 (N_11465,N_6157,N_1045);
nor U11466 (N_11466,N_1943,N_5056);
or U11467 (N_11467,N_2610,N_2185);
or U11468 (N_11468,N_2872,N_6245);
nor U11469 (N_11469,N_3402,N_5131);
nand U11470 (N_11470,N_4650,N_334);
and U11471 (N_11471,N_1071,N_2431);
xnor U11472 (N_11472,N_485,N_506);
nand U11473 (N_11473,N_4494,N_2997);
xor U11474 (N_11474,N_4652,N_3744);
nand U11475 (N_11475,N_6188,N_6042);
or U11476 (N_11476,N_4470,N_3467);
or U11477 (N_11477,N_1690,N_3552);
and U11478 (N_11478,N_5156,N_710);
and U11479 (N_11479,N_5264,N_4001);
nor U11480 (N_11480,N_3588,N_5756);
and U11481 (N_11481,N_1824,N_2289);
xor U11482 (N_11482,N_143,N_5187);
nand U11483 (N_11483,N_2569,N_439);
or U11484 (N_11484,N_2348,N_4211);
or U11485 (N_11485,N_6076,N_1202);
nor U11486 (N_11486,N_4469,N_4831);
or U11487 (N_11487,N_658,N_1581);
and U11488 (N_11488,N_4551,N_1853);
nand U11489 (N_11489,N_1014,N_4038);
or U11490 (N_11490,N_1906,N_1745);
nand U11491 (N_11491,N_2845,N_5014);
nand U11492 (N_11492,N_5541,N_2345);
xnor U11493 (N_11493,N_5134,N_1587);
or U11494 (N_11494,N_4055,N_2611);
nor U11495 (N_11495,N_2617,N_265);
nor U11496 (N_11496,N_854,N_1574);
nor U11497 (N_11497,N_3683,N_987);
and U11498 (N_11498,N_1493,N_76);
or U11499 (N_11499,N_5650,N_6085);
or U11500 (N_11500,N_1206,N_5280);
nor U11501 (N_11501,N_3397,N_3762);
nor U11502 (N_11502,N_656,N_3875);
or U11503 (N_11503,N_3609,N_316);
nor U11504 (N_11504,N_1715,N_2564);
nor U11505 (N_11505,N_3033,N_5681);
and U11506 (N_11506,N_2101,N_4366);
and U11507 (N_11507,N_2455,N_1835);
or U11508 (N_11508,N_4061,N_1918);
nor U11509 (N_11509,N_1155,N_4358);
or U11510 (N_11510,N_1632,N_1889);
xnor U11511 (N_11511,N_5509,N_297);
or U11512 (N_11512,N_2450,N_4702);
and U11513 (N_11513,N_3339,N_1525);
or U11514 (N_11514,N_1658,N_3261);
nand U11515 (N_11515,N_1942,N_5318);
nand U11516 (N_11516,N_4879,N_1716);
xor U11517 (N_11517,N_1040,N_3615);
or U11518 (N_11518,N_3410,N_3719);
nor U11519 (N_11519,N_2220,N_253);
or U11520 (N_11520,N_4811,N_4171);
or U11521 (N_11521,N_4703,N_2017);
nand U11522 (N_11522,N_3514,N_4348);
and U11523 (N_11523,N_5843,N_4192);
or U11524 (N_11524,N_3585,N_5771);
nor U11525 (N_11525,N_3479,N_2699);
nor U11526 (N_11526,N_3856,N_3178);
and U11527 (N_11527,N_5603,N_583);
and U11528 (N_11528,N_742,N_1091);
or U11529 (N_11529,N_3802,N_566);
nand U11530 (N_11530,N_4245,N_3871);
or U11531 (N_11531,N_5018,N_4250);
or U11532 (N_11532,N_4624,N_4182);
nor U11533 (N_11533,N_2083,N_480);
nand U11534 (N_11534,N_1783,N_5470);
nor U11535 (N_11535,N_815,N_1049);
or U11536 (N_11536,N_5542,N_4089);
or U11537 (N_11537,N_1321,N_4489);
nand U11538 (N_11538,N_2693,N_482);
xnor U11539 (N_11539,N_4409,N_4809);
and U11540 (N_11540,N_3764,N_4321);
nor U11541 (N_11541,N_5883,N_844);
nand U11542 (N_11542,N_4780,N_1178);
xor U11543 (N_11543,N_4500,N_3678);
nor U11544 (N_11544,N_2472,N_2163);
nor U11545 (N_11545,N_5735,N_1597);
nand U11546 (N_11546,N_3220,N_4338);
nor U11547 (N_11547,N_4696,N_4123);
nand U11548 (N_11548,N_3951,N_4028);
or U11549 (N_11549,N_1130,N_1453);
and U11550 (N_11550,N_3991,N_2908);
nand U11551 (N_11551,N_3695,N_1447);
nand U11552 (N_11552,N_5260,N_1075);
and U11553 (N_11553,N_3795,N_4608);
or U11554 (N_11554,N_5433,N_1128);
nand U11555 (N_11555,N_4003,N_3269);
or U11556 (N_11556,N_4421,N_603);
nand U11557 (N_11557,N_6152,N_3308);
nand U11558 (N_11558,N_5041,N_2719);
nand U11559 (N_11559,N_1193,N_2434);
and U11560 (N_11560,N_907,N_237);
nand U11561 (N_11561,N_4764,N_3138);
nand U11562 (N_11562,N_5139,N_2778);
nor U11563 (N_11563,N_1109,N_5155);
nand U11564 (N_11564,N_5345,N_5170);
and U11565 (N_11565,N_3069,N_1058);
and U11566 (N_11566,N_5943,N_6071);
and U11567 (N_11567,N_1240,N_5377);
nand U11568 (N_11568,N_3227,N_5577);
nor U11569 (N_11569,N_100,N_4337);
nor U11570 (N_11570,N_4086,N_3980);
nand U11571 (N_11571,N_5193,N_4965);
and U11572 (N_11572,N_5792,N_3320);
or U11573 (N_11573,N_3505,N_2262);
nor U11574 (N_11574,N_3390,N_1250);
nand U11575 (N_11575,N_1489,N_4721);
nor U11576 (N_11576,N_4453,N_2740);
nand U11577 (N_11577,N_4617,N_3121);
xor U11578 (N_11578,N_3606,N_1517);
xnor U11579 (N_11579,N_5789,N_2043);
nand U11580 (N_11580,N_275,N_4699);
nor U11581 (N_11581,N_5399,N_5662);
and U11582 (N_11582,N_4264,N_2568);
nor U11583 (N_11583,N_120,N_2953);
or U11584 (N_11584,N_2208,N_1341);
and U11585 (N_11585,N_2832,N_662);
or U11586 (N_11586,N_448,N_2794);
or U11587 (N_11587,N_3964,N_5940);
and U11588 (N_11588,N_66,N_381);
xnor U11589 (N_11589,N_2002,N_4657);
nand U11590 (N_11590,N_245,N_2884);
or U11591 (N_11591,N_2775,N_3826);
nor U11592 (N_11592,N_5185,N_3986);
nor U11593 (N_11593,N_4798,N_2116);
or U11594 (N_11594,N_3937,N_1169);
nand U11595 (N_11595,N_2849,N_4982);
or U11596 (N_11596,N_2575,N_4937);
or U11597 (N_11597,N_5017,N_183);
and U11598 (N_11598,N_5424,N_3738);
and U11599 (N_11599,N_3342,N_4278);
or U11600 (N_11600,N_3355,N_2724);
or U11601 (N_11601,N_416,N_4755);
nand U11602 (N_11602,N_6024,N_2546);
nand U11603 (N_11603,N_799,N_4635);
nor U11604 (N_11604,N_371,N_2243);
nand U11605 (N_11605,N_1129,N_3560);
and U11606 (N_11606,N_5685,N_1379);
or U11607 (N_11607,N_4247,N_4864);
or U11608 (N_11608,N_453,N_2565);
or U11609 (N_11609,N_3295,N_2776);
nor U11610 (N_11610,N_1447,N_5969);
and U11611 (N_11611,N_2568,N_5752);
nand U11612 (N_11612,N_5795,N_5017);
and U11613 (N_11613,N_746,N_1488);
nor U11614 (N_11614,N_3082,N_2639);
or U11615 (N_11615,N_4473,N_4563);
nor U11616 (N_11616,N_5015,N_2030);
xnor U11617 (N_11617,N_5407,N_3017);
nand U11618 (N_11618,N_4735,N_1333);
nand U11619 (N_11619,N_3380,N_4690);
and U11620 (N_11620,N_4800,N_627);
and U11621 (N_11621,N_1721,N_3464);
nand U11622 (N_11622,N_742,N_2841);
and U11623 (N_11623,N_1304,N_5448);
nor U11624 (N_11624,N_5662,N_3806);
xor U11625 (N_11625,N_997,N_1325);
and U11626 (N_11626,N_3486,N_3759);
or U11627 (N_11627,N_4713,N_5278);
xor U11628 (N_11628,N_3285,N_5412);
nor U11629 (N_11629,N_4743,N_6059);
xor U11630 (N_11630,N_5481,N_1099);
and U11631 (N_11631,N_1294,N_5977);
and U11632 (N_11632,N_2833,N_2738);
or U11633 (N_11633,N_2177,N_1165);
nor U11634 (N_11634,N_2310,N_2570);
xor U11635 (N_11635,N_2235,N_1058);
xnor U11636 (N_11636,N_1151,N_5536);
xor U11637 (N_11637,N_2711,N_2311);
and U11638 (N_11638,N_6029,N_1447);
or U11639 (N_11639,N_817,N_4268);
and U11640 (N_11640,N_5263,N_103);
nand U11641 (N_11641,N_2979,N_4633);
and U11642 (N_11642,N_175,N_5695);
or U11643 (N_11643,N_5288,N_1440);
or U11644 (N_11644,N_1526,N_1430);
xor U11645 (N_11645,N_2385,N_1348);
nand U11646 (N_11646,N_2474,N_6045);
and U11647 (N_11647,N_1827,N_64);
xnor U11648 (N_11648,N_4044,N_1538);
nor U11649 (N_11649,N_430,N_1518);
nor U11650 (N_11650,N_2375,N_4553);
or U11651 (N_11651,N_2245,N_3180);
and U11652 (N_11652,N_1566,N_5692);
and U11653 (N_11653,N_1723,N_4813);
and U11654 (N_11654,N_2066,N_2895);
xor U11655 (N_11655,N_5521,N_1638);
nor U11656 (N_11656,N_2800,N_4430);
nor U11657 (N_11657,N_1402,N_3072);
and U11658 (N_11658,N_5340,N_5694);
nor U11659 (N_11659,N_798,N_296);
or U11660 (N_11660,N_239,N_2333);
nor U11661 (N_11661,N_789,N_591);
xnor U11662 (N_11662,N_4761,N_4407);
or U11663 (N_11663,N_1109,N_5627);
and U11664 (N_11664,N_3046,N_468);
nand U11665 (N_11665,N_6156,N_4217);
or U11666 (N_11666,N_825,N_3736);
or U11667 (N_11667,N_2504,N_4860);
nand U11668 (N_11668,N_2803,N_3373);
or U11669 (N_11669,N_3905,N_4664);
and U11670 (N_11670,N_5557,N_394);
nor U11671 (N_11671,N_4712,N_523);
or U11672 (N_11672,N_4603,N_4360);
or U11673 (N_11673,N_3837,N_1648);
and U11674 (N_11674,N_5078,N_2621);
or U11675 (N_11675,N_2651,N_2927);
or U11676 (N_11676,N_3577,N_3681);
nor U11677 (N_11677,N_4432,N_2171);
or U11678 (N_11678,N_1127,N_2242);
nor U11679 (N_11679,N_3150,N_4735);
or U11680 (N_11680,N_4847,N_874);
or U11681 (N_11681,N_2971,N_251);
and U11682 (N_11682,N_1912,N_3326);
nor U11683 (N_11683,N_257,N_2983);
or U11684 (N_11684,N_2736,N_2542);
and U11685 (N_11685,N_4426,N_4151);
or U11686 (N_11686,N_803,N_3334);
or U11687 (N_11687,N_3626,N_1951);
or U11688 (N_11688,N_1153,N_2655);
nor U11689 (N_11689,N_645,N_466);
and U11690 (N_11690,N_3747,N_5440);
nor U11691 (N_11691,N_928,N_2669);
nand U11692 (N_11692,N_2245,N_5627);
xor U11693 (N_11693,N_287,N_1203);
or U11694 (N_11694,N_3045,N_5415);
nand U11695 (N_11695,N_1261,N_4794);
or U11696 (N_11696,N_1332,N_2124);
nor U11697 (N_11697,N_3525,N_3257);
or U11698 (N_11698,N_3482,N_4781);
xor U11699 (N_11699,N_1830,N_4062);
nor U11700 (N_11700,N_2840,N_2682);
nor U11701 (N_11701,N_1827,N_3744);
nand U11702 (N_11702,N_5563,N_3124);
nand U11703 (N_11703,N_5795,N_4274);
xnor U11704 (N_11704,N_6149,N_5028);
xor U11705 (N_11705,N_2982,N_837);
or U11706 (N_11706,N_4928,N_1711);
nor U11707 (N_11707,N_5937,N_6116);
nor U11708 (N_11708,N_4407,N_1816);
or U11709 (N_11709,N_1998,N_1433);
or U11710 (N_11710,N_3949,N_4977);
and U11711 (N_11711,N_3263,N_4524);
and U11712 (N_11712,N_3166,N_5130);
or U11713 (N_11713,N_899,N_1726);
or U11714 (N_11714,N_5892,N_4530);
or U11715 (N_11715,N_5159,N_1406);
xor U11716 (N_11716,N_5358,N_5459);
nor U11717 (N_11717,N_1879,N_3921);
nor U11718 (N_11718,N_926,N_1317);
nand U11719 (N_11719,N_4391,N_612);
and U11720 (N_11720,N_145,N_2913);
or U11721 (N_11721,N_5552,N_1754);
and U11722 (N_11722,N_8,N_367);
or U11723 (N_11723,N_1155,N_6022);
nand U11724 (N_11724,N_250,N_4864);
and U11725 (N_11725,N_2974,N_2589);
nand U11726 (N_11726,N_2312,N_4914);
nand U11727 (N_11727,N_5971,N_872);
and U11728 (N_11728,N_3412,N_3299);
or U11729 (N_11729,N_5924,N_6005);
nand U11730 (N_11730,N_1974,N_5848);
and U11731 (N_11731,N_5785,N_6066);
nor U11732 (N_11732,N_4834,N_3782);
and U11733 (N_11733,N_2538,N_5841);
and U11734 (N_11734,N_711,N_5395);
or U11735 (N_11735,N_3202,N_6046);
nand U11736 (N_11736,N_2485,N_920);
and U11737 (N_11737,N_3835,N_790);
nand U11738 (N_11738,N_4960,N_6139);
xor U11739 (N_11739,N_3046,N_350);
nor U11740 (N_11740,N_3301,N_2251);
and U11741 (N_11741,N_5837,N_3286);
nor U11742 (N_11742,N_2573,N_1133);
and U11743 (N_11743,N_1585,N_6198);
nor U11744 (N_11744,N_4443,N_491);
nand U11745 (N_11745,N_443,N_3309);
and U11746 (N_11746,N_1650,N_839);
or U11747 (N_11747,N_5290,N_3475);
nand U11748 (N_11748,N_6178,N_4352);
xnor U11749 (N_11749,N_3627,N_730);
nor U11750 (N_11750,N_3477,N_2986);
xnor U11751 (N_11751,N_3037,N_2453);
and U11752 (N_11752,N_2283,N_4271);
nor U11753 (N_11753,N_3535,N_722);
or U11754 (N_11754,N_2155,N_412);
nor U11755 (N_11755,N_4371,N_1745);
nor U11756 (N_11756,N_4969,N_2144);
or U11757 (N_11757,N_3903,N_4312);
nand U11758 (N_11758,N_1259,N_4752);
and U11759 (N_11759,N_4719,N_4644);
and U11760 (N_11760,N_4976,N_1362);
nor U11761 (N_11761,N_5504,N_2822);
nor U11762 (N_11762,N_1071,N_5985);
or U11763 (N_11763,N_1658,N_3883);
nor U11764 (N_11764,N_6240,N_1176);
or U11765 (N_11765,N_4509,N_269);
nor U11766 (N_11766,N_1610,N_6047);
nor U11767 (N_11767,N_2702,N_1261);
and U11768 (N_11768,N_1391,N_1350);
nor U11769 (N_11769,N_3153,N_1299);
nand U11770 (N_11770,N_3418,N_1244);
nor U11771 (N_11771,N_3227,N_1846);
nand U11772 (N_11772,N_2133,N_5411);
and U11773 (N_11773,N_5382,N_4352);
nor U11774 (N_11774,N_3125,N_5245);
or U11775 (N_11775,N_93,N_2574);
and U11776 (N_11776,N_1128,N_56);
and U11777 (N_11777,N_4803,N_5549);
nor U11778 (N_11778,N_6054,N_375);
nand U11779 (N_11779,N_5489,N_4643);
or U11780 (N_11780,N_1176,N_2759);
nand U11781 (N_11781,N_812,N_2247);
and U11782 (N_11782,N_3990,N_4590);
nand U11783 (N_11783,N_469,N_4881);
and U11784 (N_11784,N_5796,N_1649);
nand U11785 (N_11785,N_1760,N_5518);
and U11786 (N_11786,N_1273,N_4862);
nand U11787 (N_11787,N_588,N_1752);
nand U11788 (N_11788,N_3613,N_2029);
nor U11789 (N_11789,N_145,N_5223);
nor U11790 (N_11790,N_1951,N_4267);
or U11791 (N_11791,N_271,N_3771);
nor U11792 (N_11792,N_2037,N_4486);
nand U11793 (N_11793,N_6022,N_3062);
nand U11794 (N_11794,N_5582,N_1047);
or U11795 (N_11795,N_2693,N_4283);
nand U11796 (N_11796,N_1287,N_484);
or U11797 (N_11797,N_1096,N_967);
or U11798 (N_11798,N_1354,N_3945);
and U11799 (N_11799,N_3929,N_2829);
and U11800 (N_11800,N_465,N_2836);
nand U11801 (N_11801,N_4452,N_5591);
nor U11802 (N_11802,N_2106,N_1551);
and U11803 (N_11803,N_5604,N_1495);
nand U11804 (N_11804,N_1822,N_2685);
nand U11805 (N_11805,N_2336,N_6179);
or U11806 (N_11806,N_3183,N_122);
or U11807 (N_11807,N_6204,N_3766);
nor U11808 (N_11808,N_1811,N_5203);
xnor U11809 (N_11809,N_4545,N_3572);
or U11810 (N_11810,N_4852,N_2307);
and U11811 (N_11811,N_1573,N_677);
or U11812 (N_11812,N_212,N_533);
nand U11813 (N_11813,N_2954,N_406);
and U11814 (N_11814,N_1016,N_2871);
nand U11815 (N_11815,N_4823,N_750);
and U11816 (N_11816,N_2090,N_2546);
or U11817 (N_11817,N_4585,N_1175);
and U11818 (N_11818,N_2000,N_4052);
nand U11819 (N_11819,N_1931,N_2357);
or U11820 (N_11820,N_5968,N_2907);
nor U11821 (N_11821,N_3735,N_5878);
nor U11822 (N_11822,N_750,N_4167);
nand U11823 (N_11823,N_2343,N_416);
xor U11824 (N_11824,N_1649,N_2149);
xor U11825 (N_11825,N_2100,N_989);
nor U11826 (N_11826,N_1019,N_1778);
nand U11827 (N_11827,N_3263,N_3361);
or U11828 (N_11828,N_5924,N_864);
or U11829 (N_11829,N_4541,N_5152);
and U11830 (N_11830,N_438,N_2640);
nand U11831 (N_11831,N_5511,N_3489);
nand U11832 (N_11832,N_4470,N_316);
nor U11833 (N_11833,N_2547,N_5558);
and U11834 (N_11834,N_1603,N_1979);
and U11835 (N_11835,N_5191,N_855);
nand U11836 (N_11836,N_3448,N_4096);
and U11837 (N_11837,N_5267,N_5055);
xor U11838 (N_11838,N_645,N_1164);
or U11839 (N_11839,N_2713,N_1531);
or U11840 (N_11840,N_2380,N_3738);
or U11841 (N_11841,N_3105,N_4134);
nand U11842 (N_11842,N_1677,N_2551);
nor U11843 (N_11843,N_5183,N_495);
nand U11844 (N_11844,N_5115,N_361);
and U11845 (N_11845,N_2400,N_4535);
nand U11846 (N_11846,N_393,N_2027);
or U11847 (N_11847,N_830,N_5839);
nor U11848 (N_11848,N_4265,N_3744);
nand U11849 (N_11849,N_3789,N_4759);
nand U11850 (N_11850,N_5091,N_5048);
or U11851 (N_11851,N_1650,N_533);
or U11852 (N_11852,N_484,N_335);
nand U11853 (N_11853,N_2321,N_5143);
nor U11854 (N_11854,N_6081,N_804);
nor U11855 (N_11855,N_4365,N_4147);
or U11856 (N_11856,N_1974,N_3183);
and U11857 (N_11857,N_4437,N_949);
and U11858 (N_11858,N_1680,N_889);
and U11859 (N_11859,N_3268,N_5858);
nor U11860 (N_11860,N_1558,N_1695);
or U11861 (N_11861,N_3082,N_4565);
nor U11862 (N_11862,N_6220,N_4188);
nand U11863 (N_11863,N_198,N_3580);
nor U11864 (N_11864,N_4829,N_3814);
nor U11865 (N_11865,N_2217,N_5467);
nand U11866 (N_11866,N_1633,N_3685);
nand U11867 (N_11867,N_89,N_4532);
and U11868 (N_11868,N_2213,N_3531);
and U11869 (N_11869,N_3168,N_2906);
nand U11870 (N_11870,N_3518,N_2667);
nor U11871 (N_11871,N_1676,N_3736);
and U11872 (N_11872,N_5879,N_5099);
nand U11873 (N_11873,N_4086,N_3138);
nor U11874 (N_11874,N_1873,N_791);
nand U11875 (N_11875,N_1150,N_1184);
nand U11876 (N_11876,N_1407,N_2255);
nor U11877 (N_11877,N_2304,N_1537);
and U11878 (N_11878,N_5990,N_2688);
nand U11879 (N_11879,N_1719,N_225);
and U11880 (N_11880,N_6135,N_47);
and U11881 (N_11881,N_4356,N_5899);
or U11882 (N_11882,N_3815,N_6246);
and U11883 (N_11883,N_4977,N_3424);
and U11884 (N_11884,N_4601,N_3579);
nand U11885 (N_11885,N_264,N_5624);
nand U11886 (N_11886,N_207,N_3245);
or U11887 (N_11887,N_2525,N_695);
and U11888 (N_11888,N_1621,N_4034);
nor U11889 (N_11889,N_3213,N_3381);
and U11890 (N_11890,N_1074,N_2804);
nand U11891 (N_11891,N_963,N_4474);
and U11892 (N_11892,N_3202,N_3043);
or U11893 (N_11893,N_3667,N_4627);
nand U11894 (N_11894,N_1526,N_1594);
nor U11895 (N_11895,N_3132,N_1867);
and U11896 (N_11896,N_2362,N_4404);
and U11897 (N_11897,N_4271,N_3876);
and U11898 (N_11898,N_3814,N_5333);
and U11899 (N_11899,N_2304,N_380);
and U11900 (N_11900,N_1016,N_4624);
xnor U11901 (N_11901,N_3199,N_5857);
nor U11902 (N_11902,N_5781,N_635);
nor U11903 (N_11903,N_2701,N_3003);
nand U11904 (N_11904,N_788,N_4875);
and U11905 (N_11905,N_2478,N_525);
and U11906 (N_11906,N_3131,N_3975);
nor U11907 (N_11907,N_161,N_3731);
nor U11908 (N_11908,N_3458,N_5316);
nor U11909 (N_11909,N_5541,N_5671);
nor U11910 (N_11910,N_5330,N_5258);
xor U11911 (N_11911,N_5513,N_280);
nand U11912 (N_11912,N_228,N_2670);
nand U11913 (N_11913,N_4187,N_3082);
nor U11914 (N_11914,N_3697,N_2139);
nand U11915 (N_11915,N_4038,N_807);
nor U11916 (N_11916,N_4096,N_695);
nor U11917 (N_11917,N_191,N_2988);
nor U11918 (N_11918,N_2593,N_3759);
and U11919 (N_11919,N_4568,N_447);
or U11920 (N_11920,N_1507,N_3535);
and U11921 (N_11921,N_2109,N_4287);
and U11922 (N_11922,N_5311,N_4060);
or U11923 (N_11923,N_5797,N_1735);
nor U11924 (N_11924,N_1933,N_2854);
nand U11925 (N_11925,N_4805,N_2956);
nand U11926 (N_11926,N_514,N_81);
and U11927 (N_11927,N_3892,N_2296);
nor U11928 (N_11928,N_2418,N_5771);
nor U11929 (N_11929,N_1267,N_2059);
nor U11930 (N_11930,N_2317,N_4287);
or U11931 (N_11931,N_877,N_4734);
and U11932 (N_11932,N_2527,N_2833);
and U11933 (N_11933,N_6193,N_3078);
nor U11934 (N_11934,N_4378,N_6148);
and U11935 (N_11935,N_2876,N_419);
nor U11936 (N_11936,N_5649,N_5560);
or U11937 (N_11937,N_2937,N_5261);
nor U11938 (N_11938,N_645,N_3636);
or U11939 (N_11939,N_1106,N_1684);
nor U11940 (N_11940,N_2332,N_2199);
nor U11941 (N_11941,N_1017,N_1985);
nor U11942 (N_11942,N_5581,N_957);
nand U11943 (N_11943,N_5626,N_4348);
or U11944 (N_11944,N_570,N_4376);
nor U11945 (N_11945,N_5177,N_3238);
or U11946 (N_11946,N_3209,N_432);
nand U11947 (N_11947,N_5883,N_2449);
or U11948 (N_11948,N_865,N_1225);
nor U11949 (N_11949,N_1108,N_2187);
xor U11950 (N_11950,N_5065,N_5689);
or U11951 (N_11951,N_2955,N_5267);
and U11952 (N_11952,N_4553,N_3766);
and U11953 (N_11953,N_2824,N_3456);
nand U11954 (N_11954,N_5457,N_5033);
nor U11955 (N_11955,N_1269,N_4090);
and U11956 (N_11956,N_337,N_1027);
nand U11957 (N_11957,N_2876,N_1579);
nand U11958 (N_11958,N_4055,N_197);
nand U11959 (N_11959,N_5209,N_2235);
and U11960 (N_11960,N_2298,N_2986);
and U11961 (N_11961,N_2044,N_1297);
and U11962 (N_11962,N_4993,N_4407);
xnor U11963 (N_11963,N_3988,N_446);
and U11964 (N_11964,N_899,N_4160);
nor U11965 (N_11965,N_2553,N_6057);
and U11966 (N_11966,N_4247,N_330);
xor U11967 (N_11967,N_1084,N_84);
or U11968 (N_11968,N_1002,N_5767);
or U11969 (N_11969,N_855,N_842);
and U11970 (N_11970,N_5437,N_5251);
and U11971 (N_11971,N_164,N_1679);
and U11972 (N_11972,N_5901,N_2637);
nand U11973 (N_11973,N_97,N_5050);
or U11974 (N_11974,N_2131,N_5884);
nor U11975 (N_11975,N_6217,N_4189);
nor U11976 (N_11976,N_5250,N_4837);
xor U11977 (N_11977,N_4296,N_98);
nor U11978 (N_11978,N_3441,N_5802);
or U11979 (N_11979,N_1965,N_1946);
nor U11980 (N_11980,N_1135,N_3173);
or U11981 (N_11981,N_1247,N_35);
or U11982 (N_11982,N_3471,N_4510);
and U11983 (N_11983,N_3194,N_1414);
xor U11984 (N_11984,N_3494,N_994);
and U11985 (N_11985,N_4930,N_5595);
or U11986 (N_11986,N_4935,N_401);
nor U11987 (N_11987,N_3281,N_81);
nor U11988 (N_11988,N_5431,N_1296);
or U11989 (N_11989,N_722,N_1179);
nand U11990 (N_11990,N_2467,N_5736);
or U11991 (N_11991,N_1756,N_4111);
nand U11992 (N_11992,N_5997,N_5027);
nor U11993 (N_11993,N_5094,N_3178);
nor U11994 (N_11994,N_4382,N_2228);
nand U11995 (N_11995,N_3116,N_4103);
or U11996 (N_11996,N_3039,N_1924);
and U11997 (N_11997,N_136,N_285);
and U11998 (N_11998,N_5483,N_453);
or U11999 (N_11999,N_5250,N_5440);
nand U12000 (N_12000,N_3140,N_4972);
nand U12001 (N_12001,N_2830,N_3963);
and U12002 (N_12002,N_5780,N_3562);
or U12003 (N_12003,N_2370,N_171);
nand U12004 (N_12004,N_3116,N_3629);
xnor U12005 (N_12005,N_6129,N_3301);
or U12006 (N_12006,N_4526,N_5238);
and U12007 (N_12007,N_1326,N_4252);
nand U12008 (N_12008,N_877,N_1878);
or U12009 (N_12009,N_1982,N_565);
nor U12010 (N_12010,N_262,N_3403);
nand U12011 (N_12011,N_4179,N_4823);
nor U12012 (N_12012,N_3998,N_6003);
nand U12013 (N_12013,N_3151,N_2260);
xor U12014 (N_12014,N_4429,N_1431);
nor U12015 (N_12015,N_5917,N_4437);
xnor U12016 (N_12016,N_4420,N_582);
and U12017 (N_12017,N_205,N_2793);
xnor U12018 (N_12018,N_4570,N_823);
nor U12019 (N_12019,N_5831,N_5606);
or U12020 (N_12020,N_6228,N_1239);
nor U12021 (N_12021,N_3322,N_3140);
nor U12022 (N_12022,N_2496,N_5786);
and U12023 (N_12023,N_695,N_3799);
nor U12024 (N_12024,N_3406,N_1646);
and U12025 (N_12025,N_188,N_3399);
and U12026 (N_12026,N_4760,N_1656);
or U12027 (N_12027,N_5586,N_1983);
nand U12028 (N_12028,N_4889,N_1411);
or U12029 (N_12029,N_1527,N_1844);
or U12030 (N_12030,N_994,N_1463);
nand U12031 (N_12031,N_449,N_5114);
nor U12032 (N_12032,N_5216,N_229);
or U12033 (N_12033,N_4519,N_2684);
and U12034 (N_12034,N_3913,N_1011);
nor U12035 (N_12035,N_2006,N_1151);
nand U12036 (N_12036,N_949,N_575);
or U12037 (N_12037,N_2936,N_643);
and U12038 (N_12038,N_150,N_6219);
xor U12039 (N_12039,N_1505,N_711);
and U12040 (N_12040,N_4624,N_2684);
nand U12041 (N_12041,N_4259,N_1780);
xnor U12042 (N_12042,N_4119,N_1568);
or U12043 (N_12043,N_5836,N_4842);
or U12044 (N_12044,N_1833,N_4067);
or U12045 (N_12045,N_5898,N_2372);
nor U12046 (N_12046,N_1613,N_2739);
and U12047 (N_12047,N_3440,N_4497);
nand U12048 (N_12048,N_1257,N_1567);
and U12049 (N_12049,N_3527,N_6182);
or U12050 (N_12050,N_5235,N_1583);
xnor U12051 (N_12051,N_4915,N_3614);
or U12052 (N_12052,N_679,N_1462);
nand U12053 (N_12053,N_2524,N_46);
and U12054 (N_12054,N_6238,N_2595);
or U12055 (N_12055,N_1294,N_2578);
nand U12056 (N_12056,N_2173,N_4875);
and U12057 (N_12057,N_3879,N_1073);
or U12058 (N_12058,N_5462,N_305);
nor U12059 (N_12059,N_1597,N_5265);
xor U12060 (N_12060,N_5564,N_2830);
and U12061 (N_12061,N_4147,N_3159);
and U12062 (N_12062,N_5416,N_110);
or U12063 (N_12063,N_105,N_365);
nand U12064 (N_12064,N_4634,N_2788);
nor U12065 (N_12065,N_5280,N_3488);
nand U12066 (N_12066,N_607,N_5714);
nor U12067 (N_12067,N_5328,N_1363);
xnor U12068 (N_12068,N_5981,N_2852);
and U12069 (N_12069,N_336,N_886);
or U12070 (N_12070,N_2496,N_832);
nand U12071 (N_12071,N_477,N_54);
nor U12072 (N_12072,N_1920,N_5326);
and U12073 (N_12073,N_5619,N_5991);
and U12074 (N_12074,N_1981,N_2895);
xnor U12075 (N_12075,N_819,N_4293);
or U12076 (N_12076,N_1720,N_5176);
nor U12077 (N_12077,N_5810,N_2717);
xor U12078 (N_12078,N_2263,N_5453);
nor U12079 (N_12079,N_198,N_85);
or U12080 (N_12080,N_65,N_1520);
nand U12081 (N_12081,N_5127,N_4468);
nor U12082 (N_12082,N_6193,N_5050);
or U12083 (N_12083,N_2515,N_477);
or U12084 (N_12084,N_4593,N_863);
and U12085 (N_12085,N_2335,N_360);
nor U12086 (N_12086,N_2757,N_3242);
nand U12087 (N_12087,N_2003,N_6055);
and U12088 (N_12088,N_1095,N_4011);
and U12089 (N_12089,N_2563,N_2409);
nor U12090 (N_12090,N_3852,N_114);
nand U12091 (N_12091,N_5737,N_5832);
xnor U12092 (N_12092,N_2200,N_3634);
or U12093 (N_12093,N_2033,N_1941);
nor U12094 (N_12094,N_5028,N_3015);
nand U12095 (N_12095,N_3169,N_4612);
and U12096 (N_12096,N_2760,N_2662);
or U12097 (N_12097,N_4607,N_5091);
and U12098 (N_12098,N_5972,N_1906);
nand U12099 (N_12099,N_4398,N_4729);
and U12100 (N_12100,N_1494,N_1182);
nand U12101 (N_12101,N_2529,N_500);
nand U12102 (N_12102,N_2553,N_1678);
and U12103 (N_12103,N_1874,N_6107);
or U12104 (N_12104,N_5972,N_2869);
nand U12105 (N_12105,N_3177,N_2376);
and U12106 (N_12106,N_3914,N_990);
and U12107 (N_12107,N_4939,N_1902);
nor U12108 (N_12108,N_1843,N_3312);
or U12109 (N_12109,N_76,N_990);
nand U12110 (N_12110,N_617,N_3552);
nor U12111 (N_12111,N_4101,N_1513);
nand U12112 (N_12112,N_1701,N_3746);
xor U12113 (N_12113,N_1979,N_3513);
and U12114 (N_12114,N_2020,N_4811);
nand U12115 (N_12115,N_5567,N_802);
nor U12116 (N_12116,N_4908,N_2453);
xnor U12117 (N_12117,N_1066,N_3233);
xor U12118 (N_12118,N_4721,N_5648);
and U12119 (N_12119,N_5595,N_4796);
xor U12120 (N_12120,N_636,N_867);
or U12121 (N_12121,N_3530,N_118);
nor U12122 (N_12122,N_5071,N_960);
nand U12123 (N_12123,N_930,N_2803);
xnor U12124 (N_12124,N_804,N_4584);
xnor U12125 (N_12125,N_1016,N_3745);
nor U12126 (N_12126,N_5454,N_653);
nor U12127 (N_12127,N_5281,N_2321);
xor U12128 (N_12128,N_4190,N_5534);
nor U12129 (N_12129,N_1286,N_2844);
and U12130 (N_12130,N_1031,N_4812);
or U12131 (N_12131,N_3620,N_5495);
or U12132 (N_12132,N_5040,N_4715);
or U12133 (N_12133,N_6205,N_2081);
nand U12134 (N_12134,N_3575,N_670);
nand U12135 (N_12135,N_5089,N_2798);
nand U12136 (N_12136,N_1441,N_1947);
xnor U12137 (N_12137,N_3183,N_5666);
nand U12138 (N_12138,N_3487,N_2585);
nor U12139 (N_12139,N_2899,N_4284);
nand U12140 (N_12140,N_5696,N_3063);
nand U12141 (N_12141,N_3559,N_5341);
and U12142 (N_12142,N_2957,N_4136);
nand U12143 (N_12143,N_5630,N_5052);
and U12144 (N_12144,N_1580,N_576);
and U12145 (N_12145,N_1101,N_1694);
or U12146 (N_12146,N_1653,N_2458);
and U12147 (N_12147,N_6174,N_4506);
and U12148 (N_12148,N_2725,N_3851);
nand U12149 (N_12149,N_490,N_5509);
nor U12150 (N_12150,N_1862,N_449);
or U12151 (N_12151,N_3194,N_5880);
nor U12152 (N_12152,N_4858,N_4077);
nor U12153 (N_12153,N_5924,N_2886);
nor U12154 (N_12154,N_2613,N_4256);
nand U12155 (N_12155,N_339,N_5450);
nor U12156 (N_12156,N_523,N_5918);
or U12157 (N_12157,N_2146,N_6065);
and U12158 (N_12158,N_3609,N_2789);
nand U12159 (N_12159,N_5474,N_1812);
and U12160 (N_12160,N_3463,N_81);
nor U12161 (N_12161,N_3719,N_50);
or U12162 (N_12162,N_1366,N_269);
or U12163 (N_12163,N_831,N_2258);
or U12164 (N_12164,N_6050,N_3428);
and U12165 (N_12165,N_4260,N_5187);
nor U12166 (N_12166,N_3017,N_6098);
nor U12167 (N_12167,N_3118,N_4091);
nor U12168 (N_12168,N_3432,N_3757);
nor U12169 (N_12169,N_642,N_3900);
or U12170 (N_12170,N_5640,N_2868);
xor U12171 (N_12171,N_1474,N_5420);
or U12172 (N_12172,N_1727,N_4803);
and U12173 (N_12173,N_3228,N_2576);
nand U12174 (N_12174,N_3276,N_4203);
nand U12175 (N_12175,N_4075,N_4982);
nor U12176 (N_12176,N_2048,N_4513);
nand U12177 (N_12177,N_5240,N_313);
nor U12178 (N_12178,N_1472,N_4070);
nand U12179 (N_12179,N_2983,N_44);
and U12180 (N_12180,N_2018,N_4585);
or U12181 (N_12181,N_5055,N_5476);
nor U12182 (N_12182,N_1110,N_5350);
nand U12183 (N_12183,N_3959,N_4163);
or U12184 (N_12184,N_712,N_1442);
nor U12185 (N_12185,N_866,N_5470);
and U12186 (N_12186,N_5296,N_5589);
nor U12187 (N_12187,N_20,N_3237);
xnor U12188 (N_12188,N_4565,N_1585);
nor U12189 (N_12189,N_1237,N_3161);
nand U12190 (N_12190,N_1389,N_637);
and U12191 (N_12191,N_6104,N_208);
or U12192 (N_12192,N_4748,N_1092);
xnor U12193 (N_12193,N_794,N_1752);
xor U12194 (N_12194,N_1924,N_903);
nand U12195 (N_12195,N_2374,N_588);
nand U12196 (N_12196,N_3265,N_4268);
nand U12197 (N_12197,N_1801,N_548);
or U12198 (N_12198,N_3742,N_2451);
nor U12199 (N_12199,N_1782,N_1616);
or U12200 (N_12200,N_2972,N_3977);
nand U12201 (N_12201,N_1059,N_1526);
nand U12202 (N_12202,N_2349,N_4127);
nor U12203 (N_12203,N_3250,N_5272);
nor U12204 (N_12204,N_622,N_2612);
and U12205 (N_12205,N_3699,N_3345);
nand U12206 (N_12206,N_1868,N_4420);
and U12207 (N_12207,N_4935,N_5871);
and U12208 (N_12208,N_2279,N_77);
nor U12209 (N_12209,N_3191,N_472);
nand U12210 (N_12210,N_3619,N_3090);
nor U12211 (N_12211,N_206,N_983);
or U12212 (N_12212,N_108,N_37);
nand U12213 (N_12213,N_2738,N_3485);
nand U12214 (N_12214,N_4159,N_3146);
or U12215 (N_12215,N_4399,N_3513);
and U12216 (N_12216,N_3534,N_648);
and U12217 (N_12217,N_4061,N_4727);
and U12218 (N_12218,N_3445,N_3684);
nor U12219 (N_12219,N_953,N_551);
or U12220 (N_12220,N_573,N_3481);
xor U12221 (N_12221,N_4392,N_987);
nand U12222 (N_12222,N_5588,N_4295);
or U12223 (N_12223,N_5708,N_241);
and U12224 (N_12224,N_3304,N_2712);
nor U12225 (N_12225,N_5549,N_2233);
or U12226 (N_12226,N_4883,N_3236);
nand U12227 (N_12227,N_3721,N_2504);
or U12228 (N_12228,N_284,N_5822);
nand U12229 (N_12229,N_1959,N_2169);
or U12230 (N_12230,N_662,N_3299);
or U12231 (N_12231,N_5596,N_5375);
nor U12232 (N_12232,N_5235,N_1141);
nand U12233 (N_12233,N_4624,N_2833);
nor U12234 (N_12234,N_90,N_4246);
xor U12235 (N_12235,N_1708,N_4084);
nand U12236 (N_12236,N_3435,N_4534);
and U12237 (N_12237,N_2288,N_3172);
nor U12238 (N_12238,N_1005,N_1862);
nand U12239 (N_12239,N_1855,N_6127);
or U12240 (N_12240,N_1775,N_5641);
or U12241 (N_12241,N_1221,N_4930);
and U12242 (N_12242,N_5783,N_2709);
nand U12243 (N_12243,N_5934,N_2554);
and U12244 (N_12244,N_1585,N_4205);
and U12245 (N_12245,N_1718,N_1641);
and U12246 (N_12246,N_4409,N_5179);
and U12247 (N_12247,N_609,N_5706);
and U12248 (N_12248,N_3833,N_5204);
or U12249 (N_12249,N_2121,N_1926);
nor U12250 (N_12250,N_1855,N_1693);
nand U12251 (N_12251,N_556,N_1344);
and U12252 (N_12252,N_3048,N_5657);
and U12253 (N_12253,N_5455,N_411);
and U12254 (N_12254,N_4308,N_3799);
or U12255 (N_12255,N_1927,N_4874);
or U12256 (N_12256,N_3260,N_2149);
and U12257 (N_12257,N_2546,N_4302);
xor U12258 (N_12258,N_280,N_3541);
and U12259 (N_12259,N_1478,N_5655);
nand U12260 (N_12260,N_5720,N_4426);
xnor U12261 (N_12261,N_1156,N_3446);
nor U12262 (N_12262,N_1427,N_4222);
or U12263 (N_12263,N_1713,N_1113);
and U12264 (N_12264,N_997,N_2433);
nor U12265 (N_12265,N_2745,N_3481);
nand U12266 (N_12266,N_3405,N_2778);
or U12267 (N_12267,N_732,N_3404);
nor U12268 (N_12268,N_2656,N_1582);
nand U12269 (N_12269,N_443,N_3845);
and U12270 (N_12270,N_2001,N_2021);
nor U12271 (N_12271,N_1119,N_582);
or U12272 (N_12272,N_1501,N_4533);
and U12273 (N_12273,N_6229,N_1791);
and U12274 (N_12274,N_2915,N_1039);
xnor U12275 (N_12275,N_1376,N_799);
nor U12276 (N_12276,N_4410,N_266);
nor U12277 (N_12277,N_1015,N_3677);
and U12278 (N_12278,N_1652,N_4574);
nand U12279 (N_12279,N_1588,N_5492);
xnor U12280 (N_12280,N_3898,N_3178);
and U12281 (N_12281,N_2959,N_5262);
nor U12282 (N_12282,N_899,N_5035);
nor U12283 (N_12283,N_5353,N_314);
nand U12284 (N_12284,N_2845,N_3563);
or U12285 (N_12285,N_5980,N_6129);
nor U12286 (N_12286,N_3138,N_479);
or U12287 (N_12287,N_461,N_4488);
nor U12288 (N_12288,N_157,N_1748);
or U12289 (N_12289,N_3362,N_2536);
and U12290 (N_12290,N_5330,N_5909);
nor U12291 (N_12291,N_774,N_547);
nor U12292 (N_12292,N_3300,N_4123);
nor U12293 (N_12293,N_5651,N_4849);
nand U12294 (N_12294,N_6062,N_756);
and U12295 (N_12295,N_83,N_4462);
xor U12296 (N_12296,N_907,N_4559);
nor U12297 (N_12297,N_2857,N_3304);
and U12298 (N_12298,N_3892,N_4959);
nor U12299 (N_12299,N_6174,N_2162);
or U12300 (N_12300,N_4394,N_3449);
nor U12301 (N_12301,N_3085,N_4976);
xor U12302 (N_12302,N_4030,N_348);
or U12303 (N_12303,N_2111,N_246);
or U12304 (N_12304,N_3149,N_3578);
and U12305 (N_12305,N_5519,N_1833);
or U12306 (N_12306,N_4877,N_3745);
and U12307 (N_12307,N_5230,N_3455);
nand U12308 (N_12308,N_415,N_4044);
and U12309 (N_12309,N_5428,N_723);
and U12310 (N_12310,N_3508,N_5014);
nor U12311 (N_12311,N_281,N_1153);
nor U12312 (N_12312,N_2436,N_2356);
or U12313 (N_12313,N_5706,N_1090);
or U12314 (N_12314,N_5160,N_6148);
nand U12315 (N_12315,N_3245,N_4009);
xor U12316 (N_12316,N_1963,N_5999);
and U12317 (N_12317,N_1653,N_804);
or U12318 (N_12318,N_555,N_5147);
and U12319 (N_12319,N_4576,N_2718);
and U12320 (N_12320,N_1805,N_2341);
and U12321 (N_12321,N_705,N_4192);
or U12322 (N_12322,N_5569,N_4880);
or U12323 (N_12323,N_850,N_2941);
xor U12324 (N_12324,N_1370,N_424);
or U12325 (N_12325,N_1961,N_1027);
or U12326 (N_12326,N_3927,N_127);
and U12327 (N_12327,N_5877,N_2367);
nand U12328 (N_12328,N_2506,N_3367);
xnor U12329 (N_12329,N_2334,N_1643);
nor U12330 (N_12330,N_2545,N_630);
and U12331 (N_12331,N_3640,N_701);
and U12332 (N_12332,N_2686,N_2348);
xor U12333 (N_12333,N_869,N_2924);
xor U12334 (N_12334,N_6011,N_3108);
and U12335 (N_12335,N_4039,N_879);
nand U12336 (N_12336,N_162,N_4398);
nand U12337 (N_12337,N_1301,N_2391);
nor U12338 (N_12338,N_4413,N_5099);
nand U12339 (N_12339,N_5052,N_6205);
nand U12340 (N_12340,N_5535,N_1359);
nor U12341 (N_12341,N_3098,N_2970);
xor U12342 (N_12342,N_66,N_1135);
nor U12343 (N_12343,N_1811,N_3185);
nand U12344 (N_12344,N_800,N_897);
and U12345 (N_12345,N_2663,N_2555);
xor U12346 (N_12346,N_903,N_2615);
nand U12347 (N_12347,N_1920,N_5696);
or U12348 (N_12348,N_384,N_3564);
nor U12349 (N_12349,N_749,N_5100);
and U12350 (N_12350,N_1908,N_954);
or U12351 (N_12351,N_4571,N_3085);
nor U12352 (N_12352,N_2598,N_1611);
or U12353 (N_12353,N_4068,N_376);
xnor U12354 (N_12354,N_3664,N_2634);
nor U12355 (N_12355,N_2712,N_2808);
nand U12356 (N_12356,N_1447,N_6205);
or U12357 (N_12357,N_5001,N_1119);
nor U12358 (N_12358,N_1612,N_5628);
and U12359 (N_12359,N_3961,N_1146);
or U12360 (N_12360,N_3278,N_3490);
xnor U12361 (N_12361,N_2003,N_4932);
and U12362 (N_12362,N_3056,N_4346);
or U12363 (N_12363,N_1631,N_1153);
xor U12364 (N_12364,N_2830,N_2613);
nand U12365 (N_12365,N_2187,N_3125);
and U12366 (N_12366,N_3977,N_6245);
or U12367 (N_12367,N_461,N_1568);
nand U12368 (N_12368,N_4117,N_2380);
nand U12369 (N_12369,N_5223,N_1209);
nand U12370 (N_12370,N_2548,N_434);
or U12371 (N_12371,N_527,N_1012);
nand U12372 (N_12372,N_5478,N_891);
nand U12373 (N_12373,N_4619,N_4885);
nor U12374 (N_12374,N_3195,N_1000);
and U12375 (N_12375,N_5184,N_3268);
nor U12376 (N_12376,N_5035,N_3616);
xor U12377 (N_12377,N_5043,N_5999);
nand U12378 (N_12378,N_2806,N_832);
and U12379 (N_12379,N_4175,N_1760);
nor U12380 (N_12380,N_544,N_587);
or U12381 (N_12381,N_2378,N_707);
and U12382 (N_12382,N_5531,N_4386);
or U12383 (N_12383,N_6033,N_866);
and U12384 (N_12384,N_1600,N_3753);
and U12385 (N_12385,N_1267,N_4070);
and U12386 (N_12386,N_43,N_1913);
or U12387 (N_12387,N_2027,N_2417);
or U12388 (N_12388,N_1117,N_2511);
and U12389 (N_12389,N_3791,N_1734);
nand U12390 (N_12390,N_4630,N_4103);
nand U12391 (N_12391,N_1261,N_1130);
and U12392 (N_12392,N_3028,N_2877);
nand U12393 (N_12393,N_5475,N_1004);
nor U12394 (N_12394,N_1787,N_4301);
nand U12395 (N_12395,N_1381,N_2860);
xnor U12396 (N_12396,N_1467,N_3710);
or U12397 (N_12397,N_1200,N_798);
nor U12398 (N_12398,N_1744,N_5183);
or U12399 (N_12399,N_4796,N_345);
or U12400 (N_12400,N_5636,N_3954);
or U12401 (N_12401,N_4924,N_1120);
or U12402 (N_12402,N_2095,N_2020);
nor U12403 (N_12403,N_3095,N_4619);
nor U12404 (N_12404,N_5970,N_987);
nand U12405 (N_12405,N_661,N_8);
and U12406 (N_12406,N_2220,N_1798);
nand U12407 (N_12407,N_2879,N_787);
nand U12408 (N_12408,N_5162,N_4651);
or U12409 (N_12409,N_346,N_4163);
and U12410 (N_12410,N_5028,N_4445);
nor U12411 (N_12411,N_5501,N_1570);
or U12412 (N_12412,N_2408,N_4005);
nand U12413 (N_12413,N_4116,N_1817);
and U12414 (N_12414,N_4221,N_3944);
nand U12415 (N_12415,N_4861,N_3838);
nor U12416 (N_12416,N_2715,N_689);
xor U12417 (N_12417,N_4916,N_3140);
nand U12418 (N_12418,N_2109,N_3864);
nand U12419 (N_12419,N_200,N_2262);
and U12420 (N_12420,N_586,N_4142);
nor U12421 (N_12421,N_4815,N_1949);
nand U12422 (N_12422,N_3556,N_2007);
and U12423 (N_12423,N_807,N_5656);
or U12424 (N_12424,N_3817,N_847);
xor U12425 (N_12425,N_4011,N_2817);
and U12426 (N_12426,N_5290,N_3954);
and U12427 (N_12427,N_58,N_5684);
xor U12428 (N_12428,N_69,N_3644);
nor U12429 (N_12429,N_4178,N_2688);
and U12430 (N_12430,N_1524,N_3124);
or U12431 (N_12431,N_2644,N_4006);
and U12432 (N_12432,N_3048,N_3282);
and U12433 (N_12433,N_535,N_590);
nor U12434 (N_12434,N_3491,N_2656);
nand U12435 (N_12435,N_578,N_3355);
nand U12436 (N_12436,N_2153,N_5005);
or U12437 (N_12437,N_10,N_5122);
nand U12438 (N_12438,N_37,N_2547);
nor U12439 (N_12439,N_2212,N_5550);
nand U12440 (N_12440,N_1756,N_1800);
nor U12441 (N_12441,N_1053,N_4650);
and U12442 (N_12442,N_5929,N_179);
xor U12443 (N_12443,N_149,N_5141);
and U12444 (N_12444,N_415,N_1547);
nor U12445 (N_12445,N_5405,N_2086);
and U12446 (N_12446,N_4221,N_2299);
nor U12447 (N_12447,N_1809,N_3452);
nand U12448 (N_12448,N_4884,N_434);
nor U12449 (N_12449,N_6216,N_4900);
or U12450 (N_12450,N_2971,N_375);
nand U12451 (N_12451,N_2911,N_5667);
nor U12452 (N_12452,N_5632,N_3550);
nor U12453 (N_12453,N_2223,N_1915);
nor U12454 (N_12454,N_186,N_2992);
nor U12455 (N_12455,N_5503,N_5559);
or U12456 (N_12456,N_5296,N_5624);
nor U12457 (N_12457,N_3712,N_749);
nor U12458 (N_12458,N_4094,N_5174);
or U12459 (N_12459,N_2181,N_1853);
nor U12460 (N_12460,N_13,N_613);
nor U12461 (N_12461,N_2734,N_1645);
or U12462 (N_12462,N_3343,N_2082);
nor U12463 (N_12463,N_1393,N_1751);
xnor U12464 (N_12464,N_665,N_3295);
nor U12465 (N_12465,N_4817,N_5733);
nand U12466 (N_12466,N_2976,N_5209);
nand U12467 (N_12467,N_3988,N_353);
nand U12468 (N_12468,N_3892,N_5211);
nor U12469 (N_12469,N_1625,N_5457);
xnor U12470 (N_12470,N_248,N_4665);
nor U12471 (N_12471,N_6133,N_4303);
or U12472 (N_12472,N_6068,N_4148);
or U12473 (N_12473,N_1237,N_5846);
and U12474 (N_12474,N_1886,N_5734);
or U12475 (N_12475,N_1286,N_3169);
or U12476 (N_12476,N_3677,N_3904);
xor U12477 (N_12477,N_2693,N_720);
xor U12478 (N_12478,N_2157,N_2405);
nor U12479 (N_12479,N_3027,N_4189);
nand U12480 (N_12480,N_3231,N_722);
and U12481 (N_12481,N_2708,N_5237);
nor U12482 (N_12482,N_2740,N_1099);
and U12483 (N_12483,N_4283,N_4802);
nand U12484 (N_12484,N_314,N_4703);
xor U12485 (N_12485,N_2649,N_1753);
or U12486 (N_12486,N_5730,N_981);
xnor U12487 (N_12487,N_1111,N_3316);
nor U12488 (N_12488,N_1063,N_5921);
or U12489 (N_12489,N_1726,N_5417);
nand U12490 (N_12490,N_6111,N_3079);
and U12491 (N_12491,N_4359,N_850);
nor U12492 (N_12492,N_349,N_1598);
xnor U12493 (N_12493,N_3549,N_157);
nor U12494 (N_12494,N_3871,N_4914);
xnor U12495 (N_12495,N_388,N_5556);
and U12496 (N_12496,N_4165,N_3011);
nor U12497 (N_12497,N_131,N_4192);
xnor U12498 (N_12498,N_4242,N_2824);
nand U12499 (N_12499,N_2456,N_3117);
or U12500 (N_12500,N_8945,N_9658);
nor U12501 (N_12501,N_7332,N_11847);
xor U12502 (N_12502,N_8893,N_11233);
xnor U12503 (N_12503,N_12426,N_7546);
nor U12504 (N_12504,N_7676,N_11451);
and U12505 (N_12505,N_8823,N_11510);
nand U12506 (N_12506,N_8814,N_12291);
xor U12507 (N_12507,N_6537,N_12054);
nor U12508 (N_12508,N_12049,N_10494);
nand U12509 (N_12509,N_8970,N_12168);
and U12510 (N_12510,N_12047,N_11732);
xor U12511 (N_12511,N_11357,N_7955);
nor U12512 (N_12512,N_10215,N_11134);
or U12513 (N_12513,N_12343,N_8175);
and U12514 (N_12514,N_9030,N_7279);
xnor U12515 (N_12515,N_11093,N_10464);
and U12516 (N_12516,N_11334,N_11707);
or U12517 (N_12517,N_7277,N_9197);
xor U12518 (N_12518,N_9927,N_8515);
and U12519 (N_12519,N_10459,N_12040);
nand U12520 (N_12520,N_12165,N_7403);
or U12521 (N_12521,N_12278,N_12466);
and U12522 (N_12522,N_8055,N_11658);
and U12523 (N_12523,N_12449,N_8256);
or U12524 (N_12524,N_11508,N_11650);
nor U12525 (N_12525,N_8588,N_6747);
xnor U12526 (N_12526,N_10070,N_8167);
and U12527 (N_12527,N_6990,N_10090);
nor U12528 (N_12528,N_10607,N_8231);
nor U12529 (N_12529,N_8702,N_8137);
or U12530 (N_12530,N_8200,N_7871);
and U12531 (N_12531,N_7750,N_8343);
or U12532 (N_12532,N_10791,N_10989);
nor U12533 (N_12533,N_7926,N_9179);
and U12534 (N_12534,N_6810,N_8813);
or U12535 (N_12535,N_11395,N_10782);
xor U12536 (N_12536,N_11033,N_9499);
nor U12537 (N_12537,N_9611,N_9328);
or U12538 (N_12538,N_11772,N_8599);
and U12539 (N_12539,N_7350,N_11612);
or U12540 (N_12540,N_8082,N_11073);
or U12541 (N_12541,N_8145,N_12155);
nand U12542 (N_12542,N_8380,N_7213);
nor U12543 (N_12543,N_6974,N_11378);
nand U12544 (N_12544,N_9272,N_7587);
and U12545 (N_12545,N_8552,N_7706);
xnor U12546 (N_12546,N_11686,N_9845);
and U12547 (N_12547,N_11742,N_8192);
or U12548 (N_12548,N_6888,N_11095);
nor U12549 (N_12549,N_12363,N_8210);
or U12550 (N_12550,N_9726,N_9990);
nand U12551 (N_12551,N_9831,N_11494);
or U12552 (N_12552,N_8844,N_11101);
xor U12553 (N_12553,N_8418,N_8456);
nor U12554 (N_12554,N_11930,N_6658);
and U12555 (N_12555,N_7549,N_12354);
nor U12556 (N_12556,N_9915,N_8749);
and U12557 (N_12557,N_6822,N_12117);
and U12558 (N_12558,N_9731,N_9476);
and U12559 (N_12559,N_7057,N_8060);
nor U12560 (N_12560,N_12485,N_11043);
nand U12561 (N_12561,N_10477,N_12166);
xnor U12562 (N_12562,N_8903,N_10422);
nor U12563 (N_12563,N_12212,N_6564);
or U12564 (N_12564,N_6913,N_7615);
nor U12565 (N_12565,N_8387,N_6620);
and U12566 (N_12566,N_9366,N_10149);
nor U12567 (N_12567,N_8463,N_6274);
and U12568 (N_12568,N_10969,N_9623);
or U12569 (N_12569,N_12479,N_10768);
and U12570 (N_12570,N_8233,N_10577);
or U12571 (N_12571,N_11800,N_10666);
and U12572 (N_12572,N_7911,N_12398);
or U12573 (N_12573,N_7198,N_8936);
nand U12574 (N_12574,N_11063,N_8288);
or U12575 (N_12575,N_9784,N_7247);
and U12576 (N_12576,N_10073,N_11420);
nand U12577 (N_12577,N_7319,N_9717);
nand U12578 (N_12578,N_10805,N_6409);
or U12579 (N_12579,N_11836,N_10342);
nand U12580 (N_12580,N_8521,N_12308);
nand U12581 (N_12581,N_12246,N_8650);
and U12582 (N_12582,N_11399,N_8294);
nand U12583 (N_12583,N_9562,N_8101);
nor U12584 (N_12584,N_7987,N_7008);
nor U12585 (N_12585,N_10853,N_11606);
xor U12586 (N_12586,N_10628,N_12233);
or U12587 (N_12587,N_6824,N_8785);
xor U12588 (N_12588,N_11358,N_10418);
and U12589 (N_12589,N_7890,N_9419);
nand U12590 (N_12590,N_10462,N_11400);
nor U12591 (N_12591,N_11105,N_8701);
xor U12592 (N_12592,N_7148,N_12069);
nor U12593 (N_12593,N_10059,N_8014);
and U12594 (N_12594,N_7295,N_10207);
nand U12595 (N_12595,N_10637,N_8853);
nor U12596 (N_12596,N_11630,N_6811);
and U12597 (N_12597,N_10926,N_8135);
xnor U12598 (N_12598,N_7133,N_8609);
xnor U12599 (N_12599,N_11901,N_10844);
nand U12600 (N_12600,N_8394,N_8216);
xnor U12601 (N_12601,N_10951,N_9357);
or U12602 (N_12602,N_9038,N_10045);
nand U12603 (N_12603,N_7648,N_8023);
nor U12604 (N_12604,N_9232,N_7651);
or U12605 (N_12605,N_10238,N_12038);
nand U12606 (N_12606,N_7820,N_9669);
nand U12607 (N_12607,N_8349,N_6687);
nor U12608 (N_12608,N_6730,N_6353);
nor U12609 (N_12609,N_12442,N_10243);
or U12610 (N_12610,N_8781,N_8581);
xor U12611 (N_12611,N_12125,N_10054);
nor U12612 (N_12612,N_7830,N_12419);
nand U12613 (N_12613,N_6948,N_11480);
and U12614 (N_12614,N_6362,N_8917);
and U12615 (N_12615,N_11032,N_7765);
nor U12616 (N_12616,N_8803,N_6492);
nand U12617 (N_12617,N_10285,N_8208);
nor U12618 (N_12618,N_8492,N_9267);
nand U12619 (N_12619,N_6940,N_7055);
nor U12620 (N_12620,N_8083,N_7074);
nand U12621 (N_12621,N_8558,N_6595);
nor U12622 (N_12622,N_9959,N_10174);
nor U12623 (N_12623,N_11455,N_9180);
nor U12624 (N_12624,N_11087,N_10447);
xor U12625 (N_12625,N_6648,N_8778);
and U12626 (N_12626,N_6372,N_7265);
and U12627 (N_12627,N_9680,N_12352);
nor U12628 (N_12628,N_8190,N_6651);
and U12629 (N_12629,N_10706,N_11046);
nor U12630 (N_12630,N_10435,N_10260);
nand U12631 (N_12631,N_10956,N_8744);
nor U12632 (N_12632,N_11843,N_10959);
or U12633 (N_12633,N_11578,N_11249);
or U12634 (N_12634,N_8354,N_9593);
nand U12635 (N_12635,N_7859,N_10378);
or U12636 (N_12636,N_9710,N_9584);
and U12637 (N_12637,N_11538,N_9646);
and U12638 (N_12638,N_6330,N_8910);
nor U12639 (N_12639,N_10904,N_11565);
and U12640 (N_12640,N_9262,N_6688);
nand U12641 (N_12641,N_12245,N_8884);
or U12642 (N_12642,N_8928,N_8996);
nand U12643 (N_12643,N_12151,N_6819);
and U12644 (N_12644,N_12311,N_7438);
nor U12645 (N_12645,N_6497,N_10610);
nor U12646 (N_12646,N_8007,N_11683);
nor U12647 (N_12647,N_10503,N_11855);
nor U12648 (N_12648,N_12152,N_11220);
and U12649 (N_12649,N_10939,N_7293);
nor U12650 (N_12650,N_10894,N_8976);
xnor U12651 (N_12651,N_11318,N_11196);
and U12652 (N_12652,N_9504,N_10029);
and U12653 (N_12653,N_9853,N_11385);
and U12654 (N_12654,N_7028,N_7250);
or U12655 (N_12655,N_11921,N_8526);
nor U12656 (N_12656,N_7577,N_7856);
nand U12657 (N_12657,N_7512,N_6354);
or U12658 (N_12658,N_10937,N_11393);
nor U12659 (N_12659,N_7168,N_7827);
or U12660 (N_12660,N_9633,N_8637);
or U12661 (N_12661,N_7875,N_7780);
or U12662 (N_12662,N_9429,N_8677);
nand U12663 (N_12663,N_9746,N_10968);
xor U12664 (N_12664,N_8018,N_9064);
nor U12665 (N_12665,N_6543,N_10152);
and U12666 (N_12666,N_7164,N_9376);
nor U12667 (N_12667,N_12030,N_12131);
and U12668 (N_12668,N_6444,N_7452);
and U12669 (N_12669,N_11001,N_7855);
nand U12670 (N_12670,N_6631,N_9324);
and U12671 (N_12671,N_10144,N_6312);
and U12672 (N_12672,N_12465,N_7099);
or U12673 (N_12673,N_9399,N_11842);
and U12674 (N_12674,N_10338,N_9921);
nand U12675 (N_12675,N_8225,N_7337);
and U12676 (N_12676,N_9153,N_8093);
nand U12677 (N_12677,N_10487,N_11601);
nor U12678 (N_12678,N_9587,N_11394);
and U12679 (N_12679,N_8004,N_8261);
nand U12680 (N_12680,N_9624,N_9177);
and U12681 (N_12681,N_10393,N_8304);
or U12682 (N_12682,N_9146,N_12178);
xor U12683 (N_12683,N_8451,N_11655);
nand U12684 (N_12684,N_12108,N_11517);
and U12685 (N_12685,N_9740,N_10326);
and U12686 (N_12686,N_12217,N_7501);
nand U12687 (N_12687,N_12175,N_9302);
nand U12688 (N_12688,N_7922,N_9668);
nand U12689 (N_12689,N_7915,N_9883);
and U12690 (N_12690,N_11253,N_9341);
and U12691 (N_12691,N_7111,N_6630);
nand U12692 (N_12692,N_10450,N_11787);
or U12693 (N_12693,N_11777,N_9684);
or U12694 (N_12694,N_12411,N_8972);
nor U12695 (N_12695,N_12499,N_11229);
nand U12696 (N_12696,N_9910,N_7112);
or U12697 (N_12697,N_7027,N_6703);
nor U12698 (N_12698,N_7683,N_11066);
and U12699 (N_12699,N_7649,N_10824);
or U12700 (N_12700,N_6297,N_8035);
xor U12701 (N_12701,N_10811,N_9531);
nand U12702 (N_12702,N_10093,N_10899);
xnor U12703 (N_12703,N_11607,N_8351);
or U12704 (N_12704,N_7300,N_10961);
and U12705 (N_12705,N_11791,N_9575);
or U12706 (N_12706,N_11488,N_9778);
or U12707 (N_12707,N_11561,N_10823);
nor U12708 (N_12708,N_10298,N_10161);
nand U12709 (N_12709,N_8640,N_12110);
nor U12710 (N_12710,N_10976,N_11267);
or U12711 (N_12711,N_10919,N_6526);
or U12712 (N_12712,N_10603,N_7720);
xnor U12713 (N_12713,N_11300,N_11117);
nand U12714 (N_12714,N_9536,N_9637);
nand U12715 (N_12715,N_10341,N_11881);
xnor U12716 (N_12716,N_8523,N_11808);
nor U12717 (N_12717,N_12051,N_9889);
or U12718 (N_12718,N_11387,N_11116);
xor U12719 (N_12719,N_9068,N_11812);
nand U12720 (N_12720,N_10669,N_11124);
or U12721 (N_12721,N_6692,N_10627);
nand U12722 (N_12722,N_6760,N_6259);
nand U12723 (N_12723,N_11102,N_11265);
or U12724 (N_12724,N_12136,N_10884);
nor U12725 (N_12725,N_7609,N_7766);
and U12726 (N_12726,N_12301,N_7684);
nand U12727 (N_12727,N_6873,N_10857);
nor U12728 (N_12728,N_8671,N_10246);
nor U12729 (N_12729,N_6413,N_8052);
and U12730 (N_12730,N_10075,N_8909);
nand U12731 (N_12731,N_7659,N_10438);
nor U12732 (N_12732,N_9037,N_7785);
or U12733 (N_12733,N_10031,N_10010);
xor U12734 (N_12734,N_9574,N_10304);
nand U12735 (N_12735,N_9511,N_12360);
or U12736 (N_12736,N_9526,N_10891);
or U12737 (N_12737,N_9832,N_7774);
nand U12738 (N_12738,N_12070,N_7086);
xnor U12739 (N_12739,N_11986,N_8068);
nand U12740 (N_12740,N_6722,N_11980);
and U12741 (N_12741,N_9044,N_12272);
nand U12742 (N_12742,N_8174,N_11539);
nor U12743 (N_12743,N_10167,N_9839);
or U12744 (N_12744,N_11793,N_7625);
xnor U12745 (N_12745,N_10506,N_10016);
xnor U12746 (N_12746,N_8395,N_8595);
or U12747 (N_12747,N_7534,N_9172);
nand U12748 (N_12748,N_7018,N_12489);
nand U12749 (N_12749,N_9160,N_12028);
and U12750 (N_12750,N_8445,N_9948);
nand U12751 (N_12751,N_6551,N_9880);
nand U12752 (N_12752,N_9287,N_12474);
nand U12753 (N_12753,N_9008,N_6912);
nor U12754 (N_12754,N_10567,N_7969);
and U12755 (N_12755,N_12408,N_12043);
or U12756 (N_12756,N_9856,N_10419);
and U12757 (N_12757,N_7662,N_6707);
and U12758 (N_12758,N_9186,N_8951);
and U12759 (N_12759,N_11591,N_11215);
and U12760 (N_12760,N_11574,N_11653);
xor U12761 (N_12761,N_6861,N_7463);
nand U12762 (N_12762,N_9449,N_6773);
xor U12763 (N_12763,N_11696,N_12325);
and U12764 (N_12764,N_8504,N_9470);
nand U12765 (N_12765,N_6597,N_6344);
nor U12766 (N_12766,N_9590,N_8094);
nor U12767 (N_12767,N_10550,N_11626);
nor U12768 (N_12768,N_11388,N_7916);
and U12769 (N_12769,N_7186,N_9085);
and U12770 (N_12770,N_8587,N_7671);
and U12771 (N_12771,N_7990,N_6877);
or U12772 (N_12772,N_9781,N_12193);
or U12773 (N_12773,N_9870,N_9552);
nor U12774 (N_12774,N_11799,N_6967);
xor U12775 (N_12775,N_10694,N_9466);
xor U12776 (N_12776,N_10807,N_6643);
and U12777 (N_12777,N_11877,N_7970);
and U12778 (N_12778,N_10962,N_10986);
and U12779 (N_12779,N_11975,N_8148);
nor U12780 (N_12780,N_10454,N_11902);
nand U12781 (N_12781,N_8651,N_8839);
nand U12782 (N_12782,N_6436,N_7389);
or U12783 (N_12783,N_9607,N_7742);
or U12784 (N_12784,N_10605,N_11157);
nand U12785 (N_12785,N_9215,N_11589);
or U12786 (N_12786,N_11557,N_11919);
or U12787 (N_12787,N_8715,N_8211);
or U12788 (N_12788,N_10431,N_7644);
and U12789 (N_12789,N_7278,N_9022);
or U12790 (N_12790,N_8446,N_10017);
and U12791 (N_12791,N_10015,N_7060);
and U12792 (N_12792,N_8943,N_7179);
or U12793 (N_12793,N_10267,N_10327);
or U12794 (N_12794,N_8957,N_6418);
or U12795 (N_12795,N_9543,N_8202);
nor U12796 (N_12796,N_7009,N_9546);
nand U12797 (N_12797,N_10071,N_8835);
nor U12798 (N_12798,N_12323,N_11869);
nor U12799 (N_12799,N_8575,N_7015);
xor U12800 (N_12800,N_8087,N_8118);
nor U12801 (N_12801,N_8991,N_9007);
and U12802 (N_12802,N_8855,N_7846);
and U12803 (N_12803,N_7914,N_11104);
nor U12804 (N_12804,N_7235,N_8880);
nand U12805 (N_12805,N_10387,N_7862);
or U12806 (N_12806,N_6486,N_9534);
and U12807 (N_12807,N_10273,N_12372);
nor U12808 (N_12808,N_11007,N_9102);
nand U12809 (N_12809,N_9184,N_10983);
nand U12810 (N_12810,N_6388,N_10221);
or U12811 (N_12811,N_11513,N_8854);
or U12812 (N_12812,N_8710,N_7991);
and U12813 (N_12813,N_11103,N_11340);
nor U12814 (N_12814,N_9041,N_6415);
and U12815 (N_12815,N_9250,N_6754);
and U12816 (N_12816,N_10206,N_9181);
nor U12817 (N_12817,N_9234,N_9423);
nor U12818 (N_12818,N_9836,N_8658);
nor U12819 (N_12819,N_7394,N_11351);
and U12820 (N_12820,N_12368,N_8485);
nor U12821 (N_12821,N_8728,N_8629);
and U12822 (N_12822,N_9978,N_9887);
nor U12823 (N_12823,N_10725,N_10540);
or U12824 (N_12824,N_7132,N_12387);
xnor U12825 (N_12825,N_8383,N_7918);
nand U12826 (N_12826,N_11495,N_6624);
nor U12827 (N_12827,N_8120,N_8237);
or U12828 (N_12828,N_8967,N_10476);
nand U12829 (N_12829,N_11597,N_8904);
xnor U12830 (N_12830,N_10879,N_8826);
or U12831 (N_12831,N_8021,N_7907);
or U12832 (N_12832,N_11199,N_6917);
nor U12833 (N_12833,N_6812,N_8040);
nand U12834 (N_12834,N_6321,N_11648);
nor U12835 (N_12835,N_10060,N_10826);
nand U12836 (N_12836,N_6733,N_9226);
nor U12837 (N_12837,N_11813,N_11624);
nor U12838 (N_12838,N_7114,N_11748);
nor U12839 (N_12839,N_7902,N_10202);
or U12840 (N_12840,N_12222,N_11708);
or U12841 (N_12841,N_7307,N_8376);
nand U12842 (N_12842,N_9764,N_9338);
and U12843 (N_12843,N_12388,N_10083);
xor U12844 (N_12844,N_12230,N_11280);
and U12845 (N_12845,N_8152,N_10668);
xor U12846 (N_12846,N_9402,N_10481);
nand U12847 (N_12847,N_10589,N_7585);
nand U12848 (N_12848,N_12226,N_10907);
or U12849 (N_12849,N_10492,N_9168);
nor U12850 (N_12850,N_7531,N_10649);
nand U12851 (N_12851,N_12098,N_6355);
xnor U12852 (N_12852,N_8682,N_12185);
nor U12853 (N_12853,N_9768,N_9712);
nand U12854 (N_12854,N_8438,N_11175);
nand U12855 (N_12855,N_7783,N_10987);
or U12856 (N_12856,N_11243,N_11957);
nor U12857 (N_12857,N_11917,N_7143);
nor U12858 (N_12858,N_9025,N_7986);
or U12859 (N_12859,N_6366,N_9158);
xnor U12860 (N_12860,N_11160,N_8543);
and U12861 (N_12861,N_11210,N_11450);
nand U12862 (N_12862,N_9486,N_8414);
nand U12863 (N_12863,N_11153,N_11268);
and U12864 (N_12864,N_6263,N_8885);
nand U12865 (N_12865,N_10301,N_7078);
nor U12866 (N_12866,N_6343,N_9187);
and U12867 (N_12867,N_9620,N_11531);
nor U12868 (N_12868,N_9194,N_9891);
nand U12869 (N_12869,N_7482,N_10291);
and U12870 (N_12870,N_11810,N_9276);
nand U12871 (N_12871,N_11325,N_7269);
or U12872 (N_12872,N_7837,N_7222);
xor U12873 (N_12873,N_12303,N_9914);
nor U12874 (N_12874,N_9527,N_7681);
nand U12875 (N_12875,N_7857,N_6852);
or U12876 (N_12876,N_7272,N_10717);
nor U12877 (N_12877,N_8366,N_9282);
and U12878 (N_12878,N_10319,N_11427);
and U12879 (N_12879,N_11219,N_7029);
or U12880 (N_12880,N_12355,N_7747);
nand U12881 (N_12881,N_11365,N_7306);
nor U12882 (N_12882,N_6994,N_11804);
or U12883 (N_12883,N_10596,N_6476);
nand U12884 (N_12884,N_9212,N_10308);
nand U12885 (N_12885,N_7960,N_10057);
or U12886 (N_12886,N_7645,N_6357);
nand U12887 (N_12887,N_9174,N_11950);
nand U12888 (N_12888,N_6378,N_10139);
nor U12889 (N_12889,N_7812,N_11546);
or U12890 (N_12890,N_11060,N_9582);
nand U12891 (N_12891,N_11623,N_9991);
nand U12892 (N_12892,N_8140,N_6814);
nand U12893 (N_12893,N_8270,N_6277);
and U12894 (N_12894,N_8630,N_11471);
nand U12895 (N_12895,N_11794,N_9818);
nand U12896 (N_12896,N_7149,N_7860);
nand U12897 (N_12897,N_6850,N_9152);
and U12898 (N_12898,N_6695,N_8013);
nand U12899 (N_12899,N_11553,N_11753);
nor U12900 (N_12900,N_9062,N_11478);
or U12901 (N_12901,N_10126,N_9519);
or U12902 (N_12902,N_6448,N_9931);
and U12903 (N_12903,N_8221,N_12133);
nor U12904 (N_12904,N_6516,N_11307);
nor U12905 (N_12905,N_10084,N_9828);
nor U12906 (N_12906,N_9330,N_6629);
nand U12907 (N_12907,N_10679,N_7435);
nor U12908 (N_12908,N_7936,N_12198);
nand U12909 (N_12909,N_8706,N_12066);
nand U12910 (N_12910,N_10127,N_11465);
or U12911 (N_12911,N_7667,N_9580);
nand U12912 (N_12912,N_11074,N_8605);
nand U12913 (N_12913,N_12417,N_10365);
nor U12914 (N_12914,N_8937,N_7178);
or U12915 (N_12915,N_9191,N_10598);
nand U12916 (N_12916,N_6766,N_8325);
nor U12917 (N_12917,N_8912,N_12234);
and U12918 (N_12918,N_6751,N_9331);
nand U12919 (N_12919,N_8056,N_8328);
and U12920 (N_12920,N_12276,N_10632);
or U12921 (N_12921,N_11177,N_11867);
and U12922 (N_12922,N_8747,N_11092);
or U12923 (N_12923,N_11672,N_10032);
xor U12924 (N_12924,N_12264,N_10413);
xnor U12925 (N_12925,N_10693,N_9804);
nand U12926 (N_12926,N_9048,N_10788);
nand U12927 (N_12927,N_11911,N_7823);
nor U12928 (N_12928,N_9424,N_9583);
nand U12929 (N_12929,N_12404,N_11693);
nor U12930 (N_12930,N_11935,N_11840);
or U12931 (N_12931,N_11145,N_9610);
or U12932 (N_12932,N_8771,N_8307);
nor U12933 (N_12933,N_11809,N_8765);
nor U12934 (N_12934,N_11111,N_11470);
and U12935 (N_12935,N_6723,N_7954);
or U12936 (N_12936,N_11389,N_11963);
xor U12937 (N_12937,N_12467,N_9036);
nor U12938 (N_12938,N_11943,N_9846);
nor U12939 (N_12939,N_8670,N_7949);
nor U12940 (N_12940,N_8193,N_10027);
or U12941 (N_12941,N_11982,N_6328);
nand U12942 (N_12942,N_9865,N_8310);
nor U12943 (N_12943,N_9123,N_7993);
nor U12944 (N_12944,N_9563,N_9678);
and U12945 (N_12945,N_10467,N_6916);
nand U12946 (N_12946,N_6813,N_10617);
and U12947 (N_12947,N_7805,N_9506);
nand U12948 (N_12948,N_12441,N_7887);
and U12949 (N_12949,N_7456,N_8589);
nor U12950 (N_12950,N_8867,N_10478);
or U12951 (N_12951,N_8398,N_9029);
and U12952 (N_12952,N_11718,N_6557);
xnor U12953 (N_12953,N_8322,N_10382);
xnor U12954 (N_12954,N_8073,N_12195);
nand U12955 (N_12955,N_6608,N_8157);
nand U12956 (N_12956,N_11324,N_6927);
nand U12957 (N_12957,N_10403,N_9204);
nand U12958 (N_12958,N_7664,N_10154);
nand U12959 (N_12959,N_10284,N_12026);
or U12960 (N_12960,N_7944,N_6997);
nor U12961 (N_12961,N_9797,N_9848);
nor U12962 (N_12962,N_7570,N_7525);
xor U12963 (N_12963,N_9196,N_8738);
xor U12964 (N_12964,N_9455,N_10347);
nor U12965 (N_12965,N_7317,N_8344);
and U12966 (N_12966,N_9339,N_9723);
or U12967 (N_12967,N_9550,N_8751);
xnor U12968 (N_12968,N_10289,N_7282);
or U12969 (N_12969,N_11409,N_7711);
nor U12970 (N_12970,N_8048,N_9393);
nor U12971 (N_12971,N_10643,N_7934);
nand U12972 (N_12972,N_10854,N_8729);
or U12973 (N_12973,N_12101,N_10141);
nand U12974 (N_12974,N_6957,N_6348);
and U12975 (N_12975,N_11155,N_8986);
and U12976 (N_12976,N_11187,N_7931);
nor U12977 (N_12977,N_11934,N_9909);
nand U12978 (N_12978,N_8962,N_12395);
xor U12979 (N_12979,N_8737,N_10876);
or U12980 (N_12980,N_10774,N_7749);
or U12981 (N_12981,N_8495,N_9343);
nor U12982 (N_12982,N_8506,N_10594);
nor U12983 (N_12983,N_6909,N_7636);
nand U12984 (N_12984,N_7020,N_11706);
or U12985 (N_12985,N_12184,N_8355);
or U12986 (N_12986,N_9219,N_10885);
and U12987 (N_12987,N_11670,N_8284);
nor U12988 (N_12988,N_9941,N_11003);
nor U12989 (N_12989,N_12046,N_7848);
and U12990 (N_12990,N_11973,N_12349);
or U12991 (N_12991,N_10763,N_11885);
and U12992 (N_12992,N_8480,N_8931);
nor U12993 (N_12993,N_7666,N_10125);
nand U12994 (N_12994,N_9987,N_7260);
or U12995 (N_12995,N_6653,N_8621);
nor U12996 (N_12996,N_9368,N_8337);
nor U12997 (N_12997,N_6992,N_8339);
nor U12998 (N_12998,N_9578,N_11523);
nand U12999 (N_12999,N_7082,N_12258);
or U13000 (N_13000,N_11483,N_7733);
nand U13001 (N_13001,N_7032,N_6398);
or U13002 (N_13002,N_9016,N_11206);
nor U13003 (N_13003,N_6293,N_8948);
nor U13004 (N_13004,N_10977,N_6690);
and U13005 (N_13005,N_11178,N_7631);
xor U13006 (N_13006,N_7989,N_8817);
or U13007 (N_13007,N_8524,N_7466);
or U13008 (N_13008,N_8689,N_6567);
nand U13009 (N_13009,N_10868,N_7424);
nor U13010 (N_13010,N_7619,N_6535);
xor U13011 (N_13011,N_11512,N_6386);
nand U13012 (N_13012,N_6749,N_9609);
and U13013 (N_13013,N_8644,N_6477);
xnor U13014 (N_13014,N_9240,N_10026);
xnor U13015 (N_13015,N_7320,N_11719);
nor U13016 (N_13016,N_11089,N_12284);
and U13017 (N_13017,N_6449,N_8105);
and U13018 (N_13018,N_7243,N_10531);
or U13019 (N_13019,N_9919,N_11649);
nor U13020 (N_13020,N_7416,N_6500);
nor U13021 (N_13021,N_11348,N_6659);
xnor U13022 (N_13022,N_6901,N_7391);
nand U13023 (N_13023,N_9096,N_10275);
and U13024 (N_13024,N_9242,N_7984);
nor U13025 (N_13025,N_8549,N_9644);
nand U13026 (N_13026,N_6939,N_7948);
nor U13027 (N_13027,N_6589,N_6284);
xor U13028 (N_13028,N_12153,N_11977);
or U13029 (N_13029,N_8832,N_11675);
nor U13030 (N_13030,N_10078,N_9755);
and U13031 (N_13031,N_9632,N_10228);
nor U13032 (N_13032,N_6887,N_7520);
or U13033 (N_13033,N_6361,N_11127);
nor U13034 (N_13034,N_10195,N_12342);
and U13035 (N_13035,N_11308,N_9573);
and U13036 (N_13036,N_11688,N_9612);
nor U13037 (N_13037,N_11293,N_7497);
or U13038 (N_13038,N_10767,N_9442);
nor U13039 (N_13039,N_9689,N_8278);
and U13040 (N_13040,N_8573,N_8784);
or U13041 (N_13041,N_11964,N_6752);
nor U13042 (N_13042,N_9868,N_10177);
nand U13043 (N_13043,N_9945,N_11588);
and U13044 (N_13044,N_9178,N_9769);
nand U13045 (N_13045,N_8984,N_7346);
nand U13046 (N_13046,N_6790,N_9947);
and U13047 (N_13047,N_10019,N_8648);
and U13048 (N_13048,N_7461,N_10035);
nand U13049 (N_13049,N_11526,N_6904);
nand U13050 (N_13050,N_6718,N_10760);
nand U13051 (N_13051,N_6387,N_7000);
xnor U13052 (N_13052,N_9365,N_9130);
and U13053 (N_13053,N_7342,N_6700);
nor U13054 (N_13054,N_8722,N_11367);
and U13055 (N_13055,N_12167,N_9392);
nor U13056 (N_13056,N_11368,N_11687);
or U13057 (N_13057,N_10190,N_11671);
nor U13058 (N_13058,N_8655,N_6894);
or U13059 (N_13059,N_12298,N_11673);
xnor U13060 (N_13060,N_7703,N_6868);
xnor U13061 (N_13061,N_10164,N_10812);
or U13062 (N_13062,N_10953,N_10948);
nand U13063 (N_13063,N_8547,N_8302);
nand U13064 (N_13064,N_7448,N_8638);
and U13065 (N_13065,N_6941,N_9541);
and U13066 (N_13066,N_9452,N_10180);
or U13067 (N_13067,N_10142,N_9164);
nand U13068 (N_13068,N_6442,N_8119);
and U13069 (N_13069,N_8939,N_11129);
nand U13070 (N_13070,N_6736,N_6875);
nor U13071 (N_13071,N_9469,N_10675);
or U13072 (N_13072,N_7640,N_9697);
nor U13073 (N_13073,N_9895,N_7669);
nand U13074 (N_13074,N_10222,N_9904);
nor U13075 (N_13075,N_7994,N_10600);
nand U13076 (N_13076,N_7335,N_9375);
nor U13077 (N_13077,N_6517,N_10817);
and U13078 (N_13078,N_9690,N_11723);
nand U13079 (N_13079,N_7998,N_9000);
nor U13080 (N_13080,N_9059,N_7652);
nand U13081 (N_13081,N_9065,N_10189);
and U13082 (N_13082,N_12326,N_7634);
xor U13083 (N_13083,N_11602,N_6446);
or U13084 (N_13084,N_11222,N_12252);
and U13085 (N_13085,N_7495,N_9699);
nand U13086 (N_13086,N_6787,N_6633);
nor U13087 (N_13087,N_9679,N_9143);
or U13088 (N_13088,N_9395,N_7757);
and U13089 (N_13089,N_8820,N_7601);
or U13090 (N_13090,N_6420,N_7401);
xnor U13091 (N_13091,N_12491,N_9605);
nand U13092 (N_13092,N_11831,N_8752);
nor U13093 (N_13093,N_11923,N_7129);
or U13094 (N_13094,N_11618,N_12260);
xor U13095 (N_13095,N_7038,N_10688);
nor U13096 (N_13096,N_7831,N_9367);
nor U13097 (N_13097,N_8283,N_12237);
or U13098 (N_13098,N_11135,N_8427);
and U13099 (N_13099,N_10793,N_6403);
nand U13100 (N_13100,N_6646,N_7439);
nand U13101 (N_13101,N_8426,N_11762);
nor U13102 (N_13102,N_11757,N_8877);
nand U13103 (N_13103,N_11765,N_7578);
xnor U13104 (N_13104,N_8330,N_9087);
xor U13105 (N_13105,N_10000,N_11398);
nor U13106 (N_13106,N_10944,N_7363);
or U13107 (N_13107,N_10350,N_7417);
or U13108 (N_13108,N_12350,N_8913);
and U13109 (N_13109,N_6578,N_8363);
nor U13110 (N_13110,N_9078,N_8433);
or U13111 (N_13111,N_7369,N_8562);
xor U13112 (N_13112,N_7437,N_9493);
nand U13113 (N_13113,N_10101,N_11824);
or U13114 (N_13114,N_7537,N_6410);
nand U13115 (N_13115,N_9760,N_11994);
xor U13116 (N_13116,N_10299,N_9256);
nand U13117 (N_13117,N_11514,N_7839);
or U13118 (N_13118,N_10842,N_10936);
xnor U13119 (N_13119,N_7195,N_12451);
nand U13120 (N_13120,N_9535,N_11521);
or U13121 (N_13121,N_10111,N_9027);
xor U13122 (N_13122,N_12106,N_10484);
or U13123 (N_13123,N_9956,N_11237);
nor U13124 (N_13124,N_9465,N_10452);
or U13125 (N_13125,N_11554,N_10089);
and U13126 (N_13126,N_11774,N_11269);
nand U13127 (N_13127,N_11099,N_9283);
nand U13128 (N_13128,N_6269,N_11327);
or U13129 (N_13129,N_11294,N_12044);
nor U13130 (N_13130,N_7462,N_9901);
and U13131 (N_13131,N_6339,N_8088);
nand U13132 (N_13132,N_8533,N_11421);
and U13133 (N_13133,N_10741,N_7119);
nor U13134 (N_13134,N_10954,N_11789);
and U13135 (N_13135,N_11691,N_8528);
nand U13136 (N_13136,N_6976,N_8974);
nand U13137 (N_13137,N_10993,N_7996);
nand U13138 (N_13138,N_7327,N_6588);
and U13139 (N_13139,N_11152,N_8632);
nor U13140 (N_13140,N_9260,N_10960);
or U13141 (N_13141,N_10563,N_6506);
or U13142 (N_13142,N_6943,N_8124);
and U13143 (N_13143,N_9496,N_11681);
or U13144 (N_13144,N_10124,N_10412);
nor U13145 (N_13145,N_6823,N_11158);
nand U13146 (N_13146,N_9342,N_8009);
or U13147 (N_13147,N_11015,N_12015);
nand U13148 (N_13148,N_8846,N_12188);
nand U13149 (N_13149,N_9420,N_12369);
and U13150 (N_13150,N_7923,N_9377);
nor U13151 (N_13151,N_7406,N_11941);
and U13152 (N_13152,N_8615,N_10076);
and U13153 (N_13153,N_10242,N_6775);
xor U13154 (N_13154,N_9705,N_9604);
nor U13155 (N_13155,N_8070,N_6878);
nand U13156 (N_13156,N_7680,N_7181);
nand U13157 (N_13157,N_7113,N_10425);
nor U13158 (N_13158,N_12037,N_10008);
and U13159 (N_13159,N_8050,N_12297);
and U13160 (N_13160,N_8173,N_7787);
nor U13161 (N_13161,N_11386,N_8827);
or U13162 (N_13162,N_9933,N_6661);
and U13163 (N_13163,N_8102,N_6435);
and U13164 (N_13164,N_10985,N_8198);
or U13165 (N_13165,N_8714,N_6475);
nand U13166 (N_13166,N_8107,N_8044);
nor U13167 (N_13167,N_6380,N_11028);
nand U13168 (N_13168,N_7551,N_6266);
nand U13169 (N_13169,N_12200,N_8218);
and U13170 (N_13170,N_7627,N_8596);
nand U13171 (N_13171,N_7184,N_7853);
nand U13172 (N_13172,N_7921,N_11355);
nor U13173 (N_13173,N_7796,N_8128);
nor U13174 (N_13174,N_10369,N_10009);
nand U13175 (N_13175,N_6617,N_6673);
or U13176 (N_13176,N_11037,N_10991);
or U13177 (N_13177,N_11379,N_9790);
xor U13178 (N_13178,N_11501,N_12389);
nand U13179 (N_13179,N_7740,N_10187);
nand U13180 (N_13180,N_8305,N_10335);
and U13181 (N_13181,N_11346,N_12415);
nor U13182 (N_13182,N_11533,N_8306);
xnor U13183 (N_13183,N_9967,N_6622);
nand U13184 (N_13184,N_6804,N_11744);
or U13185 (N_13185,N_10398,N_7023);
and U13186 (N_13186,N_9791,N_11952);
nand U13187 (N_13187,N_12210,N_7790);
nand U13188 (N_13188,N_11156,N_10250);
and U13189 (N_13189,N_10529,N_10915);
nand U13190 (N_13190,N_6383,N_9325);
nand U13191 (N_13191,N_8535,N_11316);
nor U13192 (N_13192,N_7612,N_8130);
nor U13193 (N_13193,N_12261,N_8932);
and U13194 (N_13194,N_6739,N_8584);
nor U13195 (N_13195,N_11283,N_7624);
or U13196 (N_13196,N_8980,N_11834);
nor U13197 (N_13197,N_11713,N_7062);
nand U13198 (N_13198,N_11166,N_9406);
and U13199 (N_13199,N_11130,N_10931);
or U13200 (N_13200,N_10485,N_10614);
or U13201 (N_13201,N_9458,N_6426);
or U13202 (N_13202,N_7194,N_7982);
and U13203 (N_13203,N_6445,N_10847);
xor U13204 (N_13204,N_7868,N_9151);
and U13205 (N_13205,N_9088,N_9617);
or U13206 (N_13206,N_11149,N_6637);
xnor U13207 (N_13207,N_10163,N_9049);
and U13208 (N_13208,N_10066,N_9722);
and U13209 (N_13209,N_12115,N_6685);
xnor U13210 (N_13210,N_9640,N_8385);
nor U13211 (N_13211,N_10998,N_11695);
or U13212 (N_13212,N_6962,N_11761);
or U13213 (N_13213,N_12021,N_6936);
or U13214 (N_13214,N_6478,N_7388);
and U13215 (N_13215,N_10886,N_11119);
or U13216 (N_13216,N_11951,N_8126);
nor U13217 (N_13217,N_8350,N_9515);
and U13218 (N_13218,N_11555,N_7870);
and U13219 (N_13219,N_11636,N_6784);
or U13220 (N_13220,N_10570,N_8016);
nand U13221 (N_13221,N_11643,N_10262);
or U13222 (N_13222,N_9386,N_10052);
xnor U13223 (N_13223,N_10344,N_11690);
and U13224 (N_13224,N_7958,N_8663);
nand U13225 (N_13225,N_6838,N_9327);
nor U13226 (N_13226,N_9521,N_10271);
and U13227 (N_13227,N_7786,N_8406);
or U13228 (N_13228,N_9432,N_7274);
nand U13229 (N_13229,N_11694,N_9443);
and U13230 (N_13230,N_11972,N_6373);
and U13231 (N_13231,N_10942,N_6920);
and U13232 (N_13232,N_9557,N_9354);
nand U13233 (N_13233,N_9576,N_7063);
or U13234 (N_13234,N_11891,N_8894);
or U13235 (N_13235,N_6996,N_11197);
xnor U13236 (N_13236,N_12402,N_10037);
nor U13237 (N_13237,N_10354,N_6279);
and U13238 (N_13238,N_12052,N_11663);
nor U13239 (N_13239,N_11931,N_10175);
nor U13240 (N_13240,N_11890,N_8285);
and U13241 (N_13241,N_9672,N_11069);
nor U13242 (N_13242,N_11370,N_7273);
or U13243 (N_13243,N_7893,N_7858);
nor U13244 (N_13244,N_8852,N_10077);
or U13245 (N_13245,N_7153,N_7138);
nand U13246 (N_13246,N_12339,N_6769);
and U13247 (N_13247,N_8254,N_9963);
and U13248 (N_13248,N_9332,N_11615);
and U13249 (N_13249,N_7731,N_11788);
or U13250 (N_13250,N_6626,N_7555);
or U13251 (N_13251,N_9288,N_7939);
or U13252 (N_13252,N_6317,N_11710);
and U13253 (N_13253,N_8842,N_10964);
nand U13254 (N_13254,N_9958,N_8739);
and U13255 (N_13255,N_7500,N_6568);
nor U13256 (N_13256,N_9908,N_9803);
xor U13257 (N_13257,N_7535,N_7981);
nor U13258 (N_13258,N_7387,N_9547);
and U13259 (N_13259,N_9940,N_11617);
xor U13260 (N_13260,N_6358,N_12183);
and U13261 (N_13261,N_7161,N_9307);
xnor U13262 (N_13262,N_10579,N_10371);
xor U13263 (N_13263,N_12075,N_11853);
nand U13264 (N_13264,N_10690,N_7240);
and U13265 (N_13265,N_11536,N_10547);
nand U13266 (N_13266,N_7483,N_10063);
nand U13267 (N_13267,N_7019,N_7258);
nand U13268 (N_13268,N_11133,N_11321);
or U13269 (N_13269,N_8505,N_11566);
or U13270 (N_13270,N_9824,N_10443);
or U13271 (N_13271,N_10038,N_9655);
or U13272 (N_13272,N_7101,N_8356);
xnor U13273 (N_13273,N_7997,N_7568);
nor U13274 (N_13274,N_7515,N_8960);
or U13275 (N_13275,N_7377,N_10423);
nor U13276 (N_13276,N_12179,N_10616);
nor U13277 (N_13277,N_8993,N_9957);
and U13278 (N_13278,N_9254,N_6828);
or U13279 (N_13279,N_8950,N_7529);
nand U13280 (N_13280,N_10524,N_6407);
and U13281 (N_13281,N_12420,N_7177);
and U13282 (N_13282,N_11353,N_10505);
or U13283 (N_13283,N_12285,N_10896);
or U13284 (N_13284,N_7087,N_10292);
nor U13285 (N_13285,N_6925,N_7216);
or U13286 (N_13286,N_7292,N_9922);
and U13287 (N_13287,N_6563,N_10657);
or U13288 (N_13288,N_8171,N_7302);
nand U13289 (N_13289,N_10630,N_7484);
and U13290 (N_13290,N_7085,N_9453);
or U13291 (N_13291,N_12025,N_10489);
and U13292 (N_13292,N_10789,N_9378);
xnor U13293 (N_13293,N_8106,N_9539);
nor U13294 (N_13294,N_6721,N_6794);
nor U13295 (N_13295,N_6942,N_6496);
nand U13296 (N_13296,N_9484,N_7724);
nand U13297 (N_13297,N_9434,N_6559);
nor U13298 (N_13298,N_7303,N_8774);
and U13299 (N_13299,N_8390,N_12384);
nor U13300 (N_13300,N_8794,N_9685);
nor U13301 (N_13301,N_10272,N_6414);
nand U13302 (N_13302,N_8416,N_12228);
nor U13303 (N_13303,N_6309,N_7611);
and U13304 (N_13304,N_7351,N_9117);
nand U13305 (N_13305,N_11208,N_8789);
xnor U13306 (N_13306,N_9962,N_7228);
or U13307 (N_13307,N_10219,N_11550);
or U13308 (N_13308,N_9555,N_12448);
or U13309 (N_13309,N_8730,N_9682);
xnor U13310 (N_13310,N_10362,N_11279);
or U13311 (N_13311,N_6511,N_7117);
nand U13312 (N_13312,N_11310,N_6842);
and U13313 (N_13313,N_10946,N_10682);
and U13314 (N_13314,N_11096,N_8570);
and U13315 (N_13315,N_10735,N_11781);
and U13316 (N_13316,N_9097,N_9454);
or U13317 (N_13317,N_9829,N_11064);
or U13318 (N_13318,N_7459,N_10196);
and U13319 (N_13319,N_12320,N_9412);
nand U13320 (N_13320,N_8314,N_6989);
nor U13321 (N_13321,N_8411,N_10230);
nor U13322 (N_13322,N_12024,N_12199);
and U13323 (N_13323,N_9529,N_9860);
and U13324 (N_13324,N_8393,N_10379);
nor U13325 (N_13325,N_12109,N_6440);
and U13326 (N_13326,N_8359,N_6572);
nand U13327 (N_13327,N_7284,N_7241);
and U13328 (N_13328,N_10780,N_9615);
or U13329 (N_13329,N_6829,N_9659);
or U13330 (N_13330,N_12436,N_11476);
nand U13331 (N_13331,N_10809,N_12123);
nor U13332 (N_13332,N_6715,N_9071);
nand U13333 (N_13333,N_6937,N_12251);
and U13334 (N_13334,N_8684,N_12111);
nor U13335 (N_13335,N_11545,N_10343);
nand U13336 (N_13336,N_6482,N_11711);
and U13337 (N_13337,N_8611,N_7685);
nor U13338 (N_13338,N_7160,N_12270);
nor U13339 (N_13339,N_7729,N_7835);
nand U13340 (N_13340,N_11983,N_10235);
and U13341 (N_13341,N_9239,N_11477);
nand U13342 (N_13342,N_9163,N_12097);
or U13343 (N_13343,N_10783,N_7025);
nor U13344 (N_13344,N_7224,N_8251);
and U13345 (N_13345,N_7209,N_7583);
or U13346 (N_13346,N_6726,N_7908);
or U13347 (N_13347,N_12095,N_7398);
and U13348 (N_13348,N_8162,N_9193);
nor U13349 (N_13349,N_11849,N_10312);
xnor U13350 (N_13350,N_7097,N_10941);
nand U13351 (N_13351,N_6764,N_10158);
nand U13352 (N_13352,N_12223,N_11709);
xor U13353 (N_13353,N_8580,N_10434);
and U13354 (N_13354,N_9295,N_6510);
nor U13355 (N_13355,N_7832,N_6915);
or U13356 (N_13356,N_6691,N_7200);
and U13357 (N_13357,N_6923,N_6490);
and U13358 (N_13358,N_6881,N_8434);
or U13359 (N_13359,N_6374,N_10609);
nor U13360 (N_13360,N_8878,N_7980);
or U13361 (N_13361,N_12277,N_10482);
and U13362 (N_13362,N_10927,N_6561);
nor U13363 (N_13363,N_9127,N_9827);
and U13364 (N_13364,N_6285,N_11944);
nor U13365 (N_13365,N_10085,N_12105);
nand U13366 (N_13366,N_10039,N_7197);
nand U13367 (N_13367,N_8883,N_11584);
or U13368 (N_13368,N_7828,N_9537);
nand U13369 (N_13369,N_7541,N_7208);
nor U13370 (N_13370,N_9266,N_6419);
and U13371 (N_13371,N_11492,N_11487);
nand U13372 (N_13372,N_11045,N_12281);
nand U13373 (N_13373,N_7548,N_8635);
and U13374 (N_13374,N_9911,N_6865);
and U13375 (N_13375,N_7593,N_8815);
or U13376 (N_13376,N_7700,N_7358);
or U13377 (N_13377,N_8064,N_9858);
nand U13378 (N_13378,N_6254,N_11837);
and U13379 (N_13379,N_9663,N_12347);
or U13380 (N_13380,N_8736,N_12194);
nand U13381 (N_13381,N_10281,N_10205);
nor U13382 (N_13382,N_7769,N_9984);
nor U13383 (N_13383,N_11635,N_12438);
nor U13384 (N_13384,N_10699,N_11850);
nand U13385 (N_13385,N_7468,N_10072);
nand U13386 (N_13386,N_12405,N_11204);
and U13387 (N_13387,N_11100,N_6744);
nand U13388 (N_13388,N_12107,N_8753);
and U13389 (N_13389,N_9525,N_9844);
or U13390 (N_13390,N_11569,N_10297);
nand U13391 (N_13391,N_10286,N_11211);
and U13392 (N_13392,N_9892,N_6772);
nand U13393 (N_13393,N_7564,N_8591);
nand U13394 (N_13394,N_9602,N_7772);
nand U13395 (N_13395,N_8457,N_7485);
xnor U13396 (N_13396,N_9003,N_6550);
xnor U13397 (N_13397,N_7924,N_8941);
or U13398 (N_13398,N_9641,N_11148);
xnor U13399 (N_13399,N_11050,N_10633);
or U13400 (N_13400,N_7723,N_9060);
nand U13401 (N_13401,N_8988,N_8758);
nor U13402 (N_13402,N_6605,N_12391);
nand U13403 (N_13403,N_8464,N_11188);
nor U13404 (N_13404,N_11088,N_8109);
nand U13405 (N_13405,N_9654,N_8866);
or U13406 (N_13406,N_12267,N_6582);
nand U13407 (N_13407,N_11209,N_9222);
nor U13408 (N_13408,N_9490,N_12120);
or U13409 (N_13409,N_8191,N_9076);
nand U13410 (N_13410,N_11419,N_7793);
xnor U13411 (N_13411,N_9090,N_9255);
nand U13412 (N_13412,N_10798,N_9139);
and U13413 (N_13413,N_10792,N_10414);
nor U13414 (N_13414,N_12186,N_11873);
nand U13415 (N_13415,N_8282,N_9651);
nand U13416 (N_13416,N_7080,N_7472);
and U13417 (N_13417,N_7473,N_8419);
or U13418 (N_13418,N_6641,N_8405);
and U13419 (N_13419,N_6576,N_6883);
and U13420 (N_13420,N_11735,N_8271);
or U13421 (N_13421,N_10521,N_9451);
nand U13422 (N_13422,N_6738,N_10796);
and U13423 (N_13423,N_6762,N_8840);
and U13424 (N_13424,N_7775,N_12031);
or U13425 (N_13425,N_10582,N_10651);
nand U13426 (N_13426,N_7580,N_10128);
and U13427 (N_13427,N_9596,N_10498);
nor U13428 (N_13428,N_11113,N_8072);
nand U13429 (N_13429,N_10724,N_10972);
or U13430 (N_13430,N_8985,N_7450);
nand U13431 (N_13431,N_9067,N_8265);
nand U13432 (N_13432,N_7007,N_9373);
xnor U13433 (N_13433,N_11172,N_6827);
and U13434 (N_13434,N_11193,N_12310);
or U13435 (N_13435,N_8164,N_6955);
nand U13436 (N_13436,N_11179,N_7305);
or U13437 (N_13437,N_6385,N_10599);
nor U13438 (N_13438,N_7743,N_9289);
or U13439 (N_13439,N_9034,N_10933);
nand U13440 (N_13440,N_6876,N_12007);
or U13441 (N_13441,N_11537,N_11251);
nand U13442 (N_13442,N_11858,N_10509);
nor U13443 (N_13443,N_10938,N_8633);
or U13444 (N_13444,N_10541,N_8488);
nand U13445 (N_13445,N_8860,N_6984);
nand U13446 (N_13446,N_10466,N_10918);
or U13447 (N_13447,N_11530,N_10663);
nand U13448 (N_13448,N_7135,N_10320);
xor U13449 (N_13449,N_11170,N_8881);
or U13450 (N_13450,N_8027,N_9201);
or U13451 (N_13451,N_6613,N_10332);
xnor U13452 (N_13452,N_9613,N_7665);
nand U13453 (N_13453,N_6694,N_10828);
nor U13454 (N_13454,N_6884,N_10322);
or U13455 (N_13455,N_8708,N_7397);
nor U13456 (N_13456,N_9667,N_8220);
nor U13457 (N_13457,N_8697,N_7233);
xnor U13458 (N_13458,N_7088,N_10576);
nand U13459 (N_13459,N_8776,N_7380);
nand U13460 (N_13460,N_10263,N_9647);
nand U13461 (N_13461,N_7176,N_10411);
nand U13462 (N_13462,N_9788,N_10794);
or U13463 (N_13463,N_11518,N_7242);
and U13464 (N_13464,N_10537,N_7544);
nand U13465 (N_13465,N_7066,N_6710);
xor U13466 (N_13466,N_9372,N_8767);
xor U13467 (N_13467,N_7880,N_9436);
and U13468 (N_13468,N_8493,N_7232);
or U13469 (N_13469,N_9802,N_7359);
nand U13470 (N_13470,N_11689,N_8977);
nand U13471 (N_13471,N_9661,N_9730);
nand U13472 (N_13472,N_8933,N_9478);
and U13473 (N_13473,N_10024,N_9639);
or U13474 (N_13474,N_9862,N_12306);
nand U13475 (N_13475,N_12331,N_11918);
and U13476 (N_13476,N_7409,N_6777);
and U13477 (N_13477,N_12463,N_10979);
nor U13478 (N_13478,N_9943,N_9270);
or U13479 (N_13479,N_9394,N_7107);
nand U13480 (N_13480,N_8705,N_10754);
and U13481 (N_13481,N_12225,N_10331);
xnor U13482 (N_13482,N_11392,N_10134);
xnor U13483 (N_13483,N_10303,N_9635);
nor U13484 (N_13484,N_11665,N_6862);
and U13485 (N_13485,N_7836,N_6980);
or U13486 (N_13486,N_8111,N_7690);
or U13487 (N_13487,N_10978,N_11364);
or U13488 (N_13488,N_8113,N_12174);
nand U13489 (N_13489,N_11822,N_7965);
nor U13490 (N_13490,N_8871,N_9405);
or U13491 (N_13491,N_7441,N_10710);
nand U13492 (N_13492,N_9867,N_8491);
and U13493 (N_13493,N_7124,N_7714);
xnor U13494 (N_13494,N_7604,N_12182);
nand U13495 (N_13495,N_10795,N_11721);
xnor U13496 (N_13496,N_7725,N_7270);
or U13497 (N_13497,N_10023,N_8507);
nor U13498 (N_13498,N_8189,N_10359);
and U13499 (N_13499,N_8296,N_10697);
and U13500 (N_13500,N_7471,N_6945);
nor U13501 (N_13501,N_9721,N_6272);
xor U13502 (N_13502,N_6837,N_10107);
and U13503 (N_13503,N_11277,N_11301);
or U13504 (N_13504,N_8674,N_11469);
nand U13505 (N_13505,N_7048,N_9322);
nand U13506 (N_13506,N_6273,N_9009);
and U13507 (N_13507,N_11141,N_10122);
or U13508 (N_13508,N_11263,N_10043);
or U13509 (N_13509,N_6716,N_11820);
or U13510 (N_13510,N_7400,N_7106);
nand U13511 (N_13511,N_10405,N_8012);
nand U13512 (N_13512,N_12243,N_6770);
xnor U13513 (N_13513,N_6931,N_7496);
or U13514 (N_13514,N_9560,N_7146);
nand U13515 (N_13515,N_11737,N_6606);
and U13516 (N_13516,N_7928,N_11576);
xnor U13517 (N_13517,N_11183,N_12162);
nand U13518 (N_13518,N_10558,N_7108);
xor U13519 (N_13519,N_10178,N_6600);
and U13520 (N_13520,N_11520,N_11431);
nand U13521 (N_13521,N_11965,N_9540);
or U13522 (N_13522,N_10034,N_9881);
xor U13523 (N_13523,N_8911,N_6527);
xor U13524 (N_13524,N_8563,N_11645);
and U13525 (N_13525,N_6310,N_12283);
and U13526 (N_13526,N_11955,N_9894);
or U13527 (N_13527,N_10407,N_10999);
and U13528 (N_13528,N_6767,N_7657);
or U13529 (N_13529,N_7430,N_8219);
nor U13530 (N_13530,N_6457,N_8248);
xnor U13531 (N_13531,N_7042,N_10771);
and U13532 (N_13532,N_12470,N_8151);
or U13533 (N_13533,N_10349,N_7744);
and U13534 (N_13534,N_8639,N_10100);
or U13535 (N_13535,N_10160,N_7845);
or U13536 (N_13536,N_12289,N_10980);
nor U13537 (N_13537,N_6575,N_6545);
and U13538 (N_13538,N_6553,N_7806);
nor U13539 (N_13539,N_9634,N_10356);
or U13540 (N_13540,N_10495,N_11647);
or U13541 (N_13541,N_8275,N_6498);
nor U13542 (N_13542,N_10287,N_12327);
xor U13543 (N_13543,N_9149,N_10667);
nor U13544 (N_13544,N_7421,N_11802);
nand U13545 (N_13545,N_10903,N_7589);
and U13546 (N_13546,N_9026,N_8634);
nor U13547 (N_13547,N_12344,N_8641);
nor U13548 (N_13548,N_6307,N_6756);
nor U13549 (N_13549,N_6720,N_7522);
and U13550 (N_13550,N_12191,N_9448);
and U13551 (N_13551,N_12393,N_7094);
nand U13552 (N_13552,N_9066,N_7613);
nor U13553 (N_13553,N_9473,N_12096);
nor U13554 (N_13554,N_6826,N_9913);
or U13555 (N_13555,N_10924,N_6809);
and U13556 (N_13556,N_10102,N_6696);
and U13557 (N_13557,N_11425,N_8382);
nand U13558 (N_13558,N_11785,N_12227);
nor U13559 (N_13559,N_8358,N_8992);
or U13560 (N_13560,N_10940,N_11876);
and U13561 (N_13561,N_8659,N_11971);
nor U13562 (N_13562,N_9571,N_6755);
nand U13563 (N_13563,N_8342,N_7470);
xor U13564 (N_13564,N_10831,N_10266);
or U13565 (N_13565,N_8686,N_7929);
nor U13566 (N_13566,N_6351,N_7884);
xnor U13567 (N_13567,N_11974,N_8790);
nor U13568 (N_13568,N_9886,N_11908);
and U13569 (N_13569,N_7913,N_8417);
nand U13570 (N_13570,N_8822,N_8872);
nand U13571 (N_13571,N_10002,N_10088);
nor U13572 (N_13572,N_11900,N_9834);
and U13573 (N_13573,N_9977,N_10587);
and U13574 (N_13574,N_7940,N_12429);
and U13575 (N_13575,N_9728,N_7355);
and U13576 (N_13576,N_8368,N_9032);
nand U13577 (N_13577,N_11659,N_10569);
or U13578 (N_13578,N_7410,N_8707);
nand U13579 (N_13579,N_11535,N_6459);
nand U13580 (N_13580,N_7069,N_12034);
and U13581 (N_13581,N_8252,N_6712);
xor U13582 (N_13582,N_7533,N_8514);
nand U13583 (N_13583,N_10618,N_12019);
xnor U13584 (N_13584,N_7110,N_6699);
nor U13585 (N_13585,N_8043,N_6392);
or U13586 (N_13586,N_8028,N_6857);
nand U13587 (N_13587,N_12224,N_8458);
or U13588 (N_13588,N_11173,N_6472);
or U13589 (N_13589,N_11165,N_12218);
and U13590 (N_13590,N_10732,N_12287);
nand U13591 (N_13591,N_10843,N_9734);
and U13592 (N_13592,N_7571,N_10620);
and U13593 (N_13593,N_9903,N_10775);
nor U13594 (N_13594,N_7402,N_9869);
nand U13595 (N_13595,N_11005,N_9360);
xor U13596 (N_13596,N_7290,N_12197);
nor U13597 (N_13597,N_6502,N_9334);
xnor U13598 (N_13598,N_7314,N_8796);
xnor U13599 (N_13599,N_8949,N_6250);
nor U13600 (N_13600,N_11362,N_10821);
or U13601 (N_13601,N_12257,N_12266);
and U13602 (N_13602,N_6320,N_8413);
or U13603 (N_13603,N_6602,N_7354);
or U13604 (N_13604,N_11954,N_6461);
xor U13605 (N_13605,N_12335,N_9488);
xor U13606 (N_13606,N_8273,N_7876);
and U13607 (N_13607,N_8755,N_11115);
nand U13608 (N_13608,N_7340,N_6818);
nor U13609 (N_13609,N_12263,N_11415);
and U13610 (N_13610,N_7933,N_12085);
or U13611 (N_13611,N_7262,N_11722);
or U13612 (N_13612,N_8989,N_10863);
xor U13613 (N_13613,N_9572,N_6845);
xor U13614 (N_13614,N_7935,N_7202);
nand U13615 (N_13615,N_8695,N_11137);
and U13616 (N_13616,N_7079,N_8750);
nand U13617 (N_13617,N_10883,N_8527);
or U13618 (N_13618,N_8929,N_7365);
or U13619 (N_13619,N_6566,N_10892);
nor U13620 (N_13620,N_11356,N_7159);
or U13621 (N_13621,N_11377,N_7336);
nor U13622 (N_13622,N_8474,N_6389);
nor U13623 (N_13623,N_11857,N_11004);
and U13624 (N_13624,N_6778,N_6693);
and U13625 (N_13625,N_8326,N_6911);
nor U13626 (N_13626,N_8889,N_7481);
xnor U13627 (N_13627,N_7956,N_7084);
xnor U13628 (N_13628,N_9503,N_7971);
nand U13629 (N_13629,N_9785,N_8779);
and U13630 (N_13630,N_10282,N_7075);
xnor U13631 (N_13631,N_8761,N_8078);
and U13632 (N_13632,N_8460,N_10430);
nor U13633 (N_13633,N_7021,N_6758);
or U13634 (N_13634,N_7165,N_9558);
and U13635 (N_13635,N_12102,N_9681);
nand U13636 (N_13636,N_6253,N_11245);
or U13637 (N_13637,N_10117,N_7248);
xnor U13638 (N_13638,N_10472,N_11715);
xnor U13639 (N_13639,N_12156,N_12213);
and U13640 (N_13640,N_6437,N_7726);
xnor U13641 (N_13641,N_7022,N_10460);
nor U13642 (N_13642,N_9742,N_10645);
and U13643 (N_13643,N_9798,N_7395);
nand U13644 (N_13644,N_12394,N_11186);
nand U13645 (N_13645,N_7713,N_10442);
and U13646 (N_13646,N_8032,N_8169);
nor U13647 (N_13647,N_11960,N_7217);
xnor U13648 (N_13648,N_9706,N_6368);
nor U13649 (N_13649,N_9771,N_7411);
and U13650 (N_13650,N_8809,N_8586);
and U13651 (N_13651,N_6808,N_8509);
nor U13652 (N_13652,N_11080,N_7927);
nor U13653 (N_13653,N_12359,N_9400);
and U13654 (N_13654,N_8076,N_7732);
and U13655 (N_13655,N_10848,N_10932);
xor U13656 (N_13656,N_7523,N_10698);
and U13657 (N_13657,N_12065,N_11559);
nand U13658 (N_13658,N_8762,N_6474);
or U13659 (N_13659,N_11112,N_10129);
xnor U13660 (N_13660,N_7131,N_11896);
or U13661 (N_13661,N_11118,N_10213);
nand U13662 (N_13662,N_9074,N_10965);
nand U13663 (N_13663,N_9169,N_11195);
nor U13664 (N_13664,N_9554,N_6462);
or U13665 (N_13665,N_8168,N_7844);
nand U13666 (N_13666,N_7623,N_9625);
nor U13667 (N_13667,N_12088,N_8410);
and U13668 (N_13668,N_11223,N_12475);
or U13669 (N_13669,N_7428,N_11341);
nand U13670 (N_13670,N_11094,N_11482);
nand U13671 (N_13671,N_12016,N_10901);
or U13672 (N_13672,N_7514,N_12009);
nor U13673 (N_13673,N_10516,N_9950);
nand U13674 (N_13674,N_12003,N_7492);
xor U13675 (N_13675,N_11563,N_11582);
nor U13676 (N_13676,N_8453,N_8712);
nand U13677 (N_13677,N_10574,N_9816);
nor U13678 (N_13678,N_11463,N_10893);
xnor U13679 (N_13679,N_6408,N_7833);
nor U13680 (N_13680,N_9258,N_8367);
and U13681 (N_13681,N_9483,N_11323);
nand U13682 (N_13682,N_9556,N_6765);
and U13683 (N_13683,N_12140,N_10786);
or U13684 (N_13684,N_7718,N_8716);
nor U13685 (N_13685,N_7189,N_10840);
or U13686 (N_13686,N_11552,N_11567);
xnor U13687 (N_13687,N_7532,N_7259);
nor U13688 (N_13688,N_8935,N_11298);
and U13689 (N_13689,N_8723,N_8481);
nand U13690 (N_13690,N_7985,N_8646);
or U13691 (N_13691,N_9732,N_6616);
nor U13692 (N_13692,N_12333,N_9094);
or U13693 (N_13693,N_6513,N_10420);
and U13694 (N_13694,N_8975,N_11289);
or U13695 (N_13695,N_8161,N_9329);
nor U13696 (N_13696,N_8520,N_12017);
nor U13697 (N_13697,N_12386,N_8699);
or U13698 (N_13698,N_12472,N_10631);
or U13699 (N_13699,N_12392,N_11236);
nor U13700 (N_13700,N_11632,N_6815);
nand U13701 (N_13701,N_7776,N_11945);
nor U13702 (N_13702,N_11432,N_7309);
xor U13703 (N_13703,N_11084,N_12023);
or U13704 (N_13704,N_7310,N_9333);
nor U13705 (N_13705,N_7479,N_11200);
nor U13706 (N_13706,N_10606,N_11067);
nor U13707 (N_13707,N_12362,N_6356);
nor U13708 (N_13708,N_10436,N_8066);
and U13709 (N_13709,N_7379,N_12290);
nor U13710 (N_13710,N_10255,N_11870);
xnor U13711 (N_13711,N_8002,N_12458);
nand U13712 (N_13712,N_11776,N_12457);
and U13713 (N_13713,N_7658,N_7668);
nand U13714 (N_13714,N_7341,N_6900);
nor U13715 (N_13715,N_8176,N_8089);
and U13716 (N_13716,N_7538,N_6705);
nor U13717 (N_13717,N_10593,N_10113);
or U13718 (N_13718,N_7076,N_11040);
and U13719 (N_13719,N_11987,N_9166);
and U13720 (N_13720,N_10376,N_12396);
or U13721 (N_13721,N_12112,N_7162);
xnor U13722 (N_13722,N_10624,N_7204);
xor U13723 (N_13723,N_10033,N_8092);
xor U13724 (N_13724,N_11109,N_10214);
and U13725 (N_13725,N_7826,N_10386);
nand U13726 (N_13726,N_10994,N_8408);
nand U13727 (N_13727,N_6276,N_8745);
and U13728 (N_13728,N_11854,N_8841);
and U13729 (N_13729,N_10087,N_6932);
or U13730 (N_13730,N_8423,N_10982);
xnor U13731 (N_13731,N_12135,N_7253);
or U13732 (N_13732,N_8925,N_9072);
nand U13733 (N_13733,N_6565,N_9369);
nor U13734 (N_13734,N_10249,N_6678);
or U13735 (N_13735,N_12302,N_9305);
or U13736 (N_13736,N_7294,N_9973);
nand U13737 (N_13737,N_10588,N_11309);
nor U13738 (N_13738,N_8341,N_7196);
nand U13739 (N_13739,N_8598,N_10746);
and U13740 (N_13740,N_9411,N_12319);
nor U13741 (N_13741,N_10646,N_6625);
or U13742 (N_13742,N_7256,N_11086);
and U13743 (N_13743,N_11464,N_10566);
or U13744 (N_13744,N_12042,N_7207);
xor U13745 (N_13745,N_9351,N_7128);
and U13746 (N_13746,N_8250,N_8540);
nor U13747 (N_13747,N_7758,N_6585);
nand U13748 (N_13748,N_8074,N_12240);
nand U13749 (N_13749,N_10648,N_10137);
nor U13750 (N_13750,N_9687,N_11953);
and U13751 (N_13751,N_9964,N_11864);
or U13752 (N_13752,N_10231,N_11126);
and U13753 (N_13753,N_12187,N_7366);
or U13754 (N_13754,N_7268,N_7917);
nand U13755 (N_13755,N_8059,N_10833);
nand U13756 (N_13756,N_9403,N_9438);
xor U13757 (N_13757,N_7390,N_11374);
nand U13758 (N_13758,N_8698,N_7014);
xor U13759 (N_13759,N_12341,N_6791);
and U13760 (N_13760,N_7490,N_11560);
nor U13761 (N_13761,N_11131,N_8946);
and U13762 (N_13762,N_10751,N_11700);
nand U13763 (N_13763,N_9799,N_9718);
or U13764 (N_13764,N_7219,N_11946);
nor U13765 (N_13765,N_9810,N_7673);
nor U13766 (N_13766,N_7620,N_11677);
or U13767 (N_13767,N_11017,N_6929);
or U13768 (N_13768,N_10818,N_10758);
and U13769 (N_13769,N_8582,N_9918);
nand U13770 (N_13770,N_8441,N_10409);
nand U13771 (N_13771,N_9603,N_7246);
nand U13772 (N_13772,N_6998,N_11562);
nand U13773 (N_13773,N_11000,N_11763);
and U13774 (N_13774,N_9023,N_9144);
nor U13775 (N_13775,N_10155,N_10908);
nand U13776 (N_13776,N_12255,N_7420);
and U13777 (N_13777,N_11871,N_9823);
and U13778 (N_13778,N_10474,N_6843);
and U13779 (N_13779,N_8858,N_7547);
nor U13780 (N_13780,N_11948,N_8389);
or U13781 (N_13781,N_6512,N_9820);
and U13782 (N_13782,N_6780,N_9441);
or U13783 (N_13783,N_8805,N_12160);
or U13784 (N_13784,N_7800,N_11738);
and U13785 (N_13785,N_6933,N_9896);
or U13786 (N_13786,N_12078,N_9920);
nor U13787 (N_13787,N_10421,N_9758);
or U13788 (N_13788,N_9614,N_10802);
or U13789 (N_13789,N_6831,N_9595);
nand U13790 (N_13790,N_12317,N_12071);
nand U13791 (N_13791,N_10372,N_7376);
and U13792 (N_13792,N_6623,N_12440);
nor U13793 (N_13793,N_10966,N_10888);
nor U13794 (N_13794,N_10683,N_11224);
and U13795 (N_13795,N_10560,N_9765);
nand U13796 (N_13796,N_6965,N_9999);
nand U13797 (N_13797,N_7591,N_10862);
nand U13798 (N_13798,N_10488,N_11685);
and U13799 (N_13799,N_7898,N_10608);
and U13800 (N_13800,N_11500,N_9176);
xnor U13801 (N_13801,N_9150,N_6987);
nand U13802 (N_13802,N_9045,N_7072);
nor U13803 (N_13803,N_7865,N_11899);
and U13804 (N_13804,N_6628,N_11244);
nand U13805 (N_13805,N_11396,N_9426);
or U13806 (N_13806,N_7721,N_7897);
or U13807 (N_13807,N_11758,N_10532);
xor U13808 (N_13808,N_7383,N_12375);
nor U13809 (N_13809,N_6371,N_10538);
and U13810 (N_13810,N_10461,N_11053);
or U13811 (N_13811,N_9893,N_7017);
nor U13812 (N_13812,N_8653,N_9713);
nand U13813 (N_13813,N_10963,N_10288);
nand U13814 (N_13814,N_10997,N_7142);
nand U13815 (N_13815,N_11532,N_8529);
and U13816 (N_13816,N_6741,N_9505);
nand U13817 (N_13817,N_6728,N_6918);
nor U13818 (N_13818,N_12137,N_7867);
or U13819 (N_13819,N_7909,N_10162);
nor U13820 (N_13820,N_7782,N_9190);
nand U13821 (N_13821,N_12062,N_11503);
or U13822 (N_13822,N_12484,N_6836);
nand U13823 (N_13823,N_7961,N_7104);
or U13824 (N_13824,N_8158,N_9012);
nor U13825 (N_13825,N_6405,N_9569);
nor U13826 (N_13826,N_12248,N_8030);
nor U13827 (N_13827,N_10065,N_8568);
and U13828 (N_13828,N_7127,N_9811);
nor U13829 (N_13829,N_11594,N_7886);
nor U13830 (N_13830,N_9358,N_10216);
and U13831 (N_13831,N_7840,N_8371);
nor U13832 (N_13832,N_7288,N_10650);
and U13833 (N_13833,N_8981,N_6316);
nand U13834 (N_13834,N_6959,N_9813);
and U13835 (N_13835,N_9081,N_6638);
or U13836 (N_13836,N_8336,N_9985);
or U13837 (N_13837,N_6463,N_10277);
or U13838 (N_13838,N_7368,N_11106);
xnor U13839 (N_13839,N_11336,N_8969);
and U13840 (N_13840,N_10861,N_6682);
nor U13841 (N_13841,N_11845,N_10480);
or U13842 (N_13842,N_7311,N_12139);
nand U13843 (N_13843,N_7125,N_11154);
nor U13844 (N_13844,N_11817,N_10441);
xnor U13845 (N_13845,N_7118,N_8011);
and U13846 (N_13846,N_10353,N_11863);
nor U13847 (N_13847,N_9111,N_10131);
or U13848 (N_13848,N_12450,N_10455);
xor U13849 (N_13849,N_6365,N_11271);
or U13850 (N_13850,N_12462,N_10834);
nor U13851 (N_13851,N_8143,N_7225);
nor U13852 (N_13852,N_8338,N_8373);
or U13853 (N_13853,N_10340,N_12406);
nor U13854 (N_13854,N_6621,N_7550);
and U13855 (N_13855,N_8890,N_7407);
or U13856 (N_13856,N_7573,N_7952);
or U13857 (N_13857,N_10728,N_7873);
and U13858 (N_13858,N_7622,N_11023);
xnor U13859 (N_13859,N_10370,N_9463);
or U13860 (N_13860,N_7449,N_11329);
and U13861 (N_13861,N_8896,N_10191);
or U13862 (N_13862,N_7517,N_10882);
and U13863 (N_13863,N_7979,N_11335);
or U13864 (N_13864,N_6737,N_11376);
or U13865 (N_13865,N_6548,N_8746);
xor U13866 (N_13866,N_7440,N_8207);
and U13867 (N_13867,N_8618,N_9082);
nand U13868 (N_13868,N_6953,N_10123);
or U13869 (N_13869,N_6562,N_8902);
or U13870 (N_13870,N_10446,N_8652);
and U13871 (N_13871,N_11361,N_6890);
and U13872 (N_13872,N_7572,N_10661);
and U13873 (N_13873,N_7442,N_7798);
or U13874 (N_13874,N_10952,N_10112);
nor U13875 (N_13875,N_8317,N_12316);
or U13876 (N_13876,N_9224,N_9292);
nor U13877 (N_13877,N_6732,N_11551);
nor U13878 (N_13878,N_7254,N_8139);
nand U13879 (N_13879,N_8614,N_6292);
nor U13880 (N_13880,N_8713,N_6642);
nor U13881 (N_13881,N_8289,N_11461);
or U13882 (N_13882,N_8331,N_6848);
nand U13883 (N_13883,N_11254,N_7299);
xor U13884 (N_13884,N_8554,N_7699);
nor U13885 (N_13885,N_8825,N_8213);
nand U13886 (N_13886,N_11764,N_9847);
or U13887 (N_13887,N_11075,N_11391);
or U13888 (N_13888,N_12189,N_8947);
nand U13889 (N_13889,N_9857,N_7851);
and U13890 (N_13890,N_7077,N_12401);
or U13891 (N_13891,N_10584,N_9888);
nand U13892 (N_13892,N_12433,N_9231);
nand U13893 (N_13893,N_9497,N_12238);
nand U13894 (N_13894,N_6341,N_10615);
nand U13895 (N_13895,N_6803,N_11442);
nor U13896 (N_13896,N_10012,N_11027);
nand U13897 (N_13897,N_7654,N_7230);
xnor U13898 (N_13898,N_7185,N_9433);
nor U13899 (N_13899,N_6898,N_10236);
and U13900 (N_13900,N_11147,N_11481);
xor U13901 (N_13901,N_10166,N_7010);
or U13902 (N_13902,N_11108,N_11342);
nor U13903 (N_13903,N_9585,N_10549);
or U13904 (N_13904,N_10475,N_8914);
xnor U13905 (N_13905,N_11246,N_10881);
xor U13906 (N_13906,N_12249,N_9487);
xnor U13907 (N_13907,N_7748,N_6376);
and U13908 (N_13908,N_11299,N_12481);
nand U13909 (N_13909,N_11234,N_11320);
or U13910 (N_13910,N_10042,N_11185);
or U13911 (N_13911,N_11295,N_8017);
and U13912 (N_13912,N_6663,N_11619);
nand U13913 (N_13913,N_10053,N_7013);
nor U13914 (N_13914,N_7698,N_11008);
nor U13915 (N_13915,N_10448,N_11938);
nor U13916 (N_13916,N_9821,N_8512);
or U13917 (N_13917,N_10923,N_7560);
and U13918 (N_13918,N_8600,N_8308);
and U13919 (N_13919,N_9259,N_7431);
or U13920 (N_13920,N_6855,N_8720);
or U13921 (N_13921,N_9361,N_6573);
and U13922 (N_13922,N_6493,N_11338);
nor U13923 (N_13923,N_8131,N_7187);
nor U13924 (N_13924,N_9992,N_7191);
or U13925 (N_13925,N_10181,N_6640);
nor U13926 (N_13926,N_11401,N_10870);
nand U13927 (N_13927,N_12061,N_6322);
nand U13928 (N_13928,N_9304,N_9735);
nand U13929 (N_13929,N_9033,N_8361);
nor U13930 (N_13930,N_6657,N_11872);
nand U13931 (N_13931,N_6797,N_6300);
nand U13932 (N_13932,N_11319,N_10392);
and U13933 (N_13933,N_9170,N_6729);
and U13934 (N_13934,N_9673,N_7313);
nor U13935 (N_13935,N_8280,N_12424);
xnor U13936 (N_13936,N_8156,N_9492);
nor U13937 (N_13937,N_10585,N_10169);
or U13938 (N_13938,N_7353,N_11042);
or U13939 (N_13939,N_8138,N_8104);
or U13940 (N_13940,N_10552,N_7362);
or U13941 (N_13941,N_6544,N_7822);
xor U13942 (N_13942,N_11034,N_11575);
nor U13943 (N_13943,N_6950,N_11484);
nor U13944 (N_13944,N_9134,N_7516);
or U13945 (N_13945,N_11741,N_9202);
and U13946 (N_13946,N_9321,N_7182);
and U13947 (N_13947,N_10733,N_7618);
nand U13948 (N_13948,N_9542,N_11906);
nand U13949 (N_13949,N_9645,N_9278);
or U13950 (N_13950,N_11628,N_11029);
and U13951 (N_13951,N_7951,N_9124);
xor U13952 (N_13952,N_6294,N_12220);
xnor U13953 (N_13953,N_9942,N_6666);
xor U13954 (N_13954,N_12376,N_10247);
or U13955 (N_13955,N_11534,N_11180);
xnor U13956 (N_13956,N_7678,N_11278);
and U13957 (N_13957,N_12414,N_8454);
or U13958 (N_13958,N_8561,N_8773);
nor U13959 (N_13959,N_11360,N_9408);
nand U13960 (N_13960,N_6706,N_6431);
nand U13961 (N_13961,N_11547,N_12385);
nand U13962 (N_13962,N_7373,N_10575);
nand U13963 (N_13963,N_8372,N_9057);
and U13964 (N_13964,N_9069,N_7024);
or U13965 (N_13965,N_11182,N_6717);
or U13966 (N_13966,N_10981,N_12118);
nand U13967 (N_13967,N_12081,N_11637);
and U13968 (N_13968,N_6880,N_6647);
or U13969 (N_13969,N_6930,N_12036);
nand U13970 (N_13970,N_9969,N_7338);
and U13971 (N_13971,N_8147,N_8103);
or U13972 (N_13972,N_9091,N_8604);
xnor U13973 (N_13973,N_8415,N_9714);
nor U13974 (N_13974,N_7151,N_11012);
nor U13975 (N_13975,N_7334,N_11529);
nand U13976 (N_13976,N_9058,N_6745);
and U13977 (N_13977,N_11838,N_9141);
and U13978 (N_13978,N_10975,N_11571);
or U13979 (N_13979,N_10366,N_8255);
nor U13980 (N_13980,N_7446,N_10232);
or U13981 (N_13981,N_10185,N_7425);
nor U13982 (N_13982,N_7054,N_11756);
or U13983 (N_13983,N_9316,N_10859);
or U13984 (N_13984,N_8054,N_7001);
or U13985 (N_13985,N_9939,N_8907);
or U13986 (N_13986,N_7751,N_6306);
or U13987 (N_13987,N_11264,N_9643);
and U13988 (N_13988,N_11121,N_8978);
nor U13989 (N_13989,N_12483,N_6423);
nor U13990 (N_13990,N_12447,N_6609);
nand U13991 (N_13991,N_9671,N_8188);
xnor U13992 (N_13992,N_9422,N_8041);
and U13993 (N_13993,N_6345,N_10655);
nand U13994 (N_13994,N_10714,N_8117);
nand U13995 (N_13995,N_12444,N_8662);
or U13996 (N_13996,N_11805,N_7692);
or U13997 (N_13997,N_12074,N_6644);
or U13998 (N_13998,N_6396,N_9777);
nor U13999 (N_13999,N_7629,N_9520);
and U14000 (N_14000,N_6816,N_12068);
nand U14001 (N_14001,N_11916,N_7220);
or U14002 (N_14002,N_8279,N_11599);
and U14003 (N_14003,N_7460,N_11519);
nor U14004 (N_14004,N_7330,N_11333);
and U14005 (N_14005,N_10121,N_10279);
nand U14006 (N_14006,N_11052,N_9220);
nor U14007 (N_14007,N_11915,N_9119);
nand U14008 (N_14008,N_7070,N_11085);
nor U14009 (N_14009,N_7708,N_7973);
nand U14010 (N_14010,N_11978,N_11729);
nand U14011 (N_14011,N_8370,N_7423);
and U14012 (N_14012,N_10676,N_7281);
or U14013 (N_14013,N_11228,N_8530);
and U14014 (N_14014,N_11783,N_11486);
nor U14015 (N_14015,N_11525,N_7920);
xor U14016 (N_14016,N_8099,N_6363);
and U14017 (N_14017,N_9326,N_8029);
or U14018 (N_14018,N_9246,N_11354);
nor U14019 (N_14019,N_8642,N_11995);
nand U14020 (N_14020,N_11509,N_10772);
nand U14021 (N_14021,N_8360,N_8150);
nor U14022 (N_14022,N_10519,N_9380);
nor U14023 (N_14023,N_9752,N_9902);
or U14024 (N_14024,N_8311,N_6556);
and U14025 (N_14025,N_7323,N_12059);
or U14026 (N_14026,N_10742,N_8259);
or U14027 (N_14027,N_6863,N_10864);
nand U14028 (N_14028,N_10183,N_7506);
xnor U14029 (N_14029,N_8348,N_8320);
or U14030 (N_14030,N_10318,N_9953);
nor U14031 (N_14031,N_10336,N_6483);
nand U14032 (N_14032,N_10691,N_9849);
and U14033 (N_14033,N_9586,N_7276);
nor U14034 (N_14034,N_10041,N_12169);
or U14035 (N_14035,N_6315,N_11524);
nor U14036 (N_14036,N_10722,N_6332);
or U14037 (N_14037,N_11887,N_8069);
xnor U14038 (N_14038,N_10406,N_8397);
or U14039 (N_14039,N_8727,N_7705);
nand U14040 (N_14040,N_7349,N_10170);
xnor U14041 (N_14041,N_7036,N_10367);
nand U14042 (N_14042,N_8205,N_7797);
xor U14043 (N_14043,N_12216,N_6412);
or U14044 (N_14044,N_11856,N_11020);
xnor U14045 (N_14045,N_11844,N_8042);
nor U14046 (N_14046,N_11485,N_8469);
and U14047 (N_14047,N_7582,N_10463);
or U14048 (N_14048,N_9711,N_12128);
nand U14049 (N_14049,N_11959,N_12005);
or U14050 (N_14050,N_6982,N_8374);
nand U14051 (N_14051,N_10114,N_12328);
nand U14052 (N_14052,N_12149,N_10416);
nand U14053 (N_14053,N_7632,N_8287);
nand U14054 (N_14054,N_9243,N_11577);
or U14055 (N_14055,N_9203,N_11775);
xnor U14056 (N_14056,N_8995,N_12403);
and U14057 (N_14057,N_12351,N_10497);
nand U14058 (N_14058,N_11049,N_10995);
nand U14059 (N_14059,N_6301,N_10223);
xor U14060 (N_14060,N_6350,N_11143);
nand U14061 (N_14061,N_6970,N_10636);
xor U14062 (N_14062,N_6347,N_6360);
nand U14063 (N_14063,N_9754,N_7291);
and U14064 (N_14064,N_8228,N_10720);
nand U14065 (N_14065,N_9247,N_11083);
nand U14066 (N_14066,N_10565,N_11047);
or U14067 (N_14067,N_10358,N_9747);
and U14068 (N_14068,N_9929,N_8085);
and U14069 (N_14069,N_7226,N_6451);
nand U14070 (N_14070,N_8829,N_7937);
nand U14071 (N_14071,N_11903,N_10064);
xnor U14072 (N_14072,N_9664,N_7925);
nor U14073 (N_14073,N_6305,N_6834);
nor U14074 (N_14074,N_9206,N_7429);
or U14075 (N_14075,N_9826,N_11760);
nor U14076 (N_14076,N_11522,N_8484);
nor U14077 (N_14077,N_10451,N_9884);
nand U14078 (N_14078,N_8953,N_9390);
nand U14079 (N_14079,N_11138,N_11404);
and U14080 (N_14080,N_9877,N_9809);
and U14081 (N_14081,N_6634,N_6491);
nand U14082 (N_14082,N_7539,N_10351);
or U14083 (N_14083,N_8290,N_11240);
nand U14084 (N_14084,N_7728,N_8378);
nand U14085 (N_14085,N_6329,N_7697);
or U14086 (N_14086,N_10385,N_9257);
or U14087 (N_14087,N_7642,N_9075);
nor U14088 (N_14088,N_7799,N_6841);
or U14089 (N_14089,N_10227,N_12314);
or U14090 (N_14090,N_6757,N_8700);
nor U14091 (N_14091,N_12324,N_11190);
and U14092 (N_14092,N_10004,N_9890);
or U14093 (N_14093,N_11082,N_6560);
and U14094 (N_14094,N_11445,N_12274);
or U14095 (N_14095,N_10136,N_12154);
and U14096 (N_14096,N_9213,N_9782);
and U14097 (N_14097,N_11814,N_8086);
nor U14098 (N_14098,N_10659,N_10548);
or U14099 (N_14099,N_6860,N_8616);
xnor U14100 (N_14100,N_8276,N_8999);
xnor U14101 (N_14101,N_8486,N_10252);
nor U14102 (N_14102,N_7943,N_6335);
nand U14103 (N_14103,N_7433,N_7357);
and U14104 (N_14104,N_8741,N_9763);
nand U14105 (N_14105,N_10391,N_7964);
nor U14106 (N_14106,N_9015,N_8569);
nand U14107 (N_14107,N_8897,N_6840);
nor U14108 (N_14108,N_11472,N_7081);
or U14109 (N_14109,N_10218,N_11350);
nand U14110 (N_14110,N_9564,N_9871);
and U14111 (N_14111,N_10595,N_7163);
nand U14112 (N_14112,N_11473,N_6453);
or U14113 (N_14113,N_8401,N_6995);
nor U14114 (N_14114,N_8806,N_12211);
and U14115 (N_14115,N_9770,N_9666);
and U14116 (N_14116,N_9766,N_11453);
nand U14117 (N_14117,N_10201,N_9233);
and U14118 (N_14118,N_11048,N_12357);
and U14119 (N_14119,N_6369,N_8403);
nand U14120 (N_14120,N_7910,N_10898);
or U14121 (N_14121,N_9388,N_6489);
nand U14122 (N_14122,N_11734,N_8132);
or U14123 (N_14123,N_9707,N_11669);
and U14124 (N_14124,N_8870,N_10719);
nand U14125 (N_14125,N_6533,N_7576);
nor U14126 (N_14126,N_6783,N_11331);
nand U14127 (N_14127,N_11405,N_6554);
and U14128 (N_14128,N_8963,N_6488);
or U14129 (N_14129,N_9379,N_9218);
nand U14130 (N_14130,N_11949,N_9533);
or U14131 (N_14131,N_9337,N_6590);
nor U14132 (N_14132,N_7154,N_11641);
and U14133 (N_14133,N_7006,N_10687);
nor U14134 (N_14134,N_9638,N_9298);
and U14135 (N_14135,N_11726,N_7375);
nand U14136 (N_14136,N_10081,N_11506);
nand U14137 (N_14137,N_11609,N_7287);
and U14138 (N_14138,N_8392,N_9631);
nand U14139 (N_14139,N_12014,N_12330);
and U14140 (N_14140,N_10501,N_12346);
and U14141 (N_14141,N_9850,N_9932);
nor U14142 (N_14142,N_11697,N_6954);
or U14143 (N_14143,N_9657,N_11452);
and U14144 (N_14144,N_9131,N_9352);
nor U14145 (N_14145,N_11259,N_9591);
xor U14146 (N_14146,N_10240,N_8450);
or U14147 (N_14147,N_11897,N_9128);
nand U14148 (N_14148,N_10278,N_8015);
or U14149 (N_14149,N_11026,N_10264);
nor U14150 (N_14150,N_10360,N_11257);
nor U14151 (N_14151,N_8899,N_11286);
or U14152 (N_14152,N_7386,N_10712);
nor U14153 (N_14153,N_7039,N_9874);
xnor U14154 (N_14154,N_6401,N_6905);
nor U14155 (N_14155,N_6798,N_12142);
and U14156 (N_14156,N_7679,N_11402);
and U14157 (N_14157,N_12382,N_9968);
xnor U14158 (N_14158,N_10925,N_9115);
nor U14159 (N_14159,N_12366,N_10258);
xnor U14160 (N_14160,N_10514,N_10612);
and U14161 (N_14161,N_10500,N_11184);
nand U14162 (N_14162,N_12427,N_11428);
nand U14163 (N_14163,N_6835,N_6958);
and U14164 (N_14164,N_8402,N_11603);
nand U14165 (N_14165,N_7963,N_11920);
xnor U14166 (N_14166,N_6966,N_9507);
or U14167 (N_14167,N_11988,N_8312);
or U14168 (N_14168,N_11639,N_11382);
nor U14169 (N_14169,N_8110,N_12203);
and U14170 (N_14170,N_8047,N_8793);
nand U14171 (N_14171,N_10056,N_8534);
or U14172 (N_14172,N_9404,N_9662);
nor U14173 (N_14173,N_8921,N_10837);
nand U14174 (N_14174,N_7275,N_7974);
xnor U14175 (N_14175,N_8008,N_11969);
or U14176 (N_14176,N_11284,N_8542);
xor U14177 (N_14177,N_11489,N_11929);
or U14178 (N_14178,N_9925,N_10444);
nor U14179 (N_14179,N_10036,N_11217);
nand U14180 (N_14180,N_9481,N_6851);
or U14181 (N_14181,N_9294,N_10502);
and U14182 (N_14182,N_10345,N_11176);
xnor U14183 (N_14183,N_7120,N_11984);
nand U14184 (N_14184,N_7214,N_10473);
and U14185 (N_14185,N_8362,N_8574);
nor U14186 (N_14186,N_8557,N_8643);
xnor U14187 (N_14187,N_9207,N_10395);
or U14188 (N_14188,N_6314,N_8230);
nand U14189 (N_14189,N_11225,N_9636);
nor U14190 (N_14190,N_10674,N_9216);
or U14191 (N_14191,N_9736,N_6639);
nor U14192 (N_14192,N_10220,N_8661);
nor U14193 (N_14193,N_10315,N_9353);
nand U14194 (N_14194,N_9073,N_11337);
nand U14195 (N_14195,N_11433,N_11448);
nand U14196 (N_14196,N_7809,N_8246);
nor U14197 (N_14197,N_12318,N_10652);
nand U14198 (N_14198,N_9489,N_8555);
nor U14199 (N_14199,N_8020,N_9105);
nor U14200 (N_14200,N_8606,N_8483);
nor U14201 (N_14201,N_9398,N_7011);
or U14202 (N_14202,N_10851,N_6399);
and U14203 (N_14203,N_6867,N_8384);
and U14204 (N_14204,N_7091,N_10934);
and U14205 (N_14205,N_10930,N_9741);
xnor U14206 (N_14206,N_10766,N_6579);
nand U14207 (N_14207,N_11699,N_8247);
nor U14208 (N_14208,N_8955,N_7552);
or U14209 (N_14209,N_6518,N_11343);
or U14210 (N_14210,N_9313,N_6501);
nor U14211 (N_14211,N_8404,N_9559);
and U14212 (N_14212,N_10496,N_9949);
or U14213 (N_14213,N_10092,N_9425);
nor U14214 (N_14214,N_11444,N_8163);
or U14215 (N_14215,N_10397,N_8628);
nand U14216 (N_14216,N_7967,N_7696);
nor U14217 (N_14217,N_8848,N_8462);
nand U14218 (N_14218,N_10835,N_7374);
xor U14219 (N_14219,N_7047,N_9106);
nand U14220 (N_14220,N_8319,N_9116);
and U14221 (N_14221,N_12286,N_10665);
and U14222 (N_14222,N_10068,N_7414);
and U14223 (N_14223,N_8369,N_10591);
and U14224 (N_14224,N_8010,N_11580);
nor U14225 (N_14225,N_9516,N_7741);
or U14226 (N_14226,N_12214,N_11282);
nor U14227 (N_14227,N_7701,N_11770);
or U14228 (N_14228,N_10656,N_10006);
nor U14229 (N_14229,N_8938,N_7821);
or U14230 (N_14230,N_8381,N_9975);
or U14231 (N_14231,N_11430,N_11961);
nor U14232 (N_14232,N_9509,N_10626);
and U14233 (N_14233,N_9724,N_11966);
nand U14234 (N_14234,N_10820,N_12432);
nand U14235 (N_14235,N_10199,N_7067);
or U14236 (N_14236,N_10635,N_11352);
nand U14237 (N_14237,N_11139,N_10355);
or U14238 (N_14238,N_11614,N_11260);
nor U14239 (N_14239,N_7003,N_12312);
or U14240 (N_14240,N_8673,N_11568);
or U14241 (N_14241,N_12050,N_9279);
nor U14242 (N_14242,N_11306,N_12192);
nand U14243 (N_14243,N_7661,N_6549);
nor U14244 (N_14244,N_10132,N_7236);
or U14245 (N_14245,N_11564,N_8724);
and U14246 (N_14246,N_11821,N_8626);
nand U14247 (N_14247,N_7211,N_8567);
nor U14248 (N_14248,N_7434,N_11779);
nand U14249 (N_14249,N_8668,N_8025);
nor U14250 (N_14250,N_8622,N_7759);
and U14251 (N_14251,N_12132,N_12104);
xor U14252 (N_14252,N_7754,N_11114);
and U14253 (N_14253,N_10080,N_11250);
nand U14254 (N_14254,N_9297,N_7894);
or U14255 (N_14255,N_10048,N_11859);
nand U14256 (N_14256,N_9077,N_6487);
or U14257 (N_14257,N_8764,N_7575);
nor U14258 (N_14258,N_12076,N_10804);
and U14259 (N_14259,N_8922,N_7530);
nand U14260 (N_14260,N_8084,N_9056);
and U14261 (N_14261,N_8782,N_8766);
or U14262 (N_14262,N_9500,N_10504);
nor U14263 (N_14263,N_7843,N_6460);
nor U14264 (N_14264,N_8763,N_9772);
and U14265 (N_14265,N_11313,N_6264);
or U14266 (N_14266,N_12492,N_9743);
or U14267 (N_14267,N_7946,N_7735);
and U14268 (N_14268,N_11728,N_7895);
or U14269 (N_14269,N_12412,N_11201);
nor U14270 (N_14270,N_8269,N_10526);
nor U14271 (N_14271,N_10069,N_7210);
nand U14272 (N_14272,N_9013,N_6400);
and U14273 (N_14273,N_10248,N_7083);
nor U14274 (N_14274,N_8666,N_11504);
or U14275 (N_14275,N_6951,N_7371);
nand U14276 (N_14276,N_10781,N_7034);
nor U14277 (N_14277,N_9225,N_8364);
and U14278 (N_14278,N_10839,N_8511);
and U14279 (N_14279,N_7995,N_11907);
nor U14280 (N_14280,N_9132,N_12180);
and U14281 (N_14281,N_10970,N_7930);
and U14282 (N_14282,N_9835,N_6869);
nand U14283 (N_14283,N_11205,N_10328);
nand U14284 (N_14284,N_10829,N_12148);
or U14285 (N_14285,N_6654,N_8602);
nand U14286 (N_14286,N_10731,N_8407);
and U14287 (N_14287,N_10707,N_10120);
nand U14288 (N_14288,N_11880,N_7510);
nor U14289 (N_14289,N_11651,N_9336);
nand U14290 (N_14290,N_9750,N_12099);
nor U14291 (N_14291,N_11868,N_7737);
nor U14292 (N_14292,N_8321,N_6944);
or U14293 (N_14293,N_6534,N_11892);
or U14294 (N_14294,N_10256,N_7458);
and U14295 (N_14295,N_11786,N_8961);
and U14296 (N_14296,N_6507,N_11704);
or U14297 (N_14297,N_9079,N_11815);
or U14298 (N_14298,N_10377,N_11543);
or U14299 (N_14299,N_11740,N_11407);
or U14300 (N_14300,N_9347,N_6825);
or U14301 (N_14301,N_6495,N_10671);
nor U14302 (N_14302,N_9214,N_9986);
nand U14303 (N_14303,N_7328,N_6719);
xor U14304 (N_14304,N_8245,N_7586);
nor U14305 (N_14305,N_11852,N_12279);
and U14306 (N_14306,N_7445,N_7755);
and U14307 (N_14307,N_8704,N_8613);
and U14308 (N_14308,N_11825,N_9935);
nand U14309 (N_14309,N_11122,N_11055);
and U14310 (N_14310,N_6871,N_7322);
and U14311 (N_14311,N_11065,N_11462);
nor U14312 (N_14312,N_11375,N_12315);
and U14313 (N_14313,N_8177,N_9136);
nand U14314 (N_14314,N_12300,N_6280);
or U14315 (N_14315,N_9619,N_11090);
or U14316 (N_14316,N_11076,N_7331);
nor U14317 (N_14317,N_11078,N_6922);
nand U14318 (N_14318,N_7289,N_12280);
and U14319 (N_14319,N_9001,N_9995);
or U14320 (N_14320,N_9629,N_8859);
xnor U14321 (N_14321,N_8425,N_8619);
and U14322 (N_14322,N_10283,N_8253);
nor U14323 (N_14323,N_6614,N_6650);
and U14324 (N_14324,N_8440,N_6434);
nand U14325 (N_14325,N_11276,N_6503);
and U14326 (N_14326,N_8631,N_6411);
nor U14327 (N_14327,N_9938,N_6896);
nor U14328 (N_14328,N_8964,N_9185);
or U14329 (N_14329,N_8067,N_12425);
or U14330 (N_14330,N_11013,N_7695);
and U14331 (N_14331,N_9532,N_7172);
nor U14332 (N_14332,N_12332,N_11097);
or U14333 (N_14333,N_11782,N_7444);
nand U14334 (N_14334,N_6799,N_11771);
nand U14335 (N_14335,N_12446,N_6805);
and U14336 (N_14336,N_9182,N_10051);
nand U14337 (N_14337,N_7878,N_8847);
nor U14338 (N_14338,N_9627,N_8719);
or U14339 (N_14339,N_8816,N_6406);
xnor U14340 (N_14340,N_12150,N_7115);
nor U14341 (N_14341,N_6681,N_9980);
nand U14342 (N_14342,N_10910,N_8924);
nor U14343 (N_14343,N_11544,N_9011);
nand U14344 (N_14344,N_7527,N_11330);
and U14345 (N_14345,N_11884,N_8203);
nor U14346 (N_14346,N_6443,N_10104);
and U14347 (N_14347,N_10302,N_6520);
xnor U14348 (N_14348,N_8153,N_11422);
nor U14349 (N_14349,N_6586,N_12072);
nand U14350 (N_14350,N_9599,N_12299);
and U14351 (N_14351,N_9485,N_9993);
or U14352 (N_14352,N_11939,N_10245);
nand U14353 (N_14353,N_6265,N_10909);
nand U14354 (N_14354,N_6649,N_8726);
nor U14355 (N_14355,N_7223,N_8757);
and U14356 (N_14356,N_12161,N_8272);
xor U14357 (N_14357,N_9814,N_10159);
or U14358 (N_14358,N_11611,N_6370);
and U14359 (N_14359,N_12208,N_9340);
nand U14360 (N_14360,N_7382,N_9389);
or U14361 (N_14361,N_12268,N_11274);
nor U14362 (N_14362,N_7239,N_9253);
xnor U14363 (N_14363,N_8797,N_11724);
xor U14364 (N_14364,N_9268,N_8548);
nor U14365 (N_14365,N_11230,N_10380);
nand U14366 (N_14366,N_9474,N_8033);
or U14367 (N_14367,N_10013,N_7503);
xnor U14368 (N_14368,N_12304,N_12400);
xor U14369 (N_14369,N_10873,N_7842);
and U14370 (N_14370,N_10334,N_7660);
or U14371 (N_14371,N_6708,N_10517);
nor U14372 (N_14372,N_12057,N_12428);
nand U14373 (N_14373,N_9495,N_12242);
nand U14374 (N_14374,N_7141,N_9221);
nand U14375 (N_14375,N_8379,N_10432);
nand U14376 (N_14376,N_11191,N_12455);
nand U14377 (N_14377,N_9263,N_9122);
or U14378 (N_14378,N_6807,N_6326);
and U14379 (N_14379,N_11701,N_10404);
and U14380 (N_14380,N_8594,N_7900);
nand U14381 (N_14381,N_7643,N_10130);
and U14382 (N_14382,N_11752,N_12205);
and U14383 (N_14383,N_10011,N_11548);
nand U14384 (N_14384,N_8532,N_6746);
and U14385 (N_14385,N_6612,N_6349);
nor U14386 (N_14386,N_8833,N_10014);
or U14387 (N_14387,N_11423,N_7590);
xor U14388 (N_14388,N_8498,N_10623);
xor U14389 (N_14389,N_9937,N_6542);
or U14390 (N_14390,N_8136,N_7903);
and U14391 (N_14391,N_9916,N_7150);
or U14392 (N_14392,N_10399,N_9397);
and U14393 (N_14393,N_6788,N_7090);
and U14394 (N_14394,N_7819,N_10871);
nand U14395 (N_14395,N_8315,N_6615);
nor U14396 (N_14396,N_7896,N_6935);
and U14397 (N_14397,N_10755,N_6267);
or U14398 (N_14398,N_8051,N_7655);
nor U14399 (N_14399,N_10761,N_10866);
xnor U14400 (N_14400,N_12215,N_10653);
and U14401 (N_14401,N_11235,N_9482);
and U14402 (N_14402,N_12002,N_12431);
or U14403 (N_14403,N_11962,N_9311);
and U14404 (N_14404,N_7347,N_9739);
and U14405 (N_14405,N_11766,N_10740);
nand U14406 (N_14406,N_12032,N_11467);
nor U14407 (N_14407,N_11002,N_9475);
nand U14408 (N_14408,N_11942,N_9018);
nor U14409 (N_14409,N_8346,N_9513);
nand U14410 (N_14410,N_12116,N_7638);
xnor U14411 (N_14411,N_7597,N_6619);
nor U14412 (N_14412,N_10625,N_11803);
nor U14413 (N_14413,N_12307,N_12407);
or U14414 (N_14414,N_8133,N_7419);
xnor U14415 (N_14415,N_8990,N_10047);
nand U14416 (N_14416,N_7026,N_8856);
or U14417 (N_14417,N_8185,N_10528);
nor U14418 (N_14418,N_12340,N_9165);
nand U14419 (N_14419,N_9235,N_9720);
and U14420 (N_14420,N_7004,N_9796);
xor U14421 (N_14421,N_12379,N_10800);
and U14422 (N_14422,N_11682,N_11057);
nor U14423 (N_14423,N_10348,N_8323);
or U14424 (N_14424,N_6635,N_11585);
nor U14425 (N_14425,N_10310,N_8049);
or U14426 (N_14426,N_9249,N_9043);
and U14427 (N_14427,N_9450,N_6832);
nor U14428 (N_14428,N_8291,N_8824);
nor U14429 (N_14429,N_9618,N_8400);
and U14430 (N_14430,N_10523,N_12239);
nor U14431 (N_14431,N_8313,N_12143);
xnor U14432 (N_14432,N_11608,N_7396);
and U14433 (N_14433,N_7348,N_11174);
or U14434 (N_14434,N_7674,N_12430);
nor U14435 (N_14435,N_8057,N_9608);
nand U14436 (N_14436,N_6468,N_10530);
nor U14437 (N_14437,N_10118,N_10756);
nor U14438 (N_14438,N_7035,N_10784);
or U14439 (N_14439,N_12006,N_8477);
xnor U14440 (N_14440,N_11894,N_11702);
nand U14441 (N_14441,N_9912,N_11874);
or U14442 (N_14442,N_9523,N_10171);
nand U14443 (N_14443,N_10850,N_8036);
xor U14444 (N_14444,N_10208,N_9675);
nand U14445 (N_14445,N_8260,N_11366);
nand U14446 (N_14446,N_7381,N_11110);
nor U14447 (N_14447,N_9061,N_10375);
or U14448 (N_14448,N_6672,N_11627);
xor U14449 (N_14449,N_7367,N_8601);
xor U14450 (N_14450,N_11383,N_6792);
or U14451 (N_14451,N_6271,N_6251);
nand U14452 (N_14452,N_12134,N_8125);
and U14453 (N_14453,N_12089,N_7467);
and U14454 (N_14454,N_11629,N_11558);
nor U14455 (N_14455,N_6960,N_6795);
nand U14456 (N_14456,N_8886,N_11879);
nand U14457 (N_14457,N_7399,N_9427);
nand U14458 (N_14458,N_9346,N_9779);
and U14459 (N_14459,N_7677,N_12209);
or U14460 (N_14460,N_9471,N_10268);
nand U14461 (N_14461,N_12254,N_10079);
or U14462 (N_14462,N_8930,N_12434);
nor U14463 (N_14463,N_6528,N_8553);
and U14464 (N_14464,N_6956,N_9370);
nor U14465 (N_14465,N_8075,N_11862);
nand U14466 (N_14466,N_11882,N_7863);
nand U14467 (N_14467,N_12202,N_10324);
or U14468 (N_14468,N_11373,N_9138);
and U14469 (N_14469,N_9819,N_11458);
or U14470 (N_14470,N_6394,N_8473);
xnor U14471 (N_14471,N_7486,N_10323);
nand U14472 (N_14472,N_6470,N_9113);
and U14473 (N_14473,N_10921,N_10280);
nand U14474 (N_14474,N_8551,N_7736);
and U14475 (N_14475,N_10110,N_8968);
nor U14476 (N_14476,N_12171,N_6529);
xor U14477 (N_14477,N_10897,N_11886);
nand U14478 (N_14478,N_10709,N_7215);
and U14479 (N_14479,N_6866,N_10533);
nand U14480 (N_14480,N_8262,N_8258);
nand U14481 (N_14481,N_11403,N_11739);
and U14482 (N_14482,N_7384,N_11332);
xnor U14483 (N_14483,N_9053,N_6390);
and U14484 (N_14484,N_6742,N_8517);
nor U14485 (N_14485,N_6325,N_9757);
nor U14486 (N_14486,N_9118,N_8249);
or U14487 (N_14487,N_10179,N_10300);
and U14488 (N_14488,N_9364,N_9773);
and U14489 (N_14489,N_9320,N_11142);
and U14490 (N_14490,N_6686,N_8123);
or U14491 (N_14491,N_10176,N_7791);
and U14492 (N_14492,N_9981,N_7489);
nand U14493 (N_14493,N_8333,N_8821);
nand U14494 (N_14494,N_9103,N_7633);
or U14495 (N_14495,N_6618,N_10212);
nand U14496 (N_14496,N_9129,N_11848);
nor U14497 (N_14497,N_7145,N_11590);
and U14498 (N_14498,N_9040,N_6711);
nor U14499 (N_14499,N_11292,N_6874);
or U14500 (N_14500,N_11146,N_7807);
and U14501 (N_14501,N_7561,N_10748);
nor U14502 (N_14502,N_7244,N_10522);
nor U14503 (N_14503,N_10723,N_9227);
nand U14504 (N_14504,N_8340,N_6891);
and U14505 (N_14505,N_8769,N_9002);
nor U14506 (N_14506,N_9906,N_8792);
nor U14507 (N_14507,N_7513,N_9310);
nor U14508 (N_14508,N_7152,N_9767);
nand U14509 (N_14509,N_8437,N_10816);
xnor U14510 (N_14510,N_9467,N_8295);
nand U14511 (N_14511,N_6872,N_11381);
and U14512 (N_14512,N_7760,N_11216);
nand U14513 (N_14513,N_7144,N_6611);
nor U14514 (N_14514,N_11232,N_8636);
nand U14515 (N_14515,N_10641,N_8538);
xnor U14516 (N_14516,N_6596,N_11498);
and U14517 (N_14517,N_6740,N_9114);
and U14518 (N_14518,N_11132,N_11940);
xor U14519 (N_14519,N_12418,N_10470);
or U14520 (N_14520,N_7566,N_7123);
and U14521 (N_14521,N_9280,N_11363);
xnor U14522 (N_14522,N_11826,N_6571);
nand U14523 (N_14523,N_10578,N_9147);
nand U14524 (N_14524,N_7727,N_8206);
nand U14525 (N_14525,N_10204,N_7102);
xnor U14526 (N_14526,N_9875,N_8934);
and U14527 (N_14527,N_12033,N_11068);
nor U14528 (N_14528,N_7524,N_10602);
nand U14529 (N_14529,N_8448,N_10680);
or U14530 (N_14530,N_10198,N_8579);
or U14531 (N_14531,N_11371,N_6539);
or U14532 (N_14532,N_11910,N_7716);
and U14533 (N_14533,N_7778,N_11549);
nor U14534 (N_14534,N_10018,N_12029);
and U14535 (N_14535,N_10402,N_6580);
nand U14536 (N_14536,N_9806,N_9291);
and U14537 (N_14537,N_10058,N_8565);
nor U14538 (N_14538,N_11123,N_10259);
nor U14539 (N_14539,N_8687,N_11866);
nand U14540 (N_14540,N_6541,N_10715);
nand U14541 (N_14541,N_10364,N_8693);
nand U14542 (N_14542,N_11674,N_10394);
or U14543 (N_14543,N_9445,N_10681);
nand U14544 (N_14544,N_6536,N_11311);
xor U14545 (N_14545,N_9437,N_12235);
or U14546 (N_14546,N_8627,N_11913);
nand U14547 (N_14547,N_6289,N_11019);
nand U14548 (N_14548,N_9028,N_10990);
nor U14549 (N_14549,N_7370,N_10957);
nor U14550 (N_14550,N_10860,N_12250);
nor U14551 (N_14551,N_7413,N_7600);
nor U14552 (N_14552,N_9502,N_9800);
or U14553 (N_14553,N_9244,N_11581);
nor U14554 (N_14554,N_8476,N_8590);
and U14555 (N_14555,N_7405,N_8475);
and U14556 (N_14556,N_8116,N_10745);
nand U14557 (N_14557,N_10878,N_11755);
nand U14558 (N_14558,N_10762,N_8045);
nor U14559 (N_14559,N_8226,N_10912);
nor U14560 (N_14560,N_6793,N_9616);
nand U14561 (N_14561,N_6789,N_8873);
xnor U14562 (N_14562,N_10551,N_12409);
or U14563 (N_14563,N_8195,N_10808);
and U14564 (N_14564,N_8497,N_11542);
or U14565 (N_14565,N_8812,N_9792);
and U14566 (N_14566,N_10296,N_12087);
nor U14567 (N_14567,N_10244,N_8170);
xor U14568 (N_14568,N_9801,N_10329);
and U14569 (N_14569,N_9954,N_6802);
or U14570 (N_14570,N_10337,N_9248);
or U14571 (N_14571,N_7231,N_7639);
and U14572 (N_14572,N_8420,N_8690);
nand U14573 (N_14573,N_8777,N_8681);
or U14574 (N_14574,N_8329,N_8849);
nand U14575 (N_14575,N_6260,N_6677);
and U14576 (N_14576,N_6978,N_7688);
nand U14577 (N_14577,N_9175,N_7988);
or U14578 (N_14578,N_9055,N_12012);
or U14579 (N_14579,N_8422,N_7647);
or U14580 (N_14580,N_7385,N_11426);
nand U14581 (N_14581,N_12480,N_6782);
and U14582 (N_14582,N_9899,N_11022);
nor U14583 (N_14583,N_9530,N_7584);
nand U14584 (N_14584,N_8316,N_11418);
nor U14585 (N_14585,N_11999,N_8165);
or U14586 (N_14586,N_9014,N_11070);
nor U14587 (N_14587,N_9701,N_10601);
nor U14588 (N_14588,N_11018,N_11992);
xor U14589 (N_14589,N_11905,N_11928);
nor U14590 (N_14590,N_10790,N_12041);
nand U14591 (N_14591,N_6342,N_6377);
nand U14592 (N_14592,N_7073,N_8439);
xnor U14593 (N_14593,N_10673,N_7180);
or U14594 (N_14594,N_8264,N_11749);
and U14595 (N_14595,N_8711,N_11273);
nand U14596 (N_14596,N_7975,N_6441);
xnor U14597 (N_14597,N_10787,N_12141);
nor U14598 (N_14598,N_6781,N_8037);
nor U14599 (N_14599,N_10433,N_11926);
nor U14600 (N_14600,N_10658,N_12138);
or U14601 (N_14601,N_6786,N_6743);
and U14602 (N_14602,N_7686,N_7872);
nor U14603 (N_14603,N_7941,N_7715);
xnor U14604 (N_14604,N_9794,N_11161);
xnor U14605 (N_14605,N_11795,N_9019);
nor U14606 (N_14606,N_10525,N_6993);
or U14607 (N_14607,N_7709,N_11297);
xnor U14608 (N_14608,N_12079,N_8679);
and U14609 (N_14609,N_7773,N_6983);
or U14610 (N_14610,N_7866,N_8818);
or U14611 (N_14611,N_11345,N_6391);
nand U14612 (N_14612,N_8864,N_7005);
xnor U14613 (N_14613,N_11490,N_6753);
nand U14614 (N_14614,N_6684,N_10383);
xnor U14615 (N_14615,N_6508,N_9851);
and U14616 (N_14616,N_11275,N_8204);
nor U14617 (N_14617,N_8525,N_10559);
nor U14618 (N_14618,N_6806,N_10168);
and U14619 (N_14619,N_6664,N_10098);
or U14620 (N_14620,N_8787,N_10949);
and U14621 (N_14621,N_9704,N_8837);
nor U14622 (N_14622,N_8908,N_7682);
nor U14623 (N_14623,N_10534,N_7794);
xnor U14624 (N_14624,N_11846,N_10776);
nand U14625 (N_14625,N_9095,N_7829);
and U14626 (N_14626,N_9021,N_7166);
nand U14627 (N_14627,N_8592,N_8775);
or U14628 (N_14628,N_9349,N_12456);
or U14629 (N_14629,N_6975,N_8479);
and U14630 (N_14630,N_11985,N_10437);
nor U14631 (N_14631,N_8303,N_9565);
nor U14632 (N_14632,N_10253,N_9417);
nand U14633 (N_14633,N_8900,N_7653);
or U14634 (N_14634,N_7352,N_8786);
or U14635 (N_14635,N_9211,N_10542);
nor U14636 (N_14636,N_10173,N_9309);
nor U14637 (N_14637,N_7053,N_11851);
and U14638 (N_14638,N_11380,N_6333);
nor U14639 (N_14639,N_11303,N_8798);
and U14640 (N_14640,N_6359,N_12073);
or U14641 (N_14641,N_8003,N_11644);
nand U14642 (N_14642,N_8096,N_10799);
and U14643 (N_14643,N_6471,N_10203);
or U14644 (N_14644,N_6262,N_7962);
xnor U14645 (N_14645,N_10239,N_10099);
nand U14646 (N_14646,N_6748,N_11811);
nor U14647 (N_14647,N_12422,N_10449);
or U14648 (N_14648,N_11449,N_8647);
xor U14649 (N_14649,N_9653,N_7064);
nand U14650 (N_14650,N_6964,N_6540);
and U14651 (N_14651,N_9498,N_8927);
or U14652 (N_14652,N_9626,N_11717);
and U14653 (N_14653,N_8735,N_9988);
nand U14654 (N_14654,N_8669,N_12336);
nor U14655 (N_14655,N_8982,N_6379);
nand U14656 (N_14656,N_11833,N_9100);
nand U14657 (N_14657,N_11446,N_6558);
nand U14658 (N_14658,N_8144,N_7722);
nor U14659 (N_14659,N_10945,N_8942);
xor U14660 (N_14660,N_10825,N_7297);
nor U14661 (N_14661,N_12461,N_10738);
nand U14662 (N_14662,N_10801,N_10852);
nand U14663 (N_14663,N_8335,N_11036);
nand U14664 (N_14664,N_12172,N_12265);
or U14665 (N_14665,N_8919,N_10357);
nand U14666 (N_14666,N_11016,N_10457);
xnor U14667 (N_14667,N_7864,N_7393);
and U14668 (N_14668,N_9145,N_10067);
nand U14669 (N_14669,N_6531,N_11745);
or U14670 (N_14670,N_9838,N_10562);
or U14671 (N_14671,N_9928,N_7617);
and U14672 (N_14672,N_9677,N_9538);
nand U14673 (N_14673,N_10928,N_10148);
and U14674 (N_14674,N_6439,N_11796);
and U14675 (N_14675,N_7344,N_7170);
or U14676 (N_14676,N_7261,N_11661);
nor U14677 (N_14677,N_7031,N_10677);
or U14678 (N_14678,N_10539,N_6340);
and U14679 (N_14679,N_8452,N_11968);
xnor U14680 (N_14680,N_7854,N_10005);
xor U14681 (N_14681,N_11679,N_10554);
or U14682 (N_14682,N_10044,N_11801);
or U14683 (N_14683,N_10003,N_6680);
and U14684 (N_14684,N_12103,N_8386);
xor U14685 (N_14685,N_7443,N_10493);
nand U14686 (N_14686,N_11077,N_7092);
or U14687 (N_14687,N_11989,N_8223);
nand U14688 (N_14688,N_10046,N_8062);
nand U14689 (N_14689,N_6675,N_11406);
nand U14690 (N_14690,N_11716,N_6334);
or U14691 (N_14691,N_10887,N_11054);
nor U14692 (N_14692,N_8732,N_7763);
nand U14693 (N_14693,N_11620,N_12367);
nand U14694 (N_14694,N_11439,N_8352);
nor U14695 (N_14695,N_7100,N_6458);
nor U14696 (N_14696,N_7147,N_11058);
nand U14697 (N_14697,N_10511,N_10642);
nor U14698 (N_14698,N_9010,N_9700);
or U14699 (N_14699,N_9312,N_11912);
nand U14700 (N_14700,N_7432,N_12035);
nor U14701 (N_14701,N_6331,N_10622);
nor U14702 (N_14702,N_12378,N_6846);
nand U14703 (N_14703,N_8197,N_10701);
nor U14704 (N_14704,N_11372,N_8160);
or U14705 (N_14705,N_8194,N_10660);
nand U14706 (N_14706,N_9457,N_6952);
nor U14707 (N_14707,N_7710,N_9863);
nand U14708 (N_14708,N_9381,N_10543);
nand U14709 (N_14709,N_6801,N_10276);
xnor U14710 (N_14710,N_9462,N_10049);
nor U14711 (N_14711,N_9410,N_12370);
or U14712 (N_14712,N_8987,N_10396);
or U14713 (N_14713,N_11414,N_7502);
nor U14714 (N_14714,N_7889,N_11287);
or U14715 (N_14715,N_12296,N_9319);
or U14716 (N_14716,N_8071,N_8898);
nand U14717 (N_14717,N_10384,N_12469);
or U14718 (N_14718,N_6844,N_8801);
nand U14719 (N_14719,N_11819,N_11505);
and U14720 (N_14720,N_6494,N_8006);
nand U14721 (N_14721,N_11416,N_9815);
nand U14722 (N_14722,N_9356,N_12345);
or U14723 (N_14723,N_8127,N_9709);
nand U14724 (N_14724,N_7251,N_8843);
nand U14725 (N_14725,N_6552,N_11322);
and U14726 (N_14726,N_11447,N_6432);
and U14727 (N_14727,N_10974,N_11816);
nand U14728 (N_14728,N_8001,N_6604);
and U14729 (N_14729,N_6455,N_11818);
nand U14730 (N_14730,N_8545,N_7478);
nand U14731 (N_14731,N_8141,N_7983);
or U14732 (N_14732,N_9702,N_12356);
and U14733 (N_14733,N_11136,N_8956);
and U14734 (N_14734,N_7912,N_7628);
and U14735 (N_14735,N_9382,N_12045);
xnor U14736 (N_14736,N_9173,N_11434);
nand U14737 (N_14737,N_8063,N_7883);
nor U14738 (N_14738,N_9688,N_6601);
and U14739 (N_14739,N_7650,N_6683);
and U14740 (N_14740,N_8391,N_6433);
nand U14741 (N_14741,N_6302,N_10145);
nor U14742 (N_14742,N_9924,N_10486);
or U14743 (N_14743,N_8235,N_10105);
xor U14744 (N_14744,N_6921,N_6592);
or U14745 (N_14745,N_7171,N_12122);
nor U14746 (N_14746,N_8610,N_8657);
or U14747 (N_14747,N_11667,N_9314);
and U14748 (N_14748,N_10499,N_6667);
nor U14749 (N_14749,N_9965,N_6947);
nand U14750 (N_14750,N_10846,N_7841);
nor U14751 (N_14751,N_10917,N_8876);
nor U14752 (N_14752,N_10638,N_6422);
xor U14753 (N_14753,N_7670,N_8449);
and U14754 (N_14754,N_10629,N_7605);
or U14755 (N_14755,N_6859,N_6481);
nor U14756 (N_14756,N_10388,N_11305);
nor U14757 (N_14757,N_9494,N_7266);
nor U14758 (N_14758,N_8098,N_11598);
and U14759 (N_14759,N_11676,N_9205);
or U14760 (N_14760,N_9183,N_6598);
and U14761 (N_14761,N_7543,N_11904);
nand U14762 (N_14762,N_9974,N_10445);
or U14763 (N_14763,N_9444,N_9217);
or U14764 (N_14764,N_12170,N_10718);
nand U14765 (N_14765,N_9142,N_10583);
xor U14766 (N_14766,N_10465,N_7730);
or U14767 (N_14767,N_8024,N_6704);
nand U14768 (N_14768,N_10374,N_8399);
nor U14769 (N_14769,N_7607,N_7784);
or U14770 (N_14770,N_7169,N_9051);
nand U14771 (N_14771,N_10241,N_10151);
or U14772 (N_14772,N_7304,N_10210);
xor U14773 (N_14773,N_7130,N_7378);
or U14774 (N_14774,N_10647,N_7364);
nor U14775 (N_14775,N_9157,N_10684);
nor U14776 (N_14776,N_8267,N_6599);
or U14777 (N_14777,N_10958,N_12292);
or U14778 (N_14778,N_12206,N_7816);
nor U14779 (N_14779,N_9371,N_8241);
or U14780 (N_14780,N_12020,N_11218);
or U14781 (N_14781,N_7505,N_9703);
or U14782 (N_14782,N_10295,N_9317);
and U14783 (N_14783,N_11107,N_10902);
nand U14784 (N_14784,N_12114,N_9776);
and U14785 (N_14785,N_10895,N_8998);
nor U14786 (N_14786,N_9855,N_10001);
or U14787 (N_14787,N_9512,N_9277);
nor U14788 (N_14788,N_8122,N_11241);
or U14789 (N_14789,N_12288,N_10711);
xnor U14790 (N_14790,N_7882,N_9852);
and U14791 (N_14791,N_7040,N_10294);
nor U14792 (N_14792,N_10922,N_8499);
and U14793 (N_14793,N_6258,N_9031);
and U14794 (N_14794,N_9774,N_10490);
and U14795 (N_14795,N_8983,N_10103);
nor U14796 (N_14796,N_12410,N_11705);
nor U14797 (N_14797,N_6538,N_10634);
or U14798 (N_14798,N_11031,N_10867);
and U14799 (N_14799,N_8954,N_6847);
nor U14800 (N_14800,N_8718,N_8536);
or U14801 (N_14801,N_6973,N_7408);
or U14802 (N_14802,N_9686,N_10156);
nor U14803 (N_14803,N_10739,N_9414);
or U14804 (N_14804,N_7372,N_7630);
xnor U14805 (N_14805,N_7264,N_10368);
nor U14806 (N_14806,N_9551,N_7874);
nor U14807 (N_14807,N_8112,N_9885);
xor U14808 (N_14808,N_10561,N_8274);
nor U14809 (N_14809,N_8675,N_9447);
and U14810 (N_14810,N_6702,N_12365);
nand U14811 (N_14811,N_7768,N_6290);
or U14812 (N_14812,N_10143,N_10913);
or U14813 (N_14813,N_8518,N_9192);
nor U14814 (N_14814,N_11312,N_11496);
xnor U14815 (N_14815,N_7879,N_10510);
and U14816 (N_14816,N_8625,N_10305);
nand U14817 (N_14817,N_11079,N_9384);
nand U14818 (N_14818,N_8447,N_7950);
xnor U14819 (N_14819,N_8327,N_11703);
and U14820 (N_14820,N_12464,N_8178);
or U14821 (N_14821,N_10545,N_7044);
and U14822 (N_14822,N_9879,N_6839);
nor U14823 (N_14823,N_12158,N_6926);
or U14824 (N_14824,N_9749,N_7579);
nor U14825 (N_14825,N_7271,N_12321);
or U14826 (N_14826,N_9737,N_11579);
nor U14827 (N_14827,N_9374,N_6327);
nand U14828 (N_14828,N_7301,N_10225);
or U14829 (N_14829,N_8224,N_6849);
and U14830 (N_14830,N_11660,N_7767);
xor U14831 (N_14831,N_6473,N_11936);
nand U14832 (N_14832,N_10950,N_9070);
and U14833 (N_14833,N_7126,N_8691);
xnor U14834 (N_14834,N_12488,N_7885);
xor U14835 (N_14835,N_12443,N_10265);
nand U14836 (N_14836,N_10544,N_7792);
xnor U14837 (N_14837,N_9042,N_6295);
and U14838 (N_14838,N_6820,N_8238);
nand U14839 (N_14839,N_9228,N_8478);
and U14840 (N_14840,N_7972,N_9198);
nand U14841 (N_14841,N_10935,N_7480);
nor U14842 (N_14842,N_10973,N_10401);
and U14843 (N_14843,N_11516,N_7801);
or U14844 (N_14844,N_6299,N_7050);
nor U14845 (N_14845,N_10269,N_10590);
nor U14846 (N_14846,N_10381,N_7581);
xor U14847 (N_14847,N_6919,N_9107);
nor U14848 (N_14848,N_8966,N_7824);
or U14849 (N_14849,N_8559,N_9108);
nor U14850 (N_14850,N_8277,N_10237);
and U14851 (N_14851,N_9745,N_10810);
and U14852 (N_14852,N_8134,N_11021);
nand U14853 (N_14853,N_10020,N_6674);
nand U14854 (N_14854,N_9866,N_7595);
nand U14855 (N_14855,N_11714,N_10900);
or U14856 (N_14856,N_6779,N_9691);
or U14857 (N_14857,N_9391,N_7781);
or U14858 (N_14858,N_6525,N_7116);
or U14859 (N_14859,N_10400,N_10211);
nor U14860 (N_14860,N_6480,N_7095);
or U14861 (N_14861,N_8421,N_11595);
and U14862 (N_14862,N_7599,N_7992);
nor U14863 (N_14863,N_9199,N_10700);
nor U14864 (N_14864,N_6591,N_11638);
and U14865 (N_14865,N_6479,N_10274);
nor U14866 (N_14866,N_10234,N_8868);
nand U14867 (N_14867,N_6581,N_11829);
and U14868 (N_14868,N_10146,N_8293);
nand U14869 (N_14869,N_6961,N_8149);
or U14870 (N_14870,N_9508,N_11924);
and U14871 (N_14871,N_12207,N_9872);
and U14872 (N_14872,N_7415,N_10507);
and U14873 (N_14873,N_8734,N_10736);
nand U14874 (N_14874,N_11369,N_9148);
nand U14875 (N_14875,N_8958,N_7756);
xor U14876 (N_14876,N_10468,N_9126);
or U14877 (N_14877,N_10580,N_11164);
and U14878 (N_14878,N_6421,N_6796);
xor U14879 (N_14879,N_12163,N_11593);
and U14880 (N_14880,N_9271,N_7071);
or U14881 (N_14881,N_9189,N_9431);
or U14882 (N_14882,N_7229,N_8692);
and U14883 (N_14883,N_7033,N_12084);
or U14884 (N_14884,N_9383,N_8583);
nand U14885 (N_14885,N_6830,N_10150);
xor U14886 (N_14886,N_9600,N_8257);
nand U14887 (N_14887,N_11622,N_10685);
and U14888 (N_14888,N_8740,N_10750);
and U14889 (N_14889,N_6977,N_12377);
xnor U14890 (N_14890,N_6546,N_8944);
and U14891 (N_14891,N_11041,N_12486);
xnor U14892 (N_14892,N_6817,N_9648);
or U14893 (N_14893,N_9642,N_8665);
nor U14894 (N_14894,N_10785,N_8468);
nor U14895 (N_14895,N_8566,N_9290);
nor U14896 (N_14896,N_7554,N_8375);
and U14897 (N_14897,N_8516,N_6986);
nand U14898 (N_14898,N_6910,N_10916);
and U14899 (N_14899,N_11326,N_8181);
or U14900 (N_14900,N_7904,N_8114);
nor U14901 (N_14901,N_11633,N_7891);
and U14902 (N_14902,N_12364,N_6949);
or U14903 (N_14903,N_8428,N_8519);
xor U14904 (N_14904,N_12435,N_10040);
or U14905 (N_14905,N_10865,N_10703);
nor U14906 (N_14906,N_11474,N_9024);
and U14907 (N_14907,N_7646,N_7257);
xor U14908 (N_14908,N_10955,N_10557);
and U14909 (N_14909,N_9786,N_7296);
or U14910 (N_14910,N_10290,N_11692);
xnor U14911 (N_14911,N_11605,N_11937);
and U14912 (N_14912,N_6725,N_7412);
and U14913 (N_14913,N_8300,N_11680);
or U14914 (N_14914,N_6698,N_8461);
nand U14915 (N_14915,N_8709,N_9479);
nor U14916 (N_14916,N_8412,N_12027);
or U14917 (N_14917,N_7717,N_8828);
nand U14918 (N_14918,N_11743,N_10967);
nor U14919 (N_14919,N_11497,N_8973);
xor U14920 (N_14920,N_7199,N_12247);
or U14921 (N_14921,N_7188,N_8623);
nor U14922 (N_14922,N_6288,N_6416);
or U14923 (N_14923,N_10321,N_7707);
nand U14924 (N_14924,N_10757,N_10827);
nand U14925 (N_14925,N_7158,N_6291);
or U14926 (N_14926,N_9843,N_7339);
nand U14927 (N_14927,N_9553,N_7999);
and U14928 (N_14928,N_7977,N_10095);
and U14929 (N_14929,N_10097,N_10030);
or U14930 (N_14930,N_7454,N_7540);
nor U14931 (N_14931,N_6636,N_10427);
xor U14932 (N_14932,N_6282,N_7245);
and U14933 (N_14933,N_8239,N_12494);
or U14934 (N_14934,N_11424,N_10914);
or U14935 (N_14935,N_11828,N_8748);
and U14936 (N_14936,N_11733,N_6255);
or U14937 (N_14937,N_10116,N_7016);
and U14938 (N_14938,N_11712,N_10082);
or U14939 (N_14939,N_11528,N_8731);
nor U14940 (N_14940,N_7167,N_9825);
or U14941 (N_14941,N_11038,N_8034);
or U14942 (N_14942,N_9039,N_11839);
or U14943 (N_14943,N_9416,N_6991);
and U14944 (N_14944,N_12487,N_10062);
nand U14945 (N_14945,N_12399,N_9696);
nor U14946 (N_14946,N_10743,N_7849);
nand U14947 (N_14947,N_10229,N_10491);
or U14948 (N_14948,N_8940,N_11167);
nand U14949 (N_14949,N_8667,N_11213);
and U14950 (N_14950,N_11657,N_9162);
or U14951 (N_14951,N_8470,N_7193);
nand U14952 (N_14952,N_9089,N_9780);
or U14953 (N_14953,N_10689,N_11666);
and U14954 (N_14954,N_12090,N_10330);
nand U14955 (N_14955,N_6346,N_10708);
and U14956 (N_14956,N_7672,N_8959);
xor U14957 (N_14957,N_9208,N_8874);
and U14958 (N_14958,N_7881,N_11731);
nor U14959 (N_14959,N_12119,N_7598);
nor U14960 (N_14960,N_11435,N_10022);
or U14961 (N_14961,N_8240,N_9430);
nor U14962 (N_14962,N_10872,N_10664);
nand U14963 (N_14963,N_10108,N_9299);
nand U14964 (N_14964,N_8905,N_7507);
nor U14965 (N_14965,N_10314,N_6697);
nand U14966 (N_14966,N_8802,N_8760);
nand U14967 (N_14967,N_8923,N_9335);
and U14968 (N_14968,N_8166,N_7137);
xnor U14969 (N_14969,N_8850,N_11411);
nand U14970 (N_14970,N_7526,N_6530);
or U14971 (N_14971,N_7183,N_10777);
nand U14972 (N_14972,N_8501,N_6669);
nand U14973 (N_14973,N_8783,N_11014);
or U14974 (N_14974,N_9167,N_8038);
xor U14975 (N_14975,N_6679,N_9385);
and U14976 (N_14976,N_7453,N_9004);
or U14977 (N_14977,N_6485,N_8915);
and U14978 (N_14978,N_11621,N_9318);
nand U14979 (N_14979,N_10165,N_10518);
nor U14980 (N_14980,N_6676,N_8770);
and U14981 (N_14981,N_8685,N_10992);
nand U14982 (N_14982,N_11459,N_7899);
xnor U14983 (N_14983,N_7041,N_7608);
or U14984 (N_14984,N_9708,N_9936);
or U14985 (N_14985,N_7227,N_7046);
xnor U14986 (N_14986,N_9952,N_12056);
nand U14987 (N_14987,N_8121,N_6689);
nand U14988 (N_14988,N_11616,N_6456);
and U14989 (N_14989,N_10996,N_8443);
nand U14990 (N_14990,N_11640,N_8664);
nand U14991 (N_14991,N_11499,N_11266);
or U14992 (N_14992,N_8097,N_7606);
nor U14993 (N_14993,N_11247,N_11790);
xor U14994 (N_14994,N_9923,N_10713);
xor U14995 (N_14995,N_11207,N_8593);
xor U14996 (N_14996,N_8215,N_10841);
nand U14997 (N_14997,N_10573,N_12204);
and U14998 (N_14998,N_7121,N_9976);
nand U14999 (N_14999,N_9756,N_9281);
nand U15000 (N_15000,N_7938,N_12256);
nor U15001 (N_15001,N_6375,N_12309);
and U15002 (N_15002,N_11144,N_11347);
and U15003 (N_15003,N_8768,N_10233);
xnor U15004 (N_15004,N_6946,N_7476);
nand U15005 (N_15005,N_6854,N_7901);
and U15006 (N_15006,N_6897,N_11227);
and U15007 (N_15007,N_11256,N_6268);
xor U15008 (N_15008,N_11410,N_10765);
nor U15009 (N_15009,N_8263,N_7739);
nand U15010 (N_15010,N_8179,N_10311);
nand U15011 (N_15011,N_12497,N_9306);
nand U15012 (N_15012,N_9110,N_9692);
nand U15013 (N_15013,N_9840,N_8508);
nand U15014 (N_15014,N_8026,N_10905);
or U15015 (N_15015,N_6587,N_8079);
and U15016 (N_15016,N_9822,N_9409);
or U15017 (N_15017,N_12476,N_9109);
and U15018 (N_15018,N_11440,N_8108);
or U15019 (N_15019,N_10716,N_11841);
or U15020 (N_15020,N_7779,N_10553);
and U15021 (N_15021,N_6668,N_6382);
or U15022 (N_15022,N_7691,N_11727);
and U15023 (N_15023,N_12236,N_9315);
and U15024 (N_15024,N_7738,N_12083);
nor U15025 (N_15025,N_7596,N_9660);
nor U15026 (N_15026,N_10678,N_9161);
nor U15027 (N_15027,N_10581,N_10361);
nor U15028 (N_15028,N_8754,N_12126);
or U15029 (N_15029,N_12190,N_12452);
and U15030 (N_15030,N_9882,N_10855);
nor U15031 (N_15031,N_10469,N_9080);
or U15032 (N_15032,N_6450,N_11927);
nand U15033 (N_15033,N_8186,N_8061);
xnor U15034 (N_15034,N_10200,N_7103);
or U15035 (N_15035,N_7212,N_10527);
or U15036 (N_15036,N_11475,N_10734);
nand U15037 (N_15037,N_9753,N_9017);
nor U15038 (N_15038,N_6603,N_10836);
or U15039 (N_15039,N_11189,N_9387);
nand U15040 (N_15040,N_12004,N_7770);
xor U15041 (N_15041,N_11596,N_12421);
xnor U15042 (N_15042,N_11592,N_9477);
and U15043 (N_15043,N_11875,N_8345);
nor U15044 (N_15044,N_9421,N_10172);
nand U15045 (N_15045,N_11493,N_9670);
or U15046 (N_15046,N_11059,N_12478);
nor U15047 (N_15047,N_9594,N_8791);
xor U15048 (N_15048,N_8882,N_7206);
and U15049 (N_15049,N_10672,N_7788);
nor U15050 (N_15050,N_8544,N_11248);
nor U15051 (N_15051,N_7058,N_8490);
nand U15052 (N_15052,N_10662,N_12055);
and U15053 (N_15053,N_9350,N_8556);
or U15054 (N_15054,N_11429,N_12275);
nor U15055 (N_15055,N_8377,N_8266);
xor U15056 (N_15056,N_12295,N_7056);
nor U15057 (N_15057,N_11572,N_7702);
nor U15058 (N_15058,N_10157,N_7051);
nand U15059 (N_15059,N_10408,N_6424);
or U15060 (N_15060,N_7626,N_10184);
or U15061 (N_15061,N_11359,N_9446);
or U15062 (N_15062,N_12445,N_10415);
nor U15063 (N_15063,N_7218,N_8081);
or U15064 (N_15064,N_7455,N_7345);
xnor U15065 (N_15065,N_7888,N_9996);
and U15066 (N_15066,N_8466,N_9440);
nor U15067 (N_15067,N_9897,N_8862);
and U15068 (N_15068,N_9955,N_10568);
nand U15069 (N_15069,N_6521,N_6727);
xnor U15070 (N_15070,N_8863,N_8182);
and U15071 (N_15071,N_8502,N_10947);
nor U15072 (N_15072,N_7494,N_8019);
and U15073 (N_15073,N_7136,N_9005);
and U15074 (N_15074,N_12080,N_12338);
nand U15075 (N_15075,N_11784,N_10135);
nand U15076 (N_15076,N_11328,N_10096);
and U15077 (N_15077,N_9905,N_6296);
or U15078 (N_15078,N_7542,N_11344);
nand U15079 (N_15079,N_11062,N_8053);
and U15080 (N_15080,N_6662,N_6338);
or U15081 (N_15081,N_10471,N_9606);
or U15082 (N_15082,N_10007,N_12294);
nor U15083 (N_15083,N_7068,N_8347);
and U15084 (N_15084,N_9830,N_8229);
and U15085 (N_15085,N_11827,N_9407);
and U15086 (N_15086,N_6555,N_9592);
and U15087 (N_15087,N_10313,N_9983);
and U15088 (N_15088,N_12397,N_8887);
nor U15089 (N_15089,N_11194,N_6402);
nor U15090 (N_15090,N_11541,N_12196);
nor U15091 (N_15091,N_7418,N_7205);
nand U15092 (N_15092,N_10727,N_10729);
and U15093 (N_15093,N_7343,N_12181);
or U15094 (N_15094,N_10138,N_8572);
or U15095 (N_15095,N_11652,N_6505);
nor U15096 (N_15096,N_7280,N_8603);
nand U15097 (N_15097,N_9241,N_7465);
nand U15098 (N_15098,N_10061,N_8022);
and U15099 (N_15099,N_8242,N_11491);
nand U15100 (N_15100,N_9837,N_6467);
or U15101 (N_15101,N_11163,N_12374);
xnor U15102 (N_15102,N_6304,N_9665);
or U15103 (N_15103,N_11212,N_10251);
xnor U15104 (N_15104,N_10428,N_8808);
nor U15105 (N_15105,N_8733,N_9650);
nand U15106 (N_15106,N_8678,N_7814);
or U15107 (N_15107,N_7315,N_9997);
nand U15108 (N_15108,N_6655,N_8660);
nor U15109 (N_15109,N_10769,N_12269);
nor U15110 (N_15110,N_7656,N_9695);
nor U15111 (N_15111,N_9793,N_12219);
nor U15112 (N_15112,N_12130,N_10309);
and U15113 (N_15113,N_6833,N_8297);
nor U15114 (N_15114,N_6428,N_10429);
or U15115 (N_15115,N_9589,N_9775);
nand U15116 (N_15116,N_9308,N_11947);
nand U15117 (N_15117,N_8487,N_8694);
and U15118 (N_15118,N_11443,N_8286);
and U15119 (N_15119,N_10803,N_11751);
nand U15120 (N_15120,N_9579,N_8645);
nor U15121 (N_15121,N_7545,N_7947);
and U15122 (N_15122,N_8324,N_11925);
and U15123 (N_15123,N_11754,N_7687);
or U15124 (N_15124,N_8444,N_11997);
or U15125 (N_15125,N_10224,N_6252);
and U15126 (N_15126,N_7498,N_10911);
nor U15127 (N_15127,N_9719,N_6381);
nand U15128 (N_15128,N_9979,N_12000);
or U15129 (N_15129,N_8146,N_10806);
nor U15130 (N_15130,N_11861,N_8196);
nand U15131 (N_15131,N_8214,N_10695);
and U15132 (N_15132,N_8172,N_11515);
nor U15133 (N_15133,N_8564,N_10889);
xor U15134 (N_15134,N_6999,N_9998);
nor U15135 (N_15135,N_7237,N_9725);
or U15136 (N_15136,N_7704,N_6774);
or U15137 (N_15137,N_8309,N_8617);
and U15138 (N_15138,N_8301,N_7942);
nor U15139 (N_15139,N_11412,N_8585);
or U15140 (N_15140,N_6724,N_6593);
nor U15141 (N_15141,N_10822,N_8334);
and U15142 (N_15142,N_7838,N_8357);
nor U15143 (N_15143,N_10704,N_7156);
nand U15144 (N_15144,N_10424,N_6735);
nand U15145 (N_15145,N_7803,N_6278);
xnor U15146 (N_15146,N_9200,N_10316);
xor U15147 (N_15147,N_11025,N_10971);
or U15148 (N_15148,N_8696,N_8612);
nand U15149 (N_15149,N_11970,N_11778);
or U15150 (N_15150,N_7905,N_10140);
nor U15151 (N_15151,N_12086,N_6886);
or U15152 (N_15152,N_10410,N_8232);
nor U15153 (N_15153,N_6734,N_10483);
nor U15154 (N_15154,N_10021,N_9140);
and U15155 (N_15155,N_9251,N_6761);
and U15156 (N_15156,N_7810,N_9859);
nor U15157 (N_15157,N_8184,N_10106);
nor U15158 (N_15158,N_8436,N_10747);
and U15159 (N_15159,N_7263,N_9086);
nor U15160 (N_15160,N_7325,N_12157);
or U15161 (N_15161,N_8472,N_8836);
or U15162 (N_15162,N_7536,N_10692);
nand U15163 (N_15163,N_6395,N_11314);
or U15164 (N_15164,N_9264,N_8212);
or U15165 (N_15165,N_9020,N_9344);
nor U15166 (N_15166,N_12063,N_7635);
and U15167 (N_15167,N_11044,N_9960);
or U15168 (N_15168,N_7968,N_9744);
and U15169 (N_15169,N_7052,N_6776);
and U15170 (N_15170,N_7762,N_9597);
nand U15171 (N_15171,N_7869,N_6570);
nand U15172 (N_15172,N_7557,N_8865);
nor U15173 (N_15173,N_10572,N_9300);
nand U15174 (N_15174,N_7488,N_9083);
nand U15175 (N_15175,N_6509,N_8725);
or U15176 (N_15176,N_11922,N_7519);
and U15177 (N_15177,N_11613,N_9229);
nor U15178 (N_15178,N_7761,N_7203);
and U15179 (N_15179,N_10147,N_9917);
or U15180 (N_15180,N_11991,N_6397);
xor U15181 (N_15181,N_6800,N_6853);
nand U15182 (N_15182,N_11750,N_11315);
or U15183 (N_15183,N_11061,N_6971);
and U15184 (N_15184,N_10025,N_11288);
and U15185 (N_15185,N_9926,N_8721);
and U15186 (N_15186,N_11272,N_10055);
nor U15187 (N_15187,N_12293,N_9812);
and U15188 (N_15188,N_8891,N_7719);
or U15189 (N_15189,N_8541,N_6275);
and U15190 (N_15190,N_12259,N_8918);
and U15191 (N_15191,N_12423,N_7174);
nor U15192 (N_15192,N_11830,N_11540);
or U15193 (N_15193,N_10192,N_8895);
and U15194 (N_15194,N_6856,N_6645);
or U15195 (N_15195,N_7286,N_11192);
nor U15196 (N_15196,N_6652,N_11417);
or U15197 (N_15197,N_9261,N_7734);
or U15198 (N_15198,N_9154,N_9063);
and U15199 (N_15199,N_11081,N_7574);
or U15200 (N_15200,N_7493,N_12282);
xor U15201 (N_15201,N_9084,N_6438);
xor U15202 (N_15202,N_6308,N_6384);
xor U15203 (N_15203,N_7789,N_9715);
or U15204 (N_15204,N_8742,N_10479);
nor U15205 (N_15205,N_11436,N_12201);
nand U15206 (N_15206,N_11883,N_12053);
or U15207 (N_15207,N_11159,N_8268);
nor U15208 (N_15208,N_9035,N_9966);
nor U15209 (N_15209,N_10193,N_10943);
or U15210 (N_15210,N_11349,N_11807);
or U15211 (N_15211,N_6714,N_7777);
and U15212 (N_15212,N_10417,N_9348);
nor U15213 (N_15213,N_8577,N_10325);
or U15214 (N_15214,N_6858,N_8222);
nand U15215 (N_15215,N_8971,N_11979);
nor U15216 (N_15216,N_9946,N_12159);
and U15217 (N_15217,N_11996,N_9566);
nand U15218 (N_15218,N_11668,N_11198);
nor U15219 (N_15219,N_8656,N_6709);
nand U15220 (N_15220,N_9738,N_6908);
or U15221 (N_15221,N_7321,N_11317);
and U15222 (N_15222,N_11909,N_10115);
nor U15223 (N_15223,N_7105,N_9676);
and U15224 (N_15224,N_8672,N_7324);
nand U15225 (N_15225,N_11460,N_12077);
xnor U15226 (N_15226,N_8799,N_10778);
nor U15227 (N_15227,N_8550,N_10726);
nor U15228 (N_15228,N_8318,N_9006);
nor U15229 (N_15229,N_12453,N_11238);
nand U15230 (N_15230,N_7267,N_10508);
nor U15231 (N_15231,N_8465,N_7508);
nand U15232 (N_15232,N_10520,N_11242);
and U15233 (N_15233,N_9461,N_11604);
nor U15234 (N_15234,N_9054,N_9099);
and U15235 (N_15235,N_11035,N_6981);
and U15236 (N_15236,N_11958,N_9873);
and U15237 (N_15237,N_10874,N_10456);
nand U15238 (N_15238,N_9545,N_6785);
or U15239 (N_15239,N_8494,N_7096);
and U15240 (N_15240,N_9854,N_7329);
nand U15241 (N_15241,N_8244,N_7959);
and U15242 (N_15242,N_9046,N_10744);
nor U15243 (N_15243,N_8624,N_6466);
nor U15244 (N_15244,N_8926,N_9982);
xnor U15245 (N_15245,N_10028,N_7847);
nor U15246 (N_15246,N_10555,N_11631);
and U15247 (N_15247,N_8522,N_11990);
and U15248 (N_15248,N_6270,N_12113);
and U15249 (N_15249,N_6963,N_8281);
nor U15250 (N_15250,N_12229,N_6938);
or U15251 (N_15251,N_7610,N_8095);
nand U15252 (N_15252,N_9137,N_9101);
nor U15253 (N_15253,N_9092,N_10050);
xor U15254 (N_15254,N_8952,N_10611);
and U15255 (N_15255,N_9727,N_8510);
and U15256 (N_15256,N_8546,N_6879);
and U15257 (N_15257,N_7308,N_7030);
and U15258 (N_15258,N_9656,N_9245);
xor U15259 (N_15259,N_7745,N_10306);
nand U15260 (N_15260,N_8875,N_10815);
nand U15261 (N_15261,N_11468,N_11408);
and U15262 (N_15262,N_8234,N_11865);
or U15263 (N_15263,N_10293,N_9112);
nand U15264 (N_15264,N_9528,N_11438);
and U15265 (N_15265,N_9359,N_8430);
and U15266 (N_15266,N_12094,N_12313);
xnor U15267 (N_15267,N_6713,N_7804);
nand U15268 (N_15268,N_9195,N_7569);
nand U15269 (N_15269,N_9934,N_7932);
or U15270 (N_15270,N_11168,N_9518);
and U15271 (N_15271,N_11339,N_6569);
xnor U15272 (N_15272,N_7318,N_7621);
nor U15273 (N_15273,N_7588,N_11998);
or U15274 (N_15274,N_12129,N_9783);
xor U15275 (N_15275,N_9951,N_6577);
nor U15276 (N_15276,N_11730,N_10856);
xor U15277 (N_15277,N_6515,N_7978);
or U15278 (N_15278,N_9577,N_10363);
nor U15279 (N_15279,N_9188,N_6574);
nand U15280 (N_15280,N_6261,N_7122);
nand U15281 (N_15281,N_7037,N_9628);
xor U15282 (N_15282,N_8539,N_9876);
and U15283 (N_15283,N_8608,N_7475);
nor U15284 (N_15284,N_6427,N_12371);
and U15285 (N_15285,N_9524,N_7045);
nor U15286 (N_15286,N_9047,N_10988);
or U15287 (N_15287,N_11736,N_6701);
and U15288 (N_15288,N_9907,N_12001);
nand U15289 (N_15289,N_8683,N_10920);
or U15290 (N_15290,N_11231,N_10440);
or U15291 (N_15291,N_7565,N_9286);
nand U15292 (N_15292,N_12176,N_6393);
and U15293 (N_15293,N_8159,N_10753);
xnor U15294 (N_15294,N_7043,N_11720);
and U15295 (N_15295,N_7641,N_11441);
nor U15296 (N_15296,N_9209,N_7813);
and U15297 (N_15297,N_7906,N_11502);
or U15298 (N_15298,N_8396,N_10217);
nor U15299 (N_15299,N_6892,N_9125);
or U15300 (N_15300,N_11893,N_7298);
or U15301 (N_15301,N_8435,N_9561);
nand U15302 (N_15302,N_11780,N_11747);
nor U15303 (N_15303,N_8920,N_7175);
or U15304 (N_15304,N_8432,N_11586);
nand U15305 (N_15305,N_11981,N_11610);
nor U15306 (N_15306,N_8845,N_10696);
xor U15307 (N_15307,N_9401,N_12100);
and U15308 (N_15308,N_7675,N_10226);
xnor U15309 (N_15309,N_11527,N_11214);
xnor U15310 (N_15310,N_6524,N_9808);
or U15311 (N_15311,N_8800,N_11255);
nor U15312 (N_15312,N_12064,N_8298);
or U15313 (N_15313,N_10749,N_11678);
and U15314 (N_15314,N_7252,N_9514);
and U15315 (N_15315,N_9459,N_7139);
and U15316 (N_15316,N_8236,N_10869);
xor U15317 (N_15317,N_7553,N_10346);
nor U15318 (N_15318,N_7474,N_8090);
or U15319 (N_15319,N_12460,N_9155);
nand U15320 (N_15320,N_9269,N_11151);
nand U15321 (N_15321,N_11221,N_12022);
nand U15322 (N_15322,N_6902,N_9210);
or U15323 (N_15323,N_9362,N_11889);
nand U15324 (N_15324,N_9878,N_6731);
nand U15325 (N_15325,N_9961,N_12358);
and U15326 (N_15326,N_12353,N_10389);
nand U15327 (N_15327,N_9265,N_7422);
or U15328 (N_15328,N_8688,N_6257);
or U15329 (N_15329,N_8046,N_12011);
and U15330 (N_15330,N_7556,N_12058);
or U15331 (N_15331,N_9759,N_10906);
nand U15332 (N_15332,N_12482,N_9464);
or U15333 (N_15333,N_11290,N_6924);
nand U15334 (N_15334,N_7065,N_9396);
and U15335 (N_15335,N_6514,N_7012);
or U15336 (N_15336,N_9833,N_11932);
or U15337 (N_15337,N_10670,N_8455);
nand U15338 (N_15338,N_7360,N_8810);
or U15339 (N_15339,N_8459,N_9601);
and U15340 (N_15340,N_11281,N_10439);
nor U15341 (N_15341,N_10819,N_9273);
nand U15342 (N_15342,N_9098,N_12146);
xnor U15343 (N_15343,N_6298,N_7002);
nand U15344 (N_15344,N_11956,N_9544);
or U15345 (N_15345,N_9598,N_9751);
and U15346 (N_15346,N_7689,N_11072);
and U15347 (N_15347,N_6583,N_12493);
or U15348 (N_15348,N_7511,N_6425);
nor U15349 (N_15349,N_11457,N_7945);
nand U15350 (N_15350,N_7192,N_10813);
nand U15351 (N_15351,N_9230,N_10640);
nand U15352 (N_15352,N_6584,N_8227);
nand U15353 (N_15353,N_9435,N_10880);
nand U15354 (N_15354,N_7852,N_7663);
and U15355 (N_15355,N_9649,N_6594);
nand U15356 (N_15356,N_6352,N_7825);
or U15357 (N_15357,N_9900,N_11010);
xor U15358 (N_15358,N_6671,N_9093);
nand U15359 (N_15359,N_11098,N_8031);
nand U15360 (N_15360,N_7752,N_10592);
or U15361 (N_15361,N_6287,N_9568);
nor U15362 (N_15362,N_11976,N_12232);
and U15363 (N_15363,N_8807,N_11656);
nor U15364 (N_15364,N_10209,N_6750);
nor U15365 (N_15365,N_10705,N_6313);
nand U15366 (N_15366,N_8680,N_12262);
nor U15367 (N_15367,N_8129,N_11456);
nor U15368 (N_15368,N_6893,N_6670);
nand U15369 (N_15369,N_7093,N_8965);
nand U15370 (N_15370,N_12496,N_10453);
or U15371 (N_15371,N_12334,N_9363);
or U15372 (N_15372,N_11262,N_12383);
and U15373 (N_15373,N_12147,N_7089);
nor U15374 (N_15374,N_10875,N_8676);
or U15375 (N_15375,N_11895,N_7811);
and U15376 (N_15376,N_6532,N_7326);
nor U15377 (N_15377,N_10644,N_12380);
or U15378 (N_15378,N_11993,N_12361);
or U15379 (N_15379,N_12390,N_7563);
and U15380 (N_15380,N_7061,N_7746);
or U15381 (N_15381,N_11162,N_12454);
and U15382 (N_15382,N_11171,N_9693);
xor U15383 (N_15383,N_8531,N_10513);
and U15384 (N_15384,N_9694,N_7499);
nor U15385 (N_15385,N_9621,N_8080);
xor U15386 (N_15386,N_7451,N_12008);
nor U15387 (N_15387,N_12477,N_9761);
nor U15388 (N_15388,N_9236,N_8201);
or U15389 (N_15389,N_10639,N_10752);
xnor U15390 (N_15390,N_6523,N_7457);
nand U15391 (N_15391,N_8857,N_8537);
xor U15392 (N_15392,N_8888,N_9238);
nor U15393 (N_15393,N_6632,N_11662);
and U15394 (N_15394,N_10270,N_6417);
xor U15395 (N_15395,N_10153,N_6882);
nand U15396 (N_15396,N_10373,N_6337);
and U15397 (N_15397,N_9301,N_6465);
nor U15398 (N_15398,N_6660,N_10597);
xor U15399 (N_15399,N_8039,N_12121);
nand U15400 (N_15400,N_12468,N_9293);
nand U15401 (N_15401,N_12439,N_8000);
nand U15402 (N_15402,N_8217,N_9567);
xor U15403 (N_15403,N_9972,N_12082);
nand U15404 (N_15404,N_10686,N_9274);
nor U15405 (N_15405,N_6972,N_11792);
and U15406 (N_15406,N_8424,N_11011);
nor U15407 (N_15407,N_8299,N_11291);
or U15408 (N_15408,N_9345,N_7694);
or U15409 (N_15409,N_6454,N_6985);
xor U15410 (N_15410,N_8077,N_8503);
and U15411 (N_15411,N_6979,N_9415);
xnor U15412 (N_15412,N_8183,N_10773);
xor U15413 (N_15413,N_7477,N_7491);
nor U15414 (N_15414,N_8869,N_7562);
or U15415 (N_15415,N_8513,N_11390);
or U15416 (N_15416,N_11768,N_8431);
nor U15417 (N_15417,N_7861,N_9795);
nor U15418 (N_15418,N_8154,N_12093);
or U15419 (N_15419,N_9970,N_12473);
and U15420 (N_15420,N_12329,N_8005);
or U15421 (N_15421,N_11746,N_9104);
nor U15422 (N_15422,N_8916,N_10619);
or U15423 (N_15423,N_11150,N_11140);
xnor U15424 (N_15424,N_11556,N_9275);
or U15425 (N_15425,N_7333,N_9729);
nor U15426 (N_15426,N_12416,N_11051);
nor U15427 (N_15427,N_6522,N_9480);
nand U15428 (N_15428,N_10458,N_12305);
nor U15429 (N_15429,N_10194,N_8892);
or U15430 (N_15430,N_6324,N_11587);
and U15431 (N_15431,N_7221,N_11009);
or U15432 (N_15432,N_8442,N_10586);
or U15433 (N_15433,N_11798,N_7850);
nand U15434 (N_15434,N_9622,N_7157);
nor U15435 (N_15435,N_8717,N_7637);
and U15436 (N_15436,N_12273,N_11573);
or U15437 (N_15437,N_10091,N_8772);
nor U15438 (N_15438,N_11888,N_7957);
nor U15439 (N_15439,N_8831,N_12471);
nand U15440 (N_15440,N_8649,N_11759);
nand U15441 (N_15441,N_8292,N_8838);
nand U15442 (N_15442,N_6499,N_9733);
nor U15443 (N_15443,N_7592,N_11646);
nor U15444 (N_15444,N_6610,N_7469);
or U15445 (N_15445,N_6907,N_11091);
and U15446 (N_15446,N_8780,N_11823);
or U15447 (N_15447,N_9789,N_8654);
or U15448 (N_15448,N_11056,N_11898);
nand U15449 (N_15449,N_7953,N_7603);
nor U15450 (N_15450,N_7361,N_7201);
xor U15451 (N_15451,N_10086,N_8620);
nor U15452 (N_15452,N_7518,N_8607);
nand U15453 (N_15453,N_8353,N_10352);
or U15454 (N_15454,N_12495,N_12244);
and U15455 (N_15455,N_11006,N_7312);
xor U15456 (N_15456,N_10571,N_9120);
nor U15457 (N_15457,N_8861,N_8997);
xnor U15458 (N_15458,N_7558,N_6870);
and U15459 (N_15459,N_6895,N_10317);
and U15460 (N_15460,N_9439,N_9570);
nor U15461 (N_15461,N_10546,N_8830);
or U15462 (N_15462,N_8332,N_9522);
nor U15463 (N_15463,N_7285,N_8834);
or U15464 (N_15464,N_11270,N_12241);
nand U15465 (N_15465,N_7802,N_9930);
and U15466 (N_15466,N_8851,N_11664);
and U15467 (N_15467,N_6286,N_11600);
nor U15468 (N_15468,N_11202,N_6928);
or U15469 (N_15469,N_9296,N_6336);
and U15470 (N_15470,N_7753,N_11169);
nand U15471 (N_15471,N_7109,N_12173);
nand U15472 (N_15472,N_12164,N_9323);
and U15473 (N_15473,N_9460,N_8429);
and U15474 (N_15474,N_6469,N_11806);
nor U15475 (N_15475,N_8795,N_8058);
nor U15476 (N_15476,N_11466,N_10564);
and U15477 (N_15477,N_11304,N_10390);
nor U15478 (N_15478,N_6656,N_9133);
or U15479 (N_15479,N_10721,N_10814);
or U15480 (N_15480,N_11634,N_12348);
and U15481 (N_15481,N_12459,N_10094);
nand U15482 (N_15482,N_9864,N_7140);
and U15483 (N_15483,N_11252,N_8819);
xor U15484 (N_15484,N_11181,N_7892);
nand U15485 (N_15485,N_8243,N_12060);
or U15486 (N_15486,N_7795,N_10536);
and U15487 (N_15487,N_7356,N_6430);
or U15488 (N_15488,N_6864,N_10858);
nand U15489 (N_15489,N_6821,N_7877);
nand U15490 (N_15490,N_9285,N_11625);
or U15491 (N_15491,N_9994,N_8180);
and U15492 (N_15492,N_9716,N_11773);
xor U15493 (N_15493,N_7521,N_9355);
nor U15494 (N_15494,N_8496,N_8788);
nand U15495 (N_15495,N_12490,N_7238);
and U15496 (N_15496,N_7815,N_7173);
or U15497 (N_15497,N_10890,N_6627);
xor U15498 (N_15498,N_12381,N_9252);
nor U15499 (N_15499,N_11128,N_12067);
nand U15500 (N_15500,N_8571,N_11125);
or U15501 (N_15501,N_7098,N_7316);
or U15502 (N_15502,N_9237,N_7818);
nor U15503 (N_15503,N_6367,N_7808);
nand U15504 (N_15504,N_6256,N_7134);
nor U15505 (N_15505,N_8597,N_11397);
nand U15506 (N_15506,N_10133,N_10261);
nor U15507 (N_15507,N_6665,N_10770);
nor U15508 (N_15508,N_6452,N_6969);
xnor U15509 (N_15509,N_6464,N_9418);
and U15510 (N_15510,N_12048,N_12322);
nand U15511 (N_15511,N_12373,N_7602);
nand U15512 (N_15512,N_6906,N_11226);
or U15513 (N_15513,N_7594,N_11071);
and U15514 (N_15514,N_12144,N_7616);
nand U15515 (N_15515,N_6404,N_10512);
nand U15516 (N_15516,N_6429,N_12127);
or U15517 (N_15517,N_9159,N_12092);
nor U15518 (N_15518,N_8409,N_11120);
xnor U15519 (N_15519,N_12498,N_7834);
and U15520 (N_15520,N_11769,N_11258);
or U15521 (N_15521,N_7427,N_6759);
nand U15522 (N_15522,N_11860,N_11835);
or U15523 (N_15523,N_8901,N_10702);
nand U15524 (N_15524,N_6283,N_8703);
or U15525 (N_15525,N_10877,N_8199);
nor U15526 (N_15526,N_9171,N_11302);
xnor U15527 (N_15527,N_11507,N_11698);
or U15528 (N_15528,N_10984,N_7559);
xnor U15529 (N_15529,N_8560,N_6319);
nor U15530 (N_15530,N_11261,N_7447);
nand U15531 (N_15531,N_10074,N_6903);
nand U15532 (N_15532,N_11024,N_11039);
or U15533 (N_15533,N_9413,N_7614);
nand U15534 (N_15534,N_9517,N_8115);
nand U15535 (N_15535,N_9510,N_10119);
nand U15536 (N_15536,N_6968,N_11285);
nand U15537 (N_15537,N_6768,N_10182);
nand U15538 (N_15538,N_12018,N_11642);
xnor U15539 (N_15539,N_10333,N_8979);
xor U15540 (N_15540,N_6311,N_11684);
and U15541 (N_15541,N_7817,N_7487);
nand U15542 (N_15542,N_9861,N_6318);
and U15543 (N_15543,N_6771,N_8365);
nor U15544 (N_15544,N_9588,N_11296);
nor U15545 (N_15545,N_11583,N_11384);
nor U15546 (N_15546,N_7764,N_8187);
nand U15547 (N_15547,N_9050,N_10730);
nor U15548 (N_15548,N_12145,N_10426);
nor U15549 (N_15549,N_10254,N_10197);
xor U15550 (N_15550,N_11413,N_12337);
nand U15551 (N_15551,N_10613,N_10535);
nand U15552 (N_15552,N_11767,N_9630);
nor U15553 (N_15553,N_10737,N_9807);
xor U15554 (N_15554,N_6889,N_7404);
nor U15555 (N_15555,N_9683,N_12177);
xor U15556 (N_15556,N_7392,N_9428);
nor U15557 (N_15557,N_10797,N_9674);
nand U15558 (N_15558,N_12253,N_7966);
nand U15559 (N_15559,N_8209,N_9156);
nand U15560 (N_15560,N_7693,N_6988);
nand U15561 (N_15561,N_12413,N_10257);
xor U15562 (N_15562,N_6547,N_9052);
xnor U15563 (N_15563,N_9548,N_11878);
and U15564 (N_15564,N_6447,N_7919);
nor U15565 (N_15565,N_6323,N_6607);
nor U15566 (N_15566,N_12091,N_11030);
nor U15567 (N_15567,N_12437,N_6763);
or U15568 (N_15568,N_8388,N_11570);
and U15569 (N_15569,N_11797,N_8065);
or U15570 (N_15570,N_7504,N_6303);
and U15571 (N_15571,N_10621,N_10779);
nand U15572 (N_15572,N_12013,N_10339);
and U15573 (N_15573,N_11203,N_10654);
and U15574 (N_15574,N_6885,N_11914);
nor U15575 (N_15575,N_9135,N_6364);
nand U15576 (N_15576,N_7509,N_7567);
nand U15577 (N_15577,N_7249,N_10188);
or U15578 (N_15578,N_8142,N_9456);
nand U15579 (N_15579,N_8091,N_8155);
xnor U15580 (N_15580,N_9842,N_9284);
or U15581 (N_15581,N_7059,N_9817);
or U15582 (N_15582,N_6504,N_9748);
or U15583 (N_15583,N_10109,N_8578);
or U15584 (N_15584,N_8759,N_10186);
nand U15585 (N_15585,N_8743,N_10845);
nor U15586 (N_15586,N_10759,N_12039);
nor U15587 (N_15587,N_9491,N_12271);
and U15588 (N_15588,N_11654,N_7283);
nand U15589 (N_15589,N_10830,N_9898);
xnor U15590 (N_15590,N_6281,N_9805);
or U15591 (N_15591,N_8811,N_8500);
and U15592 (N_15592,N_9787,N_11725);
nand U15593 (N_15593,N_7155,N_10515);
nand U15594 (N_15594,N_9971,N_11437);
or U15595 (N_15595,N_9468,N_6934);
nor U15596 (N_15596,N_12010,N_10832);
or U15597 (N_15597,N_9841,N_10929);
or U15598 (N_15598,N_7436,N_7464);
and U15599 (N_15599,N_11454,N_9581);
nor U15600 (N_15600,N_9944,N_6519);
or U15601 (N_15601,N_7976,N_12124);
or U15602 (N_15602,N_10307,N_12231);
nand U15603 (N_15603,N_6914,N_7712);
nor U15604 (N_15604,N_11832,N_10838);
and U15605 (N_15605,N_8471,N_7049);
and U15606 (N_15606,N_9698,N_8576);
xor U15607 (N_15607,N_8994,N_9223);
or U15608 (N_15608,N_7528,N_8489);
nand U15609 (N_15609,N_8756,N_9989);
nand U15610 (N_15610,N_9121,N_10764);
nand U15611 (N_15611,N_8906,N_9762);
nor U15612 (N_15612,N_7426,N_10849);
nor U15613 (N_15613,N_8467,N_12221);
nor U15614 (N_15614,N_7255,N_6484);
xnor U15615 (N_15615,N_11967,N_7771);
or U15616 (N_15616,N_9472,N_7190);
and U15617 (N_15617,N_9652,N_11479);
nor U15618 (N_15618,N_8879,N_10556);
nand U15619 (N_15619,N_11239,N_8482);
or U15620 (N_15620,N_11933,N_10604);
nor U15621 (N_15621,N_8804,N_6899);
and U15622 (N_15622,N_11511,N_8100);
and U15623 (N_15623,N_9303,N_9549);
and U15624 (N_15624,N_9501,N_7234);
nor U15625 (N_15625,N_11528,N_11878);
or U15626 (N_15626,N_10241,N_7838);
or U15627 (N_15627,N_7761,N_8652);
nand U15628 (N_15628,N_9662,N_9597);
and U15629 (N_15629,N_8845,N_6782);
or U15630 (N_15630,N_7068,N_12428);
xnor U15631 (N_15631,N_8769,N_6289);
or U15632 (N_15632,N_9765,N_12347);
and U15633 (N_15633,N_7112,N_10156);
xnor U15634 (N_15634,N_11143,N_7411);
nor U15635 (N_15635,N_12394,N_7969);
and U15636 (N_15636,N_9794,N_8792);
nand U15637 (N_15637,N_7426,N_10361);
or U15638 (N_15638,N_9256,N_7243);
nor U15639 (N_15639,N_10970,N_9724);
nor U15640 (N_15640,N_11576,N_10252);
nor U15641 (N_15641,N_6414,N_8549);
nand U15642 (N_15642,N_10891,N_6618);
or U15643 (N_15643,N_7360,N_7372);
and U15644 (N_15644,N_11891,N_10668);
nor U15645 (N_15645,N_10593,N_8206);
nor U15646 (N_15646,N_8290,N_10533);
or U15647 (N_15647,N_7115,N_6998);
and U15648 (N_15648,N_10695,N_8996);
and U15649 (N_15649,N_12388,N_10329);
xor U15650 (N_15650,N_6460,N_8757);
nor U15651 (N_15651,N_9124,N_7069);
and U15652 (N_15652,N_10048,N_11956);
nor U15653 (N_15653,N_11698,N_7957);
and U15654 (N_15654,N_11955,N_7729);
nand U15655 (N_15655,N_11058,N_6969);
nor U15656 (N_15656,N_6782,N_8023);
and U15657 (N_15657,N_8658,N_12094);
and U15658 (N_15658,N_10888,N_7532);
nor U15659 (N_15659,N_9807,N_7649);
or U15660 (N_15660,N_10029,N_11997);
nor U15661 (N_15661,N_7063,N_11562);
nand U15662 (N_15662,N_12323,N_8506);
nand U15663 (N_15663,N_11536,N_7012);
or U15664 (N_15664,N_7977,N_8022);
or U15665 (N_15665,N_9600,N_11652);
and U15666 (N_15666,N_8951,N_10418);
nand U15667 (N_15667,N_8556,N_7628);
or U15668 (N_15668,N_7772,N_7740);
xnor U15669 (N_15669,N_11821,N_12328);
nor U15670 (N_15670,N_7498,N_8843);
or U15671 (N_15671,N_8023,N_7876);
or U15672 (N_15672,N_7949,N_6751);
nor U15673 (N_15673,N_8416,N_10968);
or U15674 (N_15674,N_6771,N_9168);
and U15675 (N_15675,N_11367,N_8204);
nor U15676 (N_15676,N_8874,N_8152);
nor U15677 (N_15677,N_11241,N_9706);
nor U15678 (N_15678,N_7911,N_7146);
and U15679 (N_15679,N_9861,N_9359);
nor U15680 (N_15680,N_12230,N_12002);
xor U15681 (N_15681,N_8264,N_12320);
or U15682 (N_15682,N_8029,N_6373);
nor U15683 (N_15683,N_9097,N_11020);
or U15684 (N_15684,N_10208,N_6758);
nand U15685 (N_15685,N_7880,N_8905);
or U15686 (N_15686,N_9147,N_7474);
nor U15687 (N_15687,N_7863,N_12020);
nor U15688 (N_15688,N_7661,N_11420);
or U15689 (N_15689,N_11190,N_11223);
or U15690 (N_15690,N_9959,N_10985);
nand U15691 (N_15691,N_7911,N_10619);
nand U15692 (N_15692,N_11965,N_7044);
xor U15693 (N_15693,N_6364,N_8562);
nor U15694 (N_15694,N_10453,N_12470);
or U15695 (N_15695,N_10102,N_9853);
nand U15696 (N_15696,N_11739,N_12114);
and U15697 (N_15697,N_10184,N_9132);
or U15698 (N_15698,N_8137,N_11866);
xor U15699 (N_15699,N_10864,N_12267);
nor U15700 (N_15700,N_6956,N_8729);
or U15701 (N_15701,N_10905,N_11217);
nand U15702 (N_15702,N_6693,N_11992);
and U15703 (N_15703,N_10502,N_10853);
nand U15704 (N_15704,N_11170,N_9839);
and U15705 (N_15705,N_7709,N_10353);
and U15706 (N_15706,N_9207,N_8894);
or U15707 (N_15707,N_9485,N_9100);
and U15708 (N_15708,N_11062,N_8077);
and U15709 (N_15709,N_9479,N_6395);
and U15710 (N_15710,N_6455,N_6373);
or U15711 (N_15711,N_10502,N_10422);
or U15712 (N_15712,N_10286,N_9792);
and U15713 (N_15713,N_9759,N_8487);
xor U15714 (N_15714,N_12414,N_9082);
and U15715 (N_15715,N_10021,N_11272);
and U15716 (N_15716,N_7518,N_10751);
nand U15717 (N_15717,N_10758,N_11454);
nand U15718 (N_15718,N_12231,N_8444);
and U15719 (N_15719,N_10132,N_10914);
xor U15720 (N_15720,N_12286,N_11875);
nand U15721 (N_15721,N_8141,N_8466);
nand U15722 (N_15722,N_6808,N_9353);
or U15723 (N_15723,N_12337,N_7548);
xnor U15724 (N_15724,N_8662,N_10152);
xor U15725 (N_15725,N_9005,N_10724);
nor U15726 (N_15726,N_9997,N_9038);
nor U15727 (N_15727,N_9956,N_11014);
or U15728 (N_15728,N_12496,N_8409);
nand U15729 (N_15729,N_6253,N_12438);
and U15730 (N_15730,N_6403,N_7692);
or U15731 (N_15731,N_9983,N_7225);
nand U15732 (N_15732,N_7864,N_9425);
nand U15733 (N_15733,N_10900,N_10907);
nand U15734 (N_15734,N_10485,N_11962);
and U15735 (N_15735,N_7183,N_12061);
and U15736 (N_15736,N_8255,N_9006);
nand U15737 (N_15737,N_9610,N_8430);
and U15738 (N_15738,N_12350,N_9336);
nor U15739 (N_15739,N_10555,N_12189);
and U15740 (N_15740,N_7718,N_10664);
nor U15741 (N_15741,N_7292,N_6782);
nor U15742 (N_15742,N_7486,N_12491);
nand U15743 (N_15743,N_8974,N_9013);
xnor U15744 (N_15744,N_12367,N_10012);
or U15745 (N_15745,N_7030,N_6755);
xnor U15746 (N_15746,N_12482,N_10918);
nand U15747 (N_15747,N_12332,N_10158);
and U15748 (N_15748,N_12043,N_11304);
and U15749 (N_15749,N_8203,N_8424);
and U15750 (N_15750,N_8371,N_9875);
nor U15751 (N_15751,N_11774,N_10808);
xnor U15752 (N_15752,N_11255,N_12190);
xor U15753 (N_15753,N_7433,N_10588);
and U15754 (N_15754,N_10253,N_9588);
and U15755 (N_15755,N_9133,N_7467);
nor U15756 (N_15756,N_10951,N_7573);
and U15757 (N_15757,N_11419,N_9441);
nand U15758 (N_15758,N_9892,N_6856);
or U15759 (N_15759,N_12412,N_6362);
and U15760 (N_15760,N_8464,N_6814);
nand U15761 (N_15761,N_9469,N_7974);
nor U15762 (N_15762,N_8103,N_9804);
nand U15763 (N_15763,N_11790,N_6258);
or U15764 (N_15764,N_10657,N_10856);
and U15765 (N_15765,N_9643,N_12259);
nor U15766 (N_15766,N_11682,N_12199);
xor U15767 (N_15767,N_9764,N_10260);
xnor U15768 (N_15768,N_10620,N_10300);
and U15769 (N_15769,N_12203,N_6432);
or U15770 (N_15770,N_9149,N_8723);
or U15771 (N_15771,N_9282,N_11963);
nor U15772 (N_15772,N_8080,N_11878);
nand U15773 (N_15773,N_7513,N_8323);
xor U15774 (N_15774,N_6331,N_11839);
and U15775 (N_15775,N_11590,N_6805);
nor U15776 (N_15776,N_8310,N_11034);
and U15777 (N_15777,N_9595,N_7519);
or U15778 (N_15778,N_12010,N_9383);
or U15779 (N_15779,N_9167,N_9429);
or U15780 (N_15780,N_10610,N_10476);
xor U15781 (N_15781,N_11526,N_8888);
and U15782 (N_15782,N_10048,N_11621);
xor U15783 (N_15783,N_6577,N_6919);
nor U15784 (N_15784,N_9941,N_11996);
or U15785 (N_15785,N_10509,N_7800);
or U15786 (N_15786,N_11618,N_10880);
xor U15787 (N_15787,N_8904,N_6570);
and U15788 (N_15788,N_11289,N_10906);
or U15789 (N_15789,N_9267,N_6500);
nand U15790 (N_15790,N_7541,N_7715);
and U15791 (N_15791,N_10585,N_6709);
nand U15792 (N_15792,N_10910,N_7739);
nor U15793 (N_15793,N_9751,N_10083);
nor U15794 (N_15794,N_7125,N_9632);
and U15795 (N_15795,N_8979,N_9538);
nand U15796 (N_15796,N_8912,N_10122);
nor U15797 (N_15797,N_12431,N_8714);
nor U15798 (N_15798,N_7758,N_9297);
or U15799 (N_15799,N_6721,N_12482);
nand U15800 (N_15800,N_7435,N_6742);
nor U15801 (N_15801,N_10031,N_12226);
nor U15802 (N_15802,N_7886,N_9129);
nand U15803 (N_15803,N_7143,N_11362);
nor U15804 (N_15804,N_7536,N_9805);
nor U15805 (N_15805,N_7882,N_9656);
xnor U15806 (N_15806,N_10892,N_10463);
nand U15807 (N_15807,N_11983,N_9828);
nand U15808 (N_15808,N_6798,N_11879);
xnor U15809 (N_15809,N_7708,N_9304);
nand U15810 (N_15810,N_8682,N_9759);
nand U15811 (N_15811,N_8556,N_10868);
nand U15812 (N_15812,N_11996,N_12012);
nor U15813 (N_15813,N_8354,N_8180);
or U15814 (N_15814,N_12347,N_10256);
or U15815 (N_15815,N_10384,N_9836);
and U15816 (N_15816,N_7670,N_10624);
and U15817 (N_15817,N_8708,N_11498);
nor U15818 (N_15818,N_12137,N_6311);
and U15819 (N_15819,N_8162,N_10611);
nor U15820 (N_15820,N_12167,N_10218);
nand U15821 (N_15821,N_11525,N_9792);
nand U15822 (N_15822,N_11585,N_12438);
nand U15823 (N_15823,N_11416,N_11842);
xor U15824 (N_15824,N_7087,N_9333);
nand U15825 (N_15825,N_8702,N_10177);
nand U15826 (N_15826,N_7891,N_9429);
nor U15827 (N_15827,N_9105,N_10668);
and U15828 (N_15828,N_9875,N_7478);
and U15829 (N_15829,N_12101,N_11067);
nor U15830 (N_15830,N_7190,N_9376);
nand U15831 (N_15831,N_7338,N_6440);
nor U15832 (N_15832,N_11511,N_11830);
nand U15833 (N_15833,N_7911,N_9114);
and U15834 (N_15834,N_6300,N_7873);
or U15835 (N_15835,N_8404,N_8100);
nand U15836 (N_15836,N_7379,N_10438);
nand U15837 (N_15837,N_9200,N_10074);
nor U15838 (N_15838,N_7233,N_7022);
or U15839 (N_15839,N_7823,N_7826);
nor U15840 (N_15840,N_9705,N_9559);
nor U15841 (N_15841,N_6337,N_7238);
xor U15842 (N_15842,N_7180,N_11742);
nand U15843 (N_15843,N_10257,N_7209);
nand U15844 (N_15844,N_8044,N_10389);
nor U15845 (N_15845,N_12005,N_8477);
nand U15846 (N_15846,N_7564,N_7857);
nor U15847 (N_15847,N_8326,N_9656);
and U15848 (N_15848,N_7072,N_8623);
nor U15849 (N_15849,N_6836,N_7675);
nor U15850 (N_15850,N_12114,N_9568);
nand U15851 (N_15851,N_10815,N_6467);
and U15852 (N_15852,N_6732,N_10793);
and U15853 (N_15853,N_8306,N_6830);
nor U15854 (N_15854,N_9681,N_6351);
nor U15855 (N_15855,N_10291,N_10866);
or U15856 (N_15856,N_7108,N_12443);
and U15857 (N_15857,N_11773,N_9788);
and U15858 (N_15858,N_8680,N_7104);
and U15859 (N_15859,N_10437,N_7667);
or U15860 (N_15860,N_7259,N_9722);
nand U15861 (N_15861,N_10143,N_11286);
nor U15862 (N_15862,N_10223,N_9240);
xor U15863 (N_15863,N_8330,N_7570);
and U15864 (N_15864,N_6551,N_8521);
nor U15865 (N_15865,N_9577,N_9172);
nand U15866 (N_15866,N_10458,N_6854);
and U15867 (N_15867,N_9625,N_6660);
and U15868 (N_15868,N_10219,N_11460);
nor U15869 (N_15869,N_9858,N_11277);
and U15870 (N_15870,N_9304,N_12090);
and U15871 (N_15871,N_10030,N_7741);
and U15872 (N_15872,N_10498,N_10208);
and U15873 (N_15873,N_11593,N_7678);
or U15874 (N_15874,N_8967,N_9314);
nor U15875 (N_15875,N_10815,N_9741);
nand U15876 (N_15876,N_9478,N_12275);
nand U15877 (N_15877,N_8198,N_7186);
or U15878 (N_15878,N_6501,N_8036);
and U15879 (N_15879,N_12471,N_7552);
nor U15880 (N_15880,N_11010,N_12348);
nor U15881 (N_15881,N_8394,N_10736);
and U15882 (N_15882,N_7289,N_6835);
nor U15883 (N_15883,N_8084,N_7038);
nor U15884 (N_15884,N_11000,N_9004);
or U15885 (N_15885,N_9301,N_9025);
or U15886 (N_15886,N_10710,N_8178);
or U15887 (N_15887,N_6445,N_6394);
nand U15888 (N_15888,N_8984,N_11443);
xor U15889 (N_15889,N_9200,N_10491);
nor U15890 (N_15890,N_9017,N_10549);
nand U15891 (N_15891,N_11798,N_6485);
xnor U15892 (N_15892,N_6658,N_11500);
nor U15893 (N_15893,N_10441,N_9918);
xor U15894 (N_15894,N_7175,N_9400);
or U15895 (N_15895,N_9443,N_11325);
nor U15896 (N_15896,N_7754,N_6345);
nand U15897 (N_15897,N_10191,N_11945);
nor U15898 (N_15898,N_6347,N_6253);
nand U15899 (N_15899,N_8058,N_9770);
nand U15900 (N_15900,N_9788,N_12422);
nor U15901 (N_15901,N_6975,N_11095);
or U15902 (N_15902,N_10585,N_12065);
or U15903 (N_15903,N_12222,N_11352);
or U15904 (N_15904,N_7444,N_9115);
nor U15905 (N_15905,N_10980,N_6465);
xnor U15906 (N_15906,N_11560,N_6841);
nand U15907 (N_15907,N_10400,N_10326);
or U15908 (N_15908,N_9601,N_8514);
and U15909 (N_15909,N_7618,N_9393);
nand U15910 (N_15910,N_9894,N_12119);
nor U15911 (N_15911,N_6581,N_8428);
nor U15912 (N_15912,N_10335,N_9792);
or U15913 (N_15913,N_7356,N_7059);
or U15914 (N_15914,N_6401,N_9389);
nand U15915 (N_15915,N_12031,N_11352);
nor U15916 (N_15916,N_11000,N_11111);
and U15917 (N_15917,N_10510,N_7951);
nor U15918 (N_15918,N_9660,N_10553);
and U15919 (N_15919,N_9189,N_8260);
nor U15920 (N_15920,N_9186,N_11870);
and U15921 (N_15921,N_6887,N_11894);
nand U15922 (N_15922,N_8245,N_9813);
and U15923 (N_15923,N_11761,N_7719);
nand U15924 (N_15924,N_9603,N_6897);
nand U15925 (N_15925,N_10294,N_11362);
nand U15926 (N_15926,N_8405,N_8439);
xnor U15927 (N_15927,N_7185,N_11600);
nand U15928 (N_15928,N_10920,N_7657);
or U15929 (N_15929,N_12134,N_11861);
xnor U15930 (N_15930,N_8187,N_10281);
xnor U15931 (N_15931,N_8962,N_7469);
nor U15932 (N_15932,N_9814,N_10731);
or U15933 (N_15933,N_6920,N_6371);
xnor U15934 (N_15934,N_8151,N_6352);
nor U15935 (N_15935,N_7430,N_7785);
xor U15936 (N_15936,N_9399,N_6664);
nand U15937 (N_15937,N_10713,N_9819);
xnor U15938 (N_15938,N_8603,N_7363);
nor U15939 (N_15939,N_10863,N_10591);
nor U15940 (N_15940,N_11972,N_6908);
and U15941 (N_15941,N_6371,N_6801);
or U15942 (N_15942,N_9754,N_9712);
nor U15943 (N_15943,N_12005,N_11617);
xnor U15944 (N_15944,N_7803,N_6870);
and U15945 (N_15945,N_10320,N_10606);
nor U15946 (N_15946,N_10721,N_9445);
and U15947 (N_15947,N_12298,N_7549);
nor U15948 (N_15948,N_10676,N_7657);
xor U15949 (N_15949,N_9993,N_10224);
nand U15950 (N_15950,N_6378,N_7511);
and U15951 (N_15951,N_9161,N_11665);
and U15952 (N_15952,N_10808,N_10282);
and U15953 (N_15953,N_6698,N_9731);
or U15954 (N_15954,N_11232,N_6573);
nor U15955 (N_15955,N_9536,N_6337);
nor U15956 (N_15956,N_9823,N_7064);
and U15957 (N_15957,N_10596,N_9977);
nand U15958 (N_15958,N_10163,N_12448);
nor U15959 (N_15959,N_7390,N_11980);
nor U15960 (N_15960,N_8230,N_8673);
nand U15961 (N_15961,N_8661,N_9845);
and U15962 (N_15962,N_7862,N_11638);
nand U15963 (N_15963,N_11916,N_6688);
or U15964 (N_15964,N_9780,N_7108);
and U15965 (N_15965,N_8745,N_7622);
and U15966 (N_15966,N_11754,N_7057);
and U15967 (N_15967,N_9582,N_9291);
and U15968 (N_15968,N_7268,N_7703);
xnor U15969 (N_15969,N_8733,N_7203);
xor U15970 (N_15970,N_9267,N_10938);
and U15971 (N_15971,N_10566,N_9336);
and U15972 (N_15972,N_9360,N_11632);
xnor U15973 (N_15973,N_10562,N_7034);
or U15974 (N_15974,N_11921,N_10365);
nor U15975 (N_15975,N_6522,N_12141);
nor U15976 (N_15976,N_12308,N_8186);
or U15977 (N_15977,N_7161,N_6661);
nand U15978 (N_15978,N_9193,N_7621);
nor U15979 (N_15979,N_10914,N_8529);
or U15980 (N_15980,N_11420,N_10176);
nand U15981 (N_15981,N_8128,N_11436);
nand U15982 (N_15982,N_6943,N_12462);
xnor U15983 (N_15983,N_9742,N_9882);
nor U15984 (N_15984,N_11642,N_7596);
nand U15985 (N_15985,N_8415,N_9133);
nor U15986 (N_15986,N_8166,N_11060);
nor U15987 (N_15987,N_8549,N_6552);
or U15988 (N_15988,N_7158,N_12360);
or U15989 (N_15989,N_10963,N_7750);
and U15990 (N_15990,N_6915,N_10513);
and U15991 (N_15991,N_12115,N_11184);
nand U15992 (N_15992,N_7683,N_7978);
nor U15993 (N_15993,N_7238,N_10559);
and U15994 (N_15994,N_12009,N_9981);
nor U15995 (N_15995,N_6639,N_10541);
or U15996 (N_15996,N_7232,N_10373);
nand U15997 (N_15997,N_10053,N_8587);
nand U15998 (N_15998,N_10884,N_12408);
or U15999 (N_15999,N_9198,N_12170);
xor U16000 (N_16000,N_10005,N_9395);
and U16001 (N_16001,N_9546,N_12456);
nand U16002 (N_16002,N_10505,N_9037);
nand U16003 (N_16003,N_11194,N_6751);
and U16004 (N_16004,N_10556,N_12340);
and U16005 (N_16005,N_9856,N_9787);
nor U16006 (N_16006,N_7351,N_9399);
or U16007 (N_16007,N_11629,N_10892);
or U16008 (N_16008,N_8813,N_9478);
nand U16009 (N_16009,N_7214,N_11160);
or U16010 (N_16010,N_9217,N_10084);
or U16011 (N_16011,N_9826,N_7589);
and U16012 (N_16012,N_7512,N_7922);
or U16013 (N_16013,N_8217,N_9097);
nand U16014 (N_16014,N_8131,N_7961);
or U16015 (N_16015,N_6621,N_11904);
nand U16016 (N_16016,N_8470,N_12027);
xnor U16017 (N_16017,N_7649,N_10785);
or U16018 (N_16018,N_10169,N_10734);
and U16019 (N_16019,N_11608,N_7029);
xor U16020 (N_16020,N_12041,N_7808);
xnor U16021 (N_16021,N_7582,N_9348);
or U16022 (N_16022,N_6660,N_9899);
nor U16023 (N_16023,N_10529,N_9962);
nand U16024 (N_16024,N_11568,N_6382);
or U16025 (N_16025,N_6566,N_9052);
nand U16026 (N_16026,N_9486,N_7259);
and U16027 (N_16027,N_7235,N_10797);
xnor U16028 (N_16028,N_12158,N_6711);
xor U16029 (N_16029,N_11841,N_8361);
or U16030 (N_16030,N_11405,N_9865);
xnor U16031 (N_16031,N_7965,N_7617);
nor U16032 (N_16032,N_10121,N_7552);
and U16033 (N_16033,N_10151,N_8439);
and U16034 (N_16034,N_6923,N_9957);
nand U16035 (N_16035,N_10326,N_7256);
or U16036 (N_16036,N_8832,N_8192);
or U16037 (N_16037,N_10632,N_11048);
or U16038 (N_16038,N_6315,N_8468);
or U16039 (N_16039,N_10337,N_9578);
and U16040 (N_16040,N_7503,N_6838);
nand U16041 (N_16041,N_9578,N_8163);
or U16042 (N_16042,N_8452,N_7920);
nor U16043 (N_16043,N_6358,N_9370);
or U16044 (N_16044,N_10688,N_6858);
or U16045 (N_16045,N_11674,N_9045);
nor U16046 (N_16046,N_9871,N_7503);
nor U16047 (N_16047,N_11626,N_10939);
nand U16048 (N_16048,N_8666,N_6340);
xor U16049 (N_16049,N_6471,N_11246);
nor U16050 (N_16050,N_10316,N_12131);
nand U16051 (N_16051,N_8380,N_6965);
or U16052 (N_16052,N_7592,N_11917);
and U16053 (N_16053,N_9201,N_10130);
nand U16054 (N_16054,N_11996,N_10648);
and U16055 (N_16055,N_6569,N_9591);
and U16056 (N_16056,N_6254,N_7704);
xor U16057 (N_16057,N_10656,N_7237);
nand U16058 (N_16058,N_8793,N_10916);
nor U16059 (N_16059,N_8235,N_9708);
nand U16060 (N_16060,N_8763,N_11892);
and U16061 (N_16061,N_7144,N_8049);
nor U16062 (N_16062,N_8154,N_8790);
or U16063 (N_16063,N_9884,N_11871);
or U16064 (N_16064,N_8554,N_11374);
or U16065 (N_16065,N_12128,N_11942);
nor U16066 (N_16066,N_6864,N_7163);
nor U16067 (N_16067,N_11443,N_6486);
and U16068 (N_16068,N_7482,N_10845);
nand U16069 (N_16069,N_10849,N_10941);
nand U16070 (N_16070,N_6798,N_9272);
and U16071 (N_16071,N_6707,N_9334);
nand U16072 (N_16072,N_10623,N_6569);
xor U16073 (N_16073,N_7418,N_11896);
or U16074 (N_16074,N_11460,N_9712);
nor U16075 (N_16075,N_10333,N_12067);
and U16076 (N_16076,N_10572,N_11149);
or U16077 (N_16077,N_9968,N_10010);
nand U16078 (N_16078,N_7672,N_12197);
nor U16079 (N_16079,N_7419,N_6345);
nand U16080 (N_16080,N_9704,N_9132);
and U16081 (N_16081,N_10547,N_9123);
or U16082 (N_16082,N_11932,N_9209);
xor U16083 (N_16083,N_10423,N_9922);
nand U16084 (N_16084,N_9272,N_11770);
or U16085 (N_16085,N_9184,N_8845);
nor U16086 (N_16086,N_9026,N_8004);
and U16087 (N_16087,N_8140,N_10596);
nor U16088 (N_16088,N_12469,N_11791);
nand U16089 (N_16089,N_10282,N_9555);
nor U16090 (N_16090,N_10144,N_6636);
nor U16091 (N_16091,N_10019,N_12430);
or U16092 (N_16092,N_6357,N_11902);
nand U16093 (N_16093,N_10071,N_11756);
nor U16094 (N_16094,N_10717,N_11254);
or U16095 (N_16095,N_10088,N_11421);
nand U16096 (N_16096,N_11594,N_10814);
nand U16097 (N_16097,N_11452,N_10209);
or U16098 (N_16098,N_7814,N_10939);
and U16099 (N_16099,N_10102,N_7688);
xnor U16100 (N_16100,N_9339,N_10681);
nor U16101 (N_16101,N_7398,N_11059);
nand U16102 (N_16102,N_8313,N_6618);
nand U16103 (N_16103,N_8988,N_9045);
nand U16104 (N_16104,N_11383,N_10327);
nand U16105 (N_16105,N_7145,N_10096);
nand U16106 (N_16106,N_9812,N_10877);
nand U16107 (N_16107,N_8806,N_8719);
and U16108 (N_16108,N_9949,N_8761);
or U16109 (N_16109,N_11358,N_10832);
nand U16110 (N_16110,N_11060,N_9275);
and U16111 (N_16111,N_7988,N_6738);
nor U16112 (N_16112,N_6575,N_10212);
nand U16113 (N_16113,N_11307,N_10679);
nor U16114 (N_16114,N_8059,N_11791);
nor U16115 (N_16115,N_9703,N_8619);
and U16116 (N_16116,N_10157,N_11249);
or U16117 (N_16117,N_12453,N_7207);
nor U16118 (N_16118,N_10764,N_9534);
or U16119 (N_16119,N_12062,N_7304);
or U16120 (N_16120,N_8267,N_10789);
nor U16121 (N_16121,N_11961,N_10218);
nor U16122 (N_16122,N_9342,N_10024);
or U16123 (N_16123,N_8946,N_12036);
nand U16124 (N_16124,N_11315,N_7474);
nand U16125 (N_16125,N_7234,N_10584);
nor U16126 (N_16126,N_9382,N_6944);
or U16127 (N_16127,N_6521,N_11346);
and U16128 (N_16128,N_11477,N_8690);
or U16129 (N_16129,N_7352,N_9622);
and U16130 (N_16130,N_8930,N_11982);
nand U16131 (N_16131,N_10652,N_9139);
nand U16132 (N_16132,N_11646,N_12499);
and U16133 (N_16133,N_6410,N_12478);
nand U16134 (N_16134,N_10979,N_7899);
and U16135 (N_16135,N_11823,N_12047);
nand U16136 (N_16136,N_11726,N_8912);
or U16137 (N_16137,N_10331,N_10512);
and U16138 (N_16138,N_10175,N_11873);
xor U16139 (N_16139,N_7982,N_12277);
nor U16140 (N_16140,N_11554,N_7412);
xor U16141 (N_16141,N_8300,N_10007);
nand U16142 (N_16142,N_9876,N_11628);
or U16143 (N_16143,N_8724,N_6865);
or U16144 (N_16144,N_10719,N_8863);
xor U16145 (N_16145,N_9594,N_7168);
or U16146 (N_16146,N_8972,N_11215);
or U16147 (N_16147,N_10834,N_12430);
nand U16148 (N_16148,N_11590,N_6660);
and U16149 (N_16149,N_7544,N_7489);
nor U16150 (N_16150,N_8306,N_9372);
xor U16151 (N_16151,N_9024,N_8610);
nand U16152 (N_16152,N_9282,N_7690);
and U16153 (N_16153,N_9616,N_7393);
nor U16154 (N_16154,N_8045,N_7600);
and U16155 (N_16155,N_10130,N_8668);
nand U16156 (N_16156,N_9638,N_7285);
and U16157 (N_16157,N_11441,N_9853);
and U16158 (N_16158,N_11107,N_12059);
nand U16159 (N_16159,N_9457,N_8794);
and U16160 (N_16160,N_8390,N_11076);
nand U16161 (N_16161,N_8525,N_6569);
nor U16162 (N_16162,N_8736,N_8863);
nand U16163 (N_16163,N_9810,N_8184);
or U16164 (N_16164,N_9717,N_10081);
or U16165 (N_16165,N_7617,N_9378);
or U16166 (N_16166,N_8376,N_6366);
xor U16167 (N_16167,N_10458,N_12174);
and U16168 (N_16168,N_10926,N_9971);
or U16169 (N_16169,N_10697,N_8407);
or U16170 (N_16170,N_12194,N_8170);
and U16171 (N_16171,N_7649,N_8004);
or U16172 (N_16172,N_10990,N_11935);
and U16173 (N_16173,N_7754,N_6794);
nand U16174 (N_16174,N_9155,N_9675);
nor U16175 (N_16175,N_6445,N_8869);
xnor U16176 (N_16176,N_9959,N_9204);
nor U16177 (N_16177,N_12024,N_9975);
and U16178 (N_16178,N_7311,N_9909);
or U16179 (N_16179,N_8595,N_12059);
nand U16180 (N_16180,N_7956,N_8564);
and U16181 (N_16181,N_10155,N_8237);
or U16182 (N_16182,N_10394,N_10589);
nand U16183 (N_16183,N_9983,N_8403);
nand U16184 (N_16184,N_11159,N_6519);
nor U16185 (N_16185,N_9807,N_7722);
nand U16186 (N_16186,N_6967,N_6985);
or U16187 (N_16187,N_12127,N_7907);
and U16188 (N_16188,N_10281,N_8747);
nor U16189 (N_16189,N_7434,N_11558);
nor U16190 (N_16190,N_12044,N_7685);
or U16191 (N_16191,N_8925,N_6528);
nand U16192 (N_16192,N_8228,N_11677);
nand U16193 (N_16193,N_10685,N_8592);
nand U16194 (N_16194,N_7551,N_11734);
nand U16195 (N_16195,N_10787,N_11263);
and U16196 (N_16196,N_9023,N_8527);
and U16197 (N_16197,N_6392,N_6450);
or U16198 (N_16198,N_7336,N_10348);
and U16199 (N_16199,N_10438,N_11850);
or U16200 (N_16200,N_10449,N_11853);
and U16201 (N_16201,N_7367,N_11164);
xor U16202 (N_16202,N_7611,N_7406);
and U16203 (N_16203,N_9052,N_8727);
nor U16204 (N_16204,N_12250,N_6466);
nand U16205 (N_16205,N_8306,N_10062);
and U16206 (N_16206,N_11202,N_9065);
or U16207 (N_16207,N_10172,N_9445);
or U16208 (N_16208,N_10848,N_10235);
xor U16209 (N_16209,N_11429,N_6359);
and U16210 (N_16210,N_7696,N_11295);
or U16211 (N_16211,N_9744,N_8361);
and U16212 (N_16212,N_11799,N_11848);
xor U16213 (N_16213,N_11335,N_9588);
or U16214 (N_16214,N_7994,N_11534);
nand U16215 (N_16215,N_9707,N_7903);
nor U16216 (N_16216,N_9822,N_8058);
xnor U16217 (N_16217,N_11712,N_12260);
nand U16218 (N_16218,N_6300,N_11536);
nand U16219 (N_16219,N_12134,N_8563);
or U16220 (N_16220,N_11879,N_10659);
nand U16221 (N_16221,N_10509,N_6335);
or U16222 (N_16222,N_11503,N_10260);
nand U16223 (N_16223,N_10169,N_8151);
or U16224 (N_16224,N_10549,N_7726);
or U16225 (N_16225,N_11350,N_7619);
and U16226 (N_16226,N_6491,N_10851);
nor U16227 (N_16227,N_8037,N_7107);
or U16228 (N_16228,N_8490,N_7925);
nor U16229 (N_16229,N_11583,N_10548);
nor U16230 (N_16230,N_8631,N_10579);
nor U16231 (N_16231,N_9954,N_7020);
or U16232 (N_16232,N_10496,N_11444);
or U16233 (N_16233,N_7760,N_11267);
and U16234 (N_16234,N_10139,N_7961);
nor U16235 (N_16235,N_6613,N_8958);
or U16236 (N_16236,N_7478,N_7681);
and U16237 (N_16237,N_6659,N_10439);
nand U16238 (N_16238,N_8442,N_10773);
nand U16239 (N_16239,N_8338,N_9392);
or U16240 (N_16240,N_9099,N_11648);
nand U16241 (N_16241,N_12132,N_8074);
nor U16242 (N_16242,N_12429,N_8953);
nor U16243 (N_16243,N_11706,N_10201);
xor U16244 (N_16244,N_12464,N_11511);
and U16245 (N_16245,N_11781,N_11243);
and U16246 (N_16246,N_10687,N_6694);
or U16247 (N_16247,N_9480,N_8863);
or U16248 (N_16248,N_7340,N_11704);
nor U16249 (N_16249,N_9101,N_9185);
or U16250 (N_16250,N_10548,N_7601);
nor U16251 (N_16251,N_6452,N_9711);
xor U16252 (N_16252,N_7817,N_6595);
or U16253 (N_16253,N_8784,N_10774);
nand U16254 (N_16254,N_6498,N_10183);
nand U16255 (N_16255,N_8975,N_9810);
nor U16256 (N_16256,N_8460,N_9959);
and U16257 (N_16257,N_10637,N_8633);
nor U16258 (N_16258,N_12146,N_11945);
nand U16259 (N_16259,N_8274,N_7265);
and U16260 (N_16260,N_10091,N_11152);
or U16261 (N_16261,N_10090,N_7096);
nor U16262 (N_16262,N_8659,N_10612);
nand U16263 (N_16263,N_6545,N_10875);
nand U16264 (N_16264,N_10230,N_6599);
nor U16265 (N_16265,N_6355,N_6259);
or U16266 (N_16266,N_10137,N_7360);
nand U16267 (N_16267,N_6631,N_8914);
nand U16268 (N_16268,N_9594,N_12063);
or U16269 (N_16269,N_7411,N_11114);
nor U16270 (N_16270,N_12131,N_7807);
nand U16271 (N_16271,N_11922,N_8191);
xnor U16272 (N_16272,N_10834,N_9887);
and U16273 (N_16273,N_7932,N_8498);
or U16274 (N_16274,N_8129,N_7046);
nand U16275 (N_16275,N_11619,N_8990);
xor U16276 (N_16276,N_11350,N_7802);
or U16277 (N_16277,N_11433,N_12208);
nor U16278 (N_16278,N_11748,N_7177);
nor U16279 (N_16279,N_11102,N_8037);
nand U16280 (N_16280,N_9574,N_6456);
or U16281 (N_16281,N_11613,N_8450);
nand U16282 (N_16282,N_8220,N_8245);
nor U16283 (N_16283,N_10607,N_8877);
nor U16284 (N_16284,N_12107,N_7735);
nand U16285 (N_16285,N_12373,N_10573);
and U16286 (N_16286,N_6591,N_12291);
nand U16287 (N_16287,N_12329,N_8514);
nand U16288 (N_16288,N_12030,N_7556);
nand U16289 (N_16289,N_10228,N_8473);
or U16290 (N_16290,N_11340,N_12322);
nand U16291 (N_16291,N_7720,N_9427);
and U16292 (N_16292,N_9372,N_6822);
nand U16293 (N_16293,N_12204,N_8720);
nand U16294 (N_16294,N_6487,N_10446);
nand U16295 (N_16295,N_7486,N_7590);
nand U16296 (N_16296,N_11575,N_9701);
nor U16297 (N_16297,N_9293,N_8597);
nor U16298 (N_16298,N_9483,N_9573);
and U16299 (N_16299,N_7846,N_12413);
and U16300 (N_16300,N_7390,N_9788);
or U16301 (N_16301,N_10846,N_11725);
nor U16302 (N_16302,N_6620,N_9939);
nand U16303 (N_16303,N_9120,N_8614);
and U16304 (N_16304,N_6455,N_6522);
or U16305 (N_16305,N_12204,N_9320);
or U16306 (N_16306,N_6927,N_6263);
nor U16307 (N_16307,N_7328,N_11138);
nand U16308 (N_16308,N_10955,N_9578);
xnor U16309 (N_16309,N_8156,N_9477);
or U16310 (N_16310,N_7504,N_8028);
nor U16311 (N_16311,N_12036,N_10012);
and U16312 (N_16312,N_9042,N_11613);
nor U16313 (N_16313,N_10471,N_7787);
and U16314 (N_16314,N_9782,N_7942);
and U16315 (N_16315,N_10243,N_9980);
nand U16316 (N_16316,N_9187,N_6675);
and U16317 (N_16317,N_7197,N_7838);
nor U16318 (N_16318,N_9071,N_7902);
or U16319 (N_16319,N_10473,N_12400);
or U16320 (N_16320,N_11098,N_6977);
or U16321 (N_16321,N_10694,N_8836);
and U16322 (N_16322,N_8115,N_6390);
xor U16323 (N_16323,N_10181,N_11840);
nor U16324 (N_16324,N_8038,N_12153);
or U16325 (N_16325,N_6560,N_7738);
nand U16326 (N_16326,N_9432,N_11042);
or U16327 (N_16327,N_6680,N_10258);
nor U16328 (N_16328,N_10355,N_7687);
or U16329 (N_16329,N_8138,N_9149);
nor U16330 (N_16330,N_6949,N_11934);
or U16331 (N_16331,N_11273,N_8626);
and U16332 (N_16332,N_7819,N_8235);
or U16333 (N_16333,N_8739,N_9696);
xor U16334 (N_16334,N_10680,N_12164);
or U16335 (N_16335,N_9162,N_11586);
and U16336 (N_16336,N_8994,N_10300);
or U16337 (N_16337,N_11087,N_6359);
and U16338 (N_16338,N_11187,N_11548);
or U16339 (N_16339,N_9556,N_11359);
or U16340 (N_16340,N_8658,N_6314);
or U16341 (N_16341,N_10451,N_6255);
and U16342 (N_16342,N_10147,N_7159);
and U16343 (N_16343,N_9002,N_7975);
and U16344 (N_16344,N_8532,N_10699);
and U16345 (N_16345,N_6778,N_8551);
nand U16346 (N_16346,N_9036,N_11832);
nand U16347 (N_16347,N_7259,N_10394);
or U16348 (N_16348,N_12202,N_9332);
nor U16349 (N_16349,N_10481,N_9122);
nand U16350 (N_16350,N_10410,N_10806);
and U16351 (N_16351,N_8520,N_10438);
or U16352 (N_16352,N_8607,N_10006);
nand U16353 (N_16353,N_7761,N_11459);
nor U16354 (N_16354,N_10571,N_9748);
nor U16355 (N_16355,N_9456,N_12344);
nand U16356 (N_16356,N_11029,N_9565);
and U16357 (N_16357,N_11722,N_6651);
nor U16358 (N_16358,N_7347,N_10541);
nor U16359 (N_16359,N_11721,N_10222);
xor U16360 (N_16360,N_11863,N_6255);
and U16361 (N_16361,N_10582,N_10082);
and U16362 (N_16362,N_12306,N_10524);
and U16363 (N_16363,N_6988,N_11141);
and U16364 (N_16364,N_10244,N_9170);
nand U16365 (N_16365,N_11513,N_8746);
xnor U16366 (N_16366,N_8047,N_10196);
nor U16367 (N_16367,N_7042,N_7988);
nor U16368 (N_16368,N_10485,N_12068);
nand U16369 (N_16369,N_11488,N_12296);
or U16370 (N_16370,N_11243,N_7309);
nand U16371 (N_16371,N_6446,N_11300);
xor U16372 (N_16372,N_8098,N_9895);
nand U16373 (N_16373,N_9016,N_6978);
and U16374 (N_16374,N_6505,N_8862);
or U16375 (N_16375,N_6767,N_12427);
xor U16376 (N_16376,N_10183,N_6598);
or U16377 (N_16377,N_8394,N_11971);
nor U16378 (N_16378,N_8942,N_11651);
xnor U16379 (N_16379,N_7478,N_12203);
nand U16380 (N_16380,N_10254,N_8776);
nor U16381 (N_16381,N_8164,N_7175);
xor U16382 (N_16382,N_8483,N_7018);
nand U16383 (N_16383,N_9883,N_12150);
nand U16384 (N_16384,N_11806,N_8754);
nor U16385 (N_16385,N_11364,N_8339);
nor U16386 (N_16386,N_7925,N_9923);
nand U16387 (N_16387,N_11642,N_9077);
and U16388 (N_16388,N_7076,N_8806);
nand U16389 (N_16389,N_9535,N_10367);
nor U16390 (N_16390,N_11667,N_8037);
nor U16391 (N_16391,N_9480,N_10154);
nor U16392 (N_16392,N_7620,N_9938);
and U16393 (N_16393,N_12390,N_11583);
nor U16394 (N_16394,N_11418,N_7129);
and U16395 (N_16395,N_8174,N_6929);
nand U16396 (N_16396,N_10696,N_8979);
and U16397 (N_16397,N_6801,N_8819);
and U16398 (N_16398,N_8371,N_11430);
and U16399 (N_16399,N_7649,N_11872);
and U16400 (N_16400,N_9513,N_10476);
or U16401 (N_16401,N_6855,N_11758);
xor U16402 (N_16402,N_8189,N_11250);
and U16403 (N_16403,N_10064,N_9866);
and U16404 (N_16404,N_6930,N_11475);
nor U16405 (N_16405,N_7069,N_8070);
xnor U16406 (N_16406,N_9308,N_11998);
or U16407 (N_16407,N_10460,N_11537);
nor U16408 (N_16408,N_6851,N_8689);
or U16409 (N_16409,N_10145,N_10360);
or U16410 (N_16410,N_12010,N_9154);
nor U16411 (N_16411,N_8017,N_6914);
and U16412 (N_16412,N_7332,N_8426);
and U16413 (N_16413,N_10306,N_10094);
and U16414 (N_16414,N_9301,N_10473);
nor U16415 (N_16415,N_7389,N_7043);
nand U16416 (N_16416,N_10088,N_6529);
xor U16417 (N_16417,N_7635,N_11262);
nand U16418 (N_16418,N_8298,N_7112);
and U16419 (N_16419,N_9492,N_11385);
and U16420 (N_16420,N_9531,N_9365);
nand U16421 (N_16421,N_10052,N_7035);
nand U16422 (N_16422,N_8917,N_9981);
or U16423 (N_16423,N_9509,N_7765);
and U16424 (N_16424,N_11588,N_10554);
and U16425 (N_16425,N_6451,N_8056);
nor U16426 (N_16426,N_8550,N_11419);
nand U16427 (N_16427,N_7054,N_9155);
nand U16428 (N_16428,N_7776,N_11347);
and U16429 (N_16429,N_8664,N_10942);
and U16430 (N_16430,N_6627,N_10962);
and U16431 (N_16431,N_11007,N_6521);
nor U16432 (N_16432,N_8062,N_10552);
nand U16433 (N_16433,N_10876,N_11063);
and U16434 (N_16434,N_9767,N_8388);
nor U16435 (N_16435,N_10269,N_9179);
nand U16436 (N_16436,N_7336,N_9816);
xor U16437 (N_16437,N_11033,N_9704);
nor U16438 (N_16438,N_7638,N_8396);
nor U16439 (N_16439,N_9300,N_7205);
xnor U16440 (N_16440,N_8845,N_7078);
nor U16441 (N_16441,N_10535,N_8898);
or U16442 (N_16442,N_6852,N_10735);
or U16443 (N_16443,N_11228,N_11624);
or U16444 (N_16444,N_9545,N_11955);
nor U16445 (N_16445,N_7154,N_11242);
or U16446 (N_16446,N_7470,N_11959);
nor U16447 (N_16447,N_6662,N_8558);
nor U16448 (N_16448,N_8353,N_7801);
or U16449 (N_16449,N_6313,N_8554);
nor U16450 (N_16450,N_9397,N_8123);
nand U16451 (N_16451,N_8256,N_6585);
nand U16452 (N_16452,N_10620,N_12212);
or U16453 (N_16453,N_6536,N_10054);
and U16454 (N_16454,N_8191,N_9472);
nor U16455 (N_16455,N_10431,N_9470);
or U16456 (N_16456,N_9506,N_9178);
nor U16457 (N_16457,N_12015,N_10173);
or U16458 (N_16458,N_9289,N_8986);
nand U16459 (N_16459,N_11001,N_9024);
and U16460 (N_16460,N_7157,N_9768);
xnor U16461 (N_16461,N_8084,N_7376);
xnor U16462 (N_16462,N_8238,N_11620);
or U16463 (N_16463,N_11548,N_11529);
and U16464 (N_16464,N_11248,N_9242);
or U16465 (N_16465,N_11964,N_9013);
nor U16466 (N_16466,N_12491,N_10487);
nand U16467 (N_16467,N_10854,N_9751);
and U16468 (N_16468,N_12498,N_12351);
and U16469 (N_16469,N_9629,N_6809);
nand U16470 (N_16470,N_10683,N_11795);
and U16471 (N_16471,N_12089,N_8278);
nand U16472 (N_16472,N_9332,N_7127);
nor U16473 (N_16473,N_9637,N_12073);
or U16474 (N_16474,N_12158,N_10228);
or U16475 (N_16475,N_7556,N_10597);
nand U16476 (N_16476,N_11296,N_10836);
and U16477 (N_16477,N_10984,N_8028);
and U16478 (N_16478,N_8609,N_7377);
nor U16479 (N_16479,N_9078,N_8278);
and U16480 (N_16480,N_11728,N_10774);
nand U16481 (N_16481,N_11274,N_12387);
and U16482 (N_16482,N_10383,N_6679);
or U16483 (N_16483,N_11722,N_7509);
or U16484 (N_16484,N_6502,N_9637);
and U16485 (N_16485,N_7412,N_7478);
nor U16486 (N_16486,N_6759,N_8013);
xor U16487 (N_16487,N_8024,N_11684);
and U16488 (N_16488,N_7023,N_7205);
or U16489 (N_16489,N_7304,N_8778);
nand U16490 (N_16490,N_12124,N_11407);
and U16491 (N_16491,N_10351,N_11634);
nand U16492 (N_16492,N_11995,N_9755);
nand U16493 (N_16493,N_12133,N_11800);
and U16494 (N_16494,N_10497,N_10985);
nand U16495 (N_16495,N_9709,N_9474);
and U16496 (N_16496,N_10279,N_11055);
nor U16497 (N_16497,N_6893,N_8093);
and U16498 (N_16498,N_7321,N_11710);
and U16499 (N_16499,N_11773,N_12499);
and U16500 (N_16500,N_11023,N_11171);
nand U16501 (N_16501,N_9592,N_11347);
and U16502 (N_16502,N_9477,N_9913);
and U16503 (N_16503,N_9401,N_11738);
nand U16504 (N_16504,N_8216,N_7946);
nor U16505 (N_16505,N_12306,N_11006);
nor U16506 (N_16506,N_8840,N_11436);
and U16507 (N_16507,N_7834,N_12211);
or U16508 (N_16508,N_10916,N_6817);
nor U16509 (N_16509,N_12041,N_7241);
nand U16510 (N_16510,N_11681,N_10762);
nor U16511 (N_16511,N_10052,N_6252);
xnor U16512 (N_16512,N_9123,N_9604);
nand U16513 (N_16513,N_6788,N_12123);
nand U16514 (N_16514,N_11855,N_6735);
and U16515 (N_16515,N_11808,N_6629);
xnor U16516 (N_16516,N_7604,N_7376);
or U16517 (N_16517,N_11128,N_11978);
xor U16518 (N_16518,N_8954,N_9439);
and U16519 (N_16519,N_6991,N_8498);
and U16520 (N_16520,N_11682,N_6866);
nor U16521 (N_16521,N_10802,N_10938);
nor U16522 (N_16522,N_8383,N_7724);
nand U16523 (N_16523,N_7643,N_11070);
and U16524 (N_16524,N_9128,N_8327);
xnor U16525 (N_16525,N_8870,N_12123);
nor U16526 (N_16526,N_11569,N_9857);
and U16527 (N_16527,N_11047,N_7056);
nor U16528 (N_16528,N_6262,N_6449);
or U16529 (N_16529,N_11838,N_11922);
or U16530 (N_16530,N_9617,N_11485);
or U16531 (N_16531,N_11363,N_6571);
and U16532 (N_16532,N_8424,N_8573);
or U16533 (N_16533,N_12179,N_10069);
nor U16534 (N_16534,N_7464,N_8701);
or U16535 (N_16535,N_11056,N_9827);
xnor U16536 (N_16536,N_10717,N_9458);
nand U16537 (N_16537,N_10655,N_12107);
or U16538 (N_16538,N_10968,N_11146);
or U16539 (N_16539,N_9380,N_8340);
and U16540 (N_16540,N_11822,N_6836);
or U16541 (N_16541,N_9490,N_7621);
or U16542 (N_16542,N_6479,N_8404);
and U16543 (N_16543,N_8057,N_9960);
or U16544 (N_16544,N_9304,N_6836);
nor U16545 (N_16545,N_10473,N_6612);
and U16546 (N_16546,N_11631,N_10384);
and U16547 (N_16547,N_11618,N_8547);
nand U16548 (N_16548,N_9587,N_8762);
nor U16549 (N_16549,N_7229,N_12497);
nand U16550 (N_16550,N_9196,N_10918);
nor U16551 (N_16551,N_11346,N_10262);
and U16552 (N_16552,N_9494,N_10323);
nor U16553 (N_16553,N_7537,N_8613);
and U16554 (N_16554,N_8854,N_11500);
nor U16555 (N_16555,N_7010,N_9650);
or U16556 (N_16556,N_9607,N_9969);
or U16557 (N_16557,N_9441,N_11686);
nor U16558 (N_16558,N_8658,N_9722);
nand U16559 (N_16559,N_7230,N_7181);
xnor U16560 (N_16560,N_11165,N_11688);
or U16561 (N_16561,N_11624,N_6599);
nand U16562 (N_16562,N_8452,N_8712);
nand U16563 (N_16563,N_10732,N_7439);
nand U16564 (N_16564,N_8780,N_6626);
xor U16565 (N_16565,N_8323,N_9596);
xor U16566 (N_16566,N_6757,N_8051);
or U16567 (N_16567,N_10392,N_11808);
and U16568 (N_16568,N_8490,N_8674);
nand U16569 (N_16569,N_6872,N_9224);
nand U16570 (N_16570,N_12243,N_7195);
xor U16571 (N_16571,N_6860,N_10661);
or U16572 (N_16572,N_10522,N_8756);
or U16573 (N_16573,N_7970,N_11434);
nand U16574 (N_16574,N_8064,N_11419);
nand U16575 (N_16575,N_7729,N_9676);
or U16576 (N_16576,N_10996,N_8518);
and U16577 (N_16577,N_7390,N_7871);
and U16578 (N_16578,N_9896,N_9494);
nand U16579 (N_16579,N_7572,N_6285);
and U16580 (N_16580,N_9448,N_8211);
or U16581 (N_16581,N_7536,N_9109);
and U16582 (N_16582,N_10642,N_8425);
xnor U16583 (N_16583,N_12453,N_9749);
and U16584 (N_16584,N_7437,N_7624);
and U16585 (N_16585,N_10232,N_12162);
and U16586 (N_16586,N_12192,N_10180);
and U16587 (N_16587,N_10871,N_7003);
nor U16588 (N_16588,N_8543,N_7052);
and U16589 (N_16589,N_11739,N_8017);
or U16590 (N_16590,N_9438,N_8483);
nand U16591 (N_16591,N_6944,N_11346);
nor U16592 (N_16592,N_6447,N_9425);
and U16593 (N_16593,N_6473,N_6650);
nor U16594 (N_16594,N_7599,N_7077);
and U16595 (N_16595,N_12207,N_6586);
nand U16596 (N_16596,N_6290,N_7116);
or U16597 (N_16597,N_6724,N_11697);
nand U16598 (N_16598,N_8493,N_12325);
and U16599 (N_16599,N_7743,N_12447);
nor U16600 (N_16600,N_11427,N_7240);
nand U16601 (N_16601,N_8381,N_8066);
and U16602 (N_16602,N_6829,N_7667);
or U16603 (N_16603,N_11537,N_7538);
xnor U16604 (N_16604,N_7290,N_8790);
nor U16605 (N_16605,N_11767,N_9904);
nor U16606 (N_16606,N_7098,N_10633);
nor U16607 (N_16607,N_9676,N_8083);
nand U16608 (N_16608,N_7310,N_11246);
nor U16609 (N_16609,N_9874,N_7502);
nand U16610 (N_16610,N_9193,N_7859);
nand U16611 (N_16611,N_9710,N_6905);
nor U16612 (N_16612,N_12141,N_8594);
nor U16613 (N_16613,N_10732,N_9421);
and U16614 (N_16614,N_9325,N_10584);
or U16615 (N_16615,N_12373,N_8474);
xor U16616 (N_16616,N_9134,N_10974);
or U16617 (N_16617,N_8540,N_9300);
xor U16618 (N_16618,N_7610,N_11272);
and U16619 (N_16619,N_9524,N_6705);
nor U16620 (N_16620,N_6518,N_11560);
or U16621 (N_16621,N_8641,N_10308);
nand U16622 (N_16622,N_9224,N_7721);
and U16623 (N_16623,N_6986,N_11954);
and U16624 (N_16624,N_8119,N_11608);
or U16625 (N_16625,N_10661,N_12341);
nand U16626 (N_16626,N_10440,N_11254);
nor U16627 (N_16627,N_10007,N_7813);
nand U16628 (N_16628,N_6332,N_12333);
nor U16629 (N_16629,N_9868,N_7993);
and U16630 (N_16630,N_7291,N_11039);
xor U16631 (N_16631,N_8154,N_12191);
nand U16632 (N_16632,N_12447,N_12437);
xnor U16633 (N_16633,N_9145,N_9126);
nand U16634 (N_16634,N_12452,N_11158);
and U16635 (N_16635,N_7788,N_8716);
and U16636 (N_16636,N_8259,N_10905);
or U16637 (N_16637,N_10625,N_7981);
nor U16638 (N_16638,N_8623,N_12404);
and U16639 (N_16639,N_6500,N_7475);
and U16640 (N_16640,N_8680,N_7544);
and U16641 (N_16641,N_9730,N_9403);
nand U16642 (N_16642,N_9330,N_8685);
or U16643 (N_16643,N_9077,N_11702);
xnor U16644 (N_16644,N_8934,N_9774);
xnor U16645 (N_16645,N_10204,N_9617);
nand U16646 (N_16646,N_6996,N_8587);
xor U16647 (N_16647,N_9743,N_7408);
and U16648 (N_16648,N_12301,N_7023);
nand U16649 (N_16649,N_10402,N_11813);
nor U16650 (N_16650,N_8323,N_6340);
nand U16651 (N_16651,N_11046,N_9317);
or U16652 (N_16652,N_9851,N_8801);
nand U16653 (N_16653,N_8913,N_9013);
nor U16654 (N_16654,N_12232,N_10211);
xnor U16655 (N_16655,N_8547,N_8620);
or U16656 (N_16656,N_11345,N_10471);
nand U16657 (N_16657,N_10507,N_6265);
nand U16658 (N_16658,N_7190,N_8866);
nand U16659 (N_16659,N_10634,N_10648);
nand U16660 (N_16660,N_12019,N_9016);
or U16661 (N_16661,N_7749,N_7915);
and U16662 (N_16662,N_7764,N_8864);
nand U16663 (N_16663,N_6809,N_11276);
nor U16664 (N_16664,N_11312,N_8053);
and U16665 (N_16665,N_9804,N_7558);
nor U16666 (N_16666,N_6676,N_9511);
and U16667 (N_16667,N_7326,N_7540);
and U16668 (N_16668,N_6408,N_12089);
nor U16669 (N_16669,N_11830,N_11428);
or U16670 (N_16670,N_11492,N_10169);
nand U16671 (N_16671,N_9238,N_8161);
or U16672 (N_16672,N_11238,N_7962);
or U16673 (N_16673,N_10451,N_11685);
or U16674 (N_16674,N_7886,N_11903);
xnor U16675 (N_16675,N_10920,N_10713);
nand U16676 (N_16676,N_7453,N_7121);
nor U16677 (N_16677,N_11977,N_12309);
nand U16678 (N_16678,N_11439,N_10017);
or U16679 (N_16679,N_11084,N_7991);
nor U16680 (N_16680,N_6824,N_12008);
xnor U16681 (N_16681,N_8365,N_7909);
or U16682 (N_16682,N_12261,N_7226);
nor U16683 (N_16683,N_11562,N_8931);
or U16684 (N_16684,N_11398,N_6912);
nor U16685 (N_16685,N_9689,N_9542);
nand U16686 (N_16686,N_10661,N_11195);
nor U16687 (N_16687,N_10476,N_10163);
or U16688 (N_16688,N_11345,N_12179);
xor U16689 (N_16689,N_10634,N_7555);
and U16690 (N_16690,N_9422,N_11892);
nor U16691 (N_16691,N_9738,N_6497);
nor U16692 (N_16692,N_12171,N_9224);
xnor U16693 (N_16693,N_7229,N_9423);
nand U16694 (N_16694,N_12481,N_9504);
nand U16695 (N_16695,N_6991,N_6688);
nand U16696 (N_16696,N_9139,N_7914);
and U16697 (N_16697,N_9993,N_10051);
nand U16698 (N_16698,N_7692,N_11704);
nand U16699 (N_16699,N_10281,N_12147);
nand U16700 (N_16700,N_10451,N_7148);
and U16701 (N_16701,N_12285,N_10417);
nand U16702 (N_16702,N_11616,N_6734);
nor U16703 (N_16703,N_6808,N_8502);
and U16704 (N_16704,N_9515,N_7448);
nor U16705 (N_16705,N_8371,N_8843);
nor U16706 (N_16706,N_7975,N_6709);
or U16707 (N_16707,N_9199,N_9302);
nor U16708 (N_16708,N_11332,N_8074);
and U16709 (N_16709,N_11799,N_8657);
nor U16710 (N_16710,N_7598,N_10901);
nand U16711 (N_16711,N_8415,N_8129);
nor U16712 (N_16712,N_7521,N_8793);
xnor U16713 (N_16713,N_11200,N_9852);
or U16714 (N_16714,N_9415,N_9054);
xor U16715 (N_16715,N_7407,N_8020);
nor U16716 (N_16716,N_11883,N_11431);
or U16717 (N_16717,N_6333,N_9551);
or U16718 (N_16718,N_8379,N_11243);
nor U16719 (N_16719,N_11625,N_9623);
and U16720 (N_16720,N_6913,N_10067);
or U16721 (N_16721,N_6571,N_10609);
xnor U16722 (N_16722,N_11247,N_11163);
and U16723 (N_16723,N_12419,N_7231);
nor U16724 (N_16724,N_8861,N_11781);
and U16725 (N_16725,N_8694,N_11491);
nor U16726 (N_16726,N_9785,N_7469);
xnor U16727 (N_16727,N_10489,N_8092);
and U16728 (N_16728,N_10331,N_6562);
or U16729 (N_16729,N_10434,N_8749);
nand U16730 (N_16730,N_6307,N_12487);
and U16731 (N_16731,N_7313,N_7766);
nor U16732 (N_16732,N_10358,N_8399);
or U16733 (N_16733,N_7651,N_8954);
or U16734 (N_16734,N_7996,N_8985);
nand U16735 (N_16735,N_10657,N_10694);
nand U16736 (N_16736,N_10805,N_10686);
and U16737 (N_16737,N_11909,N_10181);
nor U16738 (N_16738,N_6656,N_7151);
xnor U16739 (N_16739,N_11454,N_8404);
or U16740 (N_16740,N_10654,N_8317);
nand U16741 (N_16741,N_7009,N_11795);
nand U16742 (N_16742,N_6420,N_9444);
and U16743 (N_16743,N_10424,N_7202);
nand U16744 (N_16744,N_7571,N_9005);
xor U16745 (N_16745,N_10350,N_6665);
and U16746 (N_16746,N_10465,N_12025);
or U16747 (N_16747,N_9194,N_6391);
and U16748 (N_16748,N_6303,N_11425);
nor U16749 (N_16749,N_10569,N_7899);
nand U16750 (N_16750,N_10611,N_7443);
nor U16751 (N_16751,N_10162,N_11451);
or U16752 (N_16752,N_7537,N_7723);
nand U16753 (N_16753,N_8369,N_8453);
and U16754 (N_16754,N_6446,N_6864);
nor U16755 (N_16755,N_11605,N_10290);
or U16756 (N_16756,N_8047,N_8874);
nand U16757 (N_16757,N_11768,N_10435);
nand U16758 (N_16758,N_11694,N_7548);
or U16759 (N_16759,N_10317,N_6541);
nand U16760 (N_16760,N_6934,N_12031);
or U16761 (N_16761,N_7196,N_7130);
and U16762 (N_16762,N_7330,N_11094);
and U16763 (N_16763,N_10476,N_9305);
nor U16764 (N_16764,N_6387,N_8906);
or U16765 (N_16765,N_8847,N_7822);
nor U16766 (N_16766,N_9882,N_11563);
or U16767 (N_16767,N_11119,N_12038);
or U16768 (N_16768,N_9292,N_7303);
nor U16769 (N_16769,N_10212,N_11432);
nand U16770 (N_16770,N_11290,N_8023);
or U16771 (N_16771,N_8609,N_10604);
nor U16772 (N_16772,N_10828,N_8694);
nor U16773 (N_16773,N_6878,N_7490);
nor U16774 (N_16774,N_10539,N_7613);
nor U16775 (N_16775,N_9368,N_12315);
nand U16776 (N_16776,N_8014,N_11920);
or U16777 (N_16777,N_7932,N_8097);
xnor U16778 (N_16778,N_11554,N_11944);
nor U16779 (N_16779,N_6898,N_10084);
nand U16780 (N_16780,N_7449,N_10112);
nand U16781 (N_16781,N_8899,N_8864);
nor U16782 (N_16782,N_6555,N_9217);
nor U16783 (N_16783,N_11372,N_7572);
and U16784 (N_16784,N_11440,N_10951);
nand U16785 (N_16785,N_10064,N_6998);
and U16786 (N_16786,N_10391,N_7318);
or U16787 (N_16787,N_11598,N_10051);
nand U16788 (N_16788,N_8230,N_11590);
or U16789 (N_16789,N_10398,N_8982);
nand U16790 (N_16790,N_7412,N_11957);
nor U16791 (N_16791,N_9575,N_6451);
nand U16792 (N_16792,N_9115,N_10384);
nor U16793 (N_16793,N_10608,N_9738);
nor U16794 (N_16794,N_12280,N_10226);
nand U16795 (N_16795,N_6320,N_6694);
nor U16796 (N_16796,N_11357,N_10892);
or U16797 (N_16797,N_6700,N_11787);
and U16798 (N_16798,N_10658,N_11006);
nor U16799 (N_16799,N_8115,N_12027);
and U16800 (N_16800,N_10272,N_8484);
nor U16801 (N_16801,N_12238,N_6640);
or U16802 (N_16802,N_10100,N_8549);
nand U16803 (N_16803,N_9326,N_7686);
nor U16804 (N_16804,N_8576,N_11250);
or U16805 (N_16805,N_11918,N_6815);
and U16806 (N_16806,N_12338,N_6330);
and U16807 (N_16807,N_7341,N_6277);
nand U16808 (N_16808,N_6399,N_11998);
nor U16809 (N_16809,N_9259,N_11054);
and U16810 (N_16810,N_7834,N_12449);
or U16811 (N_16811,N_7457,N_11592);
nand U16812 (N_16812,N_10868,N_8569);
and U16813 (N_16813,N_6483,N_12490);
nor U16814 (N_16814,N_7041,N_10741);
or U16815 (N_16815,N_11978,N_8615);
or U16816 (N_16816,N_7986,N_7477);
and U16817 (N_16817,N_11973,N_10428);
and U16818 (N_16818,N_8608,N_11568);
and U16819 (N_16819,N_10011,N_7661);
and U16820 (N_16820,N_7572,N_8938);
and U16821 (N_16821,N_9494,N_9759);
and U16822 (N_16822,N_11679,N_9855);
xnor U16823 (N_16823,N_6309,N_10058);
and U16824 (N_16824,N_9907,N_11513);
nand U16825 (N_16825,N_10127,N_8338);
nor U16826 (N_16826,N_10754,N_7652);
or U16827 (N_16827,N_11967,N_10136);
and U16828 (N_16828,N_6768,N_8096);
xnor U16829 (N_16829,N_7541,N_8960);
xnor U16830 (N_16830,N_7791,N_11393);
nor U16831 (N_16831,N_6813,N_11541);
nand U16832 (N_16832,N_8546,N_12206);
nand U16833 (N_16833,N_8659,N_9568);
nand U16834 (N_16834,N_11748,N_12173);
nand U16835 (N_16835,N_12335,N_8673);
nand U16836 (N_16836,N_8517,N_11501);
or U16837 (N_16837,N_7339,N_8676);
nor U16838 (N_16838,N_7698,N_11575);
nor U16839 (N_16839,N_10040,N_8689);
nor U16840 (N_16840,N_9492,N_10954);
or U16841 (N_16841,N_9573,N_10356);
xnor U16842 (N_16842,N_6536,N_7089);
xor U16843 (N_16843,N_6899,N_8363);
nor U16844 (N_16844,N_10872,N_9532);
xnor U16845 (N_16845,N_9348,N_12447);
or U16846 (N_16846,N_10220,N_9490);
and U16847 (N_16847,N_9599,N_7033);
nor U16848 (N_16848,N_8492,N_11882);
or U16849 (N_16849,N_7951,N_10827);
nor U16850 (N_16850,N_9717,N_10479);
nor U16851 (N_16851,N_10196,N_8460);
nor U16852 (N_16852,N_6973,N_9242);
xnor U16853 (N_16853,N_8826,N_10328);
nor U16854 (N_16854,N_10327,N_9106);
and U16855 (N_16855,N_7163,N_7553);
nand U16856 (N_16856,N_11228,N_6722);
or U16857 (N_16857,N_9395,N_10205);
or U16858 (N_16858,N_6784,N_8337);
or U16859 (N_16859,N_9440,N_6790);
and U16860 (N_16860,N_9087,N_10908);
nand U16861 (N_16861,N_8895,N_7199);
nand U16862 (N_16862,N_11880,N_7169);
nor U16863 (N_16863,N_9015,N_6557);
or U16864 (N_16864,N_10698,N_8156);
and U16865 (N_16865,N_7330,N_11574);
nand U16866 (N_16866,N_9359,N_7639);
and U16867 (N_16867,N_8194,N_8605);
nand U16868 (N_16868,N_8081,N_9362);
and U16869 (N_16869,N_8722,N_10848);
nand U16870 (N_16870,N_9537,N_8945);
nand U16871 (N_16871,N_10020,N_7943);
and U16872 (N_16872,N_10104,N_11453);
nor U16873 (N_16873,N_6886,N_11564);
or U16874 (N_16874,N_11354,N_7937);
nor U16875 (N_16875,N_9025,N_8202);
nor U16876 (N_16876,N_11147,N_11049);
or U16877 (N_16877,N_7884,N_12417);
nand U16878 (N_16878,N_6931,N_7348);
and U16879 (N_16879,N_6289,N_10805);
or U16880 (N_16880,N_7813,N_6635);
nand U16881 (N_16881,N_12000,N_10778);
nand U16882 (N_16882,N_12428,N_8686);
or U16883 (N_16883,N_9748,N_10120);
nor U16884 (N_16884,N_9174,N_7523);
or U16885 (N_16885,N_6458,N_9720);
and U16886 (N_16886,N_8244,N_6824);
nor U16887 (N_16887,N_10329,N_8864);
xnor U16888 (N_16888,N_9278,N_10771);
nand U16889 (N_16889,N_9477,N_9222);
nor U16890 (N_16890,N_7043,N_7001);
and U16891 (N_16891,N_6712,N_12018);
nor U16892 (N_16892,N_10362,N_11795);
and U16893 (N_16893,N_9020,N_11433);
and U16894 (N_16894,N_6887,N_9673);
nor U16895 (N_16895,N_12253,N_10620);
and U16896 (N_16896,N_9417,N_10010);
nor U16897 (N_16897,N_11808,N_10652);
xnor U16898 (N_16898,N_7932,N_6380);
and U16899 (N_16899,N_8785,N_8188);
nor U16900 (N_16900,N_11008,N_7903);
and U16901 (N_16901,N_9609,N_11365);
nor U16902 (N_16902,N_11546,N_10009);
nand U16903 (N_16903,N_10374,N_11925);
and U16904 (N_16904,N_6258,N_11854);
nand U16905 (N_16905,N_8405,N_7760);
and U16906 (N_16906,N_9868,N_11351);
nand U16907 (N_16907,N_7804,N_7805);
or U16908 (N_16908,N_10958,N_6957);
and U16909 (N_16909,N_10374,N_12163);
and U16910 (N_16910,N_10644,N_6511);
or U16911 (N_16911,N_11705,N_8175);
or U16912 (N_16912,N_8673,N_7466);
or U16913 (N_16913,N_9367,N_8228);
and U16914 (N_16914,N_10411,N_10427);
and U16915 (N_16915,N_9601,N_10610);
and U16916 (N_16916,N_9071,N_6406);
nand U16917 (N_16917,N_7877,N_11459);
nand U16918 (N_16918,N_11195,N_11132);
xor U16919 (N_16919,N_9003,N_7485);
or U16920 (N_16920,N_9556,N_9891);
nand U16921 (N_16921,N_10783,N_7351);
xnor U16922 (N_16922,N_7221,N_10588);
and U16923 (N_16923,N_11147,N_12286);
nand U16924 (N_16924,N_9159,N_11776);
xor U16925 (N_16925,N_6557,N_7015);
nand U16926 (N_16926,N_7746,N_7981);
nand U16927 (N_16927,N_8803,N_10385);
nand U16928 (N_16928,N_8788,N_11116);
nand U16929 (N_16929,N_8611,N_9292);
nand U16930 (N_16930,N_9531,N_7479);
or U16931 (N_16931,N_7060,N_11782);
nor U16932 (N_16932,N_7981,N_8968);
nand U16933 (N_16933,N_11626,N_10721);
xnor U16934 (N_16934,N_8522,N_11306);
nand U16935 (N_16935,N_11633,N_7106);
nand U16936 (N_16936,N_11069,N_12139);
or U16937 (N_16937,N_9173,N_9895);
or U16938 (N_16938,N_12018,N_7232);
nor U16939 (N_16939,N_7795,N_12497);
nor U16940 (N_16940,N_7048,N_7373);
nor U16941 (N_16941,N_11677,N_6575);
or U16942 (N_16942,N_11870,N_7605);
or U16943 (N_16943,N_11623,N_6791);
and U16944 (N_16944,N_12408,N_7765);
and U16945 (N_16945,N_11361,N_7090);
xor U16946 (N_16946,N_11948,N_10301);
nor U16947 (N_16947,N_9652,N_12332);
or U16948 (N_16948,N_11200,N_11981);
nand U16949 (N_16949,N_12166,N_8201);
nand U16950 (N_16950,N_7093,N_11606);
or U16951 (N_16951,N_8599,N_10733);
and U16952 (N_16952,N_9053,N_10717);
nor U16953 (N_16953,N_10763,N_7566);
nor U16954 (N_16954,N_8047,N_11996);
nand U16955 (N_16955,N_7421,N_7746);
or U16956 (N_16956,N_10507,N_7869);
nor U16957 (N_16957,N_7958,N_8479);
or U16958 (N_16958,N_7300,N_9332);
and U16959 (N_16959,N_7927,N_6616);
nor U16960 (N_16960,N_9779,N_7209);
or U16961 (N_16961,N_7762,N_12013);
or U16962 (N_16962,N_10289,N_6573);
nand U16963 (N_16963,N_9520,N_7051);
nand U16964 (N_16964,N_11681,N_10913);
and U16965 (N_16965,N_7250,N_9808);
nand U16966 (N_16966,N_6697,N_8696);
and U16967 (N_16967,N_10740,N_8827);
or U16968 (N_16968,N_7113,N_11864);
nor U16969 (N_16969,N_10725,N_11051);
nand U16970 (N_16970,N_9993,N_7862);
nor U16971 (N_16971,N_11819,N_7774);
or U16972 (N_16972,N_7532,N_7370);
nor U16973 (N_16973,N_8354,N_6729);
nand U16974 (N_16974,N_9594,N_11165);
and U16975 (N_16975,N_9893,N_9236);
or U16976 (N_16976,N_10522,N_10987);
nor U16977 (N_16977,N_12300,N_10504);
or U16978 (N_16978,N_6708,N_12103);
nand U16979 (N_16979,N_11428,N_10435);
or U16980 (N_16980,N_8780,N_8356);
or U16981 (N_16981,N_9570,N_9878);
nor U16982 (N_16982,N_6973,N_9646);
and U16983 (N_16983,N_11487,N_11950);
nor U16984 (N_16984,N_8287,N_9019);
or U16985 (N_16985,N_6576,N_10395);
and U16986 (N_16986,N_12034,N_10662);
or U16987 (N_16987,N_12277,N_7760);
nand U16988 (N_16988,N_10900,N_10501);
xor U16989 (N_16989,N_9829,N_11115);
and U16990 (N_16990,N_11612,N_7155);
and U16991 (N_16991,N_6594,N_9396);
nand U16992 (N_16992,N_10650,N_11348);
and U16993 (N_16993,N_9796,N_11640);
nand U16994 (N_16994,N_9146,N_9268);
or U16995 (N_16995,N_9475,N_7793);
xor U16996 (N_16996,N_8064,N_11993);
or U16997 (N_16997,N_11253,N_6271);
nand U16998 (N_16998,N_11509,N_11866);
or U16999 (N_16999,N_8380,N_7966);
xor U17000 (N_17000,N_9474,N_7199);
nand U17001 (N_17001,N_9729,N_7307);
nor U17002 (N_17002,N_10123,N_9132);
or U17003 (N_17003,N_11403,N_9479);
and U17004 (N_17004,N_9737,N_11605);
and U17005 (N_17005,N_9914,N_11509);
nor U17006 (N_17006,N_8425,N_10441);
or U17007 (N_17007,N_6823,N_9647);
or U17008 (N_17008,N_8559,N_10165);
nand U17009 (N_17009,N_11326,N_11699);
and U17010 (N_17010,N_12297,N_11002);
nor U17011 (N_17011,N_10665,N_9226);
and U17012 (N_17012,N_9291,N_7913);
nor U17013 (N_17013,N_11884,N_9242);
and U17014 (N_17014,N_6935,N_7298);
xor U17015 (N_17015,N_6935,N_8096);
nand U17016 (N_17016,N_12164,N_8167);
and U17017 (N_17017,N_8995,N_9929);
nor U17018 (N_17018,N_12108,N_8636);
or U17019 (N_17019,N_11032,N_8137);
or U17020 (N_17020,N_8131,N_8270);
and U17021 (N_17021,N_9977,N_8333);
or U17022 (N_17022,N_6804,N_8862);
nor U17023 (N_17023,N_12442,N_10356);
nand U17024 (N_17024,N_8868,N_7443);
and U17025 (N_17025,N_8163,N_6776);
and U17026 (N_17026,N_12327,N_10723);
nor U17027 (N_17027,N_7030,N_12463);
or U17028 (N_17028,N_11558,N_11352);
and U17029 (N_17029,N_7143,N_11252);
nand U17030 (N_17030,N_6447,N_11647);
xnor U17031 (N_17031,N_10891,N_6910);
nand U17032 (N_17032,N_9183,N_11414);
nand U17033 (N_17033,N_9307,N_6639);
xor U17034 (N_17034,N_11805,N_6405);
or U17035 (N_17035,N_7334,N_9148);
xor U17036 (N_17036,N_11332,N_6977);
nor U17037 (N_17037,N_6977,N_9785);
xor U17038 (N_17038,N_7943,N_11333);
nor U17039 (N_17039,N_10196,N_8403);
nand U17040 (N_17040,N_7086,N_12283);
nand U17041 (N_17041,N_10368,N_8650);
nand U17042 (N_17042,N_11847,N_11638);
nor U17043 (N_17043,N_8936,N_10412);
nand U17044 (N_17044,N_10765,N_9000);
or U17045 (N_17045,N_9550,N_11847);
or U17046 (N_17046,N_10244,N_6276);
nor U17047 (N_17047,N_8311,N_10006);
nor U17048 (N_17048,N_8960,N_11538);
or U17049 (N_17049,N_10063,N_12047);
nor U17050 (N_17050,N_7144,N_12227);
and U17051 (N_17051,N_8406,N_7212);
nor U17052 (N_17052,N_9430,N_6850);
xnor U17053 (N_17053,N_10533,N_6291);
nand U17054 (N_17054,N_10069,N_10383);
nor U17055 (N_17055,N_10253,N_6896);
nor U17056 (N_17056,N_8226,N_7475);
or U17057 (N_17057,N_10362,N_9805);
nor U17058 (N_17058,N_12094,N_6704);
xor U17059 (N_17059,N_12413,N_12400);
and U17060 (N_17060,N_11990,N_8917);
or U17061 (N_17061,N_10138,N_9608);
nand U17062 (N_17062,N_6812,N_9725);
nor U17063 (N_17063,N_8734,N_10914);
and U17064 (N_17064,N_12426,N_7719);
nand U17065 (N_17065,N_9963,N_11261);
nor U17066 (N_17066,N_12292,N_8432);
nor U17067 (N_17067,N_11749,N_6402);
nand U17068 (N_17068,N_10213,N_8142);
nor U17069 (N_17069,N_9439,N_6577);
nor U17070 (N_17070,N_11442,N_11008);
nand U17071 (N_17071,N_9326,N_12086);
or U17072 (N_17072,N_6704,N_12045);
or U17073 (N_17073,N_8026,N_7526);
and U17074 (N_17074,N_8421,N_8007);
or U17075 (N_17075,N_10474,N_6741);
nand U17076 (N_17076,N_12062,N_12137);
nor U17077 (N_17077,N_12166,N_8416);
or U17078 (N_17078,N_9329,N_7780);
or U17079 (N_17079,N_7258,N_8425);
nor U17080 (N_17080,N_8082,N_8276);
xor U17081 (N_17081,N_7443,N_7095);
or U17082 (N_17082,N_6282,N_12187);
nor U17083 (N_17083,N_11612,N_11219);
nor U17084 (N_17084,N_9373,N_9078);
and U17085 (N_17085,N_10758,N_8189);
or U17086 (N_17086,N_10977,N_6379);
or U17087 (N_17087,N_12488,N_9753);
nand U17088 (N_17088,N_12345,N_7193);
nor U17089 (N_17089,N_11953,N_7750);
nand U17090 (N_17090,N_10304,N_11470);
nor U17091 (N_17091,N_7830,N_12275);
xnor U17092 (N_17092,N_8819,N_10858);
nor U17093 (N_17093,N_8884,N_7483);
or U17094 (N_17094,N_7604,N_8129);
nor U17095 (N_17095,N_9070,N_12258);
and U17096 (N_17096,N_12485,N_9930);
nand U17097 (N_17097,N_8967,N_9987);
nand U17098 (N_17098,N_10096,N_11097);
and U17099 (N_17099,N_12227,N_12263);
xnor U17100 (N_17100,N_10704,N_9680);
xnor U17101 (N_17101,N_8078,N_6762);
nor U17102 (N_17102,N_8153,N_6931);
xnor U17103 (N_17103,N_10624,N_8642);
nor U17104 (N_17104,N_8089,N_12054);
and U17105 (N_17105,N_10413,N_8934);
or U17106 (N_17106,N_10654,N_6653);
and U17107 (N_17107,N_12488,N_12404);
nor U17108 (N_17108,N_6902,N_11277);
xor U17109 (N_17109,N_6924,N_6515);
nor U17110 (N_17110,N_9208,N_8011);
and U17111 (N_17111,N_6339,N_8136);
nand U17112 (N_17112,N_12410,N_8444);
xor U17113 (N_17113,N_8767,N_12357);
nand U17114 (N_17114,N_8479,N_9222);
or U17115 (N_17115,N_10300,N_10469);
and U17116 (N_17116,N_6891,N_7834);
nor U17117 (N_17117,N_10620,N_7913);
nor U17118 (N_17118,N_6399,N_6624);
and U17119 (N_17119,N_8599,N_11540);
and U17120 (N_17120,N_10309,N_9578);
or U17121 (N_17121,N_11676,N_9949);
xnor U17122 (N_17122,N_9144,N_10690);
nand U17123 (N_17123,N_7914,N_7418);
xor U17124 (N_17124,N_11202,N_11360);
or U17125 (N_17125,N_7412,N_10564);
nand U17126 (N_17126,N_8084,N_10176);
or U17127 (N_17127,N_7134,N_9305);
nor U17128 (N_17128,N_8327,N_8383);
xor U17129 (N_17129,N_11272,N_8200);
xnor U17130 (N_17130,N_7598,N_11877);
or U17131 (N_17131,N_11402,N_9444);
or U17132 (N_17132,N_8134,N_11872);
xor U17133 (N_17133,N_9763,N_7304);
nand U17134 (N_17134,N_7557,N_10809);
and U17135 (N_17135,N_6585,N_12372);
nor U17136 (N_17136,N_9992,N_10946);
nand U17137 (N_17137,N_10595,N_11274);
nand U17138 (N_17138,N_8909,N_8147);
nor U17139 (N_17139,N_10768,N_11633);
or U17140 (N_17140,N_12179,N_9892);
and U17141 (N_17141,N_11589,N_8369);
and U17142 (N_17142,N_11400,N_6353);
and U17143 (N_17143,N_8769,N_9170);
nand U17144 (N_17144,N_7204,N_8075);
and U17145 (N_17145,N_7213,N_9949);
and U17146 (N_17146,N_12024,N_10083);
and U17147 (N_17147,N_10813,N_7111);
nor U17148 (N_17148,N_11435,N_9999);
and U17149 (N_17149,N_7829,N_10858);
nor U17150 (N_17150,N_6733,N_10804);
xor U17151 (N_17151,N_10982,N_9123);
or U17152 (N_17152,N_6764,N_7277);
nand U17153 (N_17153,N_10185,N_9340);
or U17154 (N_17154,N_8010,N_10578);
or U17155 (N_17155,N_7300,N_12461);
or U17156 (N_17156,N_7040,N_6791);
nor U17157 (N_17157,N_10986,N_7967);
and U17158 (N_17158,N_12274,N_6342);
nand U17159 (N_17159,N_6546,N_10932);
and U17160 (N_17160,N_7262,N_8966);
nand U17161 (N_17161,N_11450,N_12061);
and U17162 (N_17162,N_7422,N_11646);
and U17163 (N_17163,N_8255,N_11448);
or U17164 (N_17164,N_7107,N_9586);
xnor U17165 (N_17165,N_7200,N_11212);
nand U17166 (N_17166,N_11101,N_7220);
xor U17167 (N_17167,N_6857,N_9783);
or U17168 (N_17168,N_6443,N_6349);
nand U17169 (N_17169,N_6808,N_11772);
and U17170 (N_17170,N_8656,N_10127);
xnor U17171 (N_17171,N_9618,N_12262);
nor U17172 (N_17172,N_11309,N_8856);
nand U17173 (N_17173,N_8147,N_9782);
or U17174 (N_17174,N_9672,N_11571);
nand U17175 (N_17175,N_9406,N_6736);
nand U17176 (N_17176,N_8639,N_7288);
nand U17177 (N_17177,N_10988,N_10708);
and U17178 (N_17178,N_8977,N_11886);
and U17179 (N_17179,N_11181,N_7195);
and U17180 (N_17180,N_10506,N_7736);
or U17181 (N_17181,N_9387,N_10394);
or U17182 (N_17182,N_9730,N_6333);
nand U17183 (N_17183,N_9240,N_7030);
and U17184 (N_17184,N_7228,N_12214);
nand U17185 (N_17185,N_11709,N_11947);
and U17186 (N_17186,N_11993,N_7704);
nor U17187 (N_17187,N_10115,N_7926);
and U17188 (N_17188,N_10741,N_11225);
and U17189 (N_17189,N_6554,N_8122);
and U17190 (N_17190,N_9305,N_6979);
nand U17191 (N_17191,N_12427,N_10871);
and U17192 (N_17192,N_11583,N_8202);
nor U17193 (N_17193,N_10723,N_7908);
nand U17194 (N_17194,N_8342,N_6956);
nand U17195 (N_17195,N_8729,N_9972);
nand U17196 (N_17196,N_10354,N_10228);
nand U17197 (N_17197,N_8426,N_6792);
or U17198 (N_17198,N_6258,N_9317);
nor U17199 (N_17199,N_7332,N_6946);
nor U17200 (N_17200,N_7150,N_10986);
nand U17201 (N_17201,N_10013,N_8913);
nand U17202 (N_17202,N_8455,N_9525);
nand U17203 (N_17203,N_11545,N_8639);
xnor U17204 (N_17204,N_7661,N_11192);
and U17205 (N_17205,N_12148,N_11663);
nor U17206 (N_17206,N_8636,N_9585);
nand U17207 (N_17207,N_7451,N_11997);
nor U17208 (N_17208,N_9911,N_11009);
or U17209 (N_17209,N_6994,N_9859);
nor U17210 (N_17210,N_7058,N_8167);
and U17211 (N_17211,N_10534,N_9251);
or U17212 (N_17212,N_11332,N_11997);
and U17213 (N_17213,N_10575,N_8069);
or U17214 (N_17214,N_11790,N_6593);
and U17215 (N_17215,N_11709,N_12204);
nand U17216 (N_17216,N_8658,N_7493);
or U17217 (N_17217,N_9760,N_7843);
and U17218 (N_17218,N_8176,N_11282);
or U17219 (N_17219,N_6632,N_6609);
nor U17220 (N_17220,N_9239,N_7593);
nor U17221 (N_17221,N_10373,N_12215);
or U17222 (N_17222,N_10843,N_9460);
nand U17223 (N_17223,N_10050,N_11484);
nand U17224 (N_17224,N_10836,N_9920);
and U17225 (N_17225,N_9662,N_6279);
and U17226 (N_17226,N_8144,N_8578);
nor U17227 (N_17227,N_9568,N_10621);
nand U17228 (N_17228,N_9682,N_10903);
xnor U17229 (N_17229,N_9166,N_6952);
and U17230 (N_17230,N_8005,N_11988);
and U17231 (N_17231,N_11622,N_8741);
nand U17232 (N_17232,N_8359,N_9564);
and U17233 (N_17233,N_11627,N_8302);
nand U17234 (N_17234,N_7878,N_7354);
nor U17235 (N_17235,N_10819,N_11801);
and U17236 (N_17236,N_11709,N_8431);
and U17237 (N_17237,N_11238,N_12133);
nor U17238 (N_17238,N_7299,N_11994);
or U17239 (N_17239,N_6672,N_10772);
nand U17240 (N_17240,N_12205,N_11343);
nor U17241 (N_17241,N_10690,N_6746);
and U17242 (N_17242,N_12478,N_11348);
nand U17243 (N_17243,N_8101,N_7841);
or U17244 (N_17244,N_7717,N_11172);
xnor U17245 (N_17245,N_12404,N_11907);
nand U17246 (N_17246,N_9946,N_12440);
and U17247 (N_17247,N_6785,N_9498);
or U17248 (N_17248,N_7796,N_10193);
and U17249 (N_17249,N_11751,N_12207);
nor U17250 (N_17250,N_11605,N_12422);
and U17251 (N_17251,N_10158,N_12032);
nor U17252 (N_17252,N_11676,N_10297);
nor U17253 (N_17253,N_9065,N_8309);
and U17254 (N_17254,N_11512,N_8495);
and U17255 (N_17255,N_10295,N_7683);
or U17256 (N_17256,N_6700,N_6664);
nor U17257 (N_17257,N_8251,N_9358);
or U17258 (N_17258,N_10629,N_8869);
nor U17259 (N_17259,N_11944,N_7900);
or U17260 (N_17260,N_6311,N_12283);
nand U17261 (N_17261,N_8387,N_10391);
nand U17262 (N_17262,N_6324,N_8778);
nand U17263 (N_17263,N_6975,N_6771);
nand U17264 (N_17264,N_11718,N_9575);
nand U17265 (N_17265,N_10457,N_11522);
nor U17266 (N_17266,N_9560,N_10458);
nand U17267 (N_17267,N_10489,N_6306);
xnor U17268 (N_17268,N_12462,N_8737);
and U17269 (N_17269,N_11845,N_12479);
or U17270 (N_17270,N_11785,N_10730);
nor U17271 (N_17271,N_8805,N_12072);
xnor U17272 (N_17272,N_11701,N_9546);
nand U17273 (N_17273,N_7523,N_11333);
xnor U17274 (N_17274,N_8986,N_11889);
and U17275 (N_17275,N_8042,N_9371);
nand U17276 (N_17276,N_10919,N_6819);
and U17277 (N_17277,N_7253,N_7038);
nor U17278 (N_17278,N_9118,N_6806);
and U17279 (N_17279,N_8341,N_11235);
nand U17280 (N_17280,N_10799,N_10029);
or U17281 (N_17281,N_11351,N_6481);
xnor U17282 (N_17282,N_11569,N_8598);
or U17283 (N_17283,N_8859,N_10851);
xnor U17284 (N_17284,N_11618,N_10169);
nand U17285 (N_17285,N_9912,N_7160);
xor U17286 (N_17286,N_6485,N_6705);
or U17287 (N_17287,N_9658,N_6516);
nor U17288 (N_17288,N_7545,N_8142);
nor U17289 (N_17289,N_7635,N_11718);
or U17290 (N_17290,N_12313,N_10913);
and U17291 (N_17291,N_9621,N_7226);
nand U17292 (N_17292,N_9891,N_8104);
and U17293 (N_17293,N_10370,N_11915);
nand U17294 (N_17294,N_7266,N_11832);
xor U17295 (N_17295,N_8202,N_7264);
and U17296 (N_17296,N_6928,N_10470);
nor U17297 (N_17297,N_11170,N_10044);
nor U17298 (N_17298,N_9111,N_11893);
and U17299 (N_17299,N_8975,N_6558);
xnor U17300 (N_17300,N_8713,N_12438);
and U17301 (N_17301,N_7668,N_7629);
nor U17302 (N_17302,N_8267,N_7880);
nor U17303 (N_17303,N_6665,N_7138);
and U17304 (N_17304,N_11132,N_12039);
and U17305 (N_17305,N_12197,N_7818);
and U17306 (N_17306,N_8650,N_8911);
nand U17307 (N_17307,N_6530,N_8708);
or U17308 (N_17308,N_6964,N_11421);
or U17309 (N_17309,N_12075,N_8325);
nor U17310 (N_17310,N_11009,N_6519);
xor U17311 (N_17311,N_10498,N_10279);
and U17312 (N_17312,N_12104,N_11392);
nand U17313 (N_17313,N_11235,N_6364);
nand U17314 (N_17314,N_6841,N_7352);
and U17315 (N_17315,N_8202,N_10429);
nand U17316 (N_17316,N_6963,N_12145);
nor U17317 (N_17317,N_8392,N_11728);
and U17318 (N_17318,N_11372,N_7485);
or U17319 (N_17319,N_6769,N_10702);
xnor U17320 (N_17320,N_6583,N_6734);
and U17321 (N_17321,N_7949,N_10354);
nand U17322 (N_17322,N_7588,N_12160);
xor U17323 (N_17323,N_8140,N_7663);
and U17324 (N_17324,N_9976,N_11797);
or U17325 (N_17325,N_6700,N_11120);
or U17326 (N_17326,N_7665,N_12388);
nand U17327 (N_17327,N_11560,N_11184);
nand U17328 (N_17328,N_8947,N_11548);
or U17329 (N_17329,N_12167,N_10773);
nor U17330 (N_17330,N_12285,N_10591);
nand U17331 (N_17331,N_11777,N_12356);
nor U17332 (N_17332,N_11962,N_6858);
or U17333 (N_17333,N_7043,N_9171);
nor U17334 (N_17334,N_10561,N_7634);
xor U17335 (N_17335,N_8267,N_11605);
xor U17336 (N_17336,N_8159,N_7239);
or U17337 (N_17337,N_8486,N_7207);
nand U17338 (N_17338,N_8396,N_10667);
nand U17339 (N_17339,N_11171,N_12277);
and U17340 (N_17340,N_9195,N_7749);
and U17341 (N_17341,N_11406,N_6662);
or U17342 (N_17342,N_11826,N_7905);
nand U17343 (N_17343,N_7230,N_9717);
or U17344 (N_17344,N_9099,N_8685);
and U17345 (N_17345,N_11371,N_10210);
xnor U17346 (N_17346,N_7224,N_12113);
nor U17347 (N_17347,N_7523,N_7881);
and U17348 (N_17348,N_8133,N_11027);
nor U17349 (N_17349,N_8289,N_9521);
nor U17350 (N_17350,N_7253,N_6991);
nand U17351 (N_17351,N_10007,N_8392);
and U17352 (N_17352,N_6599,N_10513);
or U17353 (N_17353,N_6894,N_11283);
or U17354 (N_17354,N_11989,N_10493);
nor U17355 (N_17355,N_12405,N_10222);
and U17356 (N_17356,N_10518,N_8719);
and U17357 (N_17357,N_10540,N_8678);
nand U17358 (N_17358,N_8578,N_6880);
nand U17359 (N_17359,N_11448,N_10671);
nor U17360 (N_17360,N_11869,N_10909);
nand U17361 (N_17361,N_10992,N_10252);
xnor U17362 (N_17362,N_6938,N_11088);
xor U17363 (N_17363,N_8942,N_9236);
or U17364 (N_17364,N_8174,N_12471);
or U17365 (N_17365,N_10903,N_6961);
nand U17366 (N_17366,N_9637,N_11394);
or U17367 (N_17367,N_11434,N_6535);
nand U17368 (N_17368,N_8263,N_8016);
or U17369 (N_17369,N_11893,N_11024);
or U17370 (N_17370,N_12164,N_8416);
xor U17371 (N_17371,N_7653,N_9801);
and U17372 (N_17372,N_11150,N_8666);
xnor U17373 (N_17373,N_11494,N_6988);
nor U17374 (N_17374,N_7231,N_6340);
and U17375 (N_17375,N_7487,N_10982);
nand U17376 (N_17376,N_9340,N_6442);
nor U17377 (N_17377,N_11827,N_10289);
or U17378 (N_17378,N_12475,N_10907);
or U17379 (N_17379,N_12399,N_9168);
nand U17380 (N_17380,N_7513,N_9290);
or U17381 (N_17381,N_7449,N_9615);
or U17382 (N_17382,N_6510,N_7020);
nor U17383 (N_17383,N_11940,N_8069);
nor U17384 (N_17384,N_6522,N_8272);
nor U17385 (N_17385,N_6407,N_8662);
nor U17386 (N_17386,N_7368,N_8730);
nor U17387 (N_17387,N_8699,N_11755);
nand U17388 (N_17388,N_10816,N_8893);
or U17389 (N_17389,N_11420,N_9911);
nand U17390 (N_17390,N_6425,N_12184);
nor U17391 (N_17391,N_10685,N_12307);
nand U17392 (N_17392,N_10353,N_9914);
nor U17393 (N_17393,N_8742,N_8888);
nand U17394 (N_17394,N_11195,N_9254);
nor U17395 (N_17395,N_10482,N_10614);
nor U17396 (N_17396,N_7162,N_7091);
nand U17397 (N_17397,N_7489,N_11585);
and U17398 (N_17398,N_8243,N_7419);
or U17399 (N_17399,N_8940,N_11168);
nand U17400 (N_17400,N_8558,N_9472);
xor U17401 (N_17401,N_11583,N_11055);
nand U17402 (N_17402,N_8666,N_9861);
xnor U17403 (N_17403,N_11352,N_8948);
nor U17404 (N_17404,N_11558,N_6761);
nor U17405 (N_17405,N_10306,N_6992);
nor U17406 (N_17406,N_8771,N_8854);
or U17407 (N_17407,N_11947,N_11881);
nand U17408 (N_17408,N_11829,N_12237);
or U17409 (N_17409,N_7190,N_11646);
nand U17410 (N_17410,N_12326,N_10348);
xnor U17411 (N_17411,N_9975,N_6699);
and U17412 (N_17412,N_10072,N_9733);
and U17413 (N_17413,N_10916,N_11377);
nor U17414 (N_17414,N_10011,N_8357);
or U17415 (N_17415,N_11160,N_7477);
nand U17416 (N_17416,N_6706,N_7736);
nand U17417 (N_17417,N_9991,N_8089);
or U17418 (N_17418,N_7245,N_8541);
nor U17419 (N_17419,N_10863,N_11520);
and U17420 (N_17420,N_7727,N_8070);
nand U17421 (N_17421,N_7946,N_9452);
nor U17422 (N_17422,N_11036,N_10602);
or U17423 (N_17423,N_9531,N_7391);
and U17424 (N_17424,N_7648,N_8401);
or U17425 (N_17425,N_9584,N_7871);
nand U17426 (N_17426,N_11858,N_8263);
and U17427 (N_17427,N_11871,N_10339);
nor U17428 (N_17428,N_8213,N_11449);
nand U17429 (N_17429,N_11108,N_12287);
and U17430 (N_17430,N_12179,N_11951);
and U17431 (N_17431,N_9846,N_9672);
and U17432 (N_17432,N_11224,N_10131);
and U17433 (N_17433,N_12204,N_7428);
nand U17434 (N_17434,N_7508,N_10877);
and U17435 (N_17435,N_6620,N_10864);
nand U17436 (N_17436,N_9660,N_7299);
and U17437 (N_17437,N_10226,N_11567);
xnor U17438 (N_17438,N_11199,N_10055);
or U17439 (N_17439,N_11773,N_7748);
nor U17440 (N_17440,N_9518,N_6864);
nand U17441 (N_17441,N_10172,N_9151);
xor U17442 (N_17442,N_10987,N_7017);
and U17443 (N_17443,N_9136,N_8211);
and U17444 (N_17444,N_7762,N_7999);
nand U17445 (N_17445,N_6769,N_6570);
nand U17446 (N_17446,N_9506,N_6514);
nand U17447 (N_17447,N_6279,N_8151);
and U17448 (N_17448,N_7640,N_6722);
and U17449 (N_17449,N_8286,N_11519);
nand U17450 (N_17450,N_12260,N_11288);
nor U17451 (N_17451,N_6310,N_8582);
xor U17452 (N_17452,N_6719,N_8371);
or U17453 (N_17453,N_8192,N_12197);
and U17454 (N_17454,N_7161,N_7593);
xor U17455 (N_17455,N_6331,N_8463);
nor U17456 (N_17456,N_12229,N_10547);
nor U17457 (N_17457,N_12445,N_6692);
or U17458 (N_17458,N_11397,N_11536);
nor U17459 (N_17459,N_8375,N_12480);
or U17460 (N_17460,N_9215,N_7726);
and U17461 (N_17461,N_7000,N_10624);
nor U17462 (N_17462,N_12474,N_10931);
nand U17463 (N_17463,N_7691,N_9264);
or U17464 (N_17464,N_9559,N_10863);
nand U17465 (N_17465,N_10729,N_6412);
nand U17466 (N_17466,N_12155,N_7574);
nand U17467 (N_17467,N_7025,N_11498);
and U17468 (N_17468,N_11963,N_11421);
or U17469 (N_17469,N_7558,N_8708);
or U17470 (N_17470,N_8549,N_12307);
nor U17471 (N_17471,N_10481,N_10370);
or U17472 (N_17472,N_6441,N_7967);
or U17473 (N_17473,N_8764,N_11124);
nand U17474 (N_17474,N_12025,N_11713);
and U17475 (N_17475,N_8152,N_12144);
nand U17476 (N_17476,N_10894,N_7159);
nor U17477 (N_17477,N_10899,N_6542);
nand U17478 (N_17478,N_11758,N_6591);
and U17479 (N_17479,N_10782,N_10083);
nor U17480 (N_17480,N_7600,N_6786);
and U17481 (N_17481,N_6680,N_10941);
nor U17482 (N_17482,N_12383,N_10882);
nand U17483 (N_17483,N_9579,N_6892);
and U17484 (N_17484,N_8140,N_8580);
xnor U17485 (N_17485,N_9414,N_9318);
nand U17486 (N_17486,N_11444,N_9635);
nand U17487 (N_17487,N_9940,N_9256);
nor U17488 (N_17488,N_9027,N_11871);
xnor U17489 (N_17489,N_9376,N_11584);
or U17490 (N_17490,N_8521,N_12134);
or U17491 (N_17491,N_8923,N_8399);
and U17492 (N_17492,N_9006,N_6312);
and U17493 (N_17493,N_10364,N_7554);
or U17494 (N_17494,N_10600,N_11663);
or U17495 (N_17495,N_7325,N_10473);
xnor U17496 (N_17496,N_8816,N_7901);
nor U17497 (N_17497,N_7827,N_10449);
xor U17498 (N_17498,N_9906,N_8494);
xor U17499 (N_17499,N_11298,N_9794);
nor U17500 (N_17500,N_12114,N_7226);
nand U17501 (N_17501,N_8771,N_8931);
or U17502 (N_17502,N_11500,N_8118);
or U17503 (N_17503,N_10067,N_8843);
or U17504 (N_17504,N_8290,N_8505);
xnor U17505 (N_17505,N_8837,N_11617);
and U17506 (N_17506,N_8320,N_9037);
nor U17507 (N_17507,N_8892,N_10102);
nand U17508 (N_17508,N_6889,N_9258);
nor U17509 (N_17509,N_12277,N_11194);
xnor U17510 (N_17510,N_7959,N_8578);
and U17511 (N_17511,N_10158,N_6591);
nand U17512 (N_17512,N_6679,N_11054);
xnor U17513 (N_17513,N_10302,N_9417);
nor U17514 (N_17514,N_9244,N_7304);
and U17515 (N_17515,N_10433,N_11973);
or U17516 (N_17516,N_10319,N_11675);
nand U17517 (N_17517,N_7567,N_8133);
and U17518 (N_17518,N_9547,N_11664);
and U17519 (N_17519,N_11934,N_11611);
and U17520 (N_17520,N_12367,N_8075);
or U17521 (N_17521,N_7377,N_10782);
nor U17522 (N_17522,N_11674,N_12360);
nand U17523 (N_17523,N_11174,N_9379);
nor U17524 (N_17524,N_10683,N_11254);
or U17525 (N_17525,N_6856,N_10532);
nor U17526 (N_17526,N_6992,N_7109);
and U17527 (N_17527,N_7515,N_11936);
or U17528 (N_17528,N_10593,N_7720);
and U17529 (N_17529,N_10983,N_9569);
nand U17530 (N_17530,N_8476,N_11113);
or U17531 (N_17531,N_8971,N_8144);
or U17532 (N_17532,N_11833,N_12333);
or U17533 (N_17533,N_9252,N_11608);
and U17534 (N_17534,N_9660,N_12326);
nand U17535 (N_17535,N_6460,N_7547);
nand U17536 (N_17536,N_6633,N_7784);
nor U17537 (N_17537,N_10647,N_10952);
and U17538 (N_17538,N_8378,N_12235);
nand U17539 (N_17539,N_12292,N_11706);
nand U17540 (N_17540,N_11091,N_7804);
or U17541 (N_17541,N_8225,N_12454);
nor U17542 (N_17542,N_8390,N_12096);
or U17543 (N_17543,N_6565,N_9672);
and U17544 (N_17544,N_11791,N_12161);
and U17545 (N_17545,N_11232,N_11073);
nor U17546 (N_17546,N_6262,N_9446);
or U17547 (N_17547,N_7194,N_7777);
nor U17548 (N_17548,N_11831,N_8924);
and U17549 (N_17549,N_8674,N_11320);
and U17550 (N_17550,N_12210,N_7020);
nor U17551 (N_17551,N_6593,N_11815);
and U17552 (N_17552,N_9525,N_10400);
or U17553 (N_17553,N_11714,N_8548);
or U17554 (N_17554,N_6742,N_7538);
nand U17555 (N_17555,N_11569,N_11778);
xor U17556 (N_17556,N_10106,N_12309);
nand U17557 (N_17557,N_9258,N_10270);
xor U17558 (N_17558,N_6303,N_8067);
xnor U17559 (N_17559,N_7989,N_11390);
nor U17560 (N_17560,N_10022,N_7059);
nand U17561 (N_17561,N_9200,N_10091);
and U17562 (N_17562,N_7292,N_9151);
nor U17563 (N_17563,N_7708,N_10455);
and U17564 (N_17564,N_7935,N_12119);
nand U17565 (N_17565,N_9593,N_6694);
nor U17566 (N_17566,N_6311,N_8530);
nand U17567 (N_17567,N_6932,N_8859);
and U17568 (N_17568,N_12463,N_11923);
nor U17569 (N_17569,N_11008,N_9696);
nor U17570 (N_17570,N_8497,N_9500);
nand U17571 (N_17571,N_8774,N_9102);
xnor U17572 (N_17572,N_10436,N_11332);
or U17573 (N_17573,N_9478,N_6727);
and U17574 (N_17574,N_8541,N_9737);
nor U17575 (N_17575,N_11167,N_11402);
nand U17576 (N_17576,N_8449,N_9187);
nor U17577 (N_17577,N_7209,N_7136);
nor U17578 (N_17578,N_8188,N_12487);
nor U17579 (N_17579,N_12486,N_9247);
nand U17580 (N_17580,N_7694,N_9384);
nor U17581 (N_17581,N_6890,N_11097);
and U17582 (N_17582,N_6679,N_10287);
xor U17583 (N_17583,N_10331,N_8556);
and U17584 (N_17584,N_12152,N_11951);
nand U17585 (N_17585,N_10682,N_11872);
and U17586 (N_17586,N_8353,N_10899);
and U17587 (N_17587,N_8367,N_7606);
or U17588 (N_17588,N_12028,N_11872);
nand U17589 (N_17589,N_8060,N_10642);
nand U17590 (N_17590,N_11813,N_9375);
and U17591 (N_17591,N_11366,N_11010);
nand U17592 (N_17592,N_9919,N_9726);
xor U17593 (N_17593,N_6467,N_9462);
xor U17594 (N_17594,N_6782,N_11481);
nor U17595 (N_17595,N_8817,N_12256);
or U17596 (N_17596,N_10831,N_10731);
nand U17597 (N_17597,N_11928,N_11542);
or U17598 (N_17598,N_10806,N_6716);
nand U17599 (N_17599,N_10836,N_12189);
or U17600 (N_17600,N_8263,N_11255);
nor U17601 (N_17601,N_10653,N_9234);
nand U17602 (N_17602,N_9419,N_8458);
nor U17603 (N_17603,N_8637,N_7939);
nand U17604 (N_17604,N_9258,N_11388);
xor U17605 (N_17605,N_8224,N_6961);
nand U17606 (N_17606,N_9539,N_11224);
nand U17607 (N_17607,N_11963,N_8158);
nand U17608 (N_17608,N_8096,N_9122);
nand U17609 (N_17609,N_9791,N_10254);
nand U17610 (N_17610,N_6258,N_8056);
or U17611 (N_17611,N_8630,N_11307);
nor U17612 (N_17612,N_12262,N_10442);
or U17613 (N_17613,N_11780,N_7707);
or U17614 (N_17614,N_11200,N_7178);
and U17615 (N_17615,N_11095,N_11126);
or U17616 (N_17616,N_7009,N_10026);
nand U17617 (N_17617,N_12040,N_9019);
and U17618 (N_17618,N_8107,N_10455);
or U17619 (N_17619,N_11320,N_8687);
and U17620 (N_17620,N_6463,N_6404);
nand U17621 (N_17621,N_12481,N_8725);
and U17622 (N_17622,N_7474,N_8004);
and U17623 (N_17623,N_9273,N_11821);
and U17624 (N_17624,N_6872,N_11879);
or U17625 (N_17625,N_9910,N_6897);
nand U17626 (N_17626,N_9604,N_11855);
nand U17627 (N_17627,N_6615,N_10976);
nand U17628 (N_17628,N_11651,N_6498);
nand U17629 (N_17629,N_9265,N_9516);
and U17630 (N_17630,N_8106,N_10907);
nand U17631 (N_17631,N_7302,N_9041);
and U17632 (N_17632,N_11809,N_12352);
and U17633 (N_17633,N_6676,N_6504);
nor U17634 (N_17634,N_7078,N_12176);
or U17635 (N_17635,N_12087,N_6997);
or U17636 (N_17636,N_12468,N_11493);
and U17637 (N_17637,N_7300,N_8184);
xnor U17638 (N_17638,N_8193,N_12042);
or U17639 (N_17639,N_11697,N_6996);
or U17640 (N_17640,N_9150,N_11537);
xor U17641 (N_17641,N_11036,N_7733);
nand U17642 (N_17642,N_12251,N_8566);
nand U17643 (N_17643,N_11002,N_7541);
and U17644 (N_17644,N_11022,N_11874);
nor U17645 (N_17645,N_10016,N_8975);
or U17646 (N_17646,N_6436,N_11890);
nor U17647 (N_17647,N_10322,N_10348);
or U17648 (N_17648,N_10488,N_8607);
xnor U17649 (N_17649,N_7869,N_8583);
and U17650 (N_17650,N_11609,N_10011);
nor U17651 (N_17651,N_7221,N_7444);
nor U17652 (N_17652,N_6687,N_6599);
and U17653 (N_17653,N_11849,N_8414);
nor U17654 (N_17654,N_11873,N_11726);
and U17655 (N_17655,N_10341,N_12276);
nor U17656 (N_17656,N_9967,N_7654);
nor U17657 (N_17657,N_9116,N_6560);
nand U17658 (N_17658,N_6331,N_7863);
nand U17659 (N_17659,N_7112,N_11569);
or U17660 (N_17660,N_7748,N_12381);
nor U17661 (N_17661,N_6612,N_9931);
nor U17662 (N_17662,N_12442,N_6896);
nor U17663 (N_17663,N_10175,N_9346);
and U17664 (N_17664,N_9216,N_8076);
and U17665 (N_17665,N_10047,N_12058);
and U17666 (N_17666,N_11635,N_8128);
and U17667 (N_17667,N_10403,N_12434);
or U17668 (N_17668,N_11868,N_8783);
nor U17669 (N_17669,N_6677,N_10028);
and U17670 (N_17670,N_12205,N_9766);
or U17671 (N_17671,N_9933,N_8104);
or U17672 (N_17672,N_9669,N_8986);
nand U17673 (N_17673,N_6671,N_8856);
nand U17674 (N_17674,N_9972,N_7749);
nor U17675 (N_17675,N_9598,N_7040);
nor U17676 (N_17676,N_6357,N_8529);
nand U17677 (N_17677,N_8103,N_7517);
or U17678 (N_17678,N_7029,N_7970);
or U17679 (N_17679,N_9380,N_7569);
or U17680 (N_17680,N_7449,N_8850);
and U17681 (N_17681,N_8182,N_7699);
nand U17682 (N_17682,N_12039,N_8045);
nor U17683 (N_17683,N_6531,N_6486);
and U17684 (N_17684,N_10329,N_12259);
or U17685 (N_17685,N_11557,N_10635);
or U17686 (N_17686,N_6309,N_6315);
or U17687 (N_17687,N_7262,N_6496);
nand U17688 (N_17688,N_7260,N_6817);
or U17689 (N_17689,N_8208,N_8014);
and U17690 (N_17690,N_8244,N_7777);
and U17691 (N_17691,N_9911,N_7275);
or U17692 (N_17692,N_8770,N_9192);
and U17693 (N_17693,N_9735,N_11316);
or U17694 (N_17694,N_8329,N_9533);
nor U17695 (N_17695,N_6827,N_11960);
nand U17696 (N_17696,N_11475,N_10896);
and U17697 (N_17697,N_11369,N_12442);
or U17698 (N_17698,N_6262,N_12201);
or U17699 (N_17699,N_9719,N_12443);
nor U17700 (N_17700,N_10729,N_11433);
nor U17701 (N_17701,N_11289,N_9078);
and U17702 (N_17702,N_8394,N_10047);
and U17703 (N_17703,N_8635,N_6486);
nor U17704 (N_17704,N_8083,N_8650);
nand U17705 (N_17705,N_11510,N_8424);
nand U17706 (N_17706,N_10206,N_8323);
nor U17707 (N_17707,N_6944,N_7192);
and U17708 (N_17708,N_7312,N_8249);
xnor U17709 (N_17709,N_10675,N_8782);
nor U17710 (N_17710,N_7303,N_9780);
nand U17711 (N_17711,N_9834,N_8023);
nand U17712 (N_17712,N_6986,N_8305);
nand U17713 (N_17713,N_8725,N_10651);
and U17714 (N_17714,N_12151,N_7809);
nor U17715 (N_17715,N_11131,N_8112);
nand U17716 (N_17716,N_6859,N_10749);
nor U17717 (N_17717,N_7342,N_8835);
nor U17718 (N_17718,N_10106,N_9753);
and U17719 (N_17719,N_8258,N_7389);
nor U17720 (N_17720,N_8216,N_7409);
xor U17721 (N_17721,N_8665,N_11190);
or U17722 (N_17722,N_9087,N_9346);
nand U17723 (N_17723,N_10748,N_7436);
or U17724 (N_17724,N_10699,N_6464);
nor U17725 (N_17725,N_6346,N_7621);
and U17726 (N_17726,N_11925,N_7489);
or U17727 (N_17727,N_9187,N_10437);
nor U17728 (N_17728,N_10280,N_7266);
nor U17729 (N_17729,N_8892,N_10576);
or U17730 (N_17730,N_8140,N_11286);
or U17731 (N_17731,N_12189,N_9538);
and U17732 (N_17732,N_11383,N_6445);
nor U17733 (N_17733,N_11326,N_10482);
nand U17734 (N_17734,N_6723,N_7413);
and U17735 (N_17735,N_10480,N_9991);
nand U17736 (N_17736,N_8723,N_9670);
and U17737 (N_17737,N_10523,N_7605);
or U17738 (N_17738,N_8191,N_10740);
nor U17739 (N_17739,N_11065,N_10834);
nand U17740 (N_17740,N_9023,N_8934);
nand U17741 (N_17741,N_9618,N_6266);
and U17742 (N_17742,N_8035,N_9783);
nor U17743 (N_17743,N_9565,N_6925);
nor U17744 (N_17744,N_11424,N_7651);
nor U17745 (N_17745,N_7305,N_10832);
and U17746 (N_17746,N_11961,N_8023);
nor U17747 (N_17747,N_6978,N_6905);
xnor U17748 (N_17748,N_8197,N_11343);
and U17749 (N_17749,N_9392,N_8837);
nor U17750 (N_17750,N_9933,N_10565);
or U17751 (N_17751,N_12326,N_11263);
nand U17752 (N_17752,N_10962,N_7612);
nor U17753 (N_17753,N_8191,N_7334);
nand U17754 (N_17754,N_11911,N_6328);
nand U17755 (N_17755,N_10150,N_8704);
nor U17756 (N_17756,N_9035,N_7262);
or U17757 (N_17757,N_6526,N_7595);
nor U17758 (N_17758,N_9373,N_9141);
and U17759 (N_17759,N_11687,N_9326);
nand U17760 (N_17760,N_12236,N_7359);
nand U17761 (N_17761,N_12081,N_11307);
nand U17762 (N_17762,N_7808,N_6413);
nor U17763 (N_17763,N_9125,N_8948);
nor U17764 (N_17764,N_8384,N_9222);
or U17765 (N_17765,N_12032,N_12474);
nor U17766 (N_17766,N_11737,N_8490);
and U17767 (N_17767,N_9579,N_8870);
nor U17768 (N_17768,N_8511,N_8532);
nor U17769 (N_17769,N_9720,N_7730);
and U17770 (N_17770,N_6549,N_6971);
nor U17771 (N_17771,N_7807,N_9531);
and U17772 (N_17772,N_11700,N_9696);
and U17773 (N_17773,N_8343,N_9224);
nand U17774 (N_17774,N_8686,N_10505);
nor U17775 (N_17775,N_9115,N_9508);
nor U17776 (N_17776,N_10919,N_9388);
nand U17777 (N_17777,N_12127,N_6314);
or U17778 (N_17778,N_12061,N_8221);
nand U17779 (N_17779,N_10293,N_9980);
or U17780 (N_17780,N_9441,N_12445);
nand U17781 (N_17781,N_10704,N_12172);
nand U17782 (N_17782,N_10819,N_8160);
nor U17783 (N_17783,N_8370,N_6277);
nor U17784 (N_17784,N_7027,N_10454);
nand U17785 (N_17785,N_9470,N_6957);
or U17786 (N_17786,N_6534,N_8271);
nor U17787 (N_17787,N_10559,N_8302);
or U17788 (N_17788,N_10180,N_8959);
or U17789 (N_17789,N_11635,N_7773);
nor U17790 (N_17790,N_7715,N_10143);
nor U17791 (N_17791,N_10703,N_11007);
xnor U17792 (N_17792,N_8057,N_10731);
xnor U17793 (N_17793,N_7289,N_7637);
or U17794 (N_17794,N_9319,N_10908);
nand U17795 (N_17795,N_8899,N_8398);
nor U17796 (N_17796,N_10483,N_10622);
nand U17797 (N_17797,N_7557,N_7515);
and U17798 (N_17798,N_8228,N_11434);
and U17799 (N_17799,N_6883,N_10538);
nor U17800 (N_17800,N_8734,N_8267);
and U17801 (N_17801,N_7901,N_8283);
nand U17802 (N_17802,N_6580,N_7876);
or U17803 (N_17803,N_10056,N_12346);
or U17804 (N_17804,N_8251,N_12307);
nor U17805 (N_17805,N_9290,N_10011);
xnor U17806 (N_17806,N_8804,N_9485);
or U17807 (N_17807,N_9698,N_7104);
or U17808 (N_17808,N_8811,N_8765);
and U17809 (N_17809,N_9433,N_8383);
and U17810 (N_17810,N_9470,N_8505);
and U17811 (N_17811,N_9666,N_8100);
nand U17812 (N_17812,N_11999,N_11850);
nand U17813 (N_17813,N_7849,N_8729);
nor U17814 (N_17814,N_7728,N_6673);
and U17815 (N_17815,N_9319,N_7558);
nor U17816 (N_17816,N_7856,N_8474);
xnor U17817 (N_17817,N_11003,N_12235);
nor U17818 (N_17818,N_9594,N_10396);
nor U17819 (N_17819,N_12105,N_7423);
nand U17820 (N_17820,N_9453,N_8835);
xor U17821 (N_17821,N_10710,N_10510);
or U17822 (N_17822,N_8910,N_8303);
and U17823 (N_17823,N_7239,N_8570);
nor U17824 (N_17824,N_7242,N_8268);
and U17825 (N_17825,N_10870,N_6975);
or U17826 (N_17826,N_10358,N_11230);
nand U17827 (N_17827,N_8391,N_9162);
or U17828 (N_17828,N_11379,N_7782);
nand U17829 (N_17829,N_7709,N_8592);
and U17830 (N_17830,N_7945,N_11145);
or U17831 (N_17831,N_8554,N_9300);
or U17832 (N_17832,N_8567,N_7645);
or U17833 (N_17833,N_12174,N_8636);
and U17834 (N_17834,N_10979,N_10764);
nand U17835 (N_17835,N_6902,N_8052);
and U17836 (N_17836,N_9876,N_7661);
nor U17837 (N_17837,N_12459,N_7398);
nor U17838 (N_17838,N_7879,N_7719);
and U17839 (N_17839,N_6274,N_10492);
or U17840 (N_17840,N_8703,N_9430);
nand U17841 (N_17841,N_6361,N_10292);
and U17842 (N_17842,N_10440,N_9891);
nor U17843 (N_17843,N_12279,N_10663);
nand U17844 (N_17844,N_10860,N_9896);
or U17845 (N_17845,N_6694,N_6433);
and U17846 (N_17846,N_7689,N_7482);
nor U17847 (N_17847,N_7503,N_9879);
or U17848 (N_17848,N_10187,N_6456);
and U17849 (N_17849,N_11572,N_7707);
nand U17850 (N_17850,N_11526,N_10112);
and U17851 (N_17851,N_11014,N_8832);
nor U17852 (N_17852,N_7715,N_12395);
nand U17853 (N_17853,N_12328,N_11997);
nand U17854 (N_17854,N_11960,N_9439);
and U17855 (N_17855,N_8950,N_12453);
or U17856 (N_17856,N_7186,N_8812);
nor U17857 (N_17857,N_6470,N_8245);
nor U17858 (N_17858,N_7406,N_7313);
xor U17859 (N_17859,N_9729,N_10956);
xnor U17860 (N_17860,N_8135,N_11560);
or U17861 (N_17861,N_6323,N_9254);
nand U17862 (N_17862,N_8524,N_10698);
and U17863 (N_17863,N_9423,N_10608);
or U17864 (N_17864,N_11524,N_8630);
or U17865 (N_17865,N_12254,N_7632);
and U17866 (N_17866,N_10883,N_9277);
xnor U17867 (N_17867,N_8077,N_10375);
nand U17868 (N_17868,N_8143,N_7901);
xor U17869 (N_17869,N_6435,N_8108);
or U17870 (N_17870,N_10867,N_10648);
nor U17871 (N_17871,N_9862,N_7104);
nand U17872 (N_17872,N_6596,N_10338);
or U17873 (N_17873,N_9405,N_7251);
xnor U17874 (N_17874,N_9690,N_10540);
and U17875 (N_17875,N_9437,N_12144);
or U17876 (N_17876,N_7578,N_10623);
nand U17877 (N_17877,N_9446,N_11467);
or U17878 (N_17878,N_8002,N_9615);
and U17879 (N_17879,N_7239,N_8232);
nor U17880 (N_17880,N_6266,N_11138);
xnor U17881 (N_17881,N_8452,N_8443);
nand U17882 (N_17882,N_6539,N_8929);
or U17883 (N_17883,N_9984,N_10647);
nand U17884 (N_17884,N_11297,N_10074);
nand U17885 (N_17885,N_6957,N_6993);
nand U17886 (N_17886,N_10186,N_8044);
nand U17887 (N_17887,N_11728,N_7399);
nor U17888 (N_17888,N_9486,N_8934);
or U17889 (N_17889,N_7612,N_9566);
and U17890 (N_17890,N_10405,N_10689);
or U17891 (N_17891,N_10240,N_11865);
nor U17892 (N_17892,N_9262,N_11394);
and U17893 (N_17893,N_9208,N_12466);
nor U17894 (N_17894,N_7256,N_9080);
or U17895 (N_17895,N_7148,N_9388);
nand U17896 (N_17896,N_7532,N_12153);
and U17897 (N_17897,N_10843,N_11152);
nor U17898 (N_17898,N_9425,N_8444);
and U17899 (N_17899,N_8360,N_7541);
and U17900 (N_17900,N_9208,N_12490);
and U17901 (N_17901,N_6784,N_12267);
xnor U17902 (N_17902,N_10660,N_12340);
nor U17903 (N_17903,N_9450,N_10588);
nor U17904 (N_17904,N_11436,N_6859);
and U17905 (N_17905,N_8773,N_6934);
or U17906 (N_17906,N_8176,N_12448);
nand U17907 (N_17907,N_9297,N_6294);
or U17908 (N_17908,N_6284,N_11719);
and U17909 (N_17909,N_10705,N_9121);
nor U17910 (N_17910,N_10668,N_8611);
xor U17911 (N_17911,N_9249,N_9048);
or U17912 (N_17912,N_6605,N_8235);
or U17913 (N_17913,N_12386,N_10601);
nand U17914 (N_17914,N_11520,N_12006);
nor U17915 (N_17915,N_7929,N_7652);
or U17916 (N_17916,N_11454,N_10000);
nand U17917 (N_17917,N_9291,N_10486);
or U17918 (N_17918,N_10442,N_8997);
nor U17919 (N_17919,N_7092,N_11440);
and U17920 (N_17920,N_9804,N_9472);
nor U17921 (N_17921,N_8780,N_6855);
and U17922 (N_17922,N_10829,N_7824);
nand U17923 (N_17923,N_9921,N_8739);
nor U17924 (N_17924,N_10218,N_12204);
nor U17925 (N_17925,N_11054,N_8345);
and U17926 (N_17926,N_6804,N_7954);
or U17927 (N_17927,N_6480,N_8189);
and U17928 (N_17928,N_6927,N_9065);
nand U17929 (N_17929,N_11278,N_10642);
nand U17930 (N_17930,N_7899,N_10025);
xnor U17931 (N_17931,N_9825,N_10330);
nor U17932 (N_17932,N_9461,N_9601);
nand U17933 (N_17933,N_11640,N_8514);
or U17934 (N_17934,N_8529,N_6453);
and U17935 (N_17935,N_11232,N_6878);
nand U17936 (N_17936,N_8202,N_11427);
and U17937 (N_17937,N_8579,N_9486);
xor U17938 (N_17938,N_8167,N_6843);
xor U17939 (N_17939,N_11814,N_8601);
or U17940 (N_17940,N_12167,N_12124);
nand U17941 (N_17941,N_10654,N_7318);
nand U17942 (N_17942,N_11435,N_8910);
nand U17943 (N_17943,N_10725,N_9645);
and U17944 (N_17944,N_8456,N_6889);
nor U17945 (N_17945,N_9183,N_7643);
nand U17946 (N_17946,N_9349,N_11256);
and U17947 (N_17947,N_7375,N_9260);
nand U17948 (N_17948,N_7333,N_12154);
nor U17949 (N_17949,N_10269,N_10575);
nand U17950 (N_17950,N_8398,N_9765);
and U17951 (N_17951,N_7331,N_11716);
and U17952 (N_17952,N_7168,N_11010);
xnor U17953 (N_17953,N_10171,N_10217);
nor U17954 (N_17954,N_6615,N_6540);
nor U17955 (N_17955,N_12318,N_12473);
nor U17956 (N_17956,N_9910,N_6857);
or U17957 (N_17957,N_10821,N_11881);
nand U17958 (N_17958,N_7726,N_7775);
nand U17959 (N_17959,N_7264,N_7282);
and U17960 (N_17960,N_9048,N_11292);
nor U17961 (N_17961,N_7474,N_9218);
nand U17962 (N_17962,N_7268,N_9991);
nor U17963 (N_17963,N_11130,N_6925);
and U17964 (N_17964,N_9466,N_10329);
nor U17965 (N_17965,N_7752,N_11602);
nor U17966 (N_17966,N_11151,N_11270);
nor U17967 (N_17967,N_11808,N_9580);
and U17968 (N_17968,N_9395,N_7151);
nor U17969 (N_17969,N_8492,N_6927);
xor U17970 (N_17970,N_8371,N_11992);
nand U17971 (N_17971,N_7430,N_8174);
nand U17972 (N_17972,N_8222,N_8167);
or U17973 (N_17973,N_10054,N_6867);
and U17974 (N_17974,N_7398,N_12314);
and U17975 (N_17975,N_9747,N_9513);
and U17976 (N_17976,N_9970,N_6986);
or U17977 (N_17977,N_12045,N_7797);
nor U17978 (N_17978,N_12212,N_8011);
and U17979 (N_17979,N_11375,N_9734);
nand U17980 (N_17980,N_9972,N_8697);
nand U17981 (N_17981,N_7417,N_8700);
nand U17982 (N_17982,N_11162,N_9834);
or U17983 (N_17983,N_11880,N_10744);
nand U17984 (N_17984,N_10347,N_10168);
nand U17985 (N_17985,N_10348,N_7099);
and U17986 (N_17986,N_6644,N_6352);
or U17987 (N_17987,N_7322,N_10942);
xor U17988 (N_17988,N_10191,N_7277);
and U17989 (N_17989,N_7650,N_10714);
and U17990 (N_17990,N_6788,N_12345);
nor U17991 (N_17991,N_11088,N_7539);
or U17992 (N_17992,N_11994,N_10111);
or U17993 (N_17993,N_11227,N_11225);
nand U17994 (N_17994,N_9222,N_9264);
nand U17995 (N_17995,N_11580,N_12018);
xnor U17996 (N_17996,N_7618,N_9073);
or U17997 (N_17997,N_7814,N_7966);
and U17998 (N_17998,N_8954,N_7185);
nand U17999 (N_17999,N_9845,N_6250);
nor U18000 (N_18000,N_6466,N_9833);
and U18001 (N_18001,N_9481,N_11001);
nand U18002 (N_18002,N_8433,N_7655);
and U18003 (N_18003,N_9803,N_8296);
or U18004 (N_18004,N_8550,N_6323);
or U18005 (N_18005,N_7059,N_7269);
and U18006 (N_18006,N_8702,N_9259);
nor U18007 (N_18007,N_6686,N_9761);
xor U18008 (N_18008,N_6889,N_8582);
and U18009 (N_18009,N_12475,N_6739);
and U18010 (N_18010,N_8838,N_7230);
or U18011 (N_18011,N_8360,N_9719);
nor U18012 (N_18012,N_7250,N_10191);
or U18013 (N_18013,N_7070,N_8654);
or U18014 (N_18014,N_11371,N_8260);
nor U18015 (N_18015,N_11621,N_12072);
nor U18016 (N_18016,N_8847,N_10383);
and U18017 (N_18017,N_11883,N_9472);
or U18018 (N_18018,N_8332,N_11471);
nand U18019 (N_18019,N_10505,N_11405);
nand U18020 (N_18020,N_9825,N_7996);
nor U18021 (N_18021,N_9543,N_10213);
xor U18022 (N_18022,N_12322,N_7358);
nand U18023 (N_18023,N_11159,N_12073);
and U18024 (N_18024,N_11764,N_6749);
nand U18025 (N_18025,N_8333,N_11448);
or U18026 (N_18026,N_10467,N_8246);
and U18027 (N_18027,N_11787,N_7705);
nand U18028 (N_18028,N_8325,N_11465);
nand U18029 (N_18029,N_8254,N_10297);
xor U18030 (N_18030,N_9037,N_7652);
nor U18031 (N_18031,N_8522,N_7086);
nor U18032 (N_18032,N_11536,N_8478);
nor U18033 (N_18033,N_8596,N_6895);
xnor U18034 (N_18034,N_6411,N_10350);
or U18035 (N_18035,N_10454,N_12264);
nand U18036 (N_18036,N_12360,N_11886);
and U18037 (N_18037,N_12355,N_8493);
nand U18038 (N_18038,N_7407,N_7946);
nor U18039 (N_18039,N_10578,N_6988);
and U18040 (N_18040,N_9902,N_12045);
and U18041 (N_18041,N_12453,N_6559);
or U18042 (N_18042,N_10071,N_11172);
nor U18043 (N_18043,N_9765,N_6728);
nor U18044 (N_18044,N_8293,N_8890);
nand U18045 (N_18045,N_7652,N_10875);
nand U18046 (N_18046,N_11651,N_8395);
and U18047 (N_18047,N_10475,N_6339);
and U18048 (N_18048,N_11937,N_6828);
and U18049 (N_18049,N_7112,N_12462);
or U18050 (N_18050,N_10630,N_6758);
or U18051 (N_18051,N_11033,N_11784);
nor U18052 (N_18052,N_10811,N_8534);
or U18053 (N_18053,N_7654,N_11283);
or U18054 (N_18054,N_8403,N_7018);
or U18055 (N_18055,N_11373,N_8313);
nand U18056 (N_18056,N_8229,N_9400);
nand U18057 (N_18057,N_9478,N_10224);
nor U18058 (N_18058,N_6721,N_11863);
nor U18059 (N_18059,N_7765,N_9916);
nand U18060 (N_18060,N_6491,N_10196);
nor U18061 (N_18061,N_9622,N_12454);
or U18062 (N_18062,N_12105,N_11425);
and U18063 (N_18063,N_8231,N_9383);
nor U18064 (N_18064,N_8460,N_10738);
and U18065 (N_18065,N_11066,N_8358);
or U18066 (N_18066,N_11094,N_8949);
and U18067 (N_18067,N_10167,N_6680);
nor U18068 (N_18068,N_7438,N_7314);
nand U18069 (N_18069,N_6621,N_7441);
nand U18070 (N_18070,N_6822,N_7278);
nor U18071 (N_18071,N_11800,N_8745);
and U18072 (N_18072,N_6478,N_9978);
or U18073 (N_18073,N_8000,N_10296);
nand U18074 (N_18074,N_6602,N_10945);
nand U18075 (N_18075,N_10243,N_7795);
nand U18076 (N_18076,N_8708,N_8375);
and U18077 (N_18077,N_6830,N_10201);
nor U18078 (N_18078,N_8775,N_11643);
or U18079 (N_18079,N_9813,N_6642);
nand U18080 (N_18080,N_7453,N_12176);
xor U18081 (N_18081,N_11927,N_9932);
or U18082 (N_18082,N_8177,N_11351);
nor U18083 (N_18083,N_12286,N_7526);
nor U18084 (N_18084,N_7625,N_10226);
and U18085 (N_18085,N_12037,N_8459);
and U18086 (N_18086,N_9316,N_12318);
nand U18087 (N_18087,N_12171,N_10042);
or U18088 (N_18088,N_6431,N_9550);
nand U18089 (N_18089,N_7492,N_10571);
or U18090 (N_18090,N_6431,N_8276);
or U18091 (N_18091,N_8267,N_11803);
or U18092 (N_18092,N_7265,N_7650);
and U18093 (N_18093,N_11497,N_11748);
xnor U18094 (N_18094,N_12231,N_8830);
nor U18095 (N_18095,N_7152,N_8744);
nand U18096 (N_18096,N_8695,N_6655);
and U18097 (N_18097,N_10454,N_6464);
nand U18098 (N_18098,N_7734,N_6485);
nand U18099 (N_18099,N_9558,N_7823);
and U18100 (N_18100,N_7689,N_7719);
and U18101 (N_18101,N_6650,N_9925);
xor U18102 (N_18102,N_10536,N_9452);
nor U18103 (N_18103,N_8131,N_10467);
or U18104 (N_18104,N_10590,N_6839);
nor U18105 (N_18105,N_9349,N_8168);
or U18106 (N_18106,N_8400,N_12154);
and U18107 (N_18107,N_11554,N_11896);
nor U18108 (N_18108,N_8367,N_6919);
xor U18109 (N_18109,N_7968,N_10050);
or U18110 (N_18110,N_11689,N_6958);
nor U18111 (N_18111,N_8278,N_10200);
nand U18112 (N_18112,N_9130,N_12081);
nand U18113 (N_18113,N_10248,N_9027);
nor U18114 (N_18114,N_9778,N_6439);
nor U18115 (N_18115,N_6389,N_12085);
xnor U18116 (N_18116,N_6807,N_9650);
and U18117 (N_18117,N_8082,N_7325);
or U18118 (N_18118,N_6974,N_8642);
nand U18119 (N_18119,N_7402,N_10057);
nand U18120 (N_18120,N_10918,N_9233);
nor U18121 (N_18121,N_11518,N_9961);
nor U18122 (N_18122,N_10204,N_12145);
nand U18123 (N_18123,N_7296,N_9319);
and U18124 (N_18124,N_6406,N_7443);
or U18125 (N_18125,N_6313,N_7642);
nand U18126 (N_18126,N_8693,N_9331);
nand U18127 (N_18127,N_10818,N_9200);
and U18128 (N_18128,N_9666,N_12039);
nor U18129 (N_18129,N_9167,N_8109);
or U18130 (N_18130,N_8440,N_11719);
nor U18131 (N_18131,N_9306,N_8592);
nand U18132 (N_18132,N_11263,N_8521);
nand U18133 (N_18133,N_12127,N_11352);
or U18134 (N_18134,N_8064,N_8763);
and U18135 (N_18135,N_10961,N_8336);
nand U18136 (N_18136,N_11243,N_8956);
nor U18137 (N_18137,N_10914,N_8717);
and U18138 (N_18138,N_9166,N_7610);
nand U18139 (N_18139,N_9801,N_11374);
nand U18140 (N_18140,N_10635,N_10953);
xor U18141 (N_18141,N_7480,N_11195);
nor U18142 (N_18142,N_7340,N_8007);
nor U18143 (N_18143,N_6977,N_9142);
nand U18144 (N_18144,N_11750,N_9114);
or U18145 (N_18145,N_10849,N_10361);
nor U18146 (N_18146,N_10008,N_8808);
and U18147 (N_18147,N_8292,N_6386);
nor U18148 (N_18148,N_8630,N_8742);
and U18149 (N_18149,N_6815,N_10582);
nand U18150 (N_18150,N_7370,N_7895);
nand U18151 (N_18151,N_12222,N_8932);
xor U18152 (N_18152,N_11176,N_11380);
or U18153 (N_18153,N_11923,N_9273);
and U18154 (N_18154,N_11328,N_7771);
and U18155 (N_18155,N_12368,N_8264);
and U18156 (N_18156,N_10717,N_10227);
nand U18157 (N_18157,N_6937,N_8419);
or U18158 (N_18158,N_11429,N_10703);
or U18159 (N_18159,N_11338,N_10644);
xnor U18160 (N_18160,N_8232,N_8400);
and U18161 (N_18161,N_9459,N_10912);
xnor U18162 (N_18162,N_10630,N_12440);
nor U18163 (N_18163,N_12409,N_8967);
and U18164 (N_18164,N_9837,N_7275);
nand U18165 (N_18165,N_12388,N_11006);
nand U18166 (N_18166,N_12358,N_9434);
and U18167 (N_18167,N_9541,N_6445);
nor U18168 (N_18168,N_9047,N_6635);
or U18169 (N_18169,N_6741,N_8450);
nand U18170 (N_18170,N_8134,N_9186);
nand U18171 (N_18171,N_10848,N_11409);
or U18172 (N_18172,N_7937,N_6250);
nor U18173 (N_18173,N_9598,N_12079);
xnor U18174 (N_18174,N_10998,N_6482);
nor U18175 (N_18175,N_12405,N_8680);
or U18176 (N_18176,N_6960,N_6253);
and U18177 (N_18177,N_6796,N_10598);
and U18178 (N_18178,N_7495,N_7611);
and U18179 (N_18179,N_8092,N_7706);
nor U18180 (N_18180,N_9098,N_8438);
or U18181 (N_18181,N_11618,N_9544);
or U18182 (N_18182,N_9364,N_7305);
nor U18183 (N_18183,N_11542,N_11211);
and U18184 (N_18184,N_7728,N_6792);
or U18185 (N_18185,N_9209,N_8617);
nand U18186 (N_18186,N_7416,N_10000);
nor U18187 (N_18187,N_8600,N_7345);
xnor U18188 (N_18188,N_7987,N_7340);
and U18189 (N_18189,N_10078,N_9774);
nor U18190 (N_18190,N_10246,N_9659);
nor U18191 (N_18191,N_9650,N_10834);
and U18192 (N_18192,N_10952,N_11073);
nand U18193 (N_18193,N_9941,N_10350);
xnor U18194 (N_18194,N_7276,N_9125);
nor U18195 (N_18195,N_8749,N_12344);
nand U18196 (N_18196,N_9066,N_9584);
or U18197 (N_18197,N_7631,N_11271);
nand U18198 (N_18198,N_8463,N_12414);
nand U18199 (N_18199,N_9264,N_8528);
and U18200 (N_18200,N_11627,N_8977);
or U18201 (N_18201,N_9576,N_9039);
nor U18202 (N_18202,N_10698,N_9043);
nand U18203 (N_18203,N_10735,N_8790);
nor U18204 (N_18204,N_12186,N_12165);
and U18205 (N_18205,N_9085,N_10344);
xnor U18206 (N_18206,N_7391,N_10444);
nand U18207 (N_18207,N_10062,N_9905);
nand U18208 (N_18208,N_11197,N_6421);
nand U18209 (N_18209,N_7287,N_7322);
nor U18210 (N_18210,N_9947,N_8114);
and U18211 (N_18211,N_10039,N_10152);
xnor U18212 (N_18212,N_9949,N_9301);
xnor U18213 (N_18213,N_8797,N_12289);
nor U18214 (N_18214,N_10613,N_7575);
or U18215 (N_18215,N_8899,N_7659);
and U18216 (N_18216,N_10366,N_7733);
xor U18217 (N_18217,N_12056,N_11057);
or U18218 (N_18218,N_11771,N_7270);
nor U18219 (N_18219,N_9045,N_11359);
xnor U18220 (N_18220,N_9344,N_11462);
nor U18221 (N_18221,N_8414,N_11365);
or U18222 (N_18222,N_9323,N_12417);
and U18223 (N_18223,N_10043,N_6289);
nor U18224 (N_18224,N_11422,N_11186);
nand U18225 (N_18225,N_11358,N_12027);
and U18226 (N_18226,N_7112,N_8154);
and U18227 (N_18227,N_7142,N_12432);
and U18228 (N_18228,N_9054,N_8839);
nand U18229 (N_18229,N_9555,N_8990);
nor U18230 (N_18230,N_6600,N_7435);
or U18231 (N_18231,N_12148,N_7522);
and U18232 (N_18232,N_9928,N_10432);
xnor U18233 (N_18233,N_9593,N_8471);
and U18234 (N_18234,N_11724,N_12226);
nand U18235 (N_18235,N_12238,N_11811);
or U18236 (N_18236,N_6298,N_11144);
nand U18237 (N_18237,N_11718,N_9343);
xor U18238 (N_18238,N_6552,N_10637);
xnor U18239 (N_18239,N_8900,N_6586);
or U18240 (N_18240,N_11907,N_12158);
and U18241 (N_18241,N_9127,N_10719);
and U18242 (N_18242,N_6789,N_11163);
and U18243 (N_18243,N_7030,N_9457);
and U18244 (N_18244,N_12389,N_11010);
nand U18245 (N_18245,N_8202,N_8227);
nor U18246 (N_18246,N_9084,N_10598);
or U18247 (N_18247,N_11014,N_6259);
nor U18248 (N_18248,N_9926,N_6851);
or U18249 (N_18249,N_9136,N_8245);
nand U18250 (N_18250,N_10138,N_10200);
nor U18251 (N_18251,N_10655,N_9500);
nor U18252 (N_18252,N_9027,N_8800);
nand U18253 (N_18253,N_6613,N_10034);
or U18254 (N_18254,N_8103,N_12037);
nand U18255 (N_18255,N_8001,N_6801);
nor U18256 (N_18256,N_11564,N_10602);
or U18257 (N_18257,N_9396,N_7584);
nand U18258 (N_18258,N_7603,N_9008);
or U18259 (N_18259,N_9477,N_6749);
or U18260 (N_18260,N_11450,N_9668);
nor U18261 (N_18261,N_7893,N_11696);
or U18262 (N_18262,N_10900,N_10803);
or U18263 (N_18263,N_12145,N_8842);
nand U18264 (N_18264,N_8740,N_10704);
nand U18265 (N_18265,N_12305,N_8300);
or U18266 (N_18266,N_6721,N_12174);
xnor U18267 (N_18267,N_7427,N_10998);
nand U18268 (N_18268,N_11059,N_7771);
and U18269 (N_18269,N_8007,N_11663);
nand U18270 (N_18270,N_11753,N_10499);
or U18271 (N_18271,N_7515,N_9623);
nand U18272 (N_18272,N_9421,N_8363);
and U18273 (N_18273,N_9694,N_7862);
nand U18274 (N_18274,N_11429,N_6741);
and U18275 (N_18275,N_6756,N_7965);
or U18276 (N_18276,N_6840,N_7962);
or U18277 (N_18277,N_11476,N_6588);
nand U18278 (N_18278,N_6295,N_9014);
nand U18279 (N_18279,N_9748,N_8500);
or U18280 (N_18280,N_6631,N_12244);
nor U18281 (N_18281,N_10862,N_7592);
or U18282 (N_18282,N_8461,N_11840);
nor U18283 (N_18283,N_10969,N_6492);
or U18284 (N_18284,N_6325,N_10073);
or U18285 (N_18285,N_11037,N_7806);
or U18286 (N_18286,N_8170,N_11501);
and U18287 (N_18287,N_11646,N_11040);
and U18288 (N_18288,N_10649,N_7272);
or U18289 (N_18289,N_6747,N_8598);
nand U18290 (N_18290,N_9550,N_7528);
nor U18291 (N_18291,N_9110,N_11515);
nor U18292 (N_18292,N_7082,N_11781);
or U18293 (N_18293,N_8289,N_8331);
xor U18294 (N_18294,N_11107,N_9221);
and U18295 (N_18295,N_11613,N_9322);
nor U18296 (N_18296,N_9440,N_9897);
nand U18297 (N_18297,N_9801,N_6572);
nor U18298 (N_18298,N_7546,N_10758);
or U18299 (N_18299,N_7955,N_7429);
or U18300 (N_18300,N_9578,N_7780);
nand U18301 (N_18301,N_12332,N_11484);
xor U18302 (N_18302,N_11466,N_9442);
nor U18303 (N_18303,N_7849,N_10769);
and U18304 (N_18304,N_7933,N_11548);
or U18305 (N_18305,N_8277,N_8934);
or U18306 (N_18306,N_10611,N_8008);
nand U18307 (N_18307,N_8083,N_6833);
nand U18308 (N_18308,N_10492,N_7769);
or U18309 (N_18309,N_7798,N_11093);
or U18310 (N_18310,N_10788,N_10238);
nor U18311 (N_18311,N_9243,N_7645);
and U18312 (N_18312,N_8410,N_11017);
nor U18313 (N_18313,N_12277,N_11599);
xor U18314 (N_18314,N_10158,N_9076);
nand U18315 (N_18315,N_8673,N_8976);
nor U18316 (N_18316,N_10304,N_9158);
or U18317 (N_18317,N_10400,N_11557);
and U18318 (N_18318,N_7297,N_8268);
nand U18319 (N_18319,N_7045,N_9680);
nand U18320 (N_18320,N_8807,N_8932);
nor U18321 (N_18321,N_12320,N_11462);
nand U18322 (N_18322,N_8044,N_11192);
and U18323 (N_18323,N_6385,N_6901);
nor U18324 (N_18324,N_12030,N_12246);
nand U18325 (N_18325,N_11590,N_10444);
xnor U18326 (N_18326,N_11456,N_7692);
nor U18327 (N_18327,N_7133,N_8155);
nor U18328 (N_18328,N_6478,N_11417);
and U18329 (N_18329,N_10454,N_9731);
nor U18330 (N_18330,N_6552,N_8220);
or U18331 (N_18331,N_12056,N_6660);
and U18332 (N_18332,N_9048,N_8822);
or U18333 (N_18333,N_8684,N_7627);
or U18334 (N_18334,N_10452,N_11694);
nor U18335 (N_18335,N_12333,N_9444);
nand U18336 (N_18336,N_12394,N_6999);
or U18337 (N_18337,N_8790,N_10469);
or U18338 (N_18338,N_11184,N_8827);
nand U18339 (N_18339,N_7893,N_10541);
nor U18340 (N_18340,N_8501,N_6741);
nand U18341 (N_18341,N_11369,N_10382);
nand U18342 (N_18342,N_11809,N_12112);
nor U18343 (N_18343,N_6334,N_12353);
or U18344 (N_18344,N_8565,N_7787);
nor U18345 (N_18345,N_11346,N_8231);
and U18346 (N_18346,N_7784,N_11742);
nor U18347 (N_18347,N_6659,N_12157);
nand U18348 (N_18348,N_7374,N_7195);
nand U18349 (N_18349,N_8634,N_7028);
xnor U18350 (N_18350,N_7293,N_7134);
nor U18351 (N_18351,N_12189,N_8804);
xor U18352 (N_18352,N_6706,N_6650);
nor U18353 (N_18353,N_12351,N_6767);
nand U18354 (N_18354,N_9205,N_7623);
and U18355 (N_18355,N_10001,N_11151);
and U18356 (N_18356,N_7444,N_7085);
or U18357 (N_18357,N_7785,N_11195);
and U18358 (N_18358,N_9716,N_12164);
nand U18359 (N_18359,N_8604,N_9104);
nor U18360 (N_18360,N_8279,N_9178);
or U18361 (N_18361,N_10528,N_9001);
or U18362 (N_18362,N_10431,N_11249);
or U18363 (N_18363,N_7040,N_12290);
nand U18364 (N_18364,N_7999,N_8213);
or U18365 (N_18365,N_12149,N_9561);
nor U18366 (N_18366,N_8371,N_8269);
xor U18367 (N_18367,N_10174,N_8935);
nand U18368 (N_18368,N_10135,N_9872);
nand U18369 (N_18369,N_10103,N_8656);
nand U18370 (N_18370,N_7152,N_9392);
and U18371 (N_18371,N_11964,N_9517);
nor U18372 (N_18372,N_10053,N_6678);
nor U18373 (N_18373,N_9765,N_7875);
or U18374 (N_18374,N_9118,N_7461);
or U18375 (N_18375,N_9455,N_11286);
nand U18376 (N_18376,N_8122,N_12136);
and U18377 (N_18377,N_9695,N_11444);
nor U18378 (N_18378,N_8771,N_10509);
or U18379 (N_18379,N_6915,N_6537);
or U18380 (N_18380,N_11107,N_7763);
nor U18381 (N_18381,N_9213,N_7300);
nand U18382 (N_18382,N_10905,N_8400);
and U18383 (N_18383,N_10483,N_11733);
or U18384 (N_18384,N_6714,N_11984);
nand U18385 (N_18385,N_8529,N_10937);
nor U18386 (N_18386,N_12091,N_7060);
and U18387 (N_18387,N_9315,N_6497);
nand U18388 (N_18388,N_10517,N_8329);
and U18389 (N_18389,N_10426,N_11555);
nor U18390 (N_18390,N_9376,N_9091);
and U18391 (N_18391,N_8037,N_6643);
nand U18392 (N_18392,N_12478,N_12222);
nand U18393 (N_18393,N_7723,N_6680);
nand U18394 (N_18394,N_8607,N_10287);
and U18395 (N_18395,N_6806,N_11885);
nor U18396 (N_18396,N_9575,N_11904);
or U18397 (N_18397,N_8748,N_9772);
or U18398 (N_18398,N_7192,N_6569);
or U18399 (N_18399,N_8110,N_8134);
nor U18400 (N_18400,N_11828,N_7977);
or U18401 (N_18401,N_7332,N_12315);
nand U18402 (N_18402,N_11258,N_8808);
or U18403 (N_18403,N_8655,N_10659);
nor U18404 (N_18404,N_8823,N_8495);
and U18405 (N_18405,N_7204,N_10947);
and U18406 (N_18406,N_6478,N_8217);
nor U18407 (N_18407,N_9576,N_8046);
xnor U18408 (N_18408,N_7062,N_8001);
and U18409 (N_18409,N_12334,N_8002);
nand U18410 (N_18410,N_8162,N_9257);
nor U18411 (N_18411,N_11287,N_8108);
nand U18412 (N_18412,N_9928,N_8706);
or U18413 (N_18413,N_7816,N_10668);
or U18414 (N_18414,N_11418,N_7636);
xor U18415 (N_18415,N_10492,N_9305);
nor U18416 (N_18416,N_6370,N_12388);
and U18417 (N_18417,N_12105,N_7651);
nand U18418 (N_18418,N_11284,N_8373);
nor U18419 (N_18419,N_8152,N_8215);
xor U18420 (N_18420,N_9811,N_12275);
nor U18421 (N_18421,N_11353,N_9941);
nand U18422 (N_18422,N_9594,N_9149);
nor U18423 (N_18423,N_11670,N_7766);
nor U18424 (N_18424,N_7718,N_6996);
nor U18425 (N_18425,N_8510,N_6981);
or U18426 (N_18426,N_12105,N_6526);
and U18427 (N_18427,N_10410,N_12339);
nor U18428 (N_18428,N_9509,N_10759);
and U18429 (N_18429,N_7766,N_6476);
and U18430 (N_18430,N_6786,N_6263);
or U18431 (N_18431,N_11325,N_7705);
nand U18432 (N_18432,N_11537,N_11636);
nor U18433 (N_18433,N_7851,N_11624);
nand U18434 (N_18434,N_8093,N_7538);
nor U18435 (N_18435,N_9744,N_12476);
and U18436 (N_18436,N_9822,N_9503);
nor U18437 (N_18437,N_6509,N_6530);
or U18438 (N_18438,N_8864,N_12429);
or U18439 (N_18439,N_9135,N_6615);
nand U18440 (N_18440,N_7289,N_8363);
nand U18441 (N_18441,N_7243,N_10997);
nand U18442 (N_18442,N_10364,N_10517);
or U18443 (N_18443,N_7274,N_7004);
xnor U18444 (N_18444,N_8865,N_9302);
nor U18445 (N_18445,N_12353,N_8940);
and U18446 (N_18446,N_6967,N_9295);
nor U18447 (N_18447,N_10659,N_7350);
nor U18448 (N_18448,N_11115,N_11601);
xnor U18449 (N_18449,N_9043,N_8461);
or U18450 (N_18450,N_8564,N_11076);
nand U18451 (N_18451,N_9294,N_11720);
nand U18452 (N_18452,N_12097,N_7585);
nand U18453 (N_18453,N_9905,N_11061);
and U18454 (N_18454,N_6283,N_11601);
xnor U18455 (N_18455,N_8625,N_8276);
and U18456 (N_18456,N_9542,N_9350);
or U18457 (N_18457,N_10865,N_11841);
and U18458 (N_18458,N_6274,N_9225);
nor U18459 (N_18459,N_9675,N_8981);
nand U18460 (N_18460,N_10709,N_7984);
nand U18461 (N_18461,N_9781,N_10294);
nor U18462 (N_18462,N_6494,N_8545);
nand U18463 (N_18463,N_10414,N_12074);
nand U18464 (N_18464,N_10065,N_11403);
nand U18465 (N_18465,N_11617,N_9134);
nor U18466 (N_18466,N_12065,N_6969);
or U18467 (N_18467,N_8185,N_11885);
nor U18468 (N_18468,N_9091,N_10471);
or U18469 (N_18469,N_9529,N_9279);
nand U18470 (N_18470,N_10159,N_10003);
nand U18471 (N_18471,N_8829,N_9138);
nand U18472 (N_18472,N_8284,N_10321);
or U18473 (N_18473,N_9859,N_9965);
and U18474 (N_18474,N_9937,N_11090);
and U18475 (N_18475,N_11095,N_7392);
nand U18476 (N_18476,N_7947,N_11457);
nor U18477 (N_18477,N_7015,N_6934);
xnor U18478 (N_18478,N_7950,N_7256);
or U18479 (N_18479,N_8178,N_6891);
and U18480 (N_18480,N_8903,N_10443);
nand U18481 (N_18481,N_8306,N_12182);
and U18482 (N_18482,N_7343,N_12160);
or U18483 (N_18483,N_11604,N_6882);
and U18484 (N_18484,N_8355,N_11323);
or U18485 (N_18485,N_11327,N_11222);
nand U18486 (N_18486,N_6896,N_6501);
and U18487 (N_18487,N_7072,N_10585);
and U18488 (N_18488,N_12156,N_10978);
nor U18489 (N_18489,N_7581,N_7334);
or U18490 (N_18490,N_11777,N_10229);
or U18491 (N_18491,N_10544,N_9081);
nand U18492 (N_18492,N_8919,N_12472);
and U18493 (N_18493,N_6755,N_8062);
nand U18494 (N_18494,N_8395,N_7252);
nand U18495 (N_18495,N_9035,N_11501);
or U18496 (N_18496,N_10728,N_7021);
nor U18497 (N_18497,N_6991,N_6467);
nand U18498 (N_18498,N_7645,N_6534);
nand U18499 (N_18499,N_11114,N_7097);
or U18500 (N_18500,N_12053,N_7856);
nand U18501 (N_18501,N_11621,N_6284);
nor U18502 (N_18502,N_7344,N_8340);
nand U18503 (N_18503,N_6627,N_10387);
and U18504 (N_18504,N_8054,N_9134);
and U18505 (N_18505,N_8578,N_8292);
and U18506 (N_18506,N_7122,N_6982);
nor U18507 (N_18507,N_8657,N_7617);
and U18508 (N_18508,N_8513,N_9998);
nand U18509 (N_18509,N_9988,N_7634);
nor U18510 (N_18510,N_11718,N_9066);
nor U18511 (N_18511,N_7389,N_7358);
xnor U18512 (N_18512,N_11900,N_11076);
and U18513 (N_18513,N_8649,N_7775);
or U18514 (N_18514,N_11754,N_7661);
and U18515 (N_18515,N_10497,N_11389);
or U18516 (N_18516,N_8412,N_10259);
or U18517 (N_18517,N_11539,N_8803);
nor U18518 (N_18518,N_12043,N_7826);
nor U18519 (N_18519,N_8824,N_7855);
and U18520 (N_18520,N_10108,N_7462);
or U18521 (N_18521,N_8605,N_10193);
and U18522 (N_18522,N_11655,N_9002);
and U18523 (N_18523,N_11525,N_8901);
nor U18524 (N_18524,N_6624,N_9669);
nor U18525 (N_18525,N_11753,N_9132);
nor U18526 (N_18526,N_11671,N_9641);
nand U18527 (N_18527,N_9104,N_10221);
and U18528 (N_18528,N_11579,N_11377);
nor U18529 (N_18529,N_7263,N_6788);
or U18530 (N_18530,N_9199,N_9339);
or U18531 (N_18531,N_8254,N_11892);
and U18532 (N_18532,N_8232,N_10412);
or U18533 (N_18533,N_10730,N_6363);
xor U18534 (N_18534,N_9226,N_12480);
or U18535 (N_18535,N_7039,N_9295);
nor U18536 (N_18536,N_10979,N_7355);
nand U18537 (N_18537,N_9745,N_11328);
xnor U18538 (N_18538,N_7603,N_8986);
nand U18539 (N_18539,N_8027,N_7912);
nor U18540 (N_18540,N_6998,N_12005);
nand U18541 (N_18541,N_10456,N_11605);
or U18542 (N_18542,N_10664,N_12175);
nor U18543 (N_18543,N_11816,N_11280);
and U18544 (N_18544,N_6770,N_7103);
nand U18545 (N_18545,N_10070,N_12398);
nand U18546 (N_18546,N_10100,N_10473);
or U18547 (N_18547,N_9170,N_9396);
nor U18548 (N_18548,N_7255,N_8854);
and U18549 (N_18549,N_12426,N_7491);
and U18550 (N_18550,N_7699,N_11332);
nand U18551 (N_18551,N_7363,N_11982);
xnor U18552 (N_18552,N_6915,N_11529);
or U18553 (N_18553,N_10776,N_12488);
and U18554 (N_18554,N_10964,N_8561);
xor U18555 (N_18555,N_7654,N_10297);
and U18556 (N_18556,N_10926,N_7278);
nor U18557 (N_18557,N_9005,N_8958);
nor U18558 (N_18558,N_11614,N_10682);
or U18559 (N_18559,N_6329,N_7149);
nand U18560 (N_18560,N_6414,N_7147);
nand U18561 (N_18561,N_8093,N_8252);
nor U18562 (N_18562,N_10298,N_6819);
and U18563 (N_18563,N_9712,N_10737);
and U18564 (N_18564,N_9033,N_9934);
and U18565 (N_18565,N_11028,N_11595);
nor U18566 (N_18566,N_9915,N_7866);
nor U18567 (N_18567,N_10960,N_8472);
nor U18568 (N_18568,N_11213,N_8022);
nand U18569 (N_18569,N_10067,N_7520);
nor U18570 (N_18570,N_8563,N_11166);
and U18571 (N_18571,N_10414,N_11830);
and U18572 (N_18572,N_7979,N_9894);
nand U18573 (N_18573,N_7715,N_10511);
nand U18574 (N_18574,N_6577,N_10356);
nand U18575 (N_18575,N_10449,N_6613);
nand U18576 (N_18576,N_9482,N_7737);
and U18577 (N_18577,N_8446,N_10634);
xor U18578 (N_18578,N_8086,N_10879);
and U18579 (N_18579,N_8507,N_6300);
or U18580 (N_18580,N_9502,N_8211);
nand U18581 (N_18581,N_6544,N_12121);
nor U18582 (N_18582,N_6321,N_10983);
nor U18583 (N_18583,N_6472,N_12068);
xnor U18584 (N_18584,N_11701,N_9956);
and U18585 (N_18585,N_8525,N_10862);
xnor U18586 (N_18586,N_7662,N_12451);
or U18587 (N_18587,N_6938,N_6815);
and U18588 (N_18588,N_7853,N_6392);
and U18589 (N_18589,N_10480,N_12098);
nor U18590 (N_18590,N_11931,N_11829);
xnor U18591 (N_18591,N_10200,N_7623);
nor U18592 (N_18592,N_6712,N_9905);
and U18593 (N_18593,N_8609,N_10225);
or U18594 (N_18594,N_11953,N_9478);
nand U18595 (N_18595,N_10284,N_8951);
nand U18596 (N_18596,N_10780,N_10385);
xor U18597 (N_18597,N_7619,N_8272);
nand U18598 (N_18598,N_11448,N_7302);
nor U18599 (N_18599,N_6449,N_7219);
nand U18600 (N_18600,N_6893,N_11576);
nand U18601 (N_18601,N_8156,N_10508);
and U18602 (N_18602,N_7891,N_10357);
nand U18603 (N_18603,N_11319,N_8315);
xor U18604 (N_18604,N_8521,N_12276);
and U18605 (N_18605,N_9392,N_7772);
and U18606 (N_18606,N_8016,N_12357);
xnor U18607 (N_18607,N_9092,N_7431);
or U18608 (N_18608,N_9916,N_6500);
nor U18609 (N_18609,N_8326,N_6294);
and U18610 (N_18610,N_7691,N_12353);
nand U18611 (N_18611,N_11220,N_12418);
or U18612 (N_18612,N_9814,N_12315);
and U18613 (N_18613,N_9837,N_8553);
or U18614 (N_18614,N_10349,N_9453);
or U18615 (N_18615,N_11981,N_6963);
xnor U18616 (N_18616,N_7217,N_10720);
nor U18617 (N_18617,N_11237,N_8255);
or U18618 (N_18618,N_10279,N_6383);
nor U18619 (N_18619,N_9131,N_8149);
nand U18620 (N_18620,N_7283,N_7400);
nor U18621 (N_18621,N_6643,N_11791);
and U18622 (N_18622,N_7529,N_9338);
and U18623 (N_18623,N_12130,N_9617);
and U18624 (N_18624,N_10163,N_8601);
xor U18625 (N_18625,N_7416,N_9666);
nand U18626 (N_18626,N_9853,N_9407);
or U18627 (N_18627,N_9315,N_12001);
or U18628 (N_18628,N_8871,N_12415);
xor U18629 (N_18629,N_6421,N_6310);
nor U18630 (N_18630,N_7180,N_7619);
xnor U18631 (N_18631,N_8159,N_10924);
or U18632 (N_18632,N_9952,N_11963);
or U18633 (N_18633,N_8900,N_12288);
and U18634 (N_18634,N_11057,N_11448);
nand U18635 (N_18635,N_7932,N_10171);
xor U18636 (N_18636,N_12159,N_10264);
nand U18637 (N_18637,N_9108,N_9752);
nand U18638 (N_18638,N_12275,N_7142);
xnor U18639 (N_18639,N_10388,N_11602);
nand U18640 (N_18640,N_9053,N_10338);
or U18641 (N_18641,N_8163,N_7035);
or U18642 (N_18642,N_7959,N_7332);
nor U18643 (N_18643,N_9354,N_10676);
nor U18644 (N_18644,N_6857,N_9778);
or U18645 (N_18645,N_11722,N_6843);
and U18646 (N_18646,N_6924,N_11879);
or U18647 (N_18647,N_11660,N_9688);
nand U18648 (N_18648,N_9352,N_6387);
or U18649 (N_18649,N_8411,N_10749);
and U18650 (N_18650,N_10202,N_6467);
and U18651 (N_18651,N_12345,N_10368);
xor U18652 (N_18652,N_12376,N_7718);
nand U18653 (N_18653,N_12168,N_9082);
and U18654 (N_18654,N_8590,N_12084);
nor U18655 (N_18655,N_7491,N_9148);
nand U18656 (N_18656,N_10005,N_6902);
nor U18657 (N_18657,N_10004,N_11002);
nand U18658 (N_18658,N_8797,N_6370);
and U18659 (N_18659,N_8023,N_8245);
or U18660 (N_18660,N_7598,N_7910);
nand U18661 (N_18661,N_11954,N_10646);
or U18662 (N_18662,N_8132,N_9623);
nand U18663 (N_18663,N_9214,N_12339);
and U18664 (N_18664,N_8415,N_9589);
and U18665 (N_18665,N_10329,N_9834);
xor U18666 (N_18666,N_12103,N_11310);
nand U18667 (N_18667,N_8378,N_8311);
and U18668 (N_18668,N_9914,N_9070);
and U18669 (N_18669,N_8213,N_7460);
and U18670 (N_18670,N_12292,N_9288);
or U18671 (N_18671,N_11271,N_11626);
and U18672 (N_18672,N_8552,N_6287);
and U18673 (N_18673,N_9869,N_7071);
nand U18674 (N_18674,N_10611,N_8735);
nand U18675 (N_18675,N_8938,N_12015);
and U18676 (N_18676,N_7630,N_9196);
nor U18677 (N_18677,N_7895,N_7312);
and U18678 (N_18678,N_11438,N_9291);
and U18679 (N_18679,N_6709,N_12389);
nor U18680 (N_18680,N_9383,N_11427);
nor U18681 (N_18681,N_9240,N_7785);
or U18682 (N_18682,N_12271,N_9765);
or U18683 (N_18683,N_10566,N_10129);
nand U18684 (N_18684,N_9039,N_11947);
nand U18685 (N_18685,N_11542,N_7350);
and U18686 (N_18686,N_11873,N_12158);
xnor U18687 (N_18687,N_10652,N_11590);
and U18688 (N_18688,N_10310,N_10935);
and U18689 (N_18689,N_9900,N_9933);
xnor U18690 (N_18690,N_8189,N_9919);
nand U18691 (N_18691,N_10231,N_8468);
nand U18692 (N_18692,N_11084,N_7530);
and U18693 (N_18693,N_7929,N_10014);
nand U18694 (N_18694,N_6408,N_11749);
nand U18695 (N_18695,N_7808,N_11008);
nand U18696 (N_18696,N_8521,N_10805);
or U18697 (N_18697,N_7001,N_7665);
nor U18698 (N_18698,N_6561,N_11990);
or U18699 (N_18699,N_7296,N_11458);
and U18700 (N_18700,N_6988,N_7264);
nand U18701 (N_18701,N_9282,N_6409);
nand U18702 (N_18702,N_10660,N_7355);
nand U18703 (N_18703,N_11429,N_6455);
nand U18704 (N_18704,N_7450,N_11038);
and U18705 (N_18705,N_12364,N_6803);
nand U18706 (N_18706,N_7191,N_9719);
and U18707 (N_18707,N_8174,N_7954);
or U18708 (N_18708,N_7892,N_8156);
or U18709 (N_18709,N_10541,N_7599);
xor U18710 (N_18710,N_10201,N_10294);
or U18711 (N_18711,N_11757,N_8969);
nand U18712 (N_18712,N_8750,N_7692);
or U18713 (N_18713,N_11410,N_8562);
nor U18714 (N_18714,N_9863,N_11579);
or U18715 (N_18715,N_7466,N_10067);
or U18716 (N_18716,N_11833,N_10233);
or U18717 (N_18717,N_8172,N_7001);
xor U18718 (N_18718,N_6691,N_10209);
and U18719 (N_18719,N_8858,N_6286);
nand U18720 (N_18720,N_11957,N_9002);
xnor U18721 (N_18721,N_7009,N_10347);
nand U18722 (N_18722,N_11874,N_7230);
nand U18723 (N_18723,N_8669,N_9087);
nand U18724 (N_18724,N_11584,N_6862);
and U18725 (N_18725,N_10651,N_7853);
nand U18726 (N_18726,N_9698,N_11051);
nor U18727 (N_18727,N_11267,N_6289);
or U18728 (N_18728,N_9320,N_11941);
and U18729 (N_18729,N_9496,N_10353);
or U18730 (N_18730,N_10709,N_9517);
nor U18731 (N_18731,N_7501,N_9467);
or U18732 (N_18732,N_9170,N_10254);
and U18733 (N_18733,N_11838,N_8206);
nor U18734 (N_18734,N_7785,N_8253);
or U18735 (N_18735,N_11051,N_10462);
nand U18736 (N_18736,N_8791,N_10002);
nor U18737 (N_18737,N_6933,N_6715);
nor U18738 (N_18738,N_10382,N_9378);
nor U18739 (N_18739,N_10726,N_6798);
nand U18740 (N_18740,N_7843,N_8073);
and U18741 (N_18741,N_9440,N_8589);
nor U18742 (N_18742,N_9862,N_12043);
nand U18743 (N_18743,N_11328,N_9232);
nand U18744 (N_18744,N_11327,N_12432);
nor U18745 (N_18745,N_9261,N_9694);
and U18746 (N_18746,N_8821,N_10084);
nand U18747 (N_18747,N_11356,N_11057);
or U18748 (N_18748,N_9545,N_8616);
nand U18749 (N_18749,N_12278,N_11771);
or U18750 (N_18750,N_18001,N_16757);
or U18751 (N_18751,N_13126,N_15015);
nand U18752 (N_18752,N_18013,N_12779);
xor U18753 (N_18753,N_13713,N_18442);
nor U18754 (N_18754,N_17215,N_13057);
and U18755 (N_18755,N_17778,N_14376);
nand U18756 (N_18756,N_16551,N_15480);
nand U18757 (N_18757,N_16565,N_14280);
or U18758 (N_18758,N_15950,N_17538);
nand U18759 (N_18759,N_13718,N_13089);
nand U18760 (N_18760,N_17590,N_18054);
and U18761 (N_18761,N_14749,N_14578);
nor U18762 (N_18762,N_16560,N_17807);
or U18763 (N_18763,N_14351,N_13213);
nand U18764 (N_18764,N_15615,N_18746);
nor U18765 (N_18765,N_18171,N_13929);
and U18766 (N_18766,N_14235,N_18566);
and U18767 (N_18767,N_14379,N_16815);
or U18768 (N_18768,N_13990,N_12804);
nor U18769 (N_18769,N_15092,N_12818);
or U18770 (N_18770,N_15721,N_14731);
nor U18771 (N_18771,N_16221,N_12917);
nor U18772 (N_18772,N_18413,N_14173);
nor U18773 (N_18773,N_18188,N_13384);
or U18774 (N_18774,N_14354,N_16018);
and U18775 (N_18775,N_16979,N_18600);
nor U18776 (N_18776,N_18497,N_15418);
or U18777 (N_18777,N_17532,N_12553);
nand U18778 (N_18778,N_16228,N_16981);
nor U18779 (N_18779,N_16725,N_12574);
and U18780 (N_18780,N_14147,N_17574);
xor U18781 (N_18781,N_15650,N_15226);
nand U18782 (N_18782,N_14932,N_13771);
and U18783 (N_18783,N_16761,N_16220);
or U18784 (N_18784,N_17890,N_15653);
nor U18785 (N_18785,N_15891,N_18341);
or U18786 (N_18786,N_13515,N_17711);
and U18787 (N_18787,N_12714,N_12706);
xor U18788 (N_18788,N_15608,N_17994);
nor U18789 (N_18789,N_13081,N_14311);
nor U18790 (N_18790,N_15422,N_14246);
xnor U18791 (N_18791,N_14163,N_15325);
nor U18792 (N_18792,N_18129,N_14446);
or U18793 (N_18793,N_15511,N_13304);
nand U18794 (N_18794,N_16192,N_17784);
nor U18795 (N_18795,N_15172,N_13590);
nand U18796 (N_18796,N_17955,N_12911);
nor U18797 (N_18797,N_15460,N_16826);
or U18798 (N_18798,N_14229,N_16919);
nand U18799 (N_18799,N_15924,N_16145);
nor U18800 (N_18800,N_18564,N_13773);
nor U18801 (N_18801,N_16582,N_15023);
nand U18802 (N_18802,N_16686,N_15473);
and U18803 (N_18803,N_17392,N_12775);
and U18804 (N_18804,N_15256,N_18205);
nand U18805 (N_18805,N_13720,N_13215);
nand U18806 (N_18806,N_17282,N_13312);
and U18807 (N_18807,N_15934,N_18072);
and U18808 (N_18808,N_16428,N_13988);
nor U18809 (N_18809,N_15348,N_18272);
and U18810 (N_18810,N_16201,N_14650);
or U18811 (N_18811,N_18379,N_16467);
or U18812 (N_18812,N_14337,N_18715);
and U18813 (N_18813,N_13759,N_15812);
or U18814 (N_18814,N_15058,N_16967);
or U18815 (N_18815,N_14460,N_18386);
nand U18816 (N_18816,N_13667,N_18217);
nand U18817 (N_18817,N_13227,N_13795);
nor U18818 (N_18818,N_13747,N_14372);
xnor U18819 (N_18819,N_17238,N_14560);
nand U18820 (N_18820,N_12921,N_16514);
or U18821 (N_18821,N_14634,N_14730);
and U18822 (N_18822,N_15397,N_14582);
nor U18823 (N_18823,N_18690,N_18436);
xor U18824 (N_18824,N_15635,N_13102);
nand U18825 (N_18825,N_14146,N_15941);
and U18826 (N_18826,N_16375,N_18077);
nor U18827 (N_18827,N_15423,N_17750);
xnor U18828 (N_18828,N_15042,N_17325);
nor U18829 (N_18829,N_17548,N_15006);
nand U18830 (N_18830,N_14097,N_13121);
or U18831 (N_18831,N_18563,N_14444);
or U18832 (N_18832,N_13758,N_17013);
nand U18833 (N_18833,N_17329,N_16391);
xnor U18834 (N_18834,N_13365,N_14334);
and U18835 (N_18835,N_14814,N_16903);
nand U18836 (N_18836,N_15755,N_14603);
and U18837 (N_18837,N_13356,N_13722);
nor U18838 (N_18838,N_13674,N_18455);
nand U18839 (N_18839,N_15384,N_16412);
or U18840 (N_18840,N_12816,N_15328);
nand U18841 (N_18841,N_14174,N_17424);
and U18842 (N_18842,N_16676,N_18042);
xor U18843 (N_18843,N_17557,N_13306);
or U18844 (N_18844,N_13279,N_17892);
nor U18845 (N_18845,N_16935,N_15558);
xnor U18846 (N_18846,N_15477,N_14487);
nor U18847 (N_18847,N_15931,N_16341);
or U18848 (N_18848,N_13011,N_14793);
and U18849 (N_18849,N_15593,N_16732);
nand U18850 (N_18850,N_16406,N_12606);
and U18851 (N_18851,N_15377,N_16189);
or U18852 (N_18852,N_16944,N_17469);
and U18853 (N_18853,N_15508,N_12947);
nand U18854 (N_18854,N_15543,N_16961);
and U18855 (N_18855,N_15569,N_18731);
and U18856 (N_18856,N_14298,N_14131);
and U18857 (N_18857,N_18457,N_16175);
and U18858 (N_18858,N_13687,N_15989);
nand U18859 (N_18859,N_15907,N_16785);
nor U18860 (N_18860,N_13800,N_14028);
nor U18861 (N_18861,N_12658,N_13769);
and U18862 (N_18862,N_18370,N_16136);
or U18863 (N_18863,N_17034,N_14906);
and U18864 (N_18864,N_14179,N_18190);
nor U18865 (N_18865,N_16419,N_12646);
or U18866 (N_18866,N_16035,N_17655);
nor U18867 (N_18867,N_16061,N_15400);
or U18868 (N_18868,N_15548,N_16152);
and U18869 (N_18869,N_16772,N_12675);
nand U18870 (N_18870,N_17736,N_13613);
nand U18871 (N_18871,N_16150,N_18583);
nor U18872 (N_18872,N_15126,N_15114);
nor U18873 (N_18873,N_16272,N_13174);
nand U18874 (N_18874,N_14570,N_17159);
and U18875 (N_18875,N_16704,N_12830);
nand U18876 (N_18876,N_17684,N_12869);
or U18877 (N_18877,N_16767,N_16888);
nor U18878 (N_18878,N_18433,N_14054);
xor U18879 (N_18879,N_17797,N_16382);
and U18880 (N_18880,N_14273,N_13396);
nor U18881 (N_18881,N_16318,N_16075);
nand U18882 (N_18882,N_18157,N_16884);
and U18883 (N_18883,N_14881,N_14382);
and U18884 (N_18884,N_13432,N_12871);
nand U18885 (N_18885,N_16791,N_14405);
or U18886 (N_18886,N_17415,N_12694);
and U18887 (N_18887,N_15312,N_15562);
xnor U18888 (N_18888,N_14953,N_16524);
nand U18889 (N_18889,N_13302,N_17222);
or U18890 (N_18890,N_15016,N_15297);
nor U18891 (N_18891,N_18395,N_14544);
and U18892 (N_18892,N_13437,N_14787);
and U18893 (N_18893,N_12718,N_14595);
nor U18894 (N_18894,N_13748,N_14773);
nor U18895 (N_18895,N_18009,N_17136);
and U18896 (N_18896,N_13949,N_18606);
or U18897 (N_18897,N_12596,N_18582);
or U18898 (N_18898,N_14159,N_15957);
nor U18899 (N_18899,N_15174,N_14457);
nor U18900 (N_18900,N_17318,N_17187);
nand U18901 (N_18901,N_17486,N_13071);
nor U18902 (N_18902,N_15388,N_17359);
nand U18903 (N_18903,N_15579,N_16950);
nand U18904 (N_18904,N_12595,N_14277);
nor U18905 (N_18905,N_18404,N_17076);
or U18906 (N_18906,N_13831,N_18422);
nand U18907 (N_18907,N_15402,N_12860);
nor U18908 (N_18908,N_15223,N_12879);
or U18909 (N_18909,N_17959,N_14997);
and U18910 (N_18910,N_14085,N_14872);
and U18911 (N_18911,N_15049,N_13609);
nand U18912 (N_18912,N_12685,N_15251);
or U18913 (N_18913,N_17310,N_14503);
nor U18914 (N_18914,N_15401,N_13061);
or U18915 (N_18915,N_16157,N_17271);
nor U18916 (N_18916,N_14770,N_17537);
or U18917 (N_18917,N_16636,N_13222);
and U18918 (N_18918,N_14133,N_17833);
nor U18919 (N_18919,N_13110,N_13340);
or U18920 (N_18920,N_16459,N_16069);
or U18921 (N_18921,N_13267,N_16254);
and U18922 (N_18922,N_14732,N_15778);
or U18923 (N_18923,N_14200,N_14576);
xor U18924 (N_18924,N_12835,N_15913);
nor U18925 (N_18925,N_12841,N_14960);
and U18926 (N_18926,N_15280,N_15117);
nand U18927 (N_18927,N_14859,N_14109);
nor U18928 (N_18928,N_17827,N_18440);
nand U18929 (N_18929,N_16561,N_16968);
or U18930 (N_18930,N_16444,N_18514);
and U18931 (N_18931,N_17811,N_13927);
and U18932 (N_18932,N_14096,N_16352);
nor U18933 (N_18933,N_14804,N_13852);
or U18934 (N_18934,N_13010,N_14862);
and U18935 (N_18935,N_18451,N_12727);
or U18936 (N_18936,N_13042,N_16842);
or U18937 (N_18937,N_13192,N_13236);
nand U18938 (N_18938,N_16945,N_15082);
or U18939 (N_18939,N_15303,N_14031);
nor U18940 (N_18940,N_16737,N_13456);
nor U18941 (N_18941,N_13162,N_14002);
xor U18942 (N_18942,N_14661,N_13987);
and U18943 (N_18943,N_16269,N_14417);
and U18944 (N_18944,N_16777,N_18398);
nor U18945 (N_18945,N_15000,N_14583);
nor U18946 (N_18946,N_17726,N_16806);
and U18947 (N_18947,N_15761,N_15043);
xor U18948 (N_18948,N_13600,N_17733);
nand U18949 (N_18949,N_12619,N_13832);
xnor U18950 (N_18950,N_13763,N_14025);
or U18951 (N_18951,N_14126,N_13185);
nor U18952 (N_18952,N_15492,N_13893);
nand U18953 (N_18953,N_18145,N_15440);
nand U18954 (N_18954,N_16520,N_18504);
or U18955 (N_18955,N_16566,N_12704);
or U18956 (N_18956,N_14892,N_18076);
or U18957 (N_18957,N_17394,N_16040);
or U18958 (N_18958,N_12914,N_17581);
or U18959 (N_18959,N_14371,N_16258);
and U18960 (N_18960,N_18461,N_14300);
nand U18961 (N_18961,N_14389,N_17041);
and U18962 (N_18962,N_15343,N_14907);
nand U18963 (N_18963,N_13237,N_18026);
xor U18964 (N_18964,N_12577,N_14984);
xor U18965 (N_18965,N_12974,N_17279);
nand U18966 (N_18966,N_14495,N_16699);
and U18967 (N_18967,N_17080,N_15190);
nand U18968 (N_18968,N_16538,N_18527);
nor U18969 (N_18969,N_15363,N_14339);
or U18970 (N_18970,N_15969,N_14077);
or U18971 (N_18971,N_17297,N_17243);
nand U18972 (N_18972,N_15220,N_18028);
nand U18973 (N_18973,N_15025,N_14328);
nand U18974 (N_18974,N_17978,N_16782);
or U18975 (N_18975,N_17549,N_15475);
or U18976 (N_18976,N_14890,N_16581);
or U18977 (N_18977,N_14699,N_12569);
nor U18978 (N_18978,N_13064,N_13498);
or U18979 (N_18979,N_13801,N_18518);
or U18980 (N_18980,N_15541,N_16377);
and U18981 (N_18981,N_18172,N_15064);
nor U18982 (N_18982,N_17450,N_14939);
nand U18983 (N_18983,N_14817,N_17308);
or U18984 (N_18984,N_17506,N_17082);
xor U18985 (N_18985,N_14805,N_12853);
nor U18986 (N_18986,N_17613,N_13277);
or U18987 (N_18987,N_16172,N_18397);
nand U18988 (N_18988,N_18195,N_17189);
nor U18989 (N_18989,N_15102,N_13080);
nor U18990 (N_18990,N_14736,N_15740);
and U18991 (N_18991,N_17909,N_16879);
or U18992 (N_18992,N_17249,N_16568);
or U18993 (N_18993,N_16947,N_17058);
nor U18994 (N_18994,N_18718,N_18599);
nand U18995 (N_18995,N_14908,N_17993);
and U18996 (N_18996,N_17017,N_16146);
or U18997 (N_18997,N_12702,N_13673);
and U18998 (N_18998,N_13779,N_18558);
and U18999 (N_18999,N_15002,N_14998);
nand U19000 (N_19000,N_15210,N_15858);
nor U19001 (N_19001,N_15130,N_14245);
or U19002 (N_19002,N_15054,N_12758);
xor U19003 (N_19003,N_17838,N_16359);
xor U19004 (N_19004,N_18260,N_17004);
xnor U19005 (N_19005,N_16197,N_18315);
nor U19006 (N_19006,N_13149,N_12684);
nor U19007 (N_19007,N_17264,N_18732);
and U19008 (N_19008,N_15347,N_18034);
nand U19009 (N_19009,N_12651,N_13039);
and U19010 (N_19010,N_13316,N_15385);
or U19011 (N_19011,N_13416,N_13349);
and U19012 (N_19012,N_13863,N_17488);
and U19013 (N_19013,N_17155,N_14122);
nand U19014 (N_19014,N_18151,N_18048);
nand U19015 (N_19015,N_12943,N_17698);
or U19016 (N_19016,N_17651,N_13723);
or U19017 (N_19017,N_12956,N_14264);
and U19018 (N_19018,N_15727,N_18131);
nand U19019 (N_19019,N_17974,N_14427);
and U19020 (N_19020,N_14909,N_14669);
or U19021 (N_19021,N_18356,N_17597);
nand U19022 (N_19022,N_13965,N_13682);
or U19023 (N_19023,N_16182,N_16063);
and U19024 (N_19024,N_14747,N_17630);
nand U19025 (N_19025,N_18268,N_13596);
and U19026 (N_19026,N_13593,N_13344);
or U19027 (N_19027,N_13642,N_15809);
nor U19028 (N_19028,N_17812,N_14424);
nand U19029 (N_19029,N_17167,N_18029);
nor U19030 (N_19030,N_15021,N_18194);
nand U19031 (N_19031,N_17500,N_18424);
nand U19032 (N_19032,N_13226,N_17077);
or U19033 (N_19033,N_18682,N_13335);
and U19034 (N_19034,N_15779,N_17771);
nor U19035 (N_19035,N_14477,N_13211);
nand U19036 (N_19036,N_15176,N_14754);
nor U19037 (N_19037,N_15928,N_13989);
nor U19038 (N_19038,N_18317,N_18472);
nand U19039 (N_19039,N_17051,N_12898);
and U19040 (N_19040,N_17610,N_12886);
nor U19041 (N_19041,N_18307,N_13083);
xnor U19042 (N_19042,N_12550,N_13150);
and U19043 (N_19043,N_13133,N_16690);
nor U19044 (N_19044,N_14409,N_16165);
nor U19045 (N_19045,N_14256,N_17332);
nor U19046 (N_19046,N_15586,N_17104);
and U19047 (N_19047,N_15072,N_13239);
nor U19048 (N_19048,N_13631,N_13347);
or U19049 (N_19049,N_15390,N_18320);
xnor U19050 (N_19050,N_17036,N_18096);
nor U19051 (N_19051,N_13997,N_17043);
xor U19052 (N_19052,N_14589,N_15603);
nand U19053 (N_19053,N_15655,N_18209);
and U19054 (N_19054,N_13700,N_15732);
or U19055 (N_19055,N_17948,N_15182);
nor U19056 (N_19056,N_13560,N_13964);
and U19057 (N_19057,N_13789,N_15419);
nor U19058 (N_19058,N_18687,N_18154);
xor U19059 (N_19059,N_16742,N_18488);
nand U19060 (N_19060,N_14592,N_13607);
nand U19061 (N_19061,N_14462,N_18184);
nor U19062 (N_19062,N_16917,N_14130);
nand U19063 (N_19063,N_15860,N_14851);
nor U19064 (N_19064,N_17951,N_17177);
xnor U19065 (N_19065,N_18281,N_14240);
or U19066 (N_19066,N_13892,N_12861);
or U19067 (N_19067,N_14515,N_15916);
and U19068 (N_19068,N_13294,N_15451);
nor U19069 (N_19069,N_14826,N_18490);
nand U19070 (N_19070,N_14100,N_14275);
or U19071 (N_19071,N_15330,N_12541);
nor U19072 (N_19072,N_17687,N_17773);
nand U19073 (N_19073,N_17011,N_15164);
nor U19074 (N_19074,N_16353,N_14464);
and U19075 (N_19075,N_13630,N_15300);
and U19076 (N_19076,N_16971,N_13881);
and U19077 (N_19077,N_17512,N_16763);
or U19078 (N_19078,N_14492,N_17089);
nor U19079 (N_19079,N_15085,N_15096);
nand U19080 (N_19080,N_13444,N_13178);
or U19081 (N_19081,N_14050,N_17765);
nand U19082 (N_19082,N_12923,N_12753);
nor U19083 (N_19083,N_16759,N_12600);
and U19084 (N_19084,N_18729,N_14992);
and U19085 (N_19085,N_15730,N_17605);
or U19086 (N_19086,N_12647,N_17130);
nand U19087 (N_19087,N_14250,N_12994);
or U19088 (N_19088,N_17563,N_14566);
nand U19089 (N_19089,N_16092,N_14741);
nand U19090 (N_19090,N_13310,N_17591);
or U19091 (N_19091,N_15531,N_17385);
nand U19092 (N_19092,N_12629,N_14480);
nand U19093 (N_19093,N_16618,N_15571);
nor U19094 (N_19094,N_17566,N_12625);
or U19095 (N_19095,N_13287,N_13669);
and U19096 (N_19096,N_18623,N_16628);
nor U19097 (N_19097,N_13455,N_16647);
and U19098 (N_19098,N_17665,N_15867);
and U19099 (N_19099,N_17576,N_16276);
nor U19100 (N_19100,N_13562,N_16550);
nor U19101 (N_19101,N_16003,N_18266);
or U19102 (N_19102,N_14542,N_13041);
xor U19103 (N_19103,N_13292,N_17119);
xor U19104 (N_19104,N_16873,N_16946);
or U19105 (N_19105,N_17923,N_16710);
nand U19106 (N_19106,N_12538,N_14190);
nor U19107 (N_19107,N_13050,N_16768);
nand U19108 (N_19108,N_16294,N_17348);
or U19109 (N_19109,N_17409,N_16207);
or U19110 (N_19110,N_13129,N_17523);
or U19111 (N_19111,N_18705,N_12975);
nand U19112 (N_19112,N_15152,N_12616);
xnor U19113 (N_19113,N_14894,N_13357);
nor U19114 (N_19114,N_12833,N_14467);
xor U19115 (N_19115,N_13030,N_13670);
xor U19116 (N_19116,N_16702,N_15289);
or U19117 (N_19117,N_12828,N_12690);
nand U19118 (N_19118,N_17161,N_15522);
or U19119 (N_19119,N_17545,N_14105);
xnor U19120 (N_19120,N_17416,N_17455);
nand U19121 (N_19121,N_16389,N_15972);
nor U19122 (N_19122,N_15920,N_15825);
and U19123 (N_19123,N_14744,N_17776);
or U19124 (N_19124,N_15718,N_16864);
nand U19125 (N_19125,N_14185,N_17304);
and U19126 (N_19126,N_15794,N_13439);
or U19127 (N_19127,N_13821,N_18605);
or U19128 (N_19128,N_17268,N_15372);
or U19129 (N_19129,N_12854,N_17103);
and U19130 (N_19130,N_15366,N_13341);
and U19131 (N_19131,N_16408,N_18291);
nand U19132 (N_19132,N_16277,N_13691);
and U19133 (N_19133,N_17096,N_13115);
nor U19134 (N_19134,N_14587,N_14509);
and U19135 (N_19135,N_18575,N_17091);
and U19136 (N_19136,N_15748,N_13686);
nand U19137 (N_19137,N_16173,N_16425);
nand U19138 (N_19138,N_13745,N_15238);
or U19139 (N_19139,N_13399,N_16205);
and U19140 (N_19140,N_13935,N_12973);
nor U19141 (N_19141,N_17072,N_17299);
nor U19142 (N_19142,N_12958,N_14990);
nor U19143 (N_19143,N_16264,N_15613);
nor U19144 (N_19144,N_14186,N_17127);
xor U19145 (N_19145,N_15367,N_14531);
or U19146 (N_19146,N_17256,N_14365);
nand U19147 (N_19147,N_15902,N_14420);
and U19148 (N_19148,N_13876,N_12701);
xnor U19149 (N_19149,N_18537,N_18263);
nor U19150 (N_19150,N_14194,N_13838);
nor U19151 (N_19151,N_14244,N_17367);
xnor U19152 (N_19152,N_16736,N_15131);
nor U19153 (N_19153,N_15617,N_16854);
nor U19154 (N_19154,N_14392,N_13376);
nor U19155 (N_19155,N_15457,N_14434);
or U19156 (N_19156,N_18337,N_17746);
or U19157 (N_19157,N_13329,N_12597);
and U19158 (N_19158,N_14837,N_14553);
nor U19159 (N_19159,N_18158,N_17973);
and U19160 (N_19160,N_16666,N_16852);
and U19161 (N_19161,N_16999,N_13666);
or U19162 (N_19162,N_14694,N_12862);
xor U19163 (N_19163,N_17937,N_13181);
nand U19164 (N_19164,N_15693,N_14935);
nor U19165 (N_19165,N_13303,N_13201);
nor U19166 (N_19166,N_17719,N_17380);
xnor U19167 (N_19167,N_16278,N_12724);
and U19168 (N_19168,N_15573,N_16251);
xnor U19169 (N_19169,N_13262,N_16310);
nor U19170 (N_19170,N_13210,N_14317);
or U19171 (N_19171,N_18292,N_17060);
nand U19172 (N_19172,N_12990,N_16706);
xor U19173 (N_19173,N_15675,N_18432);
nand U19174 (N_19174,N_15699,N_14548);
or U19175 (N_19175,N_16536,N_17867);
and U19176 (N_19176,N_13326,N_15884);
nand U19177 (N_19177,N_17620,N_13246);
nor U19178 (N_19178,N_14400,N_17910);
nand U19179 (N_19179,N_14700,N_16698);
or U19180 (N_19180,N_14323,N_16349);
nand U19181 (N_19181,N_18668,N_17427);
xor U19182 (N_19182,N_12518,N_15476);
nor U19183 (N_19183,N_17477,N_14683);
nor U19184 (N_19184,N_17115,N_14774);
and U19185 (N_19185,N_13558,N_18528);
nand U19186 (N_19186,N_12623,N_17965);
xnor U19187 (N_19187,N_15464,N_14670);
or U19188 (N_19188,N_14219,N_14110);
nor U19189 (N_19189,N_18607,N_15956);
xor U19190 (N_19190,N_13910,N_18742);
or U19191 (N_19191,N_16273,N_18749);
and U19192 (N_19192,N_15189,N_13123);
nand U19193 (N_19193,N_14029,N_16436);
nor U19194 (N_19194,N_14234,N_15607);
nand U19195 (N_19195,N_14196,N_13904);
nor U19196 (N_19196,N_15667,N_14547);
and U19197 (N_19197,N_18290,N_14459);
nor U19198 (N_19198,N_14075,N_14534);
or U19199 (N_19199,N_15212,N_12952);
nand U19200 (N_19200,N_14880,N_14698);
nor U19201 (N_19201,N_17025,N_16841);
nor U19202 (N_19202,N_17242,N_16682);
or U19203 (N_19203,N_17558,N_16174);
and U19204 (N_19204,N_17642,N_16982);
or U19205 (N_19205,N_15873,N_17259);
nand U19206 (N_19206,N_15369,N_18373);
or U19207 (N_19207,N_14377,N_13531);
or U19208 (N_19208,N_13533,N_14713);
or U19209 (N_19209,N_18653,N_16198);
nand U19210 (N_19210,N_15029,N_15915);
and U19211 (N_19211,N_15455,N_16107);
and U19212 (N_19212,N_16091,N_15336);
and U19213 (N_19213,N_16577,N_14220);
or U19214 (N_19214,N_18596,N_15877);
or U19215 (N_19215,N_16866,N_15888);
nand U19216 (N_19216,N_14089,N_16911);
and U19217 (N_19217,N_18415,N_15012);
nand U19218 (N_19218,N_14419,N_15782);
or U19219 (N_19219,N_14211,N_18123);
nor U19220 (N_19220,N_16505,N_13621);
xor U19221 (N_19221,N_14523,N_13180);
nand U19222 (N_19222,N_14915,N_13730);
and U19223 (N_19223,N_15820,N_15099);
xnor U19224 (N_19224,N_18547,N_13905);
or U19225 (N_19225,N_14291,N_13706);
nand U19226 (N_19226,N_12846,N_14154);
nor U19227 (N_19227,N_17499,N_13858);
and U19228 (N_19228,N_13214,N_13566);
or U19229 (N_19229,N_15799,N_13233);
nand U19230 (N_19230,N_17755,N_12807);
nor U19231 (N_19231,N_13783,N_15037);
nor U19232 (N_19232,N_18008,N_13827);
or U19233 (N_19233,N_14201,N_16515);
nand U19234 (N_19234,N_13373,N_15501);
nor U19235 (N_19235,N_15081,N_13418);
and U19236 (N_19236,N_16874,N_16455);
nand U19237 (N_19237,N_15895,N_14118);
nand U19238 (N_19238,N_12893,N_13088);
xor U19239 (N_19239,N_15345,N_14175);
and U19240 (N_19240,N_13029,N_17671);
or U19241 (N_19241,N_18142,N_17519);
and U19242 (N_19242,N_13378,N_14301);
nor U19243 (N_19243,N_12649,N_18085);
or U19244 (N_19244,N_18481,N_17411);
or U19245 (N_19245,N_17122,N_13293);
xnor U19246 (N_19246,N_17033,N_17203);
nor U19247 (N_19247,N_17522,N_16062);
and U19248 (N_19248,N_12903,N_13822);
or U19249 (N_19249,N_16929,N_16103);
nor U19250 (N_19250,N_15252,N_16367);
xor U19251 (N_19251,N_12645,N_16334);
or U19252 (N_19252,N_18246,N_16064);
and U19253 (N_19253,N_16593,N_15089);
nor U19254 (N_19254,N_17992,N_15765);
or U19255 (N_19255,N_14797,N_13944);
nor U19256 (N_19256,N_12571,N_17975);
nor U19257 (N_19257,N_15070,N_14266);
and U19258 (N_19258,N_15599,N_14320);
and U19259 (N_19259,N_16877,N_14846);
nand U19260 (N_19260,N_16265,N_13836);
or U19261 (N_19261,N_16398,N_15266);
nor U19262 (N_19262,N_14384,N_14139);
or U19263 (N_19263,N_17889,N_16719);
xnor U19264 (N_19264,N_17200,N_13047);
xor U19265 (N_19265,N_17603,N_14760);
nor U19266 (N_19266,N_17403,N_16304);
and U19267 (N_19267,N_15900,N_15341);
nand U19268 (N_19268,N_13204,N_15896);
or U19269 (N_19269,N_17426,N_12928);
nor U19270 (N_19270,N_13013,N_13327);
and U19271 (N_19271,N_18423,N_15807);
nand U19272 (N_19272,N_12508,N_15241);
or U19273 (N_19273,N_14343,N_17810);
nor U19274 (N_19274,N_18574,N_16513);
nor U19275 (N_19275,N_15985,N_17042);
nor U19276 (N_19276,N_15656,N_15640);
nor U19277 (N_19277,N_14135,N_17539);
nand U19278 (N_19278,N_13971,N_18097);
and U19279 (N_19279,N_14202,N_13695);
nand U19280 (N_19280,N_14475,N_15033);
and U19281 (N_19281,N_13941,N_16009);
nor U19282 (N_19282,N_13681,N_16792);
nor U19283 (N_19283,N_14994,N_16199);
or U19284 (N_19284,N_18345,N_13726);
nor U19285 (N_19285,N_12700,N_12847);
and U19286 (N_19286,N_16282,N_16141);
and U19287 (N_19287,N_12900,N_15165);
nand U19288 (N_19288,N_16379,N_13177);
nor U19289 (N_19289,N_17633,N_12584);
nor U19290 (N_19290,N_13238,N_13054);
or U19291 (N_19291,N_14326,N_16602);
and U19292 (N_19292,N_17657,N_17204);
and U19293 (N_19293,N_17387,N_14818);
and U19294 (N_19294,N_14819,N_14092);
or U19295 (N_19295,N_18000,N_12882);
nand U19296 (N_19296,N_18383,N_14090);
or U19297 (N_19297,N_15071,N_15703);
nor U19298 (N_19298,N_18595,N_14058);
and U19299 (N_19299,N_14671,N_13074);
nor U19300 (N_19300,N_15745,N_18019);
nor U19301 (N_19301,N_17199,N_13954);
and U19302 (N_19302,N_13622,N_13724);
nand U19303 (N_19303,N_18628,N_13077);
xor U19304 (N_19304,N_15835,N_15236);
nand U19305 (N_19305,N_13475,N_16203);
and U19306 (N_19306,N_16701,N_13507);
and U19307 (N_19307,N_17421,N_15798);
nor U19308 (N_19308,N_13043,N_14068);
nor U19309 (N_19309,N_16196,N_12558);
or U19310 (N_19310,N_16717,N_13656);
and U19311 (N_19311,N_13519,N_12757);
or U19312 (N_19312,N_18725,N_18658);
and U19313 (N_19313,N_12930,N_13460);
nand U19314 (N_19314,N_13052,N_15735);
and U19315 (N_19315,N_14864,N_16769);
and U19316 (N_19316,N_15179,N_13424);
nand U19317 (N_19317,N_18274,N_13807);
and U19318 (N_19318,N_16237,N_17735);
nand U19319 (N_19319,N_15068,N_14293);
nor U19320 (N_19320,N_17090,N_13886);
nand U19321 (N_19321,N_15855,N_18526);
nor U19322 (N_19322,N_15183,N_15346);
or U19323 (N_19323,N_13764,N_12995);
xor U19324 (N_19324,N_17396,N_13583);
nor U19325 (N_19325,N_15163,N_16579);
or U19326 (N_19326,N_13488,N_17451);
nand U19327 (N_19327,N_13172,N_15041);
nand U19328 (N_19328,N_15605,N_13008);
and U19329 (N_19329,N_14584,N_17084);
nand U19330 (N_19330,N_17098,N_17398);
or U19331 (N_19331,N_18156,N_15394);
or U19332 (N_19332,N_18377,N_14466);
nor U19333 (N_19333,N_16248,N_14399);
xor U19334 (N_19334,N_16426,N_13169);
or U19335 (N_19335,N_17769,N_17626);
or U19336 (N_19336,N_14833,N_14510);
and U19337 (N_19337,N_12730,N_14313);
or U19338 (N_19338,N_16434,N_13535);
and U19339 (N_19339,N_16530,N_16998);
or U19340 (N_19340,N_17021,N_15452);
and U19341 (N_19341,N_16317,N_15491);
xor U19342 (N_19342,N_15078,N_14176);
nand U19343 (N_19343,N_17709,N_13812);
nor U19344 (N_19344,N_18136,N_16988);
nand U19345 (N_19345,N_15997,N_17117);
and U19346 (N_19346,N_18685,N_14120);
nand U19347 (N_19347,N_14786,N_14041);
or U19348 (N_19348,N_14532,N_14452);
or U19349 (N_19349,N_17712,N_17521);
or U19350 (N_19350,N_13403,N_17195);
or U19351 (N_19351,N_15219,N_18063);
xor U19352 (N_19352,N_18215,N_17815);
and U19353 (N_19353,N_16463,N_16819);
and U19354 (N_19354,N_16235,N_17835);
and U19355 (N_19355,N_14180,N_15340);
and U19356 (N_19356,N_14706,N_13529);
and U19357 (N_19357,N_16037,N_13956);
or U19358 (N_19358,N_13579,N_17913);
and U19359 (N_19359,N_17178,N_16031);
and U19360 (N_19360,N_17952,N_13765);
and U19361 (N_19361,N_18122,N_13484);
and U19362 (N_19362,N_18719,N_16052);
xor U19363 (N_19363,N_17107,N_18683);
xor U19364 (N_19364,N_17728,N_13887);
and U19365 (N_19365,N_18560,N_13623);
or U19366 (N_19366,N_14660,N_16371);
nor U19367 (N_19367,N_12672,N_13406);
nand U19368 (N_19368,N_14898,N_18103);
nor U19369 (N_19369,N_14156,N_13139);
nor U19370 (N_19370,N_18094,N_14728);
nand U19371 (N_19371,N_12732,N_18362);
and U19372 (N_19372,N_17594,N_18197);
and U19373 (N_19373,N_15709,N_17445);
nand U19374 (N_19374,N_18309,N_16246);
xnor U19375 (N_19375,N_17652,N_18506);
or U19376 (N_19376,N_12764,N_16567);
or U19377 (N_19377,N_14288,N_12663);
and U19378 (N_19378,N_15724,N_17389);
nor U19379 (N_19379,N_18421,N_17049);
and U19380 (N_19380,N_17930,N_17980);
nor U19381 (N_19381,N_15516,N_13556);
and U19382 (N_19382,N_14501,N_17154);
and U19383 (N_19383,N_13288,N_18144);
nand U19384 (N_19384,N_16102,N_16024);
nor U19385 (N_19385,N_15914,N_16559);
nand U19386 (N_19386,N_14396,N_12640);
and U19387 (N_19387,N_18116,N_18603);
xor U19388 (N_19388,N_18032,N_15028);
xnor U19389 (N_19389,N_12933,N_13386);
and U19390 (N_19390,N_17866,N_13497);
or U19391 (N_19391,N_15566,N_15517);
nor U19392 (N_19392,N_18239,N_17153);
or U19393 (N_19393,N_16525,N_17109);
and U19394 (N_19394,N_13512,N_18473);
and U19395 (N_19395,N_12576,N_15254);
nor U19396 (N_19396,N_18107,N_12992);
or U19397 (N_19397,N_14074,N_12999);
and U19398 (N_19398,N_15953,N_15846);
or U19399 (N_19399,N_18495,N_14951);
and U19400 (N_19400,N_14335,N_15018);
nor U19401 (N_19401,N_12857,N_18045);
xnor U19402 (N_19402,N_14167,N_12710);
nand U19403 (N_19403,N_14979,N_13157);
nand U19404 (N_19404,N_15290,N_14181);
nand U19405 (N_19405,N_13644,N_17723);
nor U19406 (N_19406,N_15939,N_13290);
nor U19407 (N_19407,N_13045,N_13275);
nor U19408 (N_19408,N_13842,N_14508);
or U19409 (N_19409,N_16338,N_15258);
nand U19410 (N_19410,N_13980,N_15211);
nand U19411 (N_19411,N_14605,N_13729);
and U19412 (N_19412,N_18453,N_13808);
or U19413 (N_19413,N_15919,N_17808);
nor U19414 (N_19414,N_13044,N_14449);
or U19415 (N_19415,N_18241,N_12510);
and U19416 (N_19416,N_17536,N_15502);
and U19417 (N_19417,N_17895,N_18542);
nand U19418 (N_19418,N_14016,N_17970);
nand U19419 (N_19419,N_14448,N_15880);
nand U19420 (N_19420,N_14489,N_15922);
and U19421 (N_19421,N_13120,N_13499);
nand U19422 (N_19422,N_17748,N_17849);
and U19423 (N_19423,N_17192,N_16120);
nor U19424 (N_19424,N_14921,N_17434);
and U19425 (N_19425,N_18271,N_14758);
nand U19426 (N_19426,N_17110,N_17714);
xnor U19427 (N_19427,N_16751,N_15549);
or U19428 (N_19428,N_13618,N_17295);
and U19429 (N_19429,N_18041,N_16760);
or U19430 (N_19430,N_17474,N_17544);
nor U19431 (N_19431,N_18521,N_16680);
or U19432 (N_19432,N_14640,N_14062);
nand U19433 (N_19433,N_13015,N_16508);
nor U19434 (N_19434,N_12680,N_16588);
or U19435 (N_19435,N_13707,N_14983);
and U19436 (N_19436,N_16684,N_17631);
nand U19437 (N_19437,N_16604,N_17471);
and U19438 (N_19438,N_15438,N_16905);
or U19439 (N_19439,N_14969,N_14845);
nand U19440 (N_19440,N_16601,N_14816);
nor U19441 (N_19441,N_18498,N_13021);
and U19442 (N_19442,N_18482,N_15575);
nor U19443 (N_19443,N_16315,N_12792);
nor U19444 (N_19444,N_12631,N_13539);
nand U19445 (N_19445,N_14885,N_17406);
nand U19446 (N_19446,N_15066,N_16893);
xnor U19447 (N_19447,N_16494,N_17301);
and U19448 (N_19448,N_13962,N_17917);
nor U19449 (N_19449,N_13825,N_17168);
or U19450 (N_19450,N_16626,N_15112);
xor U19451 (N_19451,N_13689,N_18580);
nor U19452 (N_19452,N_16689,N_13438);
or U19453 (N_19453,N_13259,N_16073);
and U19454 (N_19454,N_17108,N_18318);
and U19455 (N_19455,N_17938,N_12528);
or U19456 (N_19456,N_13374,N_12650);
nor U19457 (N_19457,N_14474,N_16883);
nand U19458 (N_19458,N_17250,N_17190);
nand U19459 (N_19459,N_13915,N_14204);
nor U19460 (N_19460,N_13597,N_14442);
nor U19461 (N_19461,N_17121,N_18284);
and U19462 (N_19462,N_15917,N_13522);
nor U19463 (N_19463,N_14504,N_17413);
and U19464 (N_19464,N_18407,N_13511);
and U19465 (N_19465,N_17149,N_13895);
xnor U19466 (N_19466,N_16369,N_18536);
and U19467 (N_19467,N_17710,N_18276);
or U19468 (N_19468,N_16890,N_13216);
and U19469 (N_19469,N_13477,N_15696);
nand U19470 (N_19470,N_18567,N_14649);
or U19471 (N_19471,N_14762,N_15135);
or U19472 (N_19472,N_14114,N_18448);
xor U19473 (N_19473,N_17296,N_17048);
nand U19474 (N_19474,N_15351,N_17550);
and U19475 (N_19475,N_14296,N_16480);
or U19476 (N_19476,N_15191,N_16117);
nand U19477 (N_19477,N_13370,N_16194);
nor U19478 (N_19478,N_15713,N_13629);
and U19479 (N_19479,N_18279,N_13943);
and U19480 (N_19480,N_14974,N_15636);
and U19481 (N_19481,N_16995,N_12984);
nor U19482 (N_19482,N_14558,N_17452);
or U19483 (N_19483,N_17124,N_13665);
or U19484 (N_19484,N_18556,N_13116);
nand U19485 (N_19485,N_13658,N_13035);
or U19486 (N_19486,N_18012,N_15865);
or U19487 (N_19487,N_15567,N_13717);
and U19488 (N_19488,N_16381,N_14919);
or U19489 (N_19489,N_13740,N_17966);
nand U19490 (N_19490,N_14414,N_13442);
nor U19491 (N_19491,N_13221,N_14208);
nor U19492 (N_19492,N_12653,N_17885);
nand U19493 (N_19493,N_17640,N_12585);
nor U19494 (N_19494,N_17638,N_12728);
or U19495 (N_19495,N_17448,N_13067);
and U19496 (N_19496,N_17046,N_15666);
nand U19497 (N_19497,N_17120,N_15030);
nand U19498 (N_19498,N_17717,N_17659);
nor U19499 (N_19499,N_18533,N_14009);
nand U19500 (N_19500,N_14813,N_13719);
nor U19501 (N_19501,N_17601,N_17697);
and U19502 (N_19502,N_13968,N_18445);
or U19503 (N_19503,N_17950,N_12587);
nand U19504 (N_19504,N_13614,N_17792);
or U19505 (N_19505,N_14037,N_13313);
nor U19506 (N_19506,N_13589,N_15193);
or U19507 (N_19507,N_14561,N_12970);
nand U19508 (N_19508,N_18546,N_12820);
nand U19509 (N_19509,N_15279,N_18159);
xnor U19510 (N_19510,N_15157,N_17113);
or U19511 (N_19511,N_15828,N_15519);
and U19512 (N_19512,N_13027,N_18047);
nand U19513 (N_19513,N_17210,N_17330);
nor U19514 (N_19514,N_16044,N_13880);
and U19515 (N_19515,N_15110,N_13732);
nand U19516 (N_19516,N_13855,N_18219);
and U19517 (N_19517,N_12895,N_13068);
and U19518 (N_19518,N_17939,N_18005);
or U19519 (N_19519,N_18464,N_17868);
nand U19520 (N_19520,N_13703,N_18312);
and U19521 (N_19521,N_12767,N_16786);
or U19522 (N_19522,N_14978,N_12636);
xor U19523 (N_19523,N_16557,N_16115);
nand U19524 (N_19524,N_14928,N_18437);
nor U19525 (N_19525,N_15744,N_12924);
or U19526 (N_19526,N_13864,N_14893);
or U19527 (N_19527,N_14385,N_16712);
or U19528 (N_19528,N_18745,N_16017);
or U19529 (N_19529,N_15854,N_14286);
or U19530 (N_19530,N_16664,N_17997);
and U19531 (N_19531,N_13099,N_14543);
nand U19532 (N_19532,N_17456,N_16297);
nor U19533 (N_19533,N_16004,N_17197);
xor U19534 (N_19534,N_17995,N_16693);
nor U19535 (N_19535,N_15272,N_14345);
nor U19536 (N_19536,N_18035,N_16358);
nor U19537 (N_19537,N_14004,N_16771);
nand U19538 (N_19538,N_16041,N_13069);
or U19539 (N_19539,N_16233,N_16539);
nor U19540 (N_19540,N_13433,N_14646);
or U19541 (N_19541,N_16347,N_18499);
and U19542 (N_19542,N_15927,N_15128);
nor U19543 (N_19543,N_14479,N_14237);
or U19544 (N_19544,N_15302,N_14099);
xnor U19545 (N_19545,N_16796,N_17996);
or U19546 (N_19546,N_14620,N_15637);
xor U19547 (N_19547,N_17233,N_16106);
and U19548 (N_19548,N_13854,N_16456);
nor U19549 (N_19549,N_17897,N_14324);
nor U19550 (N_19550,N_15602,N_13363);
and U19551 (N_19551,N_15119,N_18476);
or U19552 (N_19552,N_16204,N_13392);
nand U19553 (N_19553,N_16029,N_16709);
nor U19554 (N_19554,N_14665,N_17762);
xor U19555 (N_19555,N_17831,N_15966);
nor U19556 (N_19556,N_16957,N_17798);
and U19557 (N_19557,N_18275,N_14091);
or U19558 (N_19558,N_15990,N_17757);
or U19559 (N_19559,N_13853,N_13338);
nor U19560 (N_19560,N_13639,N_13449);
and U19561 (N_19561,N_16108,N_18006);
nor U19562 (N_19562,N_18367,N_12790);
nor U19563 (N_19563,N_16306,N_14453);
nand U19564 (N_19564,N_12986,N_13284);
nand U19565 (N_19565,N_14390,N_15861);
or U19566 (N_19566,N_13679,N_16683);
nand U19567 (N_19567,N_13176,N_15702);
or U19568 (N_19568,N_18092,N_13520);
xor U19569 (N_19569,N_16153,N_13038);
nor U19570 (N_19570,N_17587,N_16402);
or U19571 (N_19571,N_16824,N_15546);
xor U19572 (N_19572,N_14991,N_17781);
xor U19573 (N_19573,N_15833,N_16574);
or U19574 (N_19574,N_13528,N_13598);
nor U19575 (N_19575,N_12910,N_14076);
nor U19576 (N_19576,N_14401,N_18264);
nor U19577 (N_19577,N_12588,N_14527);
and U19578 (N_19578,N_13845,N_13517);
nor U19579 (N_19579,N_15231,N_17983);
xor U19580 (N_19580,N_17941,N_15239);
and U19581 (N_19581,N_15039,N_15529);
nand U19582 (N_19582,N_17020,N_14726);
xor U19583 (N_19583,N_16523,N_13394);
nand U19584 (N_19584,N_17014,N_16123);
nor U19585 (N_19585,N_16510,N_13435);
or U19586 (N_19586,N_14599,N_16100);
nand U19587 (N_19587,N_13375,N_13850);
xor U19588 (N_19588,N_18410,N_12659);
nand U19589 (N_19589,N_18588,N_16859);
nor U19590 (N_19590,N_14413,N_15413);
or U19591 (N_19591,N_17255,N_15622);
and U19592 (N_19592,N_18703,N_12954);
nand U19593 (N_19593,N_18738,N_15181);
or U19594 (N_19594,N_18112,N_16019);
xor U19595 (N_19595,N_16275,N_17623);
or U19596 (N_19596,N_16765,N_15149);
or U19597 (N_19597,N_12697,N_12797);
nand U19598 (N_19598,N_12866,N_14606);
and U19599 (N_19599,N_17820,N_14290);
xnor U19600 (N_19600,N_15484,N_14675);
or U19601 (N_19601,N_12745,N_14065);
or U19602 (N_19602,N_18701,N_13148);
and U19603 (N_19603,N_16054,N_13716);
and U19604 (N_19604,N_15430,N_14336);
nand U19605 (N_19605,N_16608,N_13553);
and U19606 (N_19606,N_17194,N_14412);
and U19607 (N_19607,N_15469,N_14779);
nor U19608 (N_19608,N_17699,N_13269);
and U19609 (N_19609,N_15379,N_12641);
xnor U19610 (N_19610,N_14815,N_14537);
or U19611 (N_19611,N_14418,N_15701);
nand U19612 (N_19612,N_18392,N_17378);
and U19613 (N_19613,N_18178,N_13565);
nand U19614 (N_19614,N_14823,N_14500);
nor U19615 (N_19615,N_18186,N_14151);
and U19616 (N_19616,N_13894,N_18427);
or U19617 (N_19617,N_17780,N_17030);
or U19618 (N_19618,N_17535,N_16895);
nor U19619 (N_19619,N_18146,N_18299);
nand U19620 (N_19620,N_15355,N_18474);
xnor U19621 (N_19621,N_13037,N_16969);
or U19622 (N_19622,N_15694,N_13823);
nand U19623 (N_19623,N_17097,N_15213);
xnor U19624 (N_19624,N_18565,N_13735);
nand U19625 (N_19625,N_18634,N_13508);
nand U19626 (N_19626,N_18099,N_15518);
nand U19627 (N_19627,N_13699,N_14366);
nand U19628 (N_19628,N_18381,N_17257);
xor U19629 (N_19629,N_17372,N_16361);
nor U19630 (N_19630,N_14874,N_13888);
and U19631 (N_19631,N_15726,N_13098);
nor U19632 (N_19632,N_15075,N_16378);
or U19633 (N_19633,N_18501,N_14577);
nand U19634 (N_19634,N_18170,N_16845);
or U19635 (N_19635,N_12967,N_15871);
and U19636 (N_19636,N_16164,N_17055);
nand U19637 (N_19637,N_12656,N_14198);
nand U19638 (N_19638,N_16070,N_18038);
nand U19639 (N_19639,N_14015,N_14281);
nor U19640 (N_19640,N_18295,N_18586);
nor U19641 (N_19641,N_17501,N_16748);
nand U19642 (N_19642,N_13547,N_16918);
nor U19643 (N_19643,N_13092,N_15630);
xnor U19644 (N_19644,N_15715,N_13815);
and U19645 (N_19645,N_14177,N_17350);
nor U19646 (N_19646,N_15892,N_13557);
and U19647 (N_19647,N_12561,N_18249);
nand U19648 (N_19648,N_18505,N_16687);
nand U19649 (N_19649,N_13897,N_15857);
nor U19650 (N_19650,N_13848,N_15403);
or U19651 (N_19651,N_14657,N_15781);
nor U19652 (N_19652,N_16673,N_15968);
nor U19653 (N_19653,N_13749,N_15065);
and U19654 (N_19654,N_13253,N_16169);
nand U19655 (N_19655,N_18232,N_16332);
and U19656 (N_19656,N_14072,N_15673);
nand U19657 (N_19657,N_18484,N_18278);
and U19658 (N_19658,N_13198,N_13705);
and U19659 (N_19659,N_13168,N_13627);
and U19660 (N_19660,N_13992,N_16753);
and U19661 (N_19661,N_16534,N_14249);
or U19662 (N_19662,N_14690,N_18672);
nand U19663 (N_19663,N_14554,N_14438);
and U19664 (N_19664,N_16405,N_14187);
nor U19665 (N_19665,N_14005,N_15898);
nand U19666 (N_19666,N_13398,N_16837);
or U19667 (N_19667,N_18625,N_14228);
or U19668 (N_19668,N_14536,N_13108);
and U19669 (N_19669,N_15536,N_15627);
xnor U19670 (N_19670,N_15286,N_15425);
xnor U19671 (N_19671,N_17852,N_13400);
and U19672 (N_19672,N_13354,N_13206);
or U19673 (N_19673,N_16955,N_17873);
and U19674 (N_19674,N_15244,N_15980);
xnor U19675 (N_19675,N_16143,N_14852);
nand U19676 (N_19676,N_12542,N_12749);
nor U19677 (N_19677,N_15293,N_13919);
or U19678 (N_19678,N_14188,N_13241);
or U19679 (N_19679,N_16850,N_14171);
and U19680 (N_19680,N_16002,N_14721);
and U19681 (N_19681,N_16458,N_16799);
nand U19682 (N_19682,N_17608,N_17460);
and U19683 (N_19683,N_14209,N_16443);
and U19684 (N_19684,N_16790,N_16096);
or U19685 (N_19685,N_13857,N_15247);
xnor U19686 (N_19686,N_12733,N_18500);
nand U19687 (N_19687,N_13457,N_14687);
and U19688 (N_19688,N_13397,N_16766);
or U19689 (N_19689,N_17245,N_16869);
nor U19690 (N_19690,N_13308,N_13564);
nor U19691 (N_19691,N_16393,N_14429);
nor U19692 (N_19692,N_16293,N_18185);
or U19693 (N_19693,N_15670,N_13966);
nand U19694 (N_19694,N_13661,N_16522);
nand U19695 (N_19695,N_14498,N_18532);
or U19696 (N_19696,N_12788,N_18298);
nand U19697 (N_19697,N_12759,N_15192);
and U19698 (N_19698,N_12748,N_14496);
nor U19699 (N_19699,N_14276,N_12875);
nor U19700 (N_19700,N_12781,N_16284);
nand U19701 (N_19701,N_13518,N_14403);
nor U19702 (N_19702,N_12593,N_13509);
xor U19703 (N_19703,N_18181,N_12698);
and U19704 (N_19704,N_15767,N_12872);
nor U19705 (N_19705,N_16326,N_12823);
nand U19706 (N_19706,N_17209,N_14513);
nor U19707 (N_19707,N_15937,N_17826);
or U19708 (N_19708,N_16517,N_14594);
or U19709 (N_19709,N_14000,N_15737);
nor U19710 (N_19710,N_12644,N_13391);
nand U19711 (N_19711,N_18478,N_16414);
xor U19712 (N_19712,N_12613,N_16475);
nand U19713 (N_19713,N_14021,N_14785);
nand U19714 (N_19714,N_15935,N_18166);
or U19715 (N_19715,N_18590,N_17432);
or U19716 (N_19716,N_14849,N_16622);
xnor U19717 (N_19717,N_18631,N_14958);
nor U19718 (N_19718,N_18301,N_15563);
nor U19719 (N_19719,N_14511,N_14461);
and U19720 (N_19720,N_18343,N_16831);
or U19721 (N_19721,N_13817,N_17731);
or U19722 (N_19722,N_18329,N_14772);
nand U19723 (N_19723,N_16300,N_15851);
or U19724 (N_19724,N_14468,N_17720);
nor U19725 (N_19725,N_13777,N_14473);
and U19726 (N_19726,N_13647,N_13422);
nand U19727 (N_19727,N_15834,N_16773);
and U19728 (N_19728,N_13207,N_15537);
or U19729 (N_19729,N_17912,N_13914);
nor U19730 (N_19730,N_12908,N_15230);
nor U19731 (N_19731,N_16056,N_14008);
and U19732 (N_19732,N_14265,N_14955);
nand U19733 (N_19733,N_16231,N_17261);
and U19734 (N_19734,N_14672,N_18363);
nand U19735 (N_19735,N_16200,N_13878);
and U19736 (N_19736,N_14213,N_17112);
or U19737 (N_19737,N_17526,N_17541);
or U19738 (N_19738,N_15316,N_13049);
nand U19739 (N_19739,N_18059,N_13828);
or U19740 (N_19740,N_17453,N_16177);
or U19741 (N_19741,N_18561,N_16583);
or U19742 (N_19742,N_17854,N_15878);
and U19743 (N_19743,N_18548,N_13322);
or U19744 (N_19744,N_14712,N_15453);
and U19745 (N_19745,N_16423,N_17482);
nor U19746 (N_19746,N_13834,N_14038);
or U19747 (N_19747,N_18293,N_16504);
nor U19748 (N_19748,N_18573,N_17902);
and U19749 (N_19749,N_16965,N_13833);
and U19750 (N_19750,N_13441,N_17607);
nor U19751 (N_19751,N_15383,N_12533);
xor U19752 (N_19752,N_16900,N_13584);
nor U19753 (N_19753,N_14718,N_17749);
nor U19754 (N_19754,N_13981,N_13134);
nand U19755 (N_19755,N_18508,N_17718);
and U19756 (N_19756,N_14784,N_14743);
nand U19757 (N_19757,N_13434,N_17430);
nand U19758 (N_19758,N_14347,N_12848);
or U19759 (N_19759,N_13908,N_16012);
nand U19760 (N_19760,N_16675,N_12679);
and U19761 (N_19761,N_18147,N_12839);
nor U19762 (N_19762,N_13028,N_14860);
nand U19763 (N_19763,N_17555,N_12916);
xnor U19764 (N_19764,N_18578,N_14565);
nand U19765 (N_19765,N_14042,N_15093);
and U19766 (N_19766,N_16930,N_12966);
xnor U19767 (N_19767,N_18016,N_17211);
and U19768 (N_19768,N_17656,N_18037);
xnor U19769 (N_19769,N_17667,N_14087);
nor U19770 (N_19770,N_13625,N_15626);
or U19771 (N_19771,N_16461,N_17766);
and U19772 (N_19772,N_13772,N_12961);
nand U19773 (N_19773,N_18512,N_16262);
nand U19774 (N_19774,N_15409,N_15134);
and U19775 (N_19775,N_17226,N_15269);
nor U19776 (N_19776,N_13184,N_18017);
nand U19777 (N_19777,N_16446,N_16195);
and U19778 (N_19778,N_14647,N_18626);
xnor U19779 (N_19779,N_15329,N_17228);
xnor U19780 (N_19780,N_13955,N_14057);
nor U19781 (N_19781,N_15692,N_15838);
xor U19782 (N_19782,N_15826,N_17306);
or U19783 (N_19783,N_17002,N_12655);
nor U19784 (N_19784,N_16098,N_13360);
or U19785 (N_19785,N_13819,N_15741);
or U19786 (N_19786,N_12562,N_16362);
nand U19787 (N_19787,N_18621,N_17893);
nand U19788 (N_19788,N_14045,N_15590);
or U19789 (N_19789,N_15649,N_18277);
and U19790 (N_19790,N_15339,N_17915);
nand U19791 (N_19791,N_12852,N_13445);
nand U19792 (N_19792,N_17099,N_15478);
xor U19793 (N_19793,N_12602,N_18200);
or U19794 (N_19794,N_13408,N_15248);
and U19795 (N_19795,N_14623,N_16206);
nor U19796 (N_19796,N_12935,N_18326);
xor U19797 (N_19797,N_15380,N_13608);
or U19798 (N_19798,N_13708,N_18150);
and U19799 (N_19799,N_17716,N_13882);
nor U19800 (N_19800,N_18522,N_15841);
nand U19801 (N_19801,N_13587,N_14210);
nand U19802 (N_19802,N_13250,N_14946);
and U19803 (N_19803,N_13766,N_15944);
nand U19804 (N_19804,N_15327,N_14651);
and U19805 (N_19805,N_13810,N_15708);
or U19806 (N_19806,N_15951,N_16101);
nor U19807 (N_19807,N_15322,N_16253);
nand U19808 (N_19808,N_16724,N_13591);
xor U19809 (N_19809,N_14952,N_14841);
xnor U19810 (N_19810,N_16909,N_15208);
nor U19811 (N_19811,N_15683,N_14051);
nand U19812 (N_19812,N_13568,N_16224);
and U19813 (N_19813,N_18608,N_13849);
and U19814 (N_19814,N_14010,N_15111);
nor U19815 (N_19815,N_18400,N_13417);
nor U19816 (N_19816,N_14988,N_15268);
and U19817 (N_19817,N_17625,N_17679);
nor U19818 (N_19818,N_14780,N_15648);
nor U19819 (N_19819,N_13967,N_15342);
and U19820 (N_19820,N_14575,N_12548);
nor U19821 (N_19821,N_17824,N_16503);
and U19822 (N_19822,N_17908,N_17345);
nand U19823 (N_19823,N_14676,N_17057);
or U19824 (N_19824,N_15459,N_18134);
nor U19825 (N_19825,N_12815,N_18270);
or U19826 (N_19826,N_13405,N_13229);
nor U19827 (N_19827,N_13452,N_17621);
or U19828 (N_19828,N_14538,N_14193);
nor U19829 (N_19829,N_18637,N_17087);
nor U19830 (N_19830,N_15848,N_13197);
nor U19831 (N_19831,N_14821,N_18419);
nor U19832 (N_19832,N_14007,N_17604);
nor U19833 (N_19833,N_17335,N_17752);
nand U19834 (N_19834,N_13592,N_16442);
xnor U19835 (N_19835,N_18629,N_15420);
xnor U19836 (N_19836,N_17176,N_17050);
xnor U19837 (N_19837,N_17517,N_17105);
nand U19838 (N_19838,N_16285,N_13033);
and U19839 (N_19839,N_15261,N_18082);
and U19840 (N_19840,N_14022,N_14243);
or U19841 (N_19841,N_13271,N_18022);
nor U19842 (N_19842,N_14297,N_13023);
nand U19843 (N_19843,N_17085,N_12743);
nor U19844 (N_19844,N_18297,N_14559);
nand U19845 (N_19845,N_17646,N_13230);
nor U19846 (N_19846,N_12883,N_14674);
and U19847 (N_19847,N_13482,N_12591);
nand U19848 (N_19848,N_17800,N_16090);
or U19849 (N_19849,N_12755,N_17232);
nor U19850 (N_19850,N_17674,N_13464);
or U19851 (N_19851,N_13816,N_14360);
xor U19852 (N_19852,N_16934,N_18167);
and U19853 (N_19853,N_13451,N_14497);
or U19854 (N_19854,N_12506,N_16057);
nand U19855 (N_19855,N_16010,N_13151);
or U19856 (N_19856,N_15287,N_18722);
nand U19857 (N_19857,N_14637,N_16547);
nand U19858 (N_19858,N_13381,N_18350);
or U19859 (N_19859,N_16556,N_17361);
nor U19860 (N_19860,N_14886,N_16319);
nand U19861 (N_19861,N_15813,N_16835);
nor U19862 (N_19862,N_18463,N_15314);
nor U19863 (N_19863,N_12677,N_13448);
nand U19864 (N_19864,N_13525,N_15056);
nor U19865 (N_19865,N_16644,N_18231);
xnor U19866 (N_19866,N_16966,N_16470);
nand U19867 (N_19867,N_14084,N_15147);
xnor U19868 (N_19868,N_18332,N_13390);
nor U19869 (N_19869,N_15651,N_15882);
and U19870 (N_19870,N_15789,N_15818);
nor U19871 (N_19871,N_15062,N_13542);
nand U19872 (N_19872,N_18255,N_13787);
nand U19873 (N_19873,N_18196,N_14622);
or U19874 (N_19874,N_16817,N_18148);
nor U19875 (N_19875,N_14285,N_13744);
or U19876 (N_19876,N_12639,N_16563);
or U19877 (N_19877,N_18543,N_15038);
nand U19878 (N_19878,N_16743,N_15331);
nor U19879 (N_19879,N_17419,N_15601);
nand U19880 (N_19880,N_16650,N_18191);
nor U19881 (N_19881,N_17401,N_14636);
xor U19882 (N_19882,N_13973,N_17003);
nand U19883 (N_19883,N_18641,N_17311);
nor U19884 (N_19884,N_13419,N_18327);
nor U19885 (N_19885,N_15612,N_13265);
xnor U19886 (N_19886,N_15685,N_18581);
nor U19887 (N_19887,N_16694,N_18226);
nand U19888 (N_19888,N_14251,N_16497);
nand U19889 (N_19889,N_16392,N_17188);
nand U19890 (N_19890,N_15620,N_15447);
and U19891 (N_19891,N_16952,N_16784);
and U19892 (N_19892,N_17137,N_16939);
nand U19893 (N_19893,N_17732,N_16882);
and U19894 (N_19894,N_12763,N_12531);
or U19895 (N_19895,N_16499,N_13491);
or U19896 (N_19896,N_12556,N_12583);
nand U19897 (N_19897,N_16621,N_12521);
or U19898 (N_19898,N_17400,N_16959);
nand U19899 (N_19899,N_12747,N_14039);
or U19900 (N_19900,N_18458,N_16124);
and U19901 (N_19901,N_13570,N_15596);
and U19902 (N_19902,N_13870,N_15830);
xnor U19903 (N_19903,N_16860,N_15434);
xor U19904 (N_19904,N_16088,N_18454);
or U19905 (N_19905,N_14572,N_15631);
nand U19906 (N_19906,N_16185,N_14614);
and U19907 (N_19907,N_17617,N_18015);
or U19908 (N_19908,N_14535,N_13273);
nand U19909 (N_19909,N_16139,N_17724);
and U19910 (N_19910,N_16578,N_13208);
and U19911 (N_19911,N_14269,N_16540);
or U19912 (N_19912,N_15783,N_16598);
nor U19913 (N_19913,N_12926,N_15001);
or U19914 (N_19914,N_14905,N_17365);
nor U19915 (N_19915,N_16211,N_17676);
nand U19916 (N_19916,N_18408,N_17323);
nor U19917 (N_19917,N_15399,N_16252);
nor U19918 (N_19918,N_16043,N_16339);
nand U19919 (N_19919,N_15625,N_18061);
or U19920 (N_19920,N_18180,N_18235);
nor U19921 (N_19921,N_13650,N_14752);
and U19922 (N_19922,N_18539,N_13913);
and U19923 (N_19923,N_15984,N_14685);
and U19924 (N_19924,N_15063,N_14879);
nor U19925 (N_19925,N_14902,N_14001);
nor U19926 (N_19926,N_17267,N_12793);
nor U19927 (N_19927,N_18223,N_17102);
nand U19928 (N_19928,N_18280,N_16571);
or U19929 (N_19929,N_14098,N_17967);
and U19930 (N_19930,N_16677,N_13291);
or U19931 (N_19931,N_15808,N_12611);
nand U19932 (N_19932,N_14737,N_15921);
nor U19933 (N_19933,N_13101,N_14205);
xnor U19934 (N_19934,N_18360,N_14053);
and U19935 (N_19935,N_18416,N_13778);
nand U19936 (N_19936,N_15797,N_17258);
nand U19937 (N_19937,N_18555,N_14416);
and U19938 (N_19938,N_17315,N_15308);
or U19939 (N_19939,N_14929,N_16509);
or U19940 (N_19940,N_16597,N_16015);
or U19941 (N_19941,N_18024,N_13263);
and U19942 (N_19942,N_16314,N_17028);
nor U19943 (N_19943,N_13883,N_14274);
or U19944 (N_19944,N_15270,N_12785);
and U19945 (N_19945,N_12526,N_13383);
nand U19946 (N_19946,N_15793,N_17616);
nand U19947 (N_19947,N_16920,N_16178);
or U19948 (N_19948,N_18294,N_17999);
and U19949 (N_19949,N_16097,N_13599);
nand U19950 (N_19950,N_17793,N_13124);
or U19951 (N_19951,N_15080,N_15166);
or U19952 (N_19952,N_17447,N_13963);
nand U19953 (N_19953,N_14226,N_18553);
nor U19954 (N_19954,N_18736,N_15780);
or U19955 (N_19955,N_13060,N_13412);
and U19956 (N_19956,N_17270,N_18316);
and U19957 (N_19957,N_16891,N_13153);
and U19958 (N_19958,N_14673,N_16005);
nand U19959 (N_19959,N_16569,N_13601);
nand U19960 (N_19960,N_16528,N_15171);
nand U19961 (N_19961,N_15186,N_14095);
nand U19962 (N_19962,N_13753,N_17737);
nand U19963 (N_19963,N_17461,N_17441);
and U19964 (N_19964,N_15893,N_17689);
nand U19965 (N_19965,N_15659,N_15205);
nor U19966 (N_19966,N_15665,N_13685);
or U19967 (N_19967,N_18372,N_17986);
nand U19968 (N_19968,N_15844,N_13194);
or U19969 (N_19969,N_15104,N_13200);
nor U19970 (N_19970,N_14428,N_17370);
and U19971 (N_19971,N_15671,N_15321);
xnor U19972 (N_19972,N_13025,N_15853);
nand U19973 (N_19973,N_13588,N_17770);
or U19974 (N_19974,N_14825,N_14738);
or U19975 (N_19975,N_15899,N_12965);
and U19976 (N_19976,N_18492,N_18447);
and U19977 (N_19977,N_17309,N_13296);
nand U19978 (N_19978,N_18336,N_18030);
or U19979 (N_19979,N_18622,N_15046);
nand U19980 (N_19980,N_17022,N_14318);
nand U19981 (N_19981,N_17147,N_18202);
or U19982 (N_19982,N_13657,N_13911);
nand U19983 (N_19983,N_13526,N_15291);
nand U19984 (N_19984,N_14552,N_18649);
or U19985 (N_19985,N_13285,N_16535);
or U19986 (N_19986,N_13311,N_15169);
and U19987 (N_19987,N_16723,N_16184);
or U19988 (N_19988,N_15555,N_17546);
and U19989 (N_19989,N_14368,N_16219);
and U19990 (N_19990,N_18211,N_14397);
nor U19991 (N_19991,N_15426,N_14305);
xor U19992 (N_19992,N_12579,N_13059);
or U19993 (N_19993,N_18296,N_14734);
and U19994 (N_19994,N_15792,N_15168);
nor U19995 (N_19995,N_14888,N_15494);
or U19996 (N_19996,N_16828,N_14889);
nor U19997 (N_19997,N_18228,N_17135);
and U19998 (N_19998,N_13569,N_13323);
and U19999 (N_19999,N_14580,N_15406);
or U20000 (N_20000,N_13002,N_12773);
nand U20001 (N_20001,N_16810,N_14716);
or U20002 (N_20002,N_14088,N_17498);
nand U20003 (N_20003,N_15512,N_13796);
nand U20004 (N_20004,N_15955,N_16034);
xnor U20005 (N_20005,N_18593,N_16672);
or U20006 (N_20006,N_17982,N_17740);
or U20007 (N_20007,N_14643,N_18283);
nor U20008 (N_20008,N_18406,N_16927);
nor U20009 (N_20009,N_12838,N_14341);
or U20010 (N_20010,N_16915,N_12892);
and U20011 (N_20011,N_14006,N_14155);
and U20012 (N_20012,N_17841,N_15101);
nor U20013 (N_20013,N_15768,N_14069);
xor U20014 (N_20014,N_14924,N_15175);
nor U20015 (N_20015,N_15305,N_16411);
nor U20016 (N_20016,N_18286,N_12982);
or U20017 (N_20017,N_13741,N_13541);
and U20018 (N_20018,N_16617,N_15733);
nor U20019 (N_20019,N_13190,N_12570);
nand U20020 (N_20020,N_17324,N_18088);
nor U20021 (N_20021,N_13580,N_13861);
nor U20022 (N_20022,N_17353,N_17462);
nand U20023 (N_20023,N_16298,N_18728);
or U20024 (N_20024,N_14838,N_14049);
or U20025 (N_20025,N_13974,N_18469);
nand U20026 (N_20026,N_18709,N_14950);
or U20027 (N_20027,N_14788,N_16663);
or U20028 (N_20028,N_12532,N_12610);
or U20029 (N_20029,N_17379,N_13366);
nand U20030 (N_20030,N_17971,N_17981);
nand U20031 (N_20031,N_14895,N_14847);
or U20032 (N_20032,N_15378,N_16328);
or U20033 (N_20033,N_17540,N_14873);
and U20034 (N_20034,N_18545,N_16159);
xnor U20035 (N_20035,N_16822,N_14034);
nor U20036 (N_20036,N_13111,N_16099);
xor U20037 (N_20037,N_13563,N_12783);
or U20038 (N_20038,N_14967,N_13389);
or U20039 (N_20039,N_13264,N_13333);
nand U20040 (N_20040,N_12626,N_16066);
or U20041 (N_20041,N_12618,N_14724);
and U20042 (N_20042,N_13113,N_17722);
nand U20043 (N_20043,N_17483,N_13999);
and U20044 (N_20044,N_17768,N_16437);
and U20045 (N_20045,N_17101,N_12509);
nand U20046 (N_20046,N_17489,N_15497);
and U20047 (N_20047,N_15486,N_18100);
nor U20048 (N_20048,N_14136,N_16288);
or U20049 (N_20049,N_15417,N_15788);
xor U20050 (N_20050,N_16033,N_17875);
xnor U20051 (N_20051,N_15764,N_17384);
nand U20052 (N_20052,N_12942,N_17402);
and U20053 (N_20053,N_14740,N_13586);
and U20054 (N_20054,N_18206,N_18348);
xor U20055 (N_20055,N_12628,N_18382);
nand U20056 (N_20056,N_17834,N_13469);
nor U20057 (N_20057,N_18540,N_12512);
nand U20058 (N_20058,N_15852,N_13677);
and U20059 (N_20059,N_16247,N_13170);
nor U20060 (N_20060,N_14066,N_13923);
or U20061 (N_20061,N_17516,N_17839);
or U20062 (N_20062,N_16916,N_18676);
nand U20063 (N_20063,N_12601,N_17157);
xnor U20064 (N_20064,N_14161,N_13447);
and U20065 (N_20065,N_13567,N_14525);
nand U20066 (N_20066,N_13048,N_15454);
nand U20067 (N_20067,N_15565,N_15227);
and U20068 (N_20068,N_13093,N_16580);
and U20069 (N_20069,N_18319,N_14891);
or U20070 (N_20070,N_12825,N_13903);
or U20071 (N_20071,N_14689,N_17265);
nor U20072 (N_20072,N_16649,N_16438);
and U20073 (N_20073,N_12981,N_17859);
and U20074 (N_20074,N_13320,N_12858);
or U20075 (N_20075,N_16795,N_12791);
and U20076 (N_20076,N_12503,N_18224);
and U20077 (N_20077,N_12813,N_17666);
nand U20078 (N_20078,N_18328,N_18325);
or U20079 (N_20079,N_15185,N_14970);
and U20080 (N_20080,N_12822,N_15952);
or U20081 (N_20081,N_13283,N_15901);
nand U20082 (N_20082,N_12859,N_15446);
or U20083 (N_20083,N_13867,N_13977);
xor U20084 (N_20084,N_17559,N_18066);
xor U20085 (N_20085,N_13585,N_14063);
nor U20086 (N_20086,N_12865,N_14930);
nor U20087 (N_20087,N_13465,N_12989);
and U20088 (N_20088,N_16370,N_13299);
and U20089 (N_20089,N_17877,N_15124);
nand U20090 (N_20090,N_17314,N_17567);
nor U20091 (N_20091,N_18177,N_16230);
nor U20092 (N_20092,N_15911,N_13022);
nor U20093 (N_20093,N_13219,N_13367);
and U20094 (N_20094,N_12845,N_14715);
nor U20095 (N_20095,N_16708,N_16801);
nand U20096 (N_20096,N_13007,N_13671);
or U20097 (N_20097,N_16452,N_18525);
and U20098 (N_20098,N_18344,N_17012);
or U20099 (N_20099,N_15013,N_13728);
nor U20100 (N_20100,N_16234,N_13791);
or U20101 (N_20101,N_18090,N_16754);
or U20102 (N_20102,N_17148,N_16949);
nor U20103 (N_20103,N_18036,N_12913);
or U20104 (N_20104,N_17420,N_18693);
nand U20105 (N_20105,N_17143,N_14581);
and U20106 (N_20106,N_16450,N_14938);
nand U20107 (N_20107,N_18050,N_17156);
nor U20108 (N_20108,N_14769,N_14529);
nor U20109 (N_20109,N_17001,N_16167);
and U20110 (N_20110,N_18661,N_12726);
xnor U20111 (N_20111,N_16345,N_14310);
nand U20112 (N_20112,N_12607,N_17364);
and U20113 (N_20113,N_13502,N_13548);
nand U20114 (N_20114,N_18544,N_12665);
or U20115 (N_20115,N_17023,N_15918);
nand U20116 (N_20116,N_13407,N_17919);
nor U20117 (N_20117,N_13122,N_16407);
and U20118 (N_20118,N_16421,N_13232);
nand U20119 (N_20119,N_16280,N_15926);
or U20120 (N_20120,N_13361,N_13203);
or U20121 (N_20121,N_16603,N_17944);
nand U20122 (N_20122,N_16028,N_13527);
nand U20123 (N_20123,N_18218,N_14395);
nand U20124 (N_20124,N_16711,N_14199);
or U20125 (N_20125,N_18101,N_16478);
nand U20126 (N_20126,N_14230,N_17888);
nor U20127 (N_20127,N_18075,N_18707);
nor U20128 (N_20128,N_17704,N_18694);
nor U20129 (N_20129,N_13453,N_15161);
or U20130 (N_20130,N_14602,N_17071);
nor U20131 (N_20131,N_17653,N_13739);
and U20132 (N_20132,N_13298,N_13034);
nor U20133 (N_20133,N_18431,N_17251);
xor U20134 (N_20134,N_18429,N_14782);
nand U20135 (N_20135,N_12519,N_12919);
and U20136 (N_20136,N_14325,N_15815);
nor U20137 (N_20137,N_17622,N_16876);
nor U20138 (N_20138,N_14652,N_13056);
nand U20139 (N_20139,N_13490,N_14369);
xnor U20140 (N_20140,N_18503,N_18409);
and U20141 (N_20141,N_14356,N_17677);
or U20142 (N_20142,N_17053,N_13179);
nor U20143 (N_20143,N_16910,N_15115);
xnor U20144 (N_20144,N_15482,N_17248);
nor U20145 (N_20145,N_14800,N_15752);
and U20146 (N_20146,N_14078,N_17693);
and U20147 (N_20147,N_16926,N_16216);
nand U20148 (N_20148,N_18394,N_14828);
xor U20149 (N_20149,N_14292,N_16380);
and U20150 (N_20150,N_15977,N_12604);
or U20151 (N_20151,N_14502,N_14306);
and U20152 (N_20152,N_16793,N_17884);
xnor U20153 (N_20153,N_15278,N_16738);
or U20154 (N_20154,N_18616,N_17510);
or U20155 (N_20155,N_14282,N_17891);
nand U20156 (N_20156,N_18510,N_13380);
and U20157 (N_20157,N_18220,N_17207);
or U20158 (N_20158,N_15203,N_17933);
nand U20159 (N_20159,N_17514,N_12648);
or U20160 (N_20160,N_16922,N_14834);
nand U20161 (N_20161,N_16527,N_13248);
and U20162 (N_20162,N_15458,N_13218);
or U20163 (N_20163,N_13138,N_18584);
nor U20164 (N_20164,N_16335,N_15326);
nand U20165 (N_20165,N_14876,N_13561);
or U20166 (N_20166,N_16396,N_14942);
nor U20167 (N_20167,N_14653,N_17979);
and U20168 (N_20168,N_12756,N_17804);
nand U20169 (N_20169,N_18128,N_13336);
xor U20170 (N_20170,N_15883,N_18665);
nor U20171 (N_20171,N_16624,N_15449);
and U20172 (N_20172,N_16634,N_16615);
or U20173 (N_20173,N_14840,N_13395);
nand U20174 (N_20174,N_14241,N_13620);
and U20175 (N_20175,N_18585,N_13146);
nor U20176 (N_20176,N_16619,N_14790);
nor U20177 (N_20177,N_15432,N_13874);
nor U20178 (N_20178,N_16838,N_15515);
nand U20179 (N_20179,N_16543,N_17706);
or U20180 (N_20180,N_13610,N_16512);
nor U20181 (N_20181,N_15754,N_17183);
nor U20182 (N_20182,N_18331,N_16000);
and U20183 (N_20183,N_17796,N_13847);
nand U20184 (N_20184,N_13692,N_15337);
nand U20185 (N_20185,N_14571,N_16887);
nor U20186 (N_20186,N_14358,N_13387);
or U20187 (N_20187,N_16403,N_15973);
nor U20188 (N_20188,N_15439,N_14719);
and U20189 (N_20189,N_13009,N_12522);
or U20190 (N_20190,N_14080,N_12778);
xor U20191 (N_20191,N_18079,N_13413);
nand U20192 (N_20192,N_17664,N_17145);
nand U20193 (N_20193,N_14456,N_14222);
and U20194 (N_20194,N_17126,N_13802);
nor U20195 (N_20195,N_12589,N_14402);
nor U20196 (N_20196,N_14113,N_17056);
nor U20197 (N_20197,N_13474,N_13928);
xnor U20198 (N_20198,N_12719,N_14455);
xnor U20199 (N_20199,N_13899,N_16747);
or U20200 (N_20200,N_14794,N_13070);
xnor U20201 (N_20201,N_17045,N_15624);
or U20202 (N_20202,N_15999,N_18346);
and U20203 (N_20203,N_15551,N_17585);
xor U20204 (N_20204,N_16260,N_16722);
and U20205 (N_20205,N_13104,N_17079);
and U20206 (N_20206,N_15109,N_15391);
or U20207 (N_20207,N_16800,N_16506);
nand U20208 (N_20208,N_18069,N_16271);
nor U20209 (N_20209,N_14601,N_17244);
xnor U20210 (N_20210,N_17794,N_14299);
nand U20211 (N_20211,N_14681,N_17644);
xor U20212 (N_20212,N_14321,N_17586);
nor U20213 (N_20213,N_18018,N_13902);
nor U20214 (N_20214,N_16217,N_18375);
nand U20215 (N_20215,N_16149,N_13978);
and U20216 (N_20216,N_17016,N_17850);
nor U20217 (N_20217,N_17662,N_15307);
or U20218 (N_20218,N_17475,N_16963);
and U20219 (N_20219,N_16045,N_17673);
or U20220 (N_20220,N_17789,N_12901);
nand U20221 (N_20221,N_15642,N_15050);
nand U20222 (N_20222,N_16076,N_17216);
or U20223 (N_20223,N_17836,N_16422);
and U20224 (N_20224,N_15949,N_14933);
or U20225 (N_20225,N_17730,N_18105);
nor U20226 (N_20226,N_17078,N_16733);
xor U20227 (N_20227,N_17230,N_16605);
xor U20228 (N_20228,N_14165,N_15987);
or U20229 (N_20229,N_15387,N_12800);
nand U20230 (N_20230,N_15948,N_15067);
or U20231 (N_20231,N_17303,N_17132);
nor U20232 (N_20232,N_16448,N_16229);
and U20233 (N_20233,N_14729,N_17262);
and U20234 (N_20234,N_15121,N_18699);
nor U20235 (N_20235,N_17347,N_17494);
or U20236 (N_20236,N_14267,N_18612);
nor U20237 (N_20237,N_16889,N_14014);
and U20238 (N_20238,N_14633,N_16652);
nor U20239 (N_20239,N_14378,N_13004);
xor U20240 (N_20240,N_15521,N_17739);
nor U20241 (N_20241,N_15315,N_18723);
or U20242 (N_20242,N_16829,N_14315);
or U20243 (N_20243,N_12840,N_14430);
and U20244 (N_20244,N_15660,N_17163);
nor U20245 (N_20245,N_18117,N_17492);
xnor U20246 (N_20246,N_18638,N_14612);
and U20247 (N_20247,N_15421,N_17322);
and U20248 (N_20248,N_16212,N_13688);
nor U20249 (N_20249,N_16741,N_12689);
xor U20250 (N_20250,N_16068,N_16454);
xor U20251 (N_20251,N_14162,N_16447);
xnor U20252 (N_20252,N_18598,N_14835);
xor U20253 (N_20253,N_12979,N_17465);
nand U20254 (N_20254,N_12551,N_12880);
and U20255 (N_20255,N_15441,N_17507);
nand U20256 (N_20256,N_16259,N_16081);
nor U20257 (N_20257,N_18617,N_15604);
nor U20258 (N_20258,N_14134,N_12598);
and U20259 (N_20259,N_15234,N_13696);
nor U20260 (N_20260,N_15232,N_18193);
nor U20261 (N_20261,N_14055,N_14189);
xor U20262 (N_20262,N_17700,N_17266);
nor U20263 (N_20263,N_16502,N_12670);
nand U20264 (N_20264,N_16006,N_16440);
nand U20265 (N_20265,N_14383,N_16144);
or U20266 (N_20266,N_14117,N_13959);
and U20267 (N_20267,N_13325,N_13244);
and U20268 (N_20268,N_17754,N_17745);
and U20269 (N_20269,N_14943,N_18031);
or U20270 (N_20270,N_13358,N_15004);
or U20271 (N_20271,N_13513,N_15773);
or U20272 (N_20272,N_17237,N_15574);
and U20273 (N_20273,N_14569,N_13401);
or U20274 (N_20274,N_15839,N_12713);
xor U20275 (N_20275,N_13332,N_17863);
and U20276 (N_20276,N_17407,N_16385);
nor U20277 (N_20277,N_16716,N_13161);
or U20278 (N_20278,N_18052,N_16809);
nor U20279 (N_20279,N_16126,N_15020);
nor U20280 (N_20280,N_14107,N_12617);
or U20281 (N_20281,N_14257,N_17862);
nand U20282 (N_20282,N_17786,N_14192);
nand U20283 (N_20283,N_15774,N_15444);
and U20284 (N_20284,N_12516,N_13885);
nand U20285 (N_20285,N_16135,N_18208);
or U20286 (N_20286,N_15389,N_16886);
or U20287 (N_20287,N_18700,N_16048);
and U20288 (N_20288,N_15757,N_18531);
or U20289 (N_20289,N_17343,N_14073);
or U20290 (N_20290,N_12922,N_18425);
nand U20291 (N_20291,N_13026,N_12896);
nor U20292 (N_20292,N_15156,N_14668);
xor U20293 (N_20293,N_17349,N_18708);
and U20294 (N_20294,N_13775,N_18737);
nor U20295 (N_20295,N_16240,N_17198);
xor U20296 (N_20296,N_16104,N_14806);
nor U20297 (N_20297,N_15584,N_16688);
nand U20298 (N_20298,N_16354,N_17152);
nand U20299 (N_20299,N_13785,N_18322);
nor U20300 (N_20300,N_15628,N_13256);
nand U20301 (N_20301,N_15257,N_13018);
or U20302 (N_20302,N_15958,N_17217);
or U20303 (N_20303,N_17628,N_18570);
or U20304 (N_20304,N_17871,N_18256);
nor U20305 (N_20305,N_17725,N_14644);
xor U20306 (N_20306,N_15688,N_17703);
and U20307 (N_20307,N_14854,N_15437);
and U20308 (N_20308,N_12552,N_17166);
xor U20309 (N_20309,N_14327,N_17713);
or U20310 (N_20310,N_13770,N_12744);
nor U20311 (N_20311,N_18233,N_16546);
xnor U20312 (N_20312,N_14361,N_15368);
nor U20313 (N_20313,N_17123,N_14795);
nand U20314 (N_20314,N_13307,N_17661);
nor U20315 (N_20315,N_14682,N_14720);
or U20316 (N_20316,N_13794,N_14478);
xnor U20317 (N_20317,N_17695,N_16849);
and U20318 (N_20318,N_17865,N_16366);
xor U20319 (N_20319,N_14999,N_15282);
xnor U20320 (N_20320,N_17874,N_14408);
or U20321 (N_20321,N_13276,N_18516);
or U20322 (N_20322,N_15836,N_17408);
and U20323 (N_20323,N_14663,N_17947);
nand U20324 (N_20324,N_13223,N_12925);
or U20325 (N_20325,N_14691,N_15550);
or U20326 (N_20326,N_15998,N_17253);
xnor U20327 (N_20327,N_17734,N_14512);
nor U20328 (N_20328,N_16612,N_17764);
or U20329 (N_20329,N_15019,N_17612);
or U20330 (N_20330,N_16962,N_15010);
or U20331 (N_20331,N_18611,N_17037);
nand U20332 (N_20332,N_14207,N_12814);
nand U20333 (N_20333,N_12539,N_13257);
and U20334 (N_20334,N_12789,N_18618);
nand U20335 (N_20335,N_15450,N_17333);
nand U20336 (N_20336,N_15507,N_14013);
and U20337 (N_20337,N_17943,N_15323);
nand U20338 (N_20338,N_14799,N_13352);
xor U20339 (N_20339,N_17236,N_16268);
nor U20340 (N_20340,N_17918,N_18261);
nand U20341 (N_20341,N_15711,N_18675);
nand U20342 (N_20342,N_12953,N_16871);
or U20343 (N_20343,N_18686,N_16839);
xnor U20344 (N_20344,N_18591,N_13404);
nor U20345 (N_20345,N_18572,N_13931);
and U20346 (N_20346,N_16545,N_16993);
or U20347 (N_20347,N_16109,N_13140);
xor U20348 (N_20348,N_14375,N_15120);
nand U20349 (N_20349,N_15429,N_17193);
nand U20350 (N_20350,N_12725,N_17410);
nor U20351 (N_20351,N_16161,N_15195);
nand U20352 (N_20352,N_16812,N_15229);
nand U20353 (N_20353,N_18459,N_17010);
and U20354 (N_20354,N_17490,N_17173);
nor U20355 (N_20355,N_18065,N_18210);
nand U20356 (N_20356,N_17758,N_16500);
and U20357 (N_20357,N_13105,N_18620);
nor U20358 (N_20358,N_14757,N_14236);
xor U20359 (N_20359,N_16908,N_16401);
nor U20360 (N_20360,N_12545,N_12829);
and U20361 (N_20361,N_17805,N_16471);
nand U20362 (N_20362,N_17354,N_14064);
and U20363 (N_20363,N_17575,N_14150);
nor U20364 (N_20364,N_13648,N_14899);
and U20365 (N_20365,N_16537,N_17668);
nand U20366 (N_20366,N_14083,N_16336);
or U20367 (N_20367,N_17169,N_16931);
and U20368 (N_20368,N_13862,N_16720);
and U20369 (N_20369,N_14043,N_17106);
nor U20370 (N_20370,N_15398,N_12909);
and U20371 (N_20371,N_17870,N_14184);
xnor U20372 (N_20372,N_13660,N_14844);
and U20373 (N_20373,N_16885,N_14865);
nand U20374 (N_20374,N_16542,N_14486);
nand U20375 (N_20375,N_17182,N_17901);
nor U20376 (N_20376,N_15504,N_16902);
or U20377 (N_20377,N_15710,N_14169);
and U20378 (N_20378,N_16846,N_13829);
and U20379 (N_20379,N_18335,N_18651);
nor U20380 (N_20380,N_18519,N_18213);
nand U20381 (N_20381,N_16256,N_13109);
or U20382 (N_20382,N_15324,N_17201);
nor U20383 (N_20383,N_15148,N_13017);
and U20384 (N_20384,N_16055,N_15909);
nand U20385 (N_20385,N_13097,N_13932);
nor U20386 (N_20386,N_14221,N_14776);
nor U20387 (N_20387,N_15787,N_16078);
xnor U20388 (N_20388,N_14884,N_16681);
nor U20389 (N_20389,N_18460,N_13901);
or U20390 (N_20390,N_17705,N_17922);
xor U20391 (N_20391,N_12544,N_14044);
nor U20392 (N_20392,N_18352,N_17578);
or U20393 (N_20393,N_13733,N_14761);
and U20394 (N_20394,N_15265,N_17466);
xor U20395 (N_20395,N_14717,N_15310);
or U20396 (N_20396,N_18173,N_15827);
or U20397 (N_20397,N_15862,N_15098);
nor U20398 (N_20398,N_17619,N_13046);
nand U20399 (N_20399,N_17454,N_17358);
nand U20400 (N_20400,N_17144,N_17643);
nand U20401 (N_20401,N_17508,N_12523);
nor U20402 (N_20402,N_13711,N_15734);
nor U20403 (N_20403,N_16014,N_16623);
nor U20404 (N_20404,N_17356,N_13143);
or U20405 (N_20405,N_13467,N_12715);
nand U20406 (N_20406,N_18247,N_13410);
or U20407 (N_20407,N_18314,N_15240);
nand U20408 (N_20408,N_14040,N_14451);
nor U20409 (N_20409,N_16477,N_17763);
and U20410 (N_20410,N_18380,N_16305);
or U20411 (N_20411,N_14137,N_18339);
or U20412 (N_20412,N_18613,N_13141);
and U20413 (N_20413,N_15925,N_17391);
xnor U20414 (N_20414,N_13624,N_13087);
and U20415 (N_20415,N_14160,N_15471);
xnor U20416 (N_20416,N_12667,N_14759);
or U20417 (N_20417,N_18496,N_18243);
nor U20418 (N_20418,N_12936,N_13505);
and U20419 (N_20419,N_14735,N_13918);
or U20420 (N_20420,N_18114,N_16490);
nand U20421 (N_20421,N_16331,N_14533);
or U20422 (N_20422,N_18253,N_17744);
nor U20423 (N_20423,N_14574,N_16616);
nor U20424 (N_20424,N_14484,N_13167);
xnor U20425 (N_20425,N_18056,N_12524);
nand U20426 (N_20426,N_17932,N_15180);
nand U20427 (N_20427,N_14303,N_17670);
and U20428 (N_20428,N_18127,N_13921);
and U20429 (N_20429,N_13331,N_16190);
nand U20430 (N_20430,N_13869,N_12674);
nand U20431 (N_20431,N_12915,N_17683);
nor U20432 (N_20432,N_16023,N_14655);
nand U20433 (N_20433,N_15204,N_18068);
and U20434 (N_20434,N_14491,N_16127);
nor U20435 (N_20435,N_16263,N_17551);
and U20436 (N_20436,N_15040,N_17376);
and U20437 (N_20437,N_13254,N_14152);
or U20438 (N_20438,N_16296,N_16376);
nand U20439 (N_20439,N_14611,N_12827);
and U20440 (N_20440,N_18364,N_14284);
nand U20441 (N_20441,N_16311,N_16899);
or U20442 (N_20442,N_13983,N_15360);
or U20443 (N_20443,N_17696,N_12723);
nand U20444 (N_20444,N_16990,N_15027);
or U20445 (N_20445,N_17191,N_18489);
or U20446 (N_20446,N_12948,N_16933);
or U20447 (N_20447,N_15716,N_17234);
or U20448 (N_20448,N_18039,N_13602);
or U20449 (N_20449,N_17039,N_15889);
nor U20450 (N_20450,N_17916,N_18216);
xnor U20451 (N_20451,N_16552,N_13811);
or U20452 (N_20452,N_14404,N_13510);
nand U20453 (N_20453,N_16279,N_16758);
and U20454 (N_20454,N_14329,N_12964);
and U20455 (N_20455,N_18538,N_16431);
or U20456 (N_20456,N_18004,N_17280);
or U20457 (N_20457,N_14116,N_13036);
nor U20458 (N_20458,N_14745,N_16387);
xnor U20459 (N_20459,N_13001,N_12772);
xor U20460 (N_20460,N_13790,N_13824);
nor U20461 (N_20461,N_18589,N_13131);
and U20462 (N_20462,N_15535,N_17206);
nor U20463 (N_20463,N_15370,N_15496);
nor U20464 (N_20464,N_12615,N_17690);
or U20465 (N_20465,N_16813,N_14144);
and U20466 (N_20466,N_16325,N_14861);
and U20467 (N_20467,N_18020,N_14842);
nand U20468 (N_20468,N_16821,N_18640);
nand U20469 (N_20469,N_12565,N_15559);
nor U20470 (N_20470,N_17858,N_13471);
nor U20471 (N_20471,N_18357,N_16022);
nand U20472 (N_20472,N_15489,N_14962);
or U20473 (N_20473,N_18720,N_12844);
or U20474 (N_20474,N_15505,N_17440);
nor U20475 (N_20475,N_13182,N_12511);
nor U20476 (N_20476,N_15122,N_13076);
nor U20477 (N_20477,N_13314,N_16441);
and U20478 (N_20478,N_18403,N_12832);
and U20479 (N_20479,N_17252,N_18669);
nand U20480 (N_20480,N_13492,N_13521);
xnor U20481 (N_20481,N_13898,N_14940);
nand U20482 (N_20482,N_17593,N_13443);
and U20483 (N_20483,N_17214,N_17274);
or U20484 (N_20484,N_17806,N_14856);
nand U20485 (N_20485,N_14628,N_15663);
xor U20486 (N_20486,N_13804,N_18740);
nand U20487 (N_20487,N_18138,N_15712);
nor U20488 (N_20488,N_16991,N_14679);
nand U20489 (N_20489,N_16804,N_16975);
nor U20490 (N_20490,N_17984,N_14488);
and U20491 (N_20491,N_15751,N_12770);
nand U20492 (N_20492,N_15320,N_16643);
or U20493 (N_20493,N_16997,N_18179);
nand U20494 (N_20494,N_18378,N_13342);
or U20495 (N_20495,N_16533,N_16942);
and U20496 (N_20496,N_15720,N_13793);
or U20497 (N_20497,N_16313,N_13191);
nand U20498 (N_20498,N_17075,N_14086);
nor U20499 (N_20499,N_13813,N_16848);
nand U20500 (N_20500,N_15954,N_13784);
nor U20501 (N_20501,N_14975,N_13781);
and U20502 (N_20502,N_14541,N_15298);
nand U20503 (N_20503,N_17083,N_16573);
and U20504 (N_20504,N_15470,N_15932);
xnor U20505 (N_20505,N_16958,N_12537);
or U20506 (N_20506,N_13930,N_13933);
xnor U20507 (N_20507,N_17715,N_18242);
and U20508 (N_20508,N_13300,N_13159);
xor U20509 (N_20509,N_13155,N_16287);
nor U20510 (N_20510,N_16805,N_13504);
nand U20511 (N_20511,N_12945,N_12782);
or U20512 (N_20512,N_15525,N_17449);
nor U20513 (N_20513,N_16614,N_13994);
nor U20514 (N_20514,N_16802,N_15159);
nand U20515 (N_20515,N_14957,N_18369);
nand U20516 (N_20516,N_14820,N_14231);
nand U20517 (N_20517,N_13540,N_14528);
nand U20518 (N_20518,N_14702,N_15633);
nand U20519 (N_20519,N_18354,N_18450);
xnor U20520 (N_20520,N_13549,N_16476);
or U20521 (N_20521,N_12560,N_14153);
nand U20522 (N_20522,N_14693,N_17328);
and U20523 (N_20523,N_14746,N_16484);
nand U20524 (N_20524,N_14913,N_14588);
and U20525 (N_20525,N_13643,N_18639);
nand U20526 (N_20526,N_16655,N_17485);
nor U20527 (N_20527,N_12529,N_15654);
and U20528 (N_20528,N_14127,N_18677);
nand U20529 (N_20529,N_17903,N_14108);
and U20530 (N_20530,N_12729,N_18244);
nand U20531 (N_20531,N_14980,N_16222);
or U20532 (N_20532,N_12780,N_12739);
and U20533 (N_20533,N_17926,N_16051);
xnor U20534 (N_20534,N_13506,N_12568);
or U20535 (N_20535,N_17520,N_12864);
or U20536 (N_20536,N_17088,N_14514);
or U20537 (N_20537,N_13145,N_15187);
nor U20538 (N_20538,N_17240,N_17678);
nor U20539 (N_20539,N_17081,N_17813);
nor U20540 (N_20540,N_13258,N_16489);
and U20541 (N_20541,N_17681,N_18049);
or U20542 (N_20542,N_14900,N_14937);
or U20543 (N_20543,N_14877,N_18396);
nor U20544 (N_20544,N_18667,N_14346);
and U20545 (N_20545,N_16789,N_18507);
nor U20546 (N_20546,N_18234,N_17133);
or U20547 (N_20547,N_17818,N_12850);
nor U20548 (N_20548,N_17272,N_18109);
and U20549 (N_20549,N_15897,N_18557);
nand U20550 (N_20550,N_15199,N_15008);
and U20551 (N_20551,N_15842,N_14896);
and U20552 (N_20552,N_18650,N_17637);
or U20553 (N_20553,N_18602,N_18385);
nand U20554 (N_20554,N_14342,N_12978);
nand U20555 (N_20555,N_14910,N_12993);
nor U20556 (N_20556,N_15822,N_14263);
nor U20557 (N_20557,N_16700,N_14557);
or U20558 (N_20558,N_16208,N_17064);
nand U20559 (N_20559,N_18007,N_14965);
or U20560 (N_20560,N_16674,N_16429);
and U20561 (N_20561,N_14764,N_18702);
nor U20562 (N_20562,N_14359,N_17686);
nand U20563 (N_20563,N_13154,N_18250);
or U20564 (N_20564,N_13128,N_14227);
and U20565 (N_20565,N_15090,N_15103);
and U20566 (N_20566,N_14807,N_13268);
or U20567 (N_20567,N_13605,N_17437);
nand U20568 (N_20568,N_17843,N_13651);
and U20569 (N_20569,N_18265,N_14450);
or U20570 (N_20570,N_18010,N_17320);
and U20571 (N_20571,N_15206,N_15242);
nor U20572 (N_20572,N_14093,N_13846);
nand U20573 (N_20573,N_12806,N_14616);
nor U20574 (N_20574,N_17254,N_13249);
nand U20575 (N_20575,N_13866,N_18388);
nor U20576 (N_20576,N_14869,N_14248);
and U20577 (N_20577,N_16299,N_14750);
nor U20578 (N_20578,N_16058,N_16978);
nor U20579 (N_20579,N_15026,N_16457);
nor U20580 (N_20580,N_15311,N_16625);
or U20581 (N_20581,N_15138,N_16008);
nor U20582 (N_20582,N_14352,N_16395);
nand U20583 (N_20583,N_13865,N_16735);
and U20584 (N_20584,N_14812,N_13107);
and U20585 (N_20585,N_13272,N_13574);
or U20586 (N_20586,N_14593,N_17439);
or U20587 (N_20587,N_13760,N_13485);
nor U20588 (N_20588,N_15669,N_15769);
nor U20589 (N_20589,N_17672,N_17352);
and U20590 (N_20590,N_12802,N_13144);
nand U20591 (N_20591,N_17553,N_15202);
nand U20592 (N_20592,N_15817,N_16642);
or U20593 (N_20593,N_16067,N_15188);
and U20594 (N_20594,N_18300,N_18646);
nor U20595 (N_20595,N_16021,N_12736);
or U20596 (N_20596,N_18376,N_16989);
and U20597 (N_20597,N_13953,N_15523);
nor U20598 (N_20598,N_18633,N_14526);
or U20599 (N_20599,N_17293,N_15887);
nand U20600 (N_20600,N_15113,N_16007);
nor U20601 (N_20601,N_16121,N_15832);
or U20602 (N_20602,N_17290,N_17355);
nand U20603 (N_20603,N_18534,N_17682);
nor U20604 (N_20604,N_15273,N_12605);
nand U20605 (N_20605,N_14259,N_16383);
nor U20606 (N_20606,N_14253,N_13040);
nor U20607 (N_20607,N_14447,N_17529);
or U20608 (N_20608,N_15483,N_14947);
nor U20609 (N_20609,N_17373,N_16036);
nand U20610 (N_20610,N_15344,N_18428);
nand U20611 (N_20611,N_13500,N_16168);
or U20612 (N_20612,N_14596,N_16225);
nor U20613 (N_20613,N_18025,N_18483);
and U20614 (N_20614,N_12666,N_15404);
xnor U20615 (N_20615,N_15031,N_13235);
and U20616 (N_20616,N_17382,N_15178);
nand U20617 (N_20617,N_13078,N_17027);
and U20618 (N_20618,N_18002,N_18635);
nand U20619 (N_20619,N_17584,N_13986);
nor U20620 (N_20620,N_13900,N_16594);
and U20621 (N_20621,N_18245,N_18730);
or U20622 (N_20622,N_14215,N_17288);
or U20623 (N_20623,N_12735,N_17116);
nand U20624 (N_20624,N_14518,N_17611);
and U20625 (N_20625,N_16355,N_15177);
and U20626 (N_20626,N_16156,N_16142);
xnor U20627 (N_20627,N_18091,N_13016);
nor U20628 (N_20628,N_12867,N_18446);
nor U20629 (N_20629,N_16309,N_17934);
or U20630 (N_20630,N_13871,N_14233);
or U20631 (N_20631,N_15850,N_14036);
or U20632 (N_20632,N_15904,N_16729);
and U20633 (N_20633,N_14927,N_17595);
nor U20634 (N_20634,N_12963,N_13385);
nor U20635 (N_20635,N_13014,N_14564);
and U20636 (N_20636,N_13581,N_17931);
and U20637 (N_20637,N_14875,N_14521);
nor U20638 (N_20638,N_15153,N_16696);
and U20639 (N_20639,N_13503,N_16875);
or U20640 (N_20640,N_18734,N_18303);
and U20641 (N_20641,N_15652,N_16668);
and U20642 (N_20642,N_13979,N_15906);
or U20643 (N_20643,N_15592,N_14662);
xor U20644 (N_20644,N_17383,N_13635);
and U20645 (N_20645,N_14490,N_14030);
or U20646 (N_20646,N_13466,N_14469);
nor U20647 (N_20647,N_12794,N_12887);
nor U20648 (N_20648,N_12959,N_17588);
or U20649 (N_20649,N_14811,N_16026);
and U20650 (N_20650,N_15994,N_16451);
xnor U20651 (N_20651,N_17957,N_18523);
or U20652 (N_20652,N_15528,N_12939);
or U20653 (N_20653,N_15959,N_13712);
and U20654 (N_20654,N_15386,N_13496);
nand U20655 (N_20655,N_15224,N_13188);
xor U20656 (N_20656,N_15466,N_15431);
or U20657 (N_20657,N_13554,N_17583);
nor U20658 (N_20658,N_16780,N_14262);
nor U20659 (N_20659,N_14626,N_15201);
or U20660 (N_20660,N_12554,N_16734);
nand U20661 (N_20661,N_15805,N_18592);
or U20662 (N_20662,N_14755,N_18456);
and U20663 (N_20663,N_15561,N_15292);
or U20664 (N_20664,N_17960,N_16388);
nor U20665 (N_20665,N_13840,N_14911);
and U20666 (N_20666,N_12734,N_16739);
nand U20667 (N_20667,N_15108,N_16397);
nand U20668 (N_20668,N_18466,N_13479);
nor U20669 (N_20669,N_13339,N_16084);
nand U20670 (N_20670,N_17052,N_17150);
nand U20671 (N_20671,N_17543,N_14168);
nor U20672 (N_20672,N_13844,N_13633);
xnor U20673 (N_20673,N_16752,N_15313);
nand U20674 (N_20674,N_13606,N_18132);
xnor U20675 (N_20675,N_17921,N_18207);
or U20676 (N_20676,N_17138,N_15357);
nor U20677 (N_20677,N_12762,N_15503);
nor U20678 (N_20678,N_18426,N_16972);
nand U20679 (N_20679,N_18153,N_16820);
and U20680 (N_20680,N_16154,N_16213);
or U20681 (N_20681,N_16576,N_15804);
xnor U20682 (N_20682,N_14727,N_14441);
or U20683 (N_20683,N_14218,N_14966);
and U20684 (N_20684,N_16365,N_16410);
and U20685 (N_20685,N_16133,N_16065);
nor U20686 (N_20686,N_12760,N_17799);
nand U20687 (N_20687,N_17685,N_17388);
nand U20688 (N_20688,N_14964,N_18624);
xnor U20689 (N_20689,N_18568,N_13572);
nand U20690 (N_20690,N_15510,N_17337);
nor U20691 (N_20691,N_16122,N_14433);
nand U20692 (N_20692,N_15554,N_18647);
and U20693 (N_20693,N_17317,N_15086);
or U20694 (N_20694,N_13278,N_14255);
and U20695 (N_20695,N_18502,N_15047);
nor U20696 (N_20696,N_17202,N_13873);
and U20697 (N_20697,N_13734,N_15396);
or U20698 (N_20698,N_16324,N_16479);
or U20699 (N_20699,N_16170,N_17291);
nand U20700 (N_20700,N_14830,N_14948);
or U20701 (N_20701,N_18399,N_16856);
or U20702 (N_20702,N_12738,N_18405);
and U20703 (N_20703,N_13486,N_18642);
nor U20704 (N_20704,N_16531,N_13958);
nor U20705 (N_20705,N_13100,N_17822);
and U20706 (N_20706,N_17573,N_17165);
nand U20707 (N_20707,N_13260,N_16851);
and U20708 (N_20708,N_14331,N_17174);
xnor U20709 (N_20709,N_16445,N_17172);
nand U20710 (N_20710,N_15587,N_15335);
nor U20711 (N_20711,N_16162,N_16811);
and U20712 (N_20712,N_15697,N_16659);
or U20713 (N_20713,N_12777,N_15140);
nor U20714 (N_20714,N_13924,N_15568);
nor U20715 (N_20715,N_18576,N_13051);
and U20716 (N_20716,N_15435,N_14437);
and U20717 (N_20717,N_13653,N_14901);
and U20718 (N_20718,N_15863,N_14936);
nor U20719 (N_20719,N_18475,N_16657);
or U20720 (N_20720,N_14481,N_15170);
or U20721 (N_20721,N_15600,N_16093);
and U20722 (N_20722,N_16155,N_12671);
nor U20723 (N_20723,N_16658,N_15611);
xor U20724 (N_20724,N_13147,N_13940);
nand U20725 (N_20725,N_17846,N_17779);
nor U20726 (N_20726,N_13350,N_18102);
and U20727 (N_20727,N_18355,N_13721);
and U20728 (N_20728,N_15237,N_13458);
nand U20729 (N_20729,N_13514,N_12507);
nor U20730 (N_20730,N_16030,N_16086);
and U20731 (N_20731,N_17114,N_13055);
and U20732 (N_20732,N_18401,N_17063);
nand U20733 (N_20733,N_13005,N_13767);
nand U20734 (N_20734,N_13468,N_12696);
and U20735 (N_20735,N_13476,N_16283);
nand U20736 (N_20736,N_18248,N_12962);
or U20737 (N_20737,N_18046,N_15382);
nand U20738 (N_20738,N_14631,N_18692);
nand U20739 (N_20739,N_15493,N_18071);
nand U20740 (N_20740,N_14307,N_13112);
nor U20741 (N_20741,N_18559,N_18656);
xnor U20742 (N_20742,N_17464,N_13343);
nand U20743 (N_20743,N_13427,N_16496);
or U20744 (N_20744,N_12573,N_16973);
xnor U20745 (N_20745,N_17816,N_15414);
and U20746 (N_20746,N_15073,N_17061);
or U20747 (N_20747,N_13798,N_13743);
or U20748 (N_20748,N_14545,N_16151);
or U20749 (N_20749,N_17761,N_18358);
nor U20750 (N_20750,N_16183,N_12705);
nor U20751 (N_20751,N_16640,N_15222);
nor U20752 (N_20752,N_16678,N_18113);
and U20753 (N_20753,N_17600,N_15490);
xnor U20754 (N_20754,N_18468,N_14367);
nor U20755 (N_20755,N_13961,N_14026);
and U20756 (N_20756,N_16214,N_14380);
and U20757 (N_20757,N_15736,N_15629);
xnor U20758 (N_20758,N_15474,N_14585);
or U20759 (N_20759,N_15800,N_15881);
or U20760 (N_20760,N_16705,N_16923);
and U20761 (N_20761,N_14407,N_18044);
nand U20762 (N_20762,N_13187,N_14540);
and U20763 (N_20763,N_12668,N_14792);
or U20764 (N_20764,N_14550,N_15245);
nand U20765 (N_20765,N_18681,N_18671);
xor U20766 (N_20766,N_16374,N_17949);
nor U20767 (N_20767,N_17900,N_13752);
nor U20768 (N_20768,N_14333,N_16855);
nor U20769 (N_20769,N_15580,N_12624);
xor U20770 (N_20770,N_13576,N_17073);
or U20771 (N_20771,N_17524,N_18679);
nor U20772 (N_20772,N_13090,N_16713);
xnor U20773 (N_20773,N_13317,N_14252);
xor U20774 (N_20774,N_17029,N_13106);
nor U20775 (N_20775,N_17864,N_14982);
nor U20776 (N_20776,N_14598,N_13937);
nand U20777 (N_20777,N_17229,N_17390);
xor U20778 (N_20778,N_13754,N_15876);
nand U20779 (N_20779,N_16591,N_15762);
and U20780 (N_20780,N_17791,N_12765);
xnor U20781 (N_20781,N_18735,N_15462);
xor U20782 (N_20782,N_16492,N_13428);
nor U20783 (N_20783,N_17940,N_17404);
xnor U20784 (N_20784,N_14142,N_13663);
nor U20785 (N_20785,N_18104,N_16913);
nand U20786 (N_20786,N_18288,N_14791);
or U20787 (N_20787,N_12771,N_17618);
and U20788 (N_20788,N_17158,N_16308);
or U20789 (N_20789,N_15539,N_16128);
nor U20790 (N_20790,N_17118,N_15677);
nor U20791 (N_20791,N_13195,N_16691);
or U20792 (N_20792,N_15304,N_18550);
nand U20793 (N_20793,N_18530,N_14934);
nor U20794 (N_20794,N_12703,N_16656);
or U20795 (N_20795,N_15870,N_14332);
nor U20796 (N_20796,N_16830,N_14831);
nand U20797 (N_20797,N_18251,N_16740);
nor U20798 (N_20798,N_15538,N_14733);
nand U20799 (N_20799,N_13524,N_18571);
nand U20800 (N_20800,N_17484,N_16089);
or U20801 (N_20801,N_15218,N_12661);
or U20802 (N_20802,N_17554,N_18093);
nor U20803 (N_20803,N_18214,N_18168);
and U20804 (N_20804,N_18313,N_15594);
or U20805 (N_20805,N_13084,N_13495);
or U20806 (N_20806,N_12637,N_14579);
nor U20807 (N_20807,N_14340,N_12897);
and U20808 (N_20808,N_15513,N_14827);
nor U20809 (N_20809,N_16404,N_16685);
nand U20810 (N_20810,N_13202,N_14223);
and U20811 (N_20811,N_14551,N_12904);
nor U20812 (N_20812,N_12934,N_13668);
or U20813 (N_20813,N_18282,N_18273);
and U20814 (N_20814,N_15814,N_12819);
or U20815 (N_20815,N_12692,N_14798);
and U20816 (N_20816,N_15619,N_18304);
or U20817 (N_20817,N_15763,N_15318);
nor U20818 (N_20818,N_14868,N_18139);
nor U20819 (N_20819,N_15908,N_12968);
nand U20820 (N_20820,N_16653,N_15591);
nand U20821 (N_20821,N_15668,N_16633);
nand U20822 (N_20822,N_16834,N_17393);
xor U20823 (N_20823,N_16980,N_18739);
and U20824 (N_20824,N_16661,N_12599);
or U20825 (N_20825,N_18452,N_18387);
nor U20826 (N_20826,N_16226,N_17160);
xnor U20827 (N_20827,N_16595,N_17377);
xor U20828 (N_20828,N_18302,N_18654);
and U20829 (N_20829,N_13234,N_12856);
or U20830 (N_20830,N_17218,N_15606);
nor U20831 (N_20831,N_15678,N_17972);
nor U20832 (N_20832,N_17327,N_12699);
nand U20833 (N_20833,N_13446,N_17212);
nand U20834 (N_20834,N_14471,N_18597);
nor U20835 (N_20835,N_16606,N_13318);
xor U20836 (N_20836,N_15032,N_14238);
nand U20837 (N_20837,N_17790,N_16857);
or U20838 (N_20838,N_13975,N_14458);
or U20839 (N_20839,N_14410,N_16516);
nand U20840 (N_20840,N_14125,N_16312);
nor U20841 (N_20841,N_17422,N_17658);
nor U20842 (N_20842,N_17313,N_12754);
and U20843 (N_20843,N_12517,N_17729);
nand U20844 (N_20844,N_13714,N_15173);
and U20845 (N_20845,N_15970,N_16778);
xnor U20846 (N_20846,N_14802,N_17446);
xor U20847 (N_20847,N_18477,N_15824);
nand U20848 (N_20848,N_13604,N_15564);
nand U20849 (N_20849,N_17847,N_14763);
nor U20850 (N_20850,N_13652,N_17375);
or U20851 (N_20851,N_16592,N_17302);
nor U20852 (N_20852,N_17756,N_16077);
nand U20853 (N_20853,N_17802,N_12851);
or U20854 (N_20854,N_15051,N_12683);
xor U20855 (N_20855,N_14304,N_13582);
nor U20856 (N_20856,N_13319,N_15472);
nand U20857 (N_20857,N_14555,N_12774);
nand U20858 (N_20858,N_14415,N_15294);
xor U20859 (N_20859,N_13228,N_18434);
xor U20860 (N_20860,N_17260,N_15743);
or U20861 (N_20861,N_14349,N_18517);
and U20862 (N_20862,N_12878,N_15433);
or U20863 (N_20863,N_17351,N_13388);
and U20864 (N_20864,N_15766,N_13552);
nor U20865 (N_20865,N_13715,N_15570);
nor U20866 (N_20866,N_12855,N_17018);
nand U20867 (N_20867,N_17111,N_14684);
nor U20868 (N_20868,N_18443,N_14995);
and U20869 (N_20869,N_15376,N_14197);
or U20870 (N_20870,N_12929,N_18417);
or U20871 (N_20871,N_12590,N_15576);
xnor U20872 (N_20872,N_15209,N_16238);
nand U20873 (N_20873,N_14530,N_13196);
or U20874 (N_20874,N_13637,N_18169);
or U20875 (N_20875,N_13450,N_16953);
nor U20876 (N_20876,N_13957,N_13212);
nand U20877 (N_20877,N_16337,N_14149);
and U20878 (N_20878,N_14314,N_13305);
and U20879 (N_20879,N_17213,N_13612);
nor U20880 (N_20880,N_15262,N_17783);
nand U20881 (N_20881,N_14357,N_12652);
or U20882 (N_20882,N_15723,N_16938);
nand U20883 (N_20883,N_15533,N_18615);
nor U20884 (N_20884,N_14206,N_12633);
or U20885 (N_20885,N_16468,N_15929);
nor U20886 (N_20886,N_18391,N_12824);
or U20887 (N_20887,N_16779,N_13776);
or U20888 (N_20888,N_16715,N_18491);
nand U20889 (N_20889,N_14949,N_13952);
or U20890 (N_20890,N_17817,N_18663);
nor U20891 (N_20891,N_16904,N_14642);
and U20892 (N_20892,N_18430,N_15796);
and U20893 (N_20893,N_18562,N_14322);
nand U20894 (N_20894,N_17987,N_14115);
nor U20895 (N_20895,N_15729,N_12660);
nor U20896 (N_20896,N_12906,N_17208);
or U20897 (N_20897,N_13820,N_17366);
and U20898 (N_20898,N_12971,N_16562);
nand U20899 (N_20899,N_15352,N_13982);
or U20900 (N_20900,N_16491,N_15864);
nand U20901 (N_20901,N_15207,N_15105);
nor U20902 (N_20902,N_17433,N_14848);
and U20903 (N_20903,N_18659,N_16119);
nor U20904 (N_20904,N_13091,N_16836);
nand U20905 (N_20905,N_16110,N_14781);
nand U20906 (N_20906,N_13421,N_13429);
or U20907 (N_20907,N_14904,N_12557);
nand U20908 (N_20908,N_14803,N_15595);
nor U20909 (N_20909,N_12837,N_13000);
and U20910 (N_20910,N_13309,N_16840);
nand U20911 (N_20911,N_15747,N_16094);
and U20912 (N_20912,N_13757,N_15681);
and U20913 (N_20913,N_17669,N_16832);
or U20914 (N_20914,N_15553,N_15154);
xor U20915 (N_20915,N_15260,N_15746);
nor U20916 (N_20916,N_17688,N_17606);
or U20917 (N_20917,N_17062,N_18236);
nor U20918 (N_20918,N_14507,N_14850);
or U20919 (N_20919,N_14140,N_13837);
nor U20920 (N_20920,N_17564,N_15885);
and U20921 (N_20921,N_12889,N_17702);
nor U20922 (N_20922,N_16257,N_17886);
or U20923 (N_20923,N_13346,N_17386);
nand U20924 (N_20924,N_13085,N_14916);
nand U20925 (N_20925,N_15034,N_14182);
and U20926 (N_20926,N_18712,N_16242);
nand U20927 (N_20927,N_13826,N_16400);
nor U20928 (N_20928,N_12812,N_13636);
nor U20929 (N_20929,N_17721,N_12669);
nor U20930 (N_20930,N_13066,N_17845);
or U20931 (N_20931,N_18716,N_18402);
or U20932 (N_20932,N_14102,N_13638);
xor U20933 (N_20933,N_13282,N_17753);
and U20934 (N_20934,N_14709,N_16215);
nor U20935 (N_20935,N_17239,N_18393);
and U20936 (N_20936,N_13330,N_16462);
and U20937 (N_20937,N_13632,N_18095);
nor U20938 (N_20938,N_16250,N_17459);
or U20939 (N_20939,N_13628,N_16983);
and U20940 (N_20940,N_17645,N_15506);
nand U20941 (N_20941,N_15963,N_15442);
nand U20942 (N_20942,N_16762,N_12575);
or U20943 (N_20943,N_14278,N_15662);
nor U20944 (N_20944,N_13382,N_13321);
and U20945 (N_20945,N_16466,N_12547);
nand U20946 (N_20946,N_15309,N_13917);
and U20947 (N_20947,N_15048,N_15217);
or U20948 (N_20948,N_15758,N_15024);
or U20949 (N_20949,N_15487,N_14472);
and U20950 (N_20950,N_14996,N_18695);
nand U20951 (N_20951,N_18175,N_17774);
and U20952 (N_20952,N_13175,N_13252);
and U20953 (N_20953,N_17360,N_12931);
or U20954 (N_20954,N_15364,N_16137);
and U20955 (N_20955,N_15106,N_14103);
and U20956 (N_20956,N_14639,N_13362);
and U20957 (N_20957,N_15610,N_12998);
nor U20958 (N_20958,N_18342,N_15145);
or U20959 (N_20959,N_16465,N_16600);
nand U20960 (N_20960,N_16541,N_15125);
nor U20961 (N_20961,N_15542,N_15714);
and U20962 (N_20962,N_15514,N_15132);
or U20963 (N_20963,N_18710,N_14973);
or U20964 (N_20964,N_16071,N_17146);
and U20965 (N_20965,N_14956,N_17000);
and U20966 (N_20966,N_12795,N_17241);
and U20967 (N_20967,N_17054,N_16046);
xor U20968 (N_20968,N_13611,N_17592);
or U20969 (N_20969,N_12826,N_17019);
nand U20970 (N_20970,N_14059,N_16187);
nor U20971 (N_20971,N_17164,N_16544);
nand U20972 (N_20972,N_13075,N_14573);
xnor U20973 (N_20973,N_14617,N_18696);
nor U20974 (N_20974,N_12567,N_17814);
nand U20975 (N_20975,N_16587,N_15775);
and U20976 (N_20976,N_13809,N_12540);
or U20977 (N_20977,N_17276,N_13806);
nand U20978 (N_20978,N_18420,N_12997);
nor U20979 (N_20979,N_15638,N_14316);
or U20980 (N_20980,N_17879,N_18660);
and U20981 (N_20981,N_16632,N_16295);
nor U20982 (N_20982,N_13125,N_16637);
nor U20983 (N_20983,N_12988,N_13436);
or U20984 (N_20984,N_17368,N_13019);
and U20985 (N_20985,N_13872,N_16418);
or U20986 (N_20986,N_17782,N_12612);
xor U20987 (N_20987,N_14465,N_16372);
nand U20988 (N_20988,N_14867,N_13762);
and U20989 (N_20989,N_15621,N_13454);
and U20990 (N_20990,N_17470,N_18055);
nand U20991 (N_20991,N_16853,N_13799);
nand U20992 (N_20992,N_12932,N_18033);
and U20993 (N_20993,N_15052,N_17040);
nor U20994 (N_20994,N_15598,N_18198);
nand U20995 (N_20995,N_17334,N_17341);
nand U20996 (N_20996,N_15705,N_12761);
and U20997 (N_20997,N_16827,N_15641);
nor U20998 (N_20998,N_15837,N_15706);
xnor U20999 (N_20999,N_15790,N_14941);
xnor U21000 (N_21000,N_14539,N_16249);
nand U21001 (N_21001,N_13012,N_13543);
and U21002 (N_21002,N_15868,N_13702);
xnor U21003 (N_21003,N_17175,N_12664);
nand U21004 (N_21004,N_12525,N_13948);
xor U21005 (N_21005,N_16433,N_12937);
and U21006 (N_21006,N_17294,N_17305);
and U21007 (N_21007,N_14608,N_13345);
or U21008 (N_21008,N_15795,N_15158);
nor U21009 (N_21009,N_14374,N_13641);
nor U21010 (N_21010,N_15235,N_17478);
or U21011 (N_21011,N_13841,N_16590);
nand U21012 (N_21012,N_13550,N_12582);
nor U21013 (N_21013,N_15738,N_13926);
or U21014 (N_21014,N_18141,N_16731);
nand U21015 (N_21015,N_16507,N_18074);
xor U21016 (N_21016,N_13295,N_17528);
nor U21017 (N_21017,N_17219,N_15463);
or U21018 (N_21018,N_17624,N_15995);
xor U21019 (N_21019,N_18238,N_17273);
nand U21020 (N_21020,N_18230,N_14688);
and U21021 (N_21021,N_13976,N_18003);
nand U21022 (N_21022,N_15526,N_15686);
nor U21023 (N_21023,N_13879,N_14918);
or U21024 (N_21024,N_15933,N_18130);
nand U21025 (N_21025,N_14309,N_15296);
nor U21026 (N_21026,N_14443,N_16586);
nand U21027 (N_21027,N_16519,N_18741);
nand U21028 (N_21028,N_17399,N_14568);
nand U21029 (N_21029,N_14546,N_12905);
or U21030 (N_21030,N_15657,N_12534);
or U21031 (N_21031,N_17872,N_16050);
or U21032 (N_21032,N_12750,N_12676);
nor U21033 (N_21033,N_12687,N_12946);
nor U21034 (N_21034,N_15359,N_16631);
and U21035 (N_21035,N_18487,N_17065);
xnor U21036 (N_21036,N_16610,N_14567);
nand U21037 (N_21037,N_18269,N_18721);
nand U21038 (N_21038,N_16147,N_13173);
nand U21039 (N_21039,N_16867,N_16134);
nand U21040 (N_21040,N_15271,N_17911);
nor U21041 (N_21041,N_16011,N_14011);
or U21042 (N_21042,N_16193,N_14289);
or U21043 (N_21043,N_13626,N_15585);
or U21044 (N_21044,N_14597,N_14350);
and U21045 (N_21045,N_17692,N_15129);
nor U21046 (N_21046,N_14436,N_16049);
and U21047 (N_21047,N_17319,N_17881);
or U21048 (N_21048,N_13947,N_16481);
and U21049 (N_21049,N_13351,N_14476);
nand U21050 (N_21050,N_14692,N_14020);
or U21051 (N_21051,N_15811,N_14613);
nor U21052 (N_21052,N_16554,N_13006);
nand U21053 (N_21053,N_17775,N_12786);
nand U21054 (N_21054,N_18221,N_16390);
nand U21055 (N_21055,N_13991,N_17457);
nor U21056 (N_21056,N_12635,N_15894);
and U21057 (N_21057,N_15756,N_15983);
nor U21058 (N_21058,N_16679,N_18480);
nand U21059 (N_21059,N_18389,N_15306);
nand U21060 (N_21060,N_16996,N_16179);
and U21061 (N_21061,N_15044,N_15411);
xor U21062 (N_21062,N_15742,N_13995);
nand U21063 (N_21063,N_17405,N_14302);
and U21064 (N_21064,N_14801,N_17503);
nand U21065 (N_21065,N_18368,N_16651);
and U21066 (N_21066,N_16227,N_16814);
xnor U21067 (N_21067,N_17346,N_14944);
and U21068 (N_21068,N_16027,N_15991);
or U21069 (N_21069,N_13420,N_15588);
nor U21070 (N_21070,N_17837,N_12559);
nor U21071 (N_21071,N_13616,N_17969);
or U21072 (N_21072,N_13209,N_13523);
and U21073 (N_21073,N_18366,N_17006);
or U21074 (N_21074,N_15495,N_16482);
nor U21075 (N_21075,N_15700,N_14586);
or U21076 (N_21076,N_18254,N_18349);
nor U21077 (N_21077,N_13440,N_15448);
nand U21078 (N_21078,N_12717,N_17247);
and U21079 (N_21079,N_18189,N_15445);
nand U21080 (N_21080,N_15133,N_16749);
and U21081 (N_21081,N_16707,N_14012);
or U21082 (N_21082,N_16872,N_12983);
nand U21083 (N_21083,N_15267,N_14516);
or U21084 (N_21084,N_16797,N_14989);
and U21085 (N_21085,N_18225,N_15264);
nor U21086 (N_21086,N_14767,N_16529);
xnor U21087 (N_21087,N_16413,N_14499);
nor U21088 (N_21088,N_17777,N_15136);
xor U21089 (N_21089,N_13619,N_14170);
or U21090 (N_21090,N_14132,N_17511);
and U21091 (N_21091,N_14440,N_16937);
nand U21092 (N_21092,N_12621,N_14723);
nand U21093 (N_21093,N_15527,N_15097);
xor U21094 (N_21094,N_17095,N_18201);
and U21095 (N_21095,N_17093,N_13355);
or U21096 (N_21096,N_15784,N_16384);
nand U21097 (N_21097,N_18462,N_18435);
or U21098 (N_21098,N_12527,N_12695);
nand U21099 (N_21099,N_16721,N_15986);
nor U21100 (N_21100,N_16549,N_14822);
nor U21101 (N_21101,N_14070,N_13132);
or U21102 (N_21102,N_17509,N_15498);
and U21103 (N_21103,N_17570,N_17896);
nand U21104 (N_21104,N_12809,N_12881);
nand U21105 (N_21105,N_17635,N_16343);
nor U21106 (N_21106,N_14656,N_13459);
nand U21107 (N_21107,N_17468,N_14422);
and U21108 (N_21108,N_17634,N_14796);
xnor U21109 (N_21109,N_13782,N_13649);
nand U21110 (N_21110,N_13907,N_18192);
and U21111 (N_21111,N_18390,N_15055);
or U21112 (N_21112,N_18515,N_15578);
and U21113 (N_21113,N_12578,N_15288);
or U21114 (N_21114,N_15155,N_15277);
nor U21115 (N_21115,N_13118,N_18162);
nand U21116 (N_21116,N_14836,N_16495);
or U21117 (N_21117,N_13337,N_16994);
or U21118 (N_21118,N_14645,N_13199);
nand U21119 (N_21119,N_15295,N_13701);
nand U21120 (N_21120,N_12555,N_16921);
xnor U21121 (N_21121,N_14183,N_16501);
nand U21122 (N_21122,N_18601,N_16132);
nor U21123 (N_21123,N_12566,N_13073);
xor U21124 (N_21124,N_12752,N_18084);
and U21125 (N_21125,N_12564,N_16080);
and U21126 (N_21126,N_18689,N_13678);
and U21127 (N_21127,N_18182,N_13053);
or U21128 (N_21128,N_13925,N_13884);
nand U21129 (N_21129,N_15750,N_17694);
and U21130 (N_21130,N_14032,N_13462);
and U21131 (N_21131,N_18614,N_18106);
nand U21132 (N_21132,N_14704,N_13985);
or U21133 (N_21133,N_14697,N_18289);
xor U21134 (N_21134,N_13103,N_16825);
or U21135 (N_21135,N_12787,N_17552);
and U21136 (N_21136,N_13738,N_16847);
nand U21137 (N_21137,N_17929,N_15645);
or U21138 (N_21138,N_15375,N_16667);
and U21139 (N_21139,N_12681,N_15146);
nand U21140 (N_21140,N_14225,N_12742);
and U21141 (N_21141,N_16630,N_17582);
and U21142 (N_21142,N_15582,N_16808);
xor U21143 (N_21143,N_13709,N_15059);
xor U21144 (N_21144,N_15791,N_14590);
nor U21145 (N_21145,N_18486,N_15014);
or U21146 (N_21146,N_16047,N_16163);
nor U21147 (N_21147,N_17759,N_13603);
nand U21148 (N_21148,N_18664,N_15679);
and U21149 (N_21149,N_16302,N_15616);
and U21150 (N_21150,N_12894,N_17321);
or U21151 (N_21151,N_14853,N_15938);
nand U21152 (N_21152,N_18023,N_16292);
nor U21153 (N_21153,N_13830,N_15461);
or U21154 (N_21154,N_18411,N_16016);
or U21155 (N_21155,N_17542,N_13856);
and U21156 (N_21156,N_15847,N_15614);
or U21157 (N_21157,N_18334,N_17880);
nor U21158 (N_21158,N_13119,N_16746);
xnor U21159 (N_21159,N_17292,N_16202);
and U21160 (N_21160,N_18126,N_18164);
and U21161 (N_21161,N_14961,N_12731);
and U21162 (N_21162,N_17181,N_16038);
or U21163 (N_21163,N_17829,N_16970);
nor U21164 (N_21164,N_13165,N_15687);
nand U21165 (N_21165,N_17221,N_17828);
xor U21166 (N_21166,N_13694,N_12716);
nor U21167 (N_21167,N_14615,N_17344);
nor U21168 (N_21168,N_18678,N_17369);
or U21169 (N_21169,N_16218,N_14621);
nor U21170 (N_21170,N_14308,N_15988);
nand U21171 (N_21171,N_17246,N_17803);
or U21172 (N_21172,N_13377,N_16291);
and U21173 (N_21173,N_12514,N_12831);
or U21174 (N_21174,N_14406,N_15214);
and U21175 (N_21175,N_12608,N_14124);
nor U21176 (N_21176,N_17707,N_15676);
or U21177 (N_21177,N_15350,N_14485);
nand U21178 (N_21178,N_18727,N_12638);
nand U21179 (N_21179,N_15979,N_16351);
xnor U21180 (N_21180,N_13379,N_17513);
and U21181 (N_21181,N_17074,N_12543);
nand U21182 (N_21182,N_15116,N_14641);
nor U21183 (N_21183,N_13095,N_18305);
and U21184 (N_21184,N_14549,N_14701);
nand U21185 (N_21185,N_17338,N_15707);
nor U21186 (N_21186,N_17032,N_17312);
or U21187 (N_21187,N_16105,N_14067);
nand U21188 (N_21188,N_14607,N_17418);
xor U21189 (N_21189,N_12960,N_15196);
nand U21190 (N_21190,N_17577,N_16303);
nor U21191 (N_21191,N_18479,N_18657);
or U21192 (N_21192,N_12740,N_15802);
nand U21193 (N_21193,N_17861,N_16074);
or U21194 (N_21194,N_15415,N_18471);
or U21195 (N_21195,N_16521,N_15198);
and U21196 (N_21196,N_17976,N_18439);
and U21197 (N_21197,N_15634,N_17481);
or U21198 (N_21198,N_15509,N_15142);
and U21199 (N_21199,N_13788,N_14630);
or U21200 (N_21200,N_13281,N_15993);
nor U21201 (N_21201,N_16239,N_15684);
nand U21202 (N_21202,N_14897,N_18554);
nor U21203 (N_21203,N_18569,N_17362);
nand U21204 (N_21204,N_16344,N_16654);
xor U21205 (N_21205,N_17069,N_16744);
nor U21206 (N_21206,N_14903,N_14254);
and U21207 (N_21207,N_16878,N_18115);
or U21208 (N_21208,N_13690,N_17751);
nor U21209 (N_21209,N_13402,N_15299);
and U21210 (N_21210,N_12720,N_13875);
nand U21211 (N_21211,N_16555,N_14666);
and U21212 (N_21212,N_18374,N_14987);
and U21213 (N_21213,N_16880,N_15259);
and U21214 (N_21214,N_18310,N_15137);
or U21215 (N_21215,N_17472,N_17946);
and U21216 (N_21216,N_18697,N_16703);
nand U21217 (N_21217,N_17599,N_15284);
nand U21218 (N_21218,N_14985,N_17977);
or U21219 (N_21219,N_16020,N_13538);
or U21220 (N_21220,N_12907,N_15481);
or U21221 (N_21221,N_16330,N_14445);
or U21222 (N_21222,N_14922,N_14112);
or U21223 (N_21223,N_12888,N_14283);
and U21224 (N_21224,N_13534,N_17998);
nor U21225 (N_21225,N_16892,N_17648);
and U21226 (N_21226,N_17961,N_12811);
or U21227 (N_21227,N_16171,N_15017);
nor U21228 (N_21228,N_14625,N_15151);
or U21229 (N_21229,N_14393,N_15036);
and U21230 (N_21230,N_12505,N_15373);
nand U21231 (N_21231,N_17070,N_15427);
and U21232 (N_21232,N_16307,N_15945);
nand U21233 (N_21233,N_13680,N_18594);
or U21234 (N_21234,N_14520,N_13096);
or U21235 (N_21235,N_15717,N_15753);
and U21236 (N_21236,N_17381,N_17417);
and U21237 (N_21237,N_14765,N_17518);
nor U21238 (N_21238,N_16894,N_13675);
or U21239 (N_21239,N_14048,N_16483);
nand U21240 (N_21240,N_16289,N_13286);
and U21241 (N_21241,N_13231,N_12737);
or U21242 (N_21242,N_15947,N_18051);
nor U21243 (N_21243,N_14624,N_16745);
and U21244 (N_21244,N_12944,N_17289);
xnor U21245 (N_21245,N_15069,N_18662);
nor U21246 (N_21246,N_18726,N_15581);
xnor U21247 (N_21247,N_14425,N_16025);
nor U21248 (N_21248,N_17423,N_18652);
nand U21249 (N_21249,N_18520,N_15961);
or U21250 (N_21250,N_13240,N_14019);
and U21251 (N_21251,N_18747,N_12877);
and U21252 (N_21252,N_17184,N_16060);
nor U21253 (N_21253,N_14926,N_14972);
nor U21254 (N_21254,N_14388,N_12798);
nand U21255 (N_21255,N_15361,N_18285);
xnor U21256 (N_21256,N_13414,N_13578);
or U21257 (N_21257,N_17066,N_15243);
or U21258 (N_21258,N_15524,N_17614);
and U21259 (N_21259,N_12504,N_14239);
nor U21260 (N_21260,N_18384,N_16648);
nand U21261 (N_21261,N_14563,N_17397);
and U21262 (N_21262,N_16399,N_17035);
or U21263 (N_21263,N_15821,N_17851);
or U21264 (N_21264,N_16776,N_17059);
nor U21265 (N_21265,N_16042,N_13746);
nand U21266 (N_21266,N_18604,N_15785);
nand U21267 (N_21267,N_18257,N_16474);
or U21268 (N_21268,N_16357,N_12873);
nor U21269 (N_21269,N_17788,N_16775);
xnor U21270 (N_21270,N_16532,N_15874);
or U21271 (N_21271,N_15967,N_16001);
nor U21272 (N_21272,N_17442,N_16236);
nor U21273 (N_21273,N_18043,N_16181);
and U21274 (N_21274,N_14279,N_13780);
xor U21275 (N_21275,N_15405,N_15866);
nor U21276 (N_21276,N_15936,N_12796);
nor U21277 (N_21277,N_17009,N_14722);
xnor U21278 (N_21278,N_17284,N_15246);
nand U21279 (N_21279,N_13127,N_17235);
and U21280 (N_21280,N_16316,N_18577);
nand U21281 (N_21281,N_15698,N_17627);
xnor U21282 (N_21282,N_12805,N_16435);
or U21283 (N_21283,N_17179,N_14912);
nor U21284 (N_21284,N_15353,N_18124);
nor U21285 (N_21285,N_16861,N_15690);
nor U21286 (N_21286,N_18155,N_12957);
and U21287 (N_21287,N_15776,N_15365);
nand U21288 (N_21288,N_16669,N_15930);
nor U21289 (N_21289,N_13698,N_17094);
nand U21290 (N_21290,N_13494,N_18080);
nand U21291 (N_21291,N_17316,N_18529);
nor U21292 (N_21292,N_12620,N_15285);
and U21293 (N_21293,N_18371,N_15194);
or U21294 (N_21294,N_12863,N_16111);
and U21295 (N_21295,N_14829,N_18706);
nor U21296 (N_21296,N_13993,N_12766);
nor U21297 (N_21297,N_15349,N_13411);
xor U21298 (N_21298,N_18070,N_14411);
nor U21299 (N_21299,N_17954,N_14824);
or U21300 (N_21300,N_16611,N_18549);
or U21301 (N_21301,N_13063,N_16818);
and U21302 (N_21302,N_16327,N_16360);
nand U21303 (N_21303,N_14363,N_16764);
and U21304 (N_21304,N_15160,N_18064);
and U21305 (N_21305,N_17186,N_18684);
nand U21306 (N_21306,N_18108,N_13868);
and U21307 (N_21307,N_16662,N_12842);
or U21308 (N_21308,N_15801,N_14061);
xnor U21309 (N_21309,N_13166,N_13751);
and U21310 (N_21310,N_17821,N_17907);
or U21311 (N_21311,N_14778,N_16333);
nor U21312 (N_21312,N_17609,N_17989);
nor U21313 (N_21313,N_14272,N_14977);
nand U21314 (N_21314,N_14771,N_16816);
nand U21315 (N_21315,N_15249,N_15978);
nor U21316 (N_21316,N_17848,N_18619);
and U21317 (N_21317,N_15786,N_14232);
nor U21318 (N_21318,N_14954,N_14203);
nand U21319 (N_21319,N_17504,N_16896);
and U21320 (N_21320,N_16914,N_14878);
or U21321 (N_21321,N_12581,N_17458);
xor U21322 (N_21322,N_18630,N_16858);
nor U21323 (N_21323,N_13463,N_12870);
or U21324 (N_21324,N_13163,N_14212);
and U21325 (N_21325,N_16286,N_16823);
nor U21326 (N_21326,N_16464,N_16844);
and U21327 (N_21327,N_17560,N_13970);
and U21328 (N_21328,N_16270,N_13575);
nor U21329 (N_21329,N_17170,N_12938);
nor U21330 (N_21330,N_16210,N_15127);
nand U21331 (N_21331,N_16261,N_13082);
nand U21332 (N_21332,N_16897,N_17412);
or U21333 (N_21333,N_18306,N_13544);
nand U21334 (N_21334,N_18073,N_14338);
and U21335 (N_21335,N_12707,N_16609);
and U21336 (N_21336,N_15749,N_17026);
or U21337 (N_21337,N_13912,N_18609);
and U21338 (N_21338,N_14270,N_13130);
or U21339 (N_21339,N_18743,N_18340);
and U21340 (N_21340,N_14810,N_17742);
nand U21341 (N_21341,N_15083,N_15643);
or U21342 (N_21342,N_18119,N_15819);
and U21343 (N_21343,N_13818,N_14524);
nor U21344 (N_21344,N_16558,N_14482);
and U21345 (N_21345,N_13032,N_18467);
xor U21346 (N_21346,N_16085,N_17425);
and U21347 (N_21347,N_13659,N_18163);
nand U21348 (N_21348,N_14678,N_14600);
or U21349 (N_21349,N_16348,N_13922);
nand U21350 (N_21350,N_15910,N_15499);
and U21351 (N_21351,N_14216,N_16186);
xor U21352 (N_21352,N_15283,N_17988);
nor U21353 (N_21353,N_14843,N_15485);
and U21354 (N_21354,N_14714,N_17964);
nand U21355 (N_21355,N_16166,N_17151);
nand U21356 (N_21356,N_16373,N_15829);
nor U21357 (N_21357,N_18149,N_13065);
or U21358 (N_21358,N_15974,N_14261);
nand U21359 (N_21359,N_13664,N_16112);
or U21360 (N_21360,N_14923,N_16140);
nor U21361 (N_21361,N_17092,N_13031);
or U21362 (N_21362,N_18733,N_15250);
nand U21363 (N_21363,N_13851,N_17285);
nor U21364 (N_21364,N_17530,N_15971);
nand U21365 (N_21365,N_13301,N_14268);
or U21366 (N_21366,N_15981,N_18714);
nor U21367 (N_21367,N_18227,N_12876);
xnor U21368 (N_21368,N_16432,N_14101);
nor U21369 (N_21369,N_15725,N_17278);
xnor U21370 (N_21370,N_12609,N_13693);
nor U21371 (N_21371,N_17675,N_14519);
or U21372 (N_21372,N_17326,N_14648);
and U21373 (N_21373,N_15412,N_13938);
and U21374 (N_21374,N_16863,N_12996);
nand U21375 (N_21375,N_14522,N_15395);
nor U21376 (N_21376,N_15632,N_14483);
or U21377 (N_21377,N_16936,N_15332);
nand U21378 (N_21378,N_13117,N_18748);
nand U21379 (N_21379,N_17205,N_16726);
or U21380 (N_21380,N_18644,N_18351);
and U21381 (N_21381,N_15221,N_14033);
nor U21382 (N_21382,N_14635,N_16363);
nand U21383 (N_21383,N_13951,N_15965);
nor U21384 (N_21384,N_16394,N_15139);
and U21385 (N_21385,N_17128,N_13797);
and U21386 (N_21386,N_13137,N_18704);
nand U21387 (N_21387,N_12912,N_16607);
nand U21388 (N_21388,N_16487,N_18287);
nand U21389 (N_21389,N_18711,N_16321);
and U21390 (N_21390,N_13393,N_14986);
and U21391 (N_21391,N_14659,N_12776);
xnor U21392 (N_21392,N_14703,N_17958);
nand U21393 (N_21393,N_13369,N_17894);
nand U21394 (N_21394,N_16572,N_18118);
or U21395 (N_21395,N_15150,N_12594);
nand U21396 (N_21396,N_14260,N_15976);
or U21397 (N_21397,N_15424,N_12673);
and U21398 (N_21398,N_16079,N_14319);
nand U21399 (N_21399,N_12834,N_13546);
or U21400 (N_21400,N_17496,N_15333);
nand U21401 (N_21401,N_13725,N_14517);
nand U21402 (N_21402,N_17031,N_15682);
nor U21403 (N_21403,N_18330,N_14364);
nand U21404 (N_21404,N_18535,N_12927);
xor U21405 (N_21405,N_13470,N_14832);
nand U21406 (N_21406,N_15903,N_14024);
xor U21407 (N_21407,N_17533,N_17772);
or U21408 (N_21408,N_18673,N_16498);
or U21409 (N_21409,N_15467,N_17962);
nand U21410 (N_21410,N_13164,N_18062);
or U21411 (N_21411,N_18240,N_16409);
nor U21412 (N_21412,N_15184,N_15646);
nand U21413 (N_21413,N_17479,N_18645);
or U21414 (N_21414,N_16241,N_17139);
or U21415 (N_21415,N_16783,N_16755);
or U21416 (N_21416,N_15317,N_14629);
or U21417 (N_21417,N_16013,N_17263);
nand U21418 (N_21418,N_14505,N_15281);
nand U21419 (N_21419,N_14556,N_12688);
nor U21420 (N_21420,N_15872,N_16907);
or U21421 (N_21421,N_14968,N_12630);
nand U21422 (N_21422,N_17819,N_12821);
and U21423 (N_21423,N_17785,N_14121);
nor U21424 (N_21424,N_13805,N_12520);
nor U21425 (N_21425,N_14143,N_18444);
and U21426 (N_21426,N_16976,N_17286);
nor U21427 (N_21427,N_12643,N_15680);
xor U21428 (N_21428,N_14470,N_17561);
and U21429 (N_21429,N_18204,N_17953);
nor U21430 (N_21430,N_17660,N_16613);
and U21431 (N_21431,N_13577,N_13483);
nand U21432 (N_21432,N_12502,N_17832);
nand U21433 (N_21433,N_13220,N_18308);
and U21434 (N_21434,N_16130,N_17701);
nor U21435 (N_21435,N_12810,N_18199);
and U21436 (N_21436,N_14971,N_16180);
and U21437 (N_21437,N_14664,N_14680);
and U21438 (N_21438,N_14148,N_13189);
or U21439 (N_21439,N_18717,N_14963);
nand U21440 (N_21440,N_15964,N_18438);
and U21441 (N_21441,N_13020,N_16695);
nand U21442 (N_21442,N_16209,N_16881);
and U21443 (N_21443,N_17795,N_12627);
nand U21444 (N_21444,N_13423,N_16188);
nand U21445 (N_21445,N_17823,N_12799);
or U21446 (N_21446,N_17639,N_17428);
and U21447 (N_21447,N_17363,N_13225);
nor U21448 (N_21448,N_16596,N_16599);
and U21449 (N_21449,N_14705,N_18493);
and U21450 (N_21450,N_12987,N_17853);
and U21451 (N_21451,N_15572,N_17857);
or U21452 (N_21452,N_15552,N_17899);
nor U21453 (N_21453,N_14871,N_15253);
and U21454 (N_21454,N_17269,N_12709);
nand U21455 (N_21455,N_14295,N_12784);
and U21456 (N_21456,N_18579,N_15045);
nor U21457 (N_21457,N_12884,N_16645);
or U21458 (N_21458,N_14618,N_15215);
or U21459 (N_21459,N_16511,N_13942);
nor U21460 (N_21460,N_14391,N_15996);
xnor U21461 (N_21461,N_15319,N_17565);
nand U21462 (N_21462,N_17336,N_16118);
nand U21463 (N_21463,N_17414,N_18203);
xnor U21464 (N_21464,N_16243,N_16697);
or U21465 (N_21465,N_14129,N_18229);
nand U21466 (N_21466,N_12920,N_14258);
and U21467 (N_21467,N_17436,N_13835);
or U21468 (N_21468,N_17185,N_17727);
and U21469 (N_21469,N_17497,N_18324);
and U21470 (N_21470,N_13683,N_16974);
nand U21471 (N_21471,N_16485,N_17298);
nor U21472 (N_21472,N_18067,N_14454);
nand U21473 (N_21473,N_13372,N_17691);
or U21474 (N_21474,N_13945,N_12941);
or U21475 (N_21475,N_14079,N_12549);
nand U21476 (N_21476,N_16129,N_16114);
xnor U21477 (N_21477,N_17876,N_12836);
and U21478 (N_21478,N_13242,N_14344);
nand U21479 (N_21479,N_15100,N_15661);
nand U21480 (N_21480,N_13996,N_16255);
and U21481 (N_21481,N_15770,N_13478);
or U21482 (N_21482,N_12708,N_18744);
and U21483 (N_21483,N_12817,N_12513);
nand U21484 (N_21484,N_15428,N_16368);
and U21485 (N_21485,N_16660,N_14387);
nand U21486 (N_21486,N_17473,N_18174);
or U21487 (N_21487,N_17015,N_18137);
nand U21488 (N_21488,N_16787,N_12985);
and U21489 (N_21489,N_17991,N_12712);
nand U21490 (N_21490,N_17985,N_17224);
and U21491 (N_21491,N_18713,N_12711);
nand U21492 (N_21492,N_12890,N_14195);
and U21493 (N_21493,N_13532,N_12682);
or U21494 (N_21494,N_15886,N_16781);
or U21495 (N_21495,N_15806,N_14866);
nor U21496 (N_21496,N_18161,N_16620);
or U21497 (N_21497,N_17579,N_13594);
and U21498 (N_21498,N_18643,N_13136);
nand U21499 (N_21499,N_13537,N_16424);
nand U21500 (N_21500,N_17275,N_16486);
or U21501 (N_21501,N_17562,N_17515);
nor U21502 (N_21502,N_14808,N_18418);
or U21503 (N_21503,N_12654,N_17463);
nand U21504 (N_21504,N_17480,N_17878);
nor U21505 (N_21505,N_17534,N_17287);
xnor U21506 (N_21506,N_14191,N_17680);
nand U21507 (N_21507,N_16342,N_14421);
nor U21508 (N_21508,N_16924,N_16635);
and U21509 (N_21509,N_17431,N_15960);
and U21510 (N_21510,N_14925,N_15468);
nor U21511 (N_21511,N_15777,N_16906);
nor U21512 (N_21512,N_13684,N_13646);
nor U21513 (N_21513,N_16868,N_17914);
xnor U21514 (N_21514,N_18412,N_16340);
nand U21515 (N_21515,N_16518,N_18021);
and U21516 (N_21516,N_16460,N_15577);
or U21517 (N_21517,N_18552,N_13501);
nand U21518 (N_21518,N_17196,N_13461);
or U21519 (N_21519,N_14610,N_17898);
and U21520 (N_21520,N_15255,N_18140);
nand U21521 (N_21521,N_17856,N_13472);
or U21522 (N_21522,N_16575,N_13324);
or U21523 (N_21523,N_14164,N_15840);
xor U21524 (N_21524,N_17963,N_15077);
and U21525 (N_21525,N_14141,N_16898);
or U21526 (N_21526,N_15982,N_18183);
or U21527 (N_21527,N_18509,N_17024);
and U21528 (N_21528,N_15560,N_17904);
nand U21529 (N_21529,N_15845,N_17371);
nor U21530 (N_21530,N_14658,N_13079);
nor U21531 (N_21531,N_17141,N_16323);
nand U21532 (N_21532,N_14707,N_12530);
or U21533 (N_21533,N_18636,N_13786);
nor U21534 (N_21534,N_13368,N_16439);
nor U21535 (N_21535,N_17527,N_16570);
nand U21536 (N_21536,N_12657,N_13415);
nor U21537 (N_21537,N_13353,N_12918);
and U21538 (N_21538,N_14217,N_18688);
nor U21539 (N_21539,N_17747,N_16843);
nand U21540 (N_21540,N_13655,N_17220);
or U21541 (N_21541,N_17476,N_16553);
nor U21542 (N_21542,N_15946,N_16473);
xor U21543 (N_21543,N_17223,N_17869);
nor U21544 (N_21544,N_16987,N_14976);
or U21545 (N_21545,N_15556,N_12950);
and U21546 (N_21546,N_15443,N_14959);
nand U21547 (N_21547,N_17569,N_17825);
nand U21548 (N_21548,N_15557,N_13251);
and U21549 (N_21549,N_18267,N_12721);
xnor U21550 (N_21550,N_14071,N_16638);
and U21551 (N_21551,N_13160,N_16964);
nor U21552 (N_21552,N_17990,N_13939);
and U21553 (N_21553,N_16116,N_17180);
nand U21554 (N_21554,N_18160,N_18541);
and U21555 (N_21555,N_17008,N_18655);
nor U21556 (N_21556,N_13906,N_13224);
nor U21557 (N_21557,N_18087,N_17598);
and U21558 (N_21558,N_18040,N_13634);
and U21559 (N_21559,N_15547,N_12515);
nor U21560 (N_21560,N_16750,N_14777);
nand U21561 (N_21561,N_14104,N_14172);
nor U21562 (N_21562,N_17767,N_13371);
or U21563 (N_21563,N_15162,N_14775);
xor U21564 (N_21564,N_15084,N_16453);
or U21565 (N_21565,N_13731,N_13487);
nor U21566 (N_21566,N_15849,N_17086);
xnor U21567 (N_21567,N_13266,N_13431);
nor U21568 (N_21568,N_13860,N_18347);
nand U21569 (N_21569,N_15597,N_18152);
nor U21570 (N_21570,N_15392,N_15544);
and U21571 (N_21571,N_14686,N_14166);
nand U21572 (N_21572,N_17044,N_16862);
nand U21573 (N_21573,N_12891,N_18060);
nand U21574 (N_21574,N_15228,N_16956);
nor U21575 (N_21575,N_16160,N_16488);
or U21576 (N_21576,N_14710,N_17844);
or U21577 (N_21577,N_14145,N_13142);
or U21578 (N_21578,N_18237,N_18724);
and U21579 (N_21579,N_17956,N_17842);
nand U21580 (N_21580,N_15479,N_16948);
nand U21581 (N_21581,N_12972,N_13889);
nor U21582 (N_21582,N_14023,N_15890);
or U21583 (N_21583,N_13348,N_15940);
xnor U21584 (N_21584,N_14119,N_13171);
nand U21585 (N_21585,N_15362,N_16267);
or U21586 (N_21586,N_18014,N_16870);
nor U21587 (N_21587,N_15759,N_15354);
or U21588 (N_21588,N_16932,N_17629);
or U21589 (N_21589,N_12691,N_16158);
nor U21590 (N_21590,N_17906,N_16728);
nor U21591 (N_21591,N_13755,N_15704);
nand U21592 (N_21592,N_15233,N_13430);
nand U21593 (N_21593,N_13756,N_12686);
nand U21594 (N_21594,N_15060,N_18098);
and U21595 (N_21595,N_15141,N_17905);
nor U21596 (N_21596,N_15672,N_15088);
nor U21597 (N_21597,N_16059,N_16415);
and U21598 (N_21598,N_13936,N_16727);
and U21599 (N_21599,N_16469,N_14914);
and U21600 (N_21600,N_16083,N_13950);
or U21601 (N_21601,N_16986,N_12586);
or U21602 (N_21602,N_17741,N_17882);
and U21603 (N_21603,N_17968,N_14981);
nor U21604 (N_21604,N_16807,N_13094);
nand U21605 (N_21605,N_16472,N_18353);
and U21606 (N_21606,N_18078,N_16718);
and U21607 (N_21607,N_14809,N_18365);
nand U21608 (N_21608,N_16329,N_17945);
nor U21609 (N_21609,N_15074,N_16941);
and U21610 (N_21610,N_14855,N_16386);
or U21611 (N_21611,N_14756,N_13960);
and U21612 (N_21612,N_12976,N_12572);
nand U21613 (N_21613,N_12902,N_14783);
or U21614 (N_21614,N_15274,N_15500);
nor U21615 (N_21615,N_17307,N_17162);
nor U21616 (N_21616,N_13186,N_14381);
xor U21617 (N_21617,N_16627,N_14638);
nand U21618 (N_21618,N_18125,N_15540);
or U21619 (N_21619,N_13480,N_16984);
and U21620 (N_21620,N_14373,N_17935);
or U21621 (N_21621,N_12536,N_13909);
and U21622 (N_21622,N_16629,N_17140);
nor U21623 (N_21623,N_18610,N_15371);
nor U21624 (N_21624,N_12634,N_14920);
and U21625 (N_21625,N_17067,N_18587);
or U21626 (N_21626,N_18311,N_17395);
nor U21627 (N_21627,N_17760,N_14138);
and U21628 (N_21628,N_18670,N_13969);
nand U21629 (N_21629,N_12693,N_13859);
and U21630 (N_21630,N_12940,N_15338);
nand U21631 (N_21631,N_14753,N_14493);
or U21632 (N_21632,N_14287,N_14506);
nor U21633 (N_21633,N_15035,N_14128);
nor U21634 (N_21634,N_16671,N_16548);
and U21635 (N_21635,N_18083,N_18674);
nor U21636 (N_21636,N_16756,N_14432);
and U21637 (N_21637,N_16320,N_16032);
nor U21638 (N_21638,N_12885,N_16584);
xnor U21639 (N_21639,N_16232,N_13425);
and U21640 (N_21640,N_14839,N_18513);
nand U21641 (N_21641,N_16223,N_13742);
xor U21642 (N_21642,N_14883,N_14591);
and U21643 (N_21643,N_12614,N_13261);
or U21644 (N_21644,N_14725,N_13364);
nor U21645 (N_21645,N_17339,N_16266);
nor U21646 (N_21646,N_17855,N_13896);
or U21647 (N_21647,N_15831,N_13152);
nand U21648 (N_21648,N_13003,N_13274);
xnor U21649 (N_21649,N_14035,N_16928);
nand U21650 (N_21650,N_16774,N_17708);
and U21651 (N_21651,N_14362,N_15465);
and U21652 (N_21652,N_18120,N_16072);
and U21653 (N_21653,N_15545,N_16493);
nand U21654 (N_21654,N_12501,N_13640);
or U21655 (N_21655,N_17928,N_12955);
nand U21656 (N_21656,N_15144,N_15532);
nand U21657 (N_21657,N_14214,N_16427);
or U21658 (N_21658,N_14431,N_15923);
xor U21659 (N_21659,N_17340,N_16803);
or U21660 (N_21660,N_16788,N_15589);
nor U21661 (N_21661,N_17300,N_15639);
nor U21662 (N_21662,N_16794,N_17556);
and U21663 (N_21663,N_15079,N_15609);
or U21664 (N_21664,N_13359,N_18135);
and U21665 (N_21665,N_17632,N_13972);
or U21666 (N_21666,N_18485,N_17649);
and U21667 (N_21667,N_18632,N_13803);
nand U21668 (N_21668,N_12808,N_18111);
or U21669 (N_21669,N_17342,N_17743);
xnor U21670 (N_21670,N_16420,N_13843);
and U21671 (N_21671,N_15276,N_13328);
nand U21672 (N_21672,N_14094,N_15992);
nand U21673 (N_21673,N_15664,N_14696);
or U21674 (N_21674,N_12580,N_17068);
or U21675 (N_21675,N_14711,N_14111);
or U21676 (N_21676,N_13814,N_12977);
nor U21677 (N_21677,N_16087,N_17443);
nor U21678 (N_21678,N_12563,N_17572);
and U21679 (N_21679,N_14312,N_18212);
xor U21680 (N_21680,N_16053,N_17654);
nor U21681 (N_21681,N_15803,N_14386);
nor U21682 (N_21682,N_18187,N_14106);
and U21683 (N_21683,N_14081,N_16960);
xnor U21684 (N_21684,N_14931,N_14609);
and U21685 (N_21685,N_15225,N_18053);
and U21686 (N_21686,N_13530,N_14789);
or U21687 (N_21687,N_13058,N_16125);
and U21688 (N_21688,N_16951,N_13839);
xnor U21689 (N_21689,N_16585,N_17647);
and U21690 (N_21690,N_14766,N_15091);
nor U21691 (N_21691,N_13536,N_15167);
xnor U21692 (N_21692,N_13946,N_15583);
or U21693 (N_21693,N_17281,N_15760);
nand U21694 (N_21694,N_15520,N_16639);
nand U21695 (N_21695,N_16245,N_13559);
nand U21696 (N_21696,N_12874,N_15022);
nor U21697 (N_21697,N_13792,N_15739);
nor U21698 (N_21698,N_14348,N_16113);
nor U21699 (N_21699,N_15456,N_15263);
nor U21700 (N_21700,N_18333,N_17801);
nand U21701 (N_21701,N_17125,N_17505);
or U21702 (N_21702,N_17942,N_14003);
nor U21703 (N_21703,N_17927,N_16714);
nor U21704 (N_21704,N_17887,N_14677);
nor U21705 (N_21705,N_14632,N_13697);
nor U21706 (N_21706,N_16985,N_14017);
nor U21707 (N_21707,N_16138,N_16943);
nand U21708 (N_21708,N_16430,N_14426);
nor U21709 (N_21709,N_18262,N_14398);
or U21710 (N_21710,N_15197,N_15410);
nand U21711 (N_21711,N_17809,N_14768);
nand U21712 (N_21712,N_16798,N_15691);
and U21713 (N_21713,N_12769,N_12662);
and U21714 (N_21714,N_17100,N_12951);
nand U21715 (N_21715,N_18359,N_15416);
nor U21716 (N_21716,N_13205,N_17787);
nor U21717 (N_21717,N_16665,N_17227);
nand U21718 (N_21718,N_17495,N_17487);
and U21719 (N_21719,N_17493,N_18666);
and U21720 (N_21720,N_16191,N_13114);
and U21721 (N_21721,N_14423,N_16039);
or U21722 (N_21722,N_15094,N_12546);
nor U21723 (N_21723,N_18110,N_13289);
nand U21724 (N_21724,N_14018,N_14056);
nor U21725 (N_21725,N_16449,N_14158);
and U21726 (N_21726,N_15731,N_12622);
or U21727 (N_21727,N_18470,N_13672);
or U21728 (N_21728,N_14627,N_13615);
xnor U21729 (N_21729,N_16082,N_13595);
or U21730 (N_21730,N_13645,N_14082);
or U21731 (N_21731,N_13245,N_15644);
nor U21732 (N_21732,N_14355,N_14619);
and U21733 (N_21733,N_14604,N_12642);
or U21734 (N_21734,N_13761,N_18058);
and U21735 (N_21735,N_15053,N_16148);
nand U21736 (N_21736,N_12803,N_15942);
and U21737 (N_21737,N_16865,N_15057);
nand U21738 (N_21738,N_14945,N_12949);
nor U21739 (N_21739,N_16670,N_15358);
and U21740 (N_21740,N_13727,N_13158);
nand U21741 (N_21741,N_14882,N_17007);
or U21742 (N_21742,N_13247,N_15912);
nor U21743 (N_21743,N_16244,N_12500);
nor U21744 (N_21744,N_13183,N_18627);
or U21745 (N_21745,N_14435,N_13297);
or U21746 (N_21746,N_13270,N_13493);
or U21747 (N_21747,N_12632,N_14870);
or U21748 (N_21748,N_13555,N_15087);
nand U21749 (N_21749,N_15689,N_18465);
nor U21750 (N_21750,N_13934,N_18258);
nor U21751 (N_21751,N_16364,N_15823);
nand U21752 (N_21752,N_18321,N_17435);
xor U21753 (N_21753,N_18081,N_14695);
or U21754 (N_21754,N_13877,N_16692);
and U21755 (N_21755,N_15143,N_17129);
or U21756 (N_21756,N_15061,N_15530);
nor U21757 (N_21757,N_15011,N_16954);
nor U21758 (N_21758,N_16730,N_18143);
nand U21759 (N_21759,N_15374,N_13481);
xor U21760 (N_21760,N_17580,N_18414);
nand U21761 (N_21761,N_13516,N_14463);
nor U21762 (N_21762,N_12969,N_17283);
and U21763 (N_21763,N_16646,N_18027);
nor U21764 (N_21764,N_18698,N_13890);
nor U21765 (N_21765,N_15618,N_14224);
and U21766 (N_21766,N_14242,N_13489);
nor U21767 (N_21767,N_12980,N_16833);
and U21768 (N_21768,N_13217,N_16356);
nand U21769 (N_21769,N_17571,N_17883);
or U21770 (N_21770,N_14027,N_12722);
or U21771 (N_21771,N_17225,N_13654);
or U21772 (N_21772,N_15123,N_14247);
nand U21773 (N_21773,N_14708,N_18057);
or U21774 (N_21774,N_17615,N_15009);
and U21775 (N_21775,N_18361,N_16925);
xnor U21776 (N_21776,N_15962,N_15076);
xor U21777 (N_21777,N_14494,N_15869);
or U21778 (N_21778,N_16350,N_13774);
nor U21779 (N_21779,N_15356,N_13662);
nand U21780 (N_21780,N_15407,N_12868);
or U21781 (N_21781,N_15301,N_17936);
or U21782 (N_21782,N_13426,N_17047);
nor U21783 (N_21783,N_17438,N_14562);
and U21784 (N_21784,N_17925,N_18323);
nand U21785 (N_21785,N_12899,N_18259);
or U21786 (N_21786,N_17596,N_13024);
nand U21787 (N_21787,N_13617,N_13998);
and U21788 (N_21788,N_15879,N_17650);
and U21789 (N_21789,N_18121,N_12991);
or U21790 (N_21790,N_18524,N_18691);
nor U21791 (N_21791,N_18011,N_17738);
xor U21792 (N_21792,N_15816,N_16346);
and U21793 (N_21793,N_13062,N_12768);
nor U21794 (N_21794,N_14742,N_17502);
and U21795 (N_21795,N_17602,N_17830);
nor U21796 (N_21796,N_17663,N_15408);
and U21797 (N_21797,N_14751,N_13916);
or U21798 (N_21798,N_13984,N_14060);
or U21799 (N_21799,N_15275,N_14748);
nor U21800 (N_21800,N_13676,N_17840);
and U21801 (N_21801,N_15810,N_15393);
nand U21802 (N_21802,N_16526,N_17531);
and U21803 (N_21803,N_17131,N_13891);
nor U21804 (N_21804,N_14439,N_16095);
nor U21805 (N_21805,N_13750,N_17005);
or U21806 (N_21806,N_15488,N_13768);
and U21807 (N_21807,N_14123,N_13571);
nor U21808 (N_21808,N_14353,N_18648);
nor U21809 (N_21809,N_17920,N_16290);
nand U21810 (N_21810,N_14394,N_13255);
xor U21811 (N_21811,N_17467,N_12849);
and U21812 (N_21812,N_14178,N_15107);
and U21813 (N_21813,N_12535,N_13409);
and U21814 (N_21814,N_16912,N_13135);
nand U21815 (N_21815,N_14047,N_18680);
nor U21816 (N_21816,N_16416,N_14052);
and U21817 (N_21817,N_17331,N_13710);
xnor U21818 (N_21818,N_12678,N_12741);
xor U21819 (N_21819,N_17924,N_15674);
or U21820 (N_21820,N_17444,N_17860);
or U21821 (N_21821,N_18089,N_12751);
and U21822 (N_21822,N_14917,N_15216);
and U21823 (N_21823,N_16589,N_15728);
nor U21824 (N_21824,N_15856,N_17525);
and U21825 (N_21825,N_12603,N_17568);
nand U21826 (N_21826,N_17134,N_14370);
and U21827 (N_21827,N_13737,N_14887);
nand U21828 (N_21828,N_15843,N_14654);
or U21829 (N_21829,N_15859,N_15334);
nor U21830 (N_21830,N_15772,N_13551);
and U21831 (N_21831,N_17547,N_17277);
or U21832 (N_21832,N_14739,N_12592);
or U21833 (N_21833,N_13473,N_18511);
or U21834 (N_21834,N_15095,N_15647);
nand U21835 (N_21835,N_15007,N_16770);
nor U21836 (N_21836,N_14271,N_15381);
or U21837 (N_21837,N_15943,N_13156);
nand U21838 (N_21838,N_17491,N_18449);
and U21839 (N_21839,N_17429,N_14863);
or U21840 (N_21840,N_12746,N_16564);
or U21841 (N_21841,N_17142,N_18494);
nand U21842 (N_21842,N_15200,N_15771);
nor U21843 (N_21843,N_12801,N_14667);
and U21844 (N_21844,N_15975,N_17641);
or U21845 (N_21845,N_13334,N_13736);
and U21846 (N_21846,N_14046,N_16176);
and U21847 (N_21847,N_18252,N_16281);
or U21848 (N_21848,N_17374,N_18165);
nor U21849 (N_21849,N_15118,N_15436);
and U21850 (N_21850,N_18551,N_16940);
xor U21851 (N_21851,N_15534,N_15005);
and U21852 (N_21852,N_15003,N_15905);
nand U21853 (N_21853,N_13072,N_16992);
and U21854 (N_21854,N_16641,N_16301);
and U21855 (N_21855,N_14157,N_14993);
nor U21856 (N_21856,N_18086,N_13704);
nor U21857 (N_21857,N_17171,N_13193);
nand U21858 (N_21858,N_13315,N_13545);
nand U21859 (N_21859,N_13573,N_13086);
and U21860 (N_21860,N_12843,N_16322);
and U21861 (N_21861,N_16417,N_15695);
nor U21862 (N_21862,N_18222,N_18133);
nand U21863 (N_21863,N_18441,N_16274);
nor U21864 (N_21864,N_16901,N_15875);
xor U21865 (N_21865,N_13280,N_17636);
and U21866 (N_21866,N_17231,N_17589);
xnor U21867 (N_21867,N_15719,N_16977);
and U21868 (N_21868,N_18176,N_13243);
and U21869 (N_21869,N_15658,N_14857);
nor U21870 (N_21870,N_18338,N_14294);
xnor U21871 (N_21871,N_14330,N_14858);
nand U21872 (N_21872,N_13920,N_15623);
and U21873 (N_21873,N_16131,N_15722);
xnor U21874 (N_21874,N_17038,N_17357);
nand U21875 (N_21875,N_15150,N_18747);
or U21876 (N_21876,N_15680,N_14744);
nand U21877 (N_21877,N_18730,N_15502);
nor U21878 (N_21878,N_14462,N_12827);
or U21879 (N_21879,N_18197,N_16761);
or U21880 (N_21880,N_16563,N_16878);
or U21881 (N_21881,N_15245,N_18598);
or U21882 (N_21882,N_16369,N_17862);
nor U21883 (N_21883,N_12865,N_15854);
nor U21884 (N_21884,N_18448,N_12665);
xnor U21885 (N_21885,N_14310,N_15398);
or U21886 (N_21886,N_12675,N_15849);
nand U21887 (N_21887,N_18663,N_17936);
nand U21888 (N_21888,N_15040,N_16402);
and U21889 (N_21889,N_17801,N_18735);
nand U21890 (N_21890,N_12703,N_14601);
and U21891 (N_21891,N_17594,N_13857);
nand U21892 (N_21892,N_14436,N_14130);
or U21893 (N_21893,N_16228,N_12644);
or U21894 (N_21894,N_18664,N_14127);
nor U21895 (N_21895,N_13972,N_18256);
nand U21896 (N_21896,N_18252,N_16596);
or U21897 (N_21897,N_13542,N_13227);
xor U21898 (N_21898,N_18530,N_16172);
or U21899 (N_21899,N_14173,N_12914);
and U21900 (N_21900,N_13452,N_18371);
xor U21901 (N_21901,N_17718,N_15132);
nand U21902 (N_21902,N_13413,N_14357);
and U21903 (N_21903,N_12789,N_14169);
and U21904 (N_21904,N_14070,N_14580);
and U21905 (N_21905,N_18252,N_16068);
xnor U21906 (N_21906,N_14801,N_13488);
or U21907 (N_21907,N_13860,N_13939);
xnor U21908 (N_21908,N_13838,N_13208);
nand U21909 (N_21909,N_17926,N_16813);
nand U21910 (N_21910,N_12687,N_18404);
nor U21911 (N_21911,N_14040,N_15307);
nand U21912 (N_21912,N_13473,N_14697);
nor U21913 (N_21913,N_13109,N_17825);
or U21914 (N_21914,N_14742,N_14113);
nor U21915 (N_21915,N_17451,N_14536);
nand U21916 (N_21916,N_17705,N_16562);
or U21917 (N_21917,N_14946,N_16670);
and U21918 (N_21918,N_15857,N_15044);
or U21919 (N_21919,N_16351,N_13530);
and U21920 (N_21920,N_13512,N_17338);
and U21921 (N_21921,N_17491,N_18054);
nor U21922 (N_21922,N_12745,N_16772);
nor U21923 (N_21923,N_13710,N_16430);
or U21924 (N_21924,N_12983,N_13630);
nor U21925 (N_21925,N_16249,N_13148);
nor U21926 (N_21926,N_17002,N_16290);
or U21927 (N_21927,N_17337,N_12917);
nand U21928 (N_21928,N_12772,N_13595);
nand U21929 (N_21929,N_15812,N_13910);
or U21930 (N_21930,N_13928,N_14702);
and U21931 (N_21931,N_15267,N_15328);
nor U21932 (N_21932,N_16683,N_12757);
and U21933 (N_21933,N_18327,N_17625);
nor U21934 (N_21934,N_13388,N_18111);
nand U21935 (N_21935,N_13439,N_18278);
nor U21936 (N_21936,N_12626,N_14606);
nand U21937 (N_21937,N_15292,N_15369);
and U21938 (N_21938,N_13335,N_15992);
and U21939 (N_21939,N_12525,N_16654);
or U21940 (N_21940,N_13350,N_16635);
and U21941 (N_21941,N_12598,N_14766);
nor U21942 (N_21942,N_14233,N_12525);
nor U21943 (N_21943,N_12740,N_17477);
nor U21944 (N_21944,N_18305,N_14566);
nor U21945 (N_21945,N_15975,N_14696);
nand U21946 (N_21946,N_12848,N_15972);
and U21947 (N_21947,N_12608,N_15293);
and U21948 (N_21948,N_15232,N_14353);
nand U21949 (N_21949,N_14084,N_16276);
nor U21950 (N_21950,N_17465,N_15863);
or U21951 (N_21951,N_14051,N_13950);
nand U21952 (N_21952,N_16608,N_17955);
nand U21953 (N_21953,N_13176,N_16449);
and U21954 (N_21954,N_13838,N_18746);
nor U21955 (N_21955,N_13578,N_13655);
and U21956 (N_21956,N_13470,N_15608);
nor U21957 (N_21957,N_15886,N_14399);
or U21958 (N_21958,N_16251,N_18133);
and U21959 (N_21959,N_16872,N_16892);
or U21960 (N_21960,N_13391,N_16232);
xnor U21961 (N_21961,N_13698,N_13085);
and U21962 (N_21962,N_17043,N_17965);
xor U21963 (N_21963,N_14054,N_17676);
nand U21964 (N_21964,N_15685,N_13021);
nor U21965 (N_21965,N_17949,N_17385);
or U21966 (N_21966,N_16636,N_14984);
and U21967 (N_21967,N_15572,N_15987);
and U21968 (N_21968,N_17524,N_12715);
and U21969 (N_21969,N_13615,N_15297);
or U21970 (N_21970,N_14473,N_13750);
or U21971 (N_21971,N_18687,N_14750);
nand U21972 (N_21972,N_14439,N_15182);
or U21973 (N_21973,N_14767,N_18371);
or U21974 (N_21974,N_17454,N_13561);
or U21975 (N_21975,N_13899,N_16848);
nand U21976 (N_21976,N_12749,N_18172);
and U21977 (N_21977,N_13206,N_13941);
nor U21978 (N_21978,N_14881,N_18515);
or U21979 (N_21979,N_13476,N_13149);
and U21980 (N_21980,N_15338,N_15518);
and U21981 (N_21981,N_16605,N_13290);
nand U21982 (N_21982,N_13447,N_16250);
and U21983 (N_21983,N_18139,N_13289);
or U21984 (N_21984,N_13930,N_12604);
and U21985 (N_21985,N_13932,N_13466);
and U21986 (N_21986,N_16383,N_14396);
and U21987 (N_21987,N_17482,N_14276);
and U21988 (N_21988,N_15588,N_17921);
xnor U21989 (N_21989,N_12996,N_13840);
nand U21990 (N_21990,N_16378,N_18208);
nor U21991 (N_21991,N_17700,N_14916);
or U21992 (N_21992,N_18600,N_18091);
nand U21993 (N_21993,N_14119,N_14142);
nor U21994 (N_21994,N_15730,N_14361);
nand U21995 (N_21995,N_14759,N_16788);
or U21996 (N_21996,N_18498,N_18733);
or U21997 (N_21997,N_17568,N_18671);
or U21998 (N_21998,N_16179,N_14034);
and U21999 (N_21999,N_13834,N_15706);
nor U22000 (N_22000,N_17904,N_15681);
nand U22001 (N_22001,N_15070,N_12552);
and U22002 (N_22002,N_15533,N_16710);
or U22003 (N_22003,N_18658,N_17270);
or U22004 (N_22004,N_13393,N_13135);
nor U22005 (N_22005,N_15091,N_17642);
nand U22006 (N_22006,N_13685,N_16874);
or U22007 (N_22007,N_15476,N_18513);
nand U22008 (N_22008,N_14783,N_15236);
or U22009 (N_22009,N_15347,N_13450);
nand U22010 (N_22010,N_18418,N_13658);
and U22011 (N_22011,N_13778,N_14431);
nand U22012 (N_22012,N_12686,N_17885);
or U22013 (N_22013,N_15095,N_17501);
nor U22014 (N_22014,N_15477,N_14344);
or U22015 (N_22015,N_17617,N_14154);
or U22016 (N_22016,N_15547,N_14806);
or U22017 (N_22017,N_12786,N_14075);
nor U22018 (N_22018,N_13830,N_14871);
nor U22019 (N_22019,N_17653,N_13206);
and U22020 (N_22020,N_14415,N_12772);
xnor U22021 (N_22021,N_14527,N_17627);
or U22022 (N_22022,N_13425,N_17752);
nand U22023 (N_22023,N_15807,N_12721);
or U22024 (N_22024,N_18188,N_15941);
xor U22025 (N_22025,N_13692,N_15286);
nor U22026 (N_22026,N_16131,N_13612);
xor U22027 (N_22027,N_12897,N_16335);
and U22028 (N_22028,N_12938,N_16790);
xnor U22029 (N_22029,N_16878,N_18598);
nor U22030 (N_22030,N_14427,N_14032);
nor U22031 (N_22031,N_15609,N_15026);
nor U22032 (N_22032,N_18138,N_12750);
nand U22033 (N_22033,N_18053,N_14243);
nand U22034 (N_22034,N_14999,N_13734);
or U22035 (N_22035,N_16177,N_15857);
nand U22036 (N_22036,N_14835,N_16432);
and U22037 (N_22037,N_15826,N_14261);
nand U22038 (N_22038,N_17750,N_14419);
nand U22039 (N_22039,N_13713,N_13409);
xor U22040 (N_22040,N_17803,N_17250);
or U22041 (N_22041,N_17478,N_18272);
nand U22042 (N_22042,N_16504,N_14125);
nor U22043 (N_22043,N_18730,N_14475);
and U22044 (N_22044,N_14084,N_13477);
nor U22045 (N_22045,N_16833,N_15223);
nand U22046 (N_22046,N_16745,N_16328);
or U22047 (N_22047,N_16064,N_14672);
xor U22048 (N_22048,N_14986,N_18639);
nand U22049 (N_22049,N_13111,N_14690);
or U22050 (N_22050,N_13160,N_17977);
nand U22051 (N_22051,N_12992,N_14010);
nor U22052 (N_22052,N_14679,N_14965);
or U22053 (N_22053,N_14500,N_16915);
or U22054 (N_22054,N_13648,N_18383);
nand U22055 (N_22055,N_18745,N_14235);
xor U22056 (N_22056,N_18591,N_13707);
and U22057 (N_22057,N_12841,N_15845);
or U22058 (N_22058,N_15361,N_17470);
xnor U22059 (N_22059,N_17467,N_13811);
nor U22060 (N_22060,N_14981,N_13275);
nor U22061 (N_22061,N_13683,N_13443);
and U22062 (N_22062,N_14135,N_16982);
nand U22063 (N_22063,N_15545,N_13239);
xnor U22064 (N_22064,N_15206,N_18509);
nor U22065 (N_22065,N_12568,N_16113);
nand U22066 (N_22066,N_13446,N_13506);
and U22067 (N_22067,N_14533,N_17585);
nor U22068 (N_22068,N_13899,N_12885);
or U22069 (N_22069,N_17113,N_18375);
nor U22070 (N_22070,N_18150,N_12620);
or U22071 (N_22071,N_18167,N_18402);
or U22072 (N_22072,N_15296,N_13642);
or U22073 (N_22073,N_17170,N_15858);
and U22074 (N_22074,N_15662,N_13839);
nand U22075 (N_22075,N_14445,N_17853);
and U22076 (N_22076,N_16605,N_18594);
or U22077 (N_22077,N_18478,N_18433);
and U22078 (N_22078,N_15064,N_16456);
nor U22079 (N_22079,N_13106,N_16729);
nand U22080 (N_22080,N_17992,N_17567);
nand U22081 (N_22081,N_17212,N_14784);
or U22082 (N_22082,N_13831,N_14374);
and U22083 (N_22083,N_13151,N_12831);
nand U22084 (N_22084,N_12661,N_15447);
or U22085 (N_22085,N_15193,N_16690);
xnor U22086 (N_22086,N_15832,N_14155);
nand U22087 (N_22087,N_13136,N_13011);
xor U22088 (N_22088,N_13969,N_17992);
or U22089 (N_22089,N_13820,N_17780);
or U22090 (N_22090,N_14307,N_18230);
nand U22091 (N_22091,N_15966,N_14938);
nor U22092 (N_22092,N_12846,N_16146);
nor U22093 (N_22093,N_17984,N_13831);
and U22094 (N_22094,N_14766,N_15108);
and U22095 (N_22095,N_14405,N_14479);
nand U22096 (N_22096,N_14081,N_16088);
or U22097 (N_22097,N_15343,N_17647);
nand U22098 (N_22098,N_14586,N_13771);
nand U22099 (N_22099,N_13717,N_16884);
nor U22100 (N_22100,N_13798,N_15374);
and U22101 (N_22101,N_13319,N_18646);
nor U22102 (N_22102,N_15589,N_13836);
nand U22103 (N_22103,N_15291,N_17419);
nand U22104 (N_22104,N_13548,N_15297);
nand U22105 (N_22105,N_17807,N_15494);
or U22106 (N_22106,N_14901,N_13152);
nor U22107 (N_22107,N_14275,N_14511);
nor U22108 (N_22108,N_12738,N_17705);
or U22109 (N_22109,N_17040,N_17767);
nand U22110 (N_22110,N_14807,N_15076);
or U22111 (N_22111,N_15566,N_14385);
nand U22112 (N_22112,N_17581,N_12990);
and U22113 (N_22113,N_15781,N_14300);
nor U22114 (N_22114,N_12882,N_17879);
or U22115 (N_22115,N_17533,N_14826);
and U22116 (N_22116,N_12961,N_16873);
and U22117 (N_22117,N_15487,N_15006);
or U22118 (N_22118,N_12861,N_13261);
nand U22119 (N_22119,N_12588,N_14169);
nand U22120 (N_22120,N_17992,N_18067);
xnor U22121 (N_22121,N_16219,N_15393);
or U22122 (N_22122,N_15973,N_13212);
and U22123 (N_22123,N_16404,N_13812);
nor U22124 (N_22124,N_15668,N_15111);
nand U22125 (N_22125,N_18503,N_17054);
nor U22126 (N_22126,N_14101,N_16618);
and U22127 (N_22127,N_16635,N_14169);
nor U22128 (N_22128,N_14574,N_12801);
nand U22129 (N_22129,N_16565,N_12877);
nor U22130 (N_22130,N_16627,N_14170);
nor U22131 (N_22131,N_17957,N_17324);
nor U22132 (N_22132,N_14320,N_17083);
nand U22133 (N_22133,N_17314,N_18085);
nand U22134 (N_22134,N_16444,N_13722);
and U22135 (N_22135,N_17643,N_16176);
nand U22136 (N_22136,N_16791,N_15104);
nor U22137 (N_22137,N_13309,N_18213);
nand U22138 (N_22138,N_12734,N_16144);
nor U22139 (N_22139,N_14748,N_15892);
nand U22140 (N_22140,N_12885,N_16637);
or U22141 (N_22141,N_13955,N_15506);
or U22142 (N_22142,N_16922,N_15368);
and U22143 (N_22143,N_13670,N_18217);
nor U22144 (N_22144,N_18546,N_15365);
nand U22145 (N_22145,N_17133,N_18251);
nor U22146 (N_22146,N_15474,N_13013);
nor U22147 (N_22147,N_17919,N_14575);
or U22148 (N_22148,N_17006,N_14872);
xor U22149 (N_22149,N_13201,N_17660);
and U22150 (N_22150,N_17914,N_16259);
or U22151 (N_22151,N_13583,N_13374);
nand U22152 (N_22152,N_18722,N_13871);
and U22153 (N_22153,N_12927,N_17444);
nand U22154 (N_22154,N_13584,N_14478);
and U22155 (N_22155,N_16614,N_17153);
and U22156 (N_22156,N_18095,N_16123);
or U22157 (N_22157,N_18484,N_14508);
and U22158 (N_22158,N_16388,N_14005);
xor U22159 (N_22159,N_14535,N_18492);
nor U22160 (N_22160,N_16299,N_14426);
nor U22161 (N_22161,N_15291,N_16668);
or U22162 (N_22162,N_15933,N_16447);
or U22163 (N_22163,N_14293,N_15893);
nand U22164 (N_22164,N_13866,N_18151);
or U22165 (N_22165,N_16279,N_18273);
or U22166 (N_22166,N_17424,N_12553);
and U22167 (N_22167,N_14521,N_17482);
or U22168 (N_22168,N_17163,N_13678);
and U22169 (N_22169,N_17054,N_18021);
nand U22170 (N_22170,N_14416,N_17338);
nor U22171 (N_22171,N_15973,N_12662);
and U22172 (N_22172,N_15438,N_14554);
and U22173 (N_22173,N_16383,N_16938);
and U22174 (N_22174,N_18397,N_14207);
and U22175 (N_22175,N_14560,N_13204);
nor U22176 (N_22176,N_15646,N_15121);
or U22177 (N_22177,N_17348,N_15899);
nand U22178 (N_22178,N_16031,N_16186);
and U22179 (N_22179,N_13600,N_14619);
nand U22180 (N_22180,N_13542,N_12661);
nand U22181 (N_22181,N_14327,N_13874);
nor U22182 (N_22182,N_13534,N_16872);
and U22183 (N_22183,N_12636,N_15597);
and U22184 (N_22184,N_14035,N_15581);
xnor U22185 (N_22185,N_16712,N_15123);
nand U22186 (N_22186,N_13110,N_12555);
and U22187 (N_22187,N_18311,N_16584);
or U22188 (N_22188,N_18436,N_14255);
xor U22189 (N_22189,N_13705,N_16266);
and U22190 (N_22190,N_16961,N_16768);
nor U22191 (N_22191,N_18120,N_15930);
and U22192 (N_22192,N_16905,N_15872);
nor U22193 (N_22193,N_16763,N_15528);
nand U22194 (N_22194,N_13374,N_12687);
and U22195 (N_22195,N_14841,N_12907);
or U22196 (N_22196,N_17178,N_18200);
nor U22197 (N_22197,N_14784,N_15169);
nand U22198 (N_22198,N_18252,N_18151);
xor U22199 (N_22199,N_14301,N_17962);
nor U22200 (N_22200,N_14295,N_12841);
nor U22201 (N_22201,N_14243,N_15449);
and U22202 (N_22202,N_15894,N_16687);
and U22203 (N_22203,N_12700,N_18156);
and U22204 (N_22204,N_18684,N_13521);
nor U22205 (N_22205,N_17418,N_14756);
or U22206 (N_22206,N_18738,N_16588);
nor U22207 (N_22207,N_17895,N_15128);
or U22208 (N_22208,N_17548,N_14609);
and U22209 (N_22209,N_16779,N_18041);
or U22210 (N_22210,N_15180,N_12535);
and U22211 (N_22211,N_16601,N_15444);
or U22212 (N_22212,N_16405,N_15692);
nand U22213 (N_22213,N_16750,N_15033);
or U22214 (N_22214,N_12750,N_16043);
nand U22215 (N_22215,N_14629,N_15110);
xor U22216 (N_22216,N_18176,N_15590);
and U22217 (N_22217,N_16651,N_13186);
and U22218 (N_22218,N_13597,N_15474);
or U22219 (N_22219,N_13213,N_14030);
and U22220 (N_22220,N_13256,N_18048);
and U22221 (N_22221,N_18338,N_14298);
xor U22222 (N_22222,N_13031,N_13738);
nand U22223 (N_22223,N_13432,N_18432);
nor U22224 (N_22224,N_17305,N_14034);
or U22225 (N_22225,N_17639,N_16909);
nand U22226 (N_22226,N_15870,N_17126);
nand U22227 (N_22227,N_16230,N_15479);
xor U22228 (N_22228,N_16936,N_16340);
nor U22229 (N_22229,N_15966,N_17280);
nand U22230 (N_22230,N_15942,N_17612);
nor U22231 (N_22231,N_16736,N_13146);
nor U22232 (N_22232,N_17837,N_13724);
nor U22233 (N_22233,N_12673,N_13847);
nand U22234 (N_22234,N_18420,N_15819);
nand U22235 (N_22235,N_13704,N_15303);
and U22236 (N_22236,N_14344,N_18595);
and U22237 (N_22237,N_17312,N_16847);
or U22238 (N_22238,N_16593,N_14758);
nand U22239 (N_22239,N_14968,N_12932);
and U22240 (N_22240,N_16550,N_12882);
xor U22241 (N_22241,N_18069,N_13183);
and U22242 (N_22242,N_12792,N_18744);
nand U22243 (N_22243,N_15257,N_15301);
nand U22244 (N_22244,N_13685,N_14164);
nor U22245 (N_22245,N_15463,N_14756);
nand U22246 (N_22246,N_12777,N_12785);
nand U22247 (N_22247,N_12578,N_17451);
or U22248 (N_22248,N_18455,N_16935);
and U22249 (N_22249,N_18678,N_13858);
or U22250 (N_22250,N_18671,N_12770);
nor U22251 (N_22251,N_16514,N_17889);
nor U22252 (N_22252,N_14587,N_16498);
xnor U22253 (N_22253,N_16071,N_16185);
nand U22254 (N_22254,N_14784,N_16271);
nor U22255 (N_22255,N_15386,N_14777);
nor U22256 (N_22256,N_14852,N_18112);
and U22257 (N_22257,N_13393,N_17541);
nand U22258 (N_22258,N_14321,N_18213);
xor U22259 (N_22259,N_17817,N_17548);
and U22260 (N_22260,N_13437,N_14514);
or U22261 (N_22261,N_16646,N_13733);
nand U22262 (N_22262,N_14886,N_15581);
nor U22263 (N_22263,N_16119,N_15163);
nand U22264 (N_22264,N_14751,N_17388);
and U22265 (N_22265,N_15716,N_14597);
and U22266 (N_22266,N_17177,N_16253);
nor U22267 (N_22267,N_17019,N_17584);
nor U22268 (N_22268,N_12886,N_13193);
and U22269 (N_22269,N_15883,N_13586);
nand U22270 (N_22270,N_13574,N_15398);
or U22271 (N_22271,N_17938,N_16123);
nand U22272 (N_22272,N_15633,N_17076);
nor U22273 (N_22273,N_17096,N_16695);
nor U22274 (N_22274,N_17646,N_12739);
or U22275 (N_22275,N_17264,N_13295);
nand U22276 (N_22276,N_14419,N_17803);
and U22277 (N_22277,N_16495,N_15102);
nand U22278 (N_22278,N_13558,N_15624);
xnor U22279 (N_22279,N_13056,N_15087);
nor U22280 (N_22280,N_15270,N_18545);
nand U22281 (N_22281,N_18160,N_13723);
nand U22282 (N_22282,N_12646,N_14742);
nand U22283 (N_22283,N_14587,N_17956);
and U22284 (N_22284,N_12571,N_16754);
nor U22285 (N_22285,N_16679,N_17313);
and U22286 (N_22286,N_13860,N_18608);
nor U22287 (N_22287,N_15285,N_13693);
and U22288 (N_22288,N_12724,N_16222);
nand U22289 (N_22289,N_16281,N_14220);
or U22290 (N_22290,N_15224,N_14942);
nand U22291 (N_22291,N_16089,N_13584);
and U22292 (N_22292,N_13991,N_14792);
nor U22293 (N_22293,N_14159,N_18022);
nand U22294 (N_22294,N_17638,N_14054);
and U22295 (N_22295,N_18257,N_14546);
or U22296 (N_22296,N_16191,N_12844);
nand U22297 (N_22297,N_17360,N_15672);
or U22298 (N_22298,N_16356,N_12714);
nand U22299 (N_22299,N_14351,N_14896);
or U22300 (N_22300,N_14618,N_15379);
nand U22301 (N_22301,N_13992,N_12574);
or U22302 (N_22302,N_18086,N_12828);
or U22303 (N_22303,N_13687,N_14767);
or U22304 (N_22304,N_13719,N_18628);
nor U22305 (N_22305,N_16196,N_15949);
nand U22306 (N_22306,N_14903,N_13254);
nand U22307 (N_22307,N_17519,N_13824);
or U22308 (N_22308,N_15442,N_18136);
nor U22309 (N_22309,N_17984,N_14129);
and U22310 (N_22310,N_14392,N_14843);
nand U22311 (N_22311,N_13616,N_17984);
and U22312 (N_22312,N_18177,N_18355);
xnor U22313 (N_22313,N_16169,N_16544);
and U22314 (N_22314,N_18305,N_17096);
nand U22315 (N_22315,N_13767,N_14572);
or U22316 (N_22316,N_13814,N_14838);
xnor U22317 (N_22317,N_16339,N_16623);
nor U22318 (N_22318,N_13313,N_16481);
nand U22319 (N_22319,N_17812,N_14927);
nand U22320 (N_22320,N_13397,N_17619);
nor U22321 (N_22321,N_16371,N_15135);
or U22322 (N_22322,N_13172,N_12719);
nor U22323 (N_22323,N_13260,N_13511);
nand U22324 (N_22324,N_13874,N_16105);
and U22325 (N_22325,N_12596,N_13072);
and U22326 (N_22326,N_12810,N_17855);
xor U22327 (N_22327,N_18740,N_15390);
nand U22328 (N_22328,N_13176,N_16206);
xor U22329 (N_22329,N_12661,N_17210);
and U22330 (N_22330,N_12673,N_16636);
nor U22331 (N_22331,N_17837,N_14636);
nor U22332 (N_22332,N_16498,N_13128);
nor U22333 (N_22333,N_14708,N_16973);
nor U22334 (N_22334,N_16513,N_17268);
or U22335 (N_22335,N_18374,N_16142);
nor U22336 (N_22336,N_14907,N_13188);
and U22337 (N_22337,N_14522,N_14268);
nand U22338 (N_22338,N_15007,N_15190);
nor U22339 (N_22339,N_12863,N_12532);
nand U22340 (N_22340,N_15619,N_14993);
nand U22341 (N_22341,N_16148,N_18480);
xnor U22342 (N_22342,N_13472,N_16463);
nand U22343 (N_22343,N_15715,N_16434);
and U22344 (N_22344,N_13412,N_16547);
or U22345 (N_22345,N_14222,N_13529);
and U22346 (N_22346,N_15198,N_17379);
nand U22347 (N_22347,N_16788,N_17376);
nand U22348 (N_22348,N_17593,N_12842);
or U22349 (N_22349,N_17141,N_13269);
xor U22350 (N_22350,N_12863,N_13823);
nand U22351 (N_22351,N_15238,N_18727);
and U22352 (N_22352,N_13075,N_18353);
nand U22353 (N_22353,N_16577,N_15664);
or U22354 (N_22354,N_13572,N_15469);
or U22355 (N_22355,N_13792,N_14452);
and U22356 (N_22356,N_17682,N_12530);
and U22357 (N_22357,N_17476,N_17389);
or U22358 (N_22358,N_14079,N_17680);
and U22359 (N_22359,N_14682,N_14914);
and U22360 (N_22360,N_15516,N_18040);
and U22361 (N_22361,N_14492,N_16143);
nor U22362 (N_22362,N_14985,N_14683);
or U22363 (N_22363,N_16447,N_16315);
and U22364 (N_22364,N_17422,N_16016);
and U22365 (N_22365,N_13833,N_12631);
and U22366 (N_22366,N_14852,N_17895);
and U22367 (N_22367,N_13402,N_14426);
or U22368 (N_22368,N_15513,N_17178);
nor U22369 (N_22369,N_18732,N_16861);
nor U22370 (N_22370,N_17036,N_15497);
nand U22371 (N_22371,N_17607,N_14559);
and U22372 (N_22372,N_14654,N_12677);
nand U22373 (N_22373,N_13416,N_16735);
nand U22374 (N_22374,N_16487,N_15700);
and U22375 (N_22375,N_14972,N_18600);
and U22376 (N_22376,N_18554,N_12970);
or U22377 (N_22377,N_17497,N_13414);
xnor U22378 (N_22378,N_15739,N_13354);
nor U22379 (N_22379,N_18236,N_15110);
xnor U22380 (N_22380,N_16519,N_16518);
nand U22381 (N_22381,N_14113,N_15913);
xnor U22382 (N_22382,N_13603,N_14676);
nor U22383 (N_22383,N_15332,N_16916);
and U22384 (N_22384,N_17126,N_16410);
and U22385 (N_22385,N_16402,N_15992);
and U22386 (N_22386,N_17302,N_12557);
xnor U22387 (N_22387,N_13400,N_17089);
nor U22388 (N_22388,N_13925,N_14974);
and U22389 (N_22389,N_15505,N_14272);
and U22390 (N_22390,N_13980,N_15271);
and U22391 (N_22391,N_16093,N_14749);
and U22392 (N_22392,N_13597,N_15345);
nand U22393 (N_22393,N_16901,N_17039);
nand U22394 (N_22394,N_15570,N_15930);
nor U22395 (N_22395,N_18329,N_13356);
nand U22396 (N_22396,N_13762,N_15619);
or U22397 (N_22397,N_13817,N_16121);
nor U22398 (N_22398,N_17019,N_14137);
nand U22399 (N_22399,N_18369,N_14758);
nand U22400 (N_22400,N_14578,N_17306);
xor U22401 (N_22401,N_13722,N_13962);
or U22402 (N_22402,N_18643,N_14070);
nand U22403 (N_22403,N_17910,N_14736);
nor U22404 (N_22404,N_14696,N_13351);
xnor U22405 (N_22405,N_14321,N_16685);
and U22406 (N_22406,N_16476,N_14764);
or U22407 (N_22407,N_18499,N_15816);
or U22408 (N_22408,N_14039,N_13528);
or U22409 (N_22409,N_15765,N_18357);
nor U22410 (N_22410,N_13931,N_15305);
nor U22411 (N_22411,N_15450,N_15814);
nand U22412 (N_22412,N_15323,N_15297);
and U22413 (N_22413,N_16984,N_14044);
and U22414 (N_22414,N_18586,N_14215);
nand U22415 (N_22415,N_13102,N_14524);
xnor U22416 (N_22416,N_14744,N_13084);
nor U22417 (N_22417,N_13910,N_17961);
and U22418 (N_22418,N_18025,N_18009);
nor U22419 (N_22419,N_14773,N_15285);
and U22420 (N_22420,N_17680,N_14211);
nor U22421 (N_22421,N_17957,N_16386);
and U22422 (N_22422,N_14063,N_13947);
and U22423 (N_22423,N_15398,N_16030);
nand U22424 (N_22424,N_15381,N_12844);
or U22425 (N_22425,N_12647,N_17515);
nand U22426 (N_22426,N_17728,N_13199);
xnor U22427 (N_22427,N_17676,N_17148);
nand U22428 (N_22428,N_13786,N_15467);
nand U22429 (N_22429,N_16909,N_18680);
or U22430 (N_22430,N_13707,N_18617);
or U22431 (N_22431,N_14411,N_15523);
nand U22432 (N_22432,N_17885,N_13960);
xnor U22433 (N_22433,N_16842,N_16795);
and U22434 (N_22434,N_14619,N_13053);
or U22435 (N_22435,N_12914,N_15524);
and U22436 (N_22436,N_13267,N_13502);
nor U22437 (N_22437,N_16827,N_12792);
xor U22438 (N_22438,N_15162,N_12762);
and U22439 (N_22439,N_15800,N_15290);
and U22440 (N_22440,N_13300,N_13477);
or U22441 (N_22441,N_18112,N_18072);
and U22442 (N_22442,N_14244,N_13283);
or U22443 (N_22443,N_15889,N_13263);
nor U22444 (N_22444,N_12583,N_13398);
or U22445 (N_22445,N_14789,N_15005);
xnor U22446 (N_22446,N_15267,N_15050);
and U22447 (N_22447,N_17410,N_12617);
or U22448 (N_22448,N_18476,N_14161);
and U22449 (N_22449,N_15623,N_16315);
or U22450 (N_22450,N_15462,N_17460);
and U22451 (N_22451,N_16918,N_18555);
nor U22452 (N_22452,N_13144,N_14901);
nor U22453 (N_22453,N_12825,N_12746);
and U22454 (N_22454,N_18565,N_13860);
xnor U22455 (N_22455,N_17037,N_16984);
and U22456 (N_22456,N_15217,N_17749);
nor U22457 (N_22457,N_14934,N_15470);
xor U22458 (N_22458,N_14877,N_17261);
or U22459 (N_22459,N_14731,N_16329);
or U22460 (N_22460,N_18675,N_16408);
and U22461 (N_22461,N_15776,N_15862);
and U22462 (N_22462,N_12702,N_13782);
or U22463 (N_22463,N_15513,N_13275);
nand U22464 (N_22464,N_12700,N_16061);
nor U22465 (N_22465,N_17054,N_15827);
or U22466 (N_22466,N_16012,N_13673);
nor U22467 (N_22467,N_17107,N_12719);
nand U22468 (N_22468,N_15309,N_17486);
xor U22469 (N_22469,N_17796,N_14920);
nand U22470 (N_22470,N_14485,N_13830);
nand U22471 (N_22471,N_18076,N_16908);
nand U22472 (N_22472,N_18655,N_16359);
nor U22473 (N_22473,N_15119,N_14782);
and U22474 (N_22474,N_15248,N_18332);
xnor U22475 (N_22475,N_15245,N_13332);
and U22476 (N_22476,N_18087,N_16993);
nand U22477 (N_22477,N_15856,N_15924);
and U22478 (N_22478,N_14527,N_17424);
nand U22479 (N_22479,N_14630,N_12773);
xnor U22480 (N_22480,N_13204,N_12963);
or U22481 (N_22481,N_18196,N_14855);
nor U22482 (N_22482,N_13317,N_13304);
or U22483 (N_22483,N_15069,N_14433);
nor U22484 (N_22484,N_14029,N_16992);
nor U22485 (N_22485,N_18660,N_13412);
nor U22486 (N_22486,N_18140,N_18372);
nand U22487 (N_22487,N_13300,N_15585);
nor U22488 (N_22488,N_17258,N_18712);
nor U22489 (N_22489,N_13261,N_18536);
nand U22490 (N_22490,N_15231,N_15648);
and U22491 (N_22491,N_16606,N_18133);
nand U22492 (N_22492,N_14343,N_18724);
nor U22493 (N_22493,N_15068,N_16609);
nand U22494 (N_22494,N_14751,N_17259);
nor U22495 (N_22495,N_17758,N_14262);
nand U22496 (N_22496,N_14403,N_16029);
nand U22497 (N_22497,N_17005,N_18285);
nand U22498 (N_22498,N_15505,N_16766);
xor U22499 (N_22499,N_18358,N_12892);
nor U22500 (N_22500,N_13458,N_12833);
and U22501 (N_22501,N_15871,N_18152);
or U22502 (N_22502,N_14825,N_13002);
nor U22503 (N_22503,N_13383,N_15757);
or U22504 (N_22504,N_18378,N_18124);
and U22505 (N_22505,N_17882,N_14543);
nor U22506 (N_22506,N_14781,N_13506);
nand U22507 (N_22507,N_17231,N_17307);
or U22508 (N_22508,N_16855,N_14414);
and U22509 (N_22509,N_14881,N_17646);
or U22510 (N_22510,N_17721,N_12672);
and U22511 (N_22511,N_17051,N_15810);
xor U22512 (N_22512,N_15252,N_17958);
nor U22513 (N_22513,N_12721,N_17475);
or U22514 (N_22514,N_17557,N_13246);
xnor U22515 (N_22515,N_16274,N_12804);
and U22516 (N_22516,N_14969,N_15602);
nor U22517 (N_22517,N_14827,N_14734);
xor U22518 (N_22518,N_18279,N_18742);
or U22519 (N_22519,N_16703,N_15166);
nor U22520 (N_22520,N_17336,N_16974);
or U22521 (N_22521,N_14199,N_13564);
and U22522 (N_22522,N_15196,N_18613);
and U22523 (N_22523,N_13715,N_16942);
nand U22524 (N_22524,N_14048,N_16300);
and U22525 (N_22525,N_16479,N_16061);
and U22526 (N_22526,N_13674,N_18647);
or U22527 (N_22527,N_14449,N_15313);
nor U22528 (N_22528,N_16010,N_17263);
and U22529 (N_22529,N_12928,N_18098);
nor U22530 (N_22530,N_13841,N_15900);
nor U22531 (N_22531,N_15767,N_15497);
or U22532 (N_22532,N_15946,N_17982);
or U22533 (N_22533,N_15198,N_17192);
or U22534 (N_22534,N_13072,N_15225);
xor U22535 (N_22535,N_17214,N_15339);
nand U22536 (N_22536,N_14333,N_15924);
xnor U22537 (N_22537,N_16920,N_17581);
nor U22538 (N_22538,N_16290,N_18527);
and U22539 (N_22539,N_13142,N_18262);
nand U22540 (N_22540,N_18308,N_16532);
or U22541 (N_22541,N_16530,N_18294);
or U22542 (N_22542,N_17045,N_17758);
and U22543 (N_22543,N_12864,N_12663);
nor U22544 (N_22544,N_16236,N_13845);
nand U22545 (N_22545,N_14849,N_15346);
nand U22546 (N_22546,N_17461,N_17747);
or U22547 (N_22547,N_18004,N_15656);
nand U22548 (N_22548,N_14647,N_18156);
nor U22549 (N_22549,N_14717,N_15910);
xor U22550 (N_22550,N_17380,N_12929);
nor U22551 (N_22551,N_17480,N_16159);
nand U22552 (N_22552,N_17175,N_14343);
nor U22553 (N_22553,N_15996,N_18082);
nor U22554 (N_22554,N_18318,N_14485);
nor U22555 (N_22555,N_13864,N_16253);
and U22556 (N_22556,N_15804,N_18342);
nand U22557 (N_22557,N_16736,N_16075);
xnor U22558 (N_22558,N_15934,N_14168);
or U22559 (N_22559,N_17238,N_12823);
nor U22560 (N_22560,N_18386,N_18743);
nand U22561 (N_22561,N_13671,N_14167);
nand U22562 (N_22562,N_13447,N_17859);
nand U22563 (N_22563,N_18561,N_13610);
nor U22564 (N_22564,N_16783,N_17154);
nand U22565 (N_22565,N_18123,N_13313);
nor U22566 (N_22566,N_13830,N_17139);
and U22567 (N_22567,N_17759,N_15074);
or U22568 (N_22568,N_18143,N_14352);
nand U22569 (N_22569,N_18202,N_18085);
and U22570 (N_22570,N_16173,N_18179);
nand U22571 (N_22571,N_14869,N_14071);
or U22572 (N_22572,N_16276,N_17579);
nor U22573 (N_22573,N_18681,N_17963);
or U22574 (N_22574,N_14194,N_16054);
or U22575 (N_22575,N_17097,N_18644);
nand U22576 (N_22576,N_17666,N_14548);
nor U22577 (N_22577,N_14569,N_13885);
and U22578 (N_22578,N_14637,N_16111);
xor U22579 (N_22579,N_13848,N_13793);
nor U22580 (N_22580,N_16447,N_12506);
nand U22581 (N_22581,N_16697,N_14995);
nor U22582 (N_22582,N_13336,N_15965);
and U22583 (N_22583,N_13400,N_15660);
nand U22584 (N_22584,N_13898,N_16769);
nor U22585 (N_22585,N_17541,N_17913);
or U22586 (N_22586,N_12841,N_15280);
nor U22587 (N_22587,N_13091,N_14231);
and U22588 (N_22588,N_18148,N_12510);
and U22589 (N_22589,N_18700,N_14385);
and U22590 (N_22590,N_17279,N_14335);
nor U22591 (N_22591,N_18165,N_16214);
and U22592 (N_22592,N_13320,N_17192);
nor U22593 (N_22593,N_16888,N_14299);
nor U22594 (N_22594,N_13316,N_14412);
nand U22595 (N_22595,N_14589,N_16226);
nand U22596 (N_22596,N_12764,N_17448);
or U22597 (N_22597,N_16620,N_18291);
or U22598 (N_22598,N_13603,N_16791);
and U22599 (N_22599,N_17363,N_14131);
nor U22600 (N_22600,N_16433,N_14001);
or U22601 (N_22601,N_18007,N_14286);
or U22602 (N_22602,N_15488,N_16351);
and U22603 (N_22603,N_17861,N_18734);
or U22604 (N_22604,N_17254,N_18139);
and U22605 (N_22605,N_17450,N_14802);
nand U22606 (N_22606,N_15269,N_13257);
nor U22607 (N_22607,N_17639,N_17277);
nor U22608 (N_22608,N_12791,N_12824);
or U22609 (N_22609,N_14815,N_16807);
nor U22610 (N_22610,N_17182,N_17813);
xor U22611 (N_22611,N_15534,N_15803);
nand U22612 (N_22612,N_17191,N_15531);
and U22613 (N_22613,N_14602,N_15578);
xor U22614 (N_22614,N_16048,N_13658);
nand U22615 (N_22615,N_18387,N_17678);
nor U22616 (N_22616,N_13795,N_13218);
or U22617 (N_22617,N_14466,N_18502);
and U22618 (N_22618,N_15532,N_16882);
and U22619 (N_22619,N_16365,N_16832);
nor U22620 (N_22620,N_17189,N_17992);
nand U22621 (N_22621,N_14527,N_17199);
or U22622 (N_22622,N_16241,N_15309);
nor U22623 (N_22623,N_18719,N_17674);
nand U22624 (N_22624,N_13679,N_17566);
nand U22625 (N_22625,N_17977,N_13675);
xnor U22626 (N_22626,N_14051,N_15312);
nand U22627 (N_22627,N_13953,N_13210);
or U22628 (N_22628,N_17489,N_15244);
nand U22629 (N_22629,N_13099,N_16693);
nor U22630 (N_22630,N_16484,N_12915);
and U22631 (N_22631,N_15354,N_13076);
nand U22632 (N_22632,N_18312,N_14161);
or U22633 (N_22633,N_12520,N_17966);
and U22634 (N_22634,N_14210,N_14844);
nand U22635 (N_22635,N_12645,N_12503);
and U22636 (N_22636,N_12742,N_15179);
nand U22637 (N_22637,N_14350,N_13812);
and U22638 (N_22638,N_16512,N_16629);
nor U22639 (N_22639,N_16358,N_16004);
or U22640 (N_22640,N_15476,N_18445);
nand U22641 (N_22641,N_14589,N_17096);
xor U22642 (N_22642,N_13619,N_14686);
nand U22643 (N_22643,N_16565,N_18403);
nor U22644 (N_22644,N_13974,N_12735);
and U22645 (N_22645,N_16765,N_17209);
or U22646 (N_22646,N_17328,N_16781);
nor U22647 (N_22647,N_15497,N_18723);
and U22648 (N_22648,N_15699,N_14040);
or U22649 (N_22649,N_12998,N_17229);
and U22650 (N_22650,N_17800,N_15520);
nand U22651 (N_22651,N_12697,N_14611);
nand U22652 (N_22652,N_16567,N_16105);
or U22653 (N_22653,N_18368,N_18593);
or U22654 (N_22654,N_16754,N_12707);
or U22655 (N_22655,N_14740,N_18540);
or U22656 (N_22656,N_16048,N_18283);
or U22657 (N_22657,N_13785,N_15373);
nor U22658 (N_22658,N_15069,N_14674);
nand U22659 (N_22659,N_12556,N_13852);
nand U22660 (N_22660,N_16666,N_18051);
nor U22661 (N_22661,N_12527,N_18201);
and U22662 (N_22662,N_12873,N_13940);
and U22663 (N_22663,N_14110,N_16606);
and U22664 (N_22664,N_14618,N_14799);
nor U22665 (N_22665,N_16728,N_15403);
xnor U22666 (N_22666,N_15521,N_17512);
and U22667 (N_22667,N_13422,N_13302);
xor U22668 (N_22668,N_17895,N_12936);
xnor U22669 (N_22669,N_15449,N_15810);
or U22670 (N_22670,N_14689,N_18555);
xor U22671 (N_22671,N_13808,N_14638);
nand U22672 (N_22672,N_16962,N_16769);
or U22673 (N_22673,N_16841,N_18011);
nor U22674 (N_22674,N_12652,N_18647);
xor U22675 (N_22675,N_17465,N_15136);
nand U22676 (N_22676,N_13838,N_12810);
nand U22677 (N_22677,N_13625,N_15343);
and U22678 (N_22678,N_15979,N_12868);
xnor U22679 (N_22679,N_15834,N_12838);
nor U22680 (N_22680,N_14643,N_14149);
nand U22681 (N_22681,N_16993,N_15521);
xor U22682 (N_22682,N_17251,N_16507);
or U22683 (N_22683,N_12822,N_14995);
nand U22684 (N_22684,N_16801,N_17365);
xnor U22685 (N_22685,N_17180,N_16718);
xor U22686 (N_22686,N_12644,N_15523);
and U22687 (N_22687,N_17982,N_14343);
nand U22688 (N_22688,N_16823,N_14256);
and U22689 (N_22689,N_18642,N_12662);
nand U22690 (N_22690,N_13476,N_18341);
nand U22691 (N_22691,N_14396,N_13165);
nor U22692 (N_22692,N_13452,N_17244);
nand U22693 (N_22693,N_14743,N_18746);
nand U22694 (N_22694,N_16855,N_15822);
and U22695 (N_22695,N_18166,N_18093);
xnor U22696 (N_22696,N_13968,N_17776);
nor U22697 (N_22697,N_16401,N_17533);
or U22698 (N_22698,N_17495,N_17903);
or U22699 (N_22699,N_13730,N_18138);
and U22700 (N_22700,N_13715,N_17321);
xnor U22701 (N_22701,N_13828,N_14914);
nor U22702 (N_22702,N_16770,N_17418);
or U22703 (N_22703,N_17261,N_16876);
nor U22704 (N_22704,N_15347,N_18732);
or U22705 (N_22705,N_15572,N_15329);
nor U22706 (N_22706,N_13378,N_12585);
nand U22707 (N_22707,N_18129,N_17161);
nand U22708 (N_22708,N_12624,N_18162);
nand U22709 (N_22709,N_17616,N_15675);
nand U22710 (N_22710,N_18129,N_14126);
or U22711 (N_22711,N_14164,N_13478);
xor U22712 (N_22712,N_14187,N_17574);
xor U22713 (N_22713,N_17102,N_14261);
and U22714 (N_22714,N_17819,N_18086);
nand U22715 (N_22715,N_13695,N_16033);
and U22716 (N_22716,N_17771,N_15765);
and U22717 (N_22717,N_13988,N_17627);
or U22718 (N_22718,N_18332,N_14917);
nand U22719 (N_22719,N_17951,N_12979);
xnor U22720 (N_22720,N_16762,N_14938);
and U22721 (N_22721,N_17351,N_18611);
nand U22722 (N_22722,N_18236,N_15291);
and U22723 (N_22723,N_12889,N_18043);
or U22724 (N_22724,N_13478,N_17876);
nand U22725 (N_22725,N_16779,N_16666);
or U22726 (N_22726,N_13862,N_13385);
nor U22727 (N_22727,N_16171,N_17468);
or U22728 (N_22728,N_13580,N_16078);
or U22729 (N_22729,N_16355,N_14611);
and U22730 (N_22730,N_13615,N_16335);
nand U22731 (N_22731,N_15571,N_15031);
xor U22732 (N_22732,N_16855,N_13059);
or U22733 (N_22733,N_16020,N_16929);
and U22734 (N_22734,N_16514,N_14868);
and U22735 (N_22735,N_14276,N_12806);
or U22736 (N_22736,N_15371,N_18107);
and U22737 (N_22737,N_13169,N_17794);
or U22738 (N_22738,N_16064,N_14182);
nand U22739 (N_22739,N_13399,N_14196);
or U22740 (N_22740,N_16539,N_13281);
nor U22741 (N_22741,N_16484,N_14513);
or U22742 (N_22742,N_13563,N_18398);
xor U22743 (N_22743,N_13161,N_16285);
and U22744 (N_22744,N_14155,N_15301);
nor U22745 (N_22745,N_13533,N_16523);
or U22746 (N_22746,N_12541,N_15691);
and U22747 (N_22747,N_16005,N_13691);
nand U22748 (N_22748,N_17623,N_14072);
nor U22749 (N_22749,N_13643,N_17430);
nor U22750 (N_22750,N_15957,N_14647);
or U22751 (N_22751,N_18667,N_15578);
nand U22752 (N_22752,N_13420,N_14576);
or U22753 (N_22753,N_17415,N_15464);
and U22754 (N_22754,N_12787,N_17942);
and U22755 (N_22755,N_16014,N_18030);
and U22756 (N_22756,N_14710,N_12758);
nor U22757 (N_22757,N_15140,N_13203);
or U22758 (N_22758,N_13957,N_16771);
or U22759 (N_22759,N_15874,N_17829);
nand U22760 (N_22760,N_16504,N_16659);
nand U22761 (N_22761,N_14079,N_13217);
xnor U22762 (N_22762,N_16830,N_14125);
nor U22763 (N_22763,N_18559,N_18597);
nand U22764 (N_22764,N_14077,N_16876);
and U22765 (N_22765,N_17803,N_14502);
nor U22766 (N_22766,N_13550,N_13157);
nor U22767 (N_22767,N_15452,N_18488);
nor U22768 (N_22768,N_16010,N_15214);
and U22769 (N_22769,N_12932,N_17761);
nor U22770 (N_22770,N_18034,N_18002);
nor U22771 (N_22771,N_18747,N_15953);
and U22772 (N_22772,N_12820,N_15433);
and U22773 (N_22773,N_15215,N_16650);
nand U22774 (N_22774,N_13291,N_17438);
or U22775 (N_22775,N_16186,N_14027);
and U22776 (N_22776,N_17283,N_15717);
nand U22777 (N_22777,N_17922,N_15570);
or U22778 (N_22778,N_12901,N_18619);
nand U22779 (N_22779,N_16237,N_16262);
and U22780 (N_22780,N_16575,N_14025);
xnor U22781 (N_22781,N_18329,N_16681);
nand U22782 (N_22782,N_17339,N_17595);
and U22783 (N_22783,N_13465,N_15066);
xor U22784 (N_22784,N_16874,N_12544);
and U22785 (N_22785,N_18615,N_16073);
or U22786 (N_22786,N_15265,N_17382);
nand U22787 (N_22787,N_12679,N_15651);
nand U22788 (N_22788,N_15828,N_16429);
and U22789 (N_22789,N_18509,N_16503);
nand U22790 (N_22790,N_15027,N_13516);
nand U22791 (N_22791,N_13787,N_15085);
and U22792 (N_22792,N_12626,N_18284);
or U22793 (N_22793,N_18148,N_14261);
or U22794 (N_22794,N_16883,N_13690);
nand U22795 (N_22795,N_15232,N_15654);
and U22796 (N_22796,N_15592,N_15285);
nor U22797 (N_22797,N_13718,N_16449);
nor U22798 (N_22798,N_16769,N_14010);
nor U22799 (N_22799,N_15351,N_18460);
nor U22800 (N_22800,N_13081,N_14012);
nand U22801 (N_22801,N_16314,N_13203);
nor U22802 (N_22802,N_18720,N_17148);
or U22803 (N_22803,N_17819,N_16508);
or U22804 (N_22804,N_15071,N_16337);
and U22805 (N_22805,N_14881,N_15605);
nand U22806 (N_22806,N_15134,N_16530);
and U22807 (N_22807,N_17400,N_16953);
nand U22808 (N_22808,N_13461,N_14867);
and U22809 (N_22809,N_12509,N_16021);
nand U22810 (N_22810,N_17841,N_17134);
and U22811 (N_22811,N_14455,N_15435);
or U22812 (N_22812,N_17200,N_13309);
and U22813 (N_22813,N_15308,N_16966);
or U22814 (N_22814,N_17584,N_18316);
or U22815 (N_22815,N_17236,N_15926);
nand U22816 (N_22816,N_13125,N_15077);
and U22817 (N_22817,N_13889,N_15119);
or U22818 (N_22818,N_14787,N_15935);
nor U22819 (N_22819,N_18372,N_16019);
xor U22820 (N_22820,N_17122,N_13757);
nor U22821 (N_22821,N_13334,N_16614);
xnor U22822 (N_22822,N_13456,N_16142);
and U22823 (N_22823,N_16588,N_14750);
nor U22824 (N_22824,N_14270,N_14723);
nor U22825 (N_22825,N_17706,N_15797);
nand U22826 (N_22826,N_13503,N_17213);
or U22827 (N_22827,N_15709,N_15204);
or U22828 (N_22828,N_14299,N_16512);
xor U22829 (N_22829,N_14053,N_12754);
or U22830 (N_22830,N_13162,N_16466);
nor U22831 (N_22831,N_16217,N_12529);
nor U22832 (N_22832,N_18348,N_17332);
nor U22833 (N_22833,N_16429,N_13139);
nor U22834 (N_22834,N_12530,N_15426);
nor U22835 (N_22835,N_15579,N_12590);
nand U22836 (N_22836,N_16367,N_14983);
xnor U22837 (N_22837,N_13911,N_15190);
nand U22838 (N_22838,N_13298,N_13396);
or U22839 (N_22839,N_14303,N_17523);
or U22840 (N_22840,N_17355,N_14575);
nor U22841 (N_22841,N_15102,N_15898);
nand U22842 (N_22842,N_18460,N_15685);
nor U22843 (N_22843,N_14191,N_16614);
or U22844 (N_22844,N_14060,N_18159);
and U22845 (N_22845,N_14662,N_16077);
nand U22846 (N_22846,N_18555,N_17625);
nor U22847 (N_22847,N_15332,N_18243);
xor U22848 (N_22848,N_17093,N_15916);
or U22849 (N_22849,N_17241,N_15470);
nand U22850 (N_22850,N_15102,N_12947);
or U22851 (N_22851,N_17257,N_18552);
or U22852 (N_22852,N_12843,N_16428);
or U22853 (N_22853,N_13609,N_16803);
and U22854 (N_22854,N_17676,N_15542);
nor U22855 (N_22855,N_14005,N_15783);
and U22856 (N_22856,N_16196,N_13486);
nand U22857 (N_22857,N_16834,N_15519);
or U22858 (N_22858,N_18104,N_13264);
nor U22859 (N_22859,N_14003,N_15901);
nor U22860 (N_22860,N_12632,N_14268);
xor U22861 (N_22861,N_15535,N_15310);
nor U22862 (N_22862,N_15345,N_13282);
and U22863 (N_22863,N_12552,N_13535);
nand U22864 (N_22864,N_12830,N_16191);
and U22865 (N_22865,N_14026,N_15833);
nand U22866 (N_22866,N_13058,N_16113);
and U22867 (N_22867,N_13232,N_14448);
or U22868 (N_22868,N_12577,N_15369);
or U22869 (N_22869,N_16895,N_14839);
nand U22870 (N_22870,N_14588,N_18545);
nor U22871 (N_22871,N_14102,N_17487);
nor U22872 (N_22872,N_12867,N_18368);
and U22873 (N_22873,N_17580,N_14761);
or U22874 (N_22874,N_13702,N_12925);
nor U22875 (N_22875,N_18036,N_18683);
nor U22876 (N_22876,N_17694,N_14728);
nor U22877 (N_22877,N_14624,N_15226);
and U22878 (N_22878,N_17235,N_17228);
or U22879 (N_22879,N_14510,N_14727);
nor U22880 (N_22880,N_12520,N_17080);
nor U22881 (N_22881,N_16259,N_16448);
xor U22882 (N_22882,N_15782,N_17267);
or U22883 (N_22883,N_15247,N_17398);
nand U22884 (N_22884,N_13806,N_16160);
nand U22885 (N_22885,N_16786,N_14217);
nor U22886 (N_22886,N_17028,N_17275);
and U22887 (N_22887,N_18017,N_18520);
and U22888 (N_22888,N_12947,N_17490);
or U22889 (N_22889,N_16624,N_13726);
or U22890 (N_22890,N_15411,N_17185);
nand U22891 (N_22891,N_18370,N_12653);
xor U22892 (N_22892,N_16577,N_13160);
xnor U22893 (N_22893,N_14807,N_16181);
nand U22894 (N_22894,N_15105,N_16804);
and U22895 (N_22895,N_18019,N_15098);
or U22896 (N_22896,N_13298,N_15117);
nand U22897 (N_22897,N_12991,N_12735);
xnor U22898 (N_22898,N_17745,N_17302);
nand U22899 (N_22899,N_15417,N_16794);
or U22900 (N_22900,N_13082,N_15055);
and U22901 (N_22901,N_18314,N_15605);
and U22902 (N_22902,N_13547,N_15679);
or U22903 (N_22903,N_15986,N_18610);
xnor U22904 (N_22904,N_17252,N_14031);
nand U22905 (N_22905,N_16151,N_14358);
and U22906 (N_22906,N_15759,N_13999);
nor U22907 (N_22907,N_14649,N_15412);
and U22908 (N_22908,N_15110,N_18043);
nor U22909 (N_22909,N_17788,N_14560);
and U22910 (N_22910,N_16365,N_14351);
nor U22911 (N_22911,N_17267,N_18473);
nor U22912 (N_22912,N_18371,N_16896);
xor U22913 (N_22913,N_18657,N_13140);
nand U22914 (N_22914,N_14047,N_12500);
or U22915 (N_22915,N_15264,N_18677);
nor U22916 (N_22916,N_17805,N_16382);
or U22917 (N_22917,N_18632,N_13032);
and U22918 (N_22918,N_14370,N_16110);
and U22919 (N_22919,N_15275,N_17702);
nor U22920 (N_22920,N_14159,N_15675);
and U22921 (N_22921,N_16001,N_13120);
nand U22922 (N_22922,N_17795,N_17786);
nor U22923 (N_22923,N_15628,N_16067);
and U22924 (N_22924,N_17756,N_14858);
xor U22925 (N_22925,N_14461,N_13694);
and U22926 (N_22926,N_17520,N_14556);
nand U22927 (N_22927,N_17666,N_12602);
nor U22928 (N_22928,N_17796,N_17280);
or U22929 (N_22929,N_18087,N_14863);
and U22930 (N_22930,N_13289,N_12523);
and U22931 (N_22931,N_17242,N_14010);
nand U22932 (N_22932,N_17684,N_17300);
and U22933 (N_22933,N_16219,N_18678);
nand U22934 (N_22934,N_17263,N_13629);
nand U22935 (N_22935,N_13596,N_13685);
or U22936 (N_22936,N_15257,N_13490);
or U22937 (N_22937,N_15405,N_15322);
nor U22938 (N_22938,N_17327,N_14507);
nor U22939 (N_22939,N_15291,N_18363);
nor U22940 (N_22940,N_18629,N_13263);
nand U22941 (N_22941,N_14999,N_15721);
and U22942 (N_22942,N_14273,N_16501);
and U22943 (N_22943,N_15029,N_12810);
nor U22944 (N_22944,N_16995,N_12833);
or U22945 (N_22945,N_13048,N_17051);
nand U22946 (N_22946,N_18315,N_17573);
nand U22947 (N_22947,N_17020,N_17862);
nor U22948 (N_22948,N_16330,N_15438);
xnor U22949 (N_22949,N_17461,N_18211);
nand U22950 (N_22950,N_14042,N_17228);
nand U22951 (N_22951,N_17170,N_16806);
xnor U22952 (N_22952,N_15269,N_14025);
and U22953 (N_22953,N_12962,N_12867);
nand U22954 (N_22954,N_18169,N_14231);
xor U22955 (N_22955,N_17942,N_13727);
or U22956 (N_22956,N_13599,N_13744);
xnor U22957 (N_22957,N_15580,N_13423);
nand U22958 (N_22958,N_17735,N_18653);
xnor U22959 (N_22959,N_13403,N_17121);
or U22960 (N_22960,N_17031,N_13905);
nand U22961 (N_22961,N_17600,N_14467);
xnor U22962 (N_22962,N_15620,N_18606);
and U22963 (N_22963,N_12989,N_17376);
and U22964 (N_22964,N_18714,N_12875);
and U22965 (N_22965,N_18163,N_14299);
nand U22966 (N_22966,N_13105,N_16868);
and U22967 (N_22967,N_13209,N_16928);
nor U22968 (N_22968,N_13468,N_16381);
and U22969 (N_22969,N_18226,N_18205);
or U22970 (N_22970,N_16642,N_16157);
xor U22971 (N_22971,N_15390,N_12718);
xor U22972 (N_22972,N_13306,N_12939);
nand U22973 (N_22973,N_12891,N_13482);
nor U22974 (N_22974,N_18154,N_14812);
nor U22975 (N_22975,N_15474,N_12856);
nor U22976 (N_22976,N_17076,N_14144);
and U22977 (N_22977,N_14454,N_15123);
nor U22978 (N_22978,N_18653,N_15277);
nor U22979 (N_22979,N_16959,N_14538);
nand U22980 (N_22980,N_16841,N_15060);
or U22981 (N_22981,N_13920,N_13438);
nor U22982 (N_22982,N_17179,N_18687);
xor U22983 (N_22983,N_17054,N_18570);
nand U22984 (N_22984,N_14062,N_14195);
or U22985 (N_22985,N_13238,N_16810);
nand U22986 (N_22986,N_12710,N_16626);
or U22987 (N_22987,N_15838,N_16954);
nor U22988 (N_22988,N_13846,N_12658);
nor U22989 (N_22989,N_13395,N_15209);
xor U22990 (N_22990,N_16751,N_12557);
nand U22991 (N_22991,N_14690,N_17317);
nor U22992 (N_22992,N_15384,N_15135);
or U22993 (N_22993,N_12645,N_14114);
and U22994 (N_22994,N_12806,N_14698);
nor U22995 (N_22995,N_14694,N_15330);
and U22996 (N_22996,N_12838,N_15236);
nand U22997 (N_22997,N_16047,N_18667);
nor U22998 (N_22998,N_18553,N_13334);
xnor U22999 (N_22999,N_14934,N_16710);
and U23000 (N_23000,N_13120,N_16690);
and U23001 (N_23001,N_18249,N_13201);
xnor U23002 (N_23002,N_16980,N_17622);
or U23003 (N_23003,N_15352,N_17315);
nand U23004 (N_23004,N_14162,N_18646);
nor U23005 (N_23005,N_17048,N_16825);
nand U23006 (N_23006,N_15509,N_14963);
and U23007 (N_23007,N_14089,N_15219);
nor U23008 (N_23008,N_14041,N_16502);
nor U23009 (N_23009,N_16104,N_17949);
nor U23010 (N_23010,N_16725,N_18622);
nand U23011 (N_23011,N_13573,N_13404);
and U23012 (N_23012,N_16285,N_16856);
nor U23013 (N_23013,N_15314,N_16341);
or U23014 (N_23014,N_15012,N_17160);
or U23015 (N_23015,N_13114,N_13650);
xor U23016 (N_23016,N_14326,N_18466);
and U23017 (N_23017,N_15101,N_14676);
nor U23018 (N_23018,N_14677,N_12946);
nor U23019 (N_23019,N_14926,N_18249);
or U23020 (N_23020,N_15956,N_13141);
xor U23021 (N_23021,N_13988,N_13644);
nor U23022 (N_23022,N_18721,N_16190);
nand U23023 (N_23023,N_15567,N_18194);
and U23024 (N_23024,N_15381,N_12504);
xnor U23025 (N_23025,N_15554,N_18402);
nor U23026 (N_23026,N_12668,N_12774);
nor U23027 (N_23027,N_14366,N_17712);
or U23028 (N_23028,N_17525,N_14376);
nand U23029 (N_23029,N_16767,N_16868);
and U23030 (N_23030,N_16368,N_18731);
or U23031 (N_23031,N_12713,N_15289);
and U23032 (N_23032,N_15419,N_12652);
and U23033 (N_23033,N_17359,N_17165);
nand U23034 (N_23034,N_12597,N_16333);
nand U23035 (N_23035,N_14453,N_13850);
nor U23036 (N_23036,N_12603,N_15266);
or U23037 (N_23037,N_17843,N_17421);
nor U23038 (N_23038,N_13493,N_17677);
and U23039 (N_23039,N_18032,N_13819);
xor U23040 (N_23040,N_13027,N_14376);
or U23041 (N_23041,N_18175,N_18248);
xor U23042 (N_23042,N_15160,N_15889);
and U23043 (N_23043,N_15561,N_13395);
xnor U23044 (N_23044,N_13865,N_15056);
or U23045 (N_23045,N_15255,N_16050);
or U23046 (N_23046,N_12744,N_14781);
nor U23047 (N_23047,N_13595,N_14042);
nor U23048 (N_23048,N_14852,N_14509);
and U23049 (N_23049,N_12581,N_14302);
or U23050 (N_23050,N_13361,N_17828);
or U23051 (N_23051,N_17047,N_15068);
or U23052 (N_23052,N_17101,N_13327);
nand U23053 (N_23053,N_13655,N_14225);
nor U23054 (N_23054,N_14286,N_12613);
and U23055 (N_23055,N_16954,N_17890);
or U23056 (N_23056,N_13584,N_17609);
nand U23057 (N_23057,N_18256,N_15527);
xor U23058 (N_23058,N_18145,N_15910);
or U23059 (N_23059,N_15778,N_15680);
and U23060 (N_23060,N_15845,N_13152);
nor U23061 (N_23061,N_13199,N_16494);
or U23062 (N_23062,N_13799,N_18526);
nand U23063 (N_23063,N_18016,N_18071);
or U23064 (N_23064,N_16221,N_15522);
or U23065 (N_23065,N_14322,N_16849);
or U23066 (N_23066,N_15674,N_15920);
and U23067 (N_23067,N_16310,N_16756);
nor U23068 (N_23068,N_13777,N_17212);
and U23069 (N_23069,N_16473,N_16928);
or U23070 (N_23070,N_18472,N_15601);
and U23071 (N_23071,N_17133,N_14380);
or U23072 (N_23072,N_18624,N_17066);
and U23073 (N_23073,N_16058,N_17520);
nor U23074 (N_23074,N_15169,N_16227);
or U23075 (N_23075,N_12903,N_13284);
nand U23076 (N_23076,N_14787,N_12839);
or U23077 (N_23077,N_17551,N_17191);
nand U23078 (N_23078,N_17765,N_14206);
nand U23079 (N_23079,N_15143,N_13256);
xor U23080 (N_23080,N_17582,N_16382);
nand U23081 (N_23081,N_18581,N_16124);
or U23082 (N_23082,N_13952,N_17859);
nand U23083 (N_23083,N_16165,N_15731);
xnor U23084 (N_23084,N_13283,N_17149);
nand U23085 (N_23085,N_17829,N_16245);
or U23086 (N_23086,N_17268,N_15626);
or U23087 (N_23087,N_16227,N_16503);
and U23088 (N_23088,N_15811,N_16996);
nor U23089 (N_23089,N_14094,N_18276);
xor U23090 (N_23090,N_17225,N_15650);
nand U23091 (N_23091,N_15456,N_13855);
nor U23092 (N_23092,N_18241,N_14226);
nor U23093 (N_23093,N_16328,N_18422);
nor U23094 (N_23094,N_15120,N_12513);
or U23095 (N_23095,N_18256,N_12752);
nand U23096 (N_23096,N_15428,N_14618);
nand U23097 (N_23097,N_16149,N_18475);
nand U23098 (N_23098,N_15116,N_15916);
nor U23099 (N_23099,N_17235,N_13685);
nor U23100 (N_23100,N_15635,N_12528);
and U23101 (N_23101,N_16049,N_18547);
nor U23102 (N_23102,N_15550,N_13375);
nor U23103 (N_23103,N_15222,N_15770);
and U23104 (N_23104,N_13834,N_17998);
or U23105 (N_23105,N_17253,N_12944);
and U23106 (N_23106,N_13046,N_14028);
and U23107 (N_23107,N_13089,N_14136);
or U23108 (N_23108,N_14939,N_13905);
or U23109 (N_23109,N_12778,N_16465);
and U23110 (N_23110,N_15578,N_18089);
nand U23111 (N_23111,N_14211,N_17517);
xnor U23112 (N_23112,N_14938,N_15008);
and U23113 (N_23113,N_16350,N_15768);
or U23114 (N_23114,N_16108,N_15951);
and U23115 (N_23115,N_17567,N_16918);
nand U23116 (N_23116,N_14211,N_13397);
nor U23117 (N_23117,N_17716,N_15190);
and U23118 (N_23118,N_14472,N_14162);
or U23119 (N_23119,N_17075,N_14650);
xor U23120 (N_23120,N_12870,N_15219);
nand U23121 (N_23121,N_17115,N_15587);
nand U23122 (N_23122,N_13268,N_14836);
xor U23123 (N_23123,N_16134,N_13963);
nor U23124 (N_23124,N_15043,N_18275);
xnor U23125 (N_23125,N_14476,N_15023);
xor U23126 (N_23126,N_13144,N_17605);
nand U23127 (N_23127,N_18101,N_12943);
nor U23128 (N_23128,N_15200,N_13231);
nand U23129 (N_23129,N_14286,N_18077);
and U23130 (N_23130,N_18706,N_16877);
nor U23131 (N_23131,N_16456,N_17858);
nor U23132 (N_23132,N_14319,N_16411);
nand U23133 (N_23133,N_18662,N_15760);
nand U23134 (N_23134,N_14343,N_14492);
nand U23135 (N_23135,N_17634,N_13494);
nor U23136 (N_23136,N_14979,N_14794);
nor U23137 (N_23137,N_16422,N_14092);
and U23138 (N_23138,N_17628,N_13246);
nor U23139 (N_23139,N_18686,N_17796);
nand U23140 (N_23140,N_14357,N_15601);
nor U23141 (N_23141,N_18682,N_16809);
nand U23142 (N_23142,N_17041,N_15035);
nor U23143 (N_23143,N_13308,N_18725);
and U23144 (N_23144,N_14944,N_13616);
nand U23145 (N_23145,N_14844,N_18477);
nor U23146 (N_23146,N_15192,N_14722);
or U23147 (N_23147,N_15450,N_17907);
or U23148 (N_23148,N_17961,N_18321);
nor U23149 (N_23149,N_13229,N_12671);
and U23150 (N_23150,N_17863,N_12576);
nand U23151 (N_23151,N_12952,N_16565);
or U23152 (N_23152,N_17256,N_12745);
or U23153 (N_23153,N_14360,N_14493);
nand U23154 (N_23154,N_17755,N_17144);
nand U23155 (N_23155,N_15361,N_18449);
or U23156 (N_23156,N_15971,N_12514);
nor U23157 (N_23157,N_17676,N_14296);
xor U23158 (N_23158,N_18503,N_17140);
nand U23159 (N_23159,N_17536,N_18064);
nand U23160 (N_23160,N_13774,N_15030);
nand U23161 (N_23161,N_14461,N_16015);
xnor U23162 (N_23162,N_18683,N_16745);
or U23163 (N_23163,N_18561,N_14683);
or U23164 (N_23164,N_17675,N_17765);
or U23165 (N_23165,N_17192,N_17028);
nand U23166 (N_23166,N_18075,N_13695);
nand U23167 (N_23167,N_18038,N_18730);
nand U23168 (N_23168,N_17660,N_17794);
nand U23169 (N_23169,N_15022,N_16540);
or U23170 (N_23170,N_14515,N_17183);
or U23171 (N_23171,N_14898,N_15816);
nand U23172 (N_23172,N_15879,N_13082);
nor U23173 (N_23173,N_17081,N_17104);
or U23174 (N_23174,N_16779,N_12741);
nand U23175 (N_23175,N_18242,N_18188);
xnor U23176 (N_23176,N_16732,N_18500);
nand U23177 (N_23177,N_16549,N_13622);
and U23178 (N_23178,N_13320,N_12842);
and U23179 (N_23179,N_13984,N_13303);
or U23180 (N_23180,N_13200,N_13177);
and U23181 (N_23181,N_12727,N_15629);
or U23182 (N_23182,N_12739,N_18463);
or U23183 (N_23183,N_13398,N_17140);
nand U23184 (N_23184,N_13914,N_14089);
nor U23185 (N_23185,N_18031,N_16944);
nor U23186 (N_23186,N_14314,N_17897);
or U23187 (N_23187,N_15174,N_14988);
and U23188 (N_23188,N_18423,N_16621);
or U23189 (N_23189,N_15583,N_13824);
nand U23190 (N_23190,N_17954,N_14404);
nor U23191 (N_23191,N_13739,N_13576);
nand U23192 (N_23192,N_13983,N_17862);
and U23193 (N_23193,N_14897,N_17091);
or U23194 (N_23194,N_16110,N_18649);
or U23195 (N_23195,N_16050,N_14135);
nand U23196 (N_23196,N_16566,N_15347);
nand U23197 (N_23197,N_13711,N_16670);
and U23198 (N_23198,N_17139,N_15507);
and U23199 (N_23199,N_18543,N_14436);
and U23200 (N_23200,N_17581,N_13028);
nor U23201 (N_23201,N_14237,N_14447);
or U23202 (N_23202,N_17444,N_13597);
nand U23203 (N_23203,N_12767,N_14909);
or U23204 (N_23204,N_17227,N_15370);
and U23205 (N_23205,N_16537,N_13080);
nand U23206 (N_23206,N_17467,N_16229);
or U23207 (N_23207,N_17910,N_18219);
and U23208 (N_23208,N_14661,N_15970);
or U23209 (N_23209,N_17582,N_12747);
nor U23210 (N_23210,N_16889,N_14880);
and U23211 (N_23211,N_13464,N_17841);
or U23212 (N_23212,N_12876,N_17200);
nand U23213 (N_23213,N_17699,N_12536);
nor U23214 (N_23214,N_15252,N_18602);
or U23215 (N_23215,N_18515,N_17652);
and U23216 (N_23216,N_16055,N_12651);
and U23217 (N_23217,N_14196,N_12865);
or U23218 (N_23218,N_13456,N_17656);
or U23219 (N_23219,N_12562,N_13449);
nor U23220 (N_23220,N_14525,N_18084);
or U23221 (N_23221,N_16441,N_18712);
nand U23222 (N_23222,N_16414,N_18071);
and U23223 (N_23223,N_17437,N_13250);
xnor U23224 (N_23224,N_15250,N_14108);
and U23225 (N_23225,N_14177,N_17287);
nand U23226 (N_23226,N_17336,N_13347);
nor U23227 (N_23227,N_13169,N_14692);
or U23228 (N_23228,N_15580,N_13207);
nand U23229 (N_23229,N_15592,N_18738);
and U23230 (N_23230,N_17703,N_15879);
or U23231 (N_23231,N_13370,N_12565);
nand U23232 (N_23232,N_13958,N_14226);
and U23233 (N_23233,N_16135,N_13438);
nand U23234 (N_23234,N_15779,N_16130);
nand U23235 (N_23235,N_15828,N_13227);
nand U23236 (N_23236,N_12642,N_18207);
nor U23237 (N_23237,N_18243,N_13453);
and U23238 (N_23238,N_18477,N_16878);
or U23239 (N_23239,N_15712,N_15067);
nand U23240 (N_23240,N_12857,N_13344);
nand U23241 (N_23241,N_16017,N_15186);
or U23242 (N_23242,N_14225,N_16899);
and U23243 (N_23243,N_17475,N_15086);
or U23244 (N_23244,N_15785,N_17020);
and U23245 (N_23245,N_12680,N_15334);
nand U23246 (N_23246,N_16670,N_14252);
or U23247 (N_23247,N_16741,N_18012);
nor U23248 (N_23248,N_14449,N_13210);
nand U23249 (N_23249,N_15594,N_17116);
or U23250 (N_23250,N_14504,N_18565);
nand U23251 (N_23251,N_15843,N_17045);
nor U23252 (N_23252,N_12595,N_13232);
xnor U23253 (N_23253,N_16584,N_18642);
nor U23254 (N_23254,N_15173,N_16408);
and U23255 (N_23255,N_18524,N_17452);
nor U23256 (N_23256,N_15636,N_17629);
nand U23257 (N_23257,N_12894,N_17900);
and U23258 (N_23258,N_15760,N_18001);
nor U23259 (N_23259,N_15694,N_18517);
nand U23260 (N_23260,N_14751,N_13798);
or U23261 (N_23261,N_18707,N_14795);
and U23262 (N_23262,N_14780,N_18128);
nor U23263 (N_23263,N_14123,N_15961);
xor U23264 (N_23264,N_15257,N_12758);
nand U23265 (N_23265,N_15972,N_15608);
and U23266 (N_23266,N_12720,N_13056);
or U23267 (N_23267,N_16915,N_16878);
nor U23268 (N_23268,N_12792,N_15917);
or U23269 (N_23269,N_18679,N_16436);
or U23270 (N_23270,N_15092,N_16721);
nand U23271 (N_23271,N_13248,N_18226);
nor U23272 (N_23272,N_16211,N_15857);
and U23273 (N_23273,N_15420,N_13618);
or U23274 (N_23274,N_18253,N_13620);
or U23275 (N_23275,N_18377,N_18651);
and U23276 (N_23276,N_16007,N_15741);
or U23277 (N_23277,N_14827,N_15300);
nand U23278 (N_23278,N_17650,N_13421);
nor U23279 (N_23279,N_17715,N_17117);
or U23280 (N_23280,N_16045,N_13715);
xor U23281 (N_23281,N_16709,N_15902);
nand U23282 (N_23282,N_16790,N_13448);
nor U23283 (N_23283,N_15375,N_15676);
or U23284 (N_23284,N_15994,N_16124);
nor U23285 (N_23285,N_15695,N_17556);
nor U23286 (N_23286,N_14368,N_18369);
or U23287 (N_23287,N_18063,N_17046);
or U23288 (N_23288,N_14889,N_13582);
nor U23289 (N_23289,N_14763,N_15557);
or U23290 (N_23290,N_15060,N_17737);
nor U23291 (N_23291,N_16355,N_18149);
nor U23292 (N_23292,N_14192,N_13469);
nor U23293 (N_23293,N_16398,N_13083);
xor U23294 (N_23294,N_17295,N_15658);
nand U23295 (N_23295,N_13043,N_15485);
nand U23296 (N_23296,N_15072,N_14246);
and U23297 (N_23297,N_18389,N_13416);
nor U23298 (N_23298,N_16864,N_13356);
and U23299 (N_23299,N_16889,N_15659);
nand U23300 (N_23300,N_18749,N_12578);
xor U23301 (N_23301,N_12732,N_15335);
xor U23302 (N_23302,N_14036,N_16061);
nor U23303 (N_23303,N_16892,N_17374);
xor U23304 (N_23304,N_15769,N_16963);
nor U23305 (N_23305,N_16080,N_16624);
or U23306 (N_23306,N_12888,N_17607);
or U23307 (N_23307,N_16624,N_12548);
nor U23308 (N_23308,N_13545,N_15346);
xnor U23309 (N_23309,N_12954,N_14796);
nor U23310 (N_23310,N_15644,N_13470);
xor U23311 (N_23311,N_16773,N_17210);
xor U23312 (N_23312,N_12663,N_17002);
and U23313 (N_23313,N_14428,N_13799);
and U23314 (N_23314,N_17234,N_12750);
or U23315 (N_23315,N_16194,N_17042);
nor U23316 (N_23316,N_13577,N_15589);
nand U23317 (N_23317,N_17676,N_12944);
nand U23318 (N_23318,N_16570,N_18396);
and U23319 (N_23319,N_16794,N_14886);
nand U23320 (N_23320,N_16054,N_12647);
nor U23321 (N_23321,N_13045,N_13819);
or U23322 (N_23322,N_16116,N_15394);
and U23323 (N_23323,N_14340,N_17758);
and U23324 (N_23324,N_13778,N_12939);
nand U23325 (N_23325,N_13374,N_13238);
nor U23326 (N_23326,N_18541,N_16340);
and U23327 (N_23327,N_18245,N_14264);
nor U23328 (N_23328,N_15829,N_13716);
or U23329 (N_23329,N_14742,N_18494);
nand U23330 (N_23330,N_16909,N_15077);
and U23331 (N_23331,N_17072,N_15467);
nor U23332 (N_23332,N_17456,N_15049);
nor U23333 (N_23333,N_15827,N_13821);
nor U23334 (N_23334,N_16444,N_16010);
nor U23335 (N_23335,N_14432,N_16658);
or U23336 (N_23336,N_18653,N_12541);
nand U23337 (N_23337,N_15541,N_17209);
and U23338 (N_23338,N_18470,N_18037);
xnor U23339 (N_23339,N_18609,N_17736);
nor U23340 (N_23340,N_16573,N_15310);
nor U23341 (N_23341,N_14670,N_13740);
nand U23342 (N_23342,N_16866,N_12642);
nor U23343 (N_23343,N_15591,N_13737);
nand U23344 (N_23344,N_12652,N_16449);
xor U23345 (N_23345,N_17793,N_15550);
or U23346 (N_23346,N_12939,N_18033);
and U23347 (N_23347,N_17731,N_14846);
and U23348 (N_23348,N_14315,N_16610);
nor U23349 (N_23349,N_15437,N_16113);
or U23350 (N_23350,N_13014,N_12889);
or U23351 (N_23351,N_18299,N_15727);
and U23352 (N_23352,N_13913,N_13784);
nor U23353 (N_23353,N_17621,N_15137);
nand U23354 (N_23354,N_17782,N_18218);
nand U23355 (N_23355,N_16765,N_18283);
or U23356 (N_23356,N_14817,N_15423);
nand U23357 (N_23357,N_18076,N_13992);
and U23358 (N_23358,N_14574,N_14900);
or U23359 (N_23359,N_18272,N_15991);
and U23360 (N_23360,N_15129,N_18476);
nand U23361 (N_23361,N_16195,N_14877);
and U23362 (N_23362,N_14006,N_15477);
nand U23363 (N_23363,N_12984,N_18563);
and U23364 (N_23364,N_16003,N_12688);
and U23365 (N_23365,N_12530,N_15551);
nor U23366 (N_23366,N_16624,N_13814);
nand U23367 (N_23367,N_13083,N_18179);
nor U23368 (N_23368,N_17920,N_17001);
or U23369 (N_23369,N_18560,N_16086);
or U23370 (N_23370,N_18364,N_15787);
or U23371 (N_23371,N_14145,N_13261);
nor U23372 (N_23372,N_17484,N_12606);
nand U23373 (N_23373,N_15769,N_15703);
xor U23374 (N_23374,N_15038,N_15413);
nor U23375 (N_23375,N_13536,N_17828);
nand U23376 (N_23376,N_16429,N_15279);
nand U23377 (N_23377,N_12678,N_15035);
nor U23378 (N_23378,N_17178,N_12561);
xor U23379 (N_23379,N_12682,N_12916);
and U23380 (N_23380,N_16622,N_15535);
nor U23381 (N_23381,N_17058,N_16750);
nor U23382 (N_23382,N_16133,N_15900);
nor U23383 (N_23383,N_13134,N_18304);
and U23384 (N_23384,N_16943,N_17220);
nand U23385 (N_23385,N_17795,N_16301);
nand U23386 (N_23386,N_12738,N_17315);
nand U23387 (N_23387,N_16005,N_14959);
or U23388 (N_23388,N_16269,N_17503);
or U23389 (N_23389,N_15449,N_15476);
xnor U23390 (N_23390,N_16695,N_13550);
and U23391 (N_23391,N_18562,N_17923);
nor U23392 (N_23392,N_13738,N_18306);
xor U23393 (N_23393,N_13606,N_13942);
and U23394 (N_23394,N_16026,N_14671);
nor U23395 (N_23395,N_17627,N_13308);
or U23396 (N_23396,N_13302,N_13452);
or U23397 (N_23397,N_14265,N_16705);
nor U23398 (N_23398,N_15156,N_18304);
nand U23399 (N_23399,N_13829,N_17087);
nand U23400 (N_23400,N_14968,N_14018);
nor U23401 (N_23401,N_15595,N_12932);
or U23402 (N_23402,N_18578,N_15023);
xnor U23403 (N_23403,N_12544,N_18263);
or U23404 (N_23404,N_15847,N_17153);
xor U23405 (N_23405,N_18728,N_15149);
nand U23406 (N_23406,N_18062,N_17201);
nand U23407 (N_23407,N_15932,N_18595);
nand U23408 (N_23408,N_12935,N_15409);
and U23409 (N_23409,N_15044,N_16860);
or U23410 (N_23410,N_18412,N_17051);
nor U23411 (N_23411,N_14589,N_16359);
nand U23412 (N_23412,N_16982,N_15956);
nor U23413 (N_23413,N_17034,N_14787);
nand U23414 (N_23414,N_16804,N_13610);
xor U23415 (N_23415,N_13564,N_12651);
or U23416 (N_23416,N_13733,N_17764);
and U23417 (N_23417,N_13554,N_17803);
xor U23418 (N_23418,N_14504,N_17621);
or U23419 (N_23419,N_12691,N_17239);
nand U23420 (N_23420,N_13474,N_15555);
nor U23421 (N_23421,N_17033,N_12621);
nor U23422 (N_23422,N_17958,N_13553);
xnor U23423 (N_23423,N_13742,N_17052);
nand U23424 (N_23424,N_13556,N_13073);
nand U23425 (N_23425,N_17980,N_17416);
and U23426 (N_23426,N_18141,N_16380);
nand U23427 (N_23427,N_14459,N_15578);
nor U23428 (N_23428,N_18242,N_17884);
or U23429 (N_23429,N_15665,N_15748);
nand U23430 (N_23430,N_13874,N_15776);
and U23431 (N_23431,N_13745,N_15303);
and U23432 (N_23432,N_18410,N_17400);
nand U23433 (N_23433,N_14772,N_13138);
nor U23434 (N_23434,N_12764,N_17772);
nor U23435 (N_23435,N_17804,N_18214);
nor U23436 (N_23436,N_16462,N_14403);
nor U23437 (N_23437,N_18676,N_18650);
or U23438 (N_23438,N_15195,N_17817);
and U23439 (N_23439,N_17703,N_16187);
nand U23440 (N_23440,N_16189,N_15592);
or U23441 (N_23441,N_16587,N_16310);
or U23442 (N_23442,N_17237,N_17008);
nor U23443 (N_23443,N_17655,N_15608);
nand U23444 (N_23444,N_18060,N_13537);
nand U23445 (N_23445,N_16177,N_14522);
and U23446 (N_23446,N_16038,N_13817);
or U23447 (N_23447,N_17829,N_12614);
and U23448 (N_23448,N_15980,N_15402);
and U23449 (N_23449,N_17219,N_17515);
nor U23450 (N_23450,N_16654,N_14068);
and U23451 (N_23451,N_16135,N_13140);
nor U23452 (N_23452,N_18740,N_13815);
and U23453 (N_23453,N_18513,N_16344);
nor U23454 (N_23454,N_15140,N_18021);
or U23455 (N_23455,N_13010,N_18424);
nand U23456 (N_23456,N_14109,N_16936);
nand U23457 (N_23457,N_17999,N_15409);
nand U23458 (N_23458,N_17750,N_14717);
nand U23459 (N_23459,N_15451,N_13781);
and U23460 (N_23460,N_12687,N_14687);
and U23461 (N_23461,N_15140,N_14539);
nor U23462 (N_23462,N_17824,N_17910);
and U23463 (N_23463,N_16616,N_15813);
or U23464 (N_23464,N_15840,N_13226);
and U23465 (N_23465,N_12654,N_18241);
or U23466 (N_23466,N_15660,N_12660);
or U23467 (N_23467,N_13000,N_14573);
nor U23468 (N_23468,N_13468,N_14314);
nor U23469 (N_23469,N_14676,N_14180);
xor U23470 (N_23470,N_12836,N_16022);
and U23471 (N_23471,N_14343,N_18130);
nand U23472 (N_23472,N_16661,N_18200);
nand U23473 (N_23473,N_12873,N_14506);
nor U23474 (N_23474,N_17822,N_15497);
nand U23475 (N_23475,N_15063,N_18321);
xnor U23476 (N_23476,N_12582,N_13085);
nand U23477 (N_23477,N_16751,N_14802);
or U23478 (N_23478,N_16692,N_17078);
nor U23479 (N_23479,N_17166,N_14367);
and U23480 (N_23480,N_15029,N_14464);
nor U23481 (N_23481,N_17596,N_14879);
nand U23482 (N_23482,N_13905,N_12791);
nor U23483 (N_23483,N_12897,N_13273);
nand U23484 (N_23484,N_18644,N_16096);
and U23485 (N_23485,N_17623,N_15828);
nor U23486 (N_23486,N_14143,N_17454);
and U23487 (N_23487,N_18427,N_13474);
nor U23488 (N_23488,N_16378,N_17675);
and U23489 (N_23489,N_14741,N_17673);
nor U23490 (N_23490,N_14898,N_15509);
or U23491 (N_23491,N_14336,N_15597);
and U23492 (N_23492,N_18039,N_14030);
nor U23493 (N_23493,N_15581,N_12595);
or U23494 (N_23494,N_14782,N_16229);
nor U23495 (N_23495,N_17308,N_15584);
nor U23496 (N_23496,N_17862,N_13056);
nor U23497 (N_23497,N_17140,N_12856);
or U23498 (N_23498,N_15948,N_13635);
nor U23499 (N_23499,N_16116,N_14723);
nor U23500 (N_23500,N_14190,N_17253);
or U23501 (N_23501,N_14984,N_15325);
and U23502 (N_23502,N_16446,N_12541);
nand U23503 (N_23503,N_15353,N_17681);
nand U23504 (N_23504,N_17315,N_16199);
and U23505 (N_23505,N_18670,N_16515);
nand U23506 (N_23506,N_16927,N_17271);
and U23507 (N_23507,N_16480,N_17768);
and U23508 (N_23508,N_17949,N_14728);
xnor U23509 (N_23509,N_18295,N_15570);
nor U23510 (N_23510,N_13845,N_15056);
and U23511 (N_23511,N_14206,N_15776);
nand U23512 (N_23512,N_12977,N_14623);
or U23513 (N_23513,N_16218,N_17034);
nand U23514 (N_23514,N_18013,N_17169);
or U23515 (N_23515,N_16190,N_13515);
nand U23516 (N_23516,N_15244,N_14336);
nor U23517 (N_23517,N_13025,N_17421);
or U23518 (N_23518,N_15431,N_13792);
or U23519 (N_23519,N_13097,N_12812);
nor U23520 (N_23520,N_13274,N_15033);
xnor U23521 (N_23521,N_12929,N_17733);
and U23522 (N_23522,N_18532,N_16939);
and U23523 (N_23523,N_12688,N_18249);
and U23524 (N_23524,N_17948,N_16814);
nor U23525 (N_23525,N_17815,N_16372);
and U23526 (N_23526,N_16751,N_17234);
nand U23527 (N_23527,N_14298,N_13008);
or U23528 (N_23528,N_13324,N_13875);
xor U23529 (N_23529,N_13660,N_13996);
and U23530 (N_23530,N_14618,N_15158);
nand U23531 (N_23531,N_14210,N_17244);
nor U23532 (N_23532,N_14174,N_13158);
and U23533 (N_23533,N_14738,N_17665);
nand U23534 (N_23534,N_14469,N_18070);
and U23535 (N_23535,N_18468,N_13465);
nor U23536 (N_23536,N_15479,N_12699);
or U23537 (N_23537,N_17261,N_16372);
or U23538 (N_23538,N_16462,N_12824);
and U23539 (N_23539,N_14587,N_18027);
or U23540 (N_23540,N_16431,N_15100);
and U23541 (N_23541,N_13233,N_17734);
nand U23542 (N_23542,N_15940,N_13214);
nand U23543 (N_23543,N_12826,N_13032);
nand U23544 (N_23544,N_12633,N_14810);
nand U23545 (N_23545,N_14766,N_17225);
or U23546 (N_23546,N_14412,N_13474);
nand U23547 (N_23547,N_13935,N_17291);
nand U23548 (N_23548,N_13520,N_16243);
or U23549 (N_23549,N_12594,N_17223);
nor U23550 (N_23550,N_12969,N_18195);
or U23551 (N_23551,N_14065,N_16484);
or U23552 (N_23552,N_13590,N_17685);
nor U23553 (N_23553,N_14992,N_17290);
nand U23554 (N_23554,N_13165,N_13009);
nor U23555 (N_23555,N_18326,N_17987);
and U23556 (N_23556,N_17046,N_14161);
and U23557 (N_23557,N_17743,N_12646);
nor U23558 (N_23558,N_14321,N_17911);
and U23559 (N_23559,N_18294,N_14398);
xnor U23560 (N_23560,N_17050,N_17039);
nand U23561 (N_23561,N_14001,N_15571);
and U23562 (N_23562,N_16811,N_17015);
or U23563 (N_23563,N_13512,N_16736);
or U23564 (N_23564,N_16832,N_12839);
or U23565 (N_23565,N_17756,N_12873);
and U23566 (N_23566,N_18160,N_16724);
nand U23567 (N_23567,N_17203,N_14476);
nor U23568 (N_23568,N_13261,N_15525);
nor U23569 (N_23569,N_15418,N_17289);
nor U23570 (N_23570,N_17785,N_12789);
nor U23571 (N_23571,N_13873,N_16023);
nand U23572 (N_23572,N_17075,N_16926);
or U23573 (N_23573,N_16694,N_13683);
nand U23574 (N_23574,N_18554,N_15497);
and U23575 (N_23575,N_14869,N_15543);
nor U23576 (N_23576,N_15160,N_13054);
nor U23577 (N_23577,N_15490,N_15157);
nand U23578 (N_23578,N_17838,N_13909);
nor U23579 (N_23579,N_14087,N_18492);
xnor U23580 (N_23580,N_15697,N_12645);
nand U23581 (N_23581,N_15033,N_15288);
nand U23582 (N_23582,N_17493,N_12624);
and U23583 (N_23583,N_14917,N_17641);
nor U23584 (N_23584,N_17907,N_16278);
nand U23585 (N_23585,N_16635,N_18350);
and U23586 (N_23586,N_12711,N_12722);
nand U23587 (N_23587,N_17313,N_15428);
and U23588 (N_23588,N_15746,N_15232);
nor U23589 (N_23589,N_13666,N_17997);
nor U23590 (N_23590,N_18208,N_16630);
nor U23591 (N_23591,N_16797,N_17537);
nand U23592 (N_23592,N_13881,N_13920);
xnor U23593 (N_23593,N_17341,N_18481);
nor U23594 (N_23594,N_14459,N_14604);
and U23595 (N_23595,N_17575,N_17270);
nand U23596 (N_23596,N_12970,N_15962);
nor U23597 (N_23597,N_16644,N_15465);
nor U23598 (N_23598,N_17415,N_15659);
nand U23599 (N_23599,N_14423,N_16592);
and U23600 (N_23600,N_16913,N_13991);
xor U23601 (N_23601,N_16859,N_16921);
nor U23602 (N_23602,N_15980,N_15933);
and U23603 (N_23603,N_16212,N_14851);
nor U23604 (N_23604,N_17144,N_18540);
nand U23605 (N_23605,N_17362,N_12716);
or U23606 (N_23606,N_13566,N_15154);
nor U23607 (N_23607,N_12863,N_18612);
nor U23608 (N_23608,N_13763,N_14403);
or U23609 (N_23609,N_17662,N_18503);
or U23610 (N_23610,N_12817,N_16207);
and U23611 (N_23611,N_14560,N_14779);
nand U23612 (N_23612,N_16610,N_17063);
or U23613 (N_23613,N_15651,N_13515);
xnor U23614 (N_23614,N_13866,N_16004);
nand U23615 (N_23615,N_18594,N_16046);
nand U23616 (N_23616,N_18109,N_13936);
and U23617 (N_23617,N_15206,N_16724);
and U23618 (N_23618,N_16129,N_17738);
nand U23619 (N_23619,N_13286,N_15926);
or U23620 (N_23620,N_15900,N_14809);
xnor U23621 (N_23621,N_16496,N_15287);
or U23622 (N_23622,N_16402,N_18351);
nand U23623 (N_23623,N_13029,N_14583);
or U23624 (N_23624,N_16318,N_16348);
xor U23625 (N_23625,N_14536,N_17858);
or U23626 (N_23626,N_17438,N_13551);
xor U23627 (N_23627,N_18562,N_16244);
or U23628 (N_23628,N_17686,N_17594);
nand U23629 (N_23629,N_13443,N_15089);
nand U23630 (N_23630,N_18499,N_13301);
nor U23631 (N_23631,N_16963,N_12800);
nand U23632 (N_23632,N_14719,N_13976);
nor U23633 (N_23633,N_16431,N_12883);
nand U23634 (N_23634,N_18419,N_16617);
xnor U23635 (N_23635,N_16621,N_13887);
xor U23636 (N_23636,N_12566,N_12571);
or U23637 (N_23637,N_14775,N_13456);
nand U23638 (N_23638,N_14828,N_12905);
or U23639 (N_23639,N_17633,N_14660);
xnor U23640 (N_23640,N_16778,N_14395);
nand U23641 (N_23641,N_15449,N_15639);
or U23642 (N_23642,N_17269,N_13822);
nor U23643 (N_23643,N_13152,N_13183);
nand U23644 (N_23644,N_16160,N_16336);
nand U23645 (N_23645,N_14615,N_16856);
nand U23646 (N_23646,N_13004,N_15177);
or U23647 (N_23647,N_15640,N_14065);
xnor U23648 (N_23648,N_15296,N_15051);
xnor U23649 (N_23649,N_13653,N_16292);
or U23650 (N_23650,N_17744,N_14605);
nand U23651 (N_23651,N_16232,N_17084);
or U23652 (N_23652,N_13013,N_17619);
nand U23653 (N_23653,N_14205,N_15639);
and U23654 (N_23654,N_14849,N_15975);
and U23655 (N_23655,N_14604,N_14257);
nand U23656 (N_23656,N_14865,N_13223);
xor U23657 (N_23657,N_13987,N_13148);
or U23658 (N_23658,N_12552,N_17248);
and U23659 (N_23659,N_17670,N_14703);
or U23660 (N_23660,N_18261,N_13885);
or U23661 (N_23661,N_16735,N_14172);
nand U23662 (N_23662,N_15877,N_18323);
or U23663 (N_23663,N_13906,N_14496);
or U23664 (N_23664,N_18675,N_16516);
nor U23665 (N_23665,N_16080,N_16069);
nor U23666 (N_23666,N_12565,N_13951);
or U23667 (N_23667,N_17678,N_17336);
nand U23668 (N_23668,N_14694,N_17458);
nor U23669 (N_23669,N_15134,N_14514);
and U23670 (N_23670,N_14816,N_16478);
nor U23671 (N_23671,N_13896,N_16614);
and U23672 (N_23672,N_15120,N_17304);
or U23673 (N_23673,N_13969,N_14691);
nor U23674 (N_23674,N_13689,N_15727);
or U23675 (N_23675,N_13676,N_12993);
and U23676 (N_23676,N_18685,N_14887);
or U23677 (N_23677,N_17746,N_12859);
nor U23678 (N_23678,N_14255,N_13593);
nand U23679 (N_23679,N_14249,N_12605);
xnor U23680 (N_23680,N_16658,N_15503);
or U23681 (N_23681,N_15195,N_18395);
nand U23682 (N_23682,N_16098,N_13837);
or U23683 (N_23683,N_16138,N_16562);
and U23684 (N_23684,N_15745,N_14010);
nand U23685 (N_23685,N_17518,N_14666);
xor U23686 (N_23686,N_16192,N_13658);
and U23687 (N_23687,N_14799,N_15754);
and U23688 (N_23688,N_17976,N_16449);
nor U23689 (N_23689,N_18337,N_14980);
and U23690 (N_23690,N_16143,N_18531);
nand U23691 (N_23691,N_16553,N_14812);
and U23692 (N_23692,N_17005,N_18532);
or U23693 (N_23693,N_13586,N_13531);
nand U23694 (N_23694,N_16269,N_14908);
xor U23695 (N_23695,N_18103,N_17159);
and U23696 (N_23696,N_13814,N_14191);
xnor U23697 (N_23697,N_12524,N_18409);
nor U23698 (N_23698,N_16748,N_17278);
and U23699 (N_23699,N_13671,N_12717);
or U23700 (N_23700,N_18632,N_15925);
and U23701 (N_23701,N_16771,N_12628);
nor U23702 (N_23702,N_13625,N_18739);
and U23703 (N_23703,N_13243,N_12808);
nor U23704 (N_23704,N_15874,N_16475);
or U23705 (N_23705,N_14611,N_13711);
or U23706 (N_23706,N_17364,N_16956);
or U23707 (N_23707,N_15964,N_12966);
and U23708 (N_23708,N_15444,N_16482);
nor U23709 (N_23709,N_17548,N_12557);
nor U23710 (N_23710,N_13854,N_17849);
xor U23711 (N_23711,N_14515,N_15144);
and U23712 (N_23712,N_17382,N_13274);
nor U23713 (N_23713,N_13612,N_16684);
nand U23714 (N_23714,N_15229,N_15313);
or U23715 (N_23715,N_15962,N_16100);
or U23716 (N_23716,N_15773,N_17697);
or U23717 (N_23717,N_16150,N_18333);
nand U23718 (N_23718,N_15650,N_14268);
nand U23719 (N_23719,N_14619,N_18069);
xnor U23720 (N_23720,N_12590,N_12746);
nor U23721 (N_23721,N_18111,N_14299);
and U23722 (N_23722,N_18693,N_15146);
nand U23723 (N_23723,N_14872,N_13706);
or U23724 (N_23724,N_17575,N_13202);
xor U23725 (N_23725,N_17997,N_14795);
nor U23726 (N_23726,N_14609,N_16910);
nor U23727 (N_23727,N_16928,N_12733);
nand U23728 (N_23728,N_15245,N_17049);
and U23729 (N_23729,N_12894,N_13855);
nand U23730 (N_23730,N_17500,N_16016);
or U23731 (N_23731,N_15942,N_14116);
nor U23732 (N_23732,N_14657,N_15554);
nand U23733 (N_23733,N_16052,N_17631);
or U23734 (N_23734,N_14141,N_13903);
and U23735 (N_23735,N_15515,N_17680);
or U23736 (N_23736,N_15382,N_16476);
or U23737 (N_23737,N_16376,N_18377);
xor U23738 (N_23738,N_18734,N_15271);
xnor U23739 (N_23739,N_16982,N_17058);
and U23740 (N_23740,N_17419,N_15181);
or U23741 (N_23741,N_15954,N_16761);
nand U23742 (N_23742,N_14442,N_18299);
and U23743 (N_23743,N_13989,N_18039);
nor U23744 (N_23744,N_18106,N_13073);
nand U23745 (N_23745,N_17319,N_14598);
nor U23746 (N_23746,N_15775,N_13179);
nand U23747 (N_23747,N_15242,N_13355);
or U23748 (N_23748,N_16635,N_18164);
nand U23749 (N_23749,N_18720,N_17925);
or U23750 (N_23750,N_17448,N_18294);
xnor U23751 (N_23751,N_12746,N_17678);
and U23752 (N_23752,N_13900,N_14313);
or U23753 (N_23753,N_17530,N_15297);
nand U23754 (N_23754,N_12960,N_16879);
nand U23755 (N_23755,N_16114,N_17058);
nand U23756 (N_23756,N_17072,N_12983);
or U23757 (N_23757,N_15716,N_14041);
nor U23758 (N_23758,N_13195,N_15339);
nor U23759 (N_23759,N_13960,N_16695);
and U23760 (N_23760,N_18418,N_17031);
nand U23761 (N_23761,N_18195,N_18419);
and U23762 (N_23762,N_16839,N_15851);
nand U23763 (N_23763,N_15350,N_17346);
nand U23764 (N_23764,N_17964,N_14530);
nor U23765 (N_23765,N_13302,N_14083);
or U23766 (N_23766,N_16144,N_14903);
nand U23767 (N_23767,N_17110,N_17792);
or U23768 (N_23768,N_12587,N_14702);
nand U23769 (N_23769,N_15987,N_16455);
nand U23770 (N_23770,N_13108,N_17881);
nor U23771 (N_23771,N_14308,N_14200);
nand U23772 (N_23772,N_17559,N_14279);
and U23773 (N_23773,N_16486,N_17592);
nor U23774 (N_23774,N_14772,N_14679);
nor U23775 (N_23775,N_13579,N_13050);
and U23776 (N_23776,N_16920,N_16784);
nand U23777 (N_23777,N_15316,N_16104);
or U23778 (N_23778,N_13319,N_13736);
nand U23779 (N_23779,N_18341,N_13787);
xnor U23780 (N_23780,N_16732,N_16286);
xor U23781 (N_23781,N_13051,N_16494);
nand U23782 (N_23782,N_17125,N_17545);
nor U23783 (N_23783,N_18622,N_17949);
xnor U23784 (N_23784,N_14739,N_13149);
nor U23785 (N_23785,N_17586,N_15707);
and U23786 (N_23786,N_15239,N_15103);
nand U23787 (N_23787,N_14571,N_14057);
or U23788 (N_23788,N_17115,N_16727);
and U23789 (N_23789,N_18059,N_17807);
xnor U23790 (N_23790,N_15482,N_18192);
or U23791 (N_23791,N_14874,N_17549);
xnor U23792 (N_23792,N_14138,N_16230);
and U23793 (N_23793,N_17649,N_18388);
nor U23794 (N_23794,N_15805,N_18289);
nor U23795 (N_23795,N_13762,N_17989);
or U23796 (N_23796,N_16707,N_16929);
nand U23797 (N_23797,N_12897,N_14263);
xnor U23798 (N_23798,N_14780,N_18710);
or U23799 (N_23799,N_14538,N_16375);
or U23800 (N_23800,N_17625,N_16617);
nand U23801 (N_23801,N_15529,N_14738);
and U23802 (N_23802,N_17041,N_17135);
nand U23803 (N_23803,N_14348,N_16123);
xnor U23804 (N_23804,N_15368,N_13289);
or U23805 (N_23805,N_17679,N_13844);
or U23806 (N_23806,N_16379,N_15647);
xor U23807 (N_23807,N_14874,N_13826);
xnor U23808 (N_23808,N_16753,N_14768);
nand U23809 (N_23809,N_17325,N_17598);
xor U23810 (N_23810,N_15516,N_18323);
and U23811 (N_23811,N_13025,N_13990);
or U23812 (N_23812,N_18095,N_18167);
or U23813 (N_23813,N_15269,N_15918);
nor U23814 (N_23814,N_15762,N_16952);
nor U23815 (N_23815,N_17268,N_16449);
xnor U23816 (N_23816,N_16749,N_16438);
nand U23817 (N_23817,N_15015,N_12935);
xnor U23818 (N_23818,N_13044,N_18669);
or U23819 (N_23819,N_16716,N_17394);
and U23820 (N_23820,N_14161,N_16562);
nand U23821 (N_23821,N_13395,N_14926);
or U23822 (N_23822,N_13450,N_15281);
or U23823 (N_23823,N_15248,N_15222);
or U23824 (N_23824,N_15799,N_18308);
and U23825 (N_23825,N_18403,N_18009);
and U23826 (N_23826,N_15210,N_13936);
xor U23827 (N_23827,N_16456,N_17755);
and U23828 (N_23828,N_14820,N_15975);
nor U23829 (N_23829,N_18538,N_17907);
or U23830 (N_23830,N_12563,N_17623);
or U23831 (N_23831,N_16412,N_18159);
xnor U23832 (N_23832,N_18013,N_18668);
or U23833 (N_23833,N_16248,N_16431);
xnor U23834 (N_23834,N_17524,N_17223);
nand U23835 (N_23835,N_17690,N_15226);
nand U23836 (N_23836,N_13059,N_13533);
and U23837 (N_23837,N_15037,N_17000);
nand U23838 (N_23838,N_13278,N_15748);
and U23839 (N_23839,N_17552,N_12545);
nand U23840 (N_23840,N_14734,N_14892);
nor U23841 (N_23841,N_15386,N_18310);
or U23842 (N_23842,N_17696,N_13478);
or U23843 (N_23843,N_14182,N_17406);
or U23844 (N_23844,N_15253,N_15991);
nand U23845 (N_23845,N_14286,N_16157);
or U23846 (N_23846,N_13714,N_15835);
nand U23847 (N_23847,N_14718,N_15144);
and U23848 (N_23848,N_17707,N_13908);
nor U23849 (N_23849,N_15951,N_16879);
and U23850 (N_23850,N_17540,N_17315);
nand U23851 (N_23851,N_16030,N_15361);
or U23852 (N_23852,N_18441,N_17405);
or U23853 (N_23853,N_16916,N_13885);
or U23854 (N_23854,N_13650,N_14278);
nand U23855 (N_23855,N_16607,N_13146);
and U23856 (N_23856,N_17832,N_18702);
or U23857 (N_23857,N_14842,N_15300);
nand U23858 (N_23858,N_15774,N_17260);
nor U23859 (N_23859,N_13267,N_17074);
nor U23860 (N_23860,N_18337,N_12870);
and U23861 (N_23861,N_13258,N_14199);
nor U23862 (N_23862,N_18309,N_17895);
nand U23863 (N_23863,N_17965,N_18616);
and U23864 (N_23864,N_14936,N_17100);
or U23865 (N_23865,N_15139,N_12522);
xnor U23866 (N_23866,N_13879,N_14503);
nand U23867 (N_23867,N_15846,N_13995);
or U23868 (N_23868,N_17084,N_13093);
and U23869 (N_23869,N_15689,N_18435);
and U23870 (N_23870,N_14290,N_12600);
nand U23871 (N_23871,N_16257,N_16139);
or U23872 (N_23872,N_18324,N_18271);
xnor U23873 (N_23873,N_18237,N_13534);
nand U23874 (N_23874,N_17880,N_14227);
nor U23875 (N_23875,N_16392,N_15079);
xnor U23876 (N_23876,N_13009,N_15899);
or U23877 (N_23877,N_13578,N_13883);
or U23878 (N_23878,N_12688,N_14885);
xor U23879 (N_23879,N_18361,N_15320);
xnor U23880 (N_23880,N_17888,N_14295);
or U23881 (N_23881,N_16312,N_13529);
or U23882 (N_23882,N_14594,N_18696);
or U23883 (N_23883,N_14941,N_16880);
and U23884 (N_23884,N_12953,N_12545);
nand U23885 (N_23885,N_14764,N_17192);
nor U23886 (N_23886,N_15446,N_16026);
or U23887 (N_23887,N_15371,N_18649);
and U23888 (N_23888,N_14519,N_13659);
nand U23889 (N_23889,N_13919,N_17668);
or U23890 (N_23890,N_14197,N_18413);
nand U23891 (N_23891,N_14202,N_15233);
nand U23892 (N_23892,N_13527,N_18075);
xor U23893 (N_23893,N_17121,N_17812);
or U23894 (N_23894,N_18221,N_12580);
nor U23895 (N_23895,N_17604,N_15387);
and U23896 (N_23896,N_14540,N_17273);
nor U23897 (N_23897,N_12790,N_18615);
nor U23898 (N_23898,N_16994,N_16659);
or U23899 (N_23899,N_14362,N_15546);
and U23900 (N_23900,N_14312,N_17227);
or U23901 (N_23901,N_17937,N_15834);
xnor U23902 (N_23902,N_18739,N_14824);
or U23903 (N_23903,N_14119,N_15784);
nor U23904 (N_23904,N_13834,N_15557);
nor U23905 (N_23905,N_15065,N_12600);
nand U23906 (N_23906,N_17879,N_14431);
and U23907 (N_23907,N_17211,N_16518);
and U23908 (N_23908,N_14998,N_18276);
or U23909 (N_23909,N_13107,N_18572);
and U23910 (N_23910,N_18679,N_12776);
nand U23911 (N_23911,N_17190,N_14938);
or U23912 (N_23912,N_13758,N_17415);
xnor U23913 (N_23913,N_17612,N_18385);
nand U23914 (N_23914,N_14220,N_13462);
nand U23915 (N_23915,N_18528,N_16246);
nand U23916 (N_23916,N_14411,N_13764);
xnor U23917 (N_23917,N_13665,N_16446);
or U23918 (N_23918,N_14305,N_18703);
nor U23919 (N_23919,N_15208,N_16720);
or U23920 (N_23920,N_17473,N_14278);
or U23921 (N_23921,N_14924,N_18076);
xor U23922 (N_23922,N_16349,N_18636);
nand U23923 (N_23923,N_16949,N_18215);
nor U23924 (N_23924,N_15188,N_12961);
and U23925 (N_23925,N_14686,N_14778);
or U23926 (N_23926,N_17185,N_13731);
nand U23927 (N_23927,N_13341,N_15840);
nor U23928 (N_23928,N_13421,N_14082);
nor U23929 (N_23929,N_15001,N_16519);
nor U23930 (N_23930,N_17363,N_13504);
nand U23931 (N_23931,N_16361,N_18361);
nand U23932 (N_23932,N_17892,N_12841);
nand U23933 (N_23933,N_12950,N_13964);
nor U23934 (N_23934,N_16854,N_14231);
or U23935 (N_23935,N_15073,N_18678);
nor U23936 (N_23936,N_15113,N_18218);
and U23937 (N_23937,N_15525,N_13493);
nand U23938 (N_23938,N_12571,N_13279);
nand U23939 (N_23939,N_17685,N_17690);
or U23940 (N_23940,N_16300,N_17166);
or U23941 (N_23941,N_14220,N_13557);
and U23942 (N_23942,N_12830,N_12816);
nor U23943 (N_23943,N_16584,N_18522);
or U23944 (N_23944,N_17141,N_15440);
and U23945 (N_23945,N_13013,N_15471);
nor U23946 (N_23946,N_15326,N_15224);
nor U23947 (N_23947,N_15872,N_13654);
nand U23948 (N_23948,N_15750,N_15969);
xnor U23949 (N_23949,N_13712,N_15586);
nand U23950 (N_23950,N_13455,N_18629);
or U23951 (N_23951,N_16599,N_12591);
and U23952 (N_23952,N_15722,N_18709);
nand U23953 (N_23953,N_14363,N_16927);
or U23954 (N_23954,N_13955,N_17336);
nor U23955 (N_23955,N_15122,N_18507);
nor U23956 (N_23956,N_14758,N_18507);
or U23957 (N_23957,N_16872,N_17821);
and U23958 (N_23958,N_18390,N_13510);
or U23959 (N_23959,N_15608,N_17095);
and U23960 (N_23960,N_15296,N_13390);
nand U23961 (N_23961,N_13268,N_12980);
or U23962 (N_23962,N_17773,N_18705);
nand U23963 (N_23963,N_12827,N_17770);
and U23964 (N_23964,N_15982,N_15946);
or U23965 (N_23965,N_14353,N_13142);
or U23966 (N_23966,N_12771,N_12650);
and U23967 (N_23967,N_12738,N_16262);
nor U23968 (N_23968,N_14781,N_16479);
and U23969 (N_23969,N_16166,N_13480);
or U23970 (N_23970,N_16568,N_12728);
or U23971 (N_23971,N_17699,N_15229);
nand U23972 (N_23972,N_12640,N_13380);
nor U23973 (N_23973,N_16978,N_12823);
nand U23974 (N_23974,N_17411,N_14464);
nor U23975 (N_23975,N_18164,N_14389);
nand U23976 (N_23976,N_15371,N_17913);
nor U23977 (N_23977,N_15870,N_15987);
nand U23978 (N_23978,N_15959,N_17496);
nand U23979 (N_23979,N_14893,N_14474);
nor U23980 (N_23980,N_13158,N_13537);
nand U23981 (N_23981,N_16414,N_14647);
nor U23982 (N_23982,N_16662,N_18074);
nor U23983 (N_23983,N_14366,N_16058);
nand U23984 (N_23984,N_14509,N_13079);
nand U23985 (N_23985,N_16366,N_15234);
and U23986 (N_23986,N_14740,N_14551);
and U23987 (N_23987,N_13026,N_13649);
or U23988 (N_23988,N_15431,N_15212);
nand U23989 (N_23989,N_15884,N_14677);
xnor U23990 (N_23990,N_16521,N_14228);
nand U23991 (N_23991,N_14611,N_14724);
or U23992 (N_23992,N_16818,N_17073);
and U23993 (N_23993,N_13560,N_15902);
nand U23994 (N_23994,N_12638,N_18456);
or U23995 (N_23995,N_15708,N_15935);
nor U23996 (N_23996,N_15009,N_12553);
xnor U23997 (N_23997,N_15240,N_14054);
and U23998 (N_23998,N_16836,N_18429);
xor U23999 (N_23999,N_13599,N_16921);
nand U24000 (N_24000,N_13382,N_17887);
nand U24001 (N_24001,N_16141,N_15582);
or U24002 (N_24002,N_14206,N_17682);
nor U24003 (N_24003,N_13993,N_18120);
nor U24004 (N_24004,N_18156,N_12764);
nor U24005 (N_24005,N_15878,N_14071);
or U24006 (N_24006,N_18668,N_16744);
or U24007 (N_24007,N_17632,N_15925);
and U24008 (N_24008,N_14929,N_18622);
and U24009 (N_24009,N_12888,N_12607);
and U24010 (N_24010,N_17024,N_15960);
or U24011 (N_24011,N_13115,N_12945);
or U24012 (N_24012,N_16531,N_17670);
or U24013 (N_24013,N_18159,N_13426);
and U24014 (N_24014,N_14153,N_15635);
nand U24015 (N_24015,N_15944,N_16577);
or U24016 (N_24016,N_18629,N_16770);
nand U24017 (N_24017,N_15539,N_15877);
or U24018 (N_24018,N_16161,N_14711);
xor U24019 (N_24019,N_17266,N_14104);
and U24020 (N_24020,N_16926,N_18370);
nand U24021 (N_24021,N_12842,N_17187);
nand U24022 (N_24022,N_15114,N_16822);
or U24023 (N_24023,N_17393,N_17952);
or U24024 (N_24024,N_14584,N_17700);
nor U24025 (N_24025,N_16075,N_15395);
nand U24026 (N_24026,N_14641,N_17057);
xnor U24027 (N_24027,N_16165,N_18679);
and U24028 (N_24028,N_13739,N_16213);
and U24029 (N_24029,N_15276,N_15246);
or U24030 (N_24030,N_15319,N_15099);
nor U24031 (N_24031,N_17898,N_14043);
or U24032 (N_24032,N_17195,N_14126);
xnor U24033 (N_24033,N_16150,N_13517);
or U24034 (N_24034,N_18049,N_14389);
and U24035 (N_24035,N_16497,N_18007);
nand U24036 (N_24036,N_15867,N_13915);
nor U24037 (N_24037,N_16237,N_18140);
xnor U24038 (N_24038,N_18659,N_17756);
nand U24039 (N_24039,N_15234,N_17212);
nand U24040 (N_24040,N_14290,N_18682);
or U24041 (N_24041,N_17690,N_15150);
or U24042 (N_24042,N_15500,N_17407);
or U24043 (N_24043,N_17737,N_15952);
or U24044 (N_24044,N_16174,N_15682);
nor U24045 (N_24045,N_16020,N_15472);
and U24046 (N_24046,N_13299,N_13219);
xor U24047 (N_24047,N_13152,N_17685);
or U24048 (N_24048,N_18591,N_12901);
nand U24049 (N_24049,N_13578,N_14557);
nand U24050 (N_24050,N_13031,N_15550);
nand U24051 (N_24051,N_13510,N_15015);
and U24052 (N_24052,N_15624,N_12986);
nor U24053 (N_24053,N_16928,N_13670);
nand U24054 (N_24054,N_17061,N_17067);
nor U24055 (N_24055,N_13919,N_15245);
and U24056 (N_24056,N_12834,N_13825);
xnor U24057 (N_24057,N_14071,N_15704);
or U24058 (N_24058,N_18303,N_18440);
nand U24059 (N_24059,N_13042,N_13390);
or U24060 (N_24060,N_13811,N_13432);
nand U24061 (N_24061,N_13841,N_17408);
nand U24062 (N_24062,N_13548,N_18412);
nand U24063 (N_24063,N_12982,N_17245);
nand U24064 (N_24064,N_17549,N_13487);
and U24065 (N_24065,N_14261,N_16734);
nand U24066 (N_24066,N_16779,N_13868);
nor U24067 (N_24067,N_14037,N_16137);
or U24068 (N_24068,N_14886,N_14282);
nand U24069 (N_24069,N_14025,N_16569);
or U24070 (N_24070,N_17945,N_15166);
and U24071 (N_24071,N_16173,N_18289);
nor U24072 (N_24072,N_16329,N_18217);
nand U24073 (N_24073,N_17732,N_13123);
xnor U24074 (N_24074,N_15288,N_18147);
nor U24075 (N_24075,N_17528,N_17456);
or U24076 (N_24076,N_15263,N_14951);
nand U24077 (N_24077,N_14387,N_15023);
nand U24078 (N_24078,N_15975,N_12767);
and U24079 (N_24079,N_15393,N_14445);
or U24080 (N_24080,N_13933,N_18153);
nand U24081 (N_24081,N_16250,N_16353);
nor U24082 (N_24082,N_16137,N_14010);
nand U24083 (N_24083,N_16805,N_17756);
nor U24084 (N_24084,N_13667,N_17156);
or U24085 (N_24085,N_15900,N_12625);
xor U24086 (N_24086,N_14434,N_15105);
nor U24087 (N_24087,N_17003,N_16284);
nand U24088 (N_24088,N_13243,N_13407);
and U24089 (N_24089,N_17573,N_15616);
and U24090 (N_24090,N_13471,N_18336);
nand U24091 (N_24091,N_13892,N_14494);
nand U24092 (N_24092,N_12550,N_17170);
nor U24093 (N_24093,N_17540,N_14608);
nand U24094 (N_24094,N_12851,N_15874);
nand U24095 (N_24095,N_15226,N_16551);
and U24096 (N_24096,N_13192,N_15674);
nor U24097 (N_24097,N_13998,N_15115);
nor U24098 (N_24098,N_14183,N_13820);
xor U24099 (N_24099,N_12784,N_16634);
nand U24100 (N_24100,N_16209,N_16374);
xor U24101 (N_24101,N_17599,N_18593);
and U24102 (N_24102,N_12664,N_14437);
nand U24103 (N_24103,N_16841,N_14673);
and U24104 (N_24104,N_18233,N_15755);
and U24105 (N_24105,N_15522,N_13621);
nand U24106 (N_24106,N_17769,N_17925);
or U24107 (N_24107,N_17154,N_16823);
and U24108 (N_24108,N_18749,N_15305);
nand U24109 (N_24109,N_14216,N_14170);
or U24110 (N_24110,N_14482,N_16405);
nor U24111 (N_24111,N_18548,N_14469);
nor U24112 (N_24112,N_18488,N_15975);
nor U24113 (N_24113,N_13759,N_17094);
nand U24114 (N_24114,N_12506,N_16443);
or U24115 (N_24115,N_16508,N_18474);
or U24116 (N_24116,N_18495,N_14276);
nor U24117 (N_24117,N_15802,N_18374);
or U24118 (N_24118,N_14651,N_13992);
xnor U24119 (N_24119,N_14789,N_13784);
xor U24120 (N_24120,N_13313,N_16484);
or U24121 (N_24121,N_13599,N_14901);
nand U24122 (N_24122,N_13687,N_16778);
xor U24123 (N_24123,N_14660,N_14516);
or U24124 (N_24124,N_14226,N_15746);
and U24125 (N_24125,N_18616,N_12511);
xor U24126 (N_24126,N_13166,N_17151);
nand U24127 (N_24127,N_16897,N_18363);
and U24128 (N_24128,N_14679,N_13423);
nand U24129 (N_24129,N_13001,N_16958);
xnor U24130 (N_24130,N_16225,N_14151);
or U24131 (N_24131,N_14443,N_15709);
nor U24132 (N_24132,N_18573,N_13097);
nor U24133 (N_24133,N_16205,N_15504);
and U24134 (N_24134,N_13333,N_13053);
and U24135 (N_24135,N_16751,N_17359);
xor U24136 (N_24136,N_17062,N_17183);
xor U24137 (N_24137,N_16270,N_16057);
and U24138 (N_24138,N_16589,N_13978);
nand U24139 (N_24139,N_13729,N_14441);
and U24140 (N_24140,N_13843,N_15066);
or U24141 (N_24141,N_16136,N_13198);
xnor U24142 (N_24142,N_15638,N_12822);
or U24143 (N_24143,N_15111,N_13442);
nor U24144 (N_24144,N_14050,N_13780);
xor U24145 (N_24145,N_16966,N_16852);
nand U24146 (N_24146,N_13369,N_13875);
and U24147 (N_24147,N_13782,N_12836);
nand U24148 (N_24148,N_17233,N_17627);
nand U24149 (N_24149,N_15814,N_13473);
nand U24150 (N_24150,N_18024,N_17827);
or U24151 (N_24151,N_13694,N_13583);
nand U24152 (N_24152,N_15621,N_17932);
nand U24153 (N_24153,N_13863,N_16810);
nor U24154 (N_24154,N_13176,N_15196);
and U24155 (N_24155,N_12650,N_15405);
and U24156 (N_24156,N_13116,N_18417);
nand U24157 (N_24157,N_17330,N_14999);
nor U24158 (N_24158,N_14925,N_15367);
or U24159 (N_24159,N_16528,N_14847);
or U24160 (N_24160,N_15358,N_14833);
nor U24161 (N_24161,N_15513,N_16711);
nor U24162 (N_24162,N_17230,N_16958);
or U24163 (N_24163,N_13134,N_18420);
or U24164 (N_24164,N_15286,N_16531);
nor U24165 (N_24165,N_14513,N_15159);
nor U24166 (N_24166,N_17097,N_12524);
nand U24167 (N_24167,N_13885,N_16596);
nor U24168 (N_24168,N_16026,N_16669);
or U24169 (N_24169,N_15066,N_18333);
or U24170 (N_24170,N_13649,N_15704);
nand U24171 (N_24171,N_17470,N_16950);
or U24172 (N_24172,N_15094,N_13117);
xnor U24173 (N_24173,N_18673,N_15901);
nand U24174 (N_24174,N_15942,N_17465);
nor U24175 (N_24175,N_15890,N_12582);
or U24176 (N_24176,N_18395,N_18619);
and U24177 (N_24177,N_16841,N_17235);
and U24178 (N_24178,N_18481,N_15763);
and U24179 (N_24179,N_17558,N_18609);
or U24180 (N_24180,N_12908,N_12956);
nor U24181 (N_24181,N_14055,N_13578);
nor U24182 (N_24182,N_17777,N_14886);
nor U24183 (N_24183,N_18706,N_15714);
xor U24184 (N_24184,N_15337,N_12755);
nor U24185 (N_24185,N_16877,N_14963);
nor U24186 (N_24186,N_17614,N_15101);
or U24187 (N_24187,N_17288,N_17495);
nand U24188 (N_24188,N_15413,N_16957);
or U24189 (N_24189,N_13543,N_13934);
nor U24190 (N_24190,N_14035,N_13082);
nand U24191 (N_24191,N_14665,N_13080);
and U24192 (N_24192,N_17178,N_16845);
nand U24193 (N_24193,N_15634,N_15805);
or U24194 (N_24194,N_13788,N_15356);
nor U24195 (N_24195,N_16124,N_18451);
and U24196 (N_24196,N_13276,N_15951);
nand U24197 (N_24197,N_17680,N_18535);
xnor U24198 (N_24198,N_17898,N_16892);
or U24199 (N_24199,N_16982,N_17794);
nand U24200 (N_24200,N_12663,N_14562);
nand U24201 (N_24201,N_14279,N_17552);
nor U24202 (N_24202,N_18261,N_18535);
nand U24203 (N_24203,N_15492,N_13325);
nor U24204 (N_24204,N_14541,N_14878);
or U24205 (N_24205,N_14768,N_14991);
and U24206 (N_24206,N_18143,N_13007);
nor U24207 (N_24207,N_14932,N_18613);
nor U24208 (N_24208,N_18243,N_15392);
xor U24209 (N_24209,N_14726,N_14954);
or U24210 (N_24210,N_16770,N_15836);
or U24211 (N_24211,N_17493,N_16730);
nor U24212 (N_24212,N_14395,N_13632);
or U24213 (N_24213,N_13000,N_14633);
nand U24214 (N_24214,N_14379,N_16831);
and U24215 (N_24215,N_13896,N_15084);
and U24216 (N_24216,N_17269,N_12930);
and U24217 (N_24217,N_13889,N_18620);
and U24218 (N_24218,N_12872,N_17656);
nand U24219 (N_24219,N_15405,N_14933);
nand U24220 (N_24220,N_17983,N_18299);
and U24221 (N_24221,N_16098,N_16429);
or U24222 (N_24222,N_16449,N_14763);
or U24223 (N_24223,N_17653,N_15314);
or U24224 (N_24224,N_13134,N_17808);
or U24225 (N_24225,N_12980,N_12524);
and U24226 (N_24226,N_17084,N_18743);
and U24227 (N_24227,N_13757,N_18190);
and U24228 (N_24228,N_13566,N_15856);
nor U24229 (N_24229,N_14839,N_17342);
nand U24230 (N_24230,N_15680,N_18017);
nand U24231 (N_24231,N_12901,N_14100);
and U24232 (N_24232,N_14669,N_18149);
nor U24233 (N_24233,N_13448,N_16652);
xnor U24234 (N_24234,N_18615,N_18161);
and U24235 (N_24235,N_12894,N_16099);
nand U24236 (N_24236,N_15140,N_17312);
nand U24237 (N_24237,N_18353,N_13518);
nor U24238 (N_24238,N_14997,N_18018);
or U24239 (N_24239,N_18452,N_14742);
nand U24240 (N_24240,N_13119,N_13513);
or U24241 (N_24241,N_14658,N_17204);
nor U24242 (N_24242,N_13681,N_18479);
nor U24243 (N_24243,N_18481,N_15716);
nand U24244 (N_24244,N_17722,N_17064);
nor U24245 (N_24245,N_12601,N_14302);
nand U24246 (N_24246,N_17461,N_12593);
or U24247 (N_24247,N_15882,N_18208);
nand U24248 (N_24248,N_13264,N_14696);
and U24249 (N_24249,N_13987,N_14519);
nand U24250 (N_24250,N_18325,N_18148);
or U24251 (N_24251,N_14447,N_14050);
nand U24252 (N_24252,N_13317,N_14977);
nand U24253 (N_24253,N_14004,N_14472);
xor U24254 (N_24254,N_14483,N_15812);
xor U24255 (N_24255,N_15013,N_15519);
or U24256 (N_24256,N_12938,N_16390);
nand U24257 (N_24257,N_13152,N_12605);
and U24258 (N_24258,N_14240,N_13350);
xnor U24259 (N_24259,N_18729,N_12581);
or U24260 (N_24260,N_15932,N_12517);
or U24261 (N_24261,N_14415,N_13713);
and U24262 (N_24262,N_16148,N_13172);
or U24263 (N_24263,N_14096,N_18563);
nand U24264 (N_24264,N_12636,N_14812);
nor U24265 (N_24265,N_14334,N_15466);
or U24266 (N_24266,N_14928,N_17092);
nand U24267 (N_24267,N_13676,N_14222);
or U24268 (N_24268,N_18703,N_18252);
and U24269 (N_24269,N_16085,N_18540);
xor U24270 (N_24270,N_13362,N_18109);
or U24271 (N_24271,N_15662,N_18424);
and U24272 (N_24272,N_15711,N_17518);
or U24273 (N_24273,N_14900,N_15506);
or U24274 (N_24274,N_12666,N_14789);
xnor U24275 (N_24275,N_17629,N_16608);
and U24276 (N_24276,N_15097,N_13286);
nand U24277 (N_24277,N_16537,N_14419);
nand U24278 (N_24278,N_17412,N_16890);
nor U24279 (N_24279,N_13292,N_12832);
nand U24280 (N_24280,N_14191,N_14695);
and U24281 (N_24281,N_18616,N_12675);
nor U24282 (N_24282,N_12681,N_18591);
and U24283 (N_24283,N_17893,N_18147);
nand U24284 (N_24284,N_18257,N_13774);
and U24285 (N_24285,N_17074,N_18259);
or U24286 (N_24286,N_14228,N_17034);
xnor U24287 (N_24287,N_15471,N_18425);
xor U24288 (N_24288,N_18154,N_17940);
or U24289 (N_24289,N_18105,N_15400);
nand U24290 (N_24290,N_16265,N_16005);
nand U24291 (N_24291,N_15869,N_15405);
nand U24292 (N_24292,N_17984,N_18525);
nand U24293 (N_24293,N_14375,N_13367);
nor U24294 (N_24294,N_18656,N_15160);
or U24295 (N_24295,N_15627,N_16557);
nor U24296 (N_24296,N_14112,N_14425);
or U24297 (N_24297,N_16094,N_16964);
xor U24298 (N_24298,N_18352,N_14585);
and U24299 (N_24299,N_17823,N_17457);
nand U24300 (N_24300,N_12792,N_16177);
or U24301 (N_24301,N_15598,N_17062);
nand U24302 (N_24302,N_12905,N_15772);
and U24303 (N_24303,N_13396,N_15826);
or U24304 (N_24304,N_14526,N_14829);
and U24305 (N_24305,N_15962,N_16215);
nor U24306 (N_24306,N_18177,N_15354);
nor U24307 (N_24307,N_17884,N_14147);
nand U24308 (N_24308,N_15257,N_13653);
or U24309 (N_24309,N_12554,N_18504);
xnor U24310 (N_24310,N_12758,N_17017);
and U24311 (N_24311,N_15978,N_16442);
or U24312 (N_24312,N_15677,N_12733);
nand U24313 (N_24313,N_18479,N_14970);
and U24314 (N_24314,N_17590,N_15157);
xnor U24315 (N_24315,N_17157,N_13400);
nor U24316 (N_24316,N_18574,N_16787);
and U24317 (N_24317,N_15174,N_13855);
nand U24318 (N_24318,N_17499,N_14516);
or U24319 (N_24319,N_18076,N_17136);
nor U24320 (N_24320,N_18084,N_17427);
and U24321 (N_24321,N_14604,N_15119);
nor U24322 (N_24322,N_14298,N_15469);
nor U24323 (N_24323,N_17741,N_14212);
and U24324 (N_24324,N_16804,N_16759);
nand U24325 (N_24325,N_12806,N_13064);
or U24326 (N_24326,N_18520,N_18178);
or U24327 (N_24327,N_15992,N_18525);
nand U24328 (N_24328,N_17835,N_13126);
nand U24329 (N_24329,N_13563,N_16897);
nor U24330 (N_24330,N_15345,N_14425);
nand U24331 (N_24331,N_13450,N_15176);
nor U24332 (N_24332,N_18206,N_13359);
and U24333 (N_24333,N_17992,N_16479);
nand U24334 (N_24334,N_13872,N_12585);
nor U24335 (N_24335,N_13393,N_14403);
nand U24336 (N_24336,N_14320,N_15706);
xor U24337 (N_24337,N_13546,N_16222);
or U24338 (N_24338,N_14474,N_17693);
and U24339 (N_24339,N_16436,N_14251);
nand U24340 (N_24340,N_18026,N_14803);
xnor U24341 (N_24341,N_17927,N_14246);
nor U24342 (N_24342,N_16155,N_15722);
and U24343 (N_24343,N_13342,N_13437);
or U24344 (N_24344,N_15485,N_17375);
nand U24345 (N_24345,N_17390,N_13269);
or U24346 (N_24346,N_16818,N_17731);
nand U24347 (N_24347,N_12630,N_12507);
nand U24348 (N_24348,N_13331,N_14345);
or U24349 (N_24349,N_15036,N_15383);
nand U24350 (N_24350,N_14229,N_14275);
and U24351 (N_24351,N_15077,N_14239);
and U24352 (N_24352,N_18286,N_18357);
and U24353 (N_24353,N_16537,N_16774);
and U24354 (N_24354,N_16668,N_14378);
nor U24355 (N_24355,N_15552,N_15856);
nor U24356 (N_24356,N_12554,N_14281);
or U24357 (N_24357,N_13414,N_13983);
and U24358 (N_24358,N_15677,N_16255);
or U24359 (N_24359,N_13529,N_16102);
or U24360 (N_24360,N_12935,N_16818);
or U24361 (N_24361,N_16291,N_13962);
and U24362 (N_24362,N_17763,N_15274);
nor U24363 (N_24363,N_16997,N_16143);
and U24364 (N_24364,N_17312,N_16885);
xor U24365 (N_24365,N_14817,N_15301);
xor U24366 (N_24366,N_15683,N_15356);
and U24367 (N_24367,N_15038,N_17736);
or U24368 (N_24368,N_12765,N_17439);
or U24369 (N_24369,N_17505,N_12677);
or U24370 (N_24370,N_14199,N_16247);
and U24371 (N_24371,N_13283,N_14659);
nor U24372 (N_24372,N_15753,N_16904);
or U24373 (N_24373,N_13805,N_15564);
nor U24374 (N_24374,N_17122,N_16941);
xnor U24375 (N_24375,N_15699,N_18735);
nor U24376 (N_24376,N_13970,N_15850);
nor U24377 (N_24377,N_17280,N_16304);
or U24378 (N_24378,N_17774,N_14291);
and U24379 (N_24379,N_12608,N_15111);
nor U24380 (N_24380,N_13930,N_16230);
nor U24381 (N_24381,N_14938,N_12608);
nand U24382 (N_24382,N_16399,N_15014);
or U24383 (N_24383,N_16509,N_13113);
nand U24384 (N_24384,N_18139,N_17524);
or U24385 (N_24385,N_18255,N_15198);
xnor U24386 (N_24386,N_18100,N_12913);
nand U24387 (N_24387,N_16054,N_13855);
nor U24388 (N_24388,N_14158,N_15243);
and U24389 (N_24389,N_16996,N_16411);
nand U24390 (N_24390,N_14359,N_13773);
nor U24391 (N_24391,N_12841,N_15898);
and U24392 (N_24392,N_17126,N_17595);
nand U24393 (N_24393,N_16625,N_14194);
nor U24394 (N_24394,N_15070,N_14827);
nor U24395 (N_24395,N_17854,N_17597);
and U24396 (N_24396,N_17414,N_17405);
and U24397 (N_24397,N_17018,N_12826);
nand U24398 (N_24398,N_13357,N_14250);
or U24399 (N_24399,N_18394,N_14428);
nor U24400 (N_24400,N_16795,N_13416);
or U24401 (N_24401,N_17996,N_16622);
xnor U24402 (N_24402,N_18400,N_17285);
xnor U24403 (N_24403,N_18668,N_13686);
or U24404 (N_24404,N_16982,N_12563);
xor U24405 (N_24405,N_14203,N_17556);
nor U24406 (N_24406,N_14073,N_15383);
or U24407 (N_24407,N_15049,N_13461);
nor U24408 (N_24408,N_12552,N_16378);
or U24409 (N_24409,N_13461,N_16965);
xor U24410 (N_24410,N_12864,N_18198);
xnor U24411 (N_24411,N_14972,N_16919);
and U24412 (N_24412,N_18359,N_18114);
xnor U24413 (N_24413,N_17895,N_13291);
xnor U24414 (N_24414,N_13603,N_17089);
nor U24415 (N_24415,N_17332,N_15421);
and U24416 (N_24416,N_13391,N_14702);
and U24417 (N_24417,N_12640,N_17918);
xnor U24418 (N_24418,N_15733,N_14706);
and U24419 (N_24419,N_18507,N_18296);
nand U24420 (N_24420,N_18406,N_12596);
and U24421 (N_24421,N_13117,N_15594);
and U24422 (N_24422,N_16952,N_15220);
nand U24423 (N_24423,N_13971,N_16133);
nor U24424 (N_24424,N_15324,N_14891);
and U24425 (N_24425,N_14660,N_14042);
or U24426 (N_24426,N_14373,N_16613);
and U24427 (N_24427,N_12819,N_15193);
xnor U24428 (N_24428,N_18322,N_17979);
or U24429 (N_24429,N_14140,N_15605);
nand U24430 (N_24430,N_13580,N_17468);
nor U24431 (N_24431,N_15467,N_17397);
nand U24432 (N_24432,N_13128,N_18647);
or U24433 (N_24433,N_13337,N_13222);
or U24434 (N_24434,N_17360,N_15687);
or U24435 (N_24435,N_16303,N_17347);
nor U24436 (N_24436,N_13912,N_16730);
xnor U24437 (N_24437,N_13970,N_14738);
nand U24438 (N_24438,N_16256,N_16372);
nor U24439 (N_24439,N_15584,N_18132);
nand U24440 (N_24440,N_16576,N_14507);
nor U24441 (N_24441,N_13819,N_12720);
and U24442 (N_24442,N_16639,N_15704);
xnor U24443 (N_24443,N_14156,N_17469);
nand U24444 (N_24444,N_15918,N_18651);
nand U24445 (N_24445,N_12505,N_16826);
nor U24446 (N_24446,N_15179,N_16616);
or U24447 (N_24447,N_18057,N_15070);
or U24448 (N_24448,N_14341,N_15257);
nor U24449 (N_24449,N_15560,N_15408);
nor U24450 (N_24450,N_16083,N_15914);
nor U24451 (N_24451,N_13404,N_14820);
nor U24452 (N_24452,N_18285,N_16795);
nand U24453 (N_24453,N_14055,N_14172);
or U24454 (N_24454,N_16867,N_16196);
and U24455 (N_24455,N_15088,N_18288);
or U24456 (N_24456,N_12609,N_14746);
nand U24457 (N_24457,N_16821,N_15560);
or U24458 (N_24458,N_14927,N_16150);
nor U24459 (N_24459,N_14825,N_14197);
or U24460 (N_24460,N_16168,N_13427);
and U24461 (N_24461,N_14775,N_13487);
nand U24462 (N_24462,N_14881,N_17862);
nand U24463 (N_24463,N_13516,N_14853);
or U24464 (N_24464,N_12507,N_12572);
nand U24465 (N_24465,N_14458,N_15216);
or U24466 (N_24466,N_16777,N_16700);
nor U24467 (N_24467,N_18379,N_16442);
or U24468 (N_24468,N_18276,N_13498);
nand U24469 (N_24469,N_17487,N_17389);
xor U24470 (N_24470,N_14623,N_17409);
or U24471 (N_24471,N_15327,N_13955);
or U24472 (N_24472,N_14127,N_13701);
and U24473 (N_24473,N_16168,N_17808);
or U24474 (N_24474,N_18681,N_14073);
nand U24475 (N_24475,N_15769,N_17144);
nand U24476 (N_24476,N_17714,N_18206);
or U24477 (N_24477,N_16186,N_17495);
nor U24478 (N_24478,N_15748,N_17795);
and U24479 (N_24479,N_14326,N_15026);
nand U24480 (N_24480,N_18672,N_15795);
or U24481 (N_24481,N_18355,N_15475);
and U24482 (N_24482,N_12972,N_16736);
nand U24483 (N_24483,N_17121,N_17524);
and U24484 (N_24484,N_14683,N_17103);
and U24485 (N_24485,N_12836,N_17582);
and U24486 (N_24486,N_18703,N_13980);
and U24487 (N_24487,N_14679,N_15870);
nor U24488 (N_24488,N_13415,N_12753);
or U24489 (N_24489,N_12623,N_18046);
nor U24490 (N_24490,N_18251,N_16482);
nand U24491 (N_24491,N_15582,N_15045);
and U24492 (N_24492,N_18533,N_17470);
and U24493 (N_24493,N_16960,N_14117);
and U24494 (N_24494,N_18683,N_17150);
nand U24495 (N_24495,N_16120,N_15014);
or U24496 (N_24496,N_13319,N_17349);
xnor U24497 (N_24497,N_12718,N_13145);
nand U24498 (N_24498,N_14935,N_15477);
and U24499 (N_24499,N_14458,N_16490);
and U24500 (N_24500,N_16639,N_15486);
xnor U24501 (N_24501,N_17892,N_12760);
nand U24502 (N_24502,N_17158,N_17750);
nand U24503 (N_24503,N_17723,N_16610);
and U24504 (N_24504,N_14867,N_18484);
nand U24505 (N_24505,N_18725,N_16312);
and U24506 (N_24506,N_13091,N_18267);
nor U24507 (N_24507,N_13142,N_18683);
or U24508 (N_24508,N_13727,N_16732);
and U24509 (N_24509,N_14716,N_17215);
nor U24510 (N_24510,N_17391,N_16582);
nand U24511 (N_24511,N_17510,N_14921);
or U24512 (N_24512,N_16098,N_17967);
nand U24513 (N_24513,N_13445,N_13288);
and U24514 (N_24514,N_13096,N_12699);
and U24515 (N_24515,N_17672,N_14050);
nor U24516 (N_24516,N_17769,N_13836);
nor U24517 (N_24517,N_14055,N_16732);
or U24518 (N_24518,N_13060,N_18607);
or U24519 (N_24519,N_16783,N_14014);
or U24520 (N_24520,N_13091,N_13190);
xnor U24521 (N_24521,N_14751,N_14268);
and U24522 (N_24522,N_14069,N_18306);
nand U24523 (N_24523,N_14498,N_13285);
or U24524 (N_24524,N_18745,N_18569);
and U24525 (N_24525,N_12906,N_14283);
or U24526 (N_24526,N_13078,N_16301);
nor U24527 (N_24527,N_14036,N_13824);
or U24528 (N_24528,N_14654,N_12651);
and U24529 (N_24529,N_15321,N_15009);
nand U24530 (N_24530,N_15147,N_14199);
or U24531 (N_24531,N_14144,N_14821);
nand U24532 (N_24532,N_15831,N_14008);
nand U24533 (N_24533,N_14601,N_16015);
and U24534 (N_24534,N_15274,N_15131);
and U24535 (N_24535,N_12886,N_15954);
or U24536 (N_24536,N_17313,N_16268);
and U24537 (N_24537,N_15910,N_13990);
or U24538 (N_24538,N_18740,N_18102);
and U24539 (N_24539,N_14404,N_18133);
nand U24540 (N_24540,N_17464,N_17546);
nand U24541 (N_24541,N_17744,N_15384);
or U24542 (N_24542,N_18409,N_15385);
nor U24543 (N_24543,N_17521,N_15585);
nor U24544 (N_24544,N_16836,N_13530);
nor U24545 (N_24545,N_13566,N_17948);
nor U24546 (N_24546,N_15507,N_12856);
and U24547 (N_24547,N_18400,N_12654);
or U24548 (N_24548,N_12799,N_12758);
nor U24549 (N_24549,N_16756,N_14085);
nand U24550 (N_24550,N_17183,N_15437);
or U24551 (N_24551,N_16418,N_14171);
and U24552 (N_24552,N_13431,N_13970);
nand U24553 (N_24553,N_16557,N_15370);
nor U24554 (N_24554,N_12674,N_16140);
or U24555 (N_24555,N_17647,N_15543);
nor U24556 (N_24556,N_15994,N_15807);
or U24557 (N_24557,N_18225,N_14623);
nand U24558 (N_24558,N_16583,N_16542);
nand U24559 (N_24559,N_12543,N_15918);
and U24560 (N_24560,N_15936,N_15552);
or U24561 (N_24561,N_17247,N_17961);
and U24562 (N_24562,N_18112,N_13887);
nand U24563 (N_24563,N_16664,N_17238);
nor U24564 (N_24564,N_17573,N_17947);
nand U24565 (N_24565,N_12532,N_13401);
nand U24566 (N_24566,N_16588,N_18607);
nor U24567 (N_24567,N_17071,N_16633);
nand U24568 (N_24568,N_16157,N_16598);
or U24569 (N_24569,N_13786,N_17478);
or U24570 (N_24570,N_13849,N_12666);
nand U24571 (N_24571,N_14454,N_17385);
or U24572 (N_24572,N_17928,N_15954);
and U24573 (N_24573,N_13093,N_13374);
nand U24574 (N_24574,N_15401,N_15367);
or U24575 (N_24575,N_16772,N_15837);
nor U24576 (N_24576,N_16601,N_16603);
or U24577 (N_24577,N_18147,N_13602);
and U24578 (N_24578,N_13539,N_14299);
xnor U24579 (N_24579,N_18341,N_13024);
or U24580 (N_24580,N_13252,N_12645);
nand U24581 (N_24581,N_15286,N_14798);
nor U24582 (N_24582,N_14911,N_15284);
nor U24583 (N_24583,N_17350,N_12514);
or U24584 (N_24584,N_17918,N_17832);
nor U24585 (N_24585,N_14459,N_13961);
and U24586 (N_24586,N_14691,N_15670);
nand U24587 (N_24587,N_13473,N_13981);
or U24588 (N_24588,N_18581,N_18747);
and U24589 (N_24589,N_18508,N_17289);
or U24590 (N_24590,N_17345,N_12696);
or U24591 (N_24591,N_14157,N_16168);
or U24592 (N_24592,N_15789,N_17434);
and U24593 (N_24593,N_17225,N_14518);
nor U24594 (N_24594,N_15079,N_13213);
and U24595 (N_24595,N_17951,N_13264);
xor U24596 (N_24596,N_13635,N_15508);
or U24597 (N_24597,N_12873,N_17310);
xnor U24598 (N_24598,N_14601,N_16416);
or U24599 (N_24599,N_18022,N_15088);
nor U24600 (N_24600,N_15620,N_15844);
and U24601 (N_24601,N_17109,N_12679);
xnor U24602 (N_24602,N_16005,N_14413);
nor U24603 (N_24603,N_14163,N_18508);
nor U24604 (N_24604,N_16526,N_16179);
nand U24605 (N_24605,N_14615,N_16225);
or U24606 (N_24606,N_17556,N_15334);
or U24607 (N_24607,N_18037,N_14670);
nand U24608 (N_24608,N_17562,N_14132);
xor U24609 (N_24609,N_18318,N_12893);
nor U24610 (N_24610,N_13646,N_17630);
or U24611 (N_24611,N_16100,N_13923);
nand U24612 (N_24612,N_13849,N_12719);
nor U24613 (N_24613,N_15837,N_13472);
or U24614 (N_24614,N_12583,N_14209);
or U24615 (N_24615,N_17336,N_16192);
or U24616 (N_24616,N_15089,N_14977);
or U24617 (N_24617,N_16341,N_15080);
nor U24618 (N_24618,N_14661,N_14226);
nor U24619 (N_24619,N_12767,N_16099);
nor U24620 (N_24620,N_17980,N_13260);
nor U24621 (N_24621,N_18318,N_15141);
and U24622 (N_24622,N_18062,N_17063);
or U24623 (N_24623,N_17160,N_18072);
nand U24624 (N_24624,N_15616,N_14586);
nor U24625 (N_24625,N_13829,N_17703);
or U24626 (N_24626,N_13779,N_14370);
nor U24627 (N_24627,N_18219,N_13249);
xnor U24628 (N_24628,N_15421,N_18300);
or U24629 (N_24629,N_14831,N_18287);
and U24630 (N_24630,N_15226,N_13950);
or U24631 (N_24631,N_13714,N_17540);
and U24632 (N_24632,N_18453,N_17748);
nand U24633 (N_24633,N_13189,N_16938);
or U24634 (N_24634,N_12644,N_16929);
nor U24635 (N_24635,N_16597,N_13175);
nor U24636 (N_24636,N_15042,N_16881);
xnor U24637 (N_24637,N_13805,N_18409);
or U24638 (N_24638,N_13238,N_17374);
and U24639 (N_24639,N_18444,N_15863);
and U24640 (N_24640,N_15238,N_18134);
and U24641 (N_24641,N_18659,N_14780);
nor U24642 (N_24642,N_15118,N_16640);
or U24643 (N_24643,N_15075,N_17320);
nand U24644 (N_24644,N_16115,N_13734);
and U24645 (N_24645,N_15025,N_12796);
nand U24646 (N_24646,N_14390,N_12631);
xnor U24647 (N_24647,N_16162,N_12634);
or U24648 (N_24648,N_14740,N_13433);
nor U24649 (N_24649,N_14887,N_18479);
or U24650 (N_24650,N_14128,N_15794);
or U24651 (N_24651,N_13830,N_15595);
nand U24652 (N_24652,N_15522,N_15554);
nand U24653 (N_24653,N_13079,N_17585);
nor U24654 (N_24654,N_13588,N_16801);
or U24655 (N_24655,N_18095,N_17532);
and U24656 (N_24656,N_14907,N_15139);
nor U24657 (N_24657,N_17557,N_12679);
and U24658 (N_24658,N_16889,N_17481);
xnor U24659 (N_24659,N_14162,N_18368);
and U24660 (N_24660,N_15775,N_12698);
nor U24661 (N_24661,N_17014,N_16863);
or U24662 (N_24662,N_14354,N_13132);
nor U24663 (N_24663,N_18142,N_17408);
nand U24664 (N_24664,N_17793,N_18162);
nor U24665 (N_24665,N_18661,N_14940);
and U24666 (N_24666,N_14475,N_15508);
and U24667 (N_24667,N_13406,N_13675);
nand U24668 (N_24668,N_14001,N_12931);
or U24669 (N_24669,N_15947,N_13489);
and U24670 (N_24670,N_18232,N_13964);
nor U24671 (N_24671,N_14083,N_14726);
xnor U24672 (N_24672,N_14237,N_17802);
nor U24673 (N_24673,N_13093,N_16288);
nor U24674 (N_24674,N_12626,N_17098);
and U24675 (N_24675,N_17225,N_15624);
and U24676 (N_24676,N_18521,N_15368);
nor U24677 (N_24677,N_16519,N_16725);
and U24678 (N_24678,N_12747,N_16212);
or U24679 (N_24679,N_18573,N_16276);
xor U24680 (N_24680,N_17461,N_13809);
or U24681 (N_24681,N_18341,N_14570);
nor U24682 (N_24682,N_15876,N_14152);
nand U24683 (N_24683,N_12792,N_13142);
nand U24684 (N_24684,N_15600,N_18635);
and U24685 (N_24685,N_17249,N_16066);
nand U24686 (N_24686,N_17262,N_17790);
xor U24687 (N_24687,N_12832,N_12966);
or U24688 (N_24688,N_13379,N_14531);
nand U24689 (N_24689,N_13266,N_14641);
or U24690 (N_24690,N_17661,N_14489);
and U24691 (N_24691,N_12976,N_18034);
nand U24692 (N_24692,N_16536,N_15036);
and U24693 (N_24693,N_15966,N_13581);
nor U24694 (N_24694,N_14257,N_12582);
nor U24695 (N_24695,N_17973,N_17644);
xor U24696 (N_24696,N_15841,N_18674);
and U24697 (N_24697,N_13078,N_17846);
and U24698 (N_24698,N_13140,N_16810);
nor U24699 (N_24699,N_17613,N_18591);
nor U24700 (N_24700,N_18173,N_18057);
nor U24701 (N_24701,N_13779,N_18697);
and U24702 (N_24702,N_14540,N_14960);
nand U24703 (N_24703,N_16721,N_16485);
nand U24704 (N_24704,N_18549,N_18427);
nand U24705 (N_24705,N_12927,N_13652);
and U24706 (N_24706,N_13997,N_13283);
nand U24707 (N_24707,N_16184,N_14674);
or U24708 (N_24708,N_14069,N_17517);
and U24709 (N_24709,N_16492,N_17858);
and U24710 (N_24710,N_15643,N_15431);
xor U24711 (N_24711,N_15356,N_15471);
xor U24712 (N_24712,N_14584,N_14939);
or U24713 (N_24713,N_16755,N_17465);
nor U24714 (N_24714,N_16692,N_16276);
or U24715 (N_24715,N_16426,N_16431);
and U24716 (N_24716,N_13874,N_16044);
xnor U24717 (N_24717,N_12510,N_17607);
nand U24718 (N_24718,N_18118,N_15675);
nor U24719 (N_24719,N_16810,N_15450);
or U24720 (N_24720,N_14050,N_16834);
nand U24721 (N_24721,N_14458,N_13263);
nand U24722 (N_24722,N_13517,N_13129);
nor U24723 (N_24723,N_13768,N_14159);
nand U24724 (N_24724,N_13288,N_17438);
and U24725 (N_24725,N_13996,N_17388);
or U24726 (N_24726,N_13684,N_16886);
and U24727 (N_24727,N_14540,N_17172);
or U24728 (N_24728,N_16027,N_14962);
nor U24729 (N_24729,N_14311,N_17312);
and U24730 (N_24730,N_18164,N_15024);
nor U24731 (N_24731,N_18186,N_14498);
nor U24732 (N_24732,N_13277,N_15019);
or U24733 (N_24733,N_15620,N_12839);
or U24734 (N_24734,N_17990,N_13558);
xnor U24735 (N_24735,N_15184,N_15340);
nor U24736 (N_24736,N_16899,N_15121);
nor U24737 (N_24737,N_13712,N_18659);
and U24738 (N_24738,N_16742,N_16757);
and U24739 (N_24739,N_14190,N_12606);
nor U24740 (N_24740,N_15764,N_14335);
xor U24741 (N_24741,N_15578,N_12914);
nand U24742 (N_24742,N_15709,N_12766);
or U24743 (N_24743,N_17546,N_18101);
nor U24744 (N_24744,N_14312,N_13383);
and U24745 (N_24745,N_16866,N_17252);
or U24746 (N_24746,N_16853,N_18483);
and U24747 (N_24747,N_14120,N_13506);
nor U24748 (N_24748,N_16467,N_12933);
nor U24749 (N_24749,N_16500,N_15600);
xnor U24750 (N_24750,N_17440,N_12531);
nand U24751 (N_24751,N_13682,N_14397);
and U24752 (N_24752,N_13186,N_14801);
and U24753 (N_24753,N_14871,N_15042);
and U24754 (N_24754,N_15552,N_15127);
or U24755 (N_24755,N_18243,N_17533);
or U24756 (N_24756,N_15932,N_15492);
and U24757 (N_24757,N_15458,N_18580);
nor U24758 (N_24758,N_13019,N_12969);
and U24759 (N_24759,N_18566,N_18354);
nand U24760 (N_24760,N_13806,N_18680);
xor U24761 (N_24761,N_14825,N_18489);
and U24762 (N_24762,N_18325,N_12983);
nor U24763 (N_24763,N_13999,N_17702);
nor U24764 (N_24764,N_18391,N_15831);
and U24765 (N_24765,N_13332,N_15674);
nand U24766 (N_24766,N_17308,N_17985);
nand U24767 (N_24767,N_15645,N_12571);
xnor U24768 (N_24768,N_18678,N_17125);
nor U24769 (N_24769,N_18748,N_14390);
or U24770 (N_24770,N_16503,N_15141);
xnor U24771 (N_24771,N_15015,N_13411);
nand U24772 (N_24772,N_14418,N_14042);
nand U24773 (N_24773,N_18455,N_14851);
nor U24774 (N_24774,N_17593,N_12608);
and U24775 (N_24775,N_16657,N_13658);
and U24776 (N_24776,N_17571,N_14350);
and U24777 (N_24777,N_18145,N_17608);
or U24778 (N_24778,N_14448,N_16905);
nor U24779 (N_24779,N_18450,N_17077);
nor U24780 (N_24780,N_14511,N_13096);
or U24781 (N_24781,N_17972,N_17433);
nand U24782 (N_24782,N_12628,N_13777);
or U24783 (N_24783,N_17475,N_13081);
nand U24784 (N_24784,N_12727,N_15490);
or U24785 (N_24785,N_16258,N_15056);
nor U24786 (N_24786,N_18043,N_14155);
nor U24787 (N_24787,N_14153,N_14348);
xnor U24788 (N_24788,N_13794,N_14750);
nand U24789 (N_24789,N_12814,N_16378);
nand U24790 (N_24790,N_16128,N_12584);
nand U24791 (N_24791,N_18591,N_14510);
or U24792 (N_24792,N_16034,N_17019);
xnor U24793 (N_24793,N_16574,N_16576);
or U24794 (N_24794,N_17597,N_15542);
nor U24795 (N_24795,N_15218,N_16799);
nor U24796 (N_24796,N_15790,N_12970);
xor U24797 (N_24797,N_12701,N_15081);
nand U24798 (N_24798,N_14620,N_16967);
nor U24799 (N_24799,N_14473,N_18022);
nor U24800 (N_24800,N_16549,N_14296);
nor U24801 (N_24801,N_14657,N_14661);
and U24802 (N_24802,N_15708,N_13607);
nor U24803 (N_24803,N_17678,N_18373);
xnor U24804 (N_24804,N_14599,N_14382);
nand U24805 (N_24805,N_15654,N_12893);
and U24806 (N_24806,N_17451,N_18053);
and U24807 (N_24807,N_14828,N_15854);
xnor U24808 (N_24808,N_17465,N_16956);
xnor U24809 (N_24809,N_17498,N_13789);
or U24810 (N_24810,N_13862,N_15329);
nand U24811 (N_24811,N_16798,N_17678);
or U24812 (N_24812,N_12927,N_16971);
nor U24813 (N_24813,N_17210,N_14882);
or U24814 (N_24814,N_17367,N_15571);
xnor U24815 (N_24815,N_15392,N_13630);
nand U24816 (N_24816,N_14268,N_16112);
and U24817 (N_24817,N_16458,N_15157);
nor U24818 (N_24818,N_17869,N_15543);
nand U24819 (N_24819,N_17905,N_13488);
nand U24820 (N_24820,N_14897,N_16978);
nor U24821 (N_24821,N_18228,N_15990);
and U24822 (N_24822,N_16258,N_17082);
nand U24823 (N_24823,N_14061,N_12542);
nand U24824 (N_24824,N_15180,N_16678);
xnor U24825 (N_24825,N_17994,N_18249);
or U24826 (N_24826,N_13256,N_17260);
and U24827 (N_24827,N_18027,N_14322);
or U24828 (N_24828,N_16883,N_17447);
nor U24829 (N_24829,N_14645,N_12897);
nor U24830 (N_24830,N_16935,N_14448);
nor U24831 (N_24831,N_15971,N_16714);
nand U24832 (N_24832,N_18216,N_17086);
nand U24833 (N_24833,N_17071,N_14099);
nor U24834 (N_24834,N_15762,N_14000);
or U24835 (N_24835,N_17550,N_14884);
nor U24836 (N_24836,N_18147,N_14860);
xor U24837 (N_24837,N_16970,N_14974);
nor U24838 (N_24838,N_16738,N_13061);
and U24839 (N_24839,N_16519,N_16799);
xnor U24840 (N_24840,N_14770,N_15097);
xnor U24841 (N_24841,N_14455,N_16567);
and U24842 (N_24842,N_16452,N_16982);
nor U24843 (N_24843,N_13931,N_16115);
nand U24844 (N_24844,N_14627,N_15302);
nor U24845 (N_24845,N_15560,N_15059);
nand U24846 (N_24846,N_13597,N_18240);
nor U24847 (N_24847,N_15264,N_14669);
nand U24848 (N_24848,N_12720,N_16421);
nand U24849 (N_24849,N_12925,N_16615);
nor U24850 (N_24850,N_15526,N_17851);
nor U24851 (N_24851,N_12908,N_18348);
xor U24852 (N_24852,N_18229,N_18049);
nor U24853 (N_24853,N_15584,N_18714);
nand U24854 (N_24854,N_13397,N_15681);
and U24855 (N_24855,N_18515,N_13924);
and U24856 (N_24856,N_16570,N_14101);
xnor U24857 (N_24857,N_15233,N_13595);
or U24858 (N_24858,N_13898,N_14602);
or U24859 (N_24859,N_17222,N_16669);
or U24860 (N_24860,N_15094,N_15847);
and U24861 (N_24861,N_17121,N_16138);
and U24862 (N_24862,N_18044,N_13576);
nor U24863 (N_24863,N_15922,N_15473);
and U24864 (N_24864,N_15452,N_18032);
or U24865 (N_24865,N_13398,N_12700);
or U24866 (N_24866,N_15883,N_18312);
or U24867 (N_24867,N_13270,N_12690);
and U24868 (N_24868,N_13913,N_18199);
nor U24869 (N_24869,N_18190,N_14416);
and U24870 (N_24870,N_13846,N_14435);
and U24871 (N_24871,N_17192,N_15825);
and U24872 (N_24872,N_15482,N_16132);
xnor U24873 (N_24873,N_16728,N_12952);
and U24874 (N_24874,N_13435,N_15801);
nand U24875 (N_24875,N_16354,N_13315);
and U24876 (N_24876,N_12621,N_15093);
nand U24877 (N_24877,N_18318,N_18463);
or U24878 (N_24878,N_12753,N_16835);
or U24879 (N_24879,N_13674,N_14477);
nand U24880 (N_24880,N_16636,N_12638);
nor U24881 (N_24881,N_17794,N_13281);
nand U24882 (N_24882,N_15289,N_18237);
nand U24883 (N_24883,N_17623,N_15915);
and U24884 (N_24884,N_18677,N_17426);
nor U24885 (N_24885,N_14339,N_15091);
or U24886 (N_24886,N_14998,N_13506);
or U24887 (N_24887,N_18431,N_15546);
xnor U24888 (N_24888,N_14596,N_13521);
nor U24889 (N_24889,N_17591,N_15064);
nand U24890 (N_24890,N_13279,N_15631);
or U24891 (N_24891,N_12901,N_15433);
nand U24892 (N_24892,N_16260,N_15027);
or U24893 (N_24893,N_16297,N_16793);
nand U24894 (N_24894,N_14174,N_15514);
xnor U24895 (N_24895,N_18201,N_17097);
nand U24896 (N_24896,N_16825,N_12596);
nand U24897 (N_24897,N_14928,N_18102);
and U24898 (N_24898,N_15036,N_16170);
and U24899 (N_24899,N_12695,N_16486);
nor U24900 (N_24900,N_17863,N_18570);
or U24901 (N_24901,N_15217,N_18279);
nor U24902 (N_24902,N_14747,N_14323);
nor U24903 (N_24903,N_13438,N_17267);
or U24904 (N_24904,N_18253,N_14583);
xnor U24905 (N_24905,N_13702,N_15932);
nor U24906 (N_24906,N_17173,N_15709);
and U24907 (N_24907,N_17349,N_14772);
and U24908 (N_24908,N_16094,N_13745);
and U24909 (N_24909,N_16583,N_17834);
and U24910 (N_24910,N_12720,N_17684);
or U24911 (N_24911,N_16506,N_14490);
or U24912 (N_24912,N_13812,N_17524);
nand U24913 (N_24913,N_14553,N_13971);
or U24914 (N_24914,N_14501,N_14626);
nor U24915 (N_24915,N_18354,N_14369);
xnor U24916 (N_24916,N_17193,N_16145);
xor U24917 (N_24917,N_16150,N_17114);
and U24918 (N_24918,N_14728,N_14174);
or U24919 (N_24919,N_15463,N_15365);
nor U24920 (N_24920,N_16595,N_13050);
nand U24921 (N_24921,N_18222,N_18026);
and U24922 (N_24922,N_13354,N_18483);
and U24923 (N_24923,N_16568,N_15096);
and U24924 (N_24924,N_12708,N_13069);
and U24925 (N_24925,N_15352,N_16996);
and U24926 (N_24926,N_16086,N_17056);
nor U24927 (N_24927,N_14781,N_16725);
or U24928 (N_24928,N_13428,N_16179);
nor U24929 (N_24929,N_17174,N_16806);
nor U24930 (N_24930,N_15082,N_17323);
xnor U24931 (N_24931,N_15187,N_15977);
nand U24932 (N_24932,N_17309,N_14445);
or U24933 (N_24933,N_13144,N_17368);
nand U24934 (N_24934,N_14041,N_15299);
nor U24935 (N_24935,N_17373,N_17929);
nand U24936 (N_24936,N_14887,N_12557);
nand U24937 (N_24937,N_16059,N_15892);
nand U24938 (N_24938,N_12815,N_16454);
or U24939 (N_24939,N_17886,N_12603);
or U24940 (N_24940,N_18235,N_13660);
nand U24941 (N_24941,N_18085,N_17694);
and U24942 (N_24942,N_13910,N_13934);
or U24943 (N_24943,N_13592,N_16388);
and U24944 (N_24944,N_16878,N_14068);
nand U24945 (N_24945,N_18563,N_12649);
nand U24946 (N_24946,N_17111,N_15490);
and U24947 (N_24947,N_15706,N_18709);
or U24948 (N_24948,N_17944,N_16958);
or U24949 (N_24949,N_13853,N_16160);
nand U24950 (N_24950,N_18610,N_17222);
nor U24951 (N_24951,N_15378,N_16503);
nand U24952 (N_24952,N_13574,N_18354);
nor U24953 (N_24953,N_15150,N_18059);
xnor U24954 (N_24954,N_16973,N_17515);
or U24955 (N_24955,N_17294,N_13476);
and U24956 (N_24956,N_14777,N_18635);
or U24957 (N_24957,N_17014,N_14360);
or U24958 (N_24958,N_15791,N_15778);
and U24959 (N_24959,N_13756,N_13605);
or U24960 (N_24960,N_15518,N_13348);
or U24961 (N_24961,N_17997,N_13776);
and U24962 (N_24962,N_14052,N_16645);
and U24963 (N_24963,N_15844,N_12982);
and U24964 (N_24964,N_15511,N_15789);
nand U24965 (N_24965,N_12613,N_14032);
and U24966 (N_24966,N_14615,N_16115);
or U24967 (N_24967,N_12674,N_14158);
or U24968 (N_24968,N_13060,N_18735);
or U24969 (N_24969,N_15966,N_18598);
xor U24970 (N_24970,N_16129,N_12826);
nor U24971 (N_24971,N_13209,N_16656);
nand U24972 (N_24972,N_16683,N_15077);
xor U24973 (N_24973,N_15379,N_18260);
nand U24974 (N_24974,N_14703,N_13433);
nor U24975 (N_24975,N_16905,N_13164);
or U24976 (N_24976,N_16370,N_17029);
nor U24977 (N_24977,N_13119,N_17645);
and U24978 (N_24978,N_18380,N_17652);
and U24979 (N_24979,N_17873,N_14176);
and U24980 (N_24980,N_15051,N_16398);
and U24981 (N_24981,N_15202,N_14236);
and U24982 (N_24982,N_16015,N_17991);
xor U24983 (N_24983,N_17161,N_18599);
and U24984 (N_24984,N_16815,N_13846);
nand U24985 (N_24985,N_14746,N_16838);
nor U24986 (N_24986,N_16212,N_16847);
nor U24987 (N_24987,N_17877,N_15831);
nor U24988 (N_24988,N_14293,N_12943);
nor U24989 (N_24989,N_13036,N_13887);
nor U24990 (N_24990,N_18115,N_15924);
nor U24991 (N_24991,N_18315,N_13853);
nor U24992 (N_24992,N_13552,N_15184);
and U24993 (N_24993,N_16171,N_14966);
and U24994 (N_24994,N_16888,N_13074);
and U24995 (N_24995,N_18565,N_15530);
nor U24996 (N_24996,N_16259,N_14507);
and U24997 (N_24997,N_15082,N_12529);
xor U24998 (N_24998,N_15195,N_17993);
nand U24999 (N_24999,N_18077,N_16953);
nor UO_0 (O_0,N_23187,N_22986);
nand UO_1 (O_1,N_22103,N_24694);
and UO_2 (O_2,N_24141,N_21239);
or UO_3 (O_3,N_19703,N_19585);
or UO_4 (O_4,N_23559,N_22887);
nor UO_5 (O_5,N_20151,N_18918);
or UO_6 (O_6,N_19044,N_20840);
and UO_7 (O_7,N_20883,N_22140);
nand UO_8 (O_8,N_20963,N_22019);
nor UO_9 (O_9,N_22203,N_21774);
and UO_10 (O_10,N_23826,N_24058);
or UO_11 (O_11,N_24602,N_21358);
nor UO_12 (O_12,N_21155,N_23135);
nand UO_13 (O_13,N_22966,N_22039);
or UO_14 (O_14,N_22586,N_22016);
nand UO_15 (O_15,N_19224,N_23496);
nor UO_16 (O_16,N_19090,N_23262);
xor UO_17 (O_17,N_20948,N_24879);
and UO_18 (O_18,N_23665,N_22158);
or UO_19 (O_19,N_23145,N_23983);
or UO_20 (O_20,N_21786,N_20373);
nand UO_21 (O_21,N_20177,N_23193);
and UO_22 (O_22,N_20809,N_24130);
or UO_23 (O_23,N_24746,N_24846);
and UO_24 (O_24,N_20403,N_19430);
nand UO_25 (O_25,N_23204,N_21975);
or UO_26 (O_26,N_19136,N_23605);
nor UO_27 (O_27,N_21261,N_24573);
nor UO_28 (O_28,N_23719,N_21646);
or UO_29 (O_29,N_18939,N_24240);
or UO_30 (O_30,N_20350,N_22177);
or UO_31 (O_31,N_24350,N_20123);
xnor UO_32 (O_32,N_22637,N_20641);
nand UO_33 (O_33,N_20141,N_20608);
nand UO_34 (O_34,N_22421,N_23754);
xnor UO_35 (O_35,N_22962,N_21010);
or UO_36 (O_36,N_22467,N_20895);
and UO_37 (O_37,N_18812,N_22600);
nor UO_38 (O_38,N_21596,N_22684);
nand UO_39 (O_39,N_21340,N_19126);
and UO_40 (O_40,N_22068,N_20481);
or UO_41 (O_41,N_21073,N_24120);
or UO_42 (O_42,N_20708,N_20602);
nor UO_43 (O_43,N_23906,N_22463);
and UO_44 (O_44,N_22574,N_18940);
or UO_45 (O_45,N_24124,N_22195);
and UO_46 (O_46,N_24853,N_18823);
or UO_47 (O_47,N_24668,N_22164);
and UO_48 (O_48,N_22236,N_22893);
nand UO_49 (O_49,N_23399,N_19783);
xor UO_50 (O_50,N_22226,N_23234);
or UO_51 (O_51,N_24874,N_22382);
xnor UO_52 (O_52,N_22532,N_24186);
nor UO_53 (O_53,N_18977,N_19772);
nor UO_54 (O_54,N_20558,N_19441);
or UO_55 (O_55,N_24702,N_22165);
nand UO_56 (O_56,N_24189,N_22363);
nor UO_57 (O_57,N_24510,N_24550);
and UO_58 (O_58,N_21737,N_18906);
and UO_59 (O_59,N_19171,N_20431);
nor UO_60 (O_60,N_24414,N_23289);
nand UO_61 (O_61,N_19264,N_20473);
xnor UO_62 (O_62,N_23508,N_19630);
or UO_63 (O_63,N_20607,N_19686);
nor UO_64 (O_64,N_23296,N_23800);
xnor UO_65 (O_65,N_19434,N_21272);
or UO_66 (O_66,N_19989,N_24651);
nor UO_67 (O_67,N_21680,N_23328);
and UO_68 (O_68,N_24102,N_22377);
nand UO_69 (O_69,N_20947,N_23011);
and UO_70 (O_70,N_19012,N_18774);
and UO_71 (O_71,N_19144,N_19134);
and UO_72 (O_72,N_22865,N_22362);
xor UO_73 (O_73,N_21441,N_22901);
nor UO_74 (O_74,N_19855,N_21200);
xnor UO_75 (O_75,N_23855,N_23271);
and UO_76 (O_76,N_23054,N_22052);
nor UO_77 (O_77,N_21253,N_24231);
and UO_78 (O_78,N_20986,N_21825);
and UO_79 (O_79,N_19310,N_23030);
nor UO_80 (O_80,N_19151,N_24772);
and UO_81 (O_81,N_24653,N_19575);
or UO_82 (O_82,N_22273,N_22462);
nand UO_83 (O_83,N_24543,N_22664);
nor UO_84 (O_84,N_22880,N_19545);
or UO_85 (O_85,N_23253,N_21150);
nand UO_86 (O_86,N_20785,N_19161);
nand UO_87 (O_87,N_22794,N_22656);
and UO_88 (O_88,N_23680,N_24256);
or UO_89 (O_89,N_24147,N_20108);
nor UO_90 (O_90,N_20510,N_23833);
and UO_91 (O_91,N_19771,N_20337);
nand UO_92 (O_92,N_20367,N_18942);
and UO_93 (O_93,N_21973,N_19821);
nand UO_94 (O_94,N_18963,N_22375);
nor UO_95 (O_95,N_23297,N_23498);
or UO_96 (O_96,N_22827,N_23053);
nand UO_97 (O_97,N_23035,N_21947);
and UO_98 (O_98,N_20890,N_20078);
nor UO_99 (O_99,N_20856,N_22379);
and UO_100 (O_100,N_23349,N_23924);
or UO_101 (O_101,N_24218,N_24867);
and UO_102 (O_102,N_19488,N_23424);
nor UO_103 (O_103,N_21537,N_22124);
or UO_104 (O_104,N_24321,N_21754);
and UO_105 (O_105,N_20342,N_21466);
nor UO_106 (O_106,N_20427,N_21018);
or UO_107 (O_107,N_19979,N_20376);
nor UO_108 (O_108,N_19882,N_18845);
and UO_109 (O_109,N_22270,N_24983);
nor UO_110 (O_110,N_22971,N_23616);
nor UO_111 (O_111,N_22097,N_21432);
or UO_112 (O_112,N_24126,N_22762);
nand UO_113 (O_113,N_23149,N_23392);
nand UO_114 (O_114,N_21114,N_20677);
nor UO_115 (O_115,N_23061,N_21775);
nand UO_116 (O_116,N_22255,N_22113);
nand UO_117 (O_117,N_24869,N_23344);
and UO_118 (O_118,N_20535,N_23997);
nor UO_119 (O_119,N_22450,N_24378);
or UO_120 (O_120,N_20534,N_24599);
nand UO_121 (O_121,N_22291,N_19963);
nand UO_122 (O_122,N_21778,N_18751);
nor UO_123 (O_123,N_24302,N_18800);
nor UO_124 (O_124,N_24544,N_18783);
nor UO_125 (O_125,N_22607,N_23766);
and UO_126 (O_126,N_24255,N_24684);
and UO_127 (O_127,N_24066,N_21634);
or UO_128 (O_128,N_19403,N_21969);
or UO_129 (O_129,N_21449,N_22025);
nand UO_130 (O_130,N_23884,N_21565);
xor UO_131 (O_131,N_20476,N_24394);
or UO_132 (O_132,N_23790,N_21454);
nand UO_133 (O_133,N_23904,N_22814);
or UO_134 (O_134,N_20467,N_20968);
and UO_135 (O_135,N_20432,N_23059);
and UO_136 (O_136,N_19820,N_21361);
and UO_137 (O_137,N_24665,N_19166);
nand UO_138 (O_138,N_19765,N_19459);
or UO_139 (O_139,N_24467,N_22512);
nand UO_140 (O_140,N_19365,N_20725);
nor UO_141 (O_141,N_24024,N_24208);
nand UO_142 (O_142,N_19827,N_19064);
nand UO_143 (O_143,N_19863,N_21315);
nor UO_144 (O_144,N_21267,N_21885);
and UO_145 (O_145,N_18958,N_23429);
or UO_146 (O_146,N_20485,N_21757);
nor UO_147 (O_147,N_23147,N_20949);
nand UO_148 (O_148,N_20197,N_23759);
or UO_149 (O_149,N_22083,N_20615);
nor UO_150 (O_150,N_20798,N_21077);
xor UO_151 (O_151,N_24221,N_21148);
and UO_152 (O_152,N_21620,N_19234);
or UO_153 (O_153,N_21044,N_23968);
and UO_154 (O_154,N_19032,N_24447);
and UO_155 (O_155,N_19251,N_24073);
nor UO_156 (O_156,N_19439,N_21618);
and UO_157 (O_157,N_22400,N_24490);
or UO_158 (O_158,N_19096,N_22873);
nand UO_159 (O_159,N_24607,N_22932);
or UO_160 (O_160,N_21256,N_23547);
and UO_161 (O_161,N_22636,N_20632);
nor UO_162 (O_162,N_18891,N_19074);
or UO_163 (O_163,N_24276,N_23376);
and UO_164 (O_164,N_21437,N_23890);
xor UO_165 (O_165,N_23306,N_20219);
nor UO_166 (O_166,N_24751,N_20727);
xnor UO_167 (O_167,N_23269,N_24194);
xor UO_168 (O_168,N_22397,N_22819);
nor UO_169 (O_169,N_19031,N_21401);
or UO_170 (O_170,N_22368,N_19008);
or UO_171 (O_171,N_19217,N_23258);
and UO_172 (O_172,N_22925,N_24188);
nand UO_173 (O_173,N_19726,N_22623);
or UO_174 (O_174,N_20954,N_23136);
and UO_175 (O_175,N_24369,N_24747);
nor UO_176 (O_176,N_24131,N_21731);
and UO_177 (O_177,N_20043,N_21918);
or UO_178 (O_178,N_20580,N_21497);
or UO_179 (O_179,N_21312,N_20422);
or UO_180 (O_180,N_20820,N_23368);
and UO_181 (O_181,N_20430,N_19076);
or UO_182 (O_182,N_21597,N_21727);
nand UO_183 (O_183,N_23068,N_21222);
and UO_184 (O_184,N_21021,N_20133);
or UO_185 (O_185,N_20888,N_23236);
nor UO_186 (O_186,N_21560,N_21246);
or UO_187 (O_187,N_20600,N_23599);
xnor UO_188 (O_188,N_21330,N_19174);
nand UO_189 (O_189,N_20814,N_18788);
and UO_190 (O_190,N_22565,N_21755);
nand UO_191 (O_191,N_21208,N_24775);
and UO_192 (O_192,N_23241,N_22012);
and UO_193 (O_193,N_24390,N_21343);
nor UO_194 (O_194,N_24906,N_20841);
nand UO_195 (O_195,N_19362,N_20216);
or UO_196 (O_196,N_24205,N_20598);
xnor UO_197 (O_197,N_21643,N_21666);
and UO_198 (O_198,N_22289,N_19105);
or UO_199 (O_199,N_19925,N_20316);
nor UO_200 (O_200,N_22688,N_21004);
nand UO_201 (O_201,N_22320,N_19854);
nor UO_202 (O_202,N_24667,N_19499);
and UO_203 (O_203,N_24562,N_23079);
xnor UO_204 (O_204,N_21983,N_20314);
nor UO_205 (O_205,N_23738,N_24725);
xnor UO_206 (O_206,N_19624,N_22224);
nand UO_207 (O_207,N_19707,N_23692);
nor UO_208 (O_208,N_22453,N_23503);
or UO_209 (O_209,N_23350,N_21398);
or UO_210 (O_210,N_22758,N_19535);
nand UO_211 (O_211,N_22054,N_20399);
nand UO_212 (O_212,N_19357,N_20678);
nand UO_213 (O_213,N_23808,N_19639);
nor UO_214 (O_214,N_20882,N_24076);
and UO_215 (O_215,N_21979,N_20803);
nor UO_216 (O_216,N_20696,N_21341);
nand UO_217 (O_217,N_20149,N_22437);
nor UO_218 (O_218,N_20531,N_19766);
and UO_219 (O_219,N_19822,N_20362);
and UO_220 (O_220,N_23103,N_23849);
and UO_221 (O_221,N_22634,N_23323);
nor UO_222 (O_222,N_18895,N_19001);
or UO_223 (O_223,N_22132,N_18883);
and UO_224 (O_224,N_19973,N_20952);
nor UO_225 (O_225,N_21425,N_19652);
or UO_226 (O_226,N_23173,N_20795);
or UO_227 (O_227,N_20384,N_19163);
nand UO_228 (O_228,N_21135,N_20829);
nand UO_229 (O_229,N_21237,N_18874);
nor UO_230 (O_230,N_24998,N_19648);
and UO_231 (O_231,N_24041,N_20223);
nand UO_232 (O_232,N_20157,N_18873);
xnor UO_233 (O_233,N_21418,N_21043);
nor UO_234 (O_234,N_22000,N_19106);
nand UO_235 (O_235,N_21803,N_20714);
or UO_236 (O_236,N_21507,N_21840);
or UO_237 (O_237,N_24079,N_19280);
and UO_238 (O_238,N_22020,N_18993);
nand UO_239 (O_239,N_22352,N_24252);
nor UO_240 (O_240,N_23724,N_19103);
xor UO_241 (O_241,N_21945,N_24129);
and UO_242 (O_242,N_21522,N_24848);
nor UO_243 (O_243,N_19967,N_20466);
xnor UO_244 (O_244,N_22486,N_23438);
and UO_245 (O_245,N_21877,N_18914);
nand UO_246 (O_246,N_19446,N_21961);
or UO_247 (O_247,N_21988,N_22194);
nor UO_248 (O_248,N_24555,N_20609);
nor UO_249 (O_249,N_19849,N_20769);
nor UO_250 (O_250,N_23185,N_22922);
nor UO_251 (O_251,N_19522,N_19311);
nor UO_252 (O_252,N_22065,N_22073);
nand UO_253 (O_253,N_23390,N_22214);
nor UO_254 (O_254,N_19307,N_22072);
nand UO_255 (O_255,N_22337,N_20900);
and UO_256 (O_256,N_21818,N_23412);
nor UO_257 (O_257,N_22848,N_24410);
nand UO_258 (O_258,N_21248,N_21156);
or UO_259 (O_259,N_20461,N_18839);
nor UO_260 (O_260,N_19237,N_21117);
and UO_261 (O_261,N_19406,N_22168);
nand UO_262 (O_262,N_24416,N_21911);
nor UO_263 (O_263,N_22093,N_21532);
and UO_264 (O_264,N_20731,N_22243);
or UO_265 (O_265,N_19690,N_20086);
nor UO_266 (O_266,N_23112,N_23596);
or UO_267 (O_267,N_19469,N_24105);
and UO_268 (O_268,N_20603,N_24994);
xor UO_269 (O_269,N_22745,N_22200);
nand UO_270 (O_270,N_24827,N_21500);
or UO_271 (O_271,N_18868,N_23470);
nand UO_272 (O_272,N_24572,N_23229);
or UO_273 (O_273,N_19687,N_20258);
or UO_274 (O_274,N_24293,N_20937);
xnor UO_275 (O_275,N_22185,N_23211);
or UO_276 (O_276,N_20174,N_20028);
or UO_277 (O_277,N_21240,N_21711);
nand UO_278 (O_278,N_24083,N_18784);
and UO_279 (O_279,N_20396,N_23711);
and UO_280 (O_280,N_20410,N_24303);
nor UO_281 (O_281,N_24438,N_22519);
or UO_282 (O_282,N_23100,N_19538);
or UO_283 (O_283,N_21359,N_22081);
xnor UO_284 (O_284,N_24260,N_19627);
xor UO_285 (O_285,N_21869,N_20853);
nor UO_286 (O_286,N_19711,N_19470);
nor UO_287 (O_287,N_21713,N_19879);
or UO_288 (O_288,N_22468,N_22562);
xnor UO_289 (O_289,N_18804,N_20892);
and UO_290 (O_290,N_19740,N_21798);
nor UO_291 (O_291,N_19894,N_23619);
or UO_292 (O_292,N_21893,N_23868);
and UO_293 (O_293,N_22945,N_22395);
nor UO_294 (O_294,N_23706,N_20106);
and UO_295 (O_295,N_22259,N_19988);
or UO_296 (O_296,N_23110,N_20530);
and UO_297 (O_297,N_22638,N_20266);
or UO_298 (O_298,N_23974,N_19278);
nor UO_299 (O_299,N_19729,N_21685);
xnor UO_300 (O_300,N_19125,N_22415);
or UO_301 (O_301,N_21334,N_23860);
nor UO_302 (O_302,N_20226,N_22631);
nor UO_303 (O_303,N_21704,N_23315);
or UO_304 (O_304,N_23278,N_23001);
nand UO_305 (O_305,N_22692,N_22926);
nor UO_306 (O_306,N_24581,N_19069);
xor UO_307 (O_307,N_19492,N_18997);
and UO_308 (O_308,N_20275,N_24103);
and UO_309 (O_309,N_19068,N_19444);
nor UO_310 (O_310,N_18773,N_23774);
nor UO_311 (O_311,N_20959,N_21473);
nor UO_312 (O_312,N_19270,N_19955);
and UO_313 (O_313,N_24613,N_23685);
or UO_314 (O_314,N_21699,N_22171);
or UO_315 (O_315,N_22152,N_24583);
and UO_316 (O_316,N_23891,N_19188);
xnor UO_317 (O_317,N_20298,N_23076);
nor UO_318 (O_318,N_20179,N_19142);
nand UO_319 (O_319,N_20681,N_22406);
and UO_320 (O_320,N_20493,N_21419);
and UO_321 (O_321,N_19300,N_20009);
nand UO_322 (O_322,N_23769,N_21871);
xnor UO_323 (O_323,N_24729,N_20919);
nand UO_324 (O_324,N_24898,N_21821);
nand UO_325 (O_325,N_23947,N_19655);
or UO_326 (O_326,N_21087,N_21631);
and UO_327 (O_327,N_20335,N_20006);
nor UO_328 (O_328,N_23670,N_20453);
nor UO_329 (O_329,N_19601,N_23395);
nand UO_330 (O_330,N_23535,N_19333);
nand UO_331 (O_331,N_21673,N_21576);
xor UO_332 (O_332,N_21463,N_19508);
nand UO_333 (O_333,N_24488,N_21162);
or UO_334 (O_334,N_20479,N_22475);
nand UO_335 (O_335,N_22888,N_23239);
xor UO_336 (O_336,N_21041,N_24812);
nor UO_337 (O_337,N_24249,N_24914);
or UO_338 (O_338,N_20104,N_22583);
nand UO_339 (O_339,N_22546,N_22300);
or UO_340 (O_340,N_23178,N_22197);
nor UO_341 (O_341,N_20261,N_24709);
nand UO_342 (O_342,N_21684,N_20946);
nand UO_343 (O_343,N_20733,N_23594);
nor UO_344 (O_344,N_20380,N_21534);
xor UO_345 (O_345,N_20767,N_22543);
and UO_346 (O_346,N_20903,N_19285);
xnor UO_347 (O_347,N_24346,N_21442);
nand UO_348 (O_348,N_23862,N_19341);
nand UO_349 (O_349,N_19897,N_20593);
nor UO_350 (O_350,N_20469,N_24769);
or UO_351 (O_351,N_23656,N_21622);
xnor UO_352 (O_352,N_24844,N_19301);
nand UO_353 (O_353,N_21874,N_24866);
nand UO_354 (O_354,N_24929,N_21313);
nand UO_355 (O_355,N_20322,N_24014);
or UO_356 (O_356,N_19225,N_22680);
and UO_357 (O_357,N_18984,N_23140);
xor UO_358 (O_358,N_24856,N_24800);
and UO_359 (O_359,N_22737,N_24548);
nor UO_360 (O_360,N_23827,N_23156);
and UO_361 (O_361,N_20310,N_19862);
nor UO_362 (O_362,N_22521,N_19034);
or UO_363 (O_363,N_22325,N_20827);
nand UO_364 (O_364,N_24404,N_19672);
and UO_365 (O_365,N_23322,N_24923);
nor UO_366 (O_366,N_20684,N_18875);
nand UO_367 (O_367,N_23530,N_20782);
or UO_368 (O_368,N_20450,N_20819);
or UO_369 (O_369,N_24831,N_24415);
or UO_370 (O_370,N_23727,N_22728);
xor UO_371 (O_371,N_23932,N_21963);
and UO_372 (O_372,N_22316,N_18848);
xnor UO_373 (O_373,N_24662,N_24068);
xnor UO_374 (O_374,N_21116,N_19104);
nand UO_375 (O_375,N_21245,N_23431);
nand UO_376 (O_376,N_22896,N_21306);
or UO_377 (O_377,N_21796,N_23946);
or UO_378 (O_378,N_21994,N_23374);
nand UO_379 (O_379,N_22269,N_22323);
nor UO_380 (O_380,N_19788,N_19908);
or UO_381 (O_381,N_23542,N_21736);
nand UO_382 (O_382,N_22770,N_20207);
xor UO_383 (O_383,N_24806,N_19175);
nor UO_384 (O_384,N_24095,N_23175);
nand UO_385 (O_385,N_24871,N_21502);
nand UO_386 (O_386,N_21629,N_24462);
xnor UO_387 (O_387,N_19211,N_24008);
or UO_388 (O_388,N_22454,N_24770);
nand UO_389 (O_389,N_21904,N_24495);
or UO_390 (O_390,N_21277,N_20491);
or UO_391 (O_391,N_20242,N_22934);
and UO_392 (O_392,N_21168,N_20039);
and UO_393 (O_393,N_23473,N_24383);
nand UO_394 (O_394,N_19616,N_22045);
nor UO_395 (O_395,N_20134,N_19465);
and UO_396 (O_396,N_24431,N_23357);
nand UO_397 (O_397,N_19778,N_20200);
nor UO_398 (O_398,N_24071,N_22974);
xnor UO_399 (O_399,N_20280,N_19515);
and UO_400 (O_400,N_19255,N_21601);
and UO_401 (O_401,N_20748,N_22817);
nand UO_402 (O_402,N_20867,N_22201);
and UO_403 (O_403,N_24003,N_20391);
nand UO_404 (O_404,N_19107,N_20998);
or UO_405 (O_405,N_19838,N_24969);
xor UO_406 (O_406,N_19723,N_24327);
or UO_407 (O_407,N_19329,N_22660);
xnor UO_408 (O_408,N_24408,N_24262);
or UO_409 (O_409,N_21131,N_23179);
nand UO_410 (O_410,N_23734,N_24780);
xnor UO_411 (O_411,N_20876,N_21109);
or UO_412 (O_412,N_20447,N_19699);
nor UO_413 (O_413,N_23606,N_22975);
or UO_414 (O_414,N_20750,N_19643);
nor UO_415 (O_415,N_23259,N_19885);
nand UO_416 (O_416,N_24444,N_23397);
or UO_417 (O_417,N_19927,N_19874);
or UO_418 (O_418,N_24093,N_24726);
or UO_419 (O_419,N_23139,N_22568);
or UO_420 (O_420,N_20248,N_22834);
nor UO_421 (O_421,N_20175,N_23984);
nor UO_422 (O_422,N_24403,N_19947);
nor UO_423 (O_423,N_24591,N_20113);
nor UO_424 (O_424,N_19445,N_19347);
nand UO_425 (O_425,N_24554,N_19847);
nand UO_426 (O_426,N_22078,N_20703);
or UO_427 (O_427,N_24267,N_23252);
nand UO_428 (O_428,N_23021,N_23480);
xnor UO_429 (O_429,N_22069,N_24391);
or UO_430 (O_430,N_22742,N_23064);
and UO_431 (O_431,N_19618,N_24948);
nand UO_432 (O_432,N_21280,N_23235);
and UO_433 (O_433,N_19923,N_19569);
or UO_434 (O_434,N_22866,N_21627);
nor UO_435 (O_435,N_21420,N_20165);
nor UO_436 (O_436,N_23008,N_18816);
or UO_437 (O_437,N_22869,N_24698);
or UO_438 (O_438,N_19845,N_22264);
xor UO_439 (O_439,N_23505,N_19764);
nor UO_440 (O_440,N_19016,N_23280);
xnor UO_441 (O_441,N_24900,N_21917);
or UO_442 (O_442,N_20424,N_19604);
nor UO_443 (O_443,N_19516,N_23255);
and UO_444 (O_444,N_21777,N_23115);
nor UO_445 (O_445,N_23543,N_24190);
nand UO_446 (O_446,N_23639,N_18785);
nand UO_447 (O_447,N_20548,N_18930);
nand UO_448 (O_448,N_24759,N_20771);
nand UO_449 (O_449,N_23970,N_23497);
and UO_450 (O_450,N_23799,N_21789);
and UO_451 (O_451,N_20245,N_21366);
xnor UO_452 (O_452,N_18901,N_24044);
nor UO_453 (O_453,N_21672,N_19331);
or UO_454 (O_454,N_23561,N_24811);
or UO_455 (O_455,N_20652,N_19252);
and UO_456 (O_456,N_18948,N_20796);
and UO_457 (O_457,N_22186,N_24470);
nand UO_458 (O_458,N_24485,N_19547);
xor UO_459 (O_459,N_19412,N_23483);
and UO_460 (O_460,N_20972,N_23363);
and UO_461 (O_461,N_24097,N_24807);
and UO_462 (O_462,N_21567,N_22743);
nor UO_463 (O_463,N_22145,N_24904);
nor UO_464 (O_464,N_20000,N_18910);
or UO_465 (O_465,N_23513,N_20791);
xor UO_466 (O_466,N_22891,N_20255);
nor UO_467 (O_467,N_24435,N_20260);
and UO_468 (O_468,N_24781,N_22077);
nor UO_469 (O_469,N_20507,N_19570);
and UO_470 (O_470,N_19123,N_22241);
and UO_471 (O_471,N_24642,N_24878);
nand UO_472 (O_472,N_18990,N_19548);
or UO_473 (O_473,N_21962,N_24821);
nor UO_474 (O_474,N_19004,N_24861);
nor UO_475 (O_475,N_20568,N_23251);
and UO_476 (O_476,N_22855,N_22882);
or UO_477 (O_477,N_20650,N_21323);
and UO_478 (O_478,N_20709,N_20764);
or UO_479 (O_479,N_24964,N_24582);
nand UO_480 (O_480,N_24401,N_22603);
or UO_481 (O_481,N_21065,N_23165);
or UO_482 (O_482,N_22258,N_20222);
and UO_483 (O_483,N_20336,N_22338);
nor UO_484 (O_484,N_20922,N_19842);
nand UO_485 (O_485,N_21851,N_23441);
and UO_486 (O_486,N_24320,N_19033);
and UO_487 (O_487,N_20735,N_18992);
or UO_488 (O_488,N_24398,N_19473);
nand UO_489 (O_489,N_22723,N_20127);
or UO_490 (O_490,N_24484,N_23710);
xnor UO_491 (O_491,N_22591,N_22147);
nand UO_492 (O_492,N_24818,N_20390);
and UO_493 (O_493,N_19706,N_23534);
or UO_494 (O_494,N_23773,N_22380);
nor UO_495 (O_495,N_20169,N_20073);
nor UO_496 (O_496,N_22438,N_21679);
nand UO_497 (O_497,N_22417,N_19905);
or UO_498 (O_498,N_23885,N_22604);
nor UO_499 (O_499,N_23916,N_19191);
or UO_500 (O_500,N_19019,N_23944);
nor UO_501 (O_501,N_21436,N_24739);
or UO_502 (O_502,N_22238,N_19119);
nand UO_503 (O_503,N_24509,N_23340);
or UO_504 (O_504,N_19055,N_20184);
nor UO_505 (O_505,N_22027,N_23647);
and UO_506 (O_506,N_19079,N_23214);
nor UO_507 (O_507,N_23451,N_20309);
nand UO_508 (O_508,N_22313,N_23071);
and UO_509 (O_509,N_23638,N_24937);
or UO_510 (O_510,N_22297,N_20465);
and UO_511 (O_511,N_23133,N_23143);
xor UO_512 (O_512,N_21824,N_20706);
and UO_513 (O_513,N_19865,N_23287);
or UO_514 (O_514,N_19659,N_19295);
and UO_515 (O_515,N_23915,N_21588);
nor UO_516 (O_516,N_21722,N_20938);
and UO_517 (O_517,N_20406,N_18982);
or UO_518 (O_518,N_19363,N_23264);
and UO_519 (O_519,N_21863,N_20690);
and UO_520 (O_520,N_20893,N_22480);
xor UO_521 (O_521,N_21147,N_20514);
and UO_522 (O_522,N_19760,N_21086);
and UO_523 (O_523,N_19725,N_23500);
nor UO_524 (O_524,N_24450,N_22425);
nor UO_525 (O_525,N_23669,N_22955);
nand UO_526 (O_526,N_24840,N_21104);
nor UO_527 (O_527,N_21268,N_23248);
xnor UO_528 (O_528,N_19994,N_21225);
nand UO_529 (O_529,N_23592,N_22451);
xnor UO_530 (O_530,N_22625,N_23465);
nand UO_531 (O_531,N_20092,N_23621);
or UO_532 (O_532,N_19614,N_22879);
or UO_533 (O_533,N_20717,N_23474);
nor UO_534 (O_534,N_22181,N_21668);
nand UO_535 (O_535,N_19611,N_22252);
and UO_536 (O_536,N_24342,N_21040);
nand UO_537 (O_537,N_24338,N_19399);
nor UO_538 (O_538,N_21063,N_21066);
or UO_539 (O_539,N_23476,N_24784);
xor UO_540 (O_540,N_24380,N_24692);
and UO_541 (O_541,N_18976,N_21089);
or UO_542 (O_542,N_22327,N_18912);
nand UO_543 (O_543,N_23955,N_21855);
nand UO_544 (O_544,N_23782,N_23148);
nand UO_545 (O_545,N_21886,N_19197);
nor UO_546 (O_546,N_24215,N_21281);
or UO_547 (O_547,N_21378,N_20776);
and UO_548 (O_548,N_23486,N_23370);
or UO_549 (O_549,N_20926,N_19158);
nor UO_550 (O_550,N_22153,N_19433);
nand UO_551 (O_551,N_23080,N_22047);
nand UO_552 (O_552,N_23583,N_24138);
or UO_553 (O_553,N_21585,N_18972);
nor UO_554 (O_554,N_24005,N_23440);
or UO_555 (O_555,N_21787,N_18934);
nand UO_556 (O_556,N_24296,N_21670);
or UO_557 (O_557,N_23950,N_19758);
and UO_558 (O_558,N_22487,N_19789);
nand UO_559 (O_559,N_21830,N_22393);
or UO_560 (O_560,N_19467,N_21311);
and UO_561 (O_561,N_24620,N_24991);
and UO_562 (O_562,N_20458,N_19792);
nand UO_563 (O_563,N_23401,N_18792);
xor UO_564 (O_564,N_20992,N_22948);
nand UO_565 (O_565,N_23776,N_18878);
xnor UO_566 (O_566,N_21397,N_19284);
and UO_567 (O_567,N_22614,N_23307);
nor UO_568 (O_568,N_22976,N_21235);
xnor UO_569 (O_569,N_23332,N_24084);
or UO_570 (O_570,N_19996,N_21297);
or UO_571 (O_571,N_24178,N_21897);
nor UO_572 (O_572,N_22018,N_23797);
or UO_573 (O_573,N_24713,N_24370);
nor UO_574 (O_574,N_24616,N_18824);
nand UO_575 (O_575,N_22778,N_22191);
nand UO_576 (O_576,N_20445,N_22211);
or UO_577 (O_577,N_22531,N_22346);
or UO_578 (O_578,N_19198,N_20647);
and UO_579 (O_579,N_20645,N_22391);
and UO_580 (O_580,N_20060,N_22502);
nor UO_581 (O_581,N_23137,N_22701);
and UO_582 (O_582,N_20357,N_19534);
nor UO_583 (O_583,N_21515,N_20741);
nor UO_584 (O_584,N_24858,N_21860);
nand UO_585 (O_585,N_24714,N_20942);
or UO_586 (O_586,N_22898,N_23060);
nand UO_587 (O_587,N_21260,N_22629);
nand UO_588 (O_588,N_18944,N_18936);
nand UO_589 (O_589,N_19083,N_21834);
and UO_590 (O_590,N_24718,N_21001);
or UO_591 (O_591,N_24972,N_24743);
nor UO_592 (O_592,N_19316,N_24247);
or UO_593 (O_593,N_22253,N_22996);
or UO_594 (O_594,N_19109,N_19401);
xnor UO_595 (O_595,N_20022,N_21467);
or UO_596 (O_596,N_18952,N_22445);
nor UO_597 (O_597,N_22878,N_20192);
and UO_598 (O_598,N_21265,N_23865);
nand UO_599 (O_599,N_19313,N_24314);
nand UO_600 (O_600,N_21157,N_22564);
or UO_601 (O_601,N_22263,N_20871);
or UO_602 (O_602,N_21603,N_22430);
nor UO_603 (O_603,N_19933,N_19146);
or UO_604 (O_604,N_18885,N_23341);
and UO_605 (O_605,N_24472,N_19010);
xor UO_606 (O_606,N_21472,N_21557);
and UO_607 (O_607,N_24285,N_22821);
or UO_608 (O_608,N_19828,N_22122);
and UO_609 (O_609,N_22572,N_20557);
or UO_610 (O_610,N_19246,N_22340);
and UO_611 (O_611,N_22578,N_23750);
xnor UO_612 (O_612,N_20065,N_21141);
or UO_613 (O_613,N_24516,N_24949);
and UO_614 (O_614,N_20276,N_19386);
and UO_615 (O_615,N_20910,N_22037);
or UO_616 (O_616,N_19641,N_19914);
nand UO_617 (O_617,N_24566,N_22130);
and UO_618 (O_618,N_24274,N_20295);
and UO_619 (O_619,N_22852,N_19554);
xor UO_620 (O_620,N_22677,N_24437);
xor UO_621 (O_621,N_21481,N_23533);
or UO_622 (O_622,N_23277,N_20930);
nor UO_623 (O_623,N_22344,N_20299);
and UO_624 (O_624,N_19898,N_20833);
or UO_625 (O_625,N_20752,N_23002);
or UO_626 (O_626,N_19830,N_24166);
and UO_627 (O_627,N_24728,N_23830);
xnor UO_628 (O_628,N_22429,N_23284);
nand UO_629 (O_629,N_18796,N_19065);
nor UO_630 (O_630,N_24312,N_18809);
nor UO_631 (O_631,N_22530,N_23366);
or UO_632 (O_632,N_18991,N_19635);
nor UO_633 (O_633,N_23817,N_20783);
and UO_634 (O_634,N_21295,N_23646);
nand UO_635 (O_635,N_20264,N_21412);
nor UO_636 (O_636,N_24637,N_21942);
and UO_637 (O_637,N_20766,N_19881);
xor UO_638 (O_638,N_21823,N_19322);
nand UO_639 (O_639,N_20208,N_23767);
nor UO_640 (O_640,N_21380,N_23664);
or UO_641 (O_641,N_22061,N_22123);
or UO_642 (O_642,N_24339,N_20063);
and UO_643 (O_643,N_18908,N_24783);
or UO_644 (O_644,N_18820,N_21209);
and UO_645 (O_645,N_21835,N_19887);
nand UO_646 (O_646,N_21870,N_21527);
nor UO_647 (O_647,N_24371,N_20317);
or UO_648 (O_648,N_21645,N_19588);
or UO_649 (O_649,N_19733,N_19793);
xor UO_650 (O_650,N_21199,N_21032);
nand UO_651 (O_651,N_22515,N_22353);
nor UO_652 (O_652,N_23723,N_19348);
and UO_653 (O_653,N_20421,N_24966);
nand UO_654 (O_654,N_23744,N_21671);
nor UO_655 (O_655,N_19179,N_22220);
and UO_656 (O_656,N_20232,N_20468);
nand UO_657 (O_657,N_21817,N_23293);
or UO_658 (O_658,N_21966,N_22514);
nor UO_659 (O_659,N_21039,N_20544);
xnor UO_660 (O_660,N_24456,N_23210);
nor UO_661 (O_661,N_19853,N_23092);
and UO_662 (O_662,N_18978,N_24909);
nor UO_663 (O_663,N_20662,N_21514);
or UO_664 (O_664,N_21510,N_24749);
or UO_665 (O_665,N_21163,N_19819);
nand UO_666 (O_666,N_21548,N_22212);
nor UO_667 (O_667,N_20551,N_19808);
nand UO_668 (O_668,N_24182,N_19700);
nand UO_669 (O_669,N_23690,N_19558);
and UO_670 (O_670,N_21999,N_19392);
xor UO_671 (O_671,N_21290,N_20331);
and UO_672 (O_672,N_21828,N_23877);
nor UO_673 (O_673,N_22443,N_24082);
or UO_674 (O_674,N_22485,N_20419);
or UO_675 (O_675,N_21456,N_24956);
nor UO_676 (O_676,N_22088,N_23194);
and UO_677 (O_677,N_23158,N_24805);
and UO_678 (O_678,N_19910,N_21657);
and UO_679 (O_679,N_18766,N_21660);
xnor UO_680 (O_680,N_24798,N_18995);
nand UO_681 (O_681,N_20029,N_21512);
and UO_682 (O_682,N_24887,N_22917);
or UO_683 (O_683,N_22653,N_19775);
and UO_684 (O_684,N_19380,N_23435);
nor UO_685 (O_685,N_19461,N_20739);
or UO_686 (O_686,N_22262,N_21298);
xor UO_687 (O_687,N_23801,N_22341);
and UO_688 (O_688,N_21892,N_19029);
xnor UO_689 (O_689,N_23941,N_20212);
and UO_690 (O_690,N_20756,N_22874);
nand UO_691 (O_691,N_22013,N_21201);
and UO_692 (O_692,N_24594,N_23749);
nor UO_693 (O_693,N_22911,N_21216);
nor UO_694 (O_694,N_23952,N_24774);
nand UO_695 (O_695,N_24432,N_18770);
xor UO_696 (O_696,N_21638,N_20692);
nand UO_697 (O_697,N_22918,N_20168);
nor UO_698 (O_698,N_20365,N_22120);
nor UO_699 (O_699,N_21404,N_24675);
nor UO_700 (O_700,N_21831,N_24754);
or UO_701 (O_701,N_18951,N_21765);
and UO_702 (O_702,N_19013,N_22798);
or UO_703 (O_703,N_22501,N_22483);
and UO_704 (O_704,N_24974,N_19248);
nor UO_705 (O_705,N_22099,N_24773);
and UO_706 (O_706,N_24970,N_19187);
nor UO_707 (O_707,N_23661,N_21667);
and UO_708 (O_708,N_22646,N_24671);
and UO_709 (O_709,N_22958,N_22581);
and UO_710 (O_710,N_23917,N_23628);
nand UO_711 (O_711,N_20543,N_19502);
nand UO_712 (O_712,N_24282,N_24640);
and UO_713 (O_713,N_20683,N_21048);
or UO_714 (O_714,N_20228,N_19231);
nor UO_715 (O_715,N_21938,N_20268);
nor UO_716 (O_716,N_19702,N_22085);
or UO_717 (O_717,N_21142,N_20596);
and UO_718 (O_718,N_22560,N_18762);
nor UO_719 (O_719,N_19506,N_19537);
xor UO_720 (O_720,N_20285,N_20250);
and UO_721 (O_721,N_23405,N_19277);
and UO_722 (O_722,N_18897,N_23889);
nand UO_723 (O_723,N_24360,N_20206);
and UO_724 (O_724,N_18867,N_19549);
or UO_725 (O_725,N_22679,N_23093);
and UO_726 (O_726,N_20737,N_22471);
nor UO_727 (O_727,N_23755,N_20941);
nor UO_728 (O_728,N_20762,N_21457);
or UO_729 (O_729,N_20553,N_21368);
or UO_730 (O_730,N_22863,N_19839);
and UO_731 (O_731,N_18983,N_23490);
and UO_732 (O_732,N_21365,N_22472);
or UO_733 (O_733,N_19372,N_19952);
or UO_734 (O_734,N_23678,N_23192);
nor UO_735 (O_735,N_20987,N_19113);
or UO_736 (O_736,N_24968,N_19695);
xnor UO_737 (O_737,N_24946,N_24722);
xor UO_738 (O_738,N_21173,N_19663);
and UO_739 (O_739,N_20573,N_22548);
or UO_740 (O_740,N_19156,N_21948);
nand UO_741 (O_741,N_19637,N_24741);
and UO_742 (O_742,N_23981,N_22232);
or UO_743 (O_743,N_23560,N_20560);
nor UO_744 (O_744,N_21852,N_21197);
nand UO_745 (O_745,N_24851,N_22260);
nor UO_746 (O_746,N_21319,N_23085);
or UO_747 (O_747,N_23449,N_21762);
nor UO_748 (O_748,N_24064,N_23607);
or UO_749 (O_749,N_19520,N_20701);
and UO_750 (O_750,N_24571,N_24624);
or UO_751 (O_751,N_22754,N_18923);
or UO_752 (O_752,N_24281,N_22448);
nand UO_753 (O_753,N_19982,N_22700);
or UO_754 (O_754,N_19160,N_20225);
nand UO_755 (O_755,N_22999,N_20425);
and UO_756 (O_756,N_21078,N_20685);
xnor UO_757 (O_757,N_24372,N_20492);
xor UO_758 (O_758,N_22972,N_22785);
or UO_759 (O_759,N_19122,N_22993);
and UO_760 (O_760,N_24348,N_22727);
and UO_761 (O_761,N_21730,N_18870);
nor UO_762 (O_762,N_23373,N_24719);
xor UO_763 (O_763,N_18959,N_21405);
xor UO_764 (O_764,N_21990,N_20187);
xnor UO_765 (O_765,N_21625,N_19958);
nor UO_766 (O_766,N_19903,N_24204);
xnor UO_767 (O_767,N_22577,N_24507);
and UO_768 (O_768,N_22182,N_21783);
or UO_769 (O_769,N_23087,N_21002);
or UO_770 (O_770,N_23733,N_23180);
nor UO_771 (O_771,N_23730,N_19457);
and UO_772 (O_772,N_20383,N_21242);
and UO_773 (O_773,N_19767,N_18863);
xor UO_774 (O_774,N_21493,N_18851);
nand UO_775 (O_775,N_20951,N_19039);
and UO_776 (O_776,N_20997,N_19047);
nor UO_777 (O_777,N_20556,N_24107);
and UO_778 (O_778,N_19038,N_23524);
nand UO_779 (O_779,N_20842,N_22042);
nand UO_780 (O_780,N_24515,N_24824);
xor UO_781 (O_781,N_19671,N_22523);
or UO_782 (O_782,N_24179,N_21664);
xor UO_783 (O_783,N_19373,N_24161);
nand UO_784 (O_784,N_23371,N_24931);
or UO_785 (O_785,N_24452,N_24627);
nand UO_786 (O_786,N_20407,N_20710);
nor UO_787 (O_787,N_23334,N_24421);
or UO_788 (O_788,N_21898,N_23526);
nor UO_789 (O_789,N_21399,N_24834);
nand UO_790 (O_790,N_24682,N_23131);
nand UO_791 (O_791,N_20144,N_24540);
nor UO_792 (O_792,N_18854,N_19460);
and UO_793 (O_793,N_19028,N_21027);
nor UO_794 (O_794,N_23781,N_22280);
xor UO_795 (O_795,N_22095,N_24778);
or UO_796 (O_796,N_23319,N_24436);
nand UO_797 (O_797,N_24661,N_21644);
and UO_798 (O_798,N_20509,N_20502);
nand UO_799 (O_799,N_21022,N_19978);
nor UO_800 (O_800,N_22726,N_19975);
or UO_801 (O_801,N_20105,N_23965);
nand UO_802 (O_802,N_20913,N_21849);
xor UO_803 (O_803,N_24137,N_23267);
or UO_804 (O_804,N_23058,N_19293);
nand UO_805 (O_805,N_19954,N_24108);
xnor UO_806 (O_806,N_19769,N_24689);
and UO_807 (O_807,N_19049,N_19330);
or UO_808 (O_808,N_23856,N_20633);
nand UO_809 (O_809,N_22919,N_19027);
xor UO_810 (O_810,N_23857,N_22455);
and UO_811 (O_811,N_19795,N_22051);
nand UO_812 (O_812,N_20617,N_24409);
nand UO_813 (O_813,N_20613,N_22643);
and UO_814 (O_814,N_19343,N_20030);
and UO_815 (O_815,N_19407,N_19425);
or UO_816 (O_816,N_19089,N_21621);
nor UO_817 (O_817,N_21387,N_20506);
or UO_818 (O_818,N_23098,N_23967);
and UO_819 (O_819,N_23206,N_19296);
and UO_820 (O_820,N_23295,N_19943);
nor UO_821 (O_821,N_21153,N_21703);
nor UO_822 (O_822,N_22597,N_20587);
and UO_823 (O_823,N_21332,N_21592);
or UO_824 (O_824,N_20217,N_19626);
nor UO_825 (O_825,N_19505,N_21422);
xnor UO_826 (O_826,N_21068,N_23375);
or UO_827 (O_827,N_21891,N_22518);
and UO_828 (O_828,N_21888,N_23457);
nor UO_829 (O_829,N_22695,N_20306);
and UO_830 (O_830,N_18864,N_19877);
nand UO_831 (O_831,N_18841,N_23612);
xnor UO_832 (O_832,N_23803,N_20353);
and UO_833 (O_833,N_19024,N_20523);
and UO_834 (O_834,N_21881,N_23822);
or UO_835 (O_835,N_21998,N_21071);
or UO_836 (O_836,N_21128,N_20806);
or UO_837 (O_837,N_20686,N_23292);
nand UO_838 (O_838,N_19561,N_19186);
nor UO_839 (O_839,N_20839,N_19608);
nor UO_840 (O_840,N_18763,N_19632);
nand UO_841 (O_841,N_23130,N_18966);
or UO_842 (O_842,N_22853,N_20786);
nor UO_843 (O_843,N_24389,N_22021);
or UO_844 (O_844,N_24947,N_21321);
and UO_845 (O_845,N_19291,N_19435);
or UO_846 (O_846,N_23823,N_22612);
nor UO_847 (O_847,N_20595,N_23570);
nor UO_848 (O_848,N_24860,N_24647);
nand UO_849 (O_849,N_19836,N_23804);
or UO_850 (O_850,N_22311,N_24349);
and UO_851 (O_851,N_23642,N_22690);
nand UO_852 (O_852,N_19420,N_23208);
nor UO_853 (O_853,N_21314,N_23809);
nand UO_854 (O_854,N_21628,N_24678);
nor UO_855 (O_855,N_23991,N_19215);
or UO_856 (O_856,N_19668,N_23702);
xor UO_857 (O_857,N_23729,N_19888);
nor UO_858 (O_858,N_22730,N_23576);
and UO_859 (O_859,N_20368,N_20477);
or UO_860 (O_860,N_24941,N_22739);
and UO_861 (O_861,N_18962,N_20319);
and UO_862 (O_862,N_21108,N_22101);
or UO_863 (O_863,N_24086,N_19155);
or UO_864 (O_864,N_20505,N_24121);
and UO_865 (O_865,N_24981,N_23337);
and UO_866 (O_866,N_21743,N_23063);
nor UO_867 (O_867,N_24311,N_24738);
nand UO_868 (O_868,N_24644,N_22751);
nor UO_869 (O_869,N_21674,N_20010);
nor UO_870 (O_870,N_24236,N_21637);
nand UO_871 (O_871,N_23899,N_22649);
xor UO_872 (O_872,N_19271,N_20163);
or UO_873 (O_873,N_19841,N_20415);
and UO_874 (O_874,N_22777,N_20302);
and UO_875 (O_875,N_24938,N_21551);
nor UO_876 (O_876,N_21286,N_20932);
nand UO_877 (O_877,N_22491,N_22626);
xor UO_878 (O_878,N_19490,N_21211);
xor UO_879 (O_879,N_24639,N_22167);
or UO_880 (O_880,N_21318,N_21213);
nand UO_881 (O_881,N_22332,N_24541);
xor UO_882 (O_882,N_22141,N_24924);
and UO_883 (O_883,N_18913,N_22796);
and UO_884 (O_884,N_19389,N_24796);
or UO_885 (O_885,N_22178,N_20394);
or UO_886 (O_886,N_22870,N_24576);
and UO_887 (O_887,N_22533,N_19139);
nand UO_888 (O_888,N_20896,N_24020);
and UO_889 (O_889,N_22389,N_21198);
and UO_890 (O_890,N_20788,N_19292);
and UO_891 (O_891,N_23335,N_24043);
and UO_892 (O_892,N_21850,N_23786);
xor UO_893 (O_893,N_24618,N_19649);
nand UO_894 (O_894,N_19199,N_19875);
nand UO_895 (O_895,N_22678,N_21445);
nand UO_896 (O_896,N_24238,N_20115);
or UO_897 (O_897,N_20549,N_23346);
and UO_898 (O_898,N_20720,N_20586);
nand UO_899 (O_899,N_21659,N_21455);
and UO_900 (O_900,N_19577,N_20109);
or UO_901 (O_901,N_19196,N_19646);
or UO_902 (O_902,N_19193,N_22978);
nand UO_903 (O_903,N_22304,N_21697);
nor UO_904 (O_904,N_22931,N_22937);
and UO_905 (O_905,N_22702,N_20525);
nor UO_906 (O_906,N_20744,N_24873);
xor UO_907 (O_907,N_24197,N_22776);
nand UO_908 (O_908,N_24234,N_21140);
xor UO_909 (O_909,N_24951,N_22060);
nor UO_910 (O_910,N_22815,N_19581);
xnor UO_911 (O_911,N_22707,N_20754);
nand UO_912 (O_912,N_19584,N_22528);
nor UO_913 (O_913,N_18828,N_21887);
nor UO_914 (O_914,N_19478,N_21836);
and UO_915 (O_915,N_19235,N_19661);
nor UO_916 (O_916,N_19675,N_21856);
and UO_917 (O_917,N_24092,N_24280);
or UO_918 (O_918,N_23569,N_20437);
and UO_919 (O_919,N_20136,N_21355);
nand UO_920 (O_920,N_22023,N_21270);
xor UO_921 (O_921,N_23820,N_19576);
nor UO_922 (O_922,N_18994,N_20944);
nor UO_923 (O_923,N_21204,N_22150);
nand UO_924 (O_924,N_23051,N_20182);
and UO_925 (O_925,N_19355,N_20864);
nand UO_926 (O_926,N_22160,N_24822);
nand UO_927 (O_927,N_21427,N_21059);
and UO_928 (O_928,N_23310,N_19263);
and UO_929 (O_929,N_19628,N_20813);
xor UO_930 (O_930,N_19168,N_22771);
or UO_931 (O_931,N_20198,N_20822);
nor UO_932 (O_932,N_21868,N_20480);
or UO_933 (O_933,N_19664,N_23520);
or UO_934 (O_934,N_24443,N_18985);
nor UO_935 (O_935,N_19936,N_20273);
or UO_936 (O_936,N_19689,N_20960);
or UO_937 (O_937,N_21926,N_19732);
or UO_938 (O_938,N_19371,N_24057);
xor UO_939 (O_939,N_23426,N_24705);
xnor UO_940 (O_940,N_21747,N_23960);
nand UO_941 (O_941,N_22414,N_18935);
or UO_942 (O_942,N_20312,N_24030);
xor UO_943 (O_943,N_21937,N_23387);
nor UO_944 (O_944,N_21053,N_20224);
and UO_945 (O_945,N_20794,N_22628);
nand UO_946 (O_946,N_24760,N_24522);
or UO_947 (O_947,N_24907,N_24952);
or UO_948 (O_948,N_20486,N_20728);
and UO_949 (O_949,N_21663,N_24217);
and UO_950 (O_950,N_24418,N_24468);
or UO_951 (O_951,N_22864,N_19283);
nand UO_952 (O_952,N_21386,N_24955);
and UO_953 (O_953,N_22119,N_23578);
and UO_954 (O_954,N_23871,N_18896);
or UO_955 (O_955,N_22005,N_22536);
and UO_956 (O_956,N_18876,N_19517);
or UO_957 (O_957,N_23393,N_23645);
or UO_958 (O_958,N_21907,N_24655);
nor UO_959 (O_959,N_23309,N_19086);
nor UO_960 (O_960,N_21139,N_20436);
or UO_961 (O_961,N_19734,N_20318);
nor UO_962 (O_962,N_21600,N_22115);
xor UO_963 (O_963,N_23713,N_19080);
nor UO_964 (O_964,N_20889,N_20046);
or UO_965 (O_965,N_20459,N_24250);
and UO_966 (O_966,N_19804,N_22953);
nor UO_967 (O_967,N_23461,N_18877);
nand UO_968 (O_968,N_24891,N_18819);
nor UO_969 (O_969,N_24894,N_24253);
nor UO_970 (O_970,N_20135,N_20230);
and UO_971 (O_971,N_20267,N_21956);
nor UO_972 (O_972,N_24600,N_20004);
or UO_973 (O_973,N_21015,N_22995);
xor UO_974 (O_974,N_23627,N_20071);
and UO_975 (O_975,N_21508,N_21227);
nor UO_976 (O_976,N_18927,N_23644);
nor UO_977 (O_977,N_19598,N_22404);
nand UO_978 (O_978,N_20571,N_19974);
and UO_979 (O_979,N_20101,N_19705);
and UO_980 (O_980,N_19724,N_24744);
nor UO_981 (O_981,N_23704,N_22198);
nand UO_982 (O_982,N_19281,N_24569);
nand UO_983 (O_983,N_22594,N_20209);
nand UO_984 (O_984,N_21791,N_22102);
nor UO_985 (O_985,N_20978,N_20899);
xor UO_986 (O_986,N_20088,N_20237);
or UO_987 (O_987,N_20278,N_21394);
nor UO_988 (O_988,N_19720,N_22076);
and UO_989 (O_989,N_24460,N_23693);
or UO_990 (O_990,N_20726,N_20590);
and UO_991 (O_991,N_19289,N_21271);
nor UO_992 (O_992,N_21006,N_22118);
nand UO_993 (O_993,N_23077,N_21511);
nand UO_994 (O_994,N_22315,N_23608);
xnor UO_995 (O_995,N_22541,N_24782);
nor UO_996 (O_996,N_20524,N_21951);
nor UO_997 (O_997,N_23939,N_22265);
and UO_998 (O_998,N_23231,N_21347);
nand UO_999 (O_999,N_23870,N_18960);
nand UO_1000 (O_1000,N_23272,N_20800);
xor UO_1001 (O_1001,N_21212,N_23414);
nand UO_1002 (O_1002,N_18752,N_20382);
and UO_1003 (O_1003,N_21291,N_19361);
or UO_1004 (O_1004,N_19790,N_23409);
nor UO_1005 (O_1005,N_20577,N_23568);
or UO_1006 (O_1006,N_23958,N_18888);
and UO_1007 (O_1007,N_24196,N_22750);
nor UO_1008 (O_1008,N_23218,N_23182);
xnor UO_1009 (O_1009,N_20139,N_18953);
or UO_1010 (O_1010,N_23910,N_23434);
and UO_1011 (O_1011,N_24996,N_24170);
and UO_1012 (O_1012,N_23620,N_20405);
nand UO_1013 (O_1013,N_19274,N_19665);
or UO_1014 (O_1014,N_24292,N_20355);
or UO_1015 (O_1015,N_20294,N_24040);
and UO_1016 (O_1016,N_23279,N_20277);
nor UO_1017 (O_1017,N_19157,N_19609);
nor UO_1018 (O_1018,N_19843,N_23394);
nor UO_1019 (O_1019,N_21705,N_22317);
nor UO_1020 (O_1020,N_21615,N_21719);
nand UO_1021 (O_1021,N_20359,N_20973);
or UO_1022 (O_1022,N_22067,N_19226);
and UO_1023 (O_1023,N_22245,N_24503);
and UO_1024 (O_1024,N_19636,N_21683);
and UO_1025 (O_1025,N_21882,N_22615);
nand UO_1026 (O_1026,N_20562,N_21735);
nor UO_1027 (O_1027,N_23453,N_19482);
nand UO_1028 (O_1028,N_24310,N_20122);
nor UO_1029 (O_1029,N_24034,N_21499);
xnor UO_1030 (O_1030,N_24546,N_20044);
or UO_1031 (O_1031,N_22136,N_19325);
nor UO_1032 (O_1032,N_20967,N_23338);
or UO_1033 (O_1033,N_21487,N_23780);
and UO_1034 (O_1034,N_24918,N_23106);
nand UO_1035 (O_1035,N_22580,N_22826);
nor UO_1036 (O_1036,N_21206,N_22192);
nand UO_1037 (O_1037,N_19591,N_21867);
or UO_1038 (O_1038,N_20630,N_21258);
and UO_1039 (O_1039,N_22964,N_24801);
nand UO_1040 (O_1040,N_19244,N_24046);
and UO_1041 (O_1041,N_18866,N_24654);
or UO_1042 (O_1042,N_19745,N_20724);
nor UO_1043 (O_1043,N_18900,N_20026);
xnor UO_1044 (O_1044,N_18753,N_21707);
and UO_1045 (O_1045,N_19907,N_23779);
nand UO_1046 (O_1046,N_24347,N_19901);
or UO_1047 (O_1047,N_23658,N_19261);
or UO_1048 (O_1048,N_19202,N_24802);
or UO_1049 (O_1049,N_22038,N_24636);
or UO_1050 (O_1050,N_20021,N_18826);
or UO_1051 (O_1051,N_22681,N_22170);
nand UO_1052 (O_1052,N_20661,N_18829);
nand UO_1053 (O_1053,N_18881,N_23538);
xnor UO_1054 (O_1054,N_21443,N_23299);
xor UO_1055 (O_1055,N_21526,N_22652);
nand UO_1056 (O_1056,N_20620,N_20943);
or UO_1057 (O_1057,N_24857,N_20643);
nand UO_1058 (O_1058,N_20582,N_19182);
or UO_1059 (O_1059,N_24531,N_19003);
and UO_1060 (O_1060,N_21884,N_21196);
or UO_1061 (O_1061,N_20068,N_20585);
or UO_1062 (O_1062,N_23005,N_20489);
or UO_1063 (O_1063,N_24065,N_24500);
or UO_1064 (O_1064,N_21244,N_24993);
nor UO_1065 (O_1065,N_20080,N_22696);
and UO_1066 (O_1066,N_19479,N_23783);
or UO_1067 (O_1067,N_23551,N_19017);
nor UO_1068 (O_1068,N_22459,N_19861);
xnor UO_1069 (O_1069,N_18987,N_22157);
nand UO_1070 (O_1070,N_21496,N_20854);
or UO_1071 (O_1071,N_23601,N_21203);
nand UO_1072 (O_1072,N_20326,N_19589);
xor UO_1073 (O_1073,N_21076,N_21129);
nand UO_1074 (O_1074,N_23223,N_23510);
and UO_1075 (O_1075,N_19385,N_21194);
nor UO_1076 (O_1076,N_22376,N_24935);
nand UO_1077 (O_1077,N_21528,N_21371);
nand UO_1078 (O_1078,N_22670,N_22446);
or UO_1079 (O_1079,N_22288,N_20772);
and UO_1080 (O_1080,N_20933,N_19629);
and UO_1081 (O_1081,N_19298,N_22139);
or UO_1082 (O_1082,N_23243,N_18973);
nor UO_1083 (O_1083,N_21953,N_24112);
nand UO_1084 (O_1084,N_21007,N_19183);
or UO_1085 (O_1085,N_21047,N_20848);
or UO_1086 (O_1086,N_21636,N_22507);
xor UO_1087 (O_1087,N_20051,N_19148);
nor UO_1088 (O_1088,N_18969,N_21095);
nor UO_1089 (O_1089,N_20745,N_21767);
or UO_1090 (O_1090,N_23655,N_20981);
nand UO_1091 (O_1091,N_22439,N_23124);
nor UO_1092 (O_1092,N_24978,N_21376);
and UO_1093 (O_1093,N_20738,N_20983);
or UO_1094 (O_1094,N_20005,N_23233);
or UO_1095 (O_1095,N_22645,N_23045);
and UO_1096 (O_1096,N_22161,N_23648);
and UO_1097 (O_1097,N_24159,N_24852);
nor UO_1098 (O_1098,N_22110,N_22210);
nor UO_1099 (O_1099,N_19454,N_22465);
nor UO_1100 (O_1100,N_20723,N_24165);
or UO_1101 (O_1101,N_19239,N_23501);
and UO_1102 (O_1102,N_20512,N_21269);
xnor UO_1103 (O_1103,N_22271,N_21461);
xor UO_1104 (O_1104,N_20540,N_21189);
xnor UO_1105 (O_1105,N_22939,N_24643);
or UO_1106 (O_1106,N_23485,N_24111);
nand UO_1107 (O_1107,N_20638,N_23852);
nor UO_1108 (O_1108,N_23649,N_20878);
and UO_1109 (O_1109,N_18818,N_21878);
and UO_1110 (O_1110,N_22427,N_19904);
or UO_1111 (O_1111,N_22409,N_18931);
nand UO_1112 (O_1112,N_23151,N_19484);
and UO_1113 (O_1113,N_24222,N_23456);
xnor UO_1114 (O_1114,N_19676,N_23555);
and UO_1115 (O_1115,N_22774,N_21390);
and UO_1116 (O_1116,N_19014,N_24334);
or UO_1117 (O_1117,N_20555,N_21064);
xnor UO_1118 (O_1118,N_23184,N_24716);
nand UO_1119 (O_1119,N_22461,N_22890);
xor UO_1120 (O_1120,N_23043,N_23864);
xnor UO_1121 (O_1121,N_22921,N_18794);
xor UO_1122 (O_1122,N_23753,N_20032);
and UO_1123 (O_1123,N_19115,N_23634);
nand UO_1124 (O_1124,N_20451,N_20143);
and UO_1125 (O_1125,N_23732,N_24589);
or UO_1126 (O_1126,N_20003,N_23511);
nor UO_1127 (O_1127,N_21014,N_19340);
and UO_1128 (O_1128,N_23304,N_22331);
nand UO_1129 (O_1129,N_19081,N_20648);
nand UO_1130 (O_1130,N_21729,N_23095);
and UO_1131 (O_1131,N_21424,N_24029);
or UO_1132 (O_1132,N_23763,N_19957);
nor UO_1133 (O_1133,N_20463,N_23893);
and UO_1134 (O_1134,N_19823,N_19172);
and UO_1135 (O_1135,N_19007,N_24995);
and UO_1136 (O_1136,N_22303,N_20887);
nor UO_1137 (O_1137,N_20884,N_22234);
nand UO_1138 (O_1138,N_20618,N_21790);
or UO_1139 (O_1139,N_24703,N_22595);
and UO_1140 (O_1140,N_22278,N_19384);
xnor UO_1141 (O_1141,N_21873,N_20048);
and UO_1142 (O_1142,N_20185,N_23957);
nor UO_1143 (O_1143,N_24632,N_22573);
and UO_1144 (O_1144,N_24098,N_20016);
nor UO_1145 (O_1145,N_20700,N_22788);
xor UO_1146 (O_1146,N_22718,N_21275);
nand UO_1147 (O_1147,N_24795,N_23848);
or UO_1148 (O_1148,N_19857,N_19025);
or UO_1149 (O_1149,N_22694,N_19850);
and UO_1150 (O_1150,N_19462,N_20274);
nor UO_1151 (O_1151,N_23174,N_24896);
nand UO_1152 (O_1152,N_19981,N_23937);
or UO_1153 (O_1153,N_22188,N_19455);
and UO_1154 (O_1154,N_20649,N_19993);
or UO_1155 (O_1155,N_23274,N_24748);
nand UO_1156 (O_1156,N_19143,N_23197);
or UO_1157 (O_1157,N_22330,N_24622);
xor UO_1158 (O_1158,N_24828,N_20304);
nor UO_1159 (O_1159,N_22447,N_19260);
or UO_1160 (O_1160,N_20718,N_19848);
and UO_1161 (O_1161,N_22676,N_20401);
nand UO_1162 (O_1162,N_20760,N_21751);
nor UO_1163 (O_1163,N_24373,N_20282);
nor UO_1164 (O_1164,N_18850,N_18790);
or UO_1165 (O_1165,N_19592,N_21495);
and UO_1166 (O_1166,N_22576,N_24560);
nand UO_1167 (O_1167,N_19442,N_23614);
nor UO_1168 (O_1168,N_24610,N_23525);
nand UO_1169 (O_1169,N_24645,N_19423);
nor UO_1170 (O_1170,N_21276,N_22474);
and UO_1171 (O_1171,N_24706,N_20655);
and UO_1172 (O_1172,N_23821,N_23691);
and UO_1173 (O_1173,N_22557,N_19424);
and UO_1174 (O_1174,N_24884,N_22982);
and UO_1175 (O_1175,N_19009,N_21137);
and UO_1176 (O_1176,N_18937,N_20891);
and UO_1177 (O_1177,N_22841,N_19258);
or UO_1178 (O_1178,N_24009,N_19005);
nand UO_1179 (O_1179,N_23940,N_19337);
and UO_1180 (O_1180,N_23798,N_19272);
or UO_1181 (O_1181,N_24711,N_19162);
nand UO_1182 (O_1182,N_24740,N_23736);
nand UO_1183 (O_1183,N_22089,N_18799);
nand UO_1184 (O_1184,N_19794,N_23418);
nor UO_1185 (O_1185,N_21283,N_21045);
or UO_1186 (O_1186,N_24982,N_21093);
nand UO_1187 (O_1187,N_20597,N_21296);
nand UO_1188 (O_1188,N_23120,N_23096);
nand UO_1189 (O_1189,N_18805,N_19078);
or UO_1190 (O_1190,N_24244,N_22190);
or UO_1191 (O_1191,N_20457,N_24960);
nor UO_1192 (O_1192,N_22881,N_19210);
nor UO_1193 (O_1193,N_18986,N_19935);
nor UO_1194 (O_1194,N_23586,N_24272);
nor UO_1195 (O_1195,N_23499,N_18786);
nor UO_1196 (O_1196,N_24332,N_24207);
or UO_1197 (O_1197,N_19112,N_24328);
nand UO_1198 (O_1198,N_19418,N_21484);
nand UO_1199 (O_1199,N_22687,N_21491);
nand UO_1200 (O_1200,N_19728,N_19678);
nand UO_1201 (O_1201,N_23584,N_18975);
nand UO_1202 (O_1202,N_19851,N_19228);
and UO_1203 (O_1203,N_18920,N_20130);
and UO_1204 (O_1204,N_24132,N_21575);
and UO_1205 (O_1205,N_24326,N_23402);
or UO_1206 (O_1206,N_19317,N_20594);
and UO_1207 (O_1207,N_20894,N_21056);
or UO_1208 (O_1208,N_21011,N_19082);
nand UO_1209 (O_1209,N_20680,N_21861);
nand UO_1210 (O_1210,N_23964,N_23963);
or UO_1211 (O_1211,N_23428,N_19383);
nand UO_1212 (O_1212,N_23094,N_20715);
nand UO_1213 (O_1213,N_20669,N_21130);
or UO_1214 (O_1214,N_23598,N_23741);
and UO_1215 (O_1215,N_24638,N_20147);
nand UO_1216 (O_1216,N_21217,N_24787);
and UO_1217 (O_1217,N_22811,N_20138);
or UO_1218 (O_1218,N_19288,N_24890);
xnor UO_1219 (O_1219,N_20610,N_21357);
and UO_1220 (O_1220,N_20155,N_24429);
or UO_1221 (O_1221,N_21230,N_24483);
and UO_1222 (O_1222,N_21944,N_19613);
nand UO_1223 (O_1223,N_19154,N_21158);
or UO_1224 (O_1224,N_24013,N_23659);
nand UO_1225 (O_1225,N_18852,N_20496);
xor UO_1226 (O_1226,N_20495,N_22283);
xnor UO_1227 (O_1227,N_21362,N_22916);
nor UO_1228 (O_1228,N_19054,N_22022);
and UO_1229 (O_1229,N_23502,N_19194);
nand UO_1230 (O_1230,N_22176,N_23748);
and UO_1231 (O_1231,N_21661,N_24198);
or UO_1232 (O_1232,N_19902,N_24128);
and UO_1233 (O_1233,N_20740,N_20067);
or UO_1234 (O_1234,N_19233,N_21299);
nor UO_1235 (O_1235,N_19395,N_20989);
and UO_1236 (O_1236,N_20693,N_24808);
nand UO_1237 (O_1237,N_22952,N_20695);
nor UO_1238 (O_1238,N_20835,N_24697);
or UO_1239 (O_1239,N_19750,N_24992);
nor UO_1240 (O_1240,N_22336,N_23343);
nor UO_1241 (O_1241,N_20412,N_21132);
or UO_1242 (O_1242,N_22789,N_21734);
and UO_1243 (O_1243,N_22133,N_24712);
or UO_1244 (O_1244,N_20501,N_22721);
or UO_1245 (O_1245,N_19858,N_24464);
nor UO_1246 (O_1246,N_22907,N_21030);
and UO_1247 (O_1247,N_20416,N_24180);
or UO_1248 (O_1248,N_19491,N_22943);
nor UO_1249 (O_1249,N_20015,N_18806);
nand UO_1250 (O_1250,N_24563,N_21989);
nand UO_1251 (O_1251,N_19438,N_21223);
and UO_1252 (O_1252,N_23810,N_19533);
and UO_1253 (O_1253,N_24803,N_19022);
or UO_1254 (O_1254,N_20536,N_19677);
or UO_1255 (O_1255,N_23758,N_21970);
nor UO_1256 (O_1256,N_21238,N_24407);
nand UO_1257 (O_1257,N_22641,N_19045);
nor UO_1258 (O_1258,N_21180,N_21346);
and UO_1259 (O_1259,N_21771,N_22914);
and UO_1260 (O_1260,N_23104,N_23039);
nor UO_1261 (O_1261,N_21640,N_24928);
nand UO_1262 (O_1262,N_24455,N_24720);
or UO_1263 (O_1263,N_21307,N_19574);
and UO_1264 (O_1264,N_21530,N_21233);
and UO_1265 (O_1265,N_22034,N_24486);
xnor UO_1266 (O_1266,N_19658,N_24817);
nand UO_1267 (O_1267,N_19642,N_24384);
and UO_1268 (O_1268,N_24804,N_24471);
xor UO_1269 (O_1269,N_21780,N_21138);
or UO_1270 (O_1270,N_23622,N_21352);
nor UO_1271 (O_1271,N_20291,N_22619);
and UO_1272 (O_1272,N_19067,N_20211);
and UO_1273 (O_1273,N_23708,N_23119);
nor UO_1274 (O_1274,N_20569,N_19878);
xor UO_1275 (O_1275,N_22808,N_20847);
nor UO_1276 (O_1276,N_20190,N_23756);
nor UO_1277 (O_1277,N_24823,N_24609);
and UO_1278 (O_1278,N_24038,N_23024);
and UO_1279 (O_1279,N_23523,N_23567);
nor UO_1280 (O_1280,N_23033,N_19798);
nand UO_1281 (O_1281,N_24630,N_22008);
nand UO_1282 (O_1282,N_22477,N_21439);
and UO_1283 (O_1283,N_24731,N_24868);
and UO_1284 (O_1284,N_20907,N_20605);
and UO_1285 (O_1285,N_23903,N_19072);
nand UO_1286 (O_1286,N_22001,N_20221);
nor UO_1287 (O_1287,N_18760,N_21555);
nand UO_1288 (O_1288,N_19332,N_22592);
or UO_1289 (O_1289,N_19236,N_23318);
nand UO_1290 (O_1290,N_19920,N_24673);
or UO_1291 (O_1291,N_18759,N_20828);
or UO_1292 (O_1292,N_21929,N_19249);
and UO_1293 (O_1293,N_22401,N_22908);
and UO_1294 (O_1294,N_19999,N_22949);
and UO_1295 (O_1295,N_22230,N_19685);
xnor UO_1296 (O_1296,N_21069,N_19320);
nor UO_1297 (O_1297,N_19061,N_22222);
and UO_1298 (O_1298,N_21333,N_23195);
nand UO_1299 (O_1299,N_22504,N_23935);
xor UO_1300 (O_1300,N_23127,N_21215);
nor UO_1301 (O_1301,N_22281,N_23735);
and UO_1302 (O_1302,N_22163,N_19303);
xor UO_1303 (O_1303,N_20428,N_23651);
xor UO_1304 (O_1304,N_23703,N_24049);
nand UO_1305 (O_1305,N_23949,N_23977);
or UO_1306 (O_1306,N_24258,N_18776);
and UO_1307 (O_1307,N_23609,N_21406);
or UO_1308 (O_1308,N_20178,N_21583);
or UO_1309 (O_1309,N_19571,N_21545);
nor UO_1310 (O_1310,N_20970,N_19496);
and UO_1311 (O_1311,N_22276,N_21822);
or UO_1312 (O_1312,N_20991,N_19250);
or UO_1313 (O_1313,N_22708,N_19654);
nand UO_1314 (O_1314,N_21385,N_22787);
and UO_1315 (O_1315,N_19578,N_20201);
and UO_1316 (O_1316,N_24514,N_21800);
nor UO_1317 (O_1317,N_22028,N_24876);
nor UO_1318 (O_1318,N_23854,N_20958);
or UO_1319 (O_1319,N_23896,N_21335);
or UO_1320 (O_1320,N_19230,N_22321);
nor UO_1321 (O_1321,N_24693,N_21921);
or UO_1322 (O_1322,N_19669,N_22998);
nand UO_1323 (O_1323,N_24266,N_20519);
or UO_1324 (O_1324,N_19141,N_18893);
nor UO_1325 (O_1325,N_21494,N_22899);
nand UO_1326 (O_1326,N_19030,N_24785);
or UO_1327 (O_1327,N_20801,N_19376);
nor UO_1328 (O_1328,N_24536,N_19350);
and UO_1329 (O_1329,N_21452,N_19327);
xnor UO_1330 (O_1330,N_23288,N_20462);
nand UO_1331 (O_1331,N_23013,N_23999);
nor UO_1332 (O_1332,N_19969,N_23219);
nand UO_1333 (O_1333,N_20559,N_24552);
or UO_1334 (O_1334,N_19657,N_20589);
nand UO_1335 (O_1335,N_24298,N_20606);
or UO_1336 (O_1336,N_23844,N_23049);
nor UO_1337 (O_1337,N_24757,N_22602);
and UO_1338 (O_1338,N_20653,N_19408);
nor UO_1339 (O_1339,N_19809,N_19692);
or UO_1340 (O_1340,N_23321,N_20550);
nand UO_1341 (O_1341,N_21316,N_24764);
or UO_1342 (O_1342,N_21403,N_20454);
nand UO_1343 (O_1343,N_23380,N_21862);
xor UO_1344 (O_1344,N_23650,N_19980);
nand UO_1345 (O_1345,N_21687,N_20297);
nand UO_1346 (O_1346,N_19339,N_22355);
nor UO_1347 (O_1347,N_19524,N_21300);
or UO_1348 (O_1348,N_23812,N_24977);
and UO_1349 (O_1349,N_19762,N_21819);
nor UO_1350 (O_1350,N_23270,N_21742);
or UO_1351 (O_1351,N_24210,N_20816);
nand UO_1352 (O_1352,N_23531,N_22871);
nand UO_1353 (O_1353,N_18950,N_23183);
nand UO_1354 (O_1354,N_22142,N_23565);
xnor UO_1355 (O_1355,N_22329,N_21285);
nor UO_1356 (O_1356,N_21176,N_19087);
nand UO_1357 (O_1357,N_21833,N_23895);
and UO_1358 (O_1358,N_20994,N_21381);
and UO_1359 (O_1359,N_21112,N_18795);
nand UO_1360 (O_1360,N_20629,N_22492);
and UO_1361 (O_1361,N_22876,N_21698);
nand UO_1362 (O_1362,N_20194,N_20121);
nand UO_1363 (O_1363,N_22748,N_22885);
and UO_1364 (O_1364,N_22954,N_20575);
or UO_1365 (O_1365,N_22529,N_21701);
nand UO_1366 (O_1366,N_21266,N_21407);
and UO_1367 (O_1367,N_20126,N_22121);
nand UO_1368 (O_1368,N_23447,N_24162);
or UO_1369 (O_1369,N_24724,N_20214);
or UO_1370 (O_1370,N_20508,N_23443);
and UO_1371 (O_1371,N_21395,N_24150);
or UO_1372 (O_1372,N_22946,N_21058);
nor UO_1373 (O_1373,N_24461,N_23240);
nand UO_1374 (O_1374,N_23676,N_20093);
or UO_1375 (O_1375,N_21303,N_23250);
or UO_1376 (O_1376,N_20925,N_23563);
and UO_1377 (O_1377,N_20103,N_24961);
nand UO_1378 (O_1378,N_21009,N_19046);
nand UO_1379 (O_1379,N_23037,N_19754);
xnor UO_1380 (O_1380,N_24428,N_21772);
nand UO_1381 (O_1381,N_23339,N_21536);
xnor UO_1382 (O_1382,N_21000,N_18919);
nor UO_1383 (O_1383,N_24427,N_22228);
and UO_1384 (O_1384,N_22715,N_23442);
or UO_1385 (O_1385,N_21292,N_23432);
and UO_1386 (O_1386,N_19011,N_22527);
or UO_1387 (O_1387,N_23777,N_22237);
or UO_1388 (O_1388,N_21642,N_22058);
nor UO_1389 (O_1389,N_20014,N_24220);
and UO_1390 (O_1390,N_21763,N_19753);
or UO_1391 (O_1391,N_24308,N_22833);
xor UO_1392 (O_1392,N_19189,N_21718);
or UO_1393 (O_1393,N_20808,N_22589);
xnor UO_1394 (O_1394,N_21549,N_20619);
nand UO_1395 (O_1395,N_24325,N_24294);
and UO_1396 (O_1396,N_24052,N_23920);
or UO_1397 (O_1397,N_21662,N_21941);
or UO_1398 (O_1398,N_24227,N_19176);
or UO_1399 (O_1399,N_22011,N_23746);
nor UO_1400 (O_1400,N_22734,N_21492);
nor UO_1401 (O_1401,N_19741,N_21946);
and UO_1402 (O_1402,N_22079,N_20687);
or UO_1403 (O_1403,N_20372,N_20802);
or UO_1404 (O_1404,N_24849,N_22797);
nand UO_1405 (O_1405,N_20471,N_20417);
and UO_1406 (O_1406,N_24595,N_20880);
nand UO_1407 (O_1407,N_21571,N_19984);
nand UO_1408 (O_1408,N_20885,N_20789);
and UO_1409 (O_1409,N_23618,N_19840);
and UO_1410 (O_1410,N_21284,N_21279);
xnor UO_1411 (O_1411,N_21987,N_24528);
xnor UO_1412 (O_1412,N_23495,N_22361);
and UO_1413 (O_1413,N_22587,N_19243);
and UO_1414 (O_1414,N_20879,N_22345);
xnor UO_1415 (O_1415,N_23818,N_21453);
nor UO_1416 (O_1416,N_20034,N_21913);
xor UO_1417 (O_1417,N_24158,N_23813);
nand UO_1418 (O_1418,N_22662,N_22235);
xnor UO_1419 (O_1419,N_24422,N_22398);
nand UO_1420 (O_1420,N_19756,N_19650);
nand UO_1421 (O_1421,N_19393,N_19596);
or UO_1422 (O_1422,N_19825,N_21447);
xnor UO_1423 (O_1423,N_23384,N_19834);
and UO_1424 (O_1424,N_22807,N_22359);
and UO_1425 (O_1425,N_21652,N_23427);
nand UO_1426 (O_1426,N_22672,N_21749);
or UO_1427 (O_1427,N_19456,N_24788);
and UO_1428 (O_1428,N_19345,N_23898);
and UO_1429 (O_1429,N_21421,N_23489);
nor UO_1430 (O_1430,N_21604,N_23216);
and UO_1431 (O_1431,N_23907,N_20691);
and UO_1432 (O_1432,N_18933,N_22277);
nor UO_1433 (O_1433,N_22537,N_21143);
nand UO_1434 (O_1434,N_22014,N_22567);
nor UO_1435 (O_1435,N_23667,N_21752);
or UO_1436 (O_1436,N_19370,N_21226);
nor UO_1437 (O_1437,N_23554,N_20851);
or UO_1438 (O_1438,N_24177,N_19586);
and UO_1439 (O_1439,N_24063,N_18843);
nor UO_1440 (O_1440,N_22225,N_20243);
nand UO_1441 (O_1441,N_24149,N_22571);
xor UO_1442 (O_1442,N_20565,N_23883);
or UO_1443 (O_1443,N_19856,N_23113);
nand UO_1444 (O_1444,N_21231,N_24670);
nand UO_1445 (O_1445,N_20404,N_19099);
nor UO_1446 (O_1446,N_21458,N_19396);
nor UO_1447 (O_1447,N_23161,N_21651);
nor UO_1448 (O_1448,N_23550,N_20204);
and UO_1449 (O_1449,N_20844,N_21274);
nor UO_1450 (O_1450,N_20019,N_23575);
nor UO_1451 (O_1451,N_21541,N_21122);
nand UO_1452 (O_1452,N_23107,N_23128);
nand UO_1453 (O_1453,N_21581,N_22825);
and UO_1454 (O_1454,N_20810,N_21547);
or UO_1455 (O_1455,N_23683,N_21924);
and UO_1456 (O_1456,N_24157,N_22704);
nor UO_1457 (O_1457,N_19180,N_24732);
nor UO_1458 (O_1458,N_20360,N_20834);
or UO_1459 (O_1459,N_20765,N_23894);
nor UO_1460 (O_1460,N_24979,N_22666);
or UO_1461 (O_1461,N_20241,N_21770);
nor UO_1462 (O_1462,N_20993,N_22410);
or UO_1463 (O_1463,N_20202,N_20498);
xor UO_1464 (O_1464,N_24530,N_23050);
and UO_1465 (O_1465,N_24116,N_23177);
and UO_1466 (O_1466,N_20311,N_22831);
and UO_1467 (O_1467,N_22706,N_22897);
nor UO_1468 (O_1468,N_23504,N_20570);
nor UO_1469 (O_1469,N_22274,N_22254);
and UO_1470 (O_1470,N_21816,N_22293);
and UO_1471 (O_1471,N_20110,N_21111);
nand UO_1472 (O_1472,N_22860,N_20057);
nor UO_1473 (O_1473,N_24984,N_24598);
xnor UO_1474 (O_1474,N_19815,N_19309);
nor UO_1475 (O_1475,N_24387,N_24072);
and UO_1476 (O_1476,N_19247,N_20156);
nor UO_1477 (O_1477,N_20699,N_21396);
xor UO_1478 (O_1478,N_21302,N_23411);
nor UO_1479 (O_1479,N_23220,N_19623);
and UO_1480 (O_1480,N_18772,N_23325);
or UO_1481 (O_1481,N_24185,N_22769);
and UO_1482 (O_1482,N_24100,N_20327);
xor UO_1483 (O_1483,N_20974,N_22310);
or UO_1484 (O_1484,N_22705,N_22689);
nand UO_1485 (O_1485,N_24113,N_22693);
and UO_1486 (O_1486,N_19463,N_22661);
nor UO_1487 (O_1487,N_20753,N_20729);
xor UO_1488 (O_1488,N_23845,N_19941);
nor UO_1489 (O_1489,N_20636,N_20787);
nand UO_1490 (O_1490,N_20547,N_23491);
xnor UO_1491 (O_1491,N_20934,N_19353);
and UO_1492 (O_1492,N_19922,N_21914);
nand UO_1493 (O_1493,N_22435,N_20356);
nor UO_1494 (O_1494,N_23353,N_20188);
or UO_1495 (O_1495,N_23494,N_21872);
nor UO_1496 (O_1496,N_22064,N_22339);
nor UO_1497 (O_1497,N_20875,N_18999);
nor UO_1498 (O_1498,N_24888,N_22647);
nor UO_1499 (O_1499,N_22248,N_22490);
or UO_1500 (O_1500,N_21410,N_20513);
or UO_1501 (O_1501,N_24330,N_20996);
nor UO_1502 (O_1502,N_20667,N_19883);
nor UO_1503 (O_1503,N_19227,N_22033);
nor UO_1504 (O_1504,N_21356,N_20161);
or UO_1505 (O_1505,N_20018,N_22685);
xor UO_1506 (O_1506,N_20757,N_18844);
and UO_1507 (O_1507,N_24657,N_24434);
nor UO_1508 (O_1508,N_20345,N_19382);
and UO_1509 (O_1509,N_24976,N_24473);
or UO_1510 (O_1510,N_19799,N_20321);
nor UO_1511 (O_1511,N_18832,N_23600);
nand UO_1512 (O_1512,N_22434,N_24708);
xnor UO_1513 (O_1513,N_19060,N_22875);
and UO_1514 (O_1514,N_23381,N_24962);
or UO_1515 (O_1515,N_23493,N_19483);
or UO_1516 (O_1516,N_20588,N_19114);
nand UO_1517 (O_1517,N_22713,N_23886);
or UO_1518 (O_1518,N_21374,N_21773);
nand UO_1519 (O_1519,N_20129,N_24027);
or UO_1520 (O_1520,N_19929,N_19940);
and UO_1521 (O_1521,N_19860,N_22189);
or UO_1522 (O_1522,N_24203,N_21186);
xor UO_1523 (O_1523,N_21695,N_19421);
or UO_1524 (O_1524,N_20254,N_23752);
nor UO_1525 (O_1525,N_24826,N_21539);
nand UO_1526 (O_1526,N_20173,N_24776);
nor UO_1527 (O_1527,N_19169,N_19712);
nor UO_1528 (O_1528,N_20758,N_20460);
nand UO_1529 (O_1529,N_19102,N_22627);
and UO_1530 (O_1530,N_18810,N_21606);
nor UO_1531 (O_1531,N_20061,N_21761);
nand UO_1532 (O_1532,N_22062,N_22813);
or UO_1533 (O_1533,N_22373,N_24497);
nand UO_1534 (O_1534,N_19319,N_22747);
nand UO_1535 (O_1535,N_23689,N_19513);
and UO_1536 (O_1536,N_22364,N_24123);
and UO_1537 (O_1537,N_19023,N_23415);
nor UO_1538 (O_1538,N_19621,N_22146);
and UO_1539 (O_1539,N_19667,N_22983);
or UO_1540 (O_1540,N_19826,N_23887);
and UO_1541 (O_1541,N_22031,N_21608);
and UO_1542 (O_1542,N_22535,N_24324);
and UO_1543 (O_1543,N_23892,N_24104);
xnor UO_1544 (O_1544,N_19276,N_22912);
nand UO_1545 (O_1545,N_23176,N_24212);
or UO_1546 (O_1546,N_19541,N_23221);
or UO_1547 (O_1547,N_19185,N_20637);
nand UO_1548 (O_1548,N_21144,N_23613);
nand UO_1549 (O_1549,N_21905,N_21724);
or UO_1550 (O_1550,N_20164,N_21927);
and UO_1551 (O_1551,N_22378,N_18889);
and UO_1552 (O_1552,N_20434,N_21320);
and UO_1553 (O_1553,N_24942,N_22915);
and UO_1554 (O_1554,N_19631,N_23303);
nand UO_1555 (O_1555,N_22509,N_19556);
or UO_1556 (O_1556,N_22698,N_21658);
nand UO_1557 (O_1557,N_19835,N_23125);
nor UO_1558 (O_1558,N_19111,N_24519);
or UO_1559 (O_1559,N_21590,N_23742);
xor UO_1560 (O_1560,N_24502,N_23378);
nor UO_1561 (O_1561,N_23787,N_19147);
nor UO_1562 (O_1562,N_24612,N_18996);
nand UO_1563 (O_1563,N_19917,N_19555);
or UO_1564 (O_1564,N_20995,N_24835);
nand UO_1565 (O_1565,N_19427,N_23202);
and UO_1566 (O_1566,N_19498,N_23589);
xnor UO_1567 (O_1567,N_23224,N_19229);
or UO_1568 (O_1568,N_22046,N_23142);
or UO_1569 (O_1569,N_23003,N_20763);
nor UO_1570 (O_1570,N_21993,N_23630);
nand UO_1571 (O_1571,N_20137,N_19108);
and UO_1572 (O_1572,N_21483,N_21354);
and UO_1573 (O_1573,N_22134,N_22131);
nand UO_1574 (O_1574,N_20215,N_20300);
nor UO_1575 (O_1575,N_20442,N_23004);
nand UO_1576 (O_1576,N_20698,N_20017);
nor UO_1577 (O_1577,N_19919,N_21309);
or UO_1578 (O_1578,N_21976,N_19566);
nand UO_1579 (O_1579,N_20977,N_19666);
nand UO_1580 (O_1580,N_24028,N_21558);
nor UO_1581 (O_1581,N_21440,N_18802);
xor UO_1582 (O_1582,N_19540,N_24396);
nor UO_1583 (O_1583,N_19744,N_19509);
xor UO_1584 (O_1584,N_24445,N_21760);
or UO_1585 (O_1585,N_19494,N_20659);
and UO_1586 (O_1586,N_19165,N_19736);
and UO_1587 (O_1587,N_23129,N_20341);
nand UO_1588 (O_1588,N_22354,N_20658);
and UO_1589 (O_1589,N_18954,N_22343);
or UO_1590 (O_1590,N_23362,N_21992);
nand UO_1591 (O_1591,N_22180,N_21165);
and UO_1592 (O_1592,N_23316,N_21971);
nor UO_1593 (O_1593,N_19116,N_24745);
nor UO_1594 (O_1594,N_24441,N_24226);
nand UO_1595 (O_1595,N_24264,N_23317);
or UO_1596 (O_1596,N_19458,N_21623);
or UO_1597 (O_1597,N_20979,N_24603);
and UO_1598 (O_1598,N_24115,N_19354);
and UO_1599 (O_1599,N_24183,N_20119);
nand UO_1600 (O_1600,N_20249,N_20154);
and UO_1601 (O_1601,N_22633,N_23835);
nand UO_1602 (O_1602,N_24354,N_22174);
xnor UO_1603 (O_1603,N_24892,N_21126);
nand UO_1604 (O_1604,N_23831,N_23633);
or UO_1605 (O_1605,N_21732,N_21181);
xnor UO_1606 (O_1606,N_19565,N_22617);
nor UO_1607 (O_1607,N_24243,N_22494);
nand UO_1608 (O_1608,N_22810,N_21854);
nand UO_1609 (O_1609,N_21846,N_19924);
xnor UO_1610 (O_1610,N_20089,N_24547);
nand UO_1611 (O_1611,N_20811,N_24652);
xnor UO_1612 (O_1612,N_23602,N_18779);
or UO_1613 (O_1613,N_23527,N_22138);
or UO_1614 (O_1614,N_18840,N_24056);
and UO_1615 (O_1615,N_20516,N_23888);
nand UO_1616 (O_1616,N_22473,N_21475);
nand UO_1617 (O_1617,N_21417,N_19523);
xor UO_1618 (O_1618,N_21617,N_19949);
or UO_1619 (O_1619,N_20084,N_21967);
nor UO_1620 (O_1620,N_19791,N_19976);
nor UO_1621 (O_1621,N_24959,N_19431);
or UO_1622 (O_1622,N_20140,N_22041);
and UO_1623 (O_1623,N_21127,N_19036);
xnor UO_1624 (O_1624,N_21409,N_24171);
or UO_1625 (O_1625,N_22930,N_24184);
nand UO_1626 (O_1626,N_20561,N_24813);
or UO_1627 (O_1627,N_24146,N_21005);
or UO_1628 (O_1628,N_18980,N_21544);
and UO_1629 (O_1629,N_22056,N_23863);
nand UO_1630 (O_1630,N_18968,N_21411);
or UO_1631 (O_1631,N_20579,N_24317);
and UO_1632 (O_1632,N_19075,N_22763);
and UO_1633 (O_1633,N_24286,N_24913);
and UO_1634 (O_1634,N_20444,N_24270);
or UO_1635 (O_1635,N_22753,N_20908);
nand UO_1636 (O_1636,N_22478,N_20265);
nor UO_1637 (O_1637,N_21328,N_24295);
nor UO_1638 (O_1638,N_19464,N_21940);
or UO_1639 (O_1639,N_22733,N_19050);
or UO_1640 (O_1640,N_24629,N_24492);
and UO_1641 (O_1641,N_21146,N_21568);
nor UO_1642 (O_1642,N_24139,N_21026);
nor UO_1643 (O_1643,N_22709,N_20307);
or UO_1644 (O_1644,N_21294,N_22933);
xor UO_1645 (O_1645,N_20305,N_20912);
nand UO_1646 (O_1646,N_21813,N_19268);
nor UO_1647 (O_1647,N_19056,N_22408);
nand UO_1648 (O_1648,N_19893,N_24261);
or UO_1649 (O_1649,N_22792,N_24501);
xor UO_1650 (O_1650,N_22764,N_21826);
or UO_1651 (O_1651,N_22386,N_19684);
nor UO_1652 (O_1652,N_20563,N_24309);
or UO_1653 (O_1653,N_24323,N_19557);
xor UO_1654 (O_1654,N_19755,N_23529);
or UO_1655 (O_1655,N_18926,N_20902);
nand UO_1656 (O_1656,N_22135,N_20716);
nand UO_1657 (O_1657,N_22668,N_18869);
xnor UO_1658 (O_1658,N_21079,N_21614);
xor UO_1659 (O_1659,N_20831,N_24069);
and UO_1660 (O_1660,N_21331,N_23720);
nand UO_1661 (O_1661,N_19177,N_19921);
nand UO_1662 (O_1662,N_22609,N_21665);
or UO_1663 (O_1663,N_21103,N_24364);
nand UO_1664 (O_1664,N_19572,N_21573);
or UO_1665 (O_1665,N_21653,N_21591);
nor UO_1666 (O_1666,N_24405,N_19970);
or UO_1667 (O_1667,N_19698,N_20793);
or UO_1668 (O_1668,N_24646,N_23144);
or UO_1669 (O_1669,N_20210,N_24241);
or UO_1670 (O_1670,N_19397,N_20055);
and UO_1671 (O_1671,N_24971,N_22749);
and UO_1672 (O_1672,N_22593,N_22741);
nand UO_1673 (O_1673,N_21154,N_20153);
xnor UO_1674 (O_1674,N_20220,N_23975);
and UO_1675 (O_1675,N_23986,N_20393);
and UO_1676 (O_1676,N_20545,N_22553);
or UO_1677 (O_1677,N_23425,N_18946);
nand UO_1678 (O_1678,N_23934,N_23249);
or UO_1679 (O_1679,N_21121,N_18943);
and UO_1680 (O_1680,N_24376,N_22973);
and UO_1681 (O_1681,N_20148,N_20768);
nand UO_1682 (O_1682,N_23404,N_23677);
or UO_1683 (O_1683,N_24588,N_22759);
nor UO_1684 (O_1684,N_24676,N_21688);
nor UO_1685 (O_1685,N_23580,N_19737);
and UO_1686 (O_1686,N_21716,N_19679);
or UO_1687 (O_1687,N_21647,N_19262);
and UO_1688 (O_1688,N_23770,N_19645);
or UO_1689 (O_1689,N_19696,N_21740);
or UO_1690 (O_1690,N_22938,N_23038);
xor UO_1691 (O_1691,N_20180,N_23417);
xnor UO_1692 (O_1692,N_19026,N_19582);
or UO_1693 (O_1693,N_24934,N_22481);
or UO_1694 (O_1694,N_21866,N_23564);
nor UO_1695 (O_1695,N_20081,N_23791);
or UO_1696 (O_1696,N_22980,N_19876);
and UO_1697 (O_1697,N_20279,N_20446);
or UO_1698 (O_1698,N_24568,N_22582);
or UO_1699 (O_1699,N_24229,N_19644);
and UO_1700 (O_1700,N_19583,N_19886);
nor UO_1701 (O_1701,N_23213,N_20861);
nor UO_1702 (O_1702,N_21559,N_24336);
or UO_1703 (O_1703,N_23166,N_19200);
and UO_1704 (O_1704,N_22895,N_20955);
and UO_1705 (O_1705,N_24283,N_22256);
and UO_1706 (O_1706,N_22460,N_20320);
or UO_1707 (O_1707,N_19942,N_21806);
nand UO_1708 (O_1708,N_20315,N_22496);
or UO_1709 (O_1709,N_21243,N_19710);
and UO_1710 (O_1710,N_24870,N_21503);
and UO_1711 (O_1711,N_19411,N_18909);
xor UO_1712 (O_1712,N_21920,N_22877);
and UO_1713 (O_1713,N_24448,N_23078);
xnor UO_1714 (O_1714,N_22697,N_19956);
xnor UO_1715 (O_1715,N_23552,N_21160);
and UO_1716 (O_1716,N_19625,N_21865);
nand UO_1717 (O_1717,N_23948,N_23263);
nand UO_1718 (O_1718,N_21474,N_19414);
and UO_1719 (O_1719,N_24155,N_24440);
and UO_1720 (O_1720,N_23700,N_19634);
nand UO_1721 (O_1721,N_19041,N_20873);
nand UO_1722 (O_1722,N_21690,N_24912);
nand UO_1723 (O_1723,N_20269,N_20150);
or UO_1724 (O_1724,N_21896,N_20397);
and UO_1725 (O_1725,N_21036,N_23591);
nand UO_1726 (O_1726,N_19832,N_23585);
or UO_1727 (O_1727,N_23872,N_23629);
nor UO_1728 (O_1728,N_21448,N_18787);
and UO_1729 (O_1729,N_21841,N_19149);
nor UO_1730 (O_1730,N_24919,N_19153);
nand UO_1731 (O_1731,N_22522,N_19966);
nor UO_1732 (O_1732,N_24199,N_20537);
or UO_1733 (O_1733,N_22947,N_20100);
nor UO_1734 (O_1734,N_23509,N_21712);
nor UO_1735 (O_1735,N_20077,N_18803);
or UO_1736 (O_1736,N_23925,N_24521);
or UO_1737 (O_1737,N_19990,N_24944);
nor UO_1738 (O_1738,N_21159,N_23675);
nand UO_1739 (O_1739,N_24704,N_21529);
nand UO_1740 (O_1740,N_18861,N_21102);
nor UO_1741 (O_1741,N_23215,N_21161);
or UO_1742 (O_1742,N_21745,N_20713);
xor UO_1743 (O_1743,N_20392,N_19453);
and UO_1744 (O_1744,N_21810,N_19977);
or UO_1745 (O_1745,N_18853,N_23853);
xnor UO_1746 (O_1746,N_24990,N_21017);
and UO_1747 (O_1747,N_24920,N_21229);
nand UO_1748 (O_1748,N_20120,N_20040);
or UO_1749 (O_1749,N_21134,N_20361);
nor UO_1750 (O_1750,N_21322,N_23725);
nor UO_1751 (O_1751,N_19615,N_19120);
or UO_1752 (O_1752,N_19436,N_20426);
nand UO_1753 (O_1753,N_21383,N_24752);
nor UO_1754 (O_1754,N_23168,N_19573);
or UO_1755 (O_1755,N_24777,N_20301);
nand UO_1756 (O_1756,N_21959,N_19057);
nand UO_1757 (O_1757,N_21202,N_23994);
xnor UO_1758 (O_1758,N_23825,N_21469);
or UO_1759 (O_1759,N_19896,N_19128);
xor UO_1760 (O_1760,N_23167,N_23631);
and UO_1761 (O_1761,N_23540,N_18860);
xor UO_1762 (O_1762,N_24895,N_24393);
nand UO_1763 (O_1763,N_20433,N_20386);
nand UO_1764 (O_1764,N_22624,N_20333);
and UO_1765 (O_1765,N_23921,N_21832);
nor UO_1766 (O_1766,N_21470,N_23273);
xnor UO_1767 (O_1767,N_19253,N_23020);
nand UO_1768 (O_1768,N_18780,N_22184);
nor UO_1769 (O_1769,N_22032,N_23640);
nand UO_1770 (O_1770,N_21991,N_23329);
xnor UO_1771 (O_1771,N_20239,N_21889);
nor UO_1772 (O_1772,N_22009,N_22913);
nor UO_1773 (O_1773,N_21106,N_20644);
and UO_1774 (O_1774,N_20704,N_20377);
or UO_1775 (O_1775,N_21928,N_20286);
xor UO_1776 (O_1776,N_19117,N_21599);
nand UO_1777 (O_1777,N_19048,N_22735);
or UO_1778 (O_1778,N_18955,N_21733);
xor UO_1779 (O_1779,N_19810,N_22441);
nor UO_1780 (O_1780,N_19290,N_22043);
or UO_1781 (O_1781,N_24090,N_24397);
and UO_1782 (O_1782,N_24940,N_19088);
nor UO_1783 (O_1783,N_21389,N_20634);
xor UO_1784 (O_1784,N_22772,N_23914);
and UO_1785 (O_1785,N_23829,N_20020);
nand UO_1786 (O_1786,N_22942,N_20807);
or UO_1787 (O_1787,N_24010,N_20096);
nand UO_1788 (O_1788,N_19240,N_20339);
and UO_1789 (O_1789,N_19814,N_23778);
or UO_1790 (O_1790,N_20567,N_23943);
nand UO_1791 (O_1791,N_18925,N_21910);
nor UO_1792 (O_1792,N_24674,N_18904);
nand UO_1793 (O_1793,N_24833,N_21954);
or UO_1794 (O_1794,N_24841,N_21107);
nor UO_1795 (O_1795,N_19468,N_24505);
nor UO_1796 (O_1796,N_19349,N_19328);
xnor UO_1797 (O_1797,N_21847,N_22436);
and UO_1798 (O_1798,N_23410,N_22240);
nor UO_1799 (O_1799,N_22736,N_21950);
nor UO_1800 (O_1800,N_23212,N_20244);
or UO_1801 (O_1801,N_24337,N_23162);
nand UO_1802 (O_1802,N_19610,N_21721);
nand UO_1803 (O_1803,N_22563,N_21490);
nand UO_1804 (O_1804,N_22517,N_21393);
nand UO_1805 (O_1805,N_20097,N_24715);
or UO_1806 (O_1806,N_22691,N_24988);
nand UO_1807 (O_1807,N_22444,N_24597);
nand UO_1808 (O_1808,N_20087,N_22569);
nor UO_1809 (O_1809,N_24449,N_22049);
nand UO_1810 (O_1810,N_19321,N_20845);
nor UO_1811 (O_1811,N_24614,N_22231);
or UO_1812 (O_1812,N_23775,N_20095);
nor UO_1813 (O_1813,N_19787,N_21864);
xnor UO_1814 (O_1814,N_19892,N_24133);
nor UO_1815 (O_1815,N_19542,N_19859);
and UO_1816 (O_1816,N_20663,N_24897);
or UO_1817 (O_1817,N_24290,N_21516);
or UO_1818 (O_1818,N_22804,N_24921);
or UO_1819 (O_1819,N_23062,N_20013);
or UO_1820 (O_1820,N_24621,N_23745);
nor UO_1821 (O_1821,N_21478,N_20646);
or UO_1822 (O_1822,N_19968,N_22433);
or UO_1823 (O_1823,N_24169,N_20749);
and UO_1824 (O_1824,N_18781,N_22549);
nand UO_1825 (O_1825,N_24400,N_22275);
or UO_1826 (O_1826,N_23721,N_24053);
or UO_1827 (O_1827,N_21936,N_19073);
nor UO_1828 (O_1828,N_22584,N_19487);
and UO_1829 (O_1829,N_23265,N_22775);
or UO_1830 (O_1830,N_21903,N_19344);
or UO_1831 (O_1831,N_20166,N_21224);
and UO_1832 (O_1832,N_22835,N_24533);
or UO_1833 (O_1833,N_21725,N_24691);
nand UO_1834 (O_1834,N_23172,N_24737);
or UO_1835 (O_1835,N_24273,N_21123);
xor UO_1836 (O_1836,N_22773,N_22894);
or UO_1837 (O_1837,N_22148,N_23679);
or UO_1838 (O_1838,N_22909,N_19587);
nor UO_1839 (O_1839,N_18756,N_18771);
nand UO_1840 (O_1840,N_19477,N_19238);
nand UO_1841 (O_1841,N_22063,N_22324);
nand UO_1842 (O_1842,N_20041,N_24366);
and UO_1843 (O_1843,N_21317,N_21019);
xor UO_1844 (O_1844,N_22768,N_19306);
xnor UO_1845 (O_1845,N_19937,N_24864);
or UO_1846 (O_1846,N_19521,N_24374);
xor UO_1847 (O_1847,N_21094,N_19964);
and UO_1848 (O_1848,N_20388,N_20971);
or UO_1849 (O_1849,N_20778,N_19518);
or UO_1850 (O_1850,N_22229,N_24883);
nor UO_1851 (O_1851,N_20914,N_23365);
xor UO_1852 (O_1852,N_22992,N_24305);
nand UO_1853 (O_1853,N_24466,N_19145);
or UO_1854 (O_1854,N_21336,N_21012);
nand UO_1855 (O_1855,N_22842,N_20049);
nor UO_1856 (O_1856,N_20047,N_21344);
nand UO_1857 (O_1857,N_19844,N_24872);
nor UO_1858 (O_1858,N_21696,N_20114);
or UO_1859 (O_1859,N_20612,N_21179);
or UO_1860 (O_1860,N_21435,N_20552);
xnor UO_1861 (O_1861,N_22505,N_20288);
nor UO_1862 (O_1862,N_22126,N_23574);
nand UO_1863 (O_1863,N_19245,N_24454);
nor UO_1864 (O_1864,N_21759,N_23132);
nor UO_1865 (O_1865,N_21379,N_24758);
nor UO_1866 (O_1866,N_21804,N_23302);
or UO_1867 (O_1867,N_21149,N_23579);
nor UO_1868 (O_1868,N_23739,N_24106);
and UO_1869 (O_1869,N_21714,N_24154);
or UO_1870 (O_1870,N_24558,N_24973);
nand UO_1871 (O_1871,N_21639,N_23467);
nand UO_1872 (O_1872,N_19124,N_22090);
or UO_1873 (O_1873,N_23971,N_19429);
nand UO_1874 (O_1874,N_23345,N_23275);
nor UO_1875 (O_1875,N_21029,N_24545);
nand UO_1876 (O_1876,N_20962,N_22199);
nor UO_1877 (O_1877,N_24275,N_20631);
nand UO_1878 (O_1878,N_23281,N_19870);
and UO_1879 (O_1879,N_23122,N_24399);
nor UO_1880 (O_1880,N_24224,N_19167);
or UO_1881 (O_1881,N_23487,N_22786);
or UO_1882 (O_1882,N_22036,N_24160);
or UO_1883 (O_1883,N_20284,N_20538);
or UO_1884 (O_1884,N_24917,N_23796);
nor UO_1885 (O_1885,N_24635,N_24512);
or UO_1886 (O_1886,N_21996,N_21035);
or UO_1887 (O_1887,N_22108,N_21837);
and UO_1888 (O_1888,N_21654,N_22251);
nand UO_1889 (O_1889,N_23989,N_18837);
nand UO_1890 (O_1890,N_20270,N_24459);
xor UO_1891 (O_1891,N_20455,N_22156);
or UO_1892 (O_1892,N_23276,N_19889);
nand UO_1893 (O_1893,N_23386,N_24042);
xor UO_1894 (O_1894,N_24193,N_24211);
or UO_1895 (O_1895,N_23422,N_21795);
and UO_1896 (O_1896,N_23065,N_20036);
and UO_1897 (O_1897,N_18915,N_24855);
nor UO_1898 (O_1898,N_24517,N_19495);
nand UO_1899 (O_1899,N_21717,N_24986);
nand UO_1900 (O_1900,N_18971,N_22956);
nand UO_1901 (O_1901,N_24291,N_19890);
and UO_1902 (O_1902,N_24779,N_20196);
nand UO_1903 (O_1903,N_23256,N_23452);
and UO_1904 (O_1904,N_19449,N_23044);
nand UO_1905 (O_1905,N_22044,N_20347);
or UO_1906 (O_1906,N_18858,N_18822);
or UO_1907 (O_1907,N_22308,N_19992);
or UO_1908 (O_1908,N_24191,N_21207);
nand UO_1909 (O_1909,N_24335,N_23701);
or UO_1910 (O_1910,N_23878,N_22784);
nand UO_1911 (O_1911,N_24666,N_24377);
or UO_1912 (O_1912,N_22757,N_20849);
nand UO_1913 (O_1913,N_21550,N_19913);
nor UO_1914 (O_1914,N_18814,N_19504);
nor UO_1915 (O_1915,N_19366,N_21250);
and UO_1916 (O_1916,N_19749,N_22632);
or UO_1917 (O_1917,N_21338,N_22302);
and UO_1918 (O_1918,N_21678,N_23268);
xor UO_1919 (O_1919,N_22669,N_23420);
and UO_1920 (O_1920,N_23959,N_22385);
xor UO_1921 (O_1921,N_22520,N_19305);
and UO_1922 (O_1922,N_18859,N_20354);
nand UO_1923 (O_1923,N_19721,N_23466);
nand UO_1924 (O_1924,N_21031,N_18849);
and UO_1925 (O_1925,N_23512,N_22381);
or UO_1926 (O_1926,N_19323,N_24031);
nand UO_1927 (O_1927,N_22026,N_19746);
or UO_1928 (O_1928,N_22155,N_21188);
nand UO_1929 (O_1929,N_21416,N_24457);
and UO_1930 (O_1930,N_19715,N_21968);
and UO_1931 (O_1931,N_24997,N_24885);
nor UO_1932 (O_1932,N_24617,N_20542);
nand UO_1933 (O_1933,N_20770,N_21363);
nor UO_1934 (O_1934,N_22193,N_23553);
and UO_1935 (O_1935,N_21136,N_24963);
nor UO_1936 (O_1936,N_22837,N_24664);
nand UO_1937 (O_1937,N_22384,N_23747);
nand UO_1938 (O_1938,N_23603,N_21151);
nand UO_1939 (O_1939,N_19018,N_24439);
nor UO_1940 (O_1940,N_24026,N_19394);
and UO_1941 (O_1941,N_24825,N_24710);
or UO_1942 (O_1942,N_19006,N_24424);
and UO_1943 (O_1943,N_20193,N_20142);
and UO_1944 (O_1944,N_18769,N_24006);
nand UO_1945 (O_1945,N_21249,N_20420);
nor UO_1946 (O_1946,N_21916,N_22556);
nand UO_1947 (O_1947,N_23987,N_19110);
or UO_1948 (O_1948,N_19805,N_22551);
and UO_1949 (O_1949,N_22651,N_22761);
nor UO_1950 (O_1950,N_21566,N_22910);
and UO_1951 (O_1951,N_24209,N_21342);
nand UO_1952 (O_1952,N_24228,N_23481);
and UO_1953 (O_1953,N_24386,N_19209);
xnor UO_1954 (O_1954,N_22544,N_21020);
nor UO_1955 (O_1955,N_20400,N_21289);
or UO_1956 (O_1956,N_20572,N_24164);
nand UO_1957 (O_1957,N_19066,N_19140);
and UO_1958 (O_1958,N_23674,N_23355);
and UO_1959 (O_1959,N_20702,N_23926);
and UO_1960 (O_1960,N_19137,N_23566);
and UO_1961 (O_1961,N_23882,N_21254);
nand UO_1962 (O_1962,N_23308,N_19118);
or UO_1963 (O_1963,N_24284,N_23663);
nor UO_1964 (O_1964,N_19042,N_20751);
nand UO_1965 (O_1965,N_23109,N_24980);
and UO_1966 (O_1966,N_24269,N_24839);
or UO_1967 (O_1967,N_24755,N_19359);
nor UO_1968 (O_1968,N_23982,N_23348);
nor UO_1969 (O_1969,N_22298,N_22094);
or UO_1970 (O_1970,N_21182,N_24385);
xor UO_1971 (O_1971,N_20825,N_19085);
nor UO_1972 (O_1972,N_21632,N_24750);
nor UO_1973 (O_1973,N_20832,N_24012);
nor UO_1974 (O_1974,N_21955,N_20452);
and UO_1975 (O_1975,N_24681,N_19670);
nor UO_1976 (O_1976,N_22206,N_20843);
or UO_1977 (O_1977,N_24469,N_21748);
nand UO_1978 (O_1978,N_19580,N_23548);
or UO_1979 (O_1979,N_22655,N_20272);
and UO_1980 (O_1980,N_18961,N_19918);
nor UO_1981 (O_1981,N_24419,N_22547);
nand UO_1982 (O_1982,N_20625,N_24363);
or UO_1983 (O_1983,N_20440,N_21709);
nand UO_1984 (O_1984,N_24707,N_21205);
xnor UO_1985 (O_1985,N_20773,N_23751);
nand UO_1986 (O_1986,N_23360,N_24520);
nand UO_1987 (O_1987,N_24954,N_21450);
and UO_1988 (O_1988,N_22904,N_21728);
and UO_1989 (O_1989,N_18945,N_19092);
nor UO_1990 (O_1990,N_22648,N_20923);
nand UO_1991 (O_1991,N_22412,N_23097);
nand UO_1992 (O_1992,N_24816,N_23450);
nor UO_1993 (O_1993,N_24493,N_24838);
nand UO_1994 (O_1994,N_21025,N_20409);
nand UO_1995 (O_1995,N_18882,N_22959);
nand UO_1996 (O_1996,N_24734,N_19334);
nand UO_1997 (O_1997,N_21098,N_19346);
nand UO_1998 (O_1998,N_22867,N_23995);
nor UO_1999 (O_1999,N_22851,N_19059);
nand UO_2000 (O_2000,N_19735,N_22570);
and UO_2001 (O_2001,N_21876,N_21183);
and UO_2002 (O_2002,N_19939,N_24343);
nor UO_2003 (O_2003,N_23953,N_19777);
and UO_2004 (O_2004,N_23300,N_21580);
and UO_2005 (O_2005,N_19000,N_21978);
xnor UO_2006 (O_2006,N_23283,N_19713);
or UO_2007 (O_2007,N_22296,N_21649);
and UO_2008 (O_2008,N_24721,N_23828);
or UO_2009 (O_2009,N_19475,N_21595);
nand UO_2010 (O_2010,N_20850,N_18847);
xor UO_2011 (O_2011,N_18754,N_21257);
nor UO_2012 (O_2012,N_18821,N_23018);
or UO_2013 (O_2013,N_22616,N_21935);
nor UO_2014 (O_2014,N_23843,N_22650);
and UO_2015 (O_2015,N_22929,N_22793);
and UO_2016 (O_2016,N_20518,N_22246);
nand UO_2017 (O_2017,N_23383,N_21579);
nor UO_2018 (O_2018,N_22836,N_23083);
or UO_2019 (O_2019,N_20642,N_22319);
xor UO_2020 (O_2020,N_19656,N_19551);
xor UO_2021 (O_2021,N_24542,N_20660);
nand UO_2022 (O_2022,N_20870,N_20186);
and UO_2023 (O_2023,N_22712,N_22683);
or UO_2024 (O_2024,N_21219,N_22351);
or UO_2025 (O_2025,N_24235,N_21391);
nor UO_2026 (O_2026,N_23911,N_24019);
xnor UO_2027 (O_2027,N_19287,N_23556);
xor UO_2028 (O_2028,N_23784,N_22482);
xnor UO_2029 (O_2029,N_21807,N_21677);
nor UO_2030 (O_2030,N_22720,N_21489);
or UO_2031 (O_2031,N_24002,N_24268);
and UO_2032 (O_2032,N_24987,N_23403);
or UO_2033 (O_2033,N_19946,N_24192);
xnor UO_2034 (O_2034,N_22752,N_22828);
nand UO_2035 (O_2035,N_19192,N_19998);
nand UO_2036 (O_2036,N_20125,N_24768);
or UO_2037 (O_2037,N_23587,N_19314);
nand UO_2038 (O_2038,N_21166,N_21301);
nor UO_2039 (O_2039,N_22096,N_21288);
nor UO_2040 (O_2040,N_24820,N_24736);
nand UO_2041 (O_2041,N_19930,N_19704);
and UO_2042 (O_2042,N_21236,N_24453);
nor UO_2043 (O_2043,N_20821,N_19532);
nor UO_2044 (O_2044,N_21930,N_20761);
nor UO_2045 (O_2045,N_23521,N_20324);
and UO_2046 (O_2046,N_21633,N_20035);
xnor UO_2047 (O_2047,N_22671,N_22511);
and UO_2048 (O_2048,N_19095,N_19398);
nor UO_2049 (O_2049,N_18789,N_24525);
xor UO_2050 (O_2050,N_19360,N_19662);
xnor UO_2051 (O_2051,N_24465,N_24395);
nor UO_2052 (O_2052,N_24313,N_19751);
or UO_2053 (O_2053,N_20058,N_18801);
xor UO_2054 (O_2054,N_21723,N_24242);
or UO_2055 (O_2055,N_21894,N_20117);
and UO_2056 (O_2056,N_20246,N_22322);
nand UO_2057 (O_2057,N_22143,N_18880);
nor UO_2058 (O_2058,N_22832,N_19358);
or UO_2059 (O_2059,N_20818,N_21119);
xor UO_2060 (O_2060,N_23012,N_22886);
nand UO_2061 (O_2061,N_19256,N_23075);
or UO_2062 (O_2062,N_24021,N_21259);
nor UO_2063 (O_2063,N_19170,N_19378);
nor UO_2064 (O_2064,N_23160,N_21574);
nand UO_2065 (O_2065,N_24829,N_21482);
nand UO_2066 (O_2066,N_19776,N_21915);
nor UO_2067 (O_2067,N_22367,N_23737);
nand UO_2068 (O_2068,N_22984,N_20676);
nor UO_2069 (O_2069,N_21908,N_19150);
or UO_2070 (O_2070,N_22285,N_23217);
and UO_2071 (O_2071,N_22498,N_19419);
and UO_2072 (O_2072,N_23102,N_19131);
xor UO_2073 (O_2073,N_19972,N_20008);
nand UO_2074 (O_2074,N_23962,N_24911);
nor UO_2075 (O_2075,N_20363,N_22488);
or UO_2076 (O_2076,N_24989,N_24559);
and UO_2077 (O_2077,N_23545,N_21540);
nor UO_2078 (O_2078,N_20868,N_20898);
nand UO_2079 (O_2079,N_24375,N_19390);
or UO_2080 (O_2080,N_23794,N_20511);
and UO_2081 (O_2081,N_24957,N_23101);
nor UO_2082 (O_2082,N_24379,N_22328);
nand UO_2083 (O_2083,N_20969,N_19286);
and UO_2084 (O_2084,N_21329,N_24446);
or UO_2085 (O_2085,N_24078,N_21084);
nor UO_2086 (O_2086,N_19781,N_23138);
or UO_2087 (O_2087,N_23714,N_24430);
nor UO_2088 (O_2088,N_19472,N_19159);
nor UO_2089 (O_2089,N_21613,N_24420);
nand UO_2090 (O_2090,N_23416,N_18947);
or UO_2091 (O_2091,N_19818,N_19761);
nand UO_2092 (O_2092,N_24601,N_23996);
nand UO_2093 (O_2093,N_20837,N_20158);
and UO_2094 (O_2094,N_20070,N_19747);
and UO_2095 (O_2095,N_23805,N_19326);
and UO_2096 (O_2096,N_22659,N_21287);
nor UO_2097 (O_2097,N_21686,N_23073);
nand UO_2098 (O_2098,N_23089,N_20515);
nor UO_2099 (O_2099,N_19152,N_20387);
nand UO_2100 (O_2100,N_19595,N_23203);
or UO_2101 (O_2101,N_19302,N_22665);
nor UO_2102 (O_2102,N_18836,N_22981);
nor UO_2103 (O_2103,N_20604,N_24288);
or UO_2104 (O_2104,N_23841,N_23023);
and UO_2105 (O_2105,N_20234,N_22416);
nand UO_2106 (O_2106,N_18833,N_24865);
or UO_2107 (O_2107,N_20746,N_20564);
and UO_2108 (O_2108,N_22499,N_24248);
nand UO_2109 (O_2109,N_24930,N_24382);
or UO_2110 (O_2110,N_21218,N_23246);
nor UO_2111 (O_2111,N_21085,N_23573);
nor UO_2112 (O_2112,N_22166,N_23990);
or UO_2113 (O_2113,N_20799,N_24442);
or UO_2114 (O_2114,N_19600,N_19318);
or UO_2115 (O_2115,N_23260,N_19214);
nor UO_2116 (O_2116,N_24201,N_19489);
nand UO_2117 (O_2117,N_23482,N_21693);
xnor UO_2118 (O_2118,N_22347,N_19797);
nor UO_2119 (O_2119,N_23439,N_22314);
and UO_2120 (O_2120,N_24950,N_22588);
nand UO_2121 (O_2121,N_19944,N_24498);
or UO_2122 (O_2122,N_24580,N_18903);
and UO_2123 (O_2123,N_24345,N_23846);
nor UO_2124 (O_2124,N_18965,N_24908);
nand UO_2125 (O_2125,N_23806,N_19164);
and UO_2126 (O_2126,N_23765,N_21509);
nand UO_2127 (O_2127,N_23305,N_21446);
or UO_2128 (O_2128,N_20862,N_24799);
nor UO_2129 (O_2129,N_20904,N_22470);
or UO_2130 (O_2130,N_20614,N_23459);
xnor UO_2131 (O_2131,N_19500,N_22990);
nand UO_2132 (O_2132,N_22109,N_22365);
or UO_2133 (O_2133,N_22686,N_20146);
nand UO_2134 (O_2134,N_24690,N_22326);
nand UO_2135 (O_2135,N_22383,N_22104);
nand UO_2136 (O_2136,N_19297,N_20443);
nor UO_2137 (O_2137,N_20957,N_19205);
and UO_2138 (O_2138,N_22575,N_23879);
xor UO_2139 (O_2139,N_20945,N_19965);
or UO_2140 (O_2140,N_24122,N_21214);
or UO_2141 (O_2141,N_21369,N_22642);
and UO_2142 (O_2142,N_21797,N_23226);
nor UO_2143 (O_2143,N_23668,N_19035);
nand UO_2144 (O_2144,N_20722,N_21900);
nor UO_2145 (O_2145,N_21185,N_24564);
nor UO_2146 (O_2146,N_21096,N_23230);
and UO_2147 (O_2147,N_21486,N_18898);
and UO_2148 (O_2148,N_24902,N_18808);
xnor UO_2149 (O_2149,N_20229,N_22092);
or UO_2150 (O_2150,N_24735,N_22805);
nand UO_2151 (O_2151,N_22779,N_19450);
or UO_2152 (O_2152,N_22611,N_22843);
and UO_2153 (O_2153,N_23311,N_20797);
and UO_2154 (O_2154,N_22208,N_19481);
and UO_2155 (O_2155,N_23082,N_21958);
and UO_2156 (O_2156,N_19336,N_24451);
nor UO_2157 (O_2157,N_19204,N_22111);
and UO_2158 (O_2158,N_20343,N_23954);
or UO_2159 (O_2159,N_20886,N_21977);
and UO_2160 (O_2160,N_20911,N_19983);
nand UO_2161 (O_2161,N_20497,N_23057);
nand UO_2162 (O_2162,N_24863,N_24537);
nor UO_2163 (O_2163,N_22250,N_19364);
and UO_2164 (O_2164,N_19512,N_20414);
or UO_2165 (O_2165,N_22985,N_21220);
or UO_2166 (O_2166,N_22920,N_23361);
and UO_2167 (O_2167,N_19906,N_24039);
nand UO_2168 (O_2168,N_19911,N_22839);
nand UO_2169 (O_2169,N_21682,N_20790);
and UO_2170 (O_2170,N_23562,N_22305);
nand UO_2171 (O_2171,N_24975,N_19417);
nor UO_2172 (O_2172,N_19873,N_24915);
or UO_2173 (O_2173,N_21057,N_20781);
nand UO_2174 (O_2174,N_24361,N_19986);
and UO_2175 (O_2175,N_22710,N_22991);
and UO_2176 (O_2176,N_23254,N_21974);
or UO_2177 (O_2177,N_24134,N_22858);
and UO_2178 (O_2178,N_21091,N_22585);
or UO_2179 (O_2179,N_24922,N_20398);
nand UO_2180 (O_2180,N_20611,N_21037);
nor UO_2181 (O_2181,N_22979,N_19868);
nand UO_2182 (O_2182,N_21293,N_19093);
and UO_2183 (O_2183,N_20546,N_23026);
nor UO_2184 (O_2184,N_24277,N_22756);
nor UO_2185 (O_2185,N_21232,N_19738);
nand UO_2186 (O_2186,N_20195,N_24604);
nor UO_2187 (O_2187,N_24927,N_24077);
xnor UO_2188 (O_2188,N_22961,N_21669);
nand UO_2189 (O_2189,N_21459,N_22703);
or UO_2190 (O_2190,N_21753,N_24001);
nand UO_2191 (O_2191,N_22847,N_23815);
and UO_2192 (O_2192,N_19638,N_19831);
or UO_2193 (O_2193,N_20877,N_24508);
xor UO_2194 (O_2194,N_19985,N_20056);
nor UO_2195 (O_2195,N_23040,N_23840);
nand UO_2196 (O_2196,N_18862,N_20402);
and UO_2197 (O_2197,N_20953,N_22799);
nor UO_2198 (O_2198,N_24254,N_24425);
nand UO_2199 (O_2199,N_24504,N_19647);
xor UO_2200 (O_2200,N_21517,N_23352);
and UO_2201 (O_2201,N_22724,N_22469);
or UO_2202 (O_2202,N_23084,N_22782);
nor UO_2203 (O_2203,N_20673,N_22202);
and UO_2204 (O_2204,N_19220,N_21349);
nand UO_2205 (O_2205,N_23146,N_24847);
and UO_2206 (O_2206,N_24526,N_24096);
and UO_2207 (O_2207,N_21675,N_22963);
nand UO_2208 (O_2208,N_24842,N_22923);
nor UO_2209 (O_2209,N_24099,N_20901);
and UO_2210 (O_2210,N_24587,N_23838);
nand UO_2211 (O_2211,N_21792,N_22936);
nand UO_2212 (O_2212,N_22902,N_21353);
nand UO_2213 (O_2213,N_21221,N_21377);
nand UO_2214 (O_2214,N_21655,N_20780);
nand UO_2215 (O_2215,N_19987,N_20366);
nand UO_2216 (O_2216,N_21619,N_22151);
and UO_2217 (O_2217,N_24793,N_19207);
or UO_2218 (O_2218,N_20846,N_19181);
nand UO_2219 (O_2219,N_23972,N_21812);
or UO_2220 (O_2220,N_20984,N_23478);
nor UO_2221 (O_2221,N_21169,N_24845);
nor UO_2222 (O_2222,N_20352,N_24789);
nand UO_2223 (O_2223,N_20679,N_23785);
nand UO_2224 (O_2224,N_20218,N_23625);
nor UO_2225 (O_2225,N_21460,N_23398);
xnor UO_2226 (O_2226,N_23471,N_18798);
nor UO_2227 (O_2227,N_23519,N_18932);
or UO_2228 (O_2228,N_19774,N_24669);
or UO_2229 (O_2229,N_23969,N_21431);
nor UO_2230 (O_2230,N_20411,N_22639);
xor UO_2231 (O_2231,N_20742,N_23992);
xnor UO_2232 (O_2232,N_23111,N_23358);
nand UO_2233 (O_2233,N_23626,N_21462);
xor UO_2234 (O_2234,N_23169,N_24417);
nor UO_2235 (O_2235,N_24478,N_21899);
and UO_2236 (O_2236,N_23423,N_20990);
nand UO_2237 (O_2237,N_21793,N_19530);
or UO_2238 (O_2238,N_22673,N_20921);
and UO_2239 (O_2239,N_19040,N_20860);
and UO_2240 (O_2240,N_19786,N_23448);
nor UO_2241 (O_2241,N_24631,N_20672);
nand UO_2242 (O_2242,N_22407,N_20730);
or UO_2243 (O_2243,N_22244,N_23532);
nand UO_2244 (O_2244,N_21024,N_21034);
and UO_2245 (O_2245,N_20635,N_23247);
nand UO_2246 (O_2246,N_24810,N_23354);
nand UO_2247 (O_2247,N_24557,N_23342);
nor UO_2248 (O_2248,N_20755,N_21171);
or UO_2249 (O_2249,N_23333,N_18750);
nand UO_2250 (O_2250,N_21710,N_19254);
nor UO_2251 (O_2251,N_23196,N_18922);
and UO_2252 (O_2252,N_22242,N_23923);
nor UO_2253 (O_2253,N_21082,N_23867);
and UO_2254 (O_2254,N_21187,N_22906);
nor UO_2255 (O_2255,N_19443,N_22100);
nor UO_2256 (O_2256,N_24932,N_23684);
or UO_2257 (O_2257,N_18907,N_18778);
xor UO_2258 (O_2258,N_24089,N_22849);
nor UO_2259 (O_2259,N_20759,N_22366);
nor UO_2260 (O_2260,N_19051,N_22657);
nor UO_2261 (O_2261,N_23066,N_23873);
and UO_2262 (O_2262,N_19543,N_19743);
nor UO_2263 (O_2263,N_21932,N_24035);
nand UO_2264 (O_2264,N_19763,N_23081);
and UO_2265 (O_2265,N_23406,N_22306);
nand UO_2266 (O_2266,N_19299,N_20262);
nand UO_2267 (O_2267,N_23998,N_22387);
or UO_2268 (O_2268,N_20351,N_22884);
and UO_2269 (O_2269,N_22172,N_21488);
xor UO_2270 (O_2270,N_22795,N_20624);
and UO_2271 (O_2271,N_19391,N_19480);
or UO_2272 (O_2272,N_24148,N_23407);
nor UO_2273 (O_2273,N_23717,N_23874);
or UO_2274 (O_2274,N_19400,N_22791);
or UO_2275 (O_2275,N_23814,N_18998);
xnor UO_2276 (O_2276,N_20670,N_19232);
or UO_2277 (O_2277,N_24656,N_24766);
and UO_2278 (O_2278,N_23261,N_19097);
nor UO_2279 (O_2279,N_24306,N_23400);
and UO_2280 (O_2280,N_23010,N_18871);
or UO_2281 (O_2281,N_19959,N_20287);
nand UO_2282 (O_2282,N_23792,N_20099);
and UO_2283 (O_2283,N_19759,N_24341);
xnor UO_2284 (O_2284,N_22714,N_19275);
nor UO_2285 (O_2285,N_19015,N_23929);
nor UO_2286 (O_2286,N_18970,N_20413);
nor UO_2287 (O_2287,N_21960,N_21485);
or UO_2288 (O_2288,N_22114,N_24553);
nor UO_2289 (O_2289,N_23595,N_19130);
and UO_2290 (O_2290,N_24686,N_24532);
or UO_2291 (O_2291,N_23740,N_21607);
and UO_2292 (O_2292,N_23772,N_20259);
or UO_2293 (O_2293,N_20950,N_20038);
nand UO_2294 (O_2294,N_19620,N_24762);
and UO_2295 (O_2295,N_24219,N_18989);
or UO_2296 (O_2296,N_24901,N_19909);
and UO_2297 (O_2297,N_23528,N_23577);
nand UO_2298 (O_2298,N_21177,N_24862);
nor UO_2299 (O_2299,N_22426,N_24074);
nand UO_2300 (O_2300,N_20076,N_24015);
nand UO_2301 (O_2301,N_22644,N_19899);
xor UO_2302 (O_2302,N_22968,N_23016);
or UO_2303 (O_2303,N_18894,N_24649);
and UO_2304 (O_2304,N_23762,N_20235);
nor UO_2305 (O_2305,N_21857,N_21351);
nand UO_2306 (O_2306,N_20338,N_20541);
xnor UO_2307 (O_2307,N_19768,N_20346);
or UO_2308 (O_2308,N_22766,N_20668);
xor UO_2309 (O_2309,N_18886,N_19594);
xor UO_2310 (O_2310,N_19660,N_22149);
xor UO_2311 (O_2311,N_22074,N_19932);
and UO_2312 (O_2312,N_22722,N_23869);
and UO_2313 (O_2313,N_24265,N_20500);
nor UO_2314 (O_2314,N_24815,N_22261);
nor UO_2315 (O_2315,N_18765,N_23681);
nor UO_2316 (O_2316,N_23985,N_20917);
nor UO_2317 (O_2317,N_19802,N_22003);
and UO_2318 (O_2318,N_19579,N_23979);
nor UO_2319 (O_2319,N_21413,N_24696);
nor UO_2320 (O_2320,N_23369,N_20591);
or UO_2321 (O_2321,N_20112,N_21957);
nor UO_2322 (O_2322,N_20085,N_23464);
xor UO_2323 (O_2323,N_23367,N_20964);
nand UO_2324 (O_2324,N_19448,N_22266);
or UO_2325 (O_2325,N_20639,N_24939);
and UO_2326 (O_2326,N_21827,N_22892);
xnor UO_2327 (O_2327,N_20616,N_20812);
or UO_2328 (O_2328,N_23006,N_23117);
nor UO_2329 (O_2329,N_20980,N_20059);
and UO_2330 (O_2330,N_22015,N_23359);
or UO_2331 (O_2331,N_19544,N_22820);
nand UO_2332 (O_2332,N_24263,N_19020);
or UO_2333 (O_2333,N_20592,N_20131);
nand UO_2334 (O_2334,N_24047,N_21624);
nand UO_2335 (O_2335,N_21859,N_24958);
and UO_2336 (O_2336,N_22173,N_22129);
or UO_2337 (O_2337,N_24578,N_20199);
nand UO_2338 (O_2338,N_21739,N_20079);
and UO_2339 (O_2339,N_19539,N_19195);
nand UO_2340 (O_2340,N_20348,N_22862);
or UO_2341 (O_2341,N_22935,N_19916);
or UO_2342 (O_2342,N_22466,N_20482);
or UO_2343 (O_2343,N_24790,N_19525);
and UO_2344 (O_2344,N_23488,N_20527);
or UO_2345 (O_2345,N_20792,N_23688);
or UO_2346 (O_2346,N_22004,N_20804);
and UO_2347 (O_2347,N_24000,N_19485);
nor UO_2348 (O_2348,N_23615,N_24570);
and UO_2349 (O_2349,N_22452,N_23705);
nand UO_2350 (O_2350,N_20956,N_21414);
or UO_2351 (O_2351,N_22767,N_23652);
and UO_2352 (O_2352,N_21348,N_21569);
and UO_2353 (O_2353,N_19683,N_20734);
nand UO_2354 (O_2354,N_19259,N_19568);
and UO_2355 (O_2355,N_21170,N_22566);
or UO_2356 (O_2356,N_24660,N_23266);
nand UO_2357 (O_2357,N_24156,N_24344);
nand UO_2358 (O_2358,N_21228,N_21582);
nand UO_2359 (O_2359,N_19062,N_19342);
xnor UO_2360 (O_2360,N_21247,N_24356);
nor UO_2361 (O_2361,N_23930,N_24225);
nand UO_2362 (O_2362,N_21051,N_23771);
nand UO_2363 (O_2363,N_23793,N_19813);
and UO_2364 (O_2364,N_19716,N_21099);
or UO_2365 (O_2365,N_20395,N_21605);
nand UO_2366 (O_2366,N_23811,N_20107);
or UO_2367 (O_2367,N_22284,N_23150);
or UO_2368 (O_2368,N_24549,N_24406);
nand UO_2369 (O_2369,N_22399,N_22213);
and UO_2370 (O_2370,N_24362,N_23593);
or UO_2371 (O_2371,N_22838,N_19410);
nor UO_2372 (O_2372,N_21310,N_21934);
nand UO_2373 (O_2373,N_22349,N_23298);
nand UO_2374 (O_2374,N_22716,N_21883);
nand UO_2375 (O_2375,N_23660,N_24882);
xor UO_2376 (O_2376,N_20784,N_24278);
or UO_2377 (O_2377,N_21738,N_19218);
nor UO_2378 (O_2378,N_19691,N_23816);
or UO_2379 (O_2379,N_20257,N_20817);
or UO_2380 (O_2380,N_20007,N_23709);
nor UO_2381 (O_2381,N_20578,N_20936);
and UO_2382 (O_2382,N_20358,N_23000);
or UO_2383 (O_2383,N_20448,N_23876);
and UO_2384 (O_2384,N_22599,N_22084);
nand UO_2385 (O_2385,N_18834,N_20072);
and UO_2386 (O_2386,N_21691,N_22075);
nor UO_2387 (O_2387,N_19812,N_23114);
nor UO_2388 (O_2388,N_23123,N_23189);
or UO_2389 (O_2389,N_21326,N_21788);
or UO_2390 (O_2390,N_22428,N_24011);
and UO_2391 (O_2391,N_20441,N_22217);
nor UO_2392 (O_2392,N_20874,N_21350);
nand UO_2393 (O_2393,N_24886,N_22024);
and UO_2394 (O_2394,N_23421,N_24916);
or UO_2395 (O_2395,N_19622,N_22082);
nand UO_2396 (O_2396,N_23698,N_21562);
or UO_2397 (O_2397,N_24524,N_20988);
nand UO_2398 (O_2398,N_18831,N_20240);
or UO_2399 (O_2399,N_23624,N_24628);
nor UO_2400 (O_2400,N_22040,N_21092);
nor UO_2401 (O_2401,N_23200,N_22144);
xnor UO_2402 (O_2402,N_23662,N_20128);
nor UO_2403 (O_2403,N_20920,N_24650);
nand UO_2404 (O_2404,N_21656,N_22850);
or UO_2405 (O_2405,N_22500,N_19501);
and UO_2406 (O_2406,N_19379,N_22402);
nand UO_2407 (O_2407,N_22613,N_24331);
nand UO_2408 (O_2408,N_19476,N_24534);
and UO_2409 (O_2409,N_20777,N_23170);
nor UO_2410 (O_2410,N_21195,N_22233);
and UO_2411 (O_2411,N_20712,N_19203);
or UO_2412 (O_2412,N_24368,N_24127);
and UO_2413 (O_2413,N_22356,N_20521);
or UO_2414 (O_2414,N_20167,N_21505);
nand UO_2415 (O_2415,N_24809,N_23042);
nor UO_2416 (O_2416,N_21426,N_22682);
or UO_2417 (O_2417,N_21853,N_19837);
nor UO_2418 (O_2418,N_21433,N_21616);
and UO_2419 (O_2419,N_21282,N_23153);
or UO_2420 (O_2420,N_22287,N_21779);
nand UO_2421 (O_2421,N_19071,N_22994);
nand UO_2422 (O_2422,N_19806,N_20379);
nand UO_2423 (O_2423,N_19991,N_22239);
nand UO_2424 (O_2424,N_23205,N_23834);
or UO_2425 (O_2425,N_21546,N_22187);
and UO_2426 (O_2426,N_24623,N_24659);
nand UO_2427 (O_2427,N_24733,N_21919);
nand UO_2428 (O_2428,N_23163,N_19597);
nor UO_2429 (O_2429,N_23807,N_24271);
nand UO_2430 (O_2430,N_20429,N_22606);
xnor UO_2431 (O_2431,N_19948,N_19546);
nor UO_2432 (O_2432,N_21858,N_24854);
nand UO_2433 (O_2433,N_24174,N_20435);
xor UO_2434 (O_2434,N_20053,N_23938);
and UO_2435 (O_2435,N_22801,N_21337);
and UO_2436 (O_2436,N_23901,N_21304);
nand UO_2437 (O_2437,N_23908,N_20378);
or UO_2438 (O_2438,N_18928,N_22618);
or UO_2439 (O_2439,N_22372,N_19486);
xnor UO_2440 (O_2440,N_19282,N_22997);
and UO_2441 (O_2441,N_23007,N_22117);
nand UO_2442 (O_2442,N_20488,N_21429);
and UO_2443 (O_2443,N_20329,N_21016);
and UO_2444 (O_2444,N_20236,N_24151);
nand UO_2445 (O_2445,N_18949,N_23286);
nor UO_2446 (O_2446,N_20823,N_22554);
nand UO_2447 (O_2447,N_19960,N_24475);
nand UO_2448 (O_2448,N_21013,N_24279);
nand UO_2449 (O_2449,N_21438,N_24985);
and UO_2450 (O_2450,N_24881,N_23479);
or UO_2451 (O_2451,N_24592,N_21178);
and UO_2452 (O_2452,N_20308,N_23978);
nor UO_2453 (O_2453,N_22371,N_21801);
and UO_2454 (O_2454,N_21706,N_20281);
or UO_2455 (O_2455,N_21984,N_19190);
nor UO_2456 (O_2456,N_19681,N_19717);
xnor UO_2457 (O_2457,N_21324,N_23836);
or UO_2458 (O_2458,N_24114,N_24513);
and UO_2459 (O_2459,N_18777,N_23454);
nand UO_2460 (O_2460,N_23922,N_19682);
and UO_2461 (O_2461,N_23209,N_24067);
nand UO_2462 (O_2462,N_21234,N_22010);
and UO_2463 (O_2463,N_24168,N_23155);
nor UO_2464 (O_2464,N_23712,N_22861);
nand UO_2465 (O_2465,N_21964,N_20965);
or UO_2466 (O_2466,N_21479,N_19694);
or UO_2467 (O_2467,N_24307,N_23088);
or UO_2468 (O_2468,N_21521,N_22282);
nand UO_2469 (O_2469,N_22674,N_22290);
nand UO_2470 (O_2470,N_21965,N_24832);
nand UO_2471 (O_2471,N_23851,N_19356);
nand UO_2472 (O_2472,N_23430,N_24593);
nand UO_2473 (O_2473,N_23232,N_19265);
nand UO_2474 (O_2474,N_19133,N_24172);
nand UO_2475 (O_2475,N_24163,N_23728);
xor UO_2476 (O_2476,N_23472,N_19891);
or UO_2477 (O_2477,N_23657,N_23326);
nor UO_2478 (O_2478,N_24297,N_21689);
and UO_2479 (O_2479,N_19550,N_21922);
nor UO_2480 (O_2480,N_21210,N_24680);
nor UO_2481 (O_2481,N_22080,N_23391);
xnor UO_2482 (O_2482,N_22107,N_22334);
xnor UO_2483 (O_2483,N_19563,N_22987);
nand UO_2484 (O_2484,N_22159,N_21372);
nor UO_2485 (O_2485,N_20503,N_23141);
and UO_2486 (O_2486,N_24322,N_19995);
or UO_2487 (O_2487,N_22183,N_23617);
and UO_2488 (O_2488,N_23433,N_20370);
nand UO_2489 (O_2489,N_21033,N_22086);
nand UO_2490 (O_2490,N_24539,N_20389);
and UO_2491 (O_2491,N_22053,N_23181);
nor UO_2492 (O_2492,N_21174,N_23320);
and UO_2493 (O_2493,N_23086,N_22318);
and UO_2494 (O_2494,N_20732,N_21400);
nand UO_2495 (O_2495,N_23956,N_22844);
or UO_2496 (O_2496,N_19953,N_22658);
or UO_2497 (O_2497,N_24145,N_19817);
nor UO_2498 (O_2498,N_24144,N_21808);
and UO_2499 (O_2499,N_19257,N_22105);
and UO_2500 (O_2500,N_23571,N_23207);
or UO_2501 (O_2501,N_20664,N_23671);
and UO_2502 (O_2502,N_23072,N_19871);
nor UO_2503 (O_2503,N_23372,N_21392);
nor UO_2504 (O_2504,N_19135,N_23880);
and UO_2505 (O_2505,N_23055,N_22970);
and UO_2506 (O_2506,N_22370,N_23090);
and UO_2507 (O_2507,N_24819,N_19562);
or UO_2508 (O_2508,N_20124,N_19367);
nand UO_2509 (O_2509,N_24494,N_23105);
and UO_2510 (O_2510,N_19437,N_19697);
nand UO_2511 (O_2511,N_24875,N_20042);
nand UO_2512 (O_2512,N_23993,N_22299);
nand UO_2513 (O_2513,N_21408,N_21062);
nand UO_2514 (O_2514,N_21676,N_20449);
nand UO_2515 (O_2515,N_22128,N_19338);
nand UO_2516 (O_2516,N_19266,N_24070);
and UO_2517 (O_2517,N_21364,N_20484);
nand UO_2518 (O_2518,N_23976,N_22420);
nand UO_2519 (O_2519,N_18846,N_22830);
and UO_2520 (O_2520,N_19091,N_20171);
nor UO_2521 (O_2521,N_23034,N_24358);
nand UO_2522 (O_2522,N_24933,N_20830);
and UO_2523 (O_2523,N_21476,N_20719);
or UO_2524 (O_2524,N_24717,N_20111);
nor UO_2525 (O_2525,N_23446,N_21273);
or UO_2526 (O_2526,N_24142,N_20002);
xor UO_2527 (O_2527,N_22350,N_23116);
and UO_2528 (O_2528,N_24765,N_19602);
nand UO_2529 (O_2529,N_21384,N_19605);
and UO_2530 (O_2530,N_19833,N_22312);
nor UO_2531 (O_2531,N_22654,N_22268);
and UO_2532 (O_2532,N_20581,N_18964);
or UO_2533 (O_2533,N_22857,N_23126);
nor UO_2534 (O_2534,N_24101,N_23900);
nand UO_2535 (O_2535,N_21577,N_20050);
nor UO_2536 (O_2536,N_24411,N_24611);
and UO_2537 (O_2537,N_23190,N_24301);
xor UO_2538 (O_2538,N_21074,N_19748);
xnor UO_2539 (O_2539,N_21875,N_19640);
nor UO_2540 (O_2540,N_24206,N_22218);
nand UO_2541 (O_2541,N_23242,N_24316);
nand UO_2542 (O_2542,N_20385,N_18988);
nor UO_2543 (O_2543,N_21758,N_22216);
nor UO_2544 (O_2544,N_24175,N_23282);
and UO_2545 (O_2545,N_21028,N_23522);
or UO_2546 (O_2546,N_22806,N_22175);
nand UO_2547 (O_2547,N_22295,N_21382);
nand UO_2548 (O_2548,N_20682,N_21110);
nand UO_2549 (O_2549,N_23118,N_23973);
xnor UO_2550 (O_2550,N_24482,N_24489);
nand UO_2551 (O_2551,N_21373,N_20062);
and UO_2552 (O_2552,N_18817,N_20918);
or UO_2553 (O_2553,N_21553,N_23222);
nor UO_2554 (O_2554,N_19132,N_23672);
nand UO_2555 (O_2555,N_21720,N_24087);
nor UO_2556 (O_2556,N_24574,N_20504);
or UO_2557 (O_2557,N_19507,N_21611);
or UO_2558 (O_2558,N_24037,N_20464);
nor UO_2559 (O_2559,N_22403,N_21506);
xnor UO_2560 (O_2560,N_21327,N_24672);
or UO_2561 (O_2561,N_21769,N_20566);
or UO_2562 (O_2562,N_20626,N_19867);
nor UO_2563 (O_2563,N_22620,N_23152);
and UO_2564 (O_2564,N_24135,N_24153);
nor UO_2565 (O_2565,N_20747,N_23444);
nor UO_2566 (O_2566,N_22872,N_23413);
nand UO_2567 (O_2567,N_22550,N_20736);
or UO_2568 (O_2568,N_19674,N_24176);
nor UO_2569 (O_2569,N_19852,N_21072);
or UO_2570 (O_2570,N_21708,N_19121);
nor UO_2571 (O_2571,N_24230,N_22846);
or UO_2572 (O_2572,N_21444,N_23707);
nor UO_2573 (O_2573,N_21782,N_22951);
nand UO_2574 (O_2574,N_22162,N_24699);
nor UO_2575 (O_2575,N_21805,N_19997);
xor UO_2576 (O_2576,N_20438,N_19510);
or UO_2577 (O_2577,N_20640,N_21570);
nor UO_2578 (O_2578,N_18855,N_20205);
nor UO_2579 (O_2579,N_22802,N_20213);
or UO_2580 (O_2580,N_20576,N_21986);
nand UO_2581 (O_2581,N_22524,N_21519);
nor UO_2582 (O_2582,N_24187,N_20935);
or UO_2583 (O_2583,N_20045,N_24529);
or UO_2584 (O_2584,N_18957,N_18827);
nand UO_2585 (O_2585,N_24081,N_21523);
nand UO_2586 (O_2586,N_23588,N_19869);
nor UO_2587 (O_2587,N_23228,N_21756);
nand UO_2588 (O_2588,N_23539,N_24289);
nand UO_2589 (O_2589,N_20283,N_24023);
and UO_2590 (O_2590,N_20162,N_23469);
or UO_2591 (O_2591,N_19212,N_22967);
or UO_2592 (O_2592,N_22432,N_21278);
nor UO_2593 (O_2593,N_24523,N_19773);
nand UO_2594 (O_2594,N_22257,N_19950);
nor UO_2595 (O_2595,N_21100,N_24814);
nor UO_2596 (O_2596,N_22456,N_19693);
nand UO_2597 (O_2597,N_22928,N_20872);
or UO_2598 (O_2598,N_20349,N_18905);
or UO_2599 (O_2599,N_23191,N_18929);
nor UO_2600 (O_2600,N_20657,N_20707);
or UO_2601 (O_2601,N_20189,N_22369);
or UO_2602 (O_2602,N_18830,N_19219);
and UO_2603 (O_2603,N_22579,N_24007);
nor UO_2604 (O_2604,N_24329,N_22699);
nor UO_2605 (O_2605,N_22859,N_21423);
nand UO_2606 (O_2606,N_21345,N_20532);
and UO_2607 (O_2607,N_22950,N_24287);
or UO_2608 (O_2608,N_23324,N_21923);
nand UO_2609 (O_2609,N_20628,N_21556);
xor UO_2610 (O_2610,N_21241,N_24905);
nand UO_2611 (O_2611,N_24059,N_23590);
nor UO_2612 (O_2612,N_24880,N_22394);
and UO_2613 (O_2613,N_21052,N_19279);
nand UO_2614 (O_2614,N_24625,N_24506);
nor UO_2615 (O_2615,N_22900,N_20483);
nor UO_2616 (O_2616,N_18797,N_24136);
nand UO_2617 (O_2617,N_24634,N_21003);
nand UO_2618 (O_2618,N_19208,N_22957);
xnor UO_2619 (O_2619,N_24491,N_22630);
nand UO_2620 (O_2620,N_22598,N_21785);
and UO_2621 (O_2621,N_23477,N_24088);
and UO_2622 (O_2622,N_23931,N_24061);
nand UO_2623 (O_2623,N_19633,N_20251);
xnor UO_2624 (O_2624,N_24474,N_22358);
or UO_2625 (O_2625,N_23188,N_20330);
and UO_2626 (O_2626,N_21648,N_19895);
nor UO_2627 (O_2627,N_22622,N_21880);
nor UO_2628 (O_2628,N_19926,N_21308);
and UO_2629 (O_2629,N_22783,N_24936);
xnor UO_2630 (O_2630,N_23327,N_22760);
nor UO_2631 (O_2631,N_21630,N_20439);
or UO_2632 (O_2632,N_20344,N_22960);
nand UO_2633 (O_2633,N_22854,N_20697);
nand UO_2634 (O_2634,N_23936,N_23537);
nand UO_2635 (O_2635,N_19273,N_23824);
and UO_2636 (O_2636,N_21641,N_22419);
nor UO_2637 (O_2637,N_20584,N_20494);
nor UO_2638 (O_2638,N_21088,N_22822);
xor UO_2639 (O_2639,N_24843,N_24619);
nand UO_2640 (O_2640,N_20094,N_18857);
xnor UO_2641 (O_2641,N_24753,N_20369);
nand UO_2642 (O_2642,N_23696,N_20688);
and UO_2643 (O_2643,N_21097,N_23795);
nand UO_2644 (O_2644,N_20666,N_20271);
nand UO_2645 (O_2645,N_22112,N_22816);
and UO_2646 (O_2646,N_20160,N_20961);
nand UO_2647 (O_2647,N_22204,N_24945);
or UO_2648 (O_2648,N_24877,N_22731);
or UO_2649 (O_2649,N_19426,N_20263);
nor UO_2650 (O_2650,N_23419,N_19497);
nand UO_2651 (O_2651,N_22479,N_21375);
nor UO_2652 (O_2652,N_24641,N_23159);
and UO_2653 (O_2653,N_21125,N_21120);
nor UO_2654 (O_2654,N_24062,N_22424);
nor UO_2655 (O_2655,N_19531,N_19173);
or UO_2656 (O_2656,N_22493,N_18967);
or UO_2657 (O_2657,N_18956,N_21388);
nand UO_2658 (O_2658,N_24463,N_22440);
or UO_2659 (O_2659,N_19206,N_23290);
or UO_2660 (O_2660,N_21263,N_21584);
and UO_2661 (O_2661,N_23506,N_22137);
nand UO_2662 (O_2662,N_21726,N_24590);
or UO_2663 (O_2663,N_19866,N_18892);
and UO_2664 (O_2664,N_20227,N_22516);
nor UO_2665 (O_2665,N_20554,N_20082);
nand UO_2666 (O_2666,N_19915,N_19452);
nand UO_2667 (O_2667,N_23760,N_24797);
and UO_2668 (O_2668,N_19872,N_19730);
and UO_2669 (O_2669,N_23951,N_19312);
nand UO_2670 (O_2670,N_21193,N_22423);
and UO_2671 (O_2671,N_22969,N_24859);
and UO_2672 (O_2672,N_20470,N_22457);
nand UO_2673 (O_2673,N_19369,N_20694);
xor UO_2674 (O_2674,N_21586,N_19052);
nor UO_2675 (O_2675,N_19526,N_23460);
nor UO_2676 (O_2676,N_21251,N_22988);
or UO_2677 (O_2677,N_20881,N_22066);
or UO_2678 (O_2678,N_23468,N_21008);
or UO_2679 (O_2679,N_24233,N_23687);
nor UO_2680 (O_2680,N_20075,N_24025);
and UO_2681 (O_2681,N_21578,N_20027);
or UO_2682 (O_2682,N_20152,N_23866);
or UO_2683 (O_2683,N_23134,N_19409);
nor UO_2684 (O_2684,N_20711,N_24259);
xor UO_2685 (O_2685,N_23966,N_19402);
nand UO_2686 (O_2686,N_24565,N_21820);
nand UO_2687 (O_2687,N_23201,N_19559);
nor UO_2688 (O_2688,N_23632,N_21814);
xor UO_2689 (O_2689,N_23408,N_21184);
or UO_2690 (O_2690,N_22413,N_20408);
or UO_2691 (O_2691,N_23028,N_24055);
nor UO_2692 (O_2692,N_20674,N_21542);
xnor UO_2693 (O_2693,N_23572,N_23245);
nand UO_2694 (O_2694,N_22411,N_24213);
nor UO_2695 (O_2695,N_23031,N_20517);
nand UO_2696 (O_2696,N_23291,N_20863);
nor UO_2697 (O_2697,N_23928,N_23164);
xor UO_2698 (O_2698,N_22542,N_19619);
and UO_2699 (O_2699,N_22561,N_20526);
and UO_2700 (O_2700,N_21115,N_21070);
nor UO_2701 (O_2701,N_21552,N_20325);
xnor UO_2702 (O_2702,N_19785,N_21339);
xnor UO_2703 (O_2703,N_19718,N_22545);
and UO_2704 (O_2704,N_22154,N_23516);
xor UO_2705 (O_2705,N_21434,N_24723);
and UO_2706 (O_2706,N_19519,N_24022);
and UO_2707 (O_2707,N_21451,N_21781);
nand UO_2708 (O_2708,N_24333,N_20083);
and UO_2709 (O_2709,N_19727,N_23014);
nand UO_2710 (O_2710,N_21843,N_23597);
nand UO_2711 (O_2711,N_23041,N_22780);
and UO_2712 (O_2712,N_18842,N_19938);
nand UO_2713 (O_2713,N_19719,N_23046);
and UO_2714 (O_2714,N_23458,N_19428);
or UO_2715 (O_2715,N_24850,N_19529);
nor UO_2716 (O_2716,N_18758,N_21101);
and UO_2717 (O_2717,N_20116,N_24381);
and UO_2718 (O_2718,N_20622,N_23697);
and UO_2719 (O_2719,N_24050,N_23518);
and UO_2720 (O_2720,N_20529,N_24181);
nand UO_2721 (O_2721,N_23945,N_21997);
nor UO_2722 (O_2722,N_24033,N_23850);
xnor UO_2723 (O_2723,N_19422,N_24352);
nand UO_2724 (O_2724,N_20183,N_24091);
nor UO_2725 (O_2725,N_21113,N_23927);
and UO_2726 (O_2726,N_20857,N_24889);
or UO_2727 (O_2727,N_19405,N_24173);
and UO_2728 (O_2728,N_24943,N_24967);
nand UO_2729 (O_2729,N_23933,N_23875);
and UO_2730 (O_2730,N_22605,N_22800);
nor UO_2731 (O_2731,N_21360,N_23019);
nand UO_2732 (O_2732,N_20323,N_23056);
nor UO_2733 (O_2733,N_21982,N_24016);
or UO_2734 (O_2734,N_22729,N_23653);
nor UO_2735 (O_2735,N_19377,N_19527);
and UO_2736 (O_2736,N_20231,N_20866);
nand UO_2737 (O_2737,N_21839,N_19242);
or UO_2738 (O_2738,N_24299,N_22106);
nor UO_2739 (O_2739,N_19945,N_22007);
xor UO_2740 (O_2740,N_20176,N_24018);
nand UO_2741 (O_2741,N_23462,N_22050);
nor UO_2742 (O_2742,N_24257,N_24771);
xor UO_2743 (O_2743,N_19770,N_20858);
nand UO_2744 (O_2744,N_19129,N_19961);
nor UO_2745 (O_2745,N_20855,N_20181);
or UO_2746 (O_2746,N_22555,N_22503);
nor UO_2747 (O_2747,N_19374,N_24351);
nor UO_2748 (O_2748,N_23881,N_19880);
and UO_2749 (O_2749,N_20074,N_22125);
nand UO_2750 (O_2750,N_19127,N_22392);
nor UO_2751 (O_2751,N_21995,N_20931);
nor UO_2752 (O_2752,N_20025,N_20599);
nand UO_2753 (O_2753,N_22905,N_20012);
and UO_2754 (O_2754,N_19058,N_20233);
and UO_2755 (O_2755,N_19757,N_22221);
or UO_2756 (O_2756,N_22559,N_23070);
nand UO_2757 (O_2757,N_18815,N_23285);
nor UO_2758 (O_2758,N_18890,N_24687);
nor UO_2759 (O_2759,N_23637,N_18865);
nand UO_2760 (O_2760,N_21060,N_18974);
nand UO_2761 (O_2761,N_24538,N_19335);
or UO_2762 (O_2762,N_24304,N_19536);
and UO_2763 (O_2763,N_21145,N_21054);
and UO_2764 (O_2764,N_22205,N_22215);
or UO_2765 (O_2765,N_23988,N_21531);
and UO_2766 (O_2766,N_22738,N_21081);
or UO_2767 (O_2767,N_24315,N_23581);
nor UO_2768 (O_2768,N_22640,N_24511);
and UO_2769 (O_2769,N_19528,N_20533);
or UO_2770 (O_2770,N_22418,N_21498);
or UO_2771 (O_2771,N_24575,N_21152);
xnor UO_2772 (O_2772,N_19864,N_24893);
nand UO_2773 (O_2773,N_24605,N_20066);
or UO_2774 (O_2774,N_21811,N_21692);
nand UO_2775 (O_2775,N_24413,N_23839);
and UO_2776 (O_2776,N_20940,N_20478);
nor UO_2777 (O_2777,N_18838,N_23842);
nor UO_2778 (O_2778,N_19084,N_23025);
nand UO_2779 (O_2779,N_19216,N_20203);
and UO_2780 (O_2780,N_23186,N_23623);
nor UO_2781 (O_2781,N_19375,N_18811);
and UO_2782 (O_2782,N_24118,N_20238);
nor UO_2783 (O_2783,N_21848,N_24481);
xor UO_2784 (O_2784,N_19471,N_21931);
nand UO_2785 (O_2785,N_19564,N_18813);
nand UO_2786 (O_2786,N_20838,N_18924);
or UO_2787 (O_2787,N_21563,N_24318);
or UO_2788 (O_2788,N_22484,N_18981);
nand UO_2789 (O_2789,N_23022,N_19432);
nor UO_2790 (O_2790,N_20069,N_24004);
nor UO_2791 (O_2791,N_22223,N_22868);
and UO_2792 (O_2792,N_20132,N_20826);
and UO_2793 (O_2793,N_24388,N_18825);
xnor UO_2794 (O_2794,N_19784,N_24195);
nand UO_2795 (O_2795,N_22396,N_20601);
and UO_2796 (O_2796,N_19971,N_23198);
xnor UO_2797 (O_2797,N_21764,N_20102);
nand UO_2798 (O_2798,N_22442,N_22431);
and UO_2799 (O_2799,N_24567,N_23582);
nand UO_2800 (O_2800,N_21046,N_20574);
nor UO_2801 (O_2801,N_24239,N_21594);
nor UO_2802 (O_2802,N_22489,N_24340);
nor UO_2803 (O_2803,N_22927,N_19094);
or UO_2804 (O_2804,N_22048,N_23199);
or UO_2805 (O_2805,N_19782,N_21538);
xor UO_2806 (O_2806,N_24036,N_21626);
or UO_2807 (O_2807,N_20487,N_24487);
nor UO_2808 (O_2808,N_22525,N_20583);
and UO_2809 (O_2809,N_22840,N_23154);
xor UO_2810 (O_2810,N_19701,N_22809);
and UO_2811 (O_2811,N_23905,N_21524);
or UO_2812 (O_2812,N_21741,N_24742);
nand UO_2813 (O_2813,N_24051,N_19811);
nor UO_2814 (O_2814,N_20159,N_19816);
or UO_2815 (O_2815,N_20374,N_20775);
and UO_2816 (O_2816,N_23694,N_21543);
nand UO_2817 (O_2817,N_19590,N_23604);
nand UO_2818 (O_2818,N_18755,N_20721);
nand UO_2819 (O_2819,N_23718,N_21561);
or UO_2820 (O_2820,N_20011,N_24060);
and UO_2821 (O_2821,N_19803,N_20423);
nor UO_2822 (O_2822,N_24727,N_18807);
xnor UO_2823 (O_2823,N_23514,N_24353);
and UO_2824 (O_2824,N_23382,N_24125);
xnor UO_2825 (O_2825,N_19021,N_22534);
nor UO_2826 (O_2826,N_20999,N_23437);
nor UO_2827 (O_2827,N_21564,N_22227);
and UO_2828 (O_2828,N_22116,N_18938);
and UO_2829 (O_2829,N_23237,N_19077);
nand UO_2830 (O_2830,N_24476,N_22508);
and UO_2831 (O_2831,N_19962,N_21949);
and UO_2832 (O_2832,N_23549,N_24561);
nand UO_2833 (O_2833,N_23847,N_21402);
and UO_2834 (O_2834,N_22781,N_24300);
nor UO_2835 (O_2835,N_21746,N_23919);
nor UO_2836 (O_2836,N_19731,N_23455);
nand UO_2837 (O_2837,N_23517,N_23484);
and UO_2838 (O_2838,N_24683,N_19474);
nand UO_2839 (O_2839,N_23764,N_20313);
nor UO_2840 (O_2840,N_24999,N_22179);
nand UO_2841 (O_2841,N_23673,N_20916);
nand UO_2842 (O_2842,N_22539,N_24214);
and UO_2843 (O_2843,N_23743,N_24579);
nand UO_2844 (O_2844,N_20456,N_22301);
or UO_2845 (O_2845,N_20334,N_21933);
or UO_2846 (O_2846,N_19416,N_19567);
or UO_2847 (O_2847,N_19829,N_24367);
nand UO_2848 (O_2848,N_24761,N_19807);
nand UO_2849 (O_2849,N_22006,N_24925);
nor UO_2850 (O_2850,N_22207,N_19951);
nor UO_2851 (O_2851,N_24232,N_22091);
nand UO_2852 (O_2852,N_20976,N_20033);
nand UO_2853 (O_2853,N_19612,N_20897);
xnor UO_2854 (O_2854,N_19651,N_21650);
nand UO_2855 (O_2855,N_22249,N_21829);
xnor UO_2856 (O_2856,N_19653,N_21744);
and UO_2857 (O_2857,N_24756,N_19440);
nand UO_2858 (O_2858,N_22374,N_23099);
nand UO_2859 (O_2859,N_20859,N_24830);
xnor UO_2860 (O_2860,N_21255,N_24117);
or UO_2861 (O_2861,N_20145,N_24075);
nor UO_2862 (O_2862,N_22667,N_24633);
nor UO_2863 (O_2863,N_19708,N_23301);
nor UO_2864 (O_2864,N_24365,N_20865);
and UO_2865 (O_2865,N_23726,N_22513);
nor UO_2866 (O_2866,N_19779,N_21535);
or UO_2867 (O_2867,N_24658,N_22388);
nor UO_2868 (O_2868,N_23636,N_19294);
nor UO_2869 (O_2869,N_24110,N_20779);
or UO_2870 (O_2870,N_23067,N_23036);
nor UO_2871 (O_2871,N_20091,N_20815);
nand UO_2872 (O_2872,N_21838,N_21589);
xnor UO_2873 (O_2873,N_24109,N_23544);
or UO_2874 (O_2874,N_20675,N_18941);
nand UO_2875 (O_2875,N_24319,N_22309);
nand UO_2876 (O_2876,N_23225,N_22725);
or UO_2877 (O_2877,N_20824,N_20705);
xor UO_2878 (O_2878,N_18916,N_24216);
or UO_2879 (O_2879,N_19223,N_24903);
nor UO_2880 (O_2880,N_22883,N_22087);
or UO_2881 (O_2881,N_20656,N_21681);
nor UO_2882 (O_2882,N_21972,N_20774);
nor UO_2883 (O_2883,N_24458,N_22610);
and UO_2884 (O_2884,N_21776,N_23052);
and UO_2885 (O_2885,N_22348,N_20191);
and UO_2886 (O_2886,N_21415,N_24584);
xnor UO_2887 (O_2887,N_22526,N_19514);
nor UO_2888 (O_2888,N_23819,N_22765);
nor UO_2889 (O_2889,N_19722,N_19709);
and UO_2890 (O_2890,N_20332,N_18768);
nor UO_2891 (O_2891,N_21845,N_22856);
xor UO_2892 (O_2892,N_22675,N_20927);
nand UO_2893 (O_2893,N_20915,N_19388);
and UO_2894 (O_2894,N_23388,N_19222);
or UO_2895 (O_2895,N_20247,N_19184);
nor UO_2896 (O_2896,N_21520,N_24791);
nand UO_2897 (O_2897,N_20975,N_21844);
and UO_2898 (O_2898,N_19002,N_20490);
nand UO_2899 (O_2899,N_24167,N_24426);
or UO_2900 (O_2900,N_20170,N_19934);
or UO_2901 (O_2901,N_22558,N_19447);
and UO_2902 (O_2902,N_22829,N_22267);
nor UO_2903 (O_2903,N_22540,N_19912);
nor UO_2904 (O_2904,N_21105,N_21465);
and UO_2905 (O_2905,N_24412,N_23788);
xnor UO_2906 (O_2906,N_19593,N_24677);
nor UO_2907 (O_2907,N_22055,N_22601);
or UO_2908 (O_2908,N_18757,N_22717);
or UO_2909 (O_2909,N_22464,N_21477);
nor UO_2910 (O_2910,N_24763,N_21038);
or UO_2911 (O_2911,N_21191,N_23108);
and UO_2912 (O_2912,N_23385,N_21055);
or UO_2913 (O_2913,N_20328,N_23157);
nand UO_2914 (O_2914,N_23463,N_21172);
xnor UO_2915 (O_2915,N_24479,N_20381);
nor UO_2916 (O_2916,N_20001,N_20064);
nand UO_2917 (O_2917,N_20472,N_19415);
nor UO_2918 (O_2918,N_22538,N_19043);
nand UO_2919 (O_2919,N_19511,N_21050);
xnor UO_2920 (O_2920,N_21504,N_19931);
nor UO_2921 (O_2921,N_22272,N_24535);
nor UO_2922 (O_2922,N_21252,N_19739);
xor UO_2923 (O_2923,N_24094,N_19063);
or UO_2924 (O_2924,N_24359,N_23029);
nor UO_2925 (O_2925,N_21133,N_19138);
and UO_2926 (O_2926,N_24965,N_22497);
nor UO_2927 (O_2927,N_18782,N_21090);
xor UO_2928 (O_2928,N_24237,N_20906);
or UO_2929 (O_2929,N_21612,N_19241);
and UO_2930 (O_2930,N_18764,N_19269);
xor UO_2931 (O_2931,N_21799,N_21593);
nor UO_2932 (O_2932,N_21305,N_21939);
nor UO_2933 (O_2933,N_20256,N_18887);
xor UO_2934 (O_2934,N_19680,N_21075);
nand UO_2935 (O_2935,N_24032,N_20539);
nor UO_2936 (O_2936,N_21609,N_24556);
or UO_2937 (O_2937,N_23761,N_21750);
or UO_2938 (O_2938,N_22818,N_21262);
nor UO_2939 (O_2939,N_23635,N_23832);
xor UO_2940 (O_2940,N_23347,N_22590);
nor UO_2941 (O_2941,N_24836,N_22596);
nor UO_2942 (O_2942,N_21635,N_19606);
nand UO_2943 (O_2943,N_18775,N_24392);
nand UO_2944 (O_2944,N_24152,N_23541);
nand UO_2945 (O_2945,N_21802,N_19413);
nand UO_2946 (O_2946,N_21175,N_22071);
and UO_2947 (O_2947,N_21952,N_21190);
nor UO_2948 (O_2948,N_21784,N_24786);
xnor UO_2949 (O_2949,N_23682,N_22029);
or UO_2950 (O_2950,N_23331,N_24527);
xnor UO_2951 (O_2951,N_20289,N_20475);
nand UO_2952 (O_2952,N_21610,N_24910);
nor UO_2953 (O_2953,N_24899,N_21067);
and UO_2954 (O_2954,N_23492,N_19552);
and UO_2955 (O_2955,N_21895,N_23238);
xnor UO_2956 (O_2956,N_22621,N_22755);
and UO_2957 (O_2957,N_23641,N_22989);
and UO_2958 (O_2958,N_22977,N_21700);
nand UO_2959 (O_2959,N_23902,N_24648);
nand UO_2960 (O_2960,N_20118,N_22845);
nor UO_2961 (O_2961,N_24615,N_23396);
or UO_2962 (O_2962,N_20665,N_19560);
or UO_2963 (O_2963,N_24794,N_19100);
nand UO_2964 (O_2964,N_22002,N_19796);
nor UO_2965 (O_2965,N_21049,N_20522);
nor UO_2966 (O_2966,N_22941,N_24402);
nor UO_2967 (O_2967,N_23546,N_19607);
and UO_2968 (O_2968,N_23913,N_23861);
or UO_2969 (O_2969,N_18979,N_24423);
nand UO_2970 (O_2970,N_23475,N_21980);
or UO_2971 (O_2971,N_22746,N_21794);
nor UO_2972 (O_2972,N_23699,N_23069);
or UO_2973 (O_2973,N_21925,N_23091);
nand UO_2974 (O_2974,N_24355,N_24688);
nor UO_2975 (O_2975,N_19368,N_22608);
nor UO_2976 (O_2976,N_22889,N_21192);
nor UO_2977 (O_2977,N_22405,N_24792);
nor UO_2978 (O_2978,N_20292,N_19387);
nand UO_2979 (O_2979,N_24663,N_20474);
nand UO_2980 (O_2980,N_19603,N_23611);
or UO_2981 (O_2981,N_21325,N_22335);
nand UO_2982 (O_2982,N_22719,N_24596);
and UO_2983 (O_2983,N_21890,N_23789);
and UO_2984 (O_2984,N_23558,N_19451);
and UO_2985 (O_2985,N_21981,N_20671);
or UO_2986 (O_2986,N_19714,N_23686);
nand UO_2987 (O_2987,N_22663,N_19824);
nand UO_2988 (O_2988,N_23912,N_22824);
or UO_2989 (O_2989,N_24695,N_22803);
nand UO_2990 (O_2990,N_19101,N_23257);
xor UO_2991 (O_2991,N_21370,N_23314);
and UO_2992 (O_2992,N_20869,N_24701);
nor UO_2993 (O_2993,N_21525,N_20031);
nand UO_2994 (O_2994,N_20052,N_20364);
or UO_2995 (O_2995,N_24953,N_19404);
and UO_2996 (O_2996,N_23942,N_24245);
or UO_2997 (O_2997,N_23356,N_21164);
or UO_2998 (O_2998,N_23379,N_21809);
nor UO_2999 (O_2999,N_24586,N_18921);
endmodule