module basic_1000_10000_1500_10_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_478,In_764);
and U1 (N_1,In_297,In_771);
and U2 (N_2,In_636,In_65);
nor U3 (N_3,In_546,In_282);
nor U4 (N_4,In_507,In_279);
or U5 (N_5,In_44,In_390);
and U6 (N_6,In_275,In_866);
and U7 (N_7,In_717,In_990);
nor U8 (N_8,In_105,In_694);
and U9 (N_9,In_642,In_899);
nor U10 (N_10,In_765,In_976);
nand U11 (N_11,In_502,In_79);
and U12 (N_12,In_691,In_595);
and U13 (N_13,In_808,In_85);
nor U14 (N_14,In_534,In_201);
or U15 (N_15,In_157,In_950);
and U16 (N_16,In_592,In_22);
and U17 (N_17,In_593,In_837);
or U18 (N_18,In_224,In_653);
or U19 (N_19,In_823,In_621);
nand U20 (N_20,In_613,In_999);
nand U21 (N_21,In_370,In_409);
or U22 (N_22,In_570,In_294);
and U23 (N_23,In_206,In_780);
nand U24 (N_24,In_934,In_795);
nor U25 (N_25,In_721,In_56);
nor U26 (N_26,In_715,In_188);
or U27 (N_27,In_973,In_988);
nor U28 (N_28,In_601,In_365);
and U29 (N_29,In_214,In_357);
nand U30 (N_30,In_567,In_213);
and U31 (N_31,In_371,In_217);
or U32 (N_32,In_413,In_623);
or U33 (N_33,In_920,In_865);
or U34 (N_34,In_941,In_710);
xnor U35 (N_35,In_464,In_838);
nor U36 (N_36,In_514,In_175);
and U37 (N_37,In_802,In_805);
nand U38 (N_38,In_665,In_652);
nand U39 (N_39,In_947,In_385);
and U40 (N_40,In_202,In_151);
xnor U41 (N_41,In_733,In_477);
and U42 (N_42,In_679,In_933);
nand U43 (N_43,In_907,In_504);
and U44 (N_44,In_871,In_542);
nand U45 (N_45,In_264,In_460);
or U46 (N_46,In_255,In_7);
xnor U47 (N_47,In_944,In_482);
or U48 (N_48,In_749,In_379);
or U49 (N_49,In_20,In_982);
or U50 (N_50,In_82,In_673);
xnor U51 (N_51,In_73,In_954);
and U52 (N_52,In_353,In_801);
nand U53 (N_53,In_468,In_156);
nor U54 (N_54,In_616,In_298);
xor U55 (N_55,In_868,In_195);
xnor U56 (N_56,In_760,In_955);
and U57 (N_57,In_342,In_359);
nor U58 (N_58,In_28,In_720);
and U59 (N_59,In_582,In_212);
nand U60 (N_60,In_905,In_698);
xnor U61 (N_61,In_166,In_355);
nand U62 (N_62,In_26,In_538);
or U63 (N_63,In_554,In_18);
xor U64 (N_64,In_654,In_853);
nand U65 (N_65,In_713,In_311);
nand U66 (N_66,In_927,In_740);
nor U67 (N_67,In_290,In_533);
nand U68 (N_68,In_518,In_141);
or U69 (N_69,In_626,In_800);
or U70 (N_70,In_932,In_919);
nor U71 (N_71,In_776,In_492);
nor U72 (N_72,In_576,In_544);
nor U73 (N_73,In_272,In_895);
nor U74 (N_74,In_378,In_640);
nand U75 (N_75,In_131,In_313);
or U76 (N_76,In_452,In_814);
and U77 (N_77,In_494,In_872);
and U78 (N_78,In_309,In_936);
and U79 (N_79,In_662,In_418);
nand U80 (N_80,In_364,In_742);
nor U81 (N_81,In_816,In_967);
xor U82 (N_82,In_671,In_268);
nor U83 (N_83,In_351,In_403);
xor U84 (N_84,In_47,In_387);
and U85 (N_85,In_414,In_92);
or U86 (N_86,In_590,In_322);
and U87 (N_87,In_394,In_366);
nor U88 (N_88,In_467,In_625);
nand U89 (N_89,In_685,In_83);
xnor U90 (N_90,In_968,In_909);
or U91 (N_91,In_335,In_10);
nand U92 (N_92,In_885,In_634);
and U93 (N_93,In_887,In_957);
and U94 (N_94,In_144,In_500);
and U95 (N_95,In_74,In_894);
or U96 (N_96,In_13,In_793);
nand U97 (N_97,In_64,In_90);
nand U98 (N_98,In_664,In_556);
nor U99 (N_99,In_123,In_462);
nor U100 (N_100,In_598,In_633);
nand U101 (N_101,In_273,In_856);
nand U102 (N_102,In_843,In_261);
nor U103 (N_103,In_750,In_903);
and U104 (N_104,In_263,In_741);
or U105 (N_105,In_122,In_71);
or U106 (N_106,In_532,In_864);
nand U107 (N_107,In_429,In_66);
and U108 (N_108,In_454,In_411);
nor U109 (N_109,In_343,In_812);
or U110 (N_110,In_984,In_882);
nor U111 (N_111,In_997,In_833);
xor U112 (N_112,In_483,In_228);
nand U113 (N_113,In_744,In_761);
nand U114 (N_114,In_408,In_316);
nor U115 (N_115,In_908,In_35);
nand U116 (N_116,In_945,In_381);
nand U117 (N_117,In_134,In_553);
nand U118 (N_118,In_680,In_3);
nor U119 (N_119,In_846,In_215);
nor U120 (N_120,In_998,In_325);
nor U121 (N_121,In_915,In_589);
nand U122 (N_122,In_101,In_9);
xor U123 (N_123,In_31,In_963);
xnor U124 (N_124,In_980,In_619);
nand U125 (N_125,In_398,In_471);
and U126 (N_126,In_291,In_515);
xnor U127 (N_127,In_961,In_250);
nor U128 (N_128,In_172,In_610);
and U129 (N_129,In_407,In_327);
nand U130 (N_130,In_916,In_667);
nand U131 (N_131,In_243,In_918);
and U132 (N_132,In_643,In_964);
or U133 (N_133,In_374,In_178);
or U134 (N_134,In_736,In_148);
and U135 (N_135,In_480,In_989);
and U136 (N_136,In_981,In_987);
and U137 (N_137,In_438,In_375);
nor U138 (N_138,In_937,In_17);
or U139 (N_139,In_284,In_177);
nor U140 (N_140,In_239,In_840);
and U141 (N_141,In_774,In_752);
nor U142 (N_142,In_786,In_705);
nor U143 (N_143,In_179,In_581);
nand U144 (N_144,In_266,In_149);
or U145 (N_145,In_373,In_824);
nand U146 (N_146,In_873,In_23);
and U147 (N_147,In_116,In_139);
nand U148 (N_148,In_701,In_169);
and U149 (N_149,In_707,In_946);
and U150 (N_150,In_96,In_883);
or U151 (N_151,In_182,In_29);
and U152 (N_152,In_611,In_734);
and U153 (N_153,In_524,In_726);
or U154 (N_154,In_425,In_614);
nand U155 (N_155,In_986,In_854);
and U156 (N_156,In_314,In_146);
or U157 (N_157,In_333,In_550);
nor U158 (N_158,In_221,In_227);
and U159 (N_159,In_42,In_681);
or U160 (N_160,In_531,In_706);
or U161 (N_161,In_830,In_458);
xnor U162 (N_162,In_995,In_84);
nor U163 (N_163,In_857,In_953);
or U164 (N_164,In_389,In_265);
xor U165 (N_165,In_498,In_756);
nand U166 (N_166,In_155,In_991);
nand U167 (N_167,In_847,In_310);
or U168 (N_168,In_348,In_484);
xor U169 (N_169,In_129,In_574);
nand U170 (N_170,In_645,In_39);
and U171 (N_171,In_433,In_861);
or U172 (N_172,In_216,In_49);
xnor U173 (N_173,In_815,In_490);
nor U174 (N_174,In_441,In_759);
nor U175 (N_175,In_91,In_748);
nand U176 (N_176,In_682,In_472);
nand U177 (N_177,In_575,In_296);
nand U178 (N_178,In_474,In_540);
nor U179 (N_179,In_410,In_60);
or U180 (N_180,In_395,In_925);
or U181 (N_181,In_930,In_12);
nand U182 (N_182,In_778,In_331);
nand U183 (N_183,In_597,In_246);
and U184 (N_184,In_200,In_770);
or U185 (N_185,In_822,In_676);
and U186 (N_186,In_170,In_97);
or U187 (N_187,In_627,In_184);
nor U188 (N_188,In_639,In_525);
nand U189 (N_189,In_807,In_696);
nor U190 (N_190,In_666,In_863);
and U191 (N_191,In_826,In_347);
or U192 (N_192,In_496,In_158);
and U193 (N_193,In_469,In_449);
or U194 (N_194,In_503,In_450);
nor U195 (N_195,In_160,In_768);
nand U196 (N_196,In_168,In_161);
xor U197 (N_197,In_324,In_948);
xnor U198 (N_198,In_700,In_154);
or U199 (N_199,In_399,In_361);
or U200 (N_200,In_704,In_209);
nor U201 (N_201,In_631,In_307);
nand U202 (N_202,In_448,In_612);
nand U203 (N_203,In_784,In_539);
and U204 (N_204,In_295,In_236);
or U205 (N_205,In_545,In_677);
nand U206 (N_206,In_607,In_881);
nand U207 (N_207,In_650,In_232);
or U208 (N_208,In_929,In_259);
or U209 (N_209,In_943,In_339);
nor U210 (N_210,In_505,In_152);
or U211 (N_211,In_896,In_183);
xor U212 (N_212,In_420,In_804);
xnor U213 (N_213,In_638,In_811);
nand U214 (N_214,In_110,In_779);
or U215 (N_215,In_488,In_289);
nor U216 (N_216,In_572,In_162);
nand U217 (N_217,In_360,In_497);
and U218 (N_218,In_208,In_11);
nor U219 (N_219,In_535,In_439);
nand U220 (N_220,In_893,In_218);
nand U221 (N_221,In_940,In_569);
xor U222 (N_222,In_321,In_842);
xnor U223 (N_223,In_692,In_262);
nand U224 (N_224,In_855,In_58);
and U225 (N_225,In_789,In_32);
or U226 (N_226,In_862,In_57);
and U227 (N_227,In_878,In_120);
and U228 (N_228,In_405,In_649);
nor U229 (N_229,In_495,In_41);
and U230 (N_230,In_98,In_147);
nor U231 (N_231,In_820,In_251);
nand U232 (N_232,In_53,In_536);
or U233 (N_233,In_580,In_992);
nand U234 (N_234,In_302,In_4);
or U235 (N_235,In_821,In_111);
or U236 (N_236,In_94,In_782);
nand U237 (N_237,In_848,In_668);
nand U238 (N_238,In_76,In_788);
and U239 (N_239,In_541,In_102);
nor U240 (N_240,In_70,In_318);
and U241 (N_241,In_799,In_329);
and U242 (N_242,In_876,In_248);
nor U243 (N_243,In_443,In_465);
or U244 (N_244,In_103,In_113);
nand U245 (N_245,In_978,In_605);
nand U246 (N_246,In_180,In_869);
or U247 (N_247,In_521,In_16);
and U248 (N_248,In_697,In_813);
and U249 (N_249,In_796,In_972);
or U250 (N_250,In_763,In_655);
nor U251 (N_251,In_245,In_527);
and U252 (N_252,In_253,In_529);
and U253 (N_253,In_234,In_277);
nand U254 (N_254,In_693,In_426);
or U255 (N_255,In_437,In_660);
or U256 (N_256,In_301,In_578);
and U257 (N_257,In_979,In_724);
or U258 (N_258,In_688,In_406);
nor U259 (N_259,In_501,In_376);
or U260 (N_260,In_303,In_128);
nand U261 (N_261,In_960,In_27);
or U262 (N_262,In_193,In_75);
nand U263 (N_263,In_337,In_367);
xor U264 (N_264,In_723,In_86);
and U265 (N_265,In_491,In_308);
nand U266 (N_266,In_970,In_888);
or U267 (N_267,In_328,In_127);
nand U268 (N_268,In_138,In_340);
and U269 (N_269,In_969,In_72);
and U270 (N_270,In_911,In_197);
xor U271 (N_271,In_690,In_485);
xor U272 (N_272,In_935,In_493);
or U273 (N_273,In_966,In_384);
nand U274 (N_274,In_608,In_237);
nand U275 (N_275,In_54,In_839);
and U276 (N_276,In_382,In_902);
xnor U277 (N_277,In_167,In_225);
and U278 (N_278,In_817,In_338);
and U279 (N_279,In_30,In_52);
or U280 (N_280,In_133,In_350);
nand U281 (N_281,In_326,In_269);
or U282 (N_282,In_711,In_317);
xnor U283 (N_283,In_143,In_434);
or U284 (N_284,In_928,In_850);
and U285 (N_285,In_61,In_670);
nand U286 (N_286,In_958,In_510);
and U287 (N_287,In_568,In_783);
or U288 (N_288,In_358,In_207);
nand U289 (N_289,In_620,In_596);
xor U290 (N_290,In_190,In_602);
nor U291 (N_291,In_913,In_300);
or U292 (N_292,In_684,In_583);
nor U293 (N_293,In_686,In_8);
and U294 (N_294,In_260,In_344);
nand U295 (N_295,In_479,In_731);
or U296 (N_296,In_396,In_609);
or U297 (N_297,In_118,In_994);
and U298 (N_298,In_428,In_552);
nand U299 (N_299,In_223,In_629);
xor U300 (N_300,In_663,In_456);
nor U301 (N_301,In_563,In_463);
nor U302 (N_302,In_241,In_727);
and U303 (N_303,In_24,In_689);
and U304 (N_304,In_859,In_775);
or U305 (N_305,In_354,In_244);
nand U306 (N_306,In_555,In_19);
and U307 (N_307,In_657,In_956);
and U308 (N_308,In_912,In_171);
and U309 (N_309,In_198,In_560);
and U310 (N_310,In_648,In_790);
nor U311 (N_311,In_566,In_773);
nand U312 (N_312,In_635,In_126);
or U313 (N_313,In_586,In_637);
nor U314 (N_314,In_470,In_436);
nor U315 (N_315,In_766,In_745);
or U316 (N_316,In_345,In_124);
nor U317 (N_317,In_247,In_806);
or U318 (N_318,In_798,In_142);
or U319 (N_319,In_38,In_746);
nor U320 (N_320,In_88,In_791);
and U321 (N_321,In_530,In_442);
or U322 (N_322,In_819,In_827);
or U323 (N_323,In_257,In_699);
nand U324 (N_324,In_401,In_618);
nor U325 (N_325,In_889,In_431);
nand U326 (N_326,In_644,In_831);
nand U327 (N_327,In_884,In_669);
or U328 (N_328,In_996,In_738);
xnor U329 (N_329,In_77,In_588);
nor U330 (N_330,In_537,In_794);
xnor U331 (N_331,In_509,In_63);
and U332 (N_332,In_278,In_938);
and U333 (N_333,In_708,In_286);
or U334 (N_334,In_267,In_658);
nor U335 (N_335,In_661,In_40);
xnor U336 (N_336,In_615,In_205);
and U337 (N_337,In_898,In_719);
nand U338 (N_338,In_1,In_870);
or U339 (N_339,In_346,In_599);
and U340 (N_340,In_117,In_330);
and U341 (N_341,In_192,In_606);
nand U342 (N_342,In_242,In_104);
or U343 (N_343,In_591,In_377);
nand U344 (N_344,In_624,In_274);
nand U345 (N_345,In_959,In_320);
or U346 (N_346,In_787,In_777);
nand U347 (N_347,In_336,In_186);
nand U348 (N_348,In_747,In_106);
or U349 (N_349,In_858,In_965);
nand U350 (N_350,In_412,In_204);
and U351 (N_351,In_107,In_415);
xnor U352 (N_352,In_924,In_675);
nor U353 (N_353,In_975,In_304);
xor U354 (N_354,In_299,In_196);
nor U355 (N_355,In_722,In_557);
xor U356 (N_356,In_729,In_80);
nand U357 (N_357,In_604,In_270);
or U358 (N_358,In_755,In_674);
nand U359 (N_359,In_135,In_489);
or U360 (N_360,In_380,In_319);
and U361 (N_361,In_349,In_678);
and U362 (N_362,In_985,In_287);
nand U363 (N_363,In_136,In_513);
and U364 (N_364,In_520,In_130);
and U365 (N_365,In_173,In_877);
nand U366 (N_366,In_459,In_372);
nor U367 (N_367,In_288,In_577);
and U368 (N_368,In_579,In_159);
and U369 (N_369,In_219,In_757);
nor U370 (N_370,In_137,In_400);
or U371 (N_371,In_772,In_419);
or U372 (N_372,In_115,In_87);
nor U373 (N_373,In_446,In_174);
nor U374 (N_374,In_447,In_416);
and U375 (N_375,In_455,In_939);
and U376 (N_376,In_427,In_112);
or U377 (N_377,In_952,In_547);
or U378 (N_378,In_906,In_735);
or U379 (N_379,In_249,In_453);
and U380 (N_380,In_874,In_108);
and U381 (N_381,In_875,In_730);
and U382 (N_382,In_630,In_194);
or U383 (N_383,In_559,In_517);
xnor U384 (N_384,In_362,In_305);
and U385 (N_385,In_352,In_803);
and U386 (N_386,In_2,In_523);
and U387 (N_387,In_584,In_181);
or U388 (N_388,In_392,In_397);
and U389 (N_389,In_810,In_751);
nand U390 (N_390,In_424,In_93);
or U391 (N_391,In_222,In_962);
and U392 (N_392,In_432,In_551);
and U393 (N_393,In_473,In_573);
and U394 (N_394,In_632,In_797);
nor U395 (N_395,In_829,In_511);
and U396 (N_396,In_716,In_45);
nand U397 (N_397,In_422,In_834);
nand U398 (N_398,In_191,In_444);
xor U399 (N_399,In_341,In_923);
and U400 (N_400,In_100,In_189);
nor U401 (N_401,In_739,In_543);
or U402 (N_402,In_836,In_240);
nand U403 (N_403,In_743,In_285);
nor U404 (N_404,In_230,In_564);
and U405 (N_405,In_901,In_828);
nand U406 (N_406,In_767,In_548);
nand U407 (N_407,In_368,In_891);
or U408 (N_408,In_46,In_25);
and U409 (N_409,In_841,In_421);
nor U410 (N_410,In_109,In_641);
and U411 (N_411,In_904,In_528);
nand U412 (N_412,In_672,In_792);
or U413 (N_413,In_506,In_258);
and U414 (N_414,In_48,In_271);
and U415 (N_415,In_844,In_587);
nor U416 (N_416,In_238,In_233);
nor U417 (N_417,In_67,In_220);
nor U418 (N_418,In_499,In_187);
nand U419 (N_419,In_879,In_703);
or U420 (N_420,In_451,In_62);
and U421 (N_421,In_522,In_235);
or U422 (N_422,In_683,In_656);
nor U423 (N_423,In_971,In_809);
nand U424 (N_424,In_203,In_890);
nor U425 (N_425,In_15,In_487);
nor U426 (N_426,In_356,In_702);
nor U427 (N_427,In_562,In_646);
xor U428 (N_428,In_256,In_21);
or U429 (N_429,In_229,In_737);
nor U430 (N_430,In_114,In_712);
or U431 (N_431,In_440,In_835);
or U432 (N_432,In_226,In_659);
nand U433 (N_433,In_585,In_709);
nor U434 (N_434,In_68,In_647);
nand U435 (N_435,In_293,In_732);
or U436 (N_436,In_363,In_617);
and U437 (N_437,In_163,In_818);
nor U438 (N_438,In_974,In_832);
nand U439 (N_439,In_695,In_851);
nand U440 (N_440,In_845,In_651);
nor U441 (N_441,In_849,In_402);
nand U442 (N_442,In_37,In_417);
xnor U443 (N_443,In_292,In_949);
xnor U444 (N_444,In_466,In_921);
and U445 (N_445,In_36,In_628);
nor U446 (N_446,In_69,In_164);
nor U447 (N_447,In_728,In_210);
nand U448 (N_448,In_50,In_121);
nor U449 (N_449,In_14,In_603);
and U450 (N_450,In_600,In_55);
or U451 (N_451,In_252,In_512);
nor U452 (N_452,In_860,In_549);
nand U453 (N_453,In_254,In_558);
nand U454 (N_454,In_281,In_519);
and U455 (N_455,In_565,In_993);
nor U456 (N_456,In_404,In_897);
nand U457 (N_457,In_140,In_6);
nor U458 (N_458,In_306,In_423);
nor U459 (N_459,In_718,In_231);
nor U460 (N_460,In_211,In_758);
or U461 (N_461,In_769,In_388);
and U462 (N_462,In_461,In_516);
and U463 (N_463,In_435,In_185);
and U464 (N_464,In_852,In_725);
nor U465 (N_465,In_393,In_51);
and U466 (N_466,In_785,In_334);
or U467 (N_467,In_931,In_369);
nand U468 (N_468,In_165,In_33);
nand U469 (N_469,In_622,In_526);
and U470 (N_470,In_332,In_125);
xnor U471 (N_471,In_825,In_5);
nor U472 (N_472,In_886,In_914);
nor U473 (N_473,In_977,In_476);
nor U474 (N_474,In_312,In_280);
xor U475 (N_475,In_283,In_926);
or U476 (N_476,In_922,In_753);
xnor U477 (N_477,In_43,In_910);
nand U478 (N_478,In_81,In_0);
nor U479 (N_479,In_153,In_391);
nand U480 (N_480,In_687,In_892);
or U481 (N_481,In_430,In_457);
and U482 (N_482,In_132,In_754);
nand U483 (N_483,In_145,In_276);
nand U484 (N_484,In_942,In_983);
and U485 (N_485,In_594,In_900);
xor U486 (N_486,In_917,In_486);
nor U487 (N_487,In_508,In_199);
nor U488 (N_488,In_150,In_762);
or U489 (N_489,In_445,In_481);
or U490 (N_490,In_176,In_714);
nor U491 (N_491,In_119,In_315);
and U492 (N_492,In_99,In_561);
nor U493 (N_493,In_880,In_89);
nand U494 (N_494,In_383,In_34);
xnor U495 (N_495,In_475,In_781);
nor U496 (N_496,In_951,In_95);
nand U497 (N_497,In_867,In_78);
nor U498 (N_498,In_59,In_386);
or U499 (N_499,In_323,In_571);
xnor U500 (N_500,In_420,In_949);
and U501 (N_501,In_631,In_970);
or U502 (N_502,In_218,In_666);
nand U503 (N_503,In_48,In_811);
and U504 (N_504,In_497,In_28);
nor U505 (N_505,In_164,In_684);
and U506 (N_506,In_246,In_668);
nand U507 (N_507,In_879,In_112);
or U508 (N_508,In_41,In_795);
nor U509 (N_509,In_437,In_448);
nand U510 (N_510,In_586,In_87);
and U511 (N_511,In_794,In_772);
and U512 (N_512,In_898,In_655);
and U513 (N_513,In_290,In_383);
or U514 (N_514,In_134,In_94);
nand U515 (N_515,In_63,In_604);
nand U516 (N_516,In_906,In_41);
nand U517 (N_517,In_597,In_448);
nor U518 (N_518,In_492,In_572);
nor U519 (N_519,In_805,In_128);
and U520 (N_520,In_399,In_927);
or U521 (N_521,In_243,In_204);
or U522 (N_522,In_179,In_206);
xnor U523 (N_523,In_917,In_513);
or U524 (N_524,In_628,In_897);
or U525 (N_525,In_374,In_507);
or U526 (N_526,In_498,In_386);
and U527 (N_527,In_559,In_388);
or U528 (N_528,In_901,In_696);
nand U529 (N_529,In_427,In_271);
nand U530 (N_530,In_299,In_508);
and U531 (N_531,In_819,In_762);
nand U532 (N_532,In_455,In_240);
and U533 (N_533,In_55,In_674);
and U534 (N_534,In_329,In_759);
nor U535 (N_535,In_684,In_815);
or U536 (N_536,In_798,In_466);
and U537 (N_537,In_259,In_467);
nor U538 (N_538,In_95,In_862);
or U539 (N_539,In_779,In_311);
xnor U540 (N_540,In_512,In_394);
and U541 (N_541,In_116,In_446);
nor U542 (N_542,In_834,In_22);
or U543 (N_543,In_269,In_68);
nor U544 (N_544,In_973,In_380);
and U545 (N_545,In_836,In_114);
and U546 (N_546,In_386,In_888);
and U547 (N_547,In_960,In_389);
nand U548 (N_548,In_395,In_358);
and U549 (N_549,In_482,In_991);
and U550 (N_550,In_242,In_241);
nand U551 (N_551,In_235,In_247);
and U552 (N_552,In_179,In_239);
and U553 (N_553,In_344,In_958);
xor U554 (N_554,In_992,In_297);
nand U555 (N_555,In_584,In_292);
or U556 (N_556,In_215,In_660);
nor U557 (N_557,In_894,In_423);
nand U558 (N_558,In_238,In_591);
and U559 (N_559,In_130,In_790);
nor U560 (N_560,In_752,In_447);
nor U561 (N_561,In_321,In_174);
nand U562 (N_562,In_855,In_477);
nand U563 (N_563,In_902,In_794);
xnor U564 (N_564,In_158,In_657);
or U565 (N_565,In_876,In_584);
or U566 (N_566,In_932,In_294);
xnor U567 (N_567,In_222,In_617);
nor U568 (N_568,In_896,In_47);
nor U569 (N_569,In_125,In_452);
xor U570 (N_570,In_168,In_510);
and U571 (N_571,In_414,In_907);
and U572 (N_572,In_392,In_765);
or U573 (N_573,In_632,In_10);
or U574 (N_574,In_469,In_37);
or U575 (N_575,In_438,In_336);
and U576 (N_576,In_649,In_227);
or U577 (N_577,In_512,In_513);
or U578 (N_578,In_113,In_784);
and U579 (N_579,In_905,In_444);
nand U580 (N_580,In_846,In_654);
or U581 (N_581,In_816,In_703);
xor U582 (N_582,In_764,In_788);
and U583 (N_583,In_749,In_199);
nand U584 (N_584,In_591,In_754);
nor U585 (N_585,In_157,In_309);
and U586 (N_586,In_617,In_773);
and U587 (N_587,In_759,In_841);
and U588 (N_588,In_145,In_859);
xor U589 (N_589,In_432,In_988);
or U590 (N_590,In_608,In_27);
or U591 (N_591,In_934,In_756);
and U592 (N_592,In_471,In_210);
nand U593 (N_593,In_268,In_392);
nor U594 (N_594,In_300,In_593);
and U595 (N_595,In_606,In_345);
nand U596 (N_596,In_104,In_447);
nand U597 (N_597,In_228,In_459);
or U598 (N_598,In_898,In_309);
nand U599 (N_599,In_424,In_248);
nor U600 (N_600,In_643,In_642);
xnor U601 (N_601,In_331,In_55);
and U602 (N_602,In_226,In_597);
nor U603 (N_603,In_828,In_722);
nand U604 (N_604,In_146,In_571);
or U605 (N_605,In_817,In_800);
and U606 (N_606,In_364,In_510);
nor U607 (N_607,In_315,In_120);
and U608 (N_608,In_447,In_280);
xnor U609 (N_609,In_905,In_580);
and U610 (N_610,In_967,In_226);
xor U611 (N_611,In_419,In_470);
nor U612 (N_612,In_197,In_878);
nor U613 (N_613,In_765,In_275);
nor U614 (N_614,In_37,In_575);
nand U615 (N_615,In_68,In_651);
nor U616 (N_616,In_146,In_448);
and U617 (N_617,In_417,In_300);
nor U618 (N_618,In_556,In_922);
and U619 (N_619,In_833,In_665);
or U620 (N_620,In_43,In_668);
and U621 (N_621,In_998,In_549);
and U622 (N_622,In_941,In_131);
or U623 (N_623,In_965,In_783);
or U624 (N_624,In_877,In_962);
or U625 (N_625,In_270,In_713);
nor U626 (N_626,In_867,In_938);
xor U627 (N_627,In_613,In_702);
nand U628 (N_628,In_114,In_496);
or U629 (N_629,In_333,In_762);
and U630 (N_630,In_588,In_329);
or U631 (N_631,In_228,In_902);
nor U632 (N_632,In_659,In_474);
nor U633 (N_633,In_397,In_126);
nor U634 (N_634,In_249,In_854);
nand U635 (N_635,In_565,In_358);
and U636 (N_636,In_440,In_410);
nor U637 (N_637,In_130,In_328);
nor U638 (N_638,In_137,In_628);
nor U639 (N_639,In_540,In_808);
xnor U640 (N_640,In_712,In_108);
or U641 (N_641,In_727,In_918);
nand U642 (N_642,In_98,In_461);
and U643 (N_643,In_266,In_385);
and U644 (N_644,In_540,In_50);
nor U645 (N_645,In_799,In_82);
or U646 (N_646,In_833,In_789);
xor U647 (N_647,In_248,In_492);
nor U648 (N_648,In_983,In_250);
nor U649 (N_649,In_833,In_878);
and U650 (N_650,In_491,In_109);
nor U651 (N_651,In_471,In_232);
nand U652 (N_652,In_681,In_62);
and U653 (N_653,In_731,In_391);
nand U654 (N_654,In_217,In_414);
and U655 (N_655,In_884,In_183);
and U656 (N_656,In_603,In_372);
xnor U657 (N_657,In_742,In_85);
nand U658 (N_658,In_679,In_486);
nand U659 (N_659,In_310,In_750);
or U660 (N_660,In_89,In_10);
nand U661 (N_661,In_2,In_585);
or U662 (N_662,In_748,In_658);
xnor U663 (N_663,In_116,In_495);
nand U664 (N_664,In_91,In_970);
or U665 (N_665,In_523,In_271);
nor U666 (N_666,In_441,In_2);
xor U667 (N_667,In_715,In_378);
nand U668 (N_668,In_492,In_569);
or U669 (N_669,In_907,In_988);
nand U670 (N_670,In_276,In_959);
nand U671 (N_671,In_761,In_173);
xor U672 (N_672,In_813,In_355);
nor U673 (N_673,In_731,In_663);
nand U674 (N_674,In_841,In_579);
and U675 (N_675,In_18,In_169);
nand U676 (N_676,In_172,In_283);
xnor U677 (N_677,In_311,In_699);
or U678 (N_678,In_263,In_316);
nor U679 (N_679,In_179,In_352);
or U680 (N_680,In_831,In_462);
or U681 (N_681,In_970,In_66);
or U682 (N_682,In_594,In_829);
nand U683 (N_683,In_138,In_613);
and U684 (N_684,In_743,In_170);
nor U685 (N_685,In_757,In_510);
and U686 (N_686,In_496,In_402);
and U687 (N_687,In_116,In_630);
nand U688 (N_688,In_115,In_240);
nor U689 (N_689,In_786,In_538);
xnor U690 (N_690,In_247,In_791);
nand U691 (N_691,In_182,In_732);
nor U692 (N_692,In_115,In_258);
nand U693 (N_693,In_354,In_724);
or U694 (N_694,In_852,In_117);
or U695 (N_695,In_477,In_23);
and U696 (N_696,In_188,In_114);
xnor U697 (N_697,In_481,In_334);
xnor U698 (N_698,In_423,In_544);
and U699 (N_699,In_419,In_23);
nor U700 (N_700,In_201,In_696);
and U701 (N_701,In_616,In_128);
and U702 (N_702,In_895,In_774);
xnor U703 (N_703,In_80,In_454);
nor U704 (N_704,In_422,In_613);
or U705 (N_705,In_814,In_680);
xnor U706 (N_706,In_859,In_605);
nor U707 (N_707,In_498,In_333);
or U708 (N_708,In_39,In_44);
nand U709 (N_709,In_246,In_9);
nand U710 (N_710,In_329,In_28);
xor U711 (N_711,In_246,In_482);
nor U712 (N_712,In_352,In_883);
and U713 (N_713,In_21,In_226);
nand U714 (N_714,In_472,In_833);
nand U715 (N_715,In_382,In_624);
nand U716 (N_716,In_571,In_276);
and U717 (N_717,In_942,In_901);
nor U718 (N_718,In_471,In_885);
nor U719 (N_719,In_870,In_884);
nor U720 (N_720,In_8,In_774);
and U721 (N_721,In_436,In_742);
nor U722 (N_722,In_683,In_822);
xor U723 (N_723,In_225,In_873);
and U724 (N_724,In_904,In_73);
nand U725 (N_725,In_298,In_549);
or U726 (N_726,In_217,In_754);
and U727 (N_727,In_885,In_759);
nor U728 (N_728,In_670,In_835);
nor U729 (N_729,In_501,In_225);
nand U730 (N_730,In_376,In_670);
and U731 (N_731,In_33,In_24);
nand U732 (N_732,In_167,In_195);
or U733 (N_733,In_593,In_354);
nor U734 (N_734,In_210,In_794);
nand U735 (N_735,In_769,In_287);
nand U736 (N_736,In_807,In_698);
nand U737 (N_737,In_814,In_975);
and U738 (N_738,In_109,In_729);
or U739 (N_739,In_833,In_581);
and U740 (N_740,In_172,In_314);
or U741 (N_741,In_217,In_775);
nor U742 (N_742,In_821,In_648);
xor U743 (N_743,In_87,In_934);
and U744 (N_744,In_732,In_659);
and U745 (N_745,In_530,In_118);
and U746 (N_746,In_951,In_165);
or U747 (N_747,In_940,In_684);
xnor U748 (N_748,In_837,In_673);
nand U749 (N_749,In_614,In_649);
and U750 (N_750,In_739,In_221);
nand U751 (N_751,In_231,In_253);
nor U752 (N_752,In_906,In_16);
nand U753 (N_753,In_867,In_765);
xor U754 (N_754,In_154,In_488);
nand U755 (N_755,In_180,In_9);
xnor U756 (N_756,In_468,In_252);
nand U757 (N_757,In_21,In_584);
or U758 (N_758,In_404,In_137);
or U759 (N_759,In_917,In_99);
and U760 (N_760,In_939,In_896);
nand U761 (N_761,In_141,In_771);
nand U762 (N_762,In_536,In_535);
or U763 (N_763,In_452,In_687);
xor U764 (N_764,In_653,In_449);
or U765 (N_765,In_721,In_508);
nor U766 (N_766,In_781,In_393);
xnor U767 (N_767,In_140,In_388);
and U768 (N_768,In_815,In_410);
nand U769 (N_769,In_424,In_186);
or U770 (N_770,In_771,In_110);
nand U771 (N_771,In_492,In_942);
nand U772 (N_772,In_535,In_441);
nand U773 (N_773,In_303,In_475);
xor U774 (N_774,In_867,In_806);
or U775 (N_775,In_227,In_682);
and U776 (N_776,In_355,In_102);
or U777 (N_777,In_790,In_675);
or U778 (N_778,In_436,In_632);
or U779 (N_779,In_156,In_697);
nand U780 (N_780,In_907,In_31);
and U781 (N_781,In_557,In_736);
and U782 (N_782,In_12,In_755);
and U783 (N_783,In_255,In_349);
and U784 (N_784,In_856,In_211);
nand U785 (N_785,In_268,In_74);
or U786 (N_786,In_940,In_273);
nor U787 (N_787,In_812,In_892);
nor U788 (N_788,In_816,In_304);
nor U789 (N_789,In_657,In_76);
nand U790 (N_790,In_939,In_32);
or U791 (N_791,In_636,In_82);
nor U792 (N_792,In_417,In_862);
nor U793 (N_793,In_307,In_528);
or U794 (N_794,In_280,In_370);
or U795 (N_795,In_49,In_443);
xnor U796 (N_796,In_622,In_10);
xor U797 (N_797,In_709,In_739);
nor U798 (N_798,In_174,In_102);
or U799 (N_799,In_743,In_983);
nand U800 (N_800,In_922,In_564);
nor U801 (N_801,In_589,In_269);
and U802 (N_802,In_482,In_447);
or U803 (N_803,In_810,In_12);
or U804 (N_804,In_537,In_570);
nand U805 (N_805,In_254,In_526);
xor U806 (N_806,In_246,In_568);
nor U807 (N_807,In_882,In_836);
nand U808 (N_808,In_34,In_936);
and U809 (N_809,In_852,In_652);
nor U810 (N_810,In_189,In_226);
nand U811 (N_811,In_306,In_853);
nor U812 (N_812,In_476,In_465);
nand U813 (N_813,In_147,In_994);
nor U814 (N_814,In_30,In_957);
or U815 (N_815,In_476,In_7);
nor U816 (N_816,In_703,In_819);
and U817 (N_817,In_807,In_656);
nand U818 (N_818,In_513,In_361);
nor U819 (N_819,In_11,In_323);
and U820 (N_820,In_928,In_292);
and U821 (N_821,In_580,In_39);
xnor U822 (N_822,In_760,In_454);
nand U823 (N_823,In_410,In_507);
or U824 (N_824,In_610,In_563);
nor U825 (N_825,In_145,In_195);
nor U826 (N_826,In_681,In_370);
or U827 (N_827,In_559,In_949);
nor U828 (N_828,In_647,In_762);
nand U829 (N_829,In_987,In_558);
and U830 (N_830,In_895,In_496);
and U831 (N_831,In_921,In_993);
nor U832 (N_832,In_537,In_441);
nor U833 (N_833,In_756,In_548);
xnor U834 (N_834,In_855,In_634);
or U835 (N_835,In_907,In_980);
xnor U836 (N_836,In_349,In_623);
xor U837 (N_837,In_612,In_686);
or U838 (N_838,In_1,In_229);
and U839 (N_839,In_626,In_38);
or U840 (N_840,In_138,In_120);
and U841 (N_841,In_759,In_623);
nor U842 (N_842,In_515,In_475);
and U843 (N_843,In_137,In_533);
or U844 (N_844,In_270,In_478);
xor U845 (N_845,In_67,In_500);
nor U846 (N_846,In_940,In_756);
nand U847 (N_847,In_985,In_233);
or U848 (N_848,In_325,In_385);
and U849 (N_849,In_419,In_369);
nand U850 (N_850,In_958,In_246);
or U851 (N_851,In_649,In_925);
and U852 (N_852,In_215,In_849);
nand U853 (N_853,In_783,In_708);
nand U854 (N_854,In_77,In_678);
and U855 (N_855,In_252,In_763);
nand U856 (N_856,In_600,In_338);
nor U857 (N_857,In_334,In_217);
nand U858 (N_858,In_561,In_957);
nand U859 (N_859,In_707,In_986);
or U860 (N_860,In_266,In_48);
nand U861 (N_861,In_356,In_3);
nor U862 (N_862,In_423,In_602);
nor U863 (N_863,In_567,In_67);
or U864 (N_864,In_877,In_482);
and U865 (N_865,In_757,In_742);
nand U866 (N_866,In_178,In_88);
or U867 (N_867,In_813,In_843);
xnor U868 (N_868,In_567,In_303);
nand U869 (N_869,In_714,In_547);
nand U870 (N_870,In_722,In_614);
xor U871 (N_871,In_490,In_49);
nand U872 (N_872,In_358,In_114);
xor U873 (N_873,In_986,In_283);
or U874 (N_874,In_136,In_524);
nor U875 (N_875,In_263,In_159);
nor U876 (N_876,In_734,In_753);
nor U877 (N_877,In_543,In_224);
and U878 (N_878,In_93,In_915);
and U879 (N_879,In_98,In_543);
or U880 (N_880,In_172,In_322);
nor U881 (N_881,In_919,In_662);
or U882 (N_882,In_717,In_423);
or U883 (N_883,In_779,In_425);
or U884 (N_884,In_225,In_484);
xor U885 (N_885,In_974,In_435);
nor U886 (N_886,In_993,In_202);
nor U887 (N_887,In_656,In_965);
or U888 (N_888,In_725,In_763);
xor U889 (N_889,In_857,In_148);
nor U890 (N_890,In_967,In_297);
or U891 (N_891,In_114,In_206);
nand U892 (N_892,In_716,In_235);
and U893 (N_893,In_484,In_170);
nand U894 (N_894,In_393,In_683);
nand U895 (N_895,In_413,In_182);
xnor U896 (N_896,In_824,In_467);
xor U897 (N_897,In_19,In_536);
nand U898 (N_898,In_816,In_189);
and U899 (N_899,In_711,In_475);
or U900 (N_900,In_488,In_192);
or U901 (N_901,In_616,In_365);
nand U902 (N_902,In_781,In_539);
nand U903 (N_903,In_751,In_718);
nand U904 (N_904,In_578,In_562);
nand U905 (N_905,In_171,In_474);
nand U906 (N_906,In_349,In_888);
or U907 (N_907,In_462,In_458);
or U908 (N_908,In_145,In_438);
nand U909 (N_909,In_986,In_12);
nor U910 (N_910,In_338,In_512);
nor U911 (N_911,In_475,In_652);
xor U912 (N_912,In_862,In_74);
nor U913 (N_913,In_480,In_622);
nor U914 (N_914,In_221,In_952);
nor U915 (N_915,In_403,In_90);
nand U916 (N_916,In_694,In_997);
xor U917 (N_917,In_6,In_191);
or U918 (N_918,In_474,In_511);
nor U919 (N_919,In_555,In_876);
nor U920 (N_920,In_44,In_52);
nand U921 (N_921,In_577,In_448);
and U922 (N_922,In_182,In_335);
nor U923 (N_923,In_796,In_894);
nand U924 (N_924,In_680,In_340);
xor U925 (N_925,In_789,In_466);
xor U926 (N_926,In_249,In_263);
and U927 (N_927,In_756,In_54);
nand U928 (N_928,In_599,In_916);
or U929 (N_929,In_624,In_976);
nand U930 (N_930,In_281,In_399);
xnor U931 (N_931,In_922,In_570);
and U932 (N_932,In_871,In_345);
and U933 (N_933,In_506,In_48);
or U934 (N_934,In_987,In_415);
nor U935 (N_935,In_708,In_561);
nand U936 (N_936,In_229,In_220);
and U937 (N_937,In_276,In_404);
or U938 (N_938,In_783,In_578);
or U939 (N_939,In_294,In_218);
or U940 (N_940,In_511,In_358);
nor U941 (N_941,In_486,In_841);
nor U942 (N_942,In_382,In_914);
nor U943 (N_943,In_301,In_457);
nand U944 (N_944,In_782,In_712);
or U945 (N_945,In_763,In_656);
or U946 (N_946,In_495,In_552);
or U947 (N_947,In_569,In_339);
nand U948 (N_948,In_663,In_655);
and U949 (N_949,In_976,In_441);
or U950 (N_950,In_745,In_978);
nor U951 (N_951,In_653,In_610);
or U952 (N_952,In_497,In_52);
nor U953 (N_953,In_277,In_92);
and U954 (N_954,In_765,In_284);
and U955 (N_955,In_962,In_400);
and U956 (N_956,In_388,In_893);
or U957 (N_957,In_935,In_288);
or U958 (N_958,In_273,In_724);
xor U959 (N_959,In_717,In_852);
nand U960 (N_960,In_326,In_607);
nand U961 (N_961,In_279,In_162);
nand U962 (N_962,In_455,In_743);
nor U963 (N_963,In_785,In_12);
nor U964 (N_964,In_725,In_250);
nand U965 (N_965,In_687,In_11);
and U966 (N_966,In_518,In_810);
or U967 (N_967,In_231,In_678);
or U968 (N_968,In_757,In_45);
nor U969 (N_969,In_225,In_664);
or U970 (N_970,In_700,In_281);
or U971 (N_971,In_14,In_436);
nor U972 (N_972,In_592,In_591);
xnor U973 (N_973,In_419,In_709);
xor U974 (N_974,In_970,In_454);
nand U975 (N_975,In_285,In_360);
nand U976 (N_976,In_283,In_256);
nand U977 (N_977,In_958,In_336);
nor U978 (N_978,In_785,In_70);
nand U979 (N_979,In_583,In_644);
nor U980 (N_980,In_916,In_153);
and U981 (N_981,In_526,In_173);
or U982 (N_982,In_782,In_827);
xor U983 (N_983,In_91,In_260);
nor U984 (N_984,In_305,In_855);
nand U985 (N_985,In_343,In_348);
nand U986 (N_986,In_912,In_299);
or U987 (N_987,In_927,In_817);
xnor U988 (N_988,In_445,In_568);
or U989 (N_989,In_446,In_946);
or U990 (N_990,In_605,In_648);
and U991 (N_991,In_938,In_711);
and U992 (N_992,In_656,In_373);
and U993 (N_993,In_516,In_546);
xor U994 (N_994,In_938,In_163);
xor U995 (N_995,In_213,In_446);
nor U996 (N_996,In_592,In_378);
or U997 (N_997,In_857,In_885);
nand U998 (N_998,In_664,In_790);
or U999 (N_999,In_582,In_748);
and U1000 (N_1000,N_569,N_576);
nor U1001 (N_1001,N_260,N_298);
nor U1002 (N_1002,N_751,N_51);
or U1003 (N_1003,N_623,N_18);
nor U1004 (N_1004,N_291,N_13);
nor U1005 (N_1005,N_80,N_747);
or U1006 (N_1006,N_114,N_335);
nand U1007 (N_1007,N_840,N_495);
or U1008 (N_1008,N_437,N_804);
xnor U1009 (N_1009,N_993,N_476);
nor U1010 (N_1010,N_121,N_313);
or U1011 (N_1011,N_488,N_616);
nand U1012 (N_1012,N_17,N_978);
nor U1013 (N_1013,N_737,N_195);
nor U1014 (N_1014,N_416,N_898);
nand U1015 (N_1015,N_585,N_824);
or U1016 (N_1016,N_969,N_778);
nand U1017 (N_1017,N_829,N_679);
nand U1018 (N_1018,N_149,N_656);
nand U1019 (N_1019,N_825,N_442);
or U1020 (N_1020,N_590,N_65);
nor U1021 (N_1021,N_815,N_746);
or U1022 (N_1022,N_877,N_923);
nor U1023 (N_1023,N_699,N_67);
nand U1024 (N_1024,N_161,N_721);
nand U1025 (N_1025,N_521,N_54);
nand U1026 (N_1026,N_300,N_181);
nand U1027 (N_1027,N_944,N_283);
nor U1028 (N_1028,N_199,N_591);
or U1029 (N_1029,N_246,N_318);
or U1030 (N_1030,N_535,N_608);
and U1031 (N_1031,N_96,N_409);
nor U1032 (N_1032,N_723,N_431);
nand U1033 (N_1033,N_704,N_117);
nor U1034 (N_1034,N_701,N_878);
or U1035 (N_1035,N_542,N_166);
nor U1036 (N_1036,N_487,N_578);
xor U1037 (N_1037,N_302,N_839);
nor U1038 (N_1038,N_631,N_558);
or U1039 (N_1039,N_113,N_726);
nor U1040 (N_1040,N_243,N_438);
nor U1041 (N_1041,N_189,N_383);
and U1042 (N_1042,N_727,N_802);
nor U1043 (N_1043,N_629,N_424);
or U1044 (N_1044,N_491,N_584);
and U1045 (N_1045,N_617,N_69);
or U1046 (N_1046,N_299,N_418);
xnor U1047 (N_1047,N_380,N_456);
nand U1048 (N_1048,N_84,N_970);
and U1049 (N_1049,N_885,N_915);
or U1050 (N_1050,N_996,N_141);
and U1051 (N_1051,N_465,N_962);
nand U1052 (N_1052,N_359,N_439);
nand U1053 (N_1053,N_444,N_647);
or U1054 (N_1054,N_344,N_637);
and U1055 (N_1055,N_242,N_965);
and U1056 (N_1056,N_889,N_393);
xnor U1057 (N_1057,N_44,N_512);
and U1058 (N_1058,N_781,N_796);
and U1059 (N_1059,N_486,N_78);
xor U1060 (N_1060,N_435,N_163);
nor U1061 (N_1061,N_93,N_694);
xor U1062 (N_1062,N_12,N_817);
nand U1063 (N_1063,N_618,N_866);
or U1064 (N_1064,N_66,N_29);
and U1065 (N_1065,N_441,N_508);
or U1066 (N_1066,N_959,N_333);
nand U1067 (N_1067,N_734,N_417);
or U1068 (N_1068,N_180,N_296);
nor U1069 (N_1069,N_575,N_198);
and U1070 (N_1070,N_32,N_167);
and U1071 (N_1071,N_919,N_743);
and U1072 (N_1072,N_951,N_543);
nand U1073 (N_1073,N_914,N_7);
nand U1074 (N_1074,N_317,N_365);
nor U1075 (N_1075,N_589,N_844);
and U1076 (N_1076,N_150,N_190);
and U1077 (N_1077,N_605,N_232);
nand U1078 (N_1078,N_641,N_523);
nand U1079 (N_1079,N_626,N_554);
nor U1080 (N_1080,N_251,N_819);
nand U1081 (N_1081,N_258,N_660);
and U1082 (N_1082,N_640,N_279);
or U1083 (N_1083,N_767,N_207);
xnor U1084 (N_1084,N_500,N_579);
or U1085 (N_1085,N_800,N_570);
or U1086 (N_1086,N_853,N_38);
xor U1087 (N_1087,N_902,N_686);
nor U1088 (N_1088,N_322,N_942);
nand U1089 (N_1089,N_587,N_916);
nor U1090 (N_1090,N_156,N_133);
xor U1091 (N_1091,N_176,N_284);
nor U1092 (N_1092,N_42,N_267);
or U1093 (N_1093,N_130,N_971);
or U1094 (N_1094,N_261,N_813);
and U1095 (N_1095,N_688,N_857);
xor U1096 (N_1096,N_4,N_566);
and U1097 (N_1097,N_41,N_571);
or U1098 (N_1098,N_922,N_670);
nor U1099 (N_1099,N_337,N_323);
or U1100 (N_1100,N_655,N_528);
or U1101 (N_1101,N_135,N_593);
or U1102 (N_1102,N_832,N_35);
and U1103 (N_1103,N_875,N_275);
nand U1104 (N_1104,N_999,N_55);
and U1105 (N_1105,N_645,N_956);
or U1106 (N_1106,N_168,N_818);
nand U1107 (N_1107,N_596,N_854);
or U1108 (N_1108,N_794,N_861);
and U1109 (N_1109,N_384,N_10);
nand U1110 (N_1110,N_790,N_518);
xnor U1111 (N_1111,N_609,N_27);
nor U1112 (N_1112,N_343,N_805);
nand U1113 (N_1113,N_691,N_236);
nor U1114 (N_1114,N_293,N_458);
or U1115 (N_1115,N_351,N_77);
nor U1116 (N_1116,N_464,N_178);
and U1117 (N_1117,N_801,N_724);
xnor U1118 (N_1118,N_239,N_250);
nor U1119 (N_1119,N_797,N_597);
xor U1120 (N_1120,N_931,N_663);
and U1121 (N_1121,N_780,N_990);
nor U1122 (N_1122,N_803,N_428);
or U1123 (N_1123,N_108,N_184);
nor U1124 (N_1124,N_443,N_674);
or U1125 (N_1125,N_489,N_142);
nand U1126 (N_1126,N_930,N_912);
xor U1127 (N_1127,N_635,N_779);
nand U1128 (N_1128,N_511,N_515);
or U1129 (N_1129,N_667,N_179);
nor U1130 (N_1130,N_565,N_471);
and U1131 (N_1131,N_870,N_864);
and U1132 (N_1132,N_347,N_202);
nand U1133 (N_1133,N_371,N_685);
xor U1134 (N_1134,N_771,N_177);
nor U1135 (N_1135,N_810,N_661);
nand U1136 (N_1136,N_567,N_94);
nor U1137 (N_1137,N_692,N_639);
nand U1138 (N_1138,N_262,N_665);
or U1139 (N_1139,N_231,N_58);
and U1140 (N_1140,N_376,N_643);
nor U1141 (N_1141,N_497,N_935);
and U1142 (N_1142,N_925,N_937);
nor U1143 (N_1143,N_147,N_21);
nor U1144 (N_1144,N_182,N_315);
nor U1145 (N_1145,N_325,N_361);
nand U1146 (N_1146,N_599,N_287);
nor U1147 (N_1147,N_99,N_731);
and U1148 (N_1148,N_281,N_582);
and U1149 (N_1149,N_729,N_23);
nand U1150 (N_1150,N_501,N_34);
nor U1151 (N_1151,N_282,N_826);
and U1152 (N_1152,N_847,N_95);
and U1153 (N_1153,N_115,N_711);
nor U1154 (N_1154,N_920,N_217);
or U1155 (N_1155,N_713,N_364);
nor U1156 (N_1156,N_47,N_849);
nand U1157 (N_1157,N_550,N_764);
nor U1158 (N_1158,N_346,N_226);
or U1159 (N_1159,N_259,N_194);
or U1160 (N_1160,N_940,N_256);
nor U1161 (N_1161,N_382,N_900);
and U1162 (N_1162,N_532,N_205);
nand U1163 (N_1163,N_60,N_869);
nor U1164 (N_1164,N_845,N_473);
or U1165 (N_1165,N_307,N_388);
or U1166 (N_1166,N_681,N_59);
xor U1167 (N_1167,N_917,N_534);
and U1168 (N_1168,N_433,N_379);
or U1169 (N_1169,N_633,N_556);
or U1170 (N_1170,N_338,N_911);
or U1171 (N_1171,N_835,N_118);
and U1172 (N_1172,N_310,N_122);
and U1173 (N_1173,N_657,N_559);
and U1174 (N_1174,N_837,N_110);
nor U1175 (N_1175,N_183,N_560);
nor U1176 (N_1176,N_81,N_57);
nand U1177 (N_1177,N_200,N_973);
nor U1178 (N_1178,N_714,N_316);
nand U1179 (N_1179,N_929,N_498);
nand U1180 (N_1180,N_216,N_229);
nand U1181 (N_1181,N_682,N_607);
or U1182 (N_1182,N_328,N_469);
nor U1183 (N_1183,N_329,N_948);
and U1184 (N_1184,N_834,N_934);
and U1185 (N_1185,N_994,N_98);
nor U1186 (N_1186,N_109,N_522);
or U1187 (N_1187,N_451,N_429);
nand U1188 (N_1188,N_564,N_237);
nor U1189 (N_1189,N_127,N_943);
nor U1190 (N_1190,N_209,N_881);
nand U1191 (N_1191,N_519,N_288);
and U1192 (N_1192,N_630,N_274);
and U1193 (N_1193,N_967,N_327);
nor U1194 (N_1194,N_320,N_852);
or U1195 (N_1195,N_436,N_389);
and U1196 (N_1196,N_153,N_588);
nand U1197 (N_1197,N_319,N_462);
or U1198 (N_1198,N_123,N_785);
nor U1199 (N_1199,N_705,N_947);
nand U1200 (N_1200,N_624,N_25);
nor U1201 (N_1201,N_879,N_710);
and U1202 (N_1202,N_63,N_745);
nand U1203 (N_1203,N_809,N_192);
or U1204 (N_1204,N_601,N_610);
nor U1205 (N_1205,N_676,N_505);
xnor U1206 (N_1206,N_659,N_848);
nand U1207 (N_1207,N_358,N_646);
or U1208 (N_1208,N_827,N_24);
nor U1209 (N_1209,N_330,N_482);
xor U1210 (N_1210,N_841,N_241);
and U1211 (N_1211,N_203,N_414);
nor U1212 (N_1212,N_171,N_331);
nor U1213 (N_1213,N_614,N_953);
and U1214 (N_1214,N_286,N_808);
or U1215 (N_1215,N_452,N_391);
nor U1216 (N_1216,N_503,N_873);
nor U1217 (N_1217,N_613,N_273);
or U1218 (N_1218,N_398,N_212);
or U1219 (N_1219,N_964,N_353);
xor U1220 (N_1220,N_842,N_733);
and U1221 (N_1221,N_649,N_907);
and U1222 (N_1222,N_112,N_572);
nand U1223 (N_1223,N_87,N_594);
nor U1224 (N_1224,N_604,N_908);
and U1225 (N_1225,N_134,N_413);
nand U1226 (N_1226,N_230,N_472);
nor U1227 (N_1227,N_157,N_807);
and U1228 (N_1228,N_690,N_492);
nor U1229 (N_1229,N_107,N_933);
nand U1230 (N_1230,N_524,N_88);
nand U1231 (N_1231,N_650,N_129);
nand U1232 (N_1232,N_722,N_223);
and U1233 (N_1233,N_309,N_749);
nor U1234 (N_1234,N_901,N_463);
and U1235 (N_1235,N_769,N_897);
nand U1236 (N_1236,N_972,N_26);
and U1237 (N_1237,N_981,N_125);
nand U1238 (N_1238,N_762,N_197);
and U1239 (N_1239,N_401,N_882);
nor U1240 (N_1240,N_420,N_634);
and U1241 (N_1241,N_742,N_669);
or U1242 (N_1242,N_757,N_468);
or U1243 (N_1243,N_155,N_540);
and U1244 (N_1244,N_700,N_753);
nor U1245 (N_1245,N_759,N_628);
xnor U1246 (N_1246,N_245,N_369);
and U1247 (N_1247,N_111,N_326);
or U1248 (N_1248,N_151,N_886);
or U1249 (N_1249,N_11,N_867);
nor U1250 (N_1250,N_831,N_62);
nor U1251 (N_1251,N_290,N_777);
nor U1252 (N_1252,N_301,N_228);
xor U1253 (N_1253,N_461,N_666);
xnor U1254 (N_1254,N_132,N_531);
nand U1255 (N_1255,N_76,N_139);
and U1256 (N_1256,N_860,N_352);
and U1257 (N_1257,N_684,N_255);
and U1258 (N_1258,N_74,N_173);
nand U1259 (N_1259,N_40,N_49);
and U1260 (N_1260,N_828,N_516);
xnor U1261 (N_1261,N_741,N_636);
xor U1262 (N_1262,N_213,N_960);
xor U1263 (N_1263,N_280,N_402);
or U1264 (N_1264,N_502,N_677);
xor U1265 (N_1265,N_822,N_72);
nand U1266 (N_1266,N_22,N_884);
nand U1267 (N_1267,N_381,N_549);
xor U1268 (N_1268,N_339,N_368);
or U1269 (N_1269,N_865,N_955);
and U1270 (N_1270,N_977,N_477);
nor U1271 (N_1271,N_305,N_367);
nor U1272 (N_1272,N_968,N_986);
or U1273 (N_1273,N_483,N_568);
xnor U1274 (N_1274,N_159,N_545);
nor U1275 (N_1275,N_52,N_385);
and U1276 (N_1276,N_252,N_86);
nand U1277 (N_1277,N_784,N_906);
and U1278 (N_1278,N_975,N_308);
nand U1279 (N_1279,N_592,N_905);
nor U1280 (N_1280,N_621,N_375);
nor U1281 (N_1281,N_137,N_334);
or U1282 (N_1282,N_510,N_638);
and U1283 (N_1283,N_814,N_752);
nand U1284 (N_1284,N_625,N_939);
nor U1285 (N_1285,N_648,N_548);
nor U1286 (N_1286,N_580,N_750);
or U1287 (N_1287,N_174,N_479);
nor U1288 (N_1288,N_600,N_595);
nor U1289 (N_1289,N_90,N_448);
or U1290 (N_1290,N_921,N_404);
or U1291 (N_1291,N_101,N_119);
and U1292 (N_1292,N_756,N_356);
nor U1293 (N_1293,N_526,N_421);
and U1294 (N_1294,N_362,N_165);
nor U1295 (N_1295,N_294,N_454);
nand U1296 (N_1296,N_264,N_561);
and U1297 (N_1297,N_553,N_744);
nand U1298 (N_1298,N_128,N_53);
and U1299 (N_1299,N_14,N_434);
and U1300 (N_1300,N_210,N_793);
and U1301 (N_1301,N_405,N_683);
and U1302 (N_1302,N_843,N_514);
xor U1303 (N_1303,N_83,N_46);
nand U1304 (N_1304,N_235,N_82);
nand U1305 (N_1305,N_278,N_410);
nor U1306 (N_1306,N_1,N_186);
xor U1307 (N_1307,N_211,N_680);
nand U1308 (N_1308,N_427,N_855);
and U1309 (N_1309,N_982,N_868);
nor U1310 (N_1310,N_789,N_70);
nand U1311 (N_1311,N_430,N_664);
or U1312 (N_1312,N_775,N_673);
and U1313 (N_1313,N_952,N_85);
nand U1314 (N_1314,N_791,N_812);
and U1315 (N_1315,N_707,N_33);
xor U1316 (N_1316,N_606,N_152);
nand U1317 (N_1317,N_619,N_332);
xor U1318 (N_1318,N_792,N_728);
nor U1319 (N_1319,N_520,N_577);
xnor U1320 (N_1320,N_583,N_220);
nand U1321 (N_1321,N_709,N_222);
xor U1322 (N_1322,N_782,N_697);
and U1323 (N_1323,N_340,N_924);
nor U1324 (N_1324,N_941,N_838);
nand U1325 (N_1325,N_68,N_979);
nor U1326 (N_1326,N_718,N_696);
nor U1327 (N_1327,N_716,N_976);
or U1328 (N_1328,N_899,N_225);
or U1329 (N_1329,N_146,N_946);
and U1330 (N_1330,N_527,N_529);
or U1331 (N_1331,N_412,N_883);
or U1332 (N_1332,N_552,N_862);
nand U1333 (N_1333,N_268,N_811);
and U1334 (N_1334,N_45,N_467);
and U1335 (N_1335,N_995,N_103);
nor U1336 (N_1336,N_390,N_292);
and U1337 (N_1337,N_30,N_820);
or U1338 (N_1338,N_6,N_863);
nor U1339 (N_1339,N_201,N_823);
nand U1340 (N_1340,N_772,N_887);
and U1341 (N_1341,N_773,N_16);
or U1342 (N_1342,N_446,N_509);
or U1343 (N_1343,N_485,N_547);
xor U1344 (N_1344,N_536,N_675);
nor U1345 (N_1345,N_533,N_776);
or U1346 (N_1346,N_758,N_234);
and U1347 (N_1347,N_106,N_285);
and U1348 (N_1348,N_493,N_5);
nand U1349 (N_1349,N_276,N_145);
and U1350 (N_1350,N_913,N_719);
nor U1351 (N_1351,N_363,N_658);
and U1352 (N_1352,N_932,N_432);
and U1353 (N_1353,N_126,N_806);
or U1354 (N_1354,N_191,N_311);
nand U1355 (N_1355,N_672,N_872);
and U1356 (N_1356,N_499,N_632);
nor U1357 (N_1357,N_562,N_798);
xnor U1358 (N_1358,N_366,N_991);
or U1359 (N_1359,N_143,N_360);
or U1360 (N_1360,N_158,N_642);
nand U1361 (N_1361,N_927,N_426);
or U1362 (N_1362,N_272,N_440);
and U1363 (N_1363,N_20,N_357);
nor U1364 (N_1364,N_56,N_3);
and U1365 (N_1365,N_957,N_765);
and U1366 (N_1366,N_513,N_270);
nand U1367 (N_1367,N_15,N_668);
nor U1368 (N_1368,N_466,N_397);
and U1369 (N_1369,N_983,N_374);
nand U1370 (N_1370,N_399,N_193);
and U1371 (N_1371,N_740,N_61);
and U1372 (N_1372,N_894,N_342);
or U1373 (N_1373,N_392,N_227);
and U1374 (N_1374,N_206,N_140);
nor U1375 (N_1375,N_602,N_8);
nor U1376 (N_1376,N_484,N_124);
nand U1377 (N_1377,N_891,N_890);
and U1378 (N_1378,N_208,N_100);
or U1379 (N_1379,N_214,N_954);
nand U1380 (N_1380,N_949,N_138);
and U1381 (N_1381,N_712,N_926);
or U1382 (N_1382,N_611,N_248);
or U1383 (N_1383,N_266,N_706);
nor U1384 (N_1384,N_120,N_893);
or U1385 (N_1385,N_415,N_354);
or U1386 (N_1386,N_763,N_314);
nor U1387 (N_1387,N_144,N_271);
or U1388 (N_1388,N_2,N_830);
nand U1389 (N_1389,N_989,N_858);
nor U1390 (N_1390,N_377,N_79);
and U1391 (N_1391,N_455,N_247);
nor U1392 (N_1392,N_75,N_355);
or U1393 (N_1393,N_422,N_653);
nand U1394 (N_1394,N_689,N_131);
nand U1395 (N_1395,N_892,N_732);
and U1396 (N_1396,N_244,N_530);
and U1397 (N_1397,N_370,N_394);
nor U1398 (N_1398,N_324,N_215);
xor U1399 (N_1399,N_445,N_238);
nor U1400 (N_1400,N_219,N_481);
nand U1401 (N_1401,N_50,N_475);
nand U1402 (N_1402,N_269,N_162);
xnor U1403 (N_1403,N_693,N_105);
or U1404 (N_1404,N_447,N_739);
and U1405 (N_1405,N_490,N_39);
xnor U1406 (N_1406,N_387,N_496);
or U1407 (N_1407,N_918,N_992);
nor U1408 (N_1408,N_336,N_136);
nand U1409 (N_1409,N_378,N_406);
or U1410 (N_1410,N_517,N_945);
or U1411 (N_1411,N_188,N_525);
or U1412 (N_1412,N_735,N_233);
or U1413 (N_1413,N_31,N_348);
nand U1414 (N_1414,N_904,N_9);
or U1415 (N_1415,N_644,N_89);
and U1416 (N_1416,N_249,N_874);
or U1417 (N_1417,N_754,N_936);
xor U1418 (N_1418,N_541,N_851);
or U1419 (N_1419,N_304,N_678);
or U1420 (N_1420,N_738,N_770);
nor U1421 (N_1421,N_253,N_774);
and U1422 (N_1422,N_170,N_654);
nand U1423 (N_1423,N_449,N_386);
or U1424 (N_1424,N_116,N_450);
nor U1425 (N_1425,N_504,N_0);
and U1426 (N_1426,N_651,N_551);
or U1427 (N_1427,N_204,N_984);
and U1428 (N_1428,N_652,N_703);
or U1429 (N_1429,N_185,N_555);
or U1430 (N_1430,N_459,N_28);
nand U1431 (N_1431,N_411,N_321);
nand U1432 (N_1432,N_395,N_850);
nand U1433 (N_1433,N_755,N_43);
or U1434 (N_1434,N_349,N_736);
and U1435 (N_1435,N_963,N_345);
or U1436 (N_1436,N_303,N_871);
nor U1437 (N_1437,N_257,N_903);
or U1438 (N_1438,N_154,N_408);
or U1439 (N_1439,N_373,N_494);
xor U1440 (N_1440,N_557,N_48);
or U1441 (N_1441,N_419,N_876);
or U1442 (N_1442,N_603,N_474);
and U1443 (N_1443,N_786,N_423);
and U1444 (N_1444,N_586,N_407);
or U1445 (N_1445,N_372,N_546);
and U1446 (N_1446,N_277,N_297);
or U1447 (N_1447,N_196,N_695);
and U1448 (N_1448,N_221,N_859);
and U1449 (N_1449,N_478,N_768);
or U1450 (N_1450,N_788,N_966);
nand U1451 (N_1451,N_581,N_615);
or U1452 (N_1452,N_148,N_175);
and U1453 (N_1453,N_980,N_97);
or U1454 (N_1454,N_396,N_622);
nor U1455 (N_1455,N_295,N_760);
or U1456 (N_1456,N_938,N_717);
and U1457 (N_1457,N_563,N_896);
nor U1458 (N_1458,N_909,N_341);
xor U1459 (N_1459,N_218,N_997);
nor U1460 (N_1460,N_265,N_453);
nor U1461 (N_1461,N_480,N_240);
nor U1462 (N_1462,N_662,N_537);
nand U1463 (N_1463,N_104,N_816);
nand U1464 (N_1464,N_598,N_748);
and U1465 (N_1465,N_761,N_71);
nor U1466 (N_1466,N_671,N_795);
nand U1467 (N_1467,N_507,N_928);
nor U1468 (N_1468,N_833,N_470);
or U1469 (N_1469,N_306,N_36);
or U1470 (N_1470,N_73,N_787);
nand U1471 (N_1471,N_400,N_888);
and U1472 (N_1472,N_539,N_702);
nand U1473 (N_1473,N_846,N_766);
nand U1474 (N_1474,N_350,N_836);
xnor U1475 (N_1475,N_573,N_783);
nand U1476 (N_1476,N_698,N_720);
and U1477 (N_1477,N_263,N_620);
and U1478 (N_1478,N_987,N_958);
nor U1479 (N_1479,N_224,N_425);
nor U1480 (N_1480,N_506,N_254);
nor U1481 (N_1481,N_64,N_312);
xor U1482 (N_1482,N_687,N_19);
nor U1483 (N_1483,N_612,N_574);
or U1484 (N_1484,N_460,N_538);
or U1485 (N_1485,N_725,N_289);
or U1486 (N_1486,N_37,N_799);
nor U1487 (N_1487,N_160,N_821);
nor U1488 (N_1488,N_715,N_856);
or U1489 (N_1489,N_961,N_998);
and U1490 (N_1490,N_708,N_91);
and U1491 (N_1491,N_187,N_457);
and U1492 (N_1492,N_950,N_895);
and U1493 (N_1493,N_164,N_730);
nor U1494 (N_1494,N_627,N_172);
nor U1495 (N_1495,N_910,N_169);
and U1496 (N_1496,N_92,N_544);
or U1497 (N_1497,N_974,N_880);
xor U1498 (N_1498,N_988,N_102);
nor U1499 (N_1499,N_403,N_985);
and U1500 (N_1500,N_639,N_566);
xor U1501 (N_1501,N_10,N_735);
and U1502 (N_1502,N_206,N_321);
nand U1503 (N_1503,N_444,N_449);
xor U1504 (N_1504,N_1,N_708);
or U1505 (N_1505,N_966,N_550);
or U1506 (N_1506,N_437,N_20);
nand U1507 (N_1507,N_607,N_74);
or U1508 (N_1508,N_93,N_448);
and U1509 (N_1509,N_999,N_332);
nor U1510 (N_1510,N_115,N_360);
and U1511 (N_1511,N_119,N_171);
and U1512 (N_1512,N_806,N_395);
nand U1513 (N_1513,N_691,N_86);
or U1514 (N_1514,N_509,N_833);
xnor U1515 (N_1515,N_22,N_461);
or U1516 (N_1516,N_947,N_993);
or U1517 (N_1517,N_363,N_567);
or U1518 (N_1518,N_894,N_559);
xnor U1519 (N_1519,N_581,N_636);
or U1520 (N_1520,N_588,N_152);
or U1521 (N_1521,N_600,N_341);
nor U1522 (N_1522,N_847,N_155);
or U1523 (N_1523,N_146,N_123);
or U1524 (N_1524,N_800,N_21);
xor U1525 (N_1525,N_977,N_820);
xor U1526 (N_1526,N_581,N_796);
or U1527 (N_1527,N_255,N_308);
nor U1528 (N_1528,N_944,N_233);
nor U1529 (N_1529,N_371,N_187);
nand U1530 (N_1530,N_262,N_572);
nand U1531 (N_1531,N_427,N_371);
and U1532 (N_1532,N_289,N_678);
xnor U1533 (N_1533,N_118,N_554);
and U1534 (N_1534,N_144,N_641);
nor U1535 (N_1535,N_357,N_188);
nand U1536 (N_1536,N_937,N_480);
or U1537 (N_1537,N_76,N_549);
nand U1538 (N_1538,N_827,N_766);
nand U1539 (N_1539,N_91,N_770);
nand U1540 (N_1540,N_374,N_111);
or U1541 (N_1541,N_553,N_860);
nand U1542 (N_1542,N_438,N_276);
nor U1543 (N_1543,N_621,N_681);
nand U1544 (N_1544,N_441,N_444);
nand U1545 (N_1545,N_267,N_13);
nor U1546 (N_1546,N_746,N_405);
nand U1547 (N_1547,N_612,N_654);
or U1548 (N_1548,N_800,N_458);
xor U1549 (N_1549,N_165,N_872);
nor U1550 (N_1550,N_404,N_940);
nor U1551 (N_1551,N_640,N_830);
nand U1552 (N_1552,N_687,N_128);
and U1553 (N_1553,N_122,N_680);
and U1554 (N_1554,N_533,N_675);
and U1555 (N_1555,N_14,N_32);
nor U1556 (N_1556,N_174,N_482);
or U1557 (N_1557,N_246,N_579);
or U1558 (N_1558,N_974,N_569);
nor U1559 (N_1559,N_497,N_89);
or U1560 (N_1560,N_373,N_824);
and U1561 (N_1561,N_968,N_57);
or U1562 (N_1562,N_525,N_879);
xnor U1563 (N_1563,N_759,N_970);
nand U1564 (N_1564,N_870,N_446);
or U1565 (N_1565,N_476,N_909);
nand U1566 (N_1566,N_670,N_484);
nand U1567 (N_1567,N_340,N_257);
or U1568 (N_1568,N_420,N_58);
or U1569 (N_1569,N_968,N_698);
or U1570 (N_1570,N_445,N_616);
nor U1571 (N_1571,N_593,N_327);
nor U1572 (N_1572,N_645,N_550);
nor U1573 (N_1573,N_237,N_966);
nand U1574 (N_1574,N_655,N_673);
nand U1575 (N_1575,N_120,N_307);
or U1576 (N_1576,N_284,N_988);
and U1577 (N_1577,N_522,N_570);
or U1578 (N_1578,N_277,N_223);
and U1579 (N_1579,N_24,N_279);
nand U1580 (N_1580,N_399,N_330);
and U1581 (N_1581,N_729,N_167);
or U1582 (N_1582,N_20,N_931);
nor U1583 (N_1583,N_794,N_102);
nand U1584 (N_1584,N_849,N_602);
xor U1585 (N_1585,N_79,N_172);
xnor U1586 (N_1586,N_124,N_470);
nor U1587 (N_1587,N_733,N_876);
or U1588 (N_1588,N_718,N_684);
nor U1589 (N_1589,N_716,N_431);
nand U1590 (N_1590,N_542,N_28);
xor U1591 (N_1591,N_740,N_613);
or U1592 (N_1592,N_570,N_195);
nand U1593 (N_1593,N_74,N_988);
xor U1594 (N_1594,N_467,N_293);
nand U1595 (N_1595,N_174,N_265);
nand U1596 (N_1596,N_312,N_666);
and U1597 (N_1597,N_304,N_718);
nand U1598 (N_1598,N_91,N_844);
nand U1599 (N_1599,N_375,N_632);
nor U1600 (N_1600,N_708,N_287);
nor U1601 (N_1601,N_461,N_27);
and U1602 (N_1602,N_134,N_358);
or U1603 (N_1603,N_730,N_585);
nor U1604 (N_1604,N_698,N_316);
nor U1605 (N_1605,N_746,N_119);
nand U1606 (N_1606,N_622,N_419);
or U1607 (N_1607,N_55,N_688);
nand U1608 (N_1608,N_869,N_924);
xnor U1609 (N_1609,N_426,N_946);
and U1610 (N_1610,N_314,N_738);
xnor U1611 (N_1611,N_289,N_983);
or U1612 (N_1612,N_263,N_289);
xnor U1613 (N_1613,N_915,N_511);
nand U1614 (N_1614,N_584,N_28);
or U1615 (N_1615,N_438,N_325);
and U1616 (N_1616,N_914,N_894);
or U1617 (N_1617,N_442,N_644);
and U1618 (N_1618,N_453,N_219);
nand U1619 (N_1619,N_308,N_122);
nor U1620 (N_1620,N_319,N_379);
or U1621 (N_1621,N_611,N_960);
and U1622 (N_1622,N_752,N_555);
and U1623 (N_1623,N_504,N_433);
and U1624 (N_1624,N_78,N_721);
xor U1625 (N_1625,N_126,N_309);
nand U1626 (N_1626,N_259,N_615);
or U1627 (N_1627,N_146,N_104);
nor U1628 (N_1628,N_457,N_536);
xnor U1629 (N_1629,N_888,N_932);
nand U1630 (N_1630,N_150,N_180);
nand U1631 (N_1631,N_965,N_658);
nor U1632 (N_1632,N_664,N_601);
nor U1633 (N_1633,N_360,N_729);
and U1634 (N_1634,N_697,N_160);
or U1635 (N_1635,N_608,N_133);
nor U1636 (N_1636,N_975,N_900);
nor U1637 (N_1637,N_934,N_305);
and U1638 (N_1638,N_582,N_453);
nand U1639 (N_1639,N_885,N_133);
nor U1640 (N_1640,N_119,N_574);
xor U1641 (N_1641,N_876,N_595);
and U1642 (N_1642,N_79,N_163);
or U1643 (N_1643,N_864,N_776);
and U1644 (N_1644,N_847,N_929);
nand U1645 (N_1645,N_544,N_992);
or U1646 (N_1646,N_164,N_365);
or U1647 (N_1647,N_905,N_284);
or U1648 (N_1648,N_158,N_870);
nor U1649 (N_1649,N_358,N_126);
nor U1650 (N_1650,N_32,N_291);
nand U1651 (N_1651,N_169,N_974);
and U1652 (N_1652,N_649,N_116);
xnor U1653 (N_1653,N_52,N_106);
nand U1654 (N_1654,N_881,N_447);
xnor U1655 (N_1655,N_853,N_760);
xnor U1656 (N_1656,N_694,N_669);
nor U1657 (N_1657,N_598,N_395);
or U1658 (N_1658,N_583,N_807);
or U1659 (N_1659,N_506,N_205);
or U1660 (N_1660,N_139,N_654);
and U1661 (N_1661,N_275,N_20);
or U1662 (N_1662,N_294,N_379);
and U1663 (N_1663,N_158,N_413);
or U1664 (N_1664,N_109,N_711);
nor U1665 (N_1665,N_798,N_86);
nand U1666 (N_1666,N_388,N_127);
xor U1667 (N_1667,N_883,N_927);
and U1668 (N_1668,N_191,N_594);
xor U1669 (N_1669,N_65,N_228);
xor U1670 (N_1670,N_76,N_811);
and U1671 (N_1671,N_256,N_609);
and U1672 (N_1672,N_371,N_984);
and U1673 (N_1673,N_600,N_560);
nand U1674 (N_1674,N_98,N_575);
xor U1675 (N_1675,N_563,N_807);
or U1676 (N_1676,N_347,N_522);
nand U1677 (N_1677,N_105,N_969);
nand U1678 (N_1678,N_653,N_313);
and U1679 (N_1679,N_249,N_679);
or U1680 (N_1680,N_80,N_775);
or U1681 (N_1681,N_921,N_184);
and U1682 (N_1682,N_639,N_63);
nand U1683 (N_1683,N_629,N_483);
nor U1684 (N_1684,N_786,N_622);
nor U1685 (N_1685,N_541,N_431);
nand U1686 (N_1686,N_95,N_174);
xnor U1687 (N_1687,N_923,N_974);
nand U1688 (N_1688,N_176,N_404);
or U1689 (N_1689,N_446,N_615);
nor U1690 (N_1690,N_509,N_496);
nand U1691 (N_1691,N_269,N_671);
or U1692 (N_1692,N_202,N_736);
or U1693 (N_1693,N_981,N_242);
or U1694 (N_1694,N_228,N_947);
nor U1695 (N_1695,N_692,N_426);
nor U1696 (N_1696,N_458,N_660);
and U1697 (N_1697,N_734,N_8);
nor U1698 (N_1698,N_729,N_350);
or U1699 (N_1699,N_720,N_991);
or U1700 (N_1700,N_428,N_477);
xor U1701 (N_1701,N_471,N_643);
and U1702 (N_1702,N_717,N_662);
or U1703 (N_1703,N_910,N_680);
and U1704 (N_1704,N_837,N_423);
nor U1705 (N_1705,N_198,N_112);
nand U1706 (N_1706,N_994,N_512);
xor U1707 (N_1707,N_395,N_656);
and U1708 (N_1708,N_968,N_937);
xnor U1709 (N_1709,N_149,N_202);
nand U1710 (N_1710,N_912,N_36);
nor U1711 (N_1711,N_371,N_198);
and U1712 (N_1712,N_101,N_446);
xnor U1713 (N_1713,N_58,N_150);
and U1714 (N_1714,N_7,N_564);
nand U1715 (N_1715,N_596,N_685);
nand U1716 (N_1716,N_813,N_874);
and U1717 (N_1717,N_959,N_132);
nand U1718 (N_1718,N_978,N_292);
nor U1719 (N_1719,N_353,N_923);
xor U1720 (N_1720,N_143,N_256);
or U1721 (N_1721,N_760,N_732);
nor U1722 (N_1722,N_881,N_712);
nor U1723 (N_1723,N_916,N_38);
and U1724 (N_1724,N_86,N_370);
xnor U1725 (N_1725,N_182,N_583);
and U1726 (N_1726,N_929,N_575);
nand U1727 (N_1727,N_8,N_439);
nand U1728 (N_1728,N_860,N_912);
nand U1729 (N_1729,N_124,N_988);
and U1730 (N_1730,N_672,N_130);
or U1731 (N_1731,N_465,N_496);
nand U1732 (N_1732,N_811,N_422);
and U1733 (N_1733,N_604,N_119);
and U1734 (N_1734,N_714,N_504);
xnor U1735 (N_1735,N_236,N_341);
nand U1736 (N_1736,N_845,N_279);
nor U1737 (N_1737,N_292,N_745);
nand U1738 (N_1738,N_164,N_665);
nor U1739 (N_1739,N_821,N_208);
or U1740 (N_1740,N_117,N_623);
nand U1741 (N_1741,N_44,N_46);
and U1742 (N_1742,N_319,N_913);
nand U1743 (N_1743,N_17,N_702);
nand U1744 (N_1744,N_241,N_27);
xnor U1745 (N_1745,N_677,N_473);
or U1746 (N_1746,N_515,N_395);
or U1747 (N_1747,N_403,N_507);
nand U1748 (N_1748,N_977,N_505);
and U1749 (N_1749,N_521,N_315);
or U1750 (N_1750,N_689,N_678);
or U1751 (N_1751,N_297,N_867);
xnor U1752 (N_1752,N_153,N_660);
nor U1753 (N_1753,N_406,N_267);
and U1754 (N_1754,N_820,N_865);
xnor U1755 (N_1755,N_174,N_46);
or U1756 (N_1756,N_733,N_155);
or U1757 (N_1757,N_551,N_418);
nor U1758 (N_1758,N_607,N_255);
or U1759 (N_1759,N_498,N_609);
or U1760 (N_1760,N_584,N_807);
and U1761 (N_1761,N_663,N_962);
and U1762 (N_1762,N_97,N_751);
or U1763 (N_1763,N_695,N_525);
and U1764 (N_1764,N_64,N_213);
and U1765 (N_1765,N_68,N_617);
nand U1766 (N_1766,N_377,N_240);
nand U1767 (N_1767,N_857,N_231);
and U1768 (N_1768,N_800,N_965);
nor U1769 (N_1769,N_827,N_47);
and U1770 (N_1770,N_850,N_409);
nand U1771 (N_1771,N_989,N_647);
nor U1772 (N_1772,N_609,N_504);
xnor U1773 (N_1773,N_921,N_562);
nor U1774 (N_1774,N_166,N_575);
nor U1775 (N_1775,N_78,N_806);
nand U1776 (N_1776,N_666,N_433);
nand U1777 (N_1777,N_271,N_396);
and U1778 (N_1778,N_839,N_724);
or U1779 (N_1779,N_918,N_220);
nor U1780 (N_1780,N_923,N_260);
or U1781 (N_1781,N_608,N_405);
or U1782 (N_1782,N_864,N_198);
or U1783 (N_1783,N_628,N_870);
nor U1784 (N_1784,N_529,N_937);
xnor U1785 (N_1785,N_114,N_935);
or U1786 (N_1786,N_202,N_987);
nor U1787 (N_1787,N_586,N_224);
or U1788 (N_1788,N_815,N_724);
and U1789 (N_1789,N_115,N_339);
nand U1790 (N_1790,N_270,N_668);
nand U1791 (N_1791,N_997,N_346);
nor U1792 (N_1792,N_341,N_991);
nand U1793 (N_1793,N_362,N_756);
nand U1794 (N_1794,N_107,N_925);
and U1795 (N_1795,N_683,N_546);
and U1796 (N_1796,N_359,N_186);
xnor U1797 (N_1797,N_96,N_396);
and U1798 (N_1798,N_176,N_880);
and U1799 (N_1799,N_477,N_902);
and U1800 (N_1800,N_765,N_63);
nand U1801 (N_1801,N_659,N_21);
or U1802 (N_1802,N_265,N_317);
nor U1803 (N_1803,N_65,N_238);
nand U1804 (N_1804,N_104,N_876);
or U1805 (N_1805,N_534,N_582);
xor U1806 (N_1806,N_945,N_241);
nand U1807 (N_1807,N_935,N_180);
nand U1808 (N_1808,N_1,N_54);
nand U1809 (N_1809,N_260,N_940);
nand U1810 (N_1810,N_129,N_866);
or U1811 (N_1811,N_78,N_927);
nand U1812 (N_1812,N_429,N_266);
xnor U1813 (N_1813,N_119,N_811);
and U1814 (N_1814,N_866,N_188);
nor U1815 (N_1815,N_877,N_987);
nor U1816 (N_1816,N_943,N_605);
nand U1817 (N_1817,N_114,N_538);
nand U1818 (N_1818,N_6,N_547);
or U1819 (N_1819,N_775,N_834);
nand U1820 (N_1820,N_424,N_791);
and U1821 (N_1821,N_1,N_156);
xor U1822 (N_1822,N_600,N_743);
and U1823 (N_1823,N_273,N_634);
and U1824 (N_1824,N_25,N_515);
nor U1825 (N_1825,N_223,N_696);
nand U1826 (N_1826,N_565,N_566);
nand U1827 (N_1827,N_614,N_820);
and U1828 (N_1828,N_783,N_753);
or U1829 (N_1829,N_956,N_914);
and U1830 (N_1830,N_194,N_681);
or U1831 (N_1831,N_119,N_183);
nor U1832 (N_1832,N_829,N_553);
or U1833 (N_1833,N_861,N_311);
nand U1834 (N_1834,N_658,N_390);
nor U1835 (N_1835,N_511,N_170);
and U1836 (N_1836,N_308,N_722);
nand U1837 (N_1837,N_932,N_36);
nand U1838 (N_1838,N_151,N_450);
and U1839 (N_1839,N_210,N_731);
nor U1840 (N_1840,N_74,N_932);
nand U1841 (N_1841,N_807,N_207);
and U1842 (N_1842,N_606,N_277);
and U1843 (N_1843,N_164,N_310);
or U1844 (N_1844,N_921,N_700);
or U1845 (N_1845,N_837,N_579);
and U1846 (N_1846,N_192,N_522);
and U1847 (N_1847,N_740,N_805);
xnor U1848 (N_1848,N_724,N_400);
or U1849 (N_1849,N_132,N_428);
and U1850 (N_1850,N_200,N_512);
or U1851 (N_1851,N_673,N_354);
and U1852 (N_1852,N_317,N_568);
nand U1853 (N_1853,N_137,N_601);
and U1854 (N_1854,N_962,N_25);
and U1855 (N_1855,N_865,N_448);
and U1856 (N_1856,N_418,N_533);
nand U1857 (N_1857,N_423,N_783);
nand U1858 (N_1858,N_751,N_933);
nor U1859 (N_1859,N_579,N_344);
nor U1860 (N_1860,N_698,N_399);
nor U1861 (N_1861,N_540,N_179);
nand U1862 (N_1862,N_114,N_426);
and U1863 (N_1863,N_866,N_601);
or U1864 (N_1864,N_616,N_401);
and U1865 (N_1865,N_582,N_694);
nand U1866 (N_1866,N_708,N_25);
nor U1867 (N_1867,N_477,N_422);
or U1868 (N_1868,N_141,N_497);
and U1869 (N_1869,N_257,N_587);
and U1870 (N_1870,N_891,N_94);
xor U1871 (N_1871,N_687,N_336);
xor U1872 (N_1872,N_598,N_647);
and U1873 (N_1873,N_688,N_852);
nand U1874 (N_1874,N_942,N_879);
and U1875 (N_1875,N_446,N_516);
or U1876 (N_1876,N_976,N_167);
xnor U1877 (N_1877,N_439,N_990);
xor U1878 (N_1878,N_862,N_141);
and U1879 (N_1879,N_598,N_625);
or U1880 (N_1880,N_502,N_734);
or U1881 (N_1881,N_798,N_377);
or U1882 (N_1882,N_35,N_127);
nand U1883 (N_1883,N_637,N_184);
nand U1884 (N_1884,N_457,N_833);
nand U1885 (N_1885,N_252,N_97);
nand U1886 (N_1886,N_6,N_906);
nand U1887 (N_1887,N_390,N_269);
nand U1888 (N_1888,N_310,N_626);
or U1889 (N_1889,N_383,N_184);
nor U1890 (N_1890,N_754,N_959);
nor U1891 (N_1891,N_844,N_685);
and U1892 (N_1892,N_240,N_975);
nor U1893 (N_1893,N_297,N_166);
or U1894 (N_1894,N_94,N_293);
nor U1895 (N_1895,N_848,N_617);
or U1896 (N_1896,N_782,N_427);
nand U1897 (N_1897,N_969,N_756);
nor U1898 (N_1898,N_237,N_168);
and U1899 (N_1899,N_304,N_497);
nor U1900 (N_1900,N_455,N_937);
and U1901 (N_1901,N_782,N_319);
nand U1902 (N_1902,N_619,N_778);
nand U1903 (N_1903,N_689,N_719);
xnor U1904 (N_1904,N_15,N_11);
nor U1905 (N_1905,N_934,N_236);
and U1906 (N_1906,N_351,N_404);
nor U1907 (N_1907,N_804,N_423);
and U1908 (N_1908,N_206,N_326);
nand U1909 (N_1909,N_683,N_731);
nor U1910 (N_1910,N_577,N_563);
nor U1911 (N_1911,N_474,N_143);
xnor U1912 (N_1912,N_653,N_33);
or U1913 (N_1913,N_421,N_34);
or U1914 (N_1914,N_211,N_500);
and U1915 (N_1915,N_930,N_632);
and U1916 (N_1916,N_669,N_309);
nor U1917 (N_1917,N_322,N_565);
nor U1918 (N_1918,N_254,N_262);
or U1919 (N_1919,N_388,N_788);
or U1920 (N_1920,N_175,N_627);
nor U1921 (N_1921,N_111,N_452);
and U1922 (N_1922,N_954,N_541);
or U1923 (N_1923,N_323,N_660);
or U1924 (N_1924,N_977,N_245);
xnor U1925 (N_1925,N_753,N_950);
or U1926 (N_1926,N_881,N_200);
and U1927 (N_1927,N_972,N_778);
nand U1928 (N_1928,N_837,N_660);
nor U1929 (N_1929,N_547,N_281);
or U1930 (N_1930,N_249,N_432);
and U1931 (N_1931,N_728,N_936);
and U1932 (N_1932,N_110,N_9);
and U1933 (N_1933,N_816,N_108);
or U1934 (N_1934,N_517,N_33);
nand U1935 (N_1935,N_801,N_229);
and U1936 (N_1936,N_277,N_433);
or U1937 (N_1937,N_14,N_305);
or U1938 (N_1938,N_694,N_876);
nor U1939 (N_1939,N_692,N_175);
or U1940 (N_1940,N_301,N_718);
nor U1941 (N_1941,N_444,N_653);
nand U1942 (N_1942,N_251,N_778);
nor U1943 (N_1943,N_152,N_494);
or U1944 (N_1944,N_278,N_237);
and U1945 (N_1945,N_399,N_963);
or U1946 (N_1946,N_471,N_474);
or U1947 (N_1947,N_125,N_211);
or U1948 (N_1948,N_410,N_639);
nand U1949 (N_1949,N_48,N_590);
nor U1950 (N_1950,N_545,N_375);
xnor U1951 (N_1951,N_301,N_867);
and U1952 (N_1952,N_351,N_591);
and U1953 (N_1953,N_61,N_531);
or U1954 (N_1954,N_294,N_743);
nor U1955 (N_1955,N_679,N_180);
xor U1956 (N_1956,N_462,N_438);
nand U1957 (N_1957,N_378,N_773);
or U1958 (N_1958,N_138,N_728);
and U1959 (N_1959,N_821,N_846);
nand U1960 (N_1960,N_565,N_933);
nor U1961 (N_1961,N_630,N_941);
and U1962 (N_1962,N_201,N_434);
xnor U1963 (N_1963,N_149,N_420);
and U1964 (N_1964,N_128,N_169);
nand U1965 (N_1965,N_814,N_411);
or U1966 (N_1966,N_837,N_643);
and U1967 (N_1967,N_900,N_250);
nand U1968 (N_1968,N_149,N_576);
or U1969 (N_1969,N_915,N_714);
or U1970 (N_1970,N_443,N_240);
or U1971 (N_1971,N_932,N_396);
nor U1972 (N_1972,N_183,N_637);
nor U1973 (N_1973,N_609,N_513);
and U1974 (N_1974,N_973,N_576);
nor U1975 (N_1975,N_933,N_274);
or U1976 (N_1976,N_112,N_55);
nor U1977 (N_1977,N_46,N_216);
nor U1978 (N_1978,N_623,N_358);
xnor U1979 (N_1979,N_352,N_310);
and U1980 (N_1980,N_836,N_258);
and U1981 (N_1981,N_865,N_154);
nand U1982 (N_1982,N_311,N_626);
nor U1983 (N_1983,N_587,N_520);
nor U1984 (N_1984,N_849,N_44);
and U1985 (N_1985,N_786,N_958);
and U1986 (N_1986,N_531,N_821);
or U1987 (N_1987,N_211,N_76);
and U1988 (N_1988,N_802,N_528);
nor U1989 (N_1989,N_67,N_214);
or U1990 (N_1990,N_926,N_841);
or U1991 (N_1991,N_192,N_938);
and U1992 (N_1992,N_375,N_341);
xor U1993 (N_1993,N_375,N_167);
or U1994 (N_1994,N_725,N_8);
nor U1995 (N_1995,N_804,N_580);
nor U1996 (N_1996,N_569,N_540);
or U1997 (N_1997,N_671,N_134);
nand U1998 (N_1998,N_520,N_114);
and U1999 (N_1999,N_411,N_864);
nand U2000 (N_2000,N_1889,N_1672);
or U2001 (N_2001,N_1075,N_1210);
nand U2002 (N_2002,N_1510,N_1057);
nand U2003 (N_2003,N_1228,N_1560);
nor U2004 (N_2004,N_1989,N_1163);
nand U2005 (N_2005,N_1070,N_1985);
and U2006 (N_2006,N_1820,N_1458);
or U2007 (N_2007,N_1673,N_1624);
nand U2008 (N_2008,N_1243,N_1361);
and U2009 (N_2009,N_1067,N_1226);
or U2010 (N_2010,N_1050,N_1537);
and U2011 (N_2011,N_1151,N_1431);
nand U2012 (N_2012,N_1851,N_1375);
or U2013 (N_2013,N_1507,N_1858);
nand U2014 (N_2014,N_1407,N_1659);
or U2015 (N_2015,N_1699,N_1473);
or U2016 (N_2016,N_1114,N_1710);
or U2017 (N_2017,N_1552,N_1845);
xnor U2018 (N_2018,N_1104,N_1235);
nor U2019 (N_2019,N_1541,N_1940);
and U2020 (N_2020,N_1011,N_1367);
nand U2021 (N_2021,N_1325,N_1290);
nor U2022 (N_2022,N_1358,N_1780);
or U2023 (N_2023,N_1239,N_1834);
nand U2024 (N_2024,N_1006,N_1188);
xnor U2025 (N_2025,N_1785,N_1946);
or U2026 (N_2026,N_1765,N_1562);
or U2027 (N_2027,N_1664,N_1982);
xor U2028 (N_2028,N_1878,N_1509);
and U2029 (N_2029,N_1811,N_1886);
nand U2030 (N_2030,N_1001,N_1026);
or U2031 (N_2031,N_1821,N_1744);
or U2032 (N_2032,N_1378,N_1444);
or U2033 (N_2033,N_1696,N_1606);
nand U2034 (N_2034,N_1438,N_1351);
and U2035 (N_2035,N_1663,N_1047);
or U2036 (N_2036,N_1786,N_1233);
or U2037 (N_2037,N_1455,N_1379);
nand U2038 (N_2038,N_1413,N_1700);
nand U2039 (N_2039,N_1144,N_1198);
xor U2040 (N_2040,N_1077,N_1345);
nand U2041 (N_2041,N_1495,N_1652);
and U2042 (N_2042,N_1644,N_1120);
or U2043 (N_2043,N_1733,N_1062);
nand U2044 (N_2044,N_1098,N_1279);
nand U2045 (N_2045,N_1857,N_1176);
nor U2046 (N_2046,N_1712,N_1748);
nor U2047 (N_2047,N_1156,N_1517);
and U2048 (N_2048,N_1615,N_1997);
nand U2049 (N_2049,N_1569,N_1830);
nand U2050 (N_2050,N_1819,N_1304);
xor U2051 (N_2051,N_1079,N_1585);
or U2052 (N_2052,N_1996,N_1284);
nand U2053 (N_2053,N_1271,N_1262);
and U2054 (N_2054,N_1848,N_1576);
xnor U2055 (N_2055,N_1586,N_1191);
or U2056 (N_2056,N_1686,N_1714);
and U2057 (N_2057,N_1335,N_1933);
nand U2058 (N_2058,N_1272,N_1485);
nand U2059 (N_2059,N_1386,N_1010);
nor U2060 (N_2060,N_1154,N_1557);
or U2061 (N_2061,N_1429,N_1302);
nor U2062 (N_2062,N_1501,N_1391);
nor U2063 (N_2063,N_1462,N_1148);
nor U2064 (N_2064,N_1604,N_1420);
or U2065 (N_2065,N_1954,N_1003);
or U2066 (N_2066,N_1555,N_1978);
nand U2067 (N_2067,N_1331,N_1125);
nand U2068 (N_2068,N_1334,N_1919);
nor U2069 (N_2069,N_1698,N_1625);
nand U2070 (N_2070,N_1161,N_1309);
and U2071 (N_2071,N_1986,N_1147);
nand U2072 (N_2072,N_1666,N_1425);
nand U2073 (N_2073,N_1803,N_1582);
or U2074 (N_2074,N_1701,N_1891);
and U2075 (N_2075,N_1587,N_1969);
nor U2076 (N_2076,N_1846,N_1095);
nor U2077 (N_2077,N_1256,N_1926);
or U2078 (N_2078,N_1734,N_1016);
or U2079 (N_2079,N_1491,N_1071);
nor U2080 (N_2080,N_1729,N_1289);
or U2081 (N_2081,N_1532,N_1287);
and U2082 (N_2082,N_1253,N_1382);
or U2083 (N_2083,N_1195,N_1205);
nand U2084 (N_2084,N_1190,N_1091);
or U2085 (N_2085,N_1405,N_1179);
or U2086 (N_2086,N_1577,N_1705);
or U2087 (N_2087,N_1832,N_1564);
or U2088 (N_2088,N_1634,N_1241);
nor U2089 (N_2089,N_1038,N_1101);
and U2090 (N_2090,N_1691,N_1472);
nand U2091 (N_2091,N_1324,N_1806);
xnor U2092 (N_2092,N_1910,N_1145);
xor U2093 (N_2093,N_1988,N_1981);
nand U2094 (N_2094,N_1935,N_1119);
and U2095 (N_2095,N_1048,N_1605);
or U2096 (N_2096,N_1767,N_1214);
nor U2097 (N_2097,N_1764,N_1799);
or U2098 (N_2098,N_1169,N_1034);
xor U2099 (N_2099,N_1907,N_1841);
nor U2100 (N_2100,N_1224,N_1249);
and U2101 (N_2101,N_1657,N_1974);
nand U2102 (N_2102,N_1028,N_1958);
or U2103 (N_2103,N_1877,N_1310);
and U2104 (N_2104,N_1110,N_1392);
or U2105 (N_2105,N_1860,N_1206);
nand U2106 (N_2106,N_1423,N_1208);
or U2107 (N_2107,N_1137,N_1061);
and U2108 (N_2108,N_1890,N_1181);
or U2109 (N_2109,N_1066,N_1685);
xor U2110 (N_2110,N_1893,N_1427);
nand U2111 (N_2111,N_1627,N_1017);
or U2112 (N_2112,N_1103,N_1503);
nor U2113 (N_2113,N_1064,N_1404);
or U2114 (N_2114,N_1111,N_1209);
or U2115 (N_2115,N_1313,N_1294);
or U2116 (N_2116,N_1355,N_1941);
and U2117 (N_2117,N_1393,N_1432);
nand U2118 (N_2118,N_1506,N_1092);
nand U2119 (N_2119,N_1276,N_1623);
nor U2120 (N_2120,N_1646,N_1496);
nand U2121 (N_2121,N_1757,N_1593);
nand U2122 (N_2122,N_1342,N_1187);
and U2123 (N_2123,N_1838,N_1162);
nor U2124 (N_2124,N_1245,N_1452);
nand U2125 (N_2125,N_1398,N_1166);
nor U2126 (N_2126,N_1130,N_1369);
nand U2127 (N_2127,N_1426,N_1676);
and U2128 (N_2128,N_1327,N_1372);
xor U2129 (N_2129,N_1688,N_1338);
or U2130 (N_2130,N_1109,N_1063);
xor U2131 (N_2131,N_1184,N_1683);
nor U2132 (N_2132,N_1598,N_1620);
or U2133 (N_2133,N_1059,N_1493);
xor U2134 (N_2134,N_1527,N_1315);
and U2135 (N_2135,N_1497,N_1603);
nand U2136 (N_2136,N_1424,N_1466);
nor U2137 (N_2137,N_1029,N_1645);
nor U2138 (N_2138,N_1222,N_1177);
nand U2139 (N_2139,N_1611,N_1252);
nand U2140 (N_2140,N_1597,N_1015);
and U2141 (N_2141,N_1809,N_1121);
or U2142 (N_2142,N_1217,N_1844);
or U2143 (N_2143,N_1353,N_1648);
nand U2144 (N_2144,N_1876,N_1285);
nor U2145 (N_2145,N_1913,N_1600);
or U2146 (N_2146,N_1182,N_1990);
nand U2147 (N_2147,N_1759,N_1779);
nor U2148 (N_2148,N_1875,N_1783);
nand U2149 (N_2149,N_1678,N_1430);
or U2150 (N_2150,N_1124,N_1387);
nor U2151 (N_2151,N_1229,N_1739);
nor U2152 (N_2152,N_1330,N_1127);
and U2153 (N_2153,N_1388,N_1661);
nor U2154 (N_2154,N_1321,N_1697);
nand U2155 (N_2155,N_1453,N_1972);
and U2156 (N_2156,N_1194,N_1522);
nand U2157 (N_2157,N_1728,N_1230);
nor U2158 (N_2158,N_1917,N_1930);
nand U2159 (N_2159,N_1662,N_1140);
nor U2160 (N_2160,N_1505,N_1789);
nand U2161 (N_2161,N_1174,N_1945);
nand U2162 (N_2162,N_1536,N_1867);
or U2163 (N_2163,N_1793,N_1483);
nor U2164 (N_2164,N_1628,N_1197);
and U2165 (N_2165,N_1238,N_1080);
nand U2166 (N_2166,N_1359,N_1456);
nand U2167 (N_2167,N_1277,N_1590);
nor U2168 (N_2168,N_1344,N_1074);
xor U2169 (N_2169,N_1559,N_1549);
or U2170 (N_2170,N_1533,N_1060);
nand U2171 (N_2171,N_1370,N_1283);
or U2172 (N_2172,N_1570,N_1297);
nor U2173 (N_2173,N_1923,N_1594);
nand U2174 (N_2174,N_1964,N_1305);
and U2175 (N_2175,N_1436,N_1827);
and U2176 (N_2176,N_1873,N_1949);
nand U2177 (N_2177,N_1914,N_1725);
xnor U2178 (N_2178,N_1643,N_1642);
xor U2179 (N_2179,N_1126,N_1031);
nor U2180 (N_2180,N_1944,N_1660);
or U2181 (N_2181,N_1084,N_1521);
nand U2182 (N_2182,N_1086,N_1399);
or U2183 (N_2183,N_1747,N_1952);
nand U2184 (N_2184,N_1193,N_1754);
and U2185 (N_2185,N_1682,N_1106);
nor U2186 (N_2186,N_1295,N_1215);
or U2187 (N_2187,N_1992,N_1171);
and U2188 (N_2188,N_1870,N_1030);
xnor U2189 (N_2189,N_1653,N_1036);
or U2190 (N_2190,N_1775,N_1671);
or U2191 (N_2191,N_1146,N_1102);
nand U2192 (N_2192,N_1881,N_1300);
and U2193 (N_2193,N_1143,N_1572);
or U2194 (N_2194,N_1897,N_1412);
nor U2195 (N_2195,N_1264,N_1790);
and U2196 (N_2196,N_1979,N_1609);
xor U2197 (N_2197,N_1810,N_1674);
nand U2198 (N_2198,N_1575,N_1500);
nand U2199 (N_2199,N_1356,N_1170);
nand U2200 (N_2200,N_1039,N_1680);
xnor U2201 (N_2201,N_1439,N_1180);
or U2202 (N_2202,N_1668,N_1141);
nand U2203 (N_2203,N_1513,N_1901);
nand U2204 (N_2204,N_1022,N_1406);
and U2205 (N_2205,N_1737,N_1854);
nor U2206 (N_2206,N_1390,N_1042);
and U2207 (N_2207,N_1385,N_1463);
nor U2208 (N_2208,N_1859,N_1094);
nand U2209 (N_2209,N_1526,N_1475);
and U2210 (N_2210,N_1236,N_1818);
or U2211 (N_2211,N_1902,N_1192);
nand U2212 (N_2212,N_1089,N_1723);
nor U2213 (N_2213,N_1445,N_1993);
or U2214 (N_2214,N_1855,N_1021);
and U2215 (N_2215,N_1548,N_1203);
or U2216 (N_2216,N_1839,N_1097);
and U2217 (N_2217,N_1937,N_1292);
nand U2218 (N_2218,N_1638,N_1437);
xnor U2219 (N_2219,N_1658,N_1622);
or U2220 (N_2220,N_1987,N_1449);
or U2221 (N_2221,N_1263,N_1411);
nor U2222 (N_2222,N_1363,N_1168);
and U2223 (N_2223,N_1322,N_1962);
and U2224 (N_2224,N_1178,N_1231);
and U2225 (N_2225,N_1514,N_1581);
or U2226 (N_2226,N_1395,N_1380);
or U2227 (N_2227,N_1677,N_1885);
and U2228 (N_2228,N_1694,N_1211);
nand U2229 (N_2229,N_1630,N_1976);
nand U2230 (N_2230,N_1736,N_1588);
and U2231 (N_2231,N_1113,N_1999);
and U2232 (N_2232,N_1018,N_1816);
and U2233 (N_2233,N_1099,N_1957);
or U2234 (N_2234,N_1651,N_1749);
xnor U2235 (N_2235,N_1550,N_1690);
nor U2236 (N_2236,N_1115,N_1135);
or U2237 (N_2237,N_1134,N_1254);
xor U2238 (N_2238,N_1529,N_1908);
nor U2239 (N_2239,N_1268,N_1435);
nand U2240 (N_2240,N_1428,N_1088);
nor U2241 (N_2241,N_1813,N_1471);
and U2242 (N_2242,N_1350,N_1936);
nor U2243 (N_2243,N_1152,N_1706);
or U2244 (N_2244,N_1518,N_1286);
or U2245 (N_2245,N_1963,N_1234);
nor U2246 (N_2246,N_1288,N_1200);
nand U2247 (N_2247,N_1822,N_1804);
and U2248 (N_2248,N_1616,N_1329);
nor U2249 (N_2249,N_1833,N_1481);
and U2250 (N_2250,N_1081,N_1096);
and U2251 (N_2251,N_1293,N_1421);
xnor U2252 (N_2252,N_1709,N_1414);
or U2253 (N_2253,N_1055,N_1561);
nor U2254 (N_2254,N_1869,N_1366);
or U2255 (N_2255,N_1189,N_1947);
xor U2256 (N_2256,N_1795,N_1921);
nor U2257 (N_2257,N_1912,N_1244);
xor U2258 (N_2258,N_1433,N_1631);
and U2259 (N_2259,N_1566,N_1482);
nand U2260 (N_2260,N_1043,N_1837);
nand U2261 (N_2261,N_1221,N_1237);
and U2262 (N_2262,N_1760,N_1770);
or U2263 (N_2263,N_1093,N_1232);
or U2264 (N_2264,N_1543,N_1916);
nor U2265 (N_2265,N_1013,N_1608);
nand U2266 (N_2266,N_1872,N_1565);
nand U2267 (N_2267,N_1528,N_1213);
nor U2268 (N_2268,N_1504,N_1045);
or U2269 (N_2269,N_1448,N_1925);
and U2270 (N_2270,N_1035,N_1220);
nand U2271 (N_2271,N_1332,N_1443);
or U2272 (N_2272,N_1794,N_1502);
nor U2273 (N_2273,N_1402,N_1879);
xnor U2274 (N_2274,N_1865,N_1583);
nand U2275 (N_2275,N_1512,N_1164);
and U2276 (N_2276,N_1490,N_1218);
and U2277 (N_2277,N_1201,N_1934);
and U2278 (N_2278,N_1601,N_1519);
nand U2279 (N_2279,N_1829,N_1849);
nand U2280 (N_2280,N_1798,N_1488);
or U2281 (N_2281,N_1341,N_1971);
xnor U2282 (N_2282,N_1318,N_1339);
and U2283 (N_2283,N_1508,N_1520);
or U2284 (N_2284,N_1008,N_1896);
nand U2285 (N_2285,N_1904,N_1024);
and U2286 (N_2286,N_1319,N_1722);
nand U2287 (N_2287,N_1100,N_1282);
xor U2288 (N_2288,N_1525,N_1340);
nor U2289 (N_2289,N_1418,N_1961);
and U2290 (N_2290,N_1312,N_1489);
nand U2291 (N_2291,N_1165,N_1781);
nor U2292 (N_2292,N_1635,N_1967);
and U2293 (N_2293,N_1864,N_1632);
or U2294 (N_2294,N_1808,N_1299);
nand U2295 (N_2295,N_1970,N_1025);
nand U2296 (N_2296,N_1248,N_1762);
or U2297 (N_2297,N_1599,N_1721);
nor U2298 (N_2298,N_1571,N_1000);
xnor U2299 (N_2299,N_1219,N_1082);
nor U2300 (N_2300,N_1746,N_1977);
nor U2301 (N_2301,N_1618,N_1650);
nand U2302 (N_2302,N_1742,N_1346);
nand U2303 (N_2303,N_1447,N_1727);
or U2304 (N_2304,N_1823,N_1409);
nor U2305 (N_2305,N_1975,N_1054);
nor U2306 (N_2306,N_1337,N_1713);
xnor U2307 (N_2307,N_1882,N_1446);
or U2308 (N_2308,N_1812,N_1761);
nor U2309 (N_2309,N_1128,N_1107);
xnor U2310 (N_2310,N_1900,N_1938);
and U2311 (N_2311,N_1717,N_1814);
and U2312 (N_2312,N_1968,N_1142);
and U2313 (N_2313,N_1610,N_1225);
nand U2314 (N_2314,N_1419,N_1898);
nor U2315 (N_2315,N_1397,N_1307);
and U2316 (N_2316,N_1542,N_1669);
and U2317 (N_2317,N_1665,N_1716);
and U2318 (N_2318,N_1720,N_1776);
nor U2319 (N_2319,N_1740,N_1150);
nor U2320 (N_2320,N_1874,N_1133);
nand U2321 (N_2321,N_1396,N_1384);
nor U2322 (N_2322,N_1417,N_1051);
nor U2323 (N_2323,N_1014,N_1592);
nor U2324 (N_2324,N_1540,N_1076);
nand U2325 (N_2325,N_1911,N_1053);
or U2326 (N_2326,N_1942,N_1383);
and U2327 (N_2327,N_1202,N_1862);
and U2328 (N_2328,N_1595,N_1270);
nand U2329 (N_2329,N_1389,N_1410);
xnor U2330 (N_2330,N_1948,N_1123);
and U2331 (N_2331,N_1246,N_1069);
nand U2332 (N_2332,N_1580,N_1626);
and U2333 (N_2333,N_1995,N_1012);
nand U2334 (N_2334,N_1639,N_1223);
nor U2335 (N_2335,N_1617,N_1774);
nand U2336 (N_2336,N_1807,N_1815);
nand U2337 (N_2337,N_1479,N_1703);
nor U2338 (N_2338,N_1320,N_1049);
nand U2339 (N_2339,N_1753,N_1298);
nand U2340 (N_2340,N_1087,N_1766);
nor U2341 (N_2341,N_1105,N_1362);
nor U2342 (N_2342,N_1771,N_1469);
and U2343 (N_2343,N_1574,N_1343);
xor U2344 (N_2344,N_1805,N_1040);
and U2345 (N_2345,N_1400,N_1684);
nand U2346 (N_2346,N_1554,N_1817);
and U2347 (N_2347,N_1158,N_1715);
or U2348 (N_2348,N_1044,N_1847);
nor U2349 (N_2349,N_1539,N_1499);
or U2350 (N_2350,N_1647,N_1711);
or U2351 (N_2351,N_1352,N_1614);
nor U2352 (N_2352,N_1523,N_1751);
nor U2353 (N_2353,N_1591,N_1584);
xnor U2354 (N_2354,N_1131,N_1118);
nor U2355 (N_2355,N_1732,N_1831);
or U2356 (N_2356,N_1251,N_1116);
nand U2357 (N_2357,N_1112,N_1589);
or U2358 (N_2358,N_1415,N_1667);
or U2359 (N_2359,N_1291,N_1323);
and U2360 (N_2360,N_1461,N_1731);
nor U2361 (N_2361,N_1083,N_1136);
nand U2362 (N_2362,N_1381,N_1274);
nand U2363 (N_2363,N_1129,N_1922);
and U2364 (N_2364,N_1265,N_1998);
or U2365 (N_2365,N_1843,N_1186);
or U2366 (N_2366,N_1892,N_1906);
xnor U2367 (N_2367,N_1551,N_1547);
or U2368 (N_2368,N_1656,N_1702);
nand U2369 (N_2369,N_1856,N_1451);
nand U2370 (N_2370,N_1544,N_1303);
nand U2371 (N_2371,N_1311,N_1281);
and U2372 (N_2372,N_1440,N_1950);
or U2373 (N_2373,N_1072,N_1470);
nor U2374 (N_2374,N_1476,N_1450);
nor U2375 (N_2375,N_1273,N_1840);
xor U2376 (N_2376,N_1730,N_1132);
and U2377 (N_2377,N_1743,N_1183);
nor U2378 (N_2378,N_1073,N_1464);
xor U2379 (N_2379,N_1266,N_1797);
nor U2380 (N_2380,N_1871,N_1408);
and U2381 (N_2381,N_1261,N_1960);
xor U2382 (N_2382,N_1023,N_1953);
nor U2383 (N_2383,N_1090,N_1347);
or U2384 (N_2384,N_1905,N_1929);
xnor U2385 (N_2385,N_1784,N_1741);
nand U2386 (N_2386,N_1494,N_1068);
nor U2387 (N_2387,N_1524,N_1242);
nand U2388 (N_2388,N_1927,N_1596);
or U2389 (N_2389,N_1787,N_1227);
xnor U2390 (N_2390,N_1752,N_1306);
nor U2391 (N_2391,N_1515,N_1117);
or U2392 (N_2392,N_1498,N_1621);
nand U2393 (N_2393,N_1465,N_1991);
or U2394 (N_2394,N_1357,N_1138);
nand U2395 (N_2395,N_1037,N_1149);
nand U2396 (N_2396,N_1842,N_1887);
nor U2397 (N_2397,N_1328,N_1895);
and U2398 (N_2398,N_1296,N_1314);
and U2399 (N_2399,N_1467,N_1484);
xor U2400 (N_2400,N_1172,N_1308);
or U2401 (N_2401,N_1376,N_1240);
xor U2402 (N_2402,N_1556,N_1033);
nand U2403 (N_2403,N_1041,N_1078);
nor U2404 (N_2404,N_1065,N_1516);
nor U2405 (N_2405,N_1373,N_1965);
or U2406 (N_2406,N_1160,N_1336);
and U2407 (N_2407,N_1707,N_1007);
xnor U2408 (N_2408,N_1403,N_1578);
nor U2409 (N_2409,N_1155,N_1750);
or U2410 (N_2410,N_1689,N_1792);
or U2411 (N_2411,N_1511,N_1258);
and U2412 (N_2412,N_1153,N_1157);
nor U2413 (N_2413,N_1655,N_1951);
xnor U2414 (N_2414,N_1939,N_1984);
or U2415 (N_2415,N_1301,N_1568);
and U2416 (N_2416,N_1333,N_1167);
or U2417 (N_2417,N_1317,N_1108);
nor U2418 (N_2418,N_1364,N_1538);
nand U2419 (N_2419,N_1486,N_1349);
nand U2420 (N_2420,N_1719,N_1772);
and U2421 (N_2421,N_1883,N_1966);
or U2422 (N_2422,N_1825,N_1558);
nand U2423 (N_2423,N_1852,N_1573);
xor U2424 (N_2424,N_1269,N_1704);
and U2425 (N_2425,N_1956,N_1629);
or U2426 (N_2426,N_1861,N_1782);
nand U2427 (N_2427,N_1216,N_1374);
or U2428 (N_2428,N_1778,N_1899);
and U2429 (N_2429,N_1416,N_1368);
nor U2430 (N_2430,N_1257,N_1735);
nor U2431 (N_2431,N_1579,N_1394);
nor U2432 (N_2432,N_1654,N_1058);
nor U2433 (N_2433,N_1758,N_1020);
xor U2434 (N_2434,N_1726,N_1267);
nand U2435 (N_2435,N_1531,N_1046);
xnor U2436 (N_2436,N_1260,N_1636);
or U2437 (N_2437,N_1955,N_1612);
nand U2438 (N_2438,N_1492,N_1836);
and U2439 (N_2439,N_1348,N_1718);
nor U2440 (N_2440,N_1763,N_1980);
nand U2441 (N_2441,N_1788,N_1454);
and U2442 (N_2442,N_1915,N_1708);
or U2443 (N_2443,N_1853,N_1983);
xor U2444 (N_2444,N_1724,N_1460);
or U2445 (N_2445,N_1122,N_1903);
nand U2446 (N_2446,N_1824,N_1826);
nand U2447 (N_2447,N_1250,N_1943);
nor U2448 (N_2448,N_1459,N_1755);
nor U2449 (N_2449,N_1173,N_1477);
or U2450 (N_2450,N_1863,N_1196);
nor U2451 (N_2451,N_1487,N_1530);
nand U2452 (N_2452,N_1687,N_1828);
nor U2453 (N_2453,N_1695,N_1994);
or U2454 (N_2454,N_1692,N_1175);
nand U2455 (N_2455,N_1756,N_1894);
or U2456 (N_2456,N_1546,N_1185);
nor U2457 (N_2457,N_1207,N_1637);
and U2458 (N_2458,N_1365,N_1835);
nand U2459 (N_2459,N_1567,N_1880);
or U2460 (N_2460,N_1924,N_1675);
nor U2461 (N_2461,N_1745,N_1888);
nor U2462 (N_2462,N_1868,N_1480);
or U2463 (N_2463,N_1884,N_1920);
and U2464 (N_2464,N_1247,N_1056);
or U2465 (N_2465,N_1866,N_1005);
and U2466 (N_2466,N_1931,N_1278);
and U2467 (N_2467,N_1535,N_1009);
xnor U2468 (N_2468,N_1679,N_1769);
nor U2469 (N_2469,N_1909,N_1019);
nor U2470 (N_2470,N_1139,N_1553);
or U2471 (N_2471,N_1607,N_1738);
nor U2472 (N_2472,N_1633,N_1534);
or U2473 (N_2473,N_1478,N_1474);
nor U2474 (N_2474,N_1973,N_1316);
nand U2475 (N_2475,N_1371,N_1255);
and U2476 (N_2476,N_1959,N_1932);
or U2477 (N_2477,N_1032,N_1422);
or U2478 (N_2478,N_1800,N_1468);
or U2479 (N_2479,N_1360,N_1004);
nand U2480 (N_2480,N_1354,N_1693);
or U2481 (N_2481,N_1377,N_1199);
nand U2482 (N_2482,N_1027,N_1259);
nor U2483 (N_2483,N_1670,N_1441);
or U2484 (N_2484,N_1602,N_1649);
nor U2485 (N_2485,N_1204,N_1801);
nand U2486 (N_2486,N_1613,N_1085);
and U2487 (N_2487,N_1159,N_1401);
nand U2488 (N_2488,N_1641,N_1918);
or U2489 (N_2489,N_1928,N_1850);
and U2490 (N_2490,N_1768,N_1280);
or U2491 (N_2491,N_1640,N_1434);
nor U2492 (N_2492,N_1681,N_1802);
and U2493 (N_2493,N_1275,N_1326);
nand U2494 (N_2494,N_1796,N_1457);
nand U2495 (N_2495,N_1002,N_1619);
nor U2496 (N_2496,N_1563,N_1442);
and U2497 (N_2497,N_1052,N_1212);
and U2498 (N_2498,N_1773,N_1545);
and U2499 (N_2499,N_1777,N_1791);
xor U2500 (N_2500,N_1315,N_1613);
nor U2501 (N_2501,N_1423,N_1679);
or U2502 (N_2502,N_1759,N_1833);
and U2503 (N_2503,N_1322,N_1586);
nand U2504 (N_2504,N_1401,N_1487);
nand U2505 (N_2505,N_1653,N_1359);
and U2506 (N_2506,N_1563,N_1477);
or U2507 (N_2507,N_1755,N_1645);
and U2508 (N_2508,N_1725,N_1233);
and U2509 (N_2509,N_1853,N_1344);
nand U2510 (N_2510,N_1112,N_1610);
nand U2511 (N_2511,N_1162,N_1071);
nand U2512 (N_2512,N_1102,N_1437);
or U2513 (N_2513,N_1949,N_1956);
nor U2514 (N_2514,N_1871,N_1499);
nand U2515 (N_2515,N_1831,N_1652);
nand U2516 (N_2516,N_1194,N_1416);
nand U2517 (N_2517,N_1317,N_1559);
or U2518 (N_2518,N_1273,N_1288);
or U2519 (N_2519,N_1898,N_1314);
or U2520 (N_2520,N_1451,N_1903);
or U2521 (N_2521,N_1596,N_1705);
and U2522 (N_2522,N_1493,N_1739);
nor U2523 (N_2523,N_1886,N_1618);
nand U2524 (N_2524,N_1681,N_1408);
nand U2525 (N_2525,N_1603,N_1238);
nand U2526 (N_2526,N_1465,N_1778);
or U2527 (N_2527,N_1086,N_1336);
and U2528 (N_2528,N_1222,N_1490);
or U2529 (N_2529,N_1871,N_1232);
nor U2530 (N_2530,N_1101,N_1465);
and U2531 (N_2531,N_1101,N_1614);
nor U2532 (N_2532,N_1879,N_1356);
xor U2533 (N_2533,N_1650,N_1291);
and U2534 (N_2534,N_1706,N_1279);
nor U2535 (N_2535,N_1901,N_1147);
and U2536 (N_2536,N_1379,N_1177);
and U2537 (N_2537,N_1706,N_1864);
and U2538 (N_2538,N_1564,N_1916);
nor U2539 (N_2539,N_1915,N_1416);
nand U2540 (N_2540,N_1766,N_1117);
xnor U2541 (N_2541,N_1992,N_1663);
nand U2542 (N_2542,N_1045,N_1972);
or U2543 (N_2543,N_1962,N_1564);
or U2544 (N_2544,N_1599,N_1712);
nor U2545 (N_2545,N_1284,N_1894);
nand U2546 (N_2546,N_1843,N_1543);
and U2547 (N_2547,N_1180,N_1356);
nor U2548 (N_2548,N_1226,N_1827);
and U2549 (N_2549,N_1788,N_1443);
or U2550 (N_2550,N_1658,N_1933);
or U2551 (N_2551,N_1606,N_1392);
or U2552 (N_2552,N_1331,N_1427);
and U2553 (N_2553,N_1108,N_1436);
nor U2554 (N_2554,N_1306,N_1996);
nand U2555 (N_2555,N_1411,N_1124);
nand U2556 (N_2556,N_1584,N_1774);
or U2557 (N_2557,N_1012,N_1646);
nor U2558 (N_2558,N_1632,N_1886);
or U2559 (N_2559,N_1042,N_1572);
nand U2560 (N_2560,N_1502,N_1714);
or U2561 (N_2561,N_1591,N_1206);
nor U2562 (N_2562,N_1059,N_1946);
and U2563 (N_2563,N_1441,N_1474);
xnor U2564 (N_2564,N_1270,N_1204);
and U2565 (N_2565,N_1755,N_1679);
and U2566 (N_2566,N_1248,N_1887);
nor U2567 (N_2567,N_1566,N_1152);
nand U2568 (N_2568,N_1308,N_1291);
nor U2569 (N_2569,N_1384,N_1711);
and U2570 (N_2570,N_1751,N_1504);
or U2571 (N_2571,N_1784,N_1400);
or U2572 (N_2572,N_1052,N_1993);
nand U2573 (N_2573,N_1102,N_1622);
and U2574 (N_2574,N_1310,N_1744);
nor U2575 (N_2575,N_1873,N_1545);
nand U2576 (N_2576,N_1947,N_1704);
and U2577 (N_2577,N_1967,N_1090);
and U2578 (N_2578,N_1490,N_1522);
nor U2579 (N_2579,N_1055,N_1316);
xor U2580 (N_2580,N_1502,N_1649);
and U2581 (N_2581,N_1396,N_1597);
and U2582 (N_2582,N_1543,N_1966);
and U2583 (N_2583,N_1336,N_1027);
or U2584 (N_2584,N_1469,N_1763);
or U2585 (N_2585,N_1587,N_1971);
nand U2586 (N_2586,N_1317,N_1562);
nor U2587 (N_2587,N_1369,N_1562);
nand U2588 (N_2588,N_1949,N_1637);
and U2589 (N_2589,N_1558,N_1749);
or U2590 (N_2590,N_1213,N_1482);
nand U2591 (N_2591,N_1283,N_1811);
and U2592 (N_2592,N_1269,N_1732);
nand U2593 (N_2593,N_1881,N_1084);
nor U2594 (N_2594,N_1685,N_1428);
or U2595 (N_2595,N_1199,N_1674);
nor U2596 (N_2596,N_1444,N_1228);
nand U2597 (N_2597,N_1659,N_1711);
nor U2598 (N_2598,N_1259,N_1665);
nand U2599 (N_2599,N_1683,N_1533);
nand U2600 (N_2600,N_1948,N_1337);
nor U2601 (N_2601,N_1991,N_1696);
and U2602 (N_2602,N_1000,N_1860);
and U2603 (N_2603,N_1028,N_1765);
or U2604 (N_2604,N_1189,N_1262);
or U2605 (N_2605,N_1441,N_1066);
and U2606 (N_2606,N_1957,N_1661);
xnor U2607 (N_2607,N_1582,N_1976);
nor U2608 (N_2608,N_1394,N_1276);
nand U2609 (N_2609,N_1399,N_1785);
and U2610 (N_2610,N_1534,N_1720);
nand U2611 (N_2611,N_1176,N_1435);
xnor U2612 (N_2612,N_1093,N_1524);
and U2613 (N_2613,N_1103,N_1707);
or U2614 (N_2614,N_1445,N_1088);
nand U2615 (N_2615,N_1822,N_1151);
nand U2616 (N_2616,N_1950,N_1463);
nand U2617 (N_2617,N_1974,N_1782);
nor U2618 (N_2618,N_1761,N_1902);
xnor U2619 (N_2619,N_1256,N_1282);
or U2620 (N_2620,N_1886,N_1696);
or U2621 (N_2621,N_1308,N_1809);
xnor U2622 (N_2622,N_1869,N_1987);
or U2623 (N_2623,N_1466,N_1335);
and U2624 (N_2624,N_1533,N_1526);
xor U2625 (N_2625,N_1891,N_1649);
or U2626 (N_2626,N_1760,N_1599);
or U2627 (N_2627,N_1894,N_1916);
nand U2628 (N_2628,N_1199,N_1852);
nand U2629 (N_2629,N_1580,N_1320);
and U2630 (N_2630,N_1240,N_1550);
nor U2631 (N_2631,N_1625,N_1370);
or U2632 (N_2632,N_1775,N_1250);
or U2633 (N_2633,N_1682,N_1283);
nand U2634 (N_2634,N_1973,N_1618);
and U2635 (N_2635,N_1438,N_1223);
nor U2636 (N_2636,N_1093,N_1307);
and U2637 (N_2637,N_1876,N_1573);
nand U2638 (N_2638,N_1114,N_1153);
nor U2639 (N_2639,N_1966,N_1222);
nand U2640 (N_2640,N_1447,N_1170);
nor U2641 (N_2641,N_1841,N_1021);
nor U2642 (N_2642,N_1063,N_1436);
nand U2643 (N_2643,N_1597,N_1783);
xnor U2644 (N_2644,N_1105,N_1884);
or U2645 (N_2645,N_1925,N_1701);
or U2646 (N_2646,N_1318,N_1827);
and U2647 (N_2647,N_1415,N_1120);
and U2648 (N_2648,N_1162,N_1881);
nor U2649 (N_2649,N_1429,N_1377);
and U2650 (N_2650,N_1073,N_1588);
nand U2651 (N_2651,N_1020,N_1202);
and U2652 (N_2652,N_1848,N_1364);
xor U2653 (N_2653,N_1405,N_1300);
and U2654 (N_2654,N_1256,N_1090);
nand U2655 (N_2655,N_1803,N_1549);
nor U2656 (N_2656,N_1071,N_1124);
or U2657 (N_2657,N_1679,N_1190);
or U2658 (N_2658,N_1457,N_1139);
nand U2659 (N_2659,N_1370,N_1066);
nand U2660 (N_2660,N_1940,N_1479);
nand U2661 (N_2661,N_1835,N_1269);
nand U2662 (N_2662,N_1942,N_1803);
nand U2663 (N_2663,N_1684,N_1585);
or U2664 (N_2664,N_1010,N_1735);
or U2665 (N_2665,N_1091,N_1987);
nand U2666 (N_2666,N_1411,N_1792);
or U2667 (N_2667,N_1105,N_1667);
and U2668 (N_2668,N_1003,N_1752);
and U2669 (N_2669,N_1468,N_1065);
nand U2670 (N_2670,N_1193,N_1392);
or U2671 (N_2671,N_1685,N_1521);
nor U2672 (N_2672,N_1505,N_1948);
nor U2673 (N_2673,N_1028,N_1900);
and U2674 (N_2674,N_1736,N_1795);
and U2675 (N_2675,N_1174,N_1992);
or U2676 (N_2676,N_1628,N_1849);
or U2677 (N_2677,N_1885,N_1666);
or U2678 (N_2678,N_1973,N_1564);
nor U2679 (N_2679,N_1971,N_1724);
or U2680 (N_2680,N_1183,N_1522);
or U2681 (N_2681,N_1002,N_1133);
xnor U2682 (N_2682,N_1887,N_1316);
nor U2683 (N_2683,N_1105,N_1816);
nand U2684 (N_2684,N_1569,N_1174);
nand U2685 (N_2685,N_1958,N_1792);
or U2686 (N_2686,N_1023,N_1297);
xor U2687 (N_2687,N_1887,N_1151);
nand U2688 (N_2688,N_1563,N_1525);
or U2689 (N_2689,N_1716,N_1274);
nand U2690 (N_2690,N_1154,N_1465);
and U2691 (N_2691,N_1671,N_1839);
nand U2692 (N_2692,N_1275,N_1858);
nand U2693 (N_2693,N_1813,N_1363);
or U2694 (N_2694,N_1872,N_1360);
nand U2695 (N_2695,N_1388,N_1762);
nor U2696 (N_2696,N_1552,N_1497);
nor U2697 (N_2697,N_1204,N_1761);
nand U2698 (N_2698,N_1133,N_1415);
nor U2699 (N_2699,N_1936,N_1355);
xor U2700 (N_2700,N_1266,N_1669);
nor U2701 (N_2701,N_1496,N_1344);
or U2702 (N_2702,N_1426,N_1399);
or U2703 (N_2703,N_1547,N_1069);
or U2704 (N_2704,N_1834,N_1936);
and U2705 (N_2705,N_1073,N_1171);
or U2706 (N_2706,N_1505,N_1603);
nand U2707 (N_2707,N_1803,N_1396);
and U2708 (N_2708,N_1491,N_1830);
and U2709 (N_2709,N_1009,N_1493);
or U2710 (N_2710,N_1216,N_1807);
or U2711 (N_2711,N_1613,N_1563);
xor U2712 (N_2712,N_1148,N_1198);
or U2713 (N_2713,N_1939,N_1629);
nor U2714 (N_2714,N_1244,N_1516);
or U2715 (N_2715,N_1074,N_1197);
or U2716 (N_2716,N_1089,N_1636);
xnor U2717 (N_2717,N_1636,N_1190);
and U2718 (N_2718,N_1571,N_1956);
nand U2719 (N_2719,N_1097,N_1179);
nand U2720 (N_2720,N_1220,N_1008);
xnor U2721 (N_2721,N_1679,N_1341);
or U2722 (N_2722,N_1695,N_1908);
nand U2723 (N_2723,N_1400,N_1644);
and U2724 (N_2724,N_1562,N_1709);
nor U2725 (N_2725,N_1331,N_1928);
and U2726 (N_2726,N_1944,N_1730);
nand U2727 (N_2727,N_1096,N_1257);
nor U2728 (N_2728,N_1344,N_1324);
and U2729 (N_2729,N_1968,N_1953);
nand U2730 (N_2730,N_1880,N_1106);
and U2731 (N_2731,N_1816,N_1802);
nand U2732 (N_2732,N_1696,N_1256);
and U2733 (N_2733,N_1506,N_1894);
and U2734 (N_2734,N_1427,N_1584);
and U2735 (N_2735,N_1016,N_1928);
and U2736 (N_2736,N_1026,N_1923);
nor U2737 (N_2737,N_1511,N_1796);
nor U2738 (N_2738,N_1729,N_1163);
and U2739 (N_2739,N_1586,N_1319);
nor U2740 (N_2740,N_1513,N_1677);
or U2741 (N_2741,N_1113,N_1543);
or U2742 (N_2742,N_1024,N_1970);
nand U2743 (N_2743,N_1928,N_1761);
or U2744 (N_2744,N_1633,N_1483);
and U2745 (N_2745,N_1556,N_1772);
or U2746 (N_2746,N_1723,N_1072);
nor U2747 (N_2747,N_1935,N_1642);
and U2748 (N_2748,N_1517,N_1955);
and U2749 (N_2749,N_1036,N_1089);
nand U2750 (N_2750,N_1954,N_1255);
nand U2751 (N_2751,N_1458,N_1667);
and U2752 (N_2752,N_1433,N_1125);
or U2753 (N_2753,N_1324,N_1281);
xor U2754 (N_2754,N_1476,N_1603);
or U2755 (N_2755,N_1057,N_1242);
nor U2756 (N_2756,N_1375,N_1784);
and U2757 (N_2757,N_1013,N_1463);
and U2758 (N_2758,N_1510,N_1058);
nand U2759 (N_2759,N_1178,N_1209);
nand U2760 (N_2760,N_1683,N_1925);
nor U2761 (N_2761,N_1378,N_1674);
and U2762 (N_2762,N_1434,N_1754);
and U2763 (N_2763,N_1517,N_1133);
nor U2764 (N_2764,N_1954,N_1400);
xnor U2765 (N_2765,N_1518,N_1419);
or U2766 (N_2766,N_1867,N_1467);
and U2767 (N_2767,N_1915,N_1143);
and U2768 (N_2768,N_1648,N_1108);
xor U2769 (N_2769,N_1314,N_1599);
or U2770 (N_2770,N_1606,N_1851);
nand U2771 (N_2771,N_1914,N_1124);
or U2772 (N_2772,N_1957,N_1870);
nand U2773 (N_2773,N_1106,N_1462);
or U2774 (N_2774,N_1006,N_1866);
nand U2775 (N_2775,N_1346,N_1584);
xor U2776 (N_2776,N_1082,N_1791);
or U2777 (N_2777,N_1874,N_1393);
nand U2778 (N_2778,N_1867,N_1121);
and U2779 (N_2779,N_1651,N_1160);
or U2780 (N_2780,N_1683,N_1530);
nor U2781 (N_2781,N_1372,N_1796);
nand U2782 (N_2782,N_1647,N_1263);
nand U2783 (N_2783,N_1303,N_1774);
and U2784 (N_2784,N_1726,N_1840);
xnor U2785 (N_2785,N_1354,N_1837);
and U2786 (N_2786,N_1710,N_1170);
nand U2787 (N_2787,N_1756,N_1105);
nand U2788 (N_2788,N_1434,N_1719);
nand U2789 (N_2789,N_1364,N_1466);
or U2790 (N_2790,N_1568,N_1428);
nand U2791 (N_2791,N_1900,N_1870);
nand U2792 (N_2792,N_1870,N_1973);
nor U2793 (N_2793,N_1042,N_1894);
and U2794 (N_2794,N_1171,N_1781);
nand U2795 (N_2795,N_1480,N_1578);
or U2796 (N_2796,N_1637,N_1478);
and U2797 (N_2797,N_1263,N_1915);
nand U2798 (N_2798,N_1944,N_1579);
nor U2799 (N_2799,N_1013,N_1934);
and U2800 (N_2800,N_1018,N_1121);
and U2801 (N_2801,N_1378,N_1635);
nand U2802 (N_2802,N_1211,N_1505);
nor U2803 (N_2803,N_1756,N_1552);
and U2804 (N_2804,N_1442,N_1691);
and U2805 (N_2805,N_1078,N_1430);
nor U2806 (N_2806,N_1109,N_1453);
and U2807 (N_2807,N_1612,N_1057);
or U2808 (N_2808,N_1512,N_1400);
nand U2809 (N_2809,N_1048,N_1830);
nand U2810 (N_2810,N_1659,N_1383);
and U2811 (N_2811,N_1064,N_1185);
or U2812 (N_2812,N_1150,N_1224);
or U2813 (N_2813,N_1914,N_1983);
nor U2814 (N_2814,N_1795,N_1882);
nand U2815 (N_2815,N_1942,N_1655);
or U2816 (N_2816,N_1623,N_1669);
or U2817 (N_2817,N_1226,N_1926);
or U2818 (N_2818,N_1163,N_1990);
nand U2819 (N_2819,N_1268,N_1753);
nor U2820 (N_2820,N_1003,N_1952);
or U2821 (N_2821,N_1121,N_1620);
and U2822 (N_2822,N_1405,N_1524);
nor U2823 (N_2823,N_1524,N_1840);
nand U2824 (N_2824,N_1916,N_1771);
and U2825 (N_2825,N_1525,N_1186);
and U2826 (N_2826,N_1955,N_1130);
nor U2827 (N_2827,N_1525,N_1782);
xnor U2828 (N_2828,N_1779,N_1850);
nand U2829 (N_2829,N_1777,N_1257);
xor U2830 (N_2830,N_1332,N_1886);
xnor U2831 (N_2831,N_1436,N_1374);
nor U2832 (N_2832,N_1685,N_1067);
and U2833 (N_2833,N_1692,N_1580);
or U2834 (N_2834,N_1846,N_1536);
nor U2835 (N_2835,N_1206,N_1638);
or U2836 (N_2836,N_1243,N_1625);
and U2837 (N_2837,N_1633,N_1882);
nor U2838 (N_2838,N_1919,N_1510);
and U2839 (N_2839,N_1949,N_1621);
or U2840 (N_2840,N_1223,N_1600);
or U2841 (N_2841,N_1695,N_1002);
and U2842 (N_2842,N_1042,N_1332);
nor U2843 (N_2843,N_1687,N_1715);
or U2844 (N_2844,N_1027,N_1477);
and U2845 (N_2845,N_1002,N_1513);
xor U2846 (N_2846,N_1820,N_1437);
or U2847 (N_2847,N_1510,N_1079);
or U2848 (N_2848,N_1480,N_1961);
and U2849 (N_2849,N_1850,N_1605);
or U2850 (N_2850,N_1328,N_1733);
nor U2851 (N_2851,N_1732,N_1778);
nor U2852 (N_2852,N_1931,N_1108);
nand U2853 (N_2853,N_1712,N_1681);
or U2854 (N_2854,N_1390,N_1900);
or U2855 (N_2855,N_1640,N_1364);
nand U2856 (N_2856,N_1473,N_1924);
and U2857 (N_2857,N_1898,N_1090);
xor U2858 (N_2858,N_1306,N_1929);
and U2859 (N_2859,N_1005,N_1512);
nor U2860 (N_2860,N_1160,N_1672);
xnor U2861 (N_2861,N_1599,N_1423);
nor U2862 (N_2862,N_1501,N_1865);
and U2863 (N_2863,N_1126,N_1325);
xnor U2864 (N_2864,N_1166,N_1879);
and U2865 (N_2865,N_1408,N_1643);
and U2866 (N_2866,N_1350,N_1076);
nor U2867 (N_2867,N_1523,N_1194);
nand U2868 (N_2868,N_1876,N_1483);
and U2869 (N_2869,N_1303,N_1912);
and U2870 (N_2870,N_1194,N_1764);
or U2871 (N_2871,N_1815,N_1539);
nor U2872 (N_2872,N_1199,N_1302);
or U2873 (N_2873,N_1612,N_1903);
nand U2874 (N_2874,N_1841,N_1915);
or U2875 (N_2875,N_1195,N_1562);
and U2876 (N_2876,N_1339,N_1557);
nor U2877 (N_2877,N_1625,N_1753);
nand U2878 (N_2878,N_1002,N_1401);
nand U2879 (N_2879,N_1562,N_1497);
or U2880 (N_2880,N_1259,N_1785);
nor U2881 (N_2881,N_1749,N_1596);
and U2882 (N_2882,N_1983,N_1273);
nor U2883 (N_2883,N_1046,N_1247);
or U2884 (N_2884,N_1613,N_1369);
nor U2885 (N_2885,N_1508,N_1751);
and U2886 (N_2886,N_1699,N_1994);
nand U2887 (N_2887,N_1536,N_1857);
nor U2888 (N_2888,N_1763,N_1096);
nand U2889 (N_2889,N_1875,N_1923);
or U2890 (N_2890,N_1391,N_1769);
or U2891 (N_2891,N_1329,N_1170);
or U2892 (N_2892,N_1825,N_1980);
or U2893 (N_2893,N_1348,N_1675);
and U2894 (N_2894,N_1399,N_1950);
nand U2895 (N_2895,N_1022,N_1143);
or U2896 (N_2896,N_1632,N_1553);
nand U2897 (N_2897,N_1554,N_1704);
and U2898 (N_2898,N_1119,N_1410);
nor U2899 (N_2899,N_1397,N_1489);
nand U2900 (N_2900,N_1540,N_1688);
xnor U2901 (N_2901,N_1171,N_1558);
xnor U2902 (N_2902,N_1357,N_1681);
or U2903 (N_2903,N_1869,N_1854);
and U2904 (N_2904,N_1145,N_1236);
or U2905 (N_2905,N_1879,N_1287);
xor U2906 (N_2906,N_1673,N_1119);
nor U2907 (N_2907,N_1855,N_1465);
or U2908 (N_2908,N_1351,N_1868);
nand U2909 (N_2909,N_1559,N_1429);
nor U2910 (N_2910,N_1002,N_1164);
xnor U2911 (N_2911,N_1426,N_1984);
and U2912 (N_2912,N_1146,N_1734);
nand U2913 (N_2913,N_1634,N_1753);
xnor U2914 (N_2914,N_1597,N_1711);
nor U2915 (N_2915,N_1919,N_1568);
nor U2916 (N_2916,N_1268,N_1556);
nor U2917 (N_2917,N_1187,N_1407);
xnor U2918 (N_2918,N_1766,N_1892);
xor U2919 (N_2919,N_1049,N_1012);
nor U2920 (N_2920,N_1048,N_1597);
nor U2921 (N_2921,N_1703,N_1317);
xnor U2922 (N_2922,N_1175,N_1894);
nand U2923 (N_2923,N_1709,N_1993);
and U2924 (N_2924,N_1787,N_1446);
nor U2925 (N_2925,N_1499,N_1252);
and U2926 (N_2926,N_1183,N_1767);
nand U2927 (N_2927,N_1403,N_1050);
nor U2928 (N_2928,N_1116,N_1352);
nand U2929 (N_2929,N_1393,N_1537);
nand U2930 (N_2930,N_1870,N_1008);
or U2931 (N_2931,N_1841,N_1644);
xor U2932 (N_2932,N_1110,N_1407);
nor U2933 (N_2933,N_1314,N_1956);
or U2934 (N_2934,N_1709,N_1168);
nand U2935 (N_2935,N_1807,N_1962);
or U2936 (N_2936,N_1774,N_1562);
or U2937 (N_2937,N_1631,N_1017);
nand U2938 (N_2938,N_1480,N_1631);
or U2939 (N_2939,N_1948,N_1066);
and U2940 (N_2940,N_1178,N_1437);
nand U2941 (N_2941,N_1969,N_1925);
nand U2942 (N_2942,N_1698,N_1944);
or U2943 (N_2943,N_1546,N_1544);
and U2944 (N_2944,N_1494,N_1469);
nor U2945 (N_2945,N_1196,N_1223);
or U2946 (N_2946,N_1523,N_1673);
nor U2947 (N_2947,N_1017,N_1948);
and U2948 (N_2948,N_1295,N_1631);
and U2949 (N_2949,N_1310,N_1400);
nand U2950 (N_2950,N_1162,N_1143);
or U2951 (N_2951,N_1463,N_1331);
and U2952 (N_2952,N_1017,N_1417);
or U2953 (N_2953,N_1044,N_1270);
and U2954 (N_2954,N_1657,N_1534);
nor U2955 (N_2955,N_1947,N_1963);
xnor U2956 (N_2956,N_1594,N_1796);
nor U2957 (N_2957,N_1829,N_1787);
and U2958 (N_2958,N_1564,N_1509);
and U2959 (N_2959,N_1482,N_1908);
nor U2960 (N_2960,N_1672,N_1886);
nand U2961 (N_2961,N_1126,N_1390);
xor U2962 (N_2962,N_1219,N_1916);
and U2963 (N_2963,N_1021,N_1388);
nor U2964 (N_2964,N_1532,N_1723);
or U2965 (N_2965,N_1289,N_1828);
nor U2966 (N_2966,N_1203,N_1361);
and U2967 (N_2967,N_1507,N_1259);
and U2968 (N_2968,N_1430,N_1454);
xnor U2969 (N_2969,N_1900,N_1744);
and U2970 (N_2970,N_1808,N_1820);
or U2971 (N_2971,N_1679,N_1342);
or U2972 (N_2972,N_1796,N_1376);
and U2973 (N_2973,N_1871,N_1290);
or U2974 (N_2974,N_1972,N_1149);
nand U2975 (N_2975,N_1356,N_1504);
nor U2976 (N_2976,N_1389,N_1276);
xnor U2977 (N_2977,N_1362,N_1871);
xor U2978 (N_2978,N_1037,N_1000);
nor U2979 (N_2979,N_1050,N_1654);
nand U2980 (N_2980,N_1445,N_1172);
nand U2981 (N_2981,N_1948,N_1060);
and U2982 (N_2982,N_1356,N_1571);
and U2983 (N_2983,N_1013,N_1544);
nand U2984 (N_2984,N_1594,N_1739);
nand U2985 (N_2985,N_1242,N_1762);
or U2986 (N_2986,N_1972,N_1980);
nor U2987 (N_2987,N_1781,N_1581);
nand U2988 (N_2988,N_1551,N_1504);
or U2989 (N_2989,N_1589,N_1413);
and U2990 (N_2990,N_1318,N_1947);
or U2991 (N_2991,N_1030,N_1305);
nor U2992 (N_2992,N_1901,N_1602);
nor U2993 (N_2993,N_1583,N_1777);
nand U2994 (N_2994,N_1934,N_1260);
nor U2995 (N_2995,N_1628,N_1701);
nor U2996 (N_2996,N_1273,N_1565);
or U2997 (N_2997,N_1080,N_1374);
or U2998 (N_2998,N_1723,N_1236);
nand U2999 (N_2999,N_1100,N_1083);
nand U3000 (N_3000,N_2755,N_2999);
and U3001 (N_3001,N_2442,N_2491);
or U3002 (N_3002,N_2579,N_2238);
or U3003 (N_3003,N_2583,N_2688);
or U3004 (N_3004,N_2224,N_2675);
nor U3005 (N_3005,N_2048,N_2017);
xnor U3006 (N_3006,N_2361,N_2247);
nor U3007 (N_3007,N_2452,N_2082);
or U3008 (N_3008,N_2060,N_2058);
nor U3009 (N_3009,N_2584,N_2330);
nand U3010 (N_3010,N_2981,N_2418);
nor U3011 (N_3011,N_2037,N_2391);
nor U3012 (N_3012,N_2383,N_2648);
nand U3013 (N_3013,N_2784,N_2425);
and U3014 (N_3014,N_2997,N_2557);
or U3015 (N_3015,N_2823,N_2578);
and U3016 (N_3016,N_2947,N_2762);
and U3017 (N_3017,N_2940,N_2235);
and U3018 (N_3018,N_2560,N_2149);
nand U3019 (N_3019,N_2979,N_2427);
nand U3020 (N_3020,N_2128,N_2204);
or U3021 (N_3021,N_2931,N_2594);
or U3022 (N_3022,N_2745,N_2317);
nand U3023 (N_3023,N_2325,N_2370);
nand U3024 (N_3024,N_2776,N_2739);
nand U3025 (N_3025,N_2640,N_2661);
nand U3026 (N_3026,N_2857,N_2049);
and U3027 (N_3027,N_2988,N_2731);
and U3028 (N_3028,N_2041,N_2873);
nor U3029 (N_3029,N_2216,N_2712);
or U3030 (N_3030,N_2721,N_2405);
or U3031 (N_3031,N_2194,N_2708);
nor U3032 (N_3032,N_2530,N_2856);
nand U3033 (N_3033,N_2975,N_2005);
nand U3034 (N_3034,N_2769,N_2332);
or U3035 (N_3035,N_2923,N_2765);
nand U3036 (N_3036,N_2602,N_2348);
xor U3037 (N_3037,N_2547,N_2512);
and U3038 (N_3038,N_2394,N_2110);
nand U3039 (N_3039,N_2471,N_2057);
or U3040 (N_3040,N_2927,N_2502);
or U3041 (N_3041,N_2013,N_2496);
or U3042 (N_3042,N_2131,N_2482);
nand U3043 (N_3043,N_2672,N_2770);
nor U3044 (N_3044,N_2750,N_2633);
nor U3045 (N_3045,N_2662,N_2597);
or U3046 (N_3046,N_2229,N_2957);
or U3047 (N_3047,N_2282,N_2461);
or U3048 (N_3048,N_2123,N_2186);
xor U3049 (N_3049,N_2183,N_2531);
xnor U3050 (N_3050,N_2977,N_2117);
xnor U3051 (N_3051,N_2510,N_2347);
nor U3052 (N_3052,N_2505,N_2917);
or U3053 (N_3053,N_2278,N_2922);
nor U3054 (N_3054,N_2294,N_2012);
and U3055 (N_3055,N_2078,N_2953);
nand U3056 (N_3056,N_2837,N_2965);
xnor U3057 (N_3057,N_2038,N_2001);
nor U3058 (N_3058,N_2413,N_2937);
nand U3059 (N_3059,N_2824,N_2181);
and U3060 (N_3060,N_2213,N_2036);
nor U3061 (N_3061,N_2694,N_2220);
nand U3062 (N_3062,N_2946,N_2974);
nor U3063 (N_3063,N_2145,N_2929);
nand U3064 (N_3064,N_2820,N_2409);
nor U3065 (N_3065,N_2973,N_2870);
or U3066 (N_3066,N_2003,N_2114);
nand U3067 (N_3067,N_2958,N_2174);
or U3068 (N_3068,N_2139,N_2417);
nor U3069 (N_3069,N_2326,N_2443);
and U3070 (N_3070,N_2094,N_2787);
nor U3071 (N_3071,N_2788,N_2199);
or U3072 (N_3072,N_2901,N_2380);
nor U3073 (N_3073,N_2872,N_2832);
nand U3074 (N_3074,N_2351,N_2771);
nor U3075 (N_3075,N_2950,N_2172);
or U3076 (N_3076,N_2340,N_2867);
nor U3077 (N_3077,N_2156,N_2112);
nand U3078 (N_3078,N_2244,N_2140);
and U3079 (N_3079,N_2327,N_2523);
nor U3080 (N_3080,N_2271,N_2638);
and U3081 (N_3081,N_2853,N_2737);
and U3082 (N_3082,N_2636,N_2490);
nand U3083 (N_3083,N_2470,N_2600);
and U3084 (N_3084,N_2146,N_2398);
nand U3085 (N_3085,N_2714,N_2004);
nand U3086 (N_3086,N_2534,N_2743);
nand U3087 (N_3087,N_2693,N_2385);
and U3088 (N_3088,N_2184,N_2474);
nand U3089 (N_3089,N_2160,N_2684);
nor U3090 (N_3090,N_2375,N_2834);
xnor U3091 (N_3091,N_2772,N_2255);
and U3092 (N_3092,N_2622,N_2448);
nand U3093 (N_3093,N_2242,N_2456);
nor U3094 (N_3094,N_2558,N_2800);
nor U3095 (N_3095,N_2551,N_2728);
xor U3096 (N_3096,N_2217,N_2342);
xnor U3097 (N_3097,N_2760,N_2664);
nor U3098 (N_3098,N_2933,N_2598);
and U3099 (N_3099,N_2159,N_2086);
or U3100 (N_3100,N_2978,N_2844);
or U3101 (N_3101,N_2124,N_2577);
nand U3102 (N_3102,N_2010,N_2258);
xor U3103 (N_3103,N_2307,N_2024);
or U3104 (N_3104,N_2153,N_2717);
xor U3105 (N_3105,N_2983,N_2589);
xnor U3106 (N_3106,N_2673,N_2295);
nor U3107 (N_3107,N_2550,N_2751);
nor U3108 (N_3108,N_2415,N_2059);
and U3109 (N_3109,N_2789,N_2372);
or U3110 (N_3110,N_2264,N_2000);
xnor U3111 (N_3111,N_2143,N_2311);
nand U3112 (N_3112,N_2626,N_2033);
nor U3113 (N_3113,N_2859,N_2881);
or U3114 (N_3114,N_2670,N_2913);
or U3115 (N_3115,N_2411,N_2027);
nand U3116 (N_3116,N_2949,N_2476);
nor U3117 (N_3117,N_2888,N_2346);
nor U3118 (N_3118,N_2484,N_2871);
xnor U3119 (N_3119,N_2318,N_2548);
nand U3120 (N_3120,N_2125,N_2899);
and U3121 (N_3121,N_2580,N_2574);
or U3122 (N_3122,N_2045,N_2274);
nor U3123 (N_3123,N_2043,N_2756);
or U3124 (N_3124,N_2492,N_2647);
or U3125 (N_3125,N_2379,N_2363);
nand U3126 (N_3126,N_2686,N_2168);
or U3127 (N_3127,N_2777,N_2646);
nand U3128 (N_3128,N_2039,N_2543);
and U3129 (N_3129,N_2254,N_2506);
and U3130 (N_3130,N_2862,N_2323);
nand U3131 (N_3131,N_2354,N_2104);
nand U3132 (N_3132,N_2601,N_2088);
nand U3133 (N_3133,N_2431,N_2042);
or U3134 (N_3134,N_2179,N_2542);
and U3135 (N_3135,N_2056,N_2641);
nor U3136 (N_3136,N_2455,N_2297);
nor U3137 (N_3137,N_2089,N_2754);
and U3138 (N_3138,N_2742,N_2483);
nor U3139 (N_3139,N_2964,N_2569);
xnor U3140 (N_3140,N_2462,N_2430);
xnor U3141 (N_3141,N_2669,N_2613);
and U3142 (N_3142,N_2914,N_2381);
or U3143 (N_3143,N_2989,N_2350);
nor U3144 (N_3144,N_2680,N_2666);
nand U3145 (N_3145,N_2792,N_2321);
nand U3146 (N_3146,N_2420,N_2387);
nand U3147 (N_3147,N_2449,N_2098);
or U3148 (N_3148,N_2215,N_2313);
and U3149 (N_3149,N_2487,N_2606);
nand U3150 (N_3150,N_2085,N_2252);
nand U3151 (N_3151,N_2799,N_2734);
nor U3152 (N_3152,N_2826,N_2828);
or U3153 (N_3153,N_2458,N_2816);
and U3154 (N_3154,N_2849,N_2157);
and U3155 (N_3155,N_2064,N_2833);
nand U3156 (N_3156,N_2514,N_2538);
and U3157 (N_3157,N_2778,N_2355);
nand U3158 (N_3158,N_2338,N_2465);
nor U3159 (N_3159,N_2544,N_2911);
and U3160 (N_3160,N_2695,N_2720);
xor U3161 (N_3161,N_2070,N_2130);
or U3162 (N_3162,N_2460,N_2203);
and U3163 (N_3163,N_2447,N_2031);
or U3164 (N_3164,N_2334,N_2885);
nand U3165 (N_3165,N_2464,N_2727);
nor U3166 (N_3166,N_2109,N_2619);
nor U3167 (N_3167,N_2998,N_2681);
or U3168 (N_3168,N_2876,N_2982);
nor U3169 (N_3169,N_2838,N_2034);
or U3170 (N_3170,N_2189,N_2701);
and U3171 (N_3171,N_2921,N_2142);
nand U3172 (N_3172,N_2546,N_2726);
nor U3173 (N_3173,N_2312,N_2604);
and U3174 (N_3174,N_2685,N_2422);
xnor U3175 (N_3175,N_2200,N_2709);
xor U3176 (N_3176,N_2700,N_2963);
or U3177 (N_3177,N_2540,N_2006);
nand U3178 (N_3178,N_2101,N_2938);
xor U3179 (N_3179,N_2315,N_2827);
xor U3180 (N_3180,N_2239,N_2331);
and U3181 (N_3181,N_2898,N_2253);
nor U3182 (N_3182,N_2951,N_2212);
nor U3183 (N_3183,N_2620,N_2018);
nand U3184 (N_3184,N_2658,N_2723);
and U3185 (N_3185,N_2081,N_2892);
and U3186 (N_3186,N_2352,N_2023);
nor U3187 (N_3187,N_2316,N_2865);
nand U3188 (N_3188,N_2198,N_2794);
nor U3189 (N_3189,N_2190,N_2221);
and U3190 (N_3190,N_2453,N_2301);
or U3191 (N_3191,N_2592,N_2251);
nand U3192 (N_3192,N_2151,N_2061);
or U3193 (N_3193,N_2582,N_2591);
nor U3194 (N_3194,N_2065,N_2126);
nand U3195 (N_3195,N_2093,N_2729);
xnor U3196 (N_3196,N_2858,N_2290);
and U3197 (N_3197,N_2722,N_2161);
or U3198 (N_3198,N_2611,N_2234);
nor U3199 (N_3199,N_2840,N_2225);
and U3200 (N_3200,N_2218,N_2861);
and U3201 (N_3201,N_2993,N_2781);
xnor U3202 (N_3202,N_2749,N_2481);
or U3203 (N_3203,N_2328,N_2150);
nand U3204 (N_3204,N_2062,N_2891);
and U3205 (N_3205,N_2541,N_2284);
nor U3206 (N_3206,N_2555,N_2076);
nor U3207 (N_3207,N_2300,N_2030);
nand U3208 (N_3208,N_2240,N_2191);
and U3209 (N_3209,N_2782,N_2376);
nor U3210 (N_3210,N_2444,N_2185);
nor U3211 (N_3211,N_2025,N_2015);
xnor U3212 (N_3212,N_2280,N_2026);
nor U3213 (N_3213,N_2716,N_2846);
nor U3214 (N_3214,N_2689,N_2928);
nor U3215 (N_3215,N_2395,N_2073);
and U3216 (N_3216,N_2007,N_2932);
nand U3217 (N_3217,N_2261,N_2281);
or U3218 (N_3218,N_2752,N_2451);
or U3219 (N_3219,N_2132,N_2223);
nor U3220 (N_3220,N_2116,N_2486);
nand U3221 (N_3221,N_2173,N_2304);
nor U3222 (N_3222,N_2575,N_2854);
or U3223 (N_3223,N_2986,N_2428);
or U3224 (N_3224,N_2802,N_2192);
nor U3225 (N_3225,N_2702,N_2903);
nor U3226 (N_3226,N_2570,N_2652);
or U3227 (N_3227,N_2783,N_2848);
and U3228 (N_3228,N_2054,N_2617);
nor U3229 (N_3229,N_2805,N_2270);
or U3230 (N_3230,N_2437,N_2894);
or U3231 (N_3231,N_2516,N_2764);
nand U3232 (N_3232,N_2919,N_2485);
nor U3233 (N_3233,N_2419,N_2618);
and U3234 (N_3234,N_2524,N_2051);
nand U3235 (N_3235,N_2337,N_2711);
or U3236 (N_3236,N_2275,N_2835);
nor U3237 (N_3237,N_2990,N_2353);
nor U3238 (N_3238,N_2879,N_2236);
and U3239 (N_3239,N_2364,N_2930);
nor U3240 (N_3240,N_2256,N_2528);
and U3241 (N_3241,N_2175,N_2654);
nand U3242 (N_3242,N_2904,N_2961);
nor U3243 (N_3243,N_2603,N_2494);
xnor U3244 (N_3244,N_2768,N_2980);
and U3245 (N_3245,N_2103,N_2498);
or U3246 (N_3246,N_2659,N_2852);
or U3247 (N_3247,N_2806,N_2515);
and U3248 (N_3248,N_2421,N_2801);
or U3249 (N_3249,N_2079,N_2187);
nand U3250 (N_3250,N_2905,N_2656);
nand U3251 (N_3251,N_2400,N_2948);
nand U3252 (N_3252,N_2757,N_2774);
or U3253 (N_3253,N_2955,N_2706);
or U3254 (N_3254,N_2384,N_2022);
and U3255 (N_3255,N_2021,N_2553);
nand U3256 (N_3256,N_2697,N_2211);
xor U3257 (N_3257,N_2900,N_2227);
or U3258 (N_3258,N_2305,N_2572);
or U3259 (N_3259,N_2029,N_2438);
nor U3260 (N_3260,N_2196,N_2228);
or U3261 (N_3261,N_2171,N_2306);
and U3262 (N_3262,N_2565,N_2935);
or U3263 (N_3263,N_2303,N_2108);
xnor U3264 (N_3264,N_2741,N_2841);
or U3265 (N_3265,N_2902,N_2053);
nand U3266 (N_3266,N_2365,N_2374);
or U3267 (N_3267,N_2339,N_2099);
nor U3268 (N_3268,N_2302,N_2707);
and U3269 (N_3269,N_2267,N_2653);
and U3270 (N_3270,N_2908,N_2566);
nor U3271 (N_3271,N_2889,N_2226);
and U3272 (N_3272,N_2299,N_2556);
or U3273 (N_3273,N_2944,N_2260);
or U3274 (N_3274,N_2245,N_2248);
or U3275 (N_3275,N_2473,N_2895);
xnor U3276 (N_3276,N_2105,N_2378);
and U3277 (N_3277,N_2775,N_2207);
nor U3278 (N_3278,N_2612,N_2581);
or U3279 (N_3279,N_2087,N_2050);
nor U3280 (N_3280,N_2960,N_2956);
nor U3281 (N_3281,N_2137,N_2682);
nand U3282 (N_3282,N_2610,N_2154);
nor U3283 (N_3283,N_2668,N_2075);
nand U3284 (N_3284,N_2724,N_2368);
nor U3285 (N_3285,N_2925,N_2324);
or U3286 (N_3286,N_2044,N_2644);
and U3287 (N_3287,N_2107,N_2136);
nand U3288 (N_3288,N_2786,N_2020);
or U3289 (N_3289,N_2504,N_2084);
nand U3290 (N_3290,N_2113,N_2148);
xor U3291 (N_3291,N_2230,N_2232);
and U3292 (N_3292,N_2812,N_2585);
nand U3293 (N_3293,N_2621,N_2063);
or U3294 (N_3294,N_2595,N_2441);
xor U3295 (N_3295,N_2520,N_2501);
xnor U3296 (N_3296,N_2851,N_2283);
nand U3297 (N_3297,N_2106,N_2243);
nand U3298 (N_3298,N_2279,N_2518);
or U3299 (N_3299,N_2738,N_2587);
nor U3300 (N_3300,N_2344,N_2092);
or U3301 (N_3301,N_2563,N_2069);
nor U3302 (N_3302,N_2508,N_2014);
or U3303 (N_3303,N_2127,N_2102);
nand U3304 (N_3304,N_2055,N_2819);
and U3305 (N_3305,N_2210,N_2629);
nor U3306 (N_3306,N_2537,N_2522);
nor U3307 (N_3307,N_2072,N_2567);
nand U3308 (N_3308,N_2809,N_2869);
nand U3309 (N_3309,N_2912,N_2785);
and U3310 (N_3310,N_2576,N_2402);
xnor U3311 (N_3311,N_2166,N_2817);
or U3312 (N_3312,N_2407,N_2906);
nor U3313 (N_3313,N_2571,N_2526);
or U3314 (N_3314,N_2747,N_2814);
nand U3315 (N_3315,N_2939,N_2035);
nor U3316 (N_3316,N_2118,N_2286);
or U3317 (N_3317,N_2650,N_2630);
and U3318 (N_3318,N_2634,N_2268);
or U3319 (N_3319,N_2699,N_2798);
nor U3320 (N_3320,N_2206,N_2796);
nor U3321 (N_3321,N_2360,N_2836);
xor U3322 (N_3322,N_2767,N_2773);
xor U3323 (N_3323,N_2097,N_2144);
nand U3324 (N_3324,N_2878,N_2257);
nor U3325 (N_3325,N_2645,N_2822);
nand U3326 (N_3326,N_2310,N_2133);
nand U3327 (N_3327,N_2942,N_2959);
or U3328 (N_3328,N_2434,N_2358);
nand U3329 (N_3329,N_2954,N_2366);
nor U3330 (N_3330,N_2941,N_2825);
nor U3331 (N_3331,N_2766,N_2679);
nor U3332 (N_3332,N_2122,N_2382);
nor U3333 (N_3333,N_2839,N_2525);
or U3334 (N_3334,N_2934,N_2111);
and U3335 (N_3335,N_2262,N_2665);
nand U3336 (N_3336,N_2813,N_2549);
or U3337 (N_3337,N_2343,N_2884);
and U3338 (N_3338,N_2273,N_2803);
nor U3339 (N_3339,N_2040,N_2399);
and U3340 (N_3340,N_2265,N_2195);
nand U3341 (N_3341,N_2996,N_2468);
nand U3342 (N_3342,N_2291,N_2009);
nor U3343 (N_3343,N_2733,N_2683);
nor U3344 (N_3344,N_2627,N_2924);
and U3345 (N_3345,N_2459,N_2074);
nand U3346 (N_3346,N_2067,N_2373);
and U3347 (N_3347,N_2367,N_2687);
xnor U3348 (N_3348,N_2753,N_2219);
or U3349 (N_3349,N_2655,N_2403);
nand U3350 (N_3350,N_2625,N_2052);
and U3351 (N_3351,N_2887,N_2497);
nor U3352 (N_3352,N_2847,N_2639);
xor U3353 (N_3353,N_2517,N_2298);
nor U3354 (N_3354,N_2811,N_2152);
xnor U3355 (N_3355,N_2155,N_2984);
nor U3356 (N_3356,N_2095,N_2605);
and U3357 (N_3357,N_2289,N_2488);
or U3358 (N_3358,N_2454,N_2377);
and U3359 (N_3359,N_2489,N_2002);
nor U3360 (N_3360,N_2821,N_2436);
or U3361 (N_3361,N_2393,N_2479);
and U3362 (N_3362,N_2369,N_2467);
nor U3363 (N_3363,N_2864,N_2943);
xor U3364 (N_3364,N_2882,N_2509);
nand U3365 (N_3365,N_2744,N_2971);
nor U3366 (N_3366,N_2466,N_2918);
xor U3367 (N_3367,N_2246,N_2732);
nor U3368 (N_3368,N_2469,N_2164);
nand U3369 (N_3369,N_2780,N_2616);
nor U3370 (N_3370,N_2208,N_2926);
nor U3371 (N_3371,N_2336,N_2440);
nor U3372 (N_3372,N_2077,N_2976);
and U3373 (N_3373,N_2667,N_2532);
and U3374 (N_3374,N_2609,N_2559);
nand U3375 (N_3375,N_2703,N_2791);
nand U3376 (N_3376,N_2718,N_2972);
or U3377 (N_3377,N_2830,N_2815);
nand U3378 (N_3378,N_2201,N_2607);
nor U3379 (N_3379,N_2860,N_2406);
nand U3380 (N_3380,N_2266,N_2129);
and U3381 (N_3381,N_2293,N_2414);
nor U3382 (N_3382,N_2439,N_2475);
and U3383 (N_3383,N_2263,N_2586);
or U3384 (N_3384,N_2761,N_2288);
xor U3385 (N_3385,N_2362,N_2214);
and U3386 (N_3386,N_2967,N_2573);
and U3387 (N_3387,N_2357,N_2698);
nor U3388 (N_3388,N_2410,N_2735);
and U3389 (N_3389,N_2535,N_2608);
nor U3390 (N_3390,N_2188,N_2715);
and U3391 (N_3391,N_2011,N_2068);
nor U3392 (N_3392,N_2292,N_2886);
nor U3393 (N_3393,N_2416,N_2250);
and U3394 (N_3394,N_2843,N_2725);
or U3395 (N_3395,N_2433,N_2047);
nand U3396 (N_3396,N_2100,N_2401);
or U3397 (N_3397,N_2995,N_2046);
nand U3398 (N_3398,N_2167,N_2519);
nor U3399 (N_3399,N_2945,N_2457);
nand U3400 (N_3400,N_2371,N_2810);
and U3401 (N_3401,N_2308,N_2624);
or U3402 (N_3402,N_2162,N_2920);
nor U3403 (N_3403,N_2193,N_2863);
nand U3404 (N_3404,N_2176,N_2450);
nor U3405 (N_3405,N_2588,N_2424);
nand U3406 (N_3406,N_2028,N_2423);
and U3407 (N_3407,N_2552,N_2080);
and U3408 (N_3408,N_2445,N_2163);
nor U3409 (N_3409,N_2874,N_2119);
nor U3410 (N_3410,N_2507,N_2907);
and U3411 (N_3411,N_2333,N_2615);
nand U3412 (N_3412,N_2994,N_2829);
nand U3413 (N_3413,N_2536,N_2016);
or U3414 (N_3414,N_2677,N_2241);
or U3415 (N_3415,N_2285,N_2472);
xor U3416 (N_3416,N_2736,N_2158);
or U3417 (N_3417,N_2807,N_2568);
or U3418 (N_3418,N_2818,N_2628);
nor U3419 (N_3419,N_2643,N_2272);
xnor U3420 (N_3420,N_2205,N_2209);
nor U3421 (N_3421,N_2202,N_2478);
xnor U3422 (N_3422,N_2032,N_2177);
nand U3423 (N_3423,N_2165,N_2141);
nand U3424 (N_3424,N_2952,N_2231);
nor U3425 (N_3425,N_2651,N_2795);
nand U3426 (N_3426,N_2322,N_2790);
nand U3427 (N_3427,N_2676,N_2713);
or U3428 (N_3428,N_2564,N_2883);
and U3429 (N_3429,N_2480,N_2877);
nor U3430 (N_3430,N_2875,N_2896);
nor U3431 (N_3431,N_2590,N_2987);
xnor U3432 (N_3432,N_2249,N_2429);
nor U3433 (N_3433,N_2495,N_2446);
and U3434 (N_3434,N_2710,N_2880);
or U3435 (N_3435,N_2533,N_2529);
and U3436 (N_3436,N_2599,N_2970);
or U3437 (N_3437,N_2910,N_2746);
or U3438 (N_3438,N_2276,N_2797);
nor U3439 (N_3439,N_2614,N_2341);
and U3440 (N_3440,N_2969,N_2389);
nor U3441 (N_3441,N_2631,N_2704);
or U3442 (N_3442,N_2985,N_2408);
or U3443 (N_3443,N_2287,N_2513);
and U3444 (N_3444,N_2197,N_2690);
and U3445 (N_3445,N_2319,N_2962);
nand U3446 (N_3446,N_2309,N_2120);
and U3447 (N_3447,N_2008,N_2916);
and U3448 (N_3448,N_2499,N_2096);
and U3449 (N_3449,N_2692,N_2066);
or U3450 (N_3450,N_2992,N_2850);
nand U3451 (N_3451,N_2719,N_2500);
nand U3452 (N_3452,N_2936,N_2623);
nand U3453 (N_3453,N_2503,N_2277);
nand U3454 (N_3454,N_2397,N_2169);
nand U3455 (N_3455,N_2121,N_2527);
nor U3456 (N_3456,N_2758,N_2539);
nor U3457 (N_3457,N_2696,N_2237);
nor U3458 (N_3458,N_2660,N_2866);
nor U3459 (N_3459,N_2842,N_2705);
and U3460 (N_3460,N_2657,N_2390);
nand U3461 (N_3461,N_2335,N_2545);
or U3462 (N_3462,N_2426,N_2635);
nand U3463 (N_3463,N_2632,N_2831);
nand U3464 (N_3464,N_2561,N_2493);
xor U3465 (N_3465,N_2019,N_2090);
nand U3466 (N_3466,N_2562,N_2314);
or U3467 (N_3467,N_2356,N_2968);
nor U3468 (N_3468,N_2991,N_2463);
nand U3469 (N_3469,N_2178,N_2804);
nand U3470 (N_3470,N_2404,N_2759);
and U3471 (N_3471,N_2412,N_2915);
or U3472 (N_3472,N_2678,N_2779);
nand U3473 (N_3473,N_2182,N_2138);
nor U3474 (N_3474,N_2511,N_2296);
and U3475 (N_3475,N_2329,N_2180);
nor U3476 (N_3476,N_2134,N_2269);
nand U3477 (N_3477,N_2649,N_2909);
nor U3478 (N_3478,N_2233,N_2135);
nor U3479 (N_3479,N_2845,N_2222);
and U3480 (N_3480,N_2392,N_2435);
or U3481 (N_3481,N_2083,N_2386);
and U3482 (N_3482,N_2521,N_2642);
xnor U3483 (N_3483,N_2748,N_2432);
nor U3484 (N_3484,N_2259,N_2115);
nor U3485 (N_3485,N_2663,N_2320);
or U3486 (N_3486,N_2345,N_2893);
or U3487 (N_3487,N_2396,N_2170);
nand U3488 (N_3488,N_2147,N_2793);
xor U3489 (N_3489,N_2730,N_2091);
or U3490 (N_3490,N_2763,N_2897);
and U3491 (N_3491,N_2671,N_2477);
and U3492 (N_3492,N_2359,N_2966);
xor U3493 (N_3493,N_2593,N_2388);
nand U3494 (N_3494,N_2740,N_2349);
nor U3495 (N_3495,N_2868,N_2890);
nor U3496 (N_3496,N_2071,N_2554);
nor U3497 (N_3497,N_2808,N_2855);
and U3498 (N_3498,N_2674,N_2596);
nor U3499 (N_3499,N_2691,N_2637);
nand U3500 (N_3500,N_2469,N_2560);
nor U3501 (N_3501,N_2665,N_2949);
nand U3502 (N_3502,N_2441,N_2835);
or U3503 (N_3503,N_2033,N_2193);
nand U3504 (N_3504,N_2890,N_2598);
nor U3505 (N_3505,N_2552,N_2532);
or U3506 (N_3506,N_2452,N_2910);
nor U3507 (N_3507,N_2341,N_2404);
nor U3508 (N_3508,N_2795,N_2773);
nor U3509 (N_3509,N_2370,N_2601);
and U3510 (N_3510,N_2613,N_2630);
nand U3511 (N_3511,N_2237,N_2965);
or U3512 (N_3512,N_2012,N_2248);
or U3513 (N_3513,N_2852,N_2609);
or U3514 (N_3514,N_2223,N_2117);
nor U3515 (N_3515,N_2218,N_2867);
or U3516 (N_3516,N_2098,N_2023);
or U3517 (N_3517,N_2037,N_2743);
or U3518 (N_3518,N_2333,N_2404);
and U3519 (N_3519,N_2993,N_2076);
nand U3520 (N_3520,N_2845,N_2483);
or U3521 (N_3521,N_2123,N_2400);
nand U3522 (N_3522,N_2781,N_2310);
and U3523 (N_3523,N_2151,N_2146);
or U3524 (N_3524,N_2660,N_2210);
or U3525 (N_3525,N_2045,N_2450);
xor U3526 (N_3526,N_2569,N_2105);
and U3527 (N_3527,N_2353,N_2696);
or U3528 (N_3528,N_2394,N_2711);
nand U3529 (N_3529,N_2933,N_2376);
and U3530 (N_3530,N_2074,N_2702);
nor U3531 (N_3531,N_2321,N_2574);
and U3532 (N_3532,N_2406,N_2016);
and U3533 (N_3533,N_2815,N_2855);
nor U3534 (N_3534,N_2123,N_2207);
or U3535 (N_3535,N_2521,N_2144);
and U3536 (N_3536,N_2643,N_2567);
nor U3537 (N_3537,N_2258,N_2728);
nand U3538 (N_3538,N_2747,N_2627);
and U3539 (N_3539,N_2433,N_2096);
nor U3540 (N_3540,N_2979,N_2416);
nand U3541 (N_3541,N_2561,N_2573);
nand U3542 (N_3542,N_2639,N_2351);
nand U3543 (N_3543,N_2337,N_2287);
and U3544 (N_3544,N_2922,N_2490);
or U3545 (N_3545,N_2648,N_2606);
and U3546 (N_3546,N_2947,N_2602);
xor U3547 (N_3547,N_2662,N_2896);
or U3548 (N_3548,N_2352,N_2048);
or U3549 (N_3549,N_2936,N_2637);
xnor U3550 (N_3550,N_2666,N_2836);
nand U3551 (N_3551,N_2125,N_2309);
xnor U3552 (N_3552,N_2805,N_2458);
nand U3553 (N_3553,N_2241,N_2313);
nand U3554 (N_3554,N_2281,N_2886);
or U3555 (N_3555,N_2290,N_2162);
nand U3556 (N_3556,N_2587,N_2494);
nor U3557 (N_3557,N_2431,N_2605);
or U3558 (N_3558,N_2567,N_2395);
or U3559 (N_3559,N_2329,N_2602);
and U3560 (N_3560,N_2680,N_2973);
nand U3561 (N_3561,N_2592,N_2725);
or U3562 (N_3562,N_2172,N_2122);
or U3563 (N_3563,N_2684,N_2475);
xor U3564 (N_3564,N_2296,N_2886);
and U3565 (N_3565,N_2201,N_2104);
nand U3566 (N_3566,N_2214,N_2271);
nor U3567 (N_3567,N_2898,N_2776);
nor U3568 (N_3568,N_2284,N_2042);
nand U3569 (N_3569,N_2557,N_2864);
and U3570 (N_3570,N_2380,N_2860);
or U3571 (N_3571,N_2724,N_2548);
and U3572 (N_3572,N_2615,N_2706);
or U3573 (N_3573,N_2661,N_2721);
nand U3574 (N_3574,N_2897,N_2011);
xor U3575 (N_3575,N_2826,N_2692);
or U3576 (N_3576,N_2653,N_2703);
xor U3577 (N_3577,N_2647,N_2298);
nand U3578 (N_3578,N_2369,N_2421);
and U3579 (N_3579,N_2417,N_2386);
nand U3580 (N_3580,N_2118,N_2452);
and U3581 (N_3581,N_2393,N_2060);
and U3582 (N_3582,N_2860,N_2994);
nand U3583 (N_3583,N_2103,N_2061);
nand U3584 (N_3584,N_2989,N_2897);
and U3585 (N_3585,N_2504,N_2658);
or U3586 (N_3586,N_2529,N_2971);
xnor U3587 (N_3587,N_2624,N_2546);
or U3588 (N_3588,N_2472,N_2611);
nor U3589 (N_3589,N_2950,N_2192);
nand U3590 (N_3590,N_2744,N_2511);
and U3591 (N_3591,N_2167,N_2685);
and U3592 (N_3592,N_2717,N_2663);
nor U3593 (N_3593,N_2407,N_2539);
nand U3594 (N_3594,N_2426,N_2422);
nand U3595 (N_3595,N_2641,N_2911);
and U3596 (N_3596,N_2298,N_2120);
nand U3597 (N_3597,N_2912,N_2763);
xnor U3598 (N_3598,N_2324,N_2124);
nor U3599 (N_3599,N_2027,N_2029);
and U3600 (N_3600,N_2046,N_2984);
nor U3601 (N_3601,N_2084,N_2147);
xor U3602 (N_3602,N_2915,N_2358);
nand U3603 (N_3603,N_2257,N_2800);
nor U3604 (N_3604,N_2932,N_2322);
nor U3605 (N_3605,N_2251,N_2431);
or U3606 (N_3606,N_2980,N_2535);
or U3607 (N_3607,N_2268,N_2909);
nor U3608 (N_3608,N_2200,N_2416);
nor U3609 (N_3609,N_2177,N_2344);
or U3610 (N_3610,N_2054,N_2452);
nand U3611 (N_3611,N_2546,N_2972);
nor U3612 (N_3612,N_2690,N_2794);
and U3613 (N_3613,N_2936,N_2396);
and U3614 (N_3614,N_2654,N_2955);
or U3615 (N_3615,N_2899,N_2690);
and U3616 (N_3616,N_2010,N_2198);
and U3617 (N_3617,N_2858,N_2955);
or U3618 (N_3618,N_2450,N_2884);
nand U3619 (N_3619,N_2198,N_2775);
and U3620 (N_3620,N_2832,N_2431);
or U3621 (N_3621,N_2747,N_2352);
nor U3622 (N_3622,N_2711,N_2201);
nor U3623 (N_3623,N_2840,N_2346);
or U3624 (N_3624,N_2195,N_2080);
and U3625 (N_3625,N_2745,N_2919);
and U3626 (N_3626,N_2964,N_2798);
or U3627 (N_3627,N_2014,N_2020);
nand U3628 (N_3628,N_2097,N_2447);
or U3629 (N_3629,N_2584,N_2313);
nor U3630 (N_3630,N_2514,N_2361);
nor U3631 (N_3631,N_2180,N_2101);
or U3632 (N_3632,N_2085,N_2997);
nand U3633 (N_3633,N_2202,N_2630);
or U3634 (N_3634,N_2569,N_2502);
nand U3635 (N_3635,N_2380,N_2699);
or U3636 (N_3636,N_2909,N_2083);
or U3637 (N_3637,N_2071,N_2839);
nor U3638 (N_3638,N_2404,N_2942);
nand U3639 (N_3639,N_2221,N_2731);
and U3640 (N_3640,N_2766,N_2513);
nor U3641 (N_3641,N_2847,N_2904);
and U3642 (N_3642,N_2545,N_2598);
or U3643 (N_3643,N_2554,N_2250);
nor U3644 (N_3644,N_2673,N_2920);
and U3645 (N_3645,N_2176,N_2926);
and U3646 (N_3646,N_2911,N_2978);
or U3647 (N_3647,N_2657,N_2873);
nor U3648 (N_3648,N_2873,N_2808);
or U3649 (N_3649,N_2684,N_2677);
and U3650 (N_3650,N_2122,N_2857);
and U3651 (N_3651,N_2747,N_2355);
and U3652 (N_3652,N_2461,N_2789);
or U3653 (N_3653,N_2583,N_2428);
or U3654 (N_3654,N_2227,N_2054);
and U3655 (N_3655,N_2381,N_2829);
xor U3656 (N_3656,N_2062,N_2189);
nand U3657 (N_3657,N_2528,N_2255);
and U3658 (N_3658,N_2267,N_2409);
nor U3659 (N_3659,N_2055,N_2605);
nand U3660 (N_3660,N_2034,N_2954);
or U3661 (N_3661,N_2294,N_2767);
nor U3662 (N_3662,N_2999,N_2280);
nand U3663 (N_3663,N_2170,N_2244);
or U3664 (N_3664,N_2592,N_2938);
or U3665 (N_3665,N_2280,N_2054);
nor U3666 (N_3666,N_2868,N_2139);
nand U3667 (N_3667,N_2257,N_2162);
xnor U3668 (N_3668,N_2902,N_2010);
nand U3669 (N_3669,N_2182,N_2140);
and U3670 (N_3670,N_2540,N_2085);
nand U3671 (N_3671,N_2609,N_2822);
nand U3672 (N_3672,N_2932,N_2714);
xor U3673 (N_3673,N_2333,N_2910);
and U3674 (N_3674,N_2293,N_2052);
nand U3675 (N_3675,N_2199,N_2802);
nor U3676 (N_3676,N_2626,N_2464);
and U3677 (N_3677,N_2186,N_2731);
nand U3678 (N_3678,N_2555,N_2106);
nand U3679 (N_3679,N_2045,N_2096);
and U3680 (N_3680,N_2029,N_2063);
nor U3681 (N_3681,N_2758,N_2382);
nor U3682 (N_3682,N_2200,N_2570);
nor U3683 (N_3683,N_2503,N_2773);
nand U3684 (N_3684,N_2202,N_2031);
nand U3685 (N_3685,N_2377,N_2392);
nor U3686 (N_3686,N_2816,N_2012);
or U3687 (N_3687,N_2757,N_2857);
and U3688 (N_3688,N_2221,N_2109);
nor U3689 (N_3689,N_2741,N_2159);
nand U3690 (N_3690,N_2923,N_2560);
and U3691 (N_3691,N_2289,N_2855);
or U3692 (N_3692,N_2036,N_2357);
nor U3693 (N_3693,N_2605,N_2991);
or U3694 (N_3694,N_2527,N_2240);
and U3695 (N_3695,N_2126,N_2290);
xor U3696 (N_3696,N_2604,N_2224);
and U3697 (N_3697,N_2644,N_2508);
or U3698 (N_3698,N_2896,N_2643);
and U3699 (N_3699,N_2327,N_2711);
or U3700 (N_3700,N_2308,N_2595);
nor U3701 (N_3701,N_2756,N_2130);
or U3702 (N_3702,N_2300,N_2077);
nor U3703 (N_3703,N_2326,N_2588);
and U3704 (N_3704,N_2084,N_2202);
nor U3705 (N_3705,N_2486,N_2950);
nand U3706 (N_3706,N_2288,N_2646);
nand U3707 (N_3707,N_2342,N_2516);
nand U3708 (N_3708,N_2692,N_2551);
or U3709 (N_3709,N_2315,N_2938);
or U3710 (N_3710,N_2247,N_2882);
xor U3711 (N_3711,N_2482,N_2879);
or U3712 (N_3712,N_2410,N_2274);
and U3713 (N_3713,N_2825,N_2671);
nand U3714 (N_3714,N_2944,N_2185);
nor U3715 (N_3715,N_2213,N_2595);
and U3716 (N_3716,N_2038,N_2818);
nor U3717 (N_3717,N_2869,N_2034);
nor U3718 (N_3718,N_2683,N_2121);
and U3719 (N_3719,N_2441,N_2807);
nor U3720 (N_3720,N_2082,N_2247);
or U3721 (N_3721,N_2470,N_2468);
nand U3722 (N_3722,N_2243,N_2914);
nor U3723 (N_3723,N_2913,N_2152);
and U3724 (N_3724,N_2757,N_2883);
and U3725 (N_3725,N_2235,N_2036);
nor U3726 (N_3726,N_2830,N_2588);
nand U3727 (N_3727,N_2779,N_2351);
nand U3728 (N_3728,N_2401,N_2355);
or U3729 (N_3729,N_2636,N_2065);
and U3730 (N_3730,N_2227,N_2471);
and U3731 (N_3731,N_2230,N_2011);
or U3732 (N_3732,N_2722,N_2468);
or U3733 (N_3733,N_2199,N_2720);
nand U3734 (N_3734,N_2092,N_2632);
nand U3735 (N_3735,N_2967,N_2036);
and U3736 (N_3736,N_2913,N_2396);
or U3737 (N_3737,N_2960,N_2723);
nor U3738 (N_3738,N_2518,N_2593);
nand U3739 (N_3739,N_2535,N_2614);
or U3740 (N_3740,N_2912,N_2128);
nor U3741 (N_3741,N_2285,N_2319);
nand U3742 (N_3742,N_2448,N_2803);
nand U3743 (N_3743,N_2036,N_2936);
xor U3744 (N_3744,N_2908,N_2565);
nor U3745 (N_3745,N_2474,N_2097);
nor U3746 (N_3746,N_2615,N_2420);
nor U3747 (N_3747,N_2200,N_2378);
or U3748 (N_3748,N_2049,N_2668);
nand U3749 (N_3749,N_2843,N_2437);
nand U3750 (N_3750,N_2111,N_2358);
xor U3751 (N_3751,N_2056,N_2943);
nor U3752 (N_3752,N_2056,N_2109);
or U3753 (N_3753,N_2801,N_2215);
nand U3754 (N_3754,N_2776,N_2057);
nor U3755 (N_3755,N_2783,N_2339);
or U3756 (N_3756,N_2241,N_2983);
xor U3757 (N_3757,N_2335,N_2375);
nand U3758 (N_3758,N_2407,N_2437);
or U3759 (N_3759,N_2304,N_2746);
and U3760 (N_3760,N_2233,N_2522);
or U3761 (N_3761,N_2318,N_2191);
or U3762 (N_3762,N_2458,N_2032);
nand U3763 (N_3763,N_2200,N_2591);
xnor U3764 (N_3764,N_2015,N_2215);
nand U3765 (N_3765,N_2924,N_2665);
xor U3766 (N_3766,N_2225,N_2596);
nand U3767 (N_3767,N_2834,N_2342);
or U3768 (N_3768,N_2385,N_2530);
nor U3769 (N_3769,N_2325,N_2090);
nor U3770 (N_3770,N_2741,N_2965);
xor U3771 (N_3771,N_2880,N_2671);
and U3772 (N_3772,N_2054,N_2982);
nor U3773 (N_3773,N_2780,N_2299);
nor U3774 (N_3774,N_2390,N_2643);
xnor U3775 (N_3775,N_2686,N_2755);
and U3776 (N_3776,N_2878,N_2218);
or U3777 (N_3777,N_2772,N_2903);
or U3778 (N_3778,N_2081,N_2692);
nor U3779 (N_3779,N_2732,N_2359);
nor U3780 (N_3780,N_2504,N_2923);
or U3781 (N_3781,N_2617,N_2486);
and U3782 (N_3782,N_2153,N_2421);
nand U3783 (N_3783,N_2536,N_2738);
and U3784 (N_3784,N_2256,N_2544);
nand U3785 (N_3785,N_2972,N_2176);
nand U3786 (N_3786,N_2107,N_2963);
or U3787 (N_3787,N_2674,N_2169);
nor U3788 (N_3788,N_2169,N_2747);
nand U3789 (N_3789,N_2094,N_2509);
nor U3790 (N_3790,N_2308,N_2583);
or U3791 (N_3791,N_2436,N_2162);
nor U3792 (N_3792,N_2062,N_2043);
or U3793 (N_3793,N_2591,N_2277);
nand U3794 (N_3794,N_2125,N_2319);
nor U3795 (N_3795,N_2229,N_2646);
or U3796 (N_3796,N_2831,N_2408);
nand U3797 (N_3797,N_2251,N_2034);
nand U3798 (N_3798,N_2224,N_2529);
or U3799 (N_3799,N_2229,N_2268);
nor U3800 (N_3800,N_2586,N_2566);
or U3801 (N_3801,N_2705,N_2167);
nand U3802 (N_3802,N_2185,N_2363);
or U3803 (N_3803,N_2922,N_2815);
and U3804 (N_3804,N_2196,N_2359);
or U3805 (N_3805,N_2313,N_2213);
nand U3806 (N_3806,N_2493,N_2454);
nor U3807 (N_3807,N_2446,N_2436);
nor U3808 (N_3808,N_2830,N_2765);
nand U3809 (N_3809,N_2876,N_2564);
or U3810 (N_3810,N_2437,N_2454);
and U3811 (N_3811,N_2537,N_2493);
and U3812 (N_3812,N_2450,N_2249);
nand U3813 (N_3813,N_2697,N_2206);
nand U3814 (N_3814,N_2988,N_2781);
xnor U3815 (N_3815,N_2066,N_2925);
nand U3816 (N_3816,N_2016,N_2979);
or U3817 (N_3817,N_2202,N_2845);
nor U3818 (N_3818,N_2659,N_2225);
xor U3819 (N_3819,N_2646,N_2243);
or U3820 (N_3820,N_2198,N_2924);
nand U3821 (N_3821,N_2465,N_2213);
and U3822 (N_3822,N_2028,N_2725);
nand U3823 (N_3823,N_2831,N_2258);
nand U3824 (N_3824,N_2232,N_2114);
nor U3825 (N_3825,N_2549,N_2548);
xnor U3826 (N_3826,N_2366,N_2242);
nor U3827 (N_3827,N_2652,N_2011);
or U3828 (N_3828,N_2667,N_2958);
nor U3829 (N_3829,N_2786,N_2881);
nand U3830 (N_3830,N_2242,N_2061);
or U3831 (N_3831,N_2933,N_2758);
nand U3832 (N_3832,N_2722,N_2671);
and U3833 (N_3833,N_2216,N_2580);
nand U3834 (N_3834,N_2592,N_2531);
nor U3835 (N_3835,N_2975,N_2221);
nor U3836 (N_3836,N_2386,N_2524);
nor U3837 (N_3837,N_2519,N_2715);
nor U3838 (N_3838,N_2044,N_2295);
and U3839 (N_3839,N_2208,N_2897);
or U3840 (N_3840,N_2890,N_2243);
xor U3841 (N_3841,N_2338,N_2419);
nor U3842 (N_3842,N_2464,N_2670);
and U3843 (N_3843,N_2588,N_2541);
or U3844 (N_3844,N_2483,N_2811);
nand U3845 (N_3845,N_2397,N_2985);
nor U3846 (N_3846,N_2603,N_2012);
nor U3847 (N_3847,N_2397,N_2762);
or U3848 (N_3848,N_2419,N_2913);
or U3849 (N_3849,N_2627,N_2356);
nand U3850 (N_3850,N_2254,N_2289);
and U3851 (N_3851,N_2951,N_2192);
nor U3852 (N_3852,N_2038,N_2242);
nor U3853 (N_3853,N_2883,N_2586);
or U3854 (N_3854,N_2223,N_2522);
nand U3855 (N_3855,N_2136,N_2204);
and U3856 (N_3856,N_2025,N_2947);
nand U3857 (N_3857,N_2943,N_2607);
and U3858 (N_3858,N_2788,N_2053);
and U3859 (N_3859,N_2696,N_2008);
nor U3860 (N_3860,N_2354,N_2676);
nand U3861 (N_3861,N_2246,N_2623);
or U3862 (N_3862,N_2250,N_2379);
xor U3863 (N_3863,N_2701,N_2098);
nor U3864 (N_3864,N_2189,N_2531);
nand U3865 (N_3865,N_2350,N_2414);
nor U3866 (N_3866,N_2204,N_2148);
and U3867 (N_3867,N_2959,N_2045);
xnor U3868 (N_3868,N_2780,N_2789);
nor U3869 (N_3869,N_2438,N_2394);
xor U3870 (N_3870,N_2312,N_2979);
nand U3871 (N_3871,N_2986,N_2591);
nor U3872 (N_3872,N_2880,N_2101);
or U3873 (N_3873,N_2390,N_2820);
nand U3874 (N_3874,N_2033,N_2717);
or U3875 (N_3875,N_2693,N_2387);
and U3876 (N_3876,N_2483,N_2008);
or U3877 (N_3877,N_2239,N_2295);
nor U3878 (N_3878,N_2312,N_2096);
xnor U3879 (N_3879,N_2309,N_2071);
nor U3880 (N_3880,N_2373,N_2782);
nor U3881 (N_3881,N_2691,N_2489);
nand U3882 (N_3882,N_2544,N_2342);
and U3883 (N_3883,N_2893,N_2021);
and U3884 (N_3884,N_2726,N_2972);
and U3885 (N_3885,N_2302,N_2478);
or U3886 (N_3886,N_2043,N_2620);
or U3887 (N_3887,N_2770,N_2077);
or U3888 (N_3888,N_2196,N_2739);
xnor U3889 (N_3889,N_2647,N_2920);
xnor U3890 (N_3890,N_2389,N_2967);
and U3891 (N_3891,N_2331,N_2054);
or U3892 (N_3892,N_2733,N_2836);
and U3893 (N_3893,N_2265,N_2240);
nand U3894 (N_3894,N_2196,N_2128);
nor U3895 (N_3895,N_2483,N_2791);
or U3896 (N_3896,N_2563,N_2978);
nand U3897 (N_3897,N_2028,N_2493);
nand U3898 (N_3898,N_2463,N_2490);
nor U3899 (N_3899,N_2716,N_2387);
nand U3900 (N_3900,N_2510,N_2316);
and U3901 (N_3901,N_2481,N_2115);
and U3902 (N_3902,N_2822,N_2567);
and U3903 (N_3903,N_2341,N_2130);
or U3904 (N_3904,N_2977,N_2072);
nand U3905 (N_3905,N_2822,N_2176);
or U3906 (N_3906,N_2793,N_2773);
nor U3907 (N_3907,N_2820,N_2520);
and U3908 (N_3908,N_2721,N_2146);
xor U3909 (N_3909,N_2105,N_2153);
or U3910 (N_3910,N_2305,N_2698);
nor U3911 (N_3911,N_2068,N_2906);
nor U3912 (N_3912,N_2926,N_2248);
and U3913 (N_3913,N_2606,N_2769);
and U3914 (N_3914,N_2444,N_2505);
or U3915 (N_3915,N_2751,N_2862);
or U3916 (N_3916,N_2203,N_2602);
nor U3917 (N_3917,N_2581,N_2009);
xor U3918 (N_3918,N_2953,N_2545);
xnor U3919 (N_3919,N_2711,N_2892);
xor U3920 (N_3920,N_2960,N_2881);
xor U3921 (N_3921,N_2304,N_2133);
nor U3922 (N_3922,N_2670,N_2494);
or U3923 (N_3923,N_2006,N_2952);
nor U3924 (N_3924,N_2243,N_2833);
nand U3925 (N_3925,N_2886,N_2574);
nand U3926 (N_3926,N_2587,N_2065);
or U3927 (N_3927,N_2717,N_2091);
and U3928 (N_3928,N_2184,N_2426);
nor U3929 (N_3929,N_2693,N_2892);
nor U3930 (N_3930,N_2414,N_2796);
and U3931 (N_3931,N_2082,N_2475);
nand U3932 (N_3932,N_2994,N_2874);
nor U3933 (N_3933,N_2323,N_2222);
and U3934 (N_3934,N_2384,N_2724);
and U3935 (N_3935,N_2035,N_2126);
nor U3936 (N_3936,N_2620,N_2212);
xnor U3937 (N_3937,N_2403,N_2682);
and U3938 (N_3938,N_2243,N_2446);
nand U3939 (N_3939,N_2980,N_2467);
nand U3940 (N_3940,N_2588,N_2065);
xnor U3941 (N_3941,N_2640,N_2103);
or U3942 (N_3942,N_2977,N_2272);
nor U3943 (N_3943,N_2078,N_2972);
nor U3944 (N_3944,N_2319,N_2936);
nor U3945 (N_3945,N_2146,N_2465);
or U3946 (N_3946,N_2934,N_2259);
and U3947 (N_3947,N_2307,N_2939);
xnor U3948 (N_3948,N_2017,N_2925);
or U3949 (N_3949,N_2142,N_2640);
and U3950 (N_3950,N_2305,N_2574);
or U3951 (N_3951,N_2433,N_2212);
nand U3952 (N_3952,N_2297,N_2972);
and U3953 (N_3953,N_2098,N_2135);
or U3954 (N_3954,N_2408,N_2056);
and U3955 (N_3955,N_2615,N_2192);
nand U3956 (N_3956,N_2399,N_2125);
xor U3957 (N_3957,N_2821,N_2077);
nor U3958 (N_3958,N_2018,N_2869);
or U3959 (N_3959,N_2671,N_2261);
and U3960 (N_3960,N_2314,N_2866);
nand U3961 (N_3961,N_2521,N_2585);
nand U3962 (N_3962,N_2291,N_2237);
and U3963 (N_3963,N_2499,N_2243);
nand U3964 (N_3964,N_2051,N_2084);
nand U3965 (N_3965,N_2783,N_2767);
nor U3966 (N_3966,N_2458,N_2665);
and U3967 (N_3967,N_2179,N_2648);
xor U3968 (N_3968,N_2656,N_2093);
and U3969 (N_3969,N_2177,N_2203);
nand U3970 (N_3970,N_2044,N_2590);
nor U3971 (N_3971,N_2133,N_2297);
or U3972 (N_3972,N_2779,N_2083);
xnor U3973 (N_3973,N_2552,N_2598);
nor U3974 (N_3974,N_2314,N_2548);
nor U3975 (N_3975,N_2899,N_2882);
or U3976 (N_3976,N_2527,N_2690);
and U3977 (N_3977,N_2984,N_2978);
or U3978 (N_3978,N_2532,N_2613);
nand U3979 (N_3979,N_2576,N_2510);
and U3980 (N_3980,N_2405,N_2243);
or U3981 (N_3981,N_2662,N_2162);
nand U3982 (N_3982,N_2236,N_2757);
nor U3983 (N_3983,N_2719,N_2381);
nand U3984 (N_3984,N_2126,N_2452);
nand U3985 (N_3985,N_2014,N_2666);
and U3986 (N_3986,N_2127,N_2586);
and U3987 (N_3987,N_2800,N_2599);
or U3988 (N_3988,N_2170,N_2990);
xor U3989 (N_3989,N_2942,N_2033);
nand U3990 (N_3990,N_2604,N_2097);
nor U3991 (N_3991,N_2352,N_2103);
nor U3992 (N_3992,N_2382,N_2862);
or U3993 (N_3993,N_2135,N_2315);
xor U3994 (N_3994,N_2351,N_2185);
nor U3995 (N_3995,N_2949,N_2449);
nor U3996 (N_3996,N_2340,N_2946);
nor U3997 (N_3997,N_2303,N_2211);
nand U3998 (N_3998,N_2238,N_2527);
or U3999 (N_3999,N_2419,N_2922);
nand U4000 (N_4000,N_3909,N_3341);
or U4001 (N_4001,N_3420,N_3316);
and U4002 (N_4002,N_3499,N_3588);
nor U4003 (N_4003,N_3819,N_3919);
and U4004 (N_4004,N_3167,N_3201);
and U4005 (N_4005,N_3490,N_3014);
nand U4006 (N_4006,N_3993,N_3708);
nor U4007 (N_4007,N_3905,N_3112);
nand U4008 (N_4008,N_3711,N_3918);
nor U4009 (N_4009,N_3094,N_3268);
and U4010 (N_4010,N_3569,N_3109);
or U4011 (N_4011,N_3678,N_3850);
and U4012 (N_4012,N_3320,N_3346);
xor U4013 (N_4013,N_3326,N_3968);
and U4014 (N_4014,N_3342,N_3706);
xnor U4015 (N_4015,N_3441,N_3432);
nand U4016 (N_4016,N_3923,N_3438);
and U4017 (N_4017,N_3592,N_3925);
or U4018 (N_4018,N_3748,N_3895);
nand U4019 (N_4019,N_3257,N_3104);
nand U4020 (N_4020,N_3469,N_3952);
xnor U4021 (N_4021,N_3744,N_3428);
or U4022 (N_4022,N_3681,N_3127);
nand U4023 (N_4023,N_3026,N_3194);
or U4024 (N_4024,N_3457,N_3259);
xnor U4025 (N_4025,N_3983,N_3037);
nor U4026 (N_4026,N_3199,N_3373);
nand U4027 (N_4027,N_3817,N_3862);
or U4028 (N_4028,N_3833,N_3097);
or U4029 (N_4029,N_3690,N_3527);
xnor U4030 (N_4030,N_3989,N_3178);
nand U4031 (N_4031,N_3377,N_3791);
or U4032 (N_4032,N_3726,N_3639);
or U4033 (N_4033,N_3138,N_3205);
and U4034 (N_4034,N_3736,N_3020);
xor U4035 (N_4035,N_3656,N_3828);
and U4036 (N_4036,N_3296,N_3787);
nand U4037 (N_4037,N_3766,N_3579);
nor U4038 (N_4038,N_3019,N_3657);
nor U4039 (N_4039,N_3075,N_3660);
nand U4040 (N_4040,N_3928,N_3006);
and U4041 (N_4041,N_3635,N_3816);
or U4042 (N_4042,N_3714,N_3630);
xor U4043 (N_4043,N_3841,N_3000);
and U4044 (N_4044,N_3891,N_3016);
xor U4045 (N_4045,N_3688,N_3760);
and U4046 (N_4046,N_3480,N_3260);
nor U4047 (N_4047,N_3735,N_3548);
or U4048 (N_4048,N_3506,N_3276);
or U4049 (N_4049,N_3815,N_3699);
and U4050 (N_4050,N_3572,N_3849);
nor U4051 (N_4051,N_3088,N_3466);
xnor U4052 (N_4052,N_3519,N_3429);
and U4053 (N_4053,N_3907,N_3315);
nand U4054 (N_4054,N_3482,N_3289);
and U4055 (N_4055,N_3526,N_3576);
nand U4056 (N_4056,N_3293,N_3874);
nor U4057 (N_4057,N_3436,N_3624);
nand U4058 (N_4058,N_3483,N_3876);
nand U4059 (N_4059,N_3210,N_3970);
nor U4060 (N_4060,N_3219,N_3700);
and U4061 (N_4061,N_3421,N_3434);
or U4062 (N_4062,N_3901,N_3514);
and U4063 (N_4063,N_3414,N_3050);
and U4064 (N_4064,N_3879,N_3486);
and U4065 (N_4065,N_3118,N_3800);
or U4066 (N_4066,N_3374,N_3637);
and U4067 (N_4067,N_3803,N_3213);
xnor U4068 (N_4068,N_3134,N_3324);
or U4069 (N_4069,N_3299,N_3504);
nor U4070 (N_4070,N_3021,N_3236);
nor U4071 (N_4071,N_3033,N_3369);
or U4072 (N_4072,N_3991,N_3540);
and U4073 (N_4073,N_3730,N_3971);
or U4074 (N_4074,N_3944,N_3206);
nor U4075 (N_4075,N_3193,N_3647);
nand U4076 (N_4076,N_3757,N_3687);
nor U4077 (N_4077,N_3858,N_3180);
and U4078 (N_4078,N_3645,N_3155);
or U4079 (N_4079,N_3007,N_3521);
xor U4080 (N_4080,N_3468,N_3012);
nand U4081 (N_4081,N_3055,N_3812);
or U4082 (N_4082,N_3843,N_3488);
nand U4083 (N_4083,N_3059,N_3930);
nor U4084 (N_4084,N_3545,N_3798);
or U4085 (N_4085,N_3185,N_3638);
or U4086 (N_4086,N_3286,N_3023);
nand U4087 (N_4087,N_3826,N_3424);
nor U4088 (N_4088,N_3752,N_3753);
xor U4089 (N_4089,N_3463,N_3068);
nor U4090 (N_4090,N_3776,N_3237);
nor U4091 (N_4091,N_3847,N_3011);
and U4092 (N_4092,N_3336,N_3724);
nor U4093 (N_4093,N_3216,N_3875);
nand U4094 (N_4094,N_3543,N_3518);
nand U4095 (N_4095,N_3394,N_3158);
and U4096 (N_4096,N_3444,N_3982);
xor U4097 (N_4097,N_3285,N_3973);
nor U4098 (N_4098,N_3080,N_3433);
or U4099 (N_4099,N_3121,N_3387);
nor U4100 (N_4100,N_3004,N_3261);
xnor U4101 (N_4101,N_3830,N_3651);
nand U4102 (N_4102,N_3946,N_3427);
nand U4103 (N_4103,N_3595,N_3380);
nand U4104 (N_4104,N_3529,N_3115);
nor U4105 (N_4105,N_3042,N_3298);
nand U4106 (N_4106,N_3198,N_3084);
and U4107 (N_4107,N_3462,N_3120);
nor U4108 (N_4108,N_3208,N_3620);
or U4109 (N_4109,N_3673,N_3090);
nand U4110 (N_4110,N_3101,N_3265);
or U4111 (N_4111,N_3805,N_3510);
and U4112 (N_4112,N_3732,N_3797);
or U4113 (N_4113,N_3069,N_3790);
or U4114 (N_4114,N_3857,N_3415);
or U4115 (N_4115,N_3773,N_3203);
xnor U4116 (N_4116,N_3937,N_3263);
or U4117 (N_4117,N_3535,N_3470);
and U4118 (N_4118,N_3739,N_3751);
nand U4119 (N_4119,N_3074,N_3562);
and U4120 (N_4120,N_3684,N_3940);
nand U4121 (N_4121,N_3606,N_3741);
or U4122 (N_4122,N_3402,N_3386);
and U4123 (N_4123,N_3984,N_3966);
or U4124 (N_4124,N_3253,N_3099);
or U4125 (N_4125,N_3912,N_3935);
and U4126 (N_4126,N_3956,N_3036);
xnor U4127 (N_4127,N_3052,N_3852);
and U4128 (N_4128,N_3939,N_3931);
or U4129 (N_4129,N_3996,N_3917);
or U4130 (N_4130,N_3453,N_3372);
or U4131 (N_4131,N_3487,N_3654);
and U4132 (N_4132,N_3903,N_3856);
nor U4133 (N_4133,N_3631,N_3494);
or U4134 (N_4134,N_3029,N_3008);
or U4135 (N_4135,N_3132,N_3418);
or U4136 (N_4136,N_3948,N_3929);
nor U4137 (N_4137,N_3327,N_3695);
nand U4138 (N_4138,N_3593,N_3169);
and U4139 (N_4139,N_3742,N_3615);
xor U4140 (N_4140,N_3191,N_3611);
nor U4141 (N_4141,N_3370,N_3904);
xnor U4142 (N_4142,N_3517,N_3566);
and U4143 (N_4143,N_3822,N_3239);
and U4144 (N_4144,N_3192,N_3310);
and U4145 (N_4145,N_3622,N_3933);
and U4146 (N_4146,N_3683,N_3953);
and U4147 (N_4147,N_3211,N_3788);
nand U4148 (N_4148,N_3995,N_3422);
xor U4149 (N_4149,N_3765,N_3568);
and U4150 (N_4150,N_3291,N_3117);
xor U4151 (N_4151,N_3333,N_3671);
or U4152 (N_4152,N_3783,N_3135);
or U4153 (N_4153,N_3598,N_3458);
xnor U4154 (N_4154,N_3794,N_3682);
xnor U4155 (N_4155,N_3809,N_3039);
xor U4156 (N_4156,N_3362,N_3172);
or U4157 (N_4157,N_3652,N_3570);
or U4158 (N_4158,N_3183,N_3799);
nand U4159 (N_4159,N_3754,N_3962);
and U4160 (N_4160,N_3523,N_3743);
nor U4161 (N_4161,N_3212,N_3943);
nor U4162 (N_4162,N_3703,N_3449);
nor U4163 (N_4163,N_3044,N_3159);
nand U4164 (N_4164,N_3366,N_3778);
and U4165 (N_4165,N_3848,N_3057);
nor U4166 (N_4166,N_3792,N_3391);
and U4167 (N_4167,N_3564,N_3580);
nand U4168 (N_4168,N_3475,N_3668);
and U4169 (N_4169,N_3911,N_3698);
nor U4170 (N_4170,N_3873,N_3575);
nor U4171 (N_4171,N_3869,N_3149);
nor U4172 (N_4172,N_3028,N_3240);
nor U4173 (N_4173,N_3417,N_3345);
or U4174 (N_4174,N_3758,N_3017);
xor U4175 (N_4175,N_3725,N_3602);
and U4176 (N_4176,N_3784,N_3662);
or U4177 (N_4177,N_3329,N_3279);
nor U4178 (N_4178,N_3802,N_3536);
nor U4179 (N_4179,N_3785,N_3245);
or U4180 (N_4180,N_3426,N_3610);
or U4181 (N_4181,N_3142,N_3507);
or U4182 (N_4182,N_3061,N_3077);
and U4183 (N_4183,N_3425,N_3764);
nor U4184 (N_4184,N_3309,N_3209);
and U4185 (N_4185,N_3031,N_3133);
or U4186 (N_4186,N_3886,N_3186);
and U4187 (N_4187,N_3269,N_3632);
nor U4188 (N_4188,N_3073,N_3947);
and U4189 (N_4189,N_3275,N_3339);
xnor U4190 (N_4190,N_3001,N_3363);
nand U4191 (N_4191,N_3640,N_3877);
nand U4192 (N_4192,N_3087,N_3998);
or U4193 (N_4193,N_3095,N_3950);
and U4194 (N_4194,N_3447,N_3492);
nand U4195 (N_4195,N_3675,N_3160);
or U4196 (N_4196,N_3823,N_3957);
or U4197 (N_4197,N_3539,N_3493);
nor U4198 (N_4198,N_3844,N_3405);
nand U4199 (N_4199,N_3705,N_3137);
or U4200 (N_4200,N_3623,N_3801);
and U4201 (N_4201,N_3646,N_3516);
xnor U4202 (N_4202,N_3251,N_3078);
nand U4203 (N_4203,N_3053,N_3379);
and U4204 (N_4204,N_3601,N_3878);
or U4205 (N_4205,N_3247,N_3174);
xor U4206 (N_4206,N_3018,N_3262);
nand U4207 (N_4207,N_3252,N_3608);
nand U4208 (N_4208,N_3560,N_3283);
or U4209 (N_4209,N_3614,N_3025);
nor U4210 (N_4210,N_3556,N_3184);
xnor U4211 (N_4211,N_3508,N_3596);
xor U4212 (N_4212,N_3655,N_3454);
and U4213 (N_4213,N_3300,N_3795);
nand U4214 (N_4214,N_3367,N_3416);
nand U4215 (N_4215,N_3997,N_3577);
nand U4216 (N_4216,N_3024,N_3837);
and U4217 (N_4217,N_3888,N_3491);
or U4218 (N_4218,N_3164,N_3071);
nor U4219 (N_4219,N_3578,N_3489);
and U4220 (N_4220,N_3308,N_3332);
nor U4221 (N_4221,N_3430,N_3274);
and U4222 (N_4222,N_3062,N_3520);
nand U4223 (N_4223,N_3388,N_3464);
nor U4224 (N_4224,N_3663,N_3607);
nand U4225 (N_4225,N_3824,N_3719);
nand U4226 (N_4226,N_3119,N_3270);
nand U4227 (N_4227,N_3162,N_3472);
nor U4228 (N_4228,N_3235,N_3894);
nor U4229 (N_4229,N_3188,N_3603);
nand U4230 (N_4230,N_3932,N_3148);
xor U4231 (N_4231,N_3958,N_3584);
nor U4232 (N_4232,N_3451,N_3461);
nand U4233 (N_4233,N_3406,N_3152);
nor U4234 (N_4234,N_3963,N_3108);
nand U4235 (N_4235,N_3229,N_3474);
nor U4236 (N_4236,N_3140,N_3035);
and U4237 (N_4237,N_3243,N_3027);
or U4238 (N_4238,N_3716,N_3244);
nor U4239 (N_4239,N_3256,N_3272);
or U4240 (N_4240,N_3513,N_3410);
and U4241 (N_4241,N_3818,N_3717);
nand U4242 (N_4242,N_3335,N_3022);
or U4243 (N_4243,N_3043,N_3156);
nor U4244 (N_4244,N_3459,N_3880);
or U4245 (N_4245,N_3648,N_3642);
nand U4246 (N_4246,N_3034,N_3910);
or U4247 (N_4247,N_3634,N_3343);
or U4248 (N_4248,N_3288,N_3547);
and U4249 (N_4249,N_3955,N_3522);
xnor U4250 (N_4250,N_3157,N_3173);
nand U4251 (N_4251,N_3103,N_3302);
or U4252 (N_4252,N_3181,N_3479);
and U4253 (N_4253,N_3702,N_3839);
nor U4254 (N_4254,N_3146,N_3954);
nand U4255 (N_4255,N_3450,N_3829);
nor U4256 (N_4256,N_3718,N_3538);
nand U4257 (N_4257,N_3189,N_3038);
and U4258 (N_4258,N_3446,N_3927);
nand U4259 (N_4259,N_3694,N_3002);
xor U4260 (N_4260,N_3495,N_3759);
nand U4261 (N_4261,N_3728,N_3756);
and U4262 (N_4262,N_3864,N_3860);
and U4263 (N_4263,N_3613,N_3281);
nand U4264 (N_4264,N_3769,N_3820);
or U4265 (N_4265,N_3267,N_3460);
nor U4266 (N_4266,N_3225,N_3636);
and U4267 (N_4267,N_3303,N_3419);
nor U4268 (N_4268,N_3297,N_3644);
nor U4269 (N_4269,N_3533,N_3175);
xor U4270 (N_4270,N_3060,N_3524);
nand U4271 (N_4271,N_3107,N_3782);
xnor U4272 (N_4272,N_3553,N_3915);
or U4273 (N_4273,N_3431,N_3807);
and U4274 (N_4274,N_3177,N_3354);
nand U4275 (N_4275,N_3808,N_3273);
nor U4276 (N_4276,N_3814,N_3571);
or U4277 (N_4277,N_3665,N_3977);
and U4278 (N_4278,N_3980,N_3629);
nand U4279 (N_4279,N_3842,N_3664);
nor U4280 (N_4280,N_3355,N_3804);
and U4281 (N_4281,N_3128,N_3246);
xnor U4282 (N_4282,N_3770,N_3666);
nand U4283 (N_4283,N_3054,N_3774);
nor U4284 (N_4284,N_3314,N_3122);
xnor U4285 (N_4285,N_3563,N_3945);
nand U4286 (N_4286,N_3081,N_3999);
and U4287 (N_4287,N_3290,N_3365);
nor U4288 (N_4288,N_3621,N_3241);
and U4289 (N_4289,N_3222,N_3565);
xor U4290 (N_4290,N_3693,N_3448);
nor U4291 (N_4291,N_3897,N_3992);
xnor U4292 (N_4292,N_3264,N_3767);
or U4293 (N_4293,N_3126,N_3961);
nand U4294 (N_4294,N_3301,N_3171);
nand U4295 (N_4295,N_3473,N_3452);
nor U4296 (N_4296,N_3746,N_3686);
nand U4297 (N_4297,N_3599,N_3412);
nand U4298 (N_4298,N_3658,N_3627);
or U4299 (N_4299,N_3478,N_3885);
nor U4300 (N_4300,N_3249,N_3129);
or U4301 (N_4301,N_3361,N_3887);
and U4302 (N_4302,N_3922,N_3707);
and U4303 (N_4303,N_3105,N_3985);
xor U4304 (N_4304,N_3124,N_3582);
nor U4305 (N_4305,N_3145,N_3938);
nor U4306 (N_4306,N_3093,N_3916);
nand U4307 (N_4307,N_3967,N_3626);
nand U4308 (N_4308,N_3040,N_3195);
and U4309 (N_4309,N_3233,N_3845);
nand U4310 (N_4310,N_3015,N_3277);
and U4311 (N_4311,N_3628,N_3960);
or U4312 (N_4312,N_3009,N_3975);
and U4313 (N_4313,N_3381,N_3846);
nor U4314 (N_4314,N_3976,N_3509);
and U4315 (N_4315,N_3248,N_3633);
nor U4316 (N_4316,N_3356,N_3619);
and U4317 (N_4317,N_3650,N_3914);
and U4318 (N_4318,N_3284,N_3352);
nand U4319 (N_4319,N_3677,N_3498);
nand U4320 (N_4320,N_3340,N_3051);
and U4321 (N_4321,N_3515,N_3806);
and U4322 (N_4322,N_3541,N_3853);
nand U4323 (N_4323,N_3072,N_3691);
or U4324 (N_4324,N_3542,N_3319);
nand U4325 (N_4325,N_3723,N_3322);
and U4326 (N_4326,N_3041,N_3854);
nor U4327 (N_4327,N_3200,N_3079);
or U4328 (N_4328,N_3223,N_3397);
nand U4329 (N_4329,N_3359,N_3411);
nor U4330 (N_4330,N_3749,N_3066);
and U4331 (N_4331,N_3046,N_3147);
or U4332 (N_4332,N_3476,N_3685);
nand U4333 (N_4333,N_3064,N_3585);
nor U4334 (N_4334,N_3368,N_3859);
nand U4335 (N_4335,N_3583,N_3182);
nor U4336 (N_4336,N_3537,N_3437);
nand U4337 (N_4337,N_3959,N_3697);
nand U4338 (N_4338,N_3737,N_3768);
or U4339 (N_4339,N_3835,N_3501);
nor U4340 (N_4340,N_3005,N_3196);
and U4341 (N_4341,N_3554,N_3278);
and U4342 (N_4342,N_3242,N_3396);
or U4343 (N_4343,N_3170,N_3231);
or U4344 (N_4344,N_3400,N_3065);
and U4345 (N_4345,N_3550,N_3990);
nand U4346 (N_4346,N_3465,N_3546);
or U4347 (N_4347,N_3594,N_3643);
or U4348 (N_4348,N_3825,N_3720);
or U4349 (N_4349,N_3154,N_3435);
nor U4350 (N_4350,N_3131,N_3204);
and U4351 (N_4351,N_3867,N_3969);
nand U4352 (N_4352,N_3389,N_3500);
nand U4353 (N_4353,N_3111,N_3789);
nand U4354 (N_4354,N_3713,N_3098);
nand U4355 (N_4355,N_3821,N_3317);
nor U4356 (N_4356,N_3729,N_3612);
or U4357 (N_4357,N_3763,N_3832);
xor U4358 (N_4358,N_3512,N_3941);
and U4359 (N_4359,N_3734,N_3924);
nand U4360 (N_4360,N_3680,N_3777);
nand U4361 (N_4361,N_3618,N_3573);
and U4362 (N_4362,N_3331,N_3559);
and U4363 (N_4363,N_3965,N_3130);
and U4364 (N_4364,N_3392,N_3793);
nand U4365 (N_4365,N_3926,N_3271);
nor U4366 (N_4366,N_3401,N_3557);
xor U4367 (N_4367,N_3382,N_3979);
or U4368 (N_4368,N_3871,N_3395);
or U4369 (N_4369,N_3591,N_3906);
nand U4370 (N_4370,N_3813,N_3964);
nand U4371 (N_4371,N_3836,N_3951);
and U4372 (N_4372,N_3344,N_3348);
or U4373 (N_4373,N_3772,N_3653);
nor U4374 (N_4374,N_3889,N_3709);
or U4375 (N_4375,N_3827,N_3399);
nor U4376 (N_4376,N_3013,N_3375);
nor U4377 (N_4377,N_3481,N_3771);
and U4378 (N_4378,N_3398,N_3669);
nor U4379 (N_4379,N_3731,N_3384);
nand U4380 (N_4380,N_3692,N_3338);
nor U4381 (N_4381,N_3534,N_3704);
nor U4382 (N_4382,N_3761,N_3861);
or U4383 (N_4383,N_3376,N_3715);
nor U4384 (N_4384,N_3230,N_3502);
xor U4385 (N_4385,N_3030,N_3385);
xnor U4386 (N_4386,N_3218,N_3661);
or U4387 (N_4387,N_3641,N_3551);
xnor U4388 (N_4388,N_3558,N_3987);
nand U4389 (N_4389,N_3544,N_3934);
or U4390 (N_4390,N_3780,N_3407);
and U4391 (N_4391,N_3221,N_3232);
nor U4392 (N_4392,N_3304,N_3351);
or U4393 (N_4393,N_3091,N_3913);
and U4394 (N_4394,N_3295,N_3738);
and U4395 (N_4395,N_3306,N_3161);
nor U4396 (N_4396,N_3307,N_3899);
nor U4397 (N_4397,N_3727,N_3589);
nor U4398 (N_4398,N_3755,N_3092);
nor U4399 (N_4399,N_3532,N_3949);
or U4400 (N_4400,N_3561,N_3371);
nand U4401 (N_4401,N_3740,N_3113);
nand U4402 (N_4402,N_3383,N_3667);
or U4403 (N_4403,N_3503,N_3337);
xor U4404 (N_4404,N_3674,N_3360);
nor U4405 (N_4405,N_3831,N_3136);
nor U4406 (N_4406,N_3555,N_3328);
or U4407 (N_4407,N_3010,N_3974);
nand U4408 (N_4408,N_3202,N_3586);
and U4409 (N_4409,N_3868,N_3893);
or U4410 (N_4410,N_3689,N_3851);
or U4411 (N_4411,N_3936,N_3838);
nor U4412 (N_4412,N_3102,N_3207);
and U4413 (N_4413,N_3139,N_3549);
or U4414 (N_4414,N_3762,N_3505);
xnor U4415 (N_4415,N_3659,N_3921);
nor U4416 (N_4416,N_3456,N_3311);
nand U4417 (N_4417,N_3892,N_3292);
nand U4418 (N_4418,N_3781,N_3810);
and U4419 (N_4419,N_3679,N_3165);
nor U4420 (N_4420,N_3445,N_3153);
or U4421 (N_4421,N_3439,N_3811);
and U4422 (N_4422,N_3581,N_3605);
nand U4423 (N_4423,N_3866,N_3525);
xor U4424 (N_4424,N_3413,N_3305);
nand U4425 (N_4425,N_3076,N_3393);
or U4426 (N_4426,N_3485,N_3123);
nor U4427 (N_4427,N_3323,N_3220);
nor U4428 (N_4428,N_3423,N_3168);
and U4429 (N_4429,N_3350,N_3063);
nor U4430 (N_4430,N_3179,N_3321);
nand U4431 (N_4431,N_3676,N_3471);
or U4432 (N_4432,N_3250,N_3358);
nand U4433 (N_4433,N_3215,N_3883);
nor U4434 (N_4434,N_3779,N_3881);
nand U4435 (N_4435,N_3003,N_3442);
and U4436 (N_4436,N_3187,N_3313);
and U4437 (N_4437,N_3390,N_3511);
xor U4438 (N_4438,N_3443,N_3287);
or U4439 (N_4439,N_3047,N_3528);
xor U4440 (N_4440,N_3884,N_3214);
or U4441 (N_4441,N_3409,N_3455);
nand U4442 (N_4442,N_3190,N_3865);
xnor U4443 (N_4443,N_3144,N_3086);
and U4444 (N_4444,N_3349,N_3334);
or U4445 (N_4445,N_3604,N_3151);
nor U4446 (N_4446,N_3609,N_3477);
xor U4447 (N_4447,N_3227,N_3312);
nand U4448 (N_4448,N_3786,N_3114);
or U4449 (N_4449,N_3357,N_3353);
nor U4450 (N_4450,N_3531,N_3110);
and U4451 (N_4451,N_3364,N_3497);
nand U4452 (N_4452,N_3747,N_3085);
nand U4453 (N_4453,N_3403,N_3408);
or U4454 (N_4454,N_3067,N_3141);
nor U4455 (N_4455,N_3670,N_3942);
or U4456 (N_4456,N_3855,N_3587);
nor U4457 (N_4457,N_3294,N_3710);
nor U4458 (N_4458,N_3840,N_3176);
or U4459 (N_4459,N_3902,N_3404);
or U4460 (N_4460,N_3280,N_3625);
or U4461 (N_4461,N_3863,N_3721);
nor U4462 (N_4462,N_3986,N_3890);
and U4463 (N_4463,N_3070,N_3745);
or U4464 (N_4464,N_3872,N_3045);
or U4465 (N_4465,N_3701,N_3150);
and U4466 (N_4466,N_3981,N_3056);
and U4467 (N_4467,N_3282,N_3994);
nor U4468 (N_4468,N_3896,N_3258);
and U4469 (N_4469,N_3567,N_3775);
nor U4470 (N_4470,N_3143,N_3796);
nor U4471 (N_4471,N_3224,N_3106);
xor U4472 (N_4472,N_3590,N_3217);
nor U4473 (N_4473,N_3197,N_3834);
nand U4474 (N_4474,N_3882,N_3898);
nand U4475 (N_4475,N_3616,N_3318);
or U4476 (N_4476,N_3496,N_3096);
xnor U4477 (N_4477,N_3440,N_3574);
and U4478 (N_4478,N_3920,N_3750);
nand U4479 (N_4479,N_3325,N_3082);
xor U4480 (N_4480,N_3600,N_3238);
nor U4481 (N_4481,N_3722,N_3467);
nand U4482 (N_4482,N_3330,N_3672);
or U4483 (N_4483,N_3552,N_3972);
and U4484 (N_4484,N_3978,N_3163);
and U4485 (N_4485,N_3712,N_3484);
nor U4486 (N_4486,N_3228,N_3649);
and U4487 (N_4487,N_3733,N_3089);
nand U4488 (N_4488,N_3988,N_3908);
nor U4489 (N_4489,N_3617,N_3116);
nand U4490 (N_4490,N_3058,N_3166);
and U4491 (N_4491,N_3226,N_3048);
nand U4492 (N_4492,N_3255,N_3900);
or U4493 (N_4493,N_3696,N_3049);
nor U4494 (N_4494,N_3378,N_3032);
xor U4495 (N_4495,N_3530,N_3100);
nor U4496 (N_4496,N_3266,N_3125);
nor U4497 (N_4497,N_3083,N_3254);
nor U4498 (N_4498,N_3347,N_3870);
or U4499 (N_4499,N_3234,N_3597);
and U4500 (N_4500,N_3862,N_3682);
xor U4501 (N_4501,N_3755,N_3651);
nand U4502 (N_4502,N_3218,N_3884);
and U4503 (N_4503,N_3940,N_3782);
and U4504 (N_4504,N_3065,N_3076);
or U4505 (N_4505,N_3247,N_3754);
or U4506 (N_4506,N_3919,N_3019);
nand U4507 (N_4507,N_3684,N_3936);
xnor U4508 (N_4508,N_3122,N_3129);
nand U4509 (N_4509,N_3847,N_3462);
or U4510 (N_4510,N_3751,N_3215);
and U4511 (N_4511,N_3517,N_3585);
and U4512 (N_4512,N_3969,N_3035);
nand U4513 (N_4513,N_3534,N_3879);
nand U4514 (N_4514,N_3567,N_3398);
nand U4515 (N_4515,N_3190,N_3269);
nand U4516 (N_4516,N_3715,N_3252);
and U4517 (N_4517,N_3327,N_3736);
nand U4518 (N_4518,N_3774,N_3975);
or U4519 (N_4519,N_3555,N_3177);
and U4520 (N_4520,N_3109,N_3408);
and U4521 (N_4521,N_3487,N_3209);
or U4522 (N_4522,N_3837,N_3526);
nor U4523 (N_4523,N_3793,N_3632);
and U4524 (N_4524,N_3652,N_3642);
nand U4525 (N_4525,N_3908,N_3728);
or U4526 (N_4526,N_3114,N_3661);
nand U4527 (N_4527,N_3625,N_3049);
and U4528 (N_4528,N_3747,N_3073);
nand U4529 (N_4529,N_3929,N_3043);
nand U4530 (N_4530,N_3181,N_3303);
or U4531 (N_4531,N_3532,N_3144);
nor U4532 (N_4532,N_3252,N_3756);
and U4533 (N_4533,N_3659,N_3361);
nand U4534 (N_4534,N_3083,N_3087);
xnor U4535 (N_4535,N_3658,N_3143);
nor U4536 (N_4536,N_3021,N_3611);
nor U4537 (N_4537,N_3569,N_3692);
and U4538 (N_4538,N_3070,N_3227);
nor U4539 (N_4539,N_3669,N_3254);
nand U4540 (N_4540,N_3958,N_3722);
and U4541 (N_4541,N_3413,N_3476);
and U4542 (N_4542,N_3499,N_3092);
nand U4543 (N_4543,N_3731,N_3568);
and U4544 (N_4544,N_3673,N_3626);
nand U4545 (N_4545,N_3967,N_3177);
nand U4546 (N_4546,N_3327,N_3495);
and U4547 (N_4547,N_3395,N_3488);
and U4548 (N_4548,N_3005,N_3432);
and U4549 (N_4549,N_3861,N_3614);
xor U4550 (N_4550,N_3768,N_3266);
and U4551 (N_4551,N_3232,N_3547);
nand U4552 (N_4552,N_3866,N_3059);
nand U4553 (N_4553,N_3010,N_3779);
nand U4554 (N_4554,N_3055,N_3964);
nor U4555 (N_4555,N_3633,N_3553);
nor U4556 (N_4556,N_3797,N_3542);
nor U4557 (N_4557,N_3556,N_3952);
nor U4558 (N_4558,N_3727,N_3099);
nand U4559 (N_4559,N_3819,N_3610);
nand U4560 (N_4560,N_3783,N_3638);
xnor U4561 (N_4561,N_3781,N_3687);
and U4562 (N_4562,N_3900,N_3609);
and U4563 (N_4563,N_3141,N_3189);
nand U4564 (N_4564,N_3320,N_3364);
nor U4565 (N_4565,N_3368,N_3144);
or U4566 (N_4566,N_3259,N_3640);
xor U4567 (N_4567,N_3277,N_3511);
nor U4568 (N_4568,N_3966,N_3505);
nor U4569 (N_4569,N_3703,N_3145);
nor U4570 (N_4570,N_3587,N_3528);
nand U4571 (N_4571,N_3229,N_3670);
nand U4572 (N_4572,N_3789,N_3543);
nand U4573 (N_4573,N_3720,N_3237);
or U4574 (N_4574,N_3556,N_3727);
nor U4575 (N_4575,N_3515,N_3538);
nand U4576 (N_4576,N_3756,N_3549);
or U4577 (N_4577,N_3175,N_3559);
nor U4578 (N_4578,N_3429,N_3267);
or U4579 (N_4579,N_3312,N_3896);
nand U4580 (N_4580,N_3288,N_3379);
nor U4581 (N_4581,N_3114,N_3663);
and U4582 (N_4582,N_3967,N_3934);
and U4583 (N_4583,N_3779,N_3345);
and U4584 (N_4584,N_3122,N_3126);
and U4585 (N_4585,N_3643,N_3458);
nand U4586 (N_4586,N_3846,N_3368);
nor U4587 (N_4587,N_3246,N_3087);
nand U4588 (N_4588,N_3038,N_3197);
nand U4589 (N_4589,N_3970,N_3609);
or U4590 (N_4590,N_3189,N_3494);
and U4591 (N_4591,N_3469,N_3688);
nor U4592 (N_4592,N_3858,N_3770);
nand U4593 (N_4593,N_3977,N_3951);
nand U4594 (N_4594,N_3989,N_3742);
or U4595 (N_4595,N_3346,N_3967);
nand U4596 (N_4596,N_3120,N_3822);
and U4597 (N_4597,N_3526,N_3151);
or U4598 (N_4598,N_3460,N_3903);
and U4599 (N_4599,N_3438,N_3754);
and U4600 (N_4600,N_3845,N_3986);
nor U4601 (N_4601,N_3484,N_3705);
nor U4602 (N_4602,N_3129,N_3577);
xor U4603 (N_4603,N_3662,N_3076);
xnor U4604 (N_4604,N_3634,N_3222);
nor U4605 (N_4605,N_3697,N_3463);
nand U4606 (N_4606,N_3120,N_3324);
nand U4607 (N_4607,N_3967,N_3161);
and U4608 (N_4608,N_3063,N_3754);
or U4609 (N_4609,N_3822,N_3693);
nand U4610 (N_4610,N_3824,N_3027);
nor U4611 (N_4611,N_3219,N_3655);
nor U4612 (N_4612,N_3255,N_3299);
or U4613 (N_4613,N_3352,N_3062);
and U4614 (N_4614,N_3975,N_3115);
nor U4615 (N_4615,N_3170,N_3151);
or U4616 (N_4616,N_3704,N_3482);
nor U4617 (N_4617,N_3061,N_3432);
and U4618 (N_4618,N_3881,N_3823);
xor U4619 (N_4619,N_3401,N_3509);
nand U4620 (N_4620,N_3051,N_3570);
nor U4621 (N_4621,N_3045,N_3897);
nand U4622 (N_4622,N_3360,N_3065);
nor U4623 (N_4623,N_3387,N_3134);
or U4624 (N_4624,N_3652,N_3025);
nand U4625 (N_4625,N_3260,N_3385);
or U4626 (N_4626,N_3403,N_3983);
and U4627 (N_4627,N_3856,N_3533);
nand U4628 (N_4628,N_3304,N_3782);
or U4629 (N_4629,N_3693,N_3387);
or U4630 (N_4630,N_3289,N_3444);
nand U4631 (N_4631,N_3025,N_3323);
xnor U4632 (N_4632,N_3272,N_3622);
nor U4633 (N_4633,N_3850,N_3467);
or U4634 (N_4634,N_3610,N_3922);
nand U4635 (N_4635,N_3985,N_3777);
and U4636 (N_4636,N_3569,N_3182);
and U4637 (N_4637,N_3579,N_3796);
and U4638 (N_4638,N_3913,N_3031);
nand U4639 (N_4639,N_3134,N_3101);
nor U4640 (N_4640,N_3923,N_3358);
and U4641 (N_4641,N_3806,N_3476);
and U4642 (N_4642,N_3850,N_3888);
or U4643 (N_4643,N_3389,N_3976);
nand U4644 (N_4644,N_3979,N_3670);
xnor U4645 (N_4645,N_3959,N_3804);
and U4646 (N_4646,N_3413,N_3519);
nor U4647 (N_4647,N_3319,N_3640);
nor U4648 (N_4648,N_3621,N_3171);
nor U4649 (N_4649,N_3896,N_3448);
nand U4650 (N_4650,N_3873,N_3280);
nor U4651 (N_4651,N_3372,N_3611);
or U4652 (N_4652,N_3381,N_3706);
and U4653 (N_4653,N_3787,N_3677);
or U4654 (N_4654,N_3507,N_3320);
or U4655 (N_4655,N_3235,N_3353);
nor U4656 (N_4656,N_3935,N_3412);
xnor U4657 (N_4657,N_3239,N_3105);
and U4658 (N_4658,N_3885,N_3752);
nor U4659 (N_4659,N_3230,N_3959);
or U4660 (N_4660,N_3824,N_3524);
xor U4661 (N_4661,N_3866,N_3328);
or U4662 (N_4662,N_3006,N_3289);
nand U4663 (N_4663,N_3752,N_3760);
or U4664 (N_4664,N_3262,N_3233);
or U4665 (N_4665,N_3037,N_3050);
xnor U4666 (N_4666,N_3715,N_3477);
or U4667 (N_4667,N_3044,N_3814);
and U4668 (N_4668,N_3174,N_3678);
nor U4669 (N_4669,N_3572,N_3952);
xor U4670 (N_4670,N_3576,N_3583);
or U4671 (N_4671,N_3164,N_3423);
nor U4672 (N_4672,N_3531,N_3350);
nor U4673 (N_4673,N_3942,N_3507);
and U4674 (N_4674,N_3977,N_3499);
nand U4675 (N_4675,N_3391,N_3921);
and U4676 (N_4676,N_3519,N_3638);
nand U4677 (N_4677,N_3541,N_3883);
nor U4678 (N_4678,N_3767,N_3178);
nand U4679 (N_4679,N_3186,N_3502);
and U4680 (N_4680,N_3898,N_3243);
nor U4681 (N_4681,N_3676,N_3012);
or U4682 (N_4682,N_3148,N_3132);
xnor U4683 (N_4683,N_3897,N_3635);
or U4684 (N_4684,N_3714,N_3233);
or U4685 (N_4685,N_3876,N_3510);
nand U4686 (N_4686,N_3485,N_3981);
or U4687 (N_4687,N_3352,N_3408);
xor U4688 (N_4688,N_3003,N_3144);
or U4689 (N_4689,N_3957,N_3897);
nand U4690 (N_4690,N_3224,N_3612);
or U4691 (N_4691,N_3183,N_3304);
nand U4692 (N_4692,N_3709,N_3190);
and U4693 (N_4693,N_3603,N_3965);
nand U4694 (N_4694,N_3463,N_3832);
nand U4695 (N_4695,N_3705,N_3345);
or U4696 (N_4696,N_3621,N_3615);
or U4697 (N_4697,N_3162,N_3901);
nor U4698 (N_4698,N_3308,N_3434);
nand U4699 (N_4699,N_3479,N_3754);
nor U4700 (N_4700,N_3559,N_3377);
xor U4701 (N_4701,N_3858,N_3517);
nor U4702 (N_4702,N_3749,N_3457);
nor U4703 (N_4703,N_3000,N_3755);
nand U4704 (N_4704,N_3784,N_3445);
or U4705 (N_4705,N_3244,N_3245);
nor U4706 (N_4706,N_3358,N_3655);
nand U4707 (N_4707,N_3110,N_3228);
nand U4708 (N_4708,N_3114,N_3047);
nor U4709 (N_4709,N_3541,N_3443);
or U4710 (N_4710,N_3812,N_3551);
nand U4711 (N_4711,N_3608,N_3179);
or U4712 (N_4712,N_3736,N_3690);
nor U4713 (N_4713,N_3526,N_3338);
or U4714 (N_4714,N_3262,N_3330);
xor U4715 (N_4715,N_3512,N_3858);
nor U4716 (N_4716,N_3566,N_3345);
nor U4717 (N_4717,N_3346,N_3969);
nand U4718 (N_4718,N_3582,N_3089);
or U4719 (N_4719,N_3316,N_3578);
nand U4720 (N_4720,N_3991,N_3507);
nor U4721 (N_4721,N_3593,N_3389);
xor U4722 (N_4722,N_3520,N_3721);
and U4723 (N_4723,N_3035,N_3263);
nor U4724 (N_4724,N_3156,N_3840);
or U4725 (N_4725,N_3466,N_3270);
and U4726 (N_4726,N_3863,N_3153);
nor U4727 (N_4727,N_3972,N_3906);
and U4728 (N_4728,N_3378,N_3848);
and U4729 (N_4729,N_3533,N_3997);
or U4730 (N_4730,N_3430,N_3078);
nand U4731 (N_4731,N_3382,N_3163);
nand U4732 (N_4732,N_3162,N_3235);
and U4733 (N_4733,N_3512,N_3497);
nor U4734 (N_4734,N_3556,N_3866);
nor U4735 (N_4735,N_3332,N_3542);
nand U4736 (N_4736,N_3409,N_3643);
xnor U4737 (N_4737,N_3167,N_3517);
nand U4738 (N_4738,N_3759,N_3653);
nor U4739 (N_4739,N_3842,N_3651);
and U4740 (N_4740,N_3527,N_3182);
or U4741 (N_4741,N_3995,N_3140);
or U4742 (N_4742,N_3698,N_3429);
or U4743 (N_4743,N_3622,N_3327);
nor U4744 (N_4744,N_3333,N_3618);
and U4745 (N_4745,N_3271,N_3411);
and U4746 (N_4746,N_3586,N_3726);
or U4747 (N_4747,N_3569,N_3842);
nand U4748 (N_4748,N_3665,N_3674);
nand U4749 (N_4749,N_3428,N_3489);
or U4750 (N_4750,N_3612,N_3720);
nor U4751 (N_4751,N_3993,N_3701);
nor U4752 (N_4752,N_3277,N_3623);
xor U4753 (N_4753,N_3764,N_3806);
nand U4754 (N_4754,N_3462,N_3719);
or U4755 (N_4755,N_3126,N_3921);
and U4756 (N_4756,N_3189,N_3332);
nand U4757 (N_4757,N_3432,N_3852);
nand U4758 (N_4758,N_3825,N_3176);
nor U4759 (N_4759,N_3792,N_3471);
nand U4760 (N_4760,N_3962,N_3069);
nor U4761 (N_4761,N_3530,N_3338);
or U4762 (N_4762,N_3557,N_3944);
or U4763 (N_4763,N_3438,N_3142);
and U4764 (N_4764,N_3673,N_3309);
and U4765 (N_4765,N_3736,N_3656);
and U4766 (N_4766,N_3603,N_3713);
or U4767 (N_4767,N_3841,N_3535);
and U4768 (N_4768,N_3412,N_3086);
nor U4769 (N_4769,N_3715,N_3655);
nand U4770 (N_4770,N_3805,N_3959);
xor U4771 (N_4771,N_3735,N_3269);
xor U4772 (N_4772,N_3867,N_3586);
and U4773 (N_4773,N_3282,N_3669);
and U4774 (N_4774,N_3114,N_3429);
nand U4775 (N_4775,N_3097,N_3345);
or U4776 (N_4776,N_3002,N_3033);
nand U4777 (N_4777,N_3276,N_3173);
and U4778 (N_4778,N_3715,N_3690);
and U4779 (N_4779,N_3811,N_3566);
or U4780 (N_4780,N_3013,N_3020);
nor U4781 (N_4781,N_3794,N_3591);
xnor U4782 (N_4782,N_3292,N_3442);
or U4783 (N_4783,N_3381,N_3331);
and U4784 (N_4784,N_3485,N_3166);
and U4785 (N_4785,N_3189,N_3532);
nor U4786 (N_4786,N_3775,N_3252);
nand U4787 (N_4787,N_3576,N_3650);
nand U4788 (N_4788,N_3425,N_3234);
and U4789 (N_4789,N_3304,N_3433);
or U4790 (N_4790,N_3245,N_3201);
nand U4791 (N_4791,N_3558,N_3769);
nor U4792 (N_4792,N_3661,N_3476);
nand U4793 (N_4793,N_3546,N_3443);
and U4794 (N_4794,N_3100,N_3025);
nor U4795 (N_4795,N_3080,N_3584);
or U4796 (N_4796,N_3850,N_3299);
nand U4797 (N_4797,N_3217,N_3731);
or U4798 (N_4798,N_3447,N_3607);
or U4799 (N_4799,N_3823,N_3605);
and U4800 (N_4800,N_3401,N_3828);
nand U4801 (N_4801,N_3008,N_3785);
nor U4802 (N_4802,N_3876,N_3680);
nand U4803 (N_4803,N_3061,N_3314);
and U4804 (N_4804,N_3309,N_3544);
and U4805 (N_4805,N_3639,N_3252);
and U4806 (N_4806,N_3440,N_3499);
nand U4807 (N_4807,N_3437,N_3112);
nor U4808 (N_4808,N_3398,N_3762);
and U4809 (N_4809,N_3037,N_3094);
nand U4810 (N_4810,N_3241,N_3626);
nor U4811 (N_4811,N_3147,N_3723);
and U4812 (N_4812,N_3687,N_3239);
and U4813 (N_4813,N_3551,N_3257);
nor U4814 (N_4814,N_3005,N_3711);
or U4815 (N_4815,N_3962,N_3275);
nor U4816 (N_4816,N_3994,N_3882);
and U4817 (N_4817,N_3958,N_3354);
and U4818 (N_4818,N_3821,N_3650);
or U4819 (N_4819,N_3217,N_3975);
nand U4820 (N_4820,N_3928,N_3895);
xnor U4821 (N_4821,N_3836,N_3938);
or U4822 (N_4822,N_3349,N_3751);
nor U4823 (N_4823,N_3554,N_3364);
and U4824 (N_4824,N_3182,N_3456);
xnor U4825 (N_4825,N_3488,N_3654);
and U4826 (N_4826,N_3502,N_3054);
nand U4827 (N_4827,N_3595,N_3540);
nand U4828 (N_4828,N_3488,N_3785);
nand U4829 (N_4829,N_3858,N_3330);
xnor U4830 (N_4830,N_3473,N_3068);
nor U4831 (N_4831,N_3248,N_3127);
and U4832 (N_4832,N_3044,N_3849);
nor U4833 (N_4833,N_3777,N_3747);
and U4834 (N_4834,N_3651,N_3568);
nor U4835 (N_4835,N_3929,N_3261);
or U4836 (N_4836,N_3570,N_3298);
nand U4837 (N_4837,N_3933,N_3230);
nand U4838 (N_4838,N_3099,N_3141);
and U4839 (N_4839,N_3956,N_3793);
xor U4840 (N_4840,N_3202,N_3285);
nand U4841 (N_4841,N_3902,N_3226);
and U4842 (N_4842,N_3973,N_3408);
xnor U4843 (N_4843,N_3539,N_3027);
nand U4844 (N_4844,N_3850,N_3328);
nor U4845 (N_4845,N_3093,N_3526);
xnor U4846 (N_4846,N_3924,N_3492);
or U4847 (N_4847,N_3879,N_3188);
nor U4848 (N_4848,N_3984,N_3311);
xnor U4849 (N_4849,N_3922,N_3142);
or U4850 (N_4850,N_3303,N_3188);
nand U4851 (N_4851,N_3505,N_3493);
or U4852 (N_4852,N_3381,N_3445);
nand U4853 (N_4853,N_3328,N_3701);
nand U4854 (N_4854,N_3894,N_3596);
and U4855 (N_4855,N_3800,N_3297);
or U4856 (N_4856,N_3435,N_3988);
or U4857 (N_4857,N_3539,N_3370);
or U4858 (N_4858,N_3071,N_3418);
nor U4859 (N_4859,N_3587,N_3012);
nand U4860 (N_4860,N_3549,N_3036);
or U4861 (N_4861,N_3906,N_3375);
nor U4862 (N_4862,N_3909,N_3333);
or U4863 (N_4863,N_3301,N_3034);
and U4864 (N_4864,N_3797,N_3963);
nor U4865 (N_4865,N_3202,N_3831);
or U4866 (N_4866,N_3775,N_3379);
xor U4867 (N_4867,N_3790,N_3896);
and U4868 (N_4868,N_3243,N_3114);
and U4869 (N_4869,N_3938,N_3683);
nor U4870 (N_4870,N_3074,N_3466);
or U4871 (N_4871,N_3755,N_3819);
and U4872 (N_4872,N_3014,N_3034);
nand U4873 (N_4873,N_3004,N_3968);
and U4874 (N_4874,N_3048,N_3514);
or U4875 (N_4875,N_3050,N_3568);
and U4876 (N_4876,N_3318,N_3464);
and U4877 (N_4877,N_3677,N_3595);
and U4878 (N_4878,N_3214,N_3241);
nor U4879 (N_4879,N_3635,N_3159);
and U4880 (N_4880,N_3532,N_3362);
or U4881 (N_4881,N_3659,N_3799);
or U4882 (N_4882,N_3422,N_3121);
and U4883 (N_4883,N_3155,N_3256);
nand U4884 (N_4884,N_3114,N_3712);
nand U4885 (N_4885,N_3593,N_3764);
nand U4886 (N_4886,N_3689,N_3171);
nor U4887 (N_4887,N_3252,N_3845);
nor U4888 (N_4888,N_3940,N_3910);
or U4889 (N_4889,N_3609,N_3793);
xor U4890 (N_4890,N_3154,N_3834);
nand U4891 (N_4891,N_3302,N_3390);
and U4892 (N_4892,N_3977,N_3994);
nand U4893 (N_4893,N_3829,N_3029);
or U4894 (N_4894,N_3115,N_3142);
nand U4895 (N_4895,N_3844,N_3098);
xor U4896 (N_4896,N_3604,N_3760);
nand U4897 (N_4897,N_3717,N_3512);
nor U4898 (N_4898,N_3467,N_3229);
and U4899 (N_4899,N_3731,N_3350);
and U4900 (N_4900,N_3836,N_3623);
and U4901 (N_4901,N_3859,N_3612);
xnor U4902 (N_4902,N_3961,N_3881);
xor U4903 (N_4903,N_3416,N_3545);
nor U4904 (N_4904,N_3747,N_3690);
or U4905 (N_4905,N_3876,N_3063);
nand U4906 (N_4906,N_3284,N_3381);
or U4907 (N_4907,N_3040,N_3185);
nand U4908 (N_4908,N_3590,N_3411);
nand U4909 (N_4909,N_3655,N_3338);
nand U4910 (N_4910,N_3171,N_3703);
xor U4911 (N_4911,N_3989,N_3581);
nor U4912 (N_4912,N_3257,N_3532);
and U4913 (N_4913,N_3462,N_3952);
or U4914 (N_4914,N_3606,N_3847);
nor U4915 (N_4915,N_3629,N_3130);
nand U4916 (N_4916,N_3430,N_3988);
nand U4917 (N_4917,N_3337,N_3383);
nand U4918 (N_4918,N_3603,N_3317);
and U4919 (N_4919,N_3920,N_3172);
nor U4920 (N_4920,N_3485,N_3834);
nor U4921 (N_4921,N_3863,N_3169);
nand U4922 (N_4922,N_3493,N_3117);
or U4923 (N_4923,N_3609,N_3119);
or U4924 (N_4924,N_3501,N_3517);
nand U4925 (N_4925,N_3717,N_3628);
nand U4926 (N_4926,N_3104,N_3975);
nor U4927 (N_4927,N_3049,N_3274);
nand U4928 (N_4928,N_3016,N_3928);
nand U4929 (N_4929,N_3199,N_3465);
and U4930 (N_4930,N_3688,N_3137);
nand U4931 (N_4931,N_3404,N_3212);
and U4932 (N_4932,N_3042,N_3307);
nor U4933 (N_4933,N_3307,N_3957);
or U4934 (N_4934,N_3559,N_3832);
nand U4935 (N_4935,N_3785,N_3344);
or U4936 (N_4936,N_3250,N_3679);
nand U4937 (N_4937,N_3709,N_3209);
nand U4938 (N_4938,N_3990,N_3665);
or U4939 (N_4939,N_3650,N_3168);
and U4940 (N_4940,N_3073,N_3854);
and U4941 (N_4941,N_3478,N_3497);
nand U4942 (N_4942,N_3364,N_3369);
nand U4943 (N_4943,N_3691,N_3999);
or U4944 (N_4944,N_3122,N_3124);
and U4945 (N_4945,N_3633,N_3418);
xnor U4946 (N_4946,N_3427,N_3167);
and U4947 (N_4947,N_3015,N_3585);
nor U4948 (N_4948,N_3960,N_3222);
nand U4949 (N_4949,N_3673,N_3687);
nand U4950 (N_4950,N_3572,N_3212);
and U4951 (N_4951,N_3596,N_3849);
xnor U4952 (N_4952,N_3832,N_3287);
nand U4953 (N_4953,N_3073,N_3114);
xor U4954 (N_4954,N_3870,N_3532);
or U4955 (N_4955,N_3046,N_3215);
nor U4956 (N_4956,N_3348,N_3636);
nand U4957 (N_4957,N_3598,N_3200);
and U4958 (N_4958,N_3790,N_3158);
or U4959 (N_4959,N_3408,N_3336);
xor U4960 (N_4960,N_3876,N_3148);
and U4961 (N_4961,N_3953,N_3289);
or U4962 (N_4962,N_3923,N_3727);
and U4963 (N_4963,N_3197,N_3519);
xnor U4964 (N_4964,N_3127,N_3998);
nand U4965 (N_4965,N_3357,N_3709);
nand U4966 (N_4966,N_3635,N_3083);
and U4967 (N_4967,N_3436,N_3885);
and U4968 (N_4968,N_3485,N_3799);
and U4969 (N_4969,N_3289,N_3131);
nand U4970 (N_4970,N_3358,N_3686);
nor U4971 (N_4971,N_3561,N_3076);
nand U4972 (N_4972,N_3019,N_3652);
or U4973 (N_4973,N_3967,N_3653);
nor U4974 (N_4974,N_3577,N_3999);
and U4975 (N_4975,N_3305,N_3269);
nor U4976 (N_4976,N_3440,N_3244);
xnor U4977 (N_4977,N_3303,N_3862);
or U4978 (N_4978,N_3338,N_3968);
nand U4979 (N_4979,N_3979,N_3227);
and U4980 (N_4980,N_3161,N_3334);
nand U4981 (N_4981,N_3277,N_3461);
and U4982 (N_4982,N_3851,N_3241);
nand U4983 (N_4983,N_3851,N_3704);
and U4984 (N_4984,N_3618,N_3123);
xor U4985 (N_4985,N_3206,N_3419);
and U4986 (N_4986,N_3564,N_3072);
and U4987 (N_4987,N_3382,N_3554);
nor U4988 (N_4988,N_3895,N_3483);
xnor U4989 (N_4989,N_3465,N_3494);
or U4990 (N_4990,N_3663,N_3397);
or U4991 (N_4991,N_3833,N_3199);
and U4992 (N_4992,N_3358,N_3337);
nand U4993 (N_4993,N_3965,N_3692);
nor U4994 (N_4994,N_3062,N_3300);
or U4995 (N_4995,N_3042,N_3735);
nand U4996 (N_4996,N_3204,N_3896);
and U4997 (N_4997,N_3046,N_3090);
or U4998 (N_4998,N_3681,N_3680);
and U4999 (N_4999,N_3500,N_3377);
or U5000 (N_5000,N_4030,N_4600);
nand U5001 (N_5001,N_4159,N_4811);
nand U5002 (N_5002,N_4217,N_4139);
or U5003 (N_5003,N_4950,N_4177);
nand U5004 (N_5004,N_4121,N_4781);
nor U5005 (N_5005,N_4793,N_4658);
nand U5006 (N_5006,N_4888,N_4898);
nor U5007 (N_5007,N_4709,N_4956);
xor U5008 (N_5008,N_4722,N_4918);
nand U5009 (N_5009,N_4308,N_4355);
nor U5010 (N_5010,N_4088,N_4059);
nand U5011 (N_5011,N_4093,N_4549);
nor U5012 (N_5012,N_4429,N_4981);
or U5013 (N_5013,N_4452,N_4362);
or U5014 (N_5014,N_4017,N_4304);
or U5015 (N_5015,N_4851,N_4441);
xor U5016 (N_5016,N_4557,N_4739);
and U5017 (N_5017,N_4468,N_4850);
and U5018 (N_5018,N_4735,N_4420);
nor U5019 (N_5019,N_4791,N_4741);
and U5020 (N_5020,N_4821,N_4909);
and U5021 (N_5021,N_4712,N_4652);
nor U5022 (N_5022,N_4412,N_4290);
nor U5023 (N_5023,N_4203,N_4630);
or U5024 (N_5024,N_4332,N_4757);
or U5025 (N_5025,N_4288,N_4531);
and U5026 (N_5026,N_4021,N_4767);
nor U5027 (N_5027,N_4760,N_4554);
nand U5028 (N_5028,N_4654,N_4014);
xnor U5029 (N_5029,N_4635,N_4284);
or U5030 (N_5030,N_4189,N_4108);
and U5031 (N_5031,N_4195,N_4970);
and U5032 (N_5032,N_4053,N_4939);
nor U5033 (N_5033,N_4125,N_4185);
nor U5034 (N_5034,N_4136,N_4987);
nand U5035 (N_5035,N_4782,N_4624);
and U5036 (N_5036,N_4442,N_4762);
nand U5037 (N_5037,N_4227,N_4055);
xor U5038 (N_5038,N_4102,N_4162);
nand U5039 (N_5039,N_4228,N_4020);
or U5040 (N_5040,N_4771,N_4696);
or U5041 (N_5041,N_4621,N_4153);
nand U5042 (N_5042,N_4346,N_4356);
and U5043 (N_5043,N_4359,N_4996);
nor U5044 (N_5044,N_4375,N_4345);
xor U5045 (N_5045,N_4384,N_4144);
nor U5046 (N_5046,N_4025,N_4516);
nor U5047 (N_5047,N_4647,N_4487);
or U5048 (N_5048,N_4740,N_4302);
or U5049 (N_5049,N_4210,N_4457);
nand U5050 (N_5050,N_4484,N_4891);
and U5051 (N_5051,N_4296,N_4838);
or U5052 (N_5052,N_4444,N_4150);
nor U5053 (N_5053,N_4197,N_4648);
nor U5054 (N_5054,N_4006,N_4922);
and U5055 (N_5055,N_4685,N_4618);
nor U5056 (N_5056,N_4009,N_4213);
or U5057 (N_5057,N_4573,N_4024);
nand U5058 (N_5058,N_4804,N_4868);
nand U5059 (N_5059,N_4410,N_4510);
and U5060 (N_5060,N_4016,N_4726);
and U5061 (N_5061,N_4677,N_4815);
xnor U5062 (N_5062,N_4928,N_4727);
or U5063 (N_5063,N_4094,N_4933);
and U5064 (N_5064,N_4836,N_4411);
nor U5065 (N_5065,N_4839,N_4226);
xnor U5066 (N_5066,N_4188,N_4958);
or U5067 (N_5067,N_4687,N_4978);
or U5068 (N_5068,N_4695,N_4103);
xnor U5069 (N_5069,N_4215,N_4772);
or U5070 (N_5070,N_4309,N_4329);
nand U5071 (N_5071,N_4235,N_4071);
or U5072 (N_5072,N_4634,N_4625);
xor U5073 (N_5073,N_4550,N_4074);
and U5074 (N_5074,N_4107,N_4907);
nor U5075 (N_5075,N_4609,N_4947);
and U5076 (N_5076,N_4028,N_4272);
xnor U5077 (N_5077,N_4565,N_4408);
nand U5078 (N_5078,N_4661,N_4248);
nor U5079 (N_5079,N_4916,N_4586);
or U5080 (N_5080,N_4334,N_4358);
or U5081 (N_5081,N_4876,N_4559);
nand U5082 (N_5082,N_4234,N_4867);
or U5083 (N_5083,N_4231,N_4099);
nor U5084 (N_5084,N_4287,N_4453);
xor U5085 (N_5085,N_4954,N_4090);
nand U5086 (N_5086,N_4966,N_4002);
nor U5087 (N_5087,N_4940,N_4505);
nand U5088 (N_5088,N_4973,N_4583);
xor U5089 (N_5089,N_4990,N_4493);
nor U5090 (N_5090,N_4529,N_4478);
nand U5091 (N_5091,N_4087,N_4523);
and U5092 (N_5092,N_4524,N_4174);
and U5093 (N_5093,N_4357,N_4617);
xor U5094 (N_5094,N_4083,N_4567);
nand U5095 (N_5095,N_4509,N_4657);
nor U5096 (N_5096,N_4596,N_4639);
and U5097 (N_5097,N_4388,N_4007);
nand U5098 (N_5098,N_4140,N_4642);
and U5099 (N_5099,N_4413,N_4906);
or U5100 (N_5100,N_4196,N_4001);
or U5101 (N_5101,N_4310,N_4335);
xor U5102 (N_5102,N_4731,N_4377);
or U5103 (N_5103,N_4462,N_4467);
nand U5104 (N_5104,N_4387,N_4394);
nand U5105 (N_5105,N_4466,N_4829);
or U5106 (N_5106,N_4165,N_4116);
xnor U5107 (N_5107,N_4750,N_4305);
and U5108 (N_5108,N_4459,N_4717);
and U5109 (N_5109,N_4490,N_4344);
or U5110 (N_5110,N_4029,N_4528);
nand U5111 (N_5111,N_4438,N_4240);
or U5112 (N_5112,N_4989,N_4707);
nand U5113 (N_5113,N_4572,N_4015);
xor U5114 (N_5114,N_4551,N_4570);
nand U5115 (N_5115,N_4184,N_4322);
nand U5116 (N_5116,N_4400,N_4084);
nand U5117 (N_5117,N_4667,N_4105);
nor U5118 (N_5118,N_4142,N_4341);
nand U5119 (N_5119,N_4371,N_4668);
nand U5120 (N_5120,N_4186,N_4921);
nor U5121 (N_5121,N_4859,N_4834);
or U5122 (N_5122,N_4544,N_4436);
or U5123 (N_5123,N_4167,N_4378);
nor U5124 (N_5124,N_4000,N_4830);
nor U5125 (N_5125,N_4948,N_4742);
and U5126 (N_5126,N_4983,N_4326);
or U5127 (N_5127,N_4828,N_4392);
nor U5128 (N_5128,N_4706,N_4034);
and U5129 (N_5129,N_4564,N_4884);
nor U5130 (N_5130,N_4708,N_4753);
nand U5131 (N_5131,N_4610,N_4222);
nor U5132 (N_5132,N_4044,N_4606);
or U5133 (N_5133,N_4808,N_4124);
or U5134 (N_5134,N_4612,N_4117);
and U5135 (N_5135,N_4148,N_4748);
nand U5136 (N_5136,N_4638,N_4699);
and U5137 (N_5137,N_4417,N_4869);
and U5138 (N_5138,N_4764,N_4569);
and U5139 (N_5139,N_4402,N_4279);
and U5140 (N_5140,N_4979,N_4337);
nand U5141 (N_5141,N_4004,N_4775);
xor U5142 (N_5142,N_4477,N_4019);
and U5143 (N_5143,N_4448,N_4703);
nand U5144 (N_5144,N_4443,N_4236);
and U5145 (N_5145,N_4343,N_4541);
or U5146 (N_5146,N_4128,N_4119);
nand U5147 (N_5147,N_4521,N_4373);
or U5148 (N_5148,N_4354,N_4818);
and U5149 (N_5149,N_4342,N_4246);
nand U5150 (N_5150,N_4458,N_4774);
nor U5151 (N_5151,N_4120,N_4666);
xnor U5152 (N_5152,N_4580,N_4198);
xnor U5153 (N_5153,N_4252,N_4568);
or U5154 (N_5154,N_4470,N_4330);
or U5155 (N_5155,N_4890,N_4450);
nor U5156 (N_5156,N_4698,N_4540);
and U5157 (N_5157,N_4785,N_4249);
or U5158 (N_5158,N_4321,N_4046);
nor U5159 (N_5159,N_4315,N_4212);
and U5160 (N_5160,N_4241,N_4435);
or U5161 (N_5161,N_4942,N_4447);
and U5162 (N_5162,N_4705,N_4905);
nor U5163 (N_5163,N_4862,N_4786);
nor U5164 (N_5164,N_4861,N_4843);
or U5165 (N_5165,N_4230,N_4715);
or U5166 (N_5166,N_4012,N_4840);
nand U5167 (N_5167,N_4880,N_4061);
nor U5168 (N_5168,N_4433,N_4999);
xor U5169 (N_5169,N_4454,N_4746);
or U5170 (N_5170,N_4298,N_4456);
or U5171 (N_5171,N_4533,N_4381);
and U5172 (N_5172,N_4043,N_4488);
or U5173 (N_5173,N_4945,N_4239);
and U5174 (N_5174,N_4670,N_4190);
nor U5175 (N_5175,N_4010,N_4406);
and U5176 (N_5176,N_4277,N_4409);
nand U5177 (N_5177,N_4424,N_4496);
and U5178 (N_5178,N_4995,N_4532);
nand U5179 (N_5179,N_4694,N_4702);
nor U5180 (N_5180,N_4134,N_4504);
or U5181 (N_5181,N_4201,N_4263);
and U5182 (N_5182,N_4419,N_4736);
or U5183 (N_5183,N_4486,N_4372);
and U5184 (N_5184,N_4320,N_4721);
or U5185 (N_5185,N_4115,N_4562);
or U5186 (N_5186,N_4187,N_4011);
and U5187 (N_5187,N_4156,N_4066);
or U5188 (N_5188,N_4449,N_4849);
xor U5189 (N_5189,N_4316,N_4713);
or U5190 (N_5190,N_4794,N_4542);
xor U5191 (N_5191,N_4604,N_4650);
and U5192 (N_5192,N_4615,N_4181);
or U5193 (N_5193,N_4340,N_4306);
or U5194 (N_5194,N_4660,N_4328);
nand U5195 (N_5195,N_4951,N_4395);
nand U5196 (N_5196,N_4414,N_4092);
and U5197 (N_5197,N_4991,N_4883);
nand U5198 (N_5198,N_4558,N_4506);
and U5199 (N_5199,N_4260,N_4935);
or U5200 (N_5200,N_4502,N_4060);
and U5201 (N_5201,N_4595,N_4132);
xor U5202 (N_5202,N_4976,N_4338);
and U5203 (N_5203,N_4282,N_4137);
nor U5204 (N_5204,N_4543,N_4678);
and U5205 (N_5205,N_4111,N_4257);
nor U5206 (N_5206,N_4026,N_4555);
xnor U5207 (N_5207,N_4104,N_4644);
xnor U5208 (N_5208,N_4113,N_4180);
nand U5209 (N_5209,N_4971,N_4538);
nand U5210 (N_5210,N_4582,N_4048);
and U5211 (N_5211,N_4545,N_4503);
nand U5212 (N_5212,N_4789,N_4194);
nor U5213 (N_5213,N_4518,N_4056);
and U5214 (N_5214,N_4245,N_4261);
nor U5215 (N_5215,N_4319,N_4936);
nand U5216 (N_5216,N_4199,N_4603);
nand U5217 (N_5217,N_4672,N_4626);
nor U5218 (N_5218,N_4934,N_4091);
and U5219 (N_5219,N_4943,N_4908);
or U5220 (N_5220,N_4318,N_4745);
and U5221 (N_5221,N_4258,N_4178);
nand U5222 (N_5222,N_4498,N_4856);
and U5223 (N_5223,N_4637,N_4941);
or U5224 (N_5224,N_4988,N_4895);
nor U5225 (N_5225,N_4439,N_4919);
xnor U5226 (N_5226,N_4396,N_4292);
and U5227 (N_5227,N_4313,N_4293);
and U5228 (N_5228,N_4407,N_4275);
or U5229 (N_5229,N_4110,N_4535);
and U5230 (N_5230,N_4323,N_4253);
nor U5231 (N_5231,N_4405,N_4689);
nand U5232 (N_5232,N_4118,N_4163);
and U5233 (N_5233,N_4866,N_4464);
xor U5234 (N_5234,N_4931,N_4566);
and U5235 (N_5235,N_4857,N_4809);
nand U5236 (N_5236,N_4910,N_4640);
nor U5237 (N_5237,N_4806,N_4593);
xnor U5238 (N_5238,N_4955,N_4653);
or U5239 (N_5239,N_4679,N_4147);
nor U5240 (N_5240,N_4237,N_4812);
or U5241 (N_5241,N_4845,N_4875);
nor U5242 (N_5242,N_4386,N_4175);
nor U5243 (N_5243,N_4776,N_4686);
nand U5244 (N_5244,N_4281,N_4810);
nand U5245 (N_5245,N_4796,N_4473);
and U5246 (N_5246,N_4063,N_4601);
or U5247 (N_5247,N_4805,N_4751);
nand U5248 (N_5248,N_4984,N_4511);
xor U5249 (N_5249,N_4100,N_4530);
nand U5250 (N_5250,N_4271,N_4097);
or U5251 (N_5251,N_4923,N_4968);
nand U5252 (N_5252,N_4613,N_4065);
or U5253 (N_5253,N_4446,N_4204);
nor U5254 (N_5254,N_4311,N_4733);
nor U5255 (N_5255,N_4902,N_4171);
nor U5256 (N_5256,N_4598,N_4367);
nor U5257 (N_5257,N_4636,N_4998);
nand U5258 (N_5258,N_4391,N_4837);
nor U5259 (N_5259,N_4611,N_4041);
nor U5260 (N_5260,N_4799,N_4588);
or U5261 (N_5261,N_4130,N_4858);
nor U5262 (N_5262,N_4526,N_4070);
nand U5263 (N_5263,N_4690,N_4508);
xor U5264 (N_5264,N_4813,N_4949);
or U5265 (N_5265,N_4169,N_4114);
nand U5266 (N_5266,N_4769,N_4929);
and U5267 (N_5267,N_4759,N_4040);
nor U5268 (N_5268,N_4633,N_4584);
nand U5269 (N_5269,N_4164,N_4952);
nor U5270 (N_5270,N_4824,N_4669);
nor U5271 (N_5271,N_4525,N_4427);
or U5272 (N_5272,N_4183,N_4897);
nor U5273 (N_5273,N_4623,N_4832);
nor U5274 (N_5274,N_4539,N_4045);
and U5275 (N_5275,N_4202,N_4497);
or U5276 (N_5276,N_4106,N_4461);
or U5277 (N_5277,N_4283,N_4182);
nor U5278 (N_5278,N_4961,N_4138);
nor U5279 (N_5279,N_4676,N_4432);
nand U5280 (N_5280,N_4629,N_4244);
and U5281 (N_5281,N_4513,N_4295);
nor U5282 (N_5282,N_4064,N_4398);
nand U5283 (N_5283,N_4471,N_4882);
and U5284 (N_5284,N_4141,N_4176);
nor U5285 (N_5285,N_4369,N_4822);
or U5286 (N_5286,N_4957,N_4853);
nor U5287 (N_5287,N_4756,N_4874);
nor U5288 (N_5288,N_4982,N_4294);
nor U5289 (N_5289,N_4482,N_4997);
nor U5290 (N_5290,N_4963,N_4206);
nand U5291 (N_5291,N_4380,N_4109);
nand U5292 (N_5292,N_4224,N_4548);
nand U5293 (N_5293,N_4552,N_4327);
or U5294 (N_5294,N_4974,N_4145);
nor U5295 (N_5295,N_4052,N_4827);
nand U5296 (N_5296,N_4023,N_4719);
and U5297 (N_5297,N_4209,N_4254);
nor U5298 (N_5298,N_4546,N_4415);
nor U5299 (N_5299,N_4331,N_4553);
nor U5300 (N_5300,N_4985,N_4273);
xor U5301 (N_5301,N_4428,N_4072);
nand U5302 (N_5302,N_4434,N_4501);
nor U5303 (N_5303,N_4483,N_4317);
and U5304 (N_5304,N_4057,N_4291);
and U5305 (N_5305,N_4758,N_4925);
and U5306 (N_5306,N_4080,N_4537);
and U5307 (N_5307,N_4692,N_4013);
or U5308 (N_5308,N_4737,N_4770);
and U5309 (N_5309,N_4363,N_4219);
nor U5310 (N_5310,N_4852,N_4437);
xor U5311 (N_5311,N_4659,N_4270);
nand U5312 (N_5312,N_4911,N_4238);
nand U5313 (N_5313,N_4930,N_4903);
xnor U5314 (N_5314,N_4481,N_4077);
nor U5315 (N_5315,N_4734,N_4465);
nor U5316 (N_5316,N_4243,N_4826);
nand U5317 (N_5317,N_4460,N_4364);
nor U5318 (N_5318,N_4079,N_4616);
and U5319 (N_5319,N_4297,N_4605);
nor U5320 (N_5320,N_4844,N_4247);
or U5321 (N_5321,N_4135,N_4720);
nor U5322 (N_5322,N_4783,N_4920);
or U5323 (N_5323,N_4499,N_4347);
nand U5324 (N_5324,N_4743,N_4211);
or U5325 (N_5325,N_4519,N_4896);
and U5326 (N_5326,N_4455,N_4860);
nor U5327 (N_5327,N_4887,N_4744);
nand U5328 (N_5328,N_4390,N_4370);
and U5329 (N_5329,N_4879,N_4797);
and U5330 (N_5330,N_4807,N_4366);
nand U5331 (N_5331,N_4299,N_4058);
or U5332 (N_5332,N_4475,N_4480);
nand U5333 (N_5333,N_4067,N_4368);
nor U5334 (N_5334,N_4870,N_4872);
nand U5335 (N_5335,N_4160,N_4581);
nor U5336 (N_5336,N_4445,N_4663);
nand U5337 (N_5337,N_4577,N_4068);
or U5338 (N_5338,N_4846,N_4675);
and U5339 (N_5339,N_4491,N_4969);
nor U5340 (N_5340,N_4301,N_4223);
nor U5341 (N_5341,N_4571,N_4289);
nor U5342 (N_5342,N_4730,N_4205);
or U5343 (N_5343,N_4589,N_4801);
nand U5344 (N_5344,N_4885,N_4915);
and U5345 (N_5345,N_4819,N_4312);
nand U5346 (N_5346,N_4085,N_4101);
xnor U5347 (N_5347,N_4563,N_4324);
nor U5348 (N_5348,N_4076,N_4665);
nand U5349 (N_5349,N_4701,N_4697);
and U5350 (N_5350,N_4149,N_4723);
nor U5351 (N_5351,N_4032,N_4965);
xnor U5352 (N_5352,N_4765,N_4575);
nor U5353 (N_5353,N_4401,N_4641);
nor U5354 (N_5354,N_4865,N_4353);
nand U5355 (N_5355,N_4778,N_4716);
or U5356 (N_5356,N_4833,N_4802);
nand U5357 (N_5357,N_4592,N_4926);
nand U5358 (N_5358,N_4168,N_4440);
nand U5359 (N_5359,N_4711,N_4123);
nand U5360 (N_5360,N_4924,N_4161);
and U5361 (N_5361,N_4912,N_4674);
nand U5362 (N_5362,N_4574,N_4607);
or U5363 (N_5363,N_4560,N_4738);
nand U5364 (N_5364,N_4389,N_4536);
and U5365 (N_5365,N_4766,N_4075);
and U5366 (N_5366,N_4547,N_4307);
nor U5367 (N_5367,N_4155,N_4749);
xor U5368 (N_5368,N_4350,N_4179);
or U5369 (N_5369,N_4649,N_4430);
or U5370 (N_5370,N_4233,N_4399);
and U5371 (N_5371,N_4422,N_4031);
and U5372 (N_5372,N_4208,N_4688);
nor U5373 (N_5373,N_4431,N_4779);
and U5374 (N_5374,N_4993,N_4474);
nor U5375 (N_5375,N_4873,N_4494);
nor U5376 (N_5376,N_4514,N_4938);
nor U5377 (N_5377,N_4225,N_4143);
nor U5378 (N_5378,N_4193,N_4964);
nor U5379 (N_5379,N_4421,N_4325);
nand U5380 (N_5380,N_4214,N_4038);
nor U5381 (N_5381,N_4269,N_4251);
and U5382 (N_5382,N_4780,N_4614);
nand U5383 (N_5383,N_4095,N_4655);
nor U5384 (N_5384,N_4881,N_4628);
nor U5385 (N_5385,N_4492,N_4098);
and U5386 (N_5386,N_4286,N_4729);
nand U5387 (N_5387,N_4714,N_4752);
xnor U5388 (N_5388,N_4820,N_4047);
and U5389 (N_5389,N_4517,N_4397);
nor U5390 (N_5390,N_4520,N_4792);
nor U5391 (N_5391,N_4036,N_4127);
nor U5392 (N_5392,N_4900,N_4027);
nand U5393 (N_5393,N_4280,N_4725);
or U5394 (N_5394,N_4814,N_4967);
and U5395 (N_5395,N_4587,N_4073);
nor U5396 (N_5396,N_4986,N_4773);
and U5397 (N_5397,N_4899,N_4220);
and U5398 (N_5398,N_4122,N_4927);
nor U5399 (N_5399,N_4361,N_4005);
and U5400 (N_5400,N_4864,N_4597);
xnor U5401 (N_5401,N_4485,N_4894);
nor U5402 (N_5402,N_4049,N_4917);
xor U5403 (N_5403,N_4817,N_4627);
and U5404 (N_5404,N_4823,N_4904);
nor U5405 (N_5405,N_4841,N_4728);
and U5406 (N_5406,N_4192,N_4994);
nand U5407 (N_5407,N_4037,N_4382);
xnor U5408 (N_5408,N_4704,N_4082);
and U5409 (N_5409,N_4336,N_4953);
xnor U5410 (N_5410,N_4622,N_4579);
nor U5411 (N_5411,N_4146,N_4191);
and U5412 (N_5412,N_4268,N_4877);
nand U5413 (N_5413,N_4602,N_4795);
nor U5414 (N_5414,N_4385,N_4365);
nand U5415 (N_5415,N_4300,N_4761);
nor U5416 (N_5416,N_4932,N_4096);
nand U5417 (N_5417,N_4255,N_4673);
nor U5418 (N_5418,N_4515,N_4416);
and U5419 (N_5419,N_4078,N_4278);
and U5420 (N_5420,N_4285,N_4418);
and U5421 (N_5421,N_4732,N_4423);
and U5422 (N_5422,N_4264,N_4207);
nor U5423 (N_5423,N_4878,N_4349);
and U5424 (N_5424,N_4348,N_4170);
xor U5425 (N_5425,N_4276,N_4383);
nand U5426 (N_5426,N_4803,N_4229);
and U5427 (N_5427,N_4018,N_4662);
nor U5428 (N_5428,N_4724,N_4379);
nor U5429 (N_5429,N_4784,N_4039);
nor U5430 (N_5430,N_4152,N_4946);
nor U5431 (N_5431,N_4035,N_4003);
nand U5432 (N_5432,N_4755,N_4050);
nor U5433 (N_5433,N_4608,N_4787);
and U5434 (N_5434,N_4022,N_4671);
or U5435 (N_5435,N_4218,N_4901);
xnor U5436 (N_5436,N_4835,N_4975);
or U5437 (N_5437,N_4576,N_4972);
and U5438 (N_5438,N_4374,N_4173);
or U5439 (N_5439,N_4871,N_4768);
or U5440 (N_5440,N_4578,N_4333);
and U5441 (N_5441,N_4266,N_4042);
nand U5442 (N_5442,N_4561,N_4556);
nand U5443 (N_5443,N_4632,N_4200);
xor U5444 (N_5444,N_4265,N_4274);
or U5445 (N_5445,N_4681,N_4500);
or U5446 (N_5446,N_4684,N_4351);
nand U5447 (N_5447,N_4527,N_4062);
nand U5448 (N_5448,N_4472,N_4133);
nor U5449 (N_5449,N_4594,N_4129);
and U5450 (N_5450,N_4451,N_4825);
and U5451 (N_5451,N_4403,N_4691);
nor U5452 (N_5452,N_4664,N_4816);
nor U5453 (N_5453,N_4360,N_4495);
and U5454 (N_5454,N_4081,N_4937);
and U5455 (N_5455,N_4683,N_4718);
nor U5456 (N_5456,N_4962,N_4256);
nand U5457 (N_5457,N_4259,N_4131);
nand U5458 (N_5458,N_4848,N_4680);
xor U5459 (N_5459,N_4710,N_4651);
nand U5460 (N_5460,N_4599,N_4790);
and U5461 (N_5461,N_4944,N_4631);
nor U5462 (N_5462,N_4393,N_4842);
nand U5463 (N_5463,N_4892,N_4886);
nor U5464 (N_5464,N_4585,N_4033);
and U5465 (N_5465,N_4619,N_4854);
and U5466 (N_5466,N_4158,N_4914);
nand U5467 (N_5467,N_4069,N_4847);
nor U5468 (N_5468,N_4250,N_4643);
and U5469 (N_5469,N_4425,N_4763);
or U5470 (N_5470,N_4855,N_4151);
nand U5471 (N_5471,N_4522,N_4051);
xor U5472 (N_5472,N_4893,N_4242);
and U5473 (N_5473,N_4216,N_4777);
xor U5474 (N_5474,N_4476,N_4267);
nor U5475 (N_5475,N_4960,N_4992);
nand U5476 (N_5476,N_4798,N_4889);
nand U5477 (N_5477,N_4863,N_4534);
or U5478 (N_5478,N_4656,N_4126);
or U5479 (N_5479,N_4054,N_4089);
nand U5480 (N_5480,N_4700,N_4221);
or U5481 (N_5481,N_4590,N_4507);
and U5482 (N_5482,N_4086,N_4172);
nand U5483 (N_5483,N_4166,N_4314);
nand U5484 (N_5484,N_4959,N_4112);
and U5485 (N_5485,N_4463,N_4980);
and U5486 (N_5486,N_4693,N_4232);
nand U5487 (N_5487,N_4512,N_4352);
nand U5488 (N_5488,N_4469,N_4913);
nand U5489 (N_5489,N_4404,N_4339);
or U5490 (N_5490,N_4788,N_4489);
and U5491 (N_5491,N_4157,N_4754);
or U5492 (N_5492,N_4479,N_4426);
or U5493 (N_5493,N_4303,N_4800);
xnor U5494 (N_5494,N_4831,N_4262);
nor U5495 (N_5495,N_4747,N_4646);
and U5496 (N_5496,N_4154,N_4645);
or U5497 (N_5497,N_4682,N_4591);
nor U5498 (N_5498,N_4376,N_4977);
nor U5499 (N_5499,N_4008,N_4620);
xor U5500 (N_5500,N_4991,N_4248);
or U5501 (N_5501,N_4363,N_4652);
nor U5502 (N_5502,N_4519,N_4684);
and U5503 (N_5503,N_4528,N_4179);
xor U5504 (N_5504,N_4415,N_4639);
nor U5505 (N_5505,N_4066,N_4822);
nor U5506 (N_5506,N_4243,N_4857);
and U5507 (N_5507,N_4277,N_4867);
nand U5508 (N_5508,N_4791,N_4473);
nor U5509 (N_5509,N_4147,N_4201);
nand U5510 (N_5510,N_4864,N_4613);
or U5511 (N_5511,N_4479,N_4444);
xor U5512 (N_5512,N_4538,N_4639);
or U5513 (N_5513,N_4956,N_4684);
nand U5514 (N_5514,N_4685,N_4353);
nor U5515 (N_5515,N_4598,N_4025);
xor U5516 (N_5516,N_4965,N_4885);
or U5517 (N_5517,N_4274,N_4526);
nor U5518 (N_5518,N_4199,N_4589);
nand U5519 (N_5519,N_4259,N_4330);
nand U5520 (N_5520,N_4726,N_4676);
nand U5521 (N_5521,N_4579,N_4356);
nor U5522 (N_5522,N_4510,N_4423);
nand U5523 (N_5523,N_4071,N_4795);
xnor U5524 (N_5524,N_4183,N_4235);
xor U5525 (N_5525,N_4762,N_4213);
and U5526 (N_5526,N_4436,N_4300);
or U5527 (N_5527,N_4924,N_4200);
or U5528 (N_5528,N_4774,N_4136);
nor U5529 (N_5529,N_4604,N_4902);
nand U5530 (N_5530,N_4858,N_4800);
and U5531 (N_5531,N_4739,N_4284);
nor U5532 (N_5532,N_4041,N_4321);
and U5533 (N_5533,N_4152,N_4747);
nor U5534 (N_5534,N_4723,N_4144);
nand U5535 (N_5535,N_4330,N_4185);
and U5536 (N_5536,N_4063,N_4586);
or U5537 (N_5537,N_4089,N_4596);
or U5538 (N_5538,N_4328,N_4498);
or U5539 (N_5539,N_4545,N_4244);
nand U5540 (N_5540,N_4776,N_4960);
and U5541 (N_5541,N_4644,N_4884);
nand U5542 (N_5542,N_4442,N_4637);
or U5543 (N_5543,N_4412,N_4721);
nor U5544 (N_5544,N_4755,N_4238);
or U5545 (N_5545,N_4014,N_4761);
or U5546 (N_5546,N_4359,N_4987);
nand U5547 (N_5547,N_4563,N_4430);
xor U5548 (N_5548,N_4327,N_4623);
xor U5549 (N_5549,N_4576,N_4267);
nand U5550 (N_5550,N_4437,N_4706);
nand U5551 (N_5551,N_4741,N_4892);
and U5552 (N_5552,N_4784,N_4196);
or U5553 (N_5553,N_4905,N_4072);
or U5554 (N_5554,N_4663,N_4507);
nand U5555 (N_5555,N_4031,N_4303);
and U5556 (N_5556,N_4882,N_4856);
and U5557 (N_5557,N_4092,N_4469);
or U5558 (N_5558,N_4239,N_4996);
nor U5559 (N_5559,N_4757,N_4728);
or U5560 (N_5560,N_4299,N_4286);
nand U5561 (N_5561,N_4395,N_4936);
and U5562 (N_5562,N_4118,N_4997);
and U5563 (N_5563,N_4838,N_4336);
or U5564 (N_5564,N_4882,N_4974);
and U5565 (N_5565,N_4709,N_4804);
or U5566 (N_5566,N_4417,N_4092);
or U5567 (N_5567,N_4642,N_4480);
nor U5568 (N_5568,N_4460,N_4977);
and U5569 (N_5569,N_4954,N_4844);
nor U5570 (N_5570,N_4784,N_4249);
nor U5571 (N_5571,N_4191,N_4854);
and U5572 (N_5572,N_4893,N_4913);
or U5573 (N_5573,N_4240,N_4314);
or U5574 (N_5574,N_4310,N_4133);
nor U5575 (N_5575,N_4411,N_4157);
nor U5576 (N_5576,N_4864,N_4433);
and U5577 (N_5577,N_4364,N_4233);
nand U5578 (N_5578,N_4067,N_4333);
nor U5579 (N_5579,N_4502,N_4904);
nand U5580 (N_5580,N_4581,N_4844);
nand U5581 (N_5581,N_4751,N_4151);
nand U5582 (N_5582,N_4915,N_4328);
and U5583 (N_5583,N_4811,N_4406);
or U5584 (N_5584,N_4641,N_4801);
nor U5585 (N_5585,N_4390,N_4188);
nand U5586 (N_5586,N_4197,N_4640);
or U5587 (N_5587,N_4386,N_4881);
and U5588 (N_5588,N_4251,N_4548);
or U5589 (N_5589,N_4721,N_4128);
nand U5590 (N_5590,N_4051,N_4535);
xnor U5591 (N_5591,N_4183,N_4812);
and U5592 (N_5592,N_4769,N_4196);
and U5593 (N_5593,N_4475,N_4489);
or U5594 (N_5594,N_4197,N_4339);
nor U5595 (N_5595,N_4167,N_4109);
nor U5596 (N_5596,N_4907,N_4363);
nor U5597 (N_5597,N_4586,N_4047);
nor U5598 (N_5598,N_4660,N_4073);
xnor U5599 (N_5599,N_4112,N_4663);
nor U5600 (N_5600,N_4613,N_4571);
and U5601 (N_5601,N_4485,N_4503);
or U5602 (N_5602,N_4289,N_4025);
nand U5603 (N_5603,N_4035,N_4525);
nor U5604 (N_5604,N_4838,N_4108);
and U5605 (N_5605,N_4667,N_4846);
and U5606 (N_5606,N_4941,N_4819);
and U5607 (N_5607,N_4169,N_4672);
xnor U5608 (N_5608,N_4917,N_4690);
or U5609 (N_5609,N_4268,N_4473);
and U5610 (N_5610,N_4403,N_4048);
or U5611 (N_5611,N_4515,N_4378);
xor U5612 (N_5612,N_4875,N_4242);
or U5613 (N_5613,N_4201,N_4905);
nor U5614 (N_5614,N_4608,N_4768);
nand U5615 (N_5615,N_4613,N_4377);
nor U5616 (N_5616,N_4592,N_4836);
or U5617 (N_5617,N_4809,N_4259);
xor U5618 (N_5618,N_4838,N_4224);
xnor U5619 (N_5619,N_4535,N_4028);
and U5620 (N_5620,N_4522,N_4270);
nor U5621 (N_5621,N_4576,N_4908);
xor U5622 (N_5622,N_4456,N_4259);
nand U5623 (N_5623,N_4876,N_4352);
and U5624 (N_5624,N_4014,N_4805);
xnor U5625 (N_5625,N_4887,N_4079);
nand U5626 (N_5626,N_4143,N_4078);
nor U5627 (N_5627,N_4862,N_4447);
nor U5628 (N_5628,N_4886,N_4594);
nor U5629 (N_5629,N_4748,N_4993);
nor U5630 (N_5630,N_4786,N_4763);
or U5631 (N_5631,N_4183,N_4914);
and U5632 (N_5632,N_4081,N_4861);
or U5633 (N_5633,N_4537,N_4210);
and U5634 (N_5634,N_4395,N_4269);
or U5635 (N_5635,N_4665,N_4332);
nor U5636 (N_5636,N_4981,N_4630);
nor U5637 (N_5637,N_4744,N_4659);
nand U5638 (N_5638,N_4952,N_4583);
or U5639 (N_5639,N_4727,N_4081);
nand U5640 (N_5640,N_4118,N_4814);
and U5641 (N_5641,N_4463,N_4190);
and U5642 (N_5642,N_4826,N_4645);
and U5643 (N_5643,N_4165,N_4583);
nand U5644 (N_5644,N_4922,N_4408);
and U5645 (N_5645,N_4487,N_4938);
xor U5646 (N_5646,N_4063,N_4937);
or U5647 (N_5647,N_4362,N_4297);
nor U5648 (N_5648,N_4845,N_4096);
nand U5649 (N_5649,N_4274,N_4759);
nand U5650 (N_5650,N_4615,N_4720);
and U5651 (N_5651,N_4251,N_4400);
and U5652 (N_5652,N_4271,N_4722);
xor U5653 (N_5653,N_4485,N_4111);
nor U5654 (N_5654,N_4870,N_4190);
nor U5655 (N_5655,N_4916,N_4876);
nand U5656 (N_5656,N_4794,N_4695);
and U5657 (N_5657,N_4293,N_4404);
nand U5658 (N_5658,N_4911,N_4531);
nor U5659 (N_5659,N_4711,N_4186);
nor U5660 (N_5660,N_4989,N_4086);
or U5661 (N_5661,N_4480,N_4583);
nor U5662 (N_5662,N_4216,N_4776);
nor U5663 (N_5663,N_4189,N_4525);
or U5664 (N_5664,N_4637,N_4500);
nor U5665 (N_5665,N_4513,N_4482);
nor U5666 (N_5666,N_4740,N_4942);
nor U5667 (N_5667,N_4737,N_4258);
nor U5668 (N_5668,N_4682,N_4057);
and U5669 (N_5669,N_4488,N_4935);
and U5670 (N_5670,N_4006,N_4645);
nor U5671 (N_5671,N_4335,N_4417);
and U5672 (N_5672,N_4869,N_4662);
or U5673 (N_5673,N_4271,N_4945);
nand U5674 (N_5674,N_4897,N_4534);
nor U5675 (N_5675,N_4176,N_4583);
and U5676 (N_5676,N_4410,N_4028);
or U5677 (N_5677,N_4059,N_4837);
nand U5678 (N_5678,N_4658,N_4324);
and U5679 (N_5679,N_4104,N_4684);
and U5680 (N_5680,N_4602,N_4763);
nand U5681 (N_5681,N_4133,N_4618);
or U5682 (N_5682,N_4889,N_4292);
or U5683 (N_5683,N_4335,N_4440);
or U5684 (N_5684,N_4712,N_4957);
and U5685 (N_5685,N_4363,N_4741);
or U5686 (N_5686,N_4408,N_4617);
or U5687 (N_5687,N_4291,N_4611);
or U5688 (N_5688,N_4987,N_4105);
nand U5689 (N_5689,N_4696,N_4154);
nand U5690 (N_5690,N_4728,N_4670);
nand U5691 (N_5691,N_4422,N_4911);
or U5692 (N_5692,N_4325,N_4804);
or U5693 (N_5693,N_4796,N_4205);
nand U5694 (N_5694,N_4320,N_4223);
nor U5695 (N_5695,N_4565,N_4777);
nor U5696 (N_5696,N_4134,N_4332);
nand U5697 (N_5697,N_4438,N_4645);
or U5698 (N_5698,N_4380,N_4850);
and U5699 (N_5699,N_4447,N_4060);
or U5700 (N_5700,N_4652,N_4950);
and U5701 (N_5701,N_4471,N_4555);
or U5702 (N_5702,N_4399,N_4986);
nor U5703 (N_5703,N_4986,N_4243);
xor U5704 (N_5704,N_4576,N_4061);
nor U5705 (N_5705,N_4156,N_4021);
or U5706 (N_5706,N_4549,N_4646);
nand U5707 (N_5707,N_4345,N_4645);
nand U5708 (N_5708,N_4257,N_4292);
xor U5709 (N_5709,N_4758,N_4619);
nand U5710 (N_5710,N_4228,N_4762);
or U5711 (N_5711,N_4644,N_4977);
nor U5712 (N_5712,N_4282,N_4425);
or U5713 (N_5713,N_4643,N_4418);
nor U5714 (N_5714,N_4263,N_4897);
and U5715 (N_5715,N_4591,N_4858);
xnor U5716 (N_5716,N_4715,N_4238);
or U5717 (N_5717,N_4225,N_4354);
nand U5718 (N_5718,N_4625,N_4277);
or U5719 (N_5719,N_4706,N_4772);
nor U5720 (N_5720,N_4702,N_4297);
or U5721 (N_5721,N_4311,N_4634);
nand U5722 (N_5722,N_4450,N_4555);
nand U5723 (N_5723,N_4726,N_4159);
nand U5724 (N_5724,N_4010,N_4613);
nor U5725 (N_5725,N_4584,N_4344);
and U5726 (N_5726,N_4383,N_4854);
nor U5727 (N_5727,N_4527,N_4679);
nand U5728 (N_5728,N_4878,N_4721);
nand U5729 (N_5729,N_4217,N_4463);
and U5730 (N_5730,N_4452,N_4465);
and U5731 (N_5731,N_4317,N_4052);
or U5732 (N_5732,N_4598,N_4062);
nor U5733 (N_5733,N_4992,N_4267);
nand U5734 (N_5734,N_4953,N_4962);
or U5735 (N_5735,N_4523,N_4928);
or U5736 (N_5736,N_4366,N_4233);
nor U5737 (N_5737,N_4415,N_4533);
xor U5738 (N_5738,N_4633,N_4873);
and U5739 (N_5739,N_4844,N_4904);
xnor U5740 (N_5740,N_4378,N_4740);
nand U5741 (N_5741,N_4263,N_4593);
nand U5742 (N_5742,N_4501,N_4858);
nand U5743 (N_5743,N_4076,N_4814);
and U5744 (N_5744,N_4035,N_4896);
or U5745 (N_5745,N_4706,N_4051);
or U5746 (N_5746,N_4839,N_4493);
xnor U5747 (N_5747,N_4266,N_4091);
or U5748 (N_5748,N_4163,N_4608);
nor U5749 (N_5749,N_4903,N_4736);
and U5750 (N_5750,N_4354,N_4032);
or U5751 (N_5751,N_4919,N_4006);
and U5752 (N_5752,N_4374,N_4716);
nor U5753 (N_5753,N_4751,N_4078);
and U5754 (N_5754,N_4325,N_4954);
nand U5755 (N_5755,N_4560,N_4325);
nor U5756 (N_5756,N_4695,N_4557);
xor U5757 (N_5757,N_4117,N_4075);
nor U5758 (N_5758,N_4454,N_4528);
nand U5759 (N_5759,N_4669,N_4673);
and U5760 (N_5760,N_4593,N_4163);
nor U5761 (N_5761,N_4029,N_4625);
or U5762 (N_5762,N_4949,N_4849);
and U5763 (N_5763,N_4940,N_4622);
and U5764 (N_5764,N_4412,N_4014);
nand U5765 (N_5765,N_4788,N_4225);
or U5766 (N_5766,N_4111,N_4532);
nand U5767 (N_5767,N_4531,N_4635);
nor U5768 (N_5768,N_4774,N_4177);
nand U5769 (N_5769,N_4723,N_4362);
and U5770 (N_5770,N_4919,N_4178);
nor U5771 (N_5771,N_4725,N_4045);
or U5772 (N_5772,N_4712,N_4888);
or U5773 (N_5773,N_4586,N_4228);
or U5774 (N_5774,N_4198,N_4144);
or U5775 (N_5775,N_4504,N_4059);
nand U5776 (N_5776,N_4697,N_4178);
xnor U5777 (N_5777,N_4986,N_4494);
nor U5778 (N_5778,N_4133,N_4336);
nand U5779 (N_5779,N_4064,N_4858);
and U5780 (N_5780,N_4355,N_4408);
nand U5781 (N_5781,N_4740,N_4982);
nor U5782 (N_5782,N_4836,N_4762);
and U5783 (N_5783,N_4861,N_4713);
or U5784 (N_5784,N_4122,N_4968);
and U5785 (N_5785,N_4364,N_4922);
and U5786 (N_5786,N_4700,N_4892);
and U5787 (N_5787,N_4499,N_4206);
xor U5788 (N_5788,N_4002,N_4947);
xor U5789 (N_5789,N_4490,N_4671);
or U5790 (N_5790,N_4549,N_4028);
or U5791 (N_5791,N_4713,N_4982);
nor U5792 (N_5792,N_4826,N_4506);
and U5793 (N_5793,N_4466,N_4258);
or U5794 (N_5794,N_4985,N_4594);
and U5795 (N_5795,N_4887,N_4268);
or U5796 (N_5796,N_4712,N_4884);
nor U5797 (N_5797,N_4416,N_4086);
xor U5798 (N_5798,N_4624,N_4805);
xor U5799 (N_5799,N_4240,N_4867);
nor U5800 (N_5800,N_4968,N_4065);
nor U5801 (N_5801,N_4133,N_4498);
nand U5802 (N_5802,N_4265,N_4625);
nor U5803 (N_5803,N_4829,N_4268);
and U5804 (N_5804,N_4077,N_4601);
or U5805 (N_5805,N_4663,N_4132);
and U5806 (N_5806,N_4362,N_4480);
xor U5807 (N_5807,N_4327,N_4023);
nand U5808 (N_5808,N_4468,N_4177);
or U5809 (N_5809,N_4675,N_4590);
nor U5810 (N_5810,N_4059,N_4801);
nand U5811 (N_5811,N_4855,N_4280);
nor U5812 (N_5812,N_4620,N_4401);
or U5813 (N_5813,N_4879,N_4151);
and U5814 (N_5814,N_4641,N_4578);
nand U5815 (N_5815,N_4704,N_4961);
nor U5816 (N_5816,N_4981,N_4701);
nor U5817 (N_5817,N_4336,N_4579);
and U5818 (N_5818,N_4575,N_4454);
or U5819 (N_5819,N_4745,N_4888);
xnor U5820 (N_5820,N_4353,N_4238);
nand U5821 (N_5821,N_4824,N_4803);
xor U5822 (N_5822,N_4959,N_4700);
xor U5823 (N_5823,N_4921,N_4396);
xnor U5824 (N_5824,N_4780,N_4342);
and U5825 (N_5825,N_4030,N_4442);
nand U5826 (N_5826,N_4164,N_4702);
xnor U5827 (N_5827,N_4302,N_4411);
and U5828 (N_5828,N_4462,N_4679);
nand U5829 (N_5829,N_4349,N_4792);
or U5830 (N_5830,N_4546,N_4998);
nand U5831 (N_5831,N_4059,N_4701);
nand U5832 (N_5832,N_4936,N_4046);
and U5833 (N_5833,N_4286,N_4285);
nor U5834 (N_5834,N_4060,N_4605);
nand U5835 (N_5835,N_4499,N_4235);
nor U5836 (N_5836,N_4587,N_4393);
and U5837 (N_5837,N_4102,N_4445);
or U5838 (N_5838,N_4075,N_4053);
nand U5839 (N_5839,N_4217,N_4472);
or U5840 (N_5840,N_4641,N_4078);
and U5841 (N_5841,N_4149,N_4644);
nor U5842 (N_5842,N_4409,N_4878);
nor U5843 (N_5843,N_4480,N_4317);
xnor U5844 (N_5844,N_4045,N_4063);
nor U5845 (N_5845,N_4436,N_4854);
nor U5846 (N_5846,N_4153,N_4687);
nand U5847 (N_5847,N_4882,N_4903);
nor U5848 (N_5848,N_4458,N_4079);
and U5849 (N_5849,N_4973,N_4722);
xor U5850 (N_5850,N_4543,N_4894);
and U5851 (N_5851,N_4543,N_4117);
nand U5852 (N_5852,N_4279,N_4774);
nor U5853 (N_5853,N_4716,N_4049);
or U5854 (N_5854,N_4047,N_4305);
and U5855 (N_5855,N_4362,N_4855);
nand U5856 (N_5856,N_4627,N_4119);
or U5857 (N_5857,N_4172,N_4256);
nor U5858 (N_5858,N_4212,N_4019);
nor U5859 (N_5859,N_4577,N_4975);
nor U5860 (N_5860,N_4197,N_4093);
nor U5861 (N_5861,N_4189,N_4301);
or U5862 (N_5862,N_4857,N_4151);
and U5863 (N_5863,N_4155,N_4244);
and U5864 (N_5864,N_4689,N_4792);
or U5865 (N_5865,N_4838,N_4011);
nor U5866 (N_5866,N_4909,N_4551);
nand U5867 (N_5867,N_4718,N_4016);
and U5868 (N_5868,N_4776,N_4438);
nor U5869 (N_5869,N_4260,N_4555);
and U5870 (N_5870,N_4438,N_4260);
nand U5871 (N_5871,N_4548,N_4719);
or U5872 (N_5872,N_4629,N_4737);
nor U5873 (N_5873,N_4455,N_4914);
or U5874 (N_5874,N_4036,N_4038);
or U5875 (N_5875,N_4567,N_4258);
or U5876 (N_5876,N_4499,N_4750);
and U5877 (N_5877,N_4008,N_4573);
nand U5878 (N_5878,N_4460,N_4701);
nor U5879 (N_5879,N_4161,N_4430);
and U5880 (N_5880,N_4586,N_4723);
or U5881 (N_5881,N_4291,N_4149);
xnor U5882 (N_5882,N_4432,N_4488);
nor U5883 (N_5883,N_4899,N_4620);
or U5884 (N_5884,N_4560,N_4853);
nand U5885 (N_5885,N_4754,N_4646);
and U5886 (N_5886,N_4560,N_4571);
nand U5887 (N_5887,N_4146,N_4515);
nor U5888 (N_5888,N_4033,N_4051);
and U5889 (N_5889,N_4657,N_4235);
nand U5890 (N_5890,N_4021,N_4708);
nor U5891 (N_5891,N_4975,N_4391);
and U5892 (N_5892,N_4513,N_4306);
nand U5893 (N_5893,N_4011,N_4463);
nand U5894 (N_5894,N_4413,N_4363);
or U5895 (N_5895,N_4196,N_4530);
nand U5896 (N_5896,N_4703,N_4309);
nor U5897 (N_5897,N_4126,N_4155);
and U5898 (N_5898,N_4840,N_4134);
nor U5899 (N_5899,N_4083,N_4583);
xnor U5900 (N_5900,N_4384,N_4097);
nor U5901 (N_5901,N_4017,N_4083);
nand U5902 (N_5902,N_4597,N_4735);
and U5903 (N_5903,N_4651,N_4214);
or U5904 (N_5904,N_4098,N_4151);
and U5905 (N_5905,N_4525,N_4530);
nand U5906 (N_5906,N_4486,N_4634);
and U5907 (N_5907,N_4888,N_4859);
xnor U5908 (N_5908,N_4348,N_4780);
or U5909 (N_5909,N_4717,N_4573);
xnor U5910 (N_5910,N_4743,N_4224);
xor U5911 (N_5911,N_4390,N_4248);
nand U5912 (N_5912,N_4359,N_4758);
nand U5913 (N_5913,N_4217,N_4106);
or U5914 (N_5914,N_4871,N_4196);
nor U5915 (N_5915,N_4927,N_4916);
or U5916 (N_5916,N_4958,N_4582);
and U5917 (N_5917,N_4795,N_4662);
nor U5918 (N_5918,N_4607,N_4345);
nand U5919 (N_5919,N_4618,N_4954);
nor U5920 (N_5920,N_4033,N_4590);
and U5921 (N_5921,N_4551,N_4839);
nand U5922 (N_5922,N_4865,N_4300);
nor U5923 (N_5923,N_4758,N_4109);
nor U5924 (N_5924,N_4559,N_4936);
or U5925 (N_5925,N_4644,N_4265);
and U5926 (N_5926,N_4545,N_4060);
and U5927 (N_5927,N_4952,N_4681);
and U5928 (N_5928,N_4318,N_4307);
nand U5929 (N_5929,N_4545,N_4517);
nor U5930 (N_5930,N_4975,N_4167);
nor U5931 (N_5931,N_4711,N_4769);
nand U5932 (N_5932,N_4386,N_4679);
or U5933 (N_5933,N_4596,N_4616);
nor U5934 (N_5934,N_4303,N_4255);
nand U5935 (N_5935,N_4454,N_4989);
and U5936 (N_5936,N_4662,N_4820);
nor U5937 (N_5937,N_4717,N_4870);
and U5938 (N_5938,N_4814,N_4467);
nand U5939 (N_5939,N_4837,N_4477);
nand U5940 (N_5940,N_4995,N_4035);
or U5941 (N_5941,N_4990,N_4937);
or U5942 (N_5942,N_4640,N_4517);
nand U5943 (N_5943,N_4294,N_4134);
and U5944 (N_5944,N_4238,N_4047);
nor U5945 (N_5945,N_4817,N_4702);
nand U5946 (N_5946,N_4303,N_4469);
and U5947 (N_5947,N_4776,N_4519);
and U5948 (N_5948,N_4812,N_4117);
or U5949 (N_5949,N_4783,N_4337);
nor U5950 (N_5950,N_4755,N_4400);
and U5951 (N_5951,N_4165,N_4342);
or U5952 (N_5952,N_4957,N_4162);
nor U5953 (N_5953,N_4715,N_4309);
and U5954 (N_5954,N_4683,N_4659);
and U5955 (N_5955,N_4454,N_4363);
nor U5956 (N_5956,N_4643,N_4260);
and U5957 (N_5957,N_4461,N_4276);
and U5958 (N_5958,N_4734,N_4132);
nand U5959 (N_5959,N_4987,N_4291);
or U5960 (N_5960,N_4777,N_4966);
and U5961 (N_5961,N_4881,N_4518);
or U5962 (N_5962,N_4446,N_4828);
nand U5963 (N_5963,N_4183,N_4267);
xor U5964 (N_5964,N_4941,N_4018);
nor U5965 (N_5965,N_4767,N_4673);
nor U5966 (N_5966,N_4287,N_4627);
nand U5967 (N_5967,N_4221,N_4670);
xnor U5968 (N_5968,N_4342,N_4258);
or U5969 (N_5969,N_4400,N_4611);
nand U5970 (N_5970,N_4242,N_4584);
xnor U5971 (N_5971,N_4406,N_4135);
xnor U5972 (N_5972,N_4905,N_4864);
nand U5973 (N_5973,N_4426,N_4132);
nand U5974 (N_5974,N_4740,N_4039);
or U5975 (N_5975,N_4969,N_4774);
and U5976 (N_5976,N_4848,N_4910);
nor U5977 (N_5977,N_4297,N_4186);
xnor U5978 (N_5978,N_4025,N_4629);
nand U5979 (N_5979,N_4738,N_4430);
nor U5980 (N_5980,N_4087,N_4930);
xor U5981 (N_5981,N_4932,N_4188);
nand U5982 (N_5982,N_4985,N_4682);
nor U5983 (N_5983,N_4263,N_4792);
nor U5984 (N_5984,N_4728,N_4910);
or U5985 (N_5985,N_4416,N_4790);
nand U5986 (N_5986,N_4004,N_4612);
nor U5987 (N_5987,N_4254,N_4987);
nand U5988 (N_5988,N_4359,N_4396);
and U5989 (N_5989,N_4833,N_4994);
nor U5990 (N_5990,N_4805,N_4852);
or U5991 (N_5991,N_4256,N_4549);
nor U5992 (N_5992,N_4479,N_4080);
and U5993 (N_5993,N_4826,N_4129);
or U5994 (N_5994,N_4819,N_4328);
or U5995 (N_5995,N_4863,N_4882);
or U5996 (N_5996,N_4651,N_4639);
and U5997 (N_5997,N_4201,N_4961);
and U5998 (N_5998,N_4436,N_4313);
and U5999 (N_5999,N_4669,N_4795);
or U6000 (N_6000,N_5317,N_5666);
nor U6001 (N_6001,N_5848,N_5897);
nand U6002 (N_6002,N_5827,N_5031);
nor U6003 (N_6003,N_5047,N_5923);
and U6004 (N_6004,N_5575,N_5696);
or U6005 (N_6005,N_5995,N_5570);
and U6006 (N_6006,N_5680,N_5427);
or U6007 (N_6007,N_5414,N_5488);
and U6008 (N_6008,N_5523,N_5416);
nor U6009 (N_6009,N_5049,N_5147);
nor U6010 (N_6010,N_5653,N_5249);
or U6011 (N_6011,N_5567,N_5189);
nand U6012 (N_6012,N_5333,N_5522);
or U6013 (N_6013,N_5557,N_5423);
or U6014 (N_6014,N_5664,N_5002);
or U6015 (N_6015,N_5734,N_5795);
and U6016 (N_6016,N_5603,N_5063);
nor U6017 (N_6017,N_5999,N_5106);
xnor U6018 (N_6018,N_5324,N_5041);
and U6019 (N_6019,N_5449,N_5238);
nor U6020 (N_6020,N_5320,N_5405);
and U6021 (N_6021,N_5170,N_5313);
nor U6022 (N_6022,N_5837,N_5937);
nand U6023 (N_6023,N_5747,N_5291);
and U6024 (N_6024,N_5207,N_5472);
xor U6025 (N_6025,N_5658,N_5213);
nor U6026 (N_6026,N_5023,N_5620);
and U6027 (N_6027,N_5683,N_5770);
nand U6028 (N_6028,N_5516,N_5726);
nor U6029 (N_6029,N_5276,N_5219);
nand U6030 (N_6030,N_5681,N_5661);
or U6031 (N_6031,N_5407,N_5775);
and U6032 (N_6032,N_5275,N_5673);
nor U6033 (N_6033,N_5075,N_5255);
or U6034 (N_6034,N_5555,N_5201);
and U6035 (N_6035,N_5781,N_5045);
nand U6036 (N_6036,N_5037,N_5505);
or U6037 (N_6037,N_5057,N_5233);
or U6038 (N_6038,N_5076,N_5993);
and U6039 (N_6039,N_5308,N_5182);
xor U6040 (N_6040,N_5660,N_5107);
xnor U6041 (N_6041,N_5436,N_5003);
and U6042 (N_6042,N_5105,N_5264);
nor U6043 (N_6043,N_5828,N_5062);
or U6044 (N_6044,N_5569,N_5445);
or U6045 (N_6045,N_5392,N_5192);
xor U6046 (N_6046,N_5038,N_5117);
and U6047 (N_6047,N_5307,N_5145);
and U6048 (N_6048,N_5872,N_5403);
and U6049 (N_6049,N_5527,N_5724);
or U6050 (N_6050,N_5549,N_5826);
and U6051 (N_6051,N_5292,N_5492);
nand U6052 (N_6052,N_5645,N_5080);
nand U6053 (N_6053,N_5118,N_5210);
nor U6054 (N_6054,N_5791,N_5929);
nand U6055 (N_6055,N_5256,N_5875);
and U6056 (N_6056,N_5285,N_5853);
and U6057 (N_6057,N_5074,N_5232);
nand U6058 (N_6058,N_5573,N_5565);
or U6059 (N_6059,N_5688,N_5939);
or U6060 (N_6060,N_5882,N_5874);
and U6061 (N_6061,N_5335,N_5040);
nand U6062 (N_6062,N_5919,N_5936);
or U6063 (N_6063,N_5452,N_5027);
and U6064 (N_6064,N_5904,N_5352);
nor U6065 (N_6065,N_5588,N_5617);
or U6066 (N_6066,N_5315,N_5166);
nor U6067 (N_6067,N_5363,N_5813);
or U6068 (N_6068,N_5772,N_5873);
nor U6069 (N_6069,N_5446,N_5239);
or U6070 (N_6070,N_5650,N_5996);
or U6071 (N_6071,N_5950,N_5404);
nand U6072 (N_6072,N_5191,N_5598);
or U6073 (N_6073,N_5641,N_5672);
nand U6074 (N_6074,N_5684,N_5913);
nand U6075 (N_6075,N_5685,N_5532);
xor U6076 (N_6076,N_5022,N_5938);
or U6077 (N_6077,N_5224,N_5431);
or U6078 (N_6078,N_5587,N_5218);
xnor U6079 (N_6079,N_5368,N_5310);
or U6080 (N_6080,N_5528,N_5530);
nand U6081 (N_6081,N_5349,N_5695);
or U6082 (N_6082,N_5958,N_5116);
nor U6083 (N_6083,N_5907,N_5659);
nor U6084 (N_6084,N_5364,N_5010);
or U6085 (N_6085,N_5082,N_5410);
and U6086 (N_6086,N_5894,N_5111);
and U6087 (N_6087,N_5036,N_5931);
nand U6088 (N_6088,N_5718,N_5148);
nor U6089 (N_6089,N_5595,N_5776);
nand U6090 (N_6090,N_5044,N_5177);
and U6091 (N_6091,N_5584,N_5017);
and U6092 (N_6092,N_5924,N_5453);
and U6093 (N_6093,N_5836,N_5130);
nor U6094 (N_6094,N_5289,N_5294);
and U6095 (N_6095,N_5822,N_5927);
nand U6096 (N_6096,N_5091,N_5640);
or U6097 (N_6097,N_5120,N_5521);
and U6098 (N_6098,N_5139,N_5835);
and U6099 (N_6099,N_5069,N_5771);
and U6100 (N_6100,N_5839,N_5710);
and U6101 (N_6101,N_5476,N_5773);
and U6102 (N_6102,N_5329,N_5845);
and U6103 (N_6103,N_5341,N_5325);
or U6104 (N_6104,N_5042,N_5344);
nand U6105 (N_6105,N_5375,N_5277);
nand U6106 (N_6106,N_5388,N_5783);
xnor U6107 (N_6107,N_5437,N_5541);
nor U6108 (N_6108,N_5860,N_5486);
or U6109 (N_6109,N_5000,N_5953);
or U6110 (N_6110,N_5579,N_5322);
or U6111 (N_6111,N_5008,N_5803);
or U6112 (N_6112,N_5149,N_5367);
or U6113 (N_6113,N_5831,N_5493);
or U6114 (N_6114,N_5297,N_5581);
or U6115 (N_6115,N_5078,N_5430);
nand U6116 (N_6116,N_5426,N_5462);
or U6117 (N_6117,N_5127,N_5752);
nor U6118 (N_6118,N_5735,N_5691);
nor U6119 (N_6119,N_5095,N_5764);
or U6120 (N_6120,N_5172,N_5881);
nor U6121 (N_6121,N_5682,N_5585);
nand U6122 (N_6122,N_5073,N_5215);
and U6123 (N_6123,N_5035,N_5384);
nand U6124 (N_6124,N_5347,N_5840);
or U6125 (N_6125,N_5843,N_5917);
nand U6126 (N_6126,N_5459,N_5343);
xor U6127 (N_6127,N_5195,N_5976);
xor U6128 (N_6128,N_5876,N_5287);
or U6129 (N_6129,N_5101,N_5456);
nand U6130 (N_6130,N_5693,N_5054);
or U6131 (N_6131,N_5634,N_5507);
nand U6132 (N_6132,N_5305,N_5217);
or U6133 (N_6133,N_5885,N_5360);
or U6134 (N_6134,N_5274,N_5494);
nand U6135 (N_6135,N_5975,N_5478);
nor U6136 (N_6136,N_5815,N_5789);
nor U6137 (N_6137,N_5371,N_5266);
and U6138 (N_6138,N_5737,N_5121);
and U6139 (N_6139,N_5396,N_5269);
or U6140 (N_6140,N_5786,N_5173);
or U6141 (N_6141,N_5674,N_5484);
xnor U6142 (N_6142,N_5546,N_5060);
and U6143 (N_6143,N_5161,N_5338);
or U6144 (N_6144,N_5155,N_5960);
nor U6145 (N_6145,N_5778,N_5841);
or U6146 (N_6146,N_5804,N_5460);
nor U6147 (N_6147,N_5479,N_5918);
or U6148 (N_6148,N_5671,N_5471);
or U6149 (N_6149,N_5663,N_5957);
nand U6150 (N_6150,N_5817,N_5176);
nor U6151 (N_6151,N_5808,N_5390);
or U6152 (N_6152,N_5065,N_5200);
xnor U6153 (N_6153,N_5756,N_5151);
and U6154 (N_6154,N_5531,N_5928);
nor U6155 (N_6155,N_5337,N_5857);
nand U6156 (N_6156,N_5336,N_5199);
and U6157 (N_6157,N_5518,N_5879);
and U6158 (N_6158,N_5119,N_5485);
nand U6159 (N_6159,N_5643,N_5668);
nor U6160 (N_6160,N_5366,N_5758);
and U6161 (N_6161,N_5513,N_5965);
or U6162 (N_6162,N_5212,N_5989);
and U6163 (N_6163,N_5970,N_5769);
and U6164 (N_6164,N_5805,N_5690);
or U6165 (N_6165,N_5382,N_5866);
and U6166 (N_6166,N_5158,N_5015);
xor U6167 (N_6167,N_5739,N_5689);
and U6168 (N_6168,N_5052,N_5342);
nor U6169 (N_6169,N_5417,N_5296);
xor U6170 (N_6170,N_5900,N_5606);
nor U6171 (N_6171,N_5226,N_5257);
nand U6172 (N_6172,N_5464,N_5766);
nor U6173 (N_6173,N_5056,N_5092);
nor U6174 (N_6174,N_5635,N_5589);
or U6175 (N_6175,N_5252,N_5951);
nand U6176 (N_6176,N_5141,N_5438);
nor U6177 (N_6177,N_5153,N_5021);
nor U6178 (N_6178,N_5601,N_5009);
and U6179 (N_6179,N_5451,N_5812);
nor U6180 (N_6180,N_5966,N_5798);
and U6181 (N_6181,N_5030,N_5702);
or U6182 (N_6182,N_5962,N_5748);
nor U6183 (N_6183,N_5448,N_5895);
and U6184 (N_6184,N_5072,N_5309);
and U6185 (N_6185,N_5593,N_5997);
and U6186 (N_6186,N_5259,N_5649);
xnor U6187 (N_6187,N_5556,N_5590);
and U6188 (N_6188,N_5229,N_5942);
nand U6189 (N_6189,N_5892,N_5946);
or U6190 (N_6190,N_5744,N_5051);
nand U6191 (N_6191,N_5420,N_5301);
or U6192 (N_6192,N_5415,N_5655);
nor U6193 (N_6193,N_5699,N_5190);
xor U6194 (N_6194,N_5519,N_5605);
nand U6195 (N_6195,N_5741,N_5851);
nor U6196 (N_6196,N_5834,N_5858);
nor U6197 (N_6197,N_5466,N_5183);
nand U6198 (N_6198,N_5461,N_5214);
nor U6199 (N_6199,N_5323,N_5355);
or U6200 (N_6200,N_5043,N_5794);
or U6201 (N_6201,N_5001,N_5779);
xor U6202 (N_6202,N_5914,N_5811);
nand U6203 (N_6203,N_5284,N_5004);
and U6204 (N_6204,N_5441,N_5562);
xnor U6205 (N_6205,N_5524,N_5094);
and U6206 (N_6206,N_5319,N_5429);
or U6207 (N_6207,N_5497,N_5994);
and U6208 (N_6208,N_5508,N_5891);
nor U6209 (N_6209,N_5450,N_5220);
xnor U6210 (N_6210,N_5945,N_5638);
nand U6211 (N_6211,N_5386,N_5361);
and U6212 (N_6212,N_5893,N_5502);
or U6213 (N_6213,N_5328,N_5458);
and U6214 (N_6214,N_5053,N_5399);
xnor U6215 (N_6215,N_5402,N_5868);
or U6216 (N_6216,N_5221,N_5236);
nor U6217 (N_6217,N_5412,N_5700);
or U6218 (N_6218,N_5991,N_5086);
nor U6219 (N_6219,N_5596,N_5108);
nand U6220 (N_6220,N_5012,N_5934);
xor U6221 (N_6221,N_5963,N_5644);
nor U6222 (N_6222,N_5187,N_5064);
and U6223 (N_6223,N_5548,N_5122);
or U6224 (N_6224,N_5085,N_5646);
nand U6225 (N_6225,N_5967,N_5662);
nand U6226 (N_6226,N_5708,N_5818);
nor U6227 (N_6227,N_5146,N_5964);
and U6228 (N_6228,N_5428,N_5171);
nand U6229 (N_6229,N_5819,N_5852);
or U6230 (N_6230,N_5165,N_5642);
nor U6231 (N_6231,N_5088,N_5314);
nand U6232 (N_6232,N_5160,N_5612);
or U6233 (N_6233,N_5457,N_5408);
nand U6234 (N_6234,N_5767,N_5586);
nor U6235 (N_6235,N_5365,N_5824);
and U6236 (N_6236,N_5114,N_5348);
and U6237 (N_6237,N_5554,N_5793);
xnor U6238 (N_6238,N_5247,N_5254);
or U6239 (N_6239,N_5722,N_5880);
or U6240 (N_6240,N_5330,N_5526);
and U6241 (N_6241,N_5334,N_5385);
nand U6242 (N_6242,N_5616,N_5503);
nor U6243 (N_6243,N_5514,N_5351);
nor U6244 (N_6244,N_5736,N_5915);
and U6245 (N_6245,N_5952,N_5847);
nand U6246 (N_6246,N_5574,N_5669);
or U6247 (N_6247,N_5714,N_5283);
or U6248 (N_6248,N_5228,N_5547);
nand U6249 (N_6249,N_5512,N_5704);
and U6250 (N_6250,N_5707,N_5757);
and U6251 (N_6251,N_5357,N_5765);
nor U6252 (N_6252,N_5482,N_5622);
nand U6253 (N_6253,N_5988,N_5205);
nor U6254 (N_6254,N_5679,N_5186);
nor U6255 (N_6255,N_5667,N_5721);
nand U6256 (N_6256,N_5697,N_5084);
nand U6257 (N_6257,N_5899,N_5856);
nand U6258 (N_6258,N_5079,N_5943);
and U6259 (N_6259,N_5792,N_5340);
nor U6260 (N_6260,N_5398,N_5169);
or U6261 (N_6261,N_5312,N_5395);
nand U6262 (N_6262,N_5142,N_5369);
nand U6263 (N_6263,N_5763,N_5090);
or U6264 (N_6264,N_5443,N_5240);
and U6265 (N_6265,N_5018,N_5820);
and U6266 (N_6266,N_5933,N_5124);
nand U6267 (N_6267,N_5947,N_5552);
and U6268 (N_6268,N_5944,N_5903);
or U6269 (N_6269,N_5103,N_5258);
nand U6270 (N_6270,N_5273,N_5339);
nand U6271 (N_6271,N_5926,N_5611);
nor U6272 (N_6272,N_5354,N_5067);
nor U6273 (N_6273,N_5814,N_5675);
or U6274 (N_6274,N_5849,N_5159);
or U6275 (N_6275,N_5123,N_5833);
nor U6276 (N_6276,N_5925,N_5318);
nor U6277 (N_6277,N_5539,N_5433);
or U6278 (N_6278,N_5209,N_5203);
nor U6279 (N_6279,N_5393,N_5627);
and U6280 (N_6280,N_5235,N_5790);
nor U6281 (N_6281,N_5442,N_5738);
nor U6282 (N_6282,N_5796,N_5614);
or U6283 (N_6283,N_5633,N_5916);
nor U6284 (N_6284,N_5846,N_5353);
or U6285 (N_6285,N_5089,N_5138);
nor U6286 (N_6286,N_5136,N_5906);
nor U6287 (N_6287,N_5715,N_5571);
nor U6288 (N_6288,N_5972,N_5949);
or U6289 (N_6289,N_5394,N_5961);
nor U6290 (N_6290,N_5740,N_5987);
nand U6291 (N_6291,N_5582,N_5474);
or U6292 (N_6292,N_5855,N_5729);
or U6293 (N_6293,N_5941,N_5711);
xnor U6294 (N_6294,N_5954,N_5743);
nor U6295 (N_6295,N_5432,N_5577);
or U6296 (N_6296,N_5332,N_5720);
and U6297 (N_6297,N_5162,N_5609);
xnor U6298 (N_6298,N_5538,N_5447);
and U6299 (N_6299,N_5306,N_5801);
nand U6300 (N_6300,N_5745,N_5629);
nand U6301 (N_6301,N_5179,N_5241);
and U6302 (N_6302,N_5288,N_5025);
nand U6303 (N_6303,N_5129,N_5534);
and U6304 (N_6304,N_5409,N_5345);
nand U6305 (N_6305,N_5782,N_5498);
and U6306 (N_6306,N_5016,N_5560);
and U6307 (N_6307,N_5270,N_5359);
and U6308 (N_6308,N_5424,N_5419);
and U6309 (N_6309,N_5185,N_5754);
nand U6310 (N_6310,N_5039,N_5637);
or U6311 (N_6311,N_5104,N_5865);
nor U6312 (N_6312,N_5143,N_5180);
nor U6313 (N_6313,N_5413,N_5356);
nor U6314 (N_6314,N_5712,N_5135);
or U6315 (N_6315,N_5376,N_5973);
nor U6316 (N_6316,N_5391,N_5243);
nor U6317 (N_6317,N_5750,N_5971);
or U6318 (N_6318,N_5193,N_5558);
and U6319 (N_6319,N_5290,N_5703);
or U6320 (N_6320,N_5777,N_5517);
or U6321 (N_6321,N_5483,N_5265);
nand U6322 (N_6322,N_5033,N_5863);
and U6323 (N_6323,N_5525,N_5678);
and U6324 (N_6324,N_5204,N_5751);
nand U6325 (N_6325,N_5597,N_5550);
xnor U6326 (N_6326,N_5807,N_5346);
nand U6327 (N_6327,N_5261,N_5959);
nand U6328 (N_6328,N_5006,N_5373);
nand U6329 (N_6329,N_5990,N_5639);
or U6330 (N_6330,N_5687,N_5379);
and U6331 (N_6331,N_5623,N_5746);
or U6332 (N_6332,N_5480,N_5955);
xor U6333 (N_6333,N_5245,N_5400);
and U6334 (N_6334,N_5383,N_5665);
xor U6335 (N_6335,N_5850,N_5761);
or U6336 (N_6336,N_5061,N_5867);
and U6337 (N_6337,N_5974,N_5133);
nand U6338 (N_6338,N_5607,N_5491);
or U6339 (N_6339,N_5861,N_5029);
nor U6340 (N_6340,N_5048,N_5227);
or U6341 (N_6341,N_5592,N_5272);
or U6342 (N_6342,N_5096,N_5293);
or U6343 (N_6343,N_5097,N_5331);
nor U6344 (N_6344,N_5178,N_5206);
and U6345 (N_6345,N_5225,N_5600);
or U6346 (N_6346,N_5401,N_5501);
nand U6347 (N_6347,N_5830,N_5223);
nand U6348 (N_6348,N_5864,N_5742);
nand U6349 (N_6349,N_5081,N_5568);
nand U6350 (N_6350,N_5537,N_5599);
or U6351 (N_6351,N_5071,N_5544);
and U6352 (N_6352,N_5250,N_5780);
or U6353 (N_6353,N_5760,N_5905);
nor U6354 (N_6354,N_5490,N_5087);
xor U6355 (N_6355,N_5198,N_5878);
or U6356 (N_6356,N_5618,N_5175);
and U6357 (N_6357,N_5140,N_5869);
and U6358 (N_6358,N_5421,N_5098);
and U6359 (N_6359,N_5150,N_5896);
nand U6360 (N_6360,N_5477,N_5887);
nor U6361 (N_6361,N_5231,N_5467);
and U6362 (N_6362,N_5099,N_5890);
or U6363 (N_6363,N_5604,N_5469);
xnor U6364 (N_6364,N_5908,N_5630);
and U6365 (N_6365,N_5730,N_5034);
nand U6366 (N_6366,N_5920,N_5529);
nor U6367 (N_6367,N_5709,N_5268);
nor U6368 (N_6368,N_5475,N_5020);
or U6369 (N_6369,N_5248,N_5216);
nor U6370 (N_6370,N_5998,N_5083);
nor U6371 (N_6371,N_5838,N_5984);
nor U6372 (N_6372,N_5912,N_5434);
nand U6373 (N_6373,N_5188,N_5610);
or U6374 (N_6374,N_5370,N_5888);
and U6375 (N_6375,N_5632,N_5281);
nand U6376 (N_6376,N_5326,N_5468);
xnor U6377 (N_6377,N_5732,N_5759);
and U6378 (N_6378,N_5626,N_5059);
nand U6379 (N_6379,N_5473,N_5591);
or U6380 (N_6380,N_5444,N_5762);
nor U6381 (N_6381,N_5686,N_5982);
nor U6382 (N_6382,N_5489,N_5652);
nand U6383 (N_6383,N_5321,N_5230);
nand U6384 (N_6384,N_5350,N_5797);
or U6385 (N_6385,N_5411,N_5208);
and U6386 (N_6386,N_5316,N_5435);
and U6387 (N_6387,N_5271,N_5125);
xnor U6388 (N_6388,N_5280,N_5551);
nand U6389 (N_6389,N_5676,N_5511);
nor U6390 (N_6390,N_5768,N_5692);
or U6391 (N_6391,N_5168,N_5901);
or U6392 (N_6392,N_5911,N_5728);
nor U6393 (N_6393,N_5608,N_5594);
or U6394 (N_6394,N_5300,N_5564);
or U6395 (N_6395,N_5774,N_5628);
or U6396 (N_6396,N_5279,N_5540);
nand U6397 (N_6397,N_5303,N_5563);
nor U6398 (N_6398,N_5026,N_5253);
and U6399 (N_6399,N_5509,N_5948);
or U6400 (N_6400,N_5237,N_5242);
nor U6401 (N_6401,N_5028,N_5749);
nor U6402 (N_6402,N_5621,N_5810);
nand U6403 (N_6403,N_5282,N_5506);
or U6404 (N_6404,N_5439,N_5977);
xor U6405 (N_6405,N_5504,N_5755);
nor U6406 (N_6406,N_5134,N_5753);
and U6407 (N_6407,N_5295,N_5883);
nor U6408 (N_6408,N_5992,N_5387);
and U6409 (N_6409,N_5922,N_5286);
and U6410 (N_6410,N_5802,N_5533);
nand U6411 (N_6411,N_5184,N_5727);
and U6412 (N_6412,N_5377,N_5131);
xor U6413 (N_6413,N_5656,N_5799);
and U6414 (N_6414,N_5543,N_5495);
or U6415 (N_6415,N_5418,N_5113);
xnor U6416 (N_6416,N_5921,N_5372);
and U6417 (N_6417,N_5935,N_5785);
and U6418 (N_6418,N_5499,N_5378);
or U6419 (N_6419,N_5299,N_5093);
and U6420 (N_6420,N_5066,N_5234);
nor U6421 (N_6421,N_5164,N_5454);
xor U6422 (N_6422,N_5670,N_5007);
nand U6423 (N_6423,N_5898,N_5058);
or U6424 (N_6424,N_5077,N_5070);
nand U6425 (N_6425,N_5809,N_5909);
nand U6426 (N_6426,N_5583,N_5545);
nor U6427 (N_6427,N_5302,N_5859);
and U6428 (N_6428,N_5154,N_5157);
nand U6429 (N_6429,N_5536,N_5717);
nor U6430 (N_6430,N_5196,N_5102);
nor U6431 (N_6431,N_5397,N_5535);
or U6432 (N_6432,N_5985,N_5625);
nor U6433 (N_6433,N_5406,N_5829);
xnor U6434 (N_6434,N_5654,N_5055);
and U6435 (N_6435,N_5870,N_5211);
or U6436 (N_6436,N_5481,N_5262);
nand U6437 (N_6437,N_5602,N_5787);
nand U6438 (N_6438,N_5422,N_5024);
nor U6439 (N_6439,N_5716,N_5005);
xor U6440 (N_6440,N_5821,N_5278);
or U6441 (N_6441,N_5520,N_5806);
or U6442 (N_6442,N_5886,N_5463);
nand U6443 (N_6443,N_5983,N_5733);
xor U6444 (N_6444,N_5978,N_5251);
xnor U6445 (N_6445,N_5362,N_5013);
nor U6446 (N_6446,N_5677,N_5425);
and U6447 (N_6447,N_5311,N_5152);
nand U6448 (N_6448,N_5842,N_5487);
nor U6449 (N_6449,N_5126,N_5380);
and U6450 (N_6450,N_5222,N_5014);
nand U6451 (N_6451,N_5167,N_5174);
xor U6452 (N_6452,N_5260,N_5496);
xnor U6453 (N_6453,N_5884,N_5011);
or U6454 (N_6454,N_5561,N_5455);
nand U6455 (N_6455,N_5019,N_5647);
nor U6456 (N_6456,N_5515,N_5862);
or U6457 (N_6457,N_5969,N_5381);
xor U6458 (N_6458,N_5542,N_5844);
and U6459 (N_6459,N_5636,N_5578);
nor U6460 (N_6460,N_5576,N_5816);
or U6461 (N_6461,N_5613,N_5832);
nor U6462 (N_6462,N_5800,N_5050);
or U6463 (N_6463,N_5374,N_5719);
nor U6464 (N_6464,N_5559,N_5784);
or U6465 (N_6465,N_5510,N_5110);
and U6466 (N_6466,N_5854,N_5877);
or U6467 (N_6467,N_5788,N_5694);
nor U6468 (N_6468,N_5705,N_5202);
or U6469 (N_6469,N_5619,N_5465);
or U6470 (N_6470,N_5871,N_5930);
and U6471 (N_6471,N_5197,N_5500);
and U6472 (N_6472,N_5304,N_5902);
xor U6473 (N_6473,N_5389,N_5657);
and U6474 (N_6474,N_5932,N_5706);
or U6475 (N_6475,N_5246,N_5440);
and U6476 (N_6476,N_5553,N_5132);
and U6477 (N_6477,N_5032,N_5194);
or U6478 (N_6478,N_5651,N_5327);
xor U6479 (N_6479,N_5358,N_5115);
or U6480 (N_6480,N_5701,N_5163);
nor U6481 (N_6481,N_5615,N_5631);
nor U6482 (N_6482,N_5979,N_5580);
and U6483 (N_6483,N_5156,N_5713);
nor U6484 (N_6484,N_5731,N_5109);
and U6485 (N_6485,N_5100,N_5980);
and U6486 (N_6486,N_5698,N_5956);
and U6487 (N_6487,N_5910,N_5244);
or U6488 (N_6488,N_5267,N_5624);
nor U6489 (N_6489,N_5940,N_5725);
nor U6490 (N_6490,N_5723,N_5128);
nor U6491 (N_6491,N_5986,N_5298);
nor U6492 (N_6492,N_5181,N_5046);
nor U6493 (N_6493,N_5112,N_5470);
nor U6494 (N_6494,N_5825,N_5648);
or U6495 (N_6495,N_5823,N_5572);
and U6496 (N_6496,N_5889,N_5068);
nor U6497 (N_6497,N_5144,N_5137);
or U6498 (N_6498,N_5566,N_5263);
xor U6499 (N_6499,N_5981,N_5968);
and U6500 (N_6500,N_5591,N_5318);
nand U6501 (N_6501,N_5338,N_5354);
and U6502 (N_6502,N_5815,N_5394);
nor U6503 (N_6503,N_5246,N_5967);
and U6504 (N_6504,N_5088,N_5052);
or U6505 (N_6505,N_5619,N_5536);
and U6506 (N_6506,N_5949,N_5894);
and U6507 (N_6507,N_5650,N_5057);
or U6508 (N_6508,N_5144,N_5094);
nor U6509 (N_6509,N_5232,N_5166);
or U6510 (N_6510,N_5153,N_5039);
xor U6511 (N_6511,N_5967,N_5915);
nor U6512 (N_6512,N_5511,N_5897);
nand U6513 (N_6513,N_5031,N_5249);
or U6514 (N_6514,N_5329,N_5868);
or U6515 (N_6515,N_5529,N_5927);
xor U6516 (N_6516,N_5137,N_5189);
nor U6517 (N_6517,N_5566,N_5017);
xor U6518 (N_6518,N_5581,N_5367);
xor U6519 (N_6519,N_5382,N_5953);
or U6520 (N_6520,N_5445,N_5350);
and U6521 (N_6521,N_5384,N_5655);
nand U6522 (N_6522,N_5657,N_5534);
nor U6523 (N_6523,N_5849,N_5814);
or U6524 (N_6524,N_5569,N_5438);
and U6525 (N_6525,N_5316,N_5993);
and U6526 (N_6526,N_5835,N_5158);
nor U6527 (N_6527,N_5418,N_5317);
nor U6528 (N_6528,N_5631,N_5940);
or U6529 (N_6529,N_5702,N_5540);
nand U6530 (N_6530,N_5391,N_5324);
xor U6531 (N_6531,N_5122,N_5025);
nor U6532 (N_6532,N_5099,N_5520);
or U6533 (N_6533,N_5962,N_5288);
nand U6534 (N_6534,N_5536,N_5760);
and U6535 (N_6535,N_5453,N_5916);
nand U6536 (N_6536,N_5458,N_5098);
or U6537 (N_6537,N_5954,N_5409);
nor U6538 (N_6538,N_5811,N_5265);
or U6539 (N_6539,N_5579,N_5539);
or U6540 (N_6540,N_5577,N_5788);
or U6541 (N_6541,N_5010,N_5374);
or U6542 (N_6542,N_5222,N_5033);
or U6543 (N_6543,N_5482,N_5155);
nand U6544 (N_6544,N_5465,N_5737);
or U6545 (N_6545,N_5730,N_5869);
nand U6546 (N_6546,N_5638,N_5735);
nor U6547 (N_6547,N_5448,N_5726);
and U6548 (N_6548,N_5682,N_5073);
and U6549 (N_6549,N_5597,N_5854);
nor U6550 (N_6550,N_5067,N_5843);
or U6551 (N_6551,N_5045,N_5780);
and U6552 (N_6552,N_5234,N_5721);
nor U6553 (N_6553,N_5064,N_5960);
or U6554 (N_6554,N_5619,N_5761);
and U6555 (N_6555,N_5082,N_5716);
nor U6556 (N_6556,N_5824,N_5550);
or U6557 (N_6557,N_5651,N_5196);
or U6558 (N_6558,N_5874,N_5159);
nor U6559 (N_6559,N_5188,N_5985);
nand U6560 (N_6560,N_5107,N_5935);
nand U6561 (N_6561,N_5611,N_5221);
and U6562 (N_6562,N_5082,N_5523);
nand U6563 (N_6563,N_5164,N_5913);
nand U6564 (N_6564,N_5742,N_5612);
or U6565 (N_6565,N_5125,N_5745);
nor U6566 (N_6566,N_5667,N_5773);
xor U6567 (N_6567,N_5434,N_5297);
nand U6568 (N_6568,N_5289,N_5633);
nor U6569 (N_6569,N_5590,N_5405);
and U6570 (N_6570,N_5074,N_5439);
nand U6571 (N_6571,N_5513,N_5885);
nor U6572 (N_6572,N_5817,N_5180);
and U6573 (N_6573,N_5569,N_5340);
nor U6574 (N_6574,N_5082,N_5889);
and U6575 (N_6575,N_5822,N_5737);
or U6576 (N_6576,N_5578,N_5501);
nand U6577 (N_6577,N_5289,N_5797);
nor U6578 (N_6578,N_5278,N_5102);
nor U6579 (N_6579,N_5839,N_5682);
and U6580 (N_6580,N_5472,N_5175);
nor U6581 (N_6581,N_5619,N_5722);
and U6582 (N_6582,N_5939,N_5062);
nor U6583 (N_6583,N_5633,N_5728);
nor U6584 (N_6584,N_5165,N_5891);
xor U6585 (N_6585,N_5433,N_5618);
or U6586 (N_6586,N_5868,N_5305);
or U6587 (N_6587,N_5287,N_5611);
and U6588 (N_6588,N_5635,N_5133);
nand U6589 (N_6589,N_5597,N_5996);
and U6590 (N_6590,N_5214,N_5464);
and U6591 (N_6591,N_5153,N_5130);
nand U6592 (N_6592,N_5947,N_5754);
and U6593 (N_6593,N_5607,N_5118);
or U6594 (N_6594,N_5293,N_5840);
nand U6595 (N_6595,N_5499,N_5089);
nor U6596 (N_6596,N_5678,N_5829);
or U6597 (N_6597,N_5111,N_5693);
nand U6598 (N_6598,N_5917,N_5842);
nor U6599 (N_6599,N_5607,N_5562);
nor U6600 (N_6600,N_5505,N_5758);
or U6601 (N_6601,N_5139,N_5393);
or U6602 (N_6602,N_5596,N_5447);
nor U6603 (N_6603,N_5869,N_5703);
or U6604 (N_6604,N_5018,N_5982);
nand U6605 (N_6605,N_5902,N_5495);
nand U6606 (N_6606,N_5918,N_5192);
or U6607 (N_6607,N_5461,N_5524);
or U6608 (N_6608,N_5225,N_5460);
nor U6609 (N_6609,N_5252,N_5161);
nand U6610 (N_6610,N_5981,N_5977);
nand U6611 (N_6611,N_5727,N_5449);
nand U6612 (N_6612,N_5639,N_5516);
nand U6613 (N_6613,N_5131,N_5376);
xor U6614 (N_6614,N_5493,N_5196);
nand U6615 (N_6615,N_5194,N_5930);
nand U6616 (N_6616,N_5858,N_5405);
and U6617 (N_6617,N_5052,N_5696);
and U6618 (N_6618,N_5694,N_5869);
or U6619 (N_6619,N_5419,N_5627);
nand U6620 (N_6620,N_5300,N_5526);
nand U6621 (N_6621,N_5964,N_5776);
xor U6622 (N_6622,N_5452,N_5229);
nor U6623 (N_6623,N_5858,N_5798);
and U6624 (N_6624,N_5530,N_5386);
and U6625 (N_6625,N_5667,N_5439);
nor U6626 (N_6626,N_5269,N_5051);
xnor U6627 (N_6627,N_5338,N_5318);
xor U6628 (N_6628,N_5262,N_5811);
xor U6629 (N_6629,N_5573,N_5239);
nand U6630 (N_6630,N_5516,N_5209);
nand U6631 (N_6631,N_5201,N_5149);
and U6632 (N_6632,N_5492,N_5682);
nor U6633 (N_6633,N_5859,N_5686);
nor U6634 (N_6634,N_5595,N_5040);
and U6635 (N_6635,N_5816,N_5450);
and U6636 (N_6636,N_5799,N_5257);
nand U6637 (N_6637,N_5677,N_5213);
and U6638 (N_6638,N_5576,N_5475);
and U6639 (N_6639,N_5935,N_5938);
xnor U6640 (N_6640,N_5477,N_5353);
nand U6641 (N_6641,N_5493,N_5467);
and U6642 (N_6642,N_5563,N_5956);
nand U6643 (N_6643,N_5352,N_5012);
nand U6644 (N_6644,N_5964,N_5538);
xnor U6645 (N_6645,N_5336,N_5096);
and U6646 (N_6646,N_5684,N_5589);
xnor U6647 (N_6647,N_5598,N_5390);
nor U6648 (N_6648,N_5804,N_5896);
nand U6649 (N_6649,N_5054,N_5375);
or U6650 (N_6650,N_5189,N_5906);
and U6651 (N_6651,N_5408,N_5435);
nor U6652 (N_6652,N_5613,N_5203);
and U6653 (N_6653,N_5015,N_5152);
or U6654 (N_6654,N_5365,N_5871);
or U6655 (N_6655,N_5333,N_5426);
nand U6656 (N_6656,N_5369,N_5236);
and U6657 (N_6657,N_5582,N_5024);
or U6658 (N_6658,N_5393,N_5193);
and U6659 (N_6659,N_5279,N_5624);
nor U6660 (N_6660,N_5412,N_5250);
xor U6661 (N_6661,N_5051,N_5445);
and U6662 (N_6662,N_5892,N_5244);
xor U6663 (N_6663,N_5325,N_5428);
and U6664 (N_6664,N_5662,N_5902);
or U6665 (N_6665,N_5288,N_5678);
and U6666 (N_6666,N_5394,N_5842);
or U6667 (N_6667,N_5528,N_5718);
and U6668 (N_6668,N_5527,N_5370);
nor U6669 (N_6669,N_5787,N_5445);
nor U6670 (N_6670,N_5616,N_5031);
and U6671 (N_6671,N_5260,N_5397);
nor U6672 (N_6672,N_5476,N_5203);
nor U6673 (N_6673,N_5002,N_5151);
nand U6674 (N_6674,N_5562,N_5106);
nor U6675 (N_6675,N_5734,N_5082);
or U6676 (N_6676,N_5246,N_5745);
or U6677 (N_6677,N_5482,N_5256);
nor U6678 (N_6678,N_5326,N_5775);
nor U6679 (N_6679,N_5513,N_5560);
and U6680 (N_6680,N_5558,N_5545);
or U6681 (N_6681,N_5087,N_5574);
nor U6682 (N_6682,N_5913,N_5620);
xor U6683 (N_6683,N_5009,N_5077);
and U6684 (N_6684,N_5684,N_5236);
and U6685 (N_6685,N_5592,N_5904);
nor U6686 (N_6686,N_5395,N_5164);
nor U6687 (N_6687,N_5862,N_5483);
xnor U6688 (N_6688,N_5694,N_5744);
and U6689 (N_6689,N_5994,N_5482);
and U6690 (N_6690,N_5461,N_5583);
and U6691 (N_6691,N_5339,N_5917);
xor U6692 (N_6692,N_5067,N_5497);
xnor U6693 (N_6693,N_5809,N_5156);
xor U6694 (N_6694,N_5126,N_5889);
nor U6695 (N_6695,N_5247,N_5549);
nand U6696 (N_6696,N_5041,N_5867);
xor U6697 (N_6697,N_5525,N_5921);
and U6698 (N_6698,N_5686,N_5655);
nand U6699 (N_6699,N_5151,N_5796);
nand U6700 (N_6700,N_5692,N_5108);
nand U6701 (N_6701,N_5879,N_5288);
xnor U6702 (N_6702,N_5442,N_5289);
nand U6703 (N_6703,N_5324,N_5658);
nor U6704 (N_6704,N_5703,N_5226);
nor U6705 (N_6705,N_5911,N_5776);
nand U6706 (N_6706,N_5159,N_5842);
or U6707 (N_6707,N_5606,N_5158);
and U6708 (N_6708,N_5793,N_5537);
or U6709 (N_6709,N_5451,N_5066);
and U6710 (N_6710,N_5161,N_5938);
nor U6711 (N_6711,N_5571,N_5612);
and U6712 (N_6712,N_5419,N_5410);
nand U6713 (N_6713,N_5259,N_5292);
nand U6714 (N_6714,N_5211,N_5225);
and U6715 (N_6715,N_5160,N_5844);
nor U6716 (N_6716,N_5132,N_5197);
nand U6717 (N_6717,N_5930,N_5891);
xor U6718 (N_6718,N_5370,N_5587);
or U6719 (N_6719,N_5528,N_5669);
and U6720 (N_6720,N_5473,N_5110);
nor U6721 (N_6721,N_5158,N_5773);
nor U6722 (N_6722,N_5468,N_5366);
nand U6723 (N_6723,N_5445,N_5092);
and U6724 (N_6724,N_5438,N_5112);
and U6725 (N_6725,N_5824,N_5150);
and U6726 (N_6726,N_5692,N_5990);
nand U6727 (N_6727,N_5010,N_5359);
and U6728 (N_6728,N_5137,N_5015);
or U6729 (N_6729,N_5490,N_5259);
and U6730 (N_6730,N_5790,N_5229);
and U6731 (N_6731,N_5459,N_5061);
nor U6732 (N_6732,N_5595,N_5215);
nor U6733 (N_6733,N_5197,N_5838);
and U6734 (N_6734,N_5832,N_5666);
and U6735 (N_6735,N_5521,N_5179);
or U6736 (N_6736,N_5543,N_5175);
nand U6737 (N_6737,N_5684,N_5549);
nand U6738 (N_6738,N_5401,N_5286);
or U6739 (N_6739,N_5617,N_5465);
nand U6740 (N_6740,N_5132,N_5551);
nand U6741 (N_6741,N_5318,N_5653);
xnor U6742 (N_6742,N_5193,N_5690);
nor U6743 (N_6743,N_5841,N_5863);
nand U6744 (N_6744,N_5802,N_5998);
or U6745 (N_6745,N_5571,N_5201);
nor U6746 (N_6746,N_5630,N_5884);
nand U6747 (N_6747,N_5312,N_5363);
xnor U6748 (N_6748,N_5685,N_5736);
nor U6749 (N_6749,N_5851,N_5971);
xnor U6750 (N_6750,N_5717,N_5283);
and U6751 (N_6751,N_5391,N_5853);
or U6752 (N_6752,N_5216,N_5802);
nand U6753 (N_6753,N_5600,N_5824);
xor U6754 (N_6754,N_5013,N_5489);
nor U6755 (N_6755,N_5453,N_5790);
nand U6756 (N_6756,N_5718,N_5180);
and U6757 (N_6757,N_5590,N_5433);
nor U6758 (N_6758,N_5396,N_5527);
nand U6759 (N_6759,N_5186,N_5259);
nor U6760 (N_6760,N_5222,N_5459);
and U6761 (N_6761,N_5336,N_5737);
or U6762 (N_6762,N_5684,N_5255);
nor U6763 (N_6763,N_5997,N_5397);
nand U6764 (N_6764,N_5875,N_5558);
or U6765 (N_6765,N_5882,N_5551);
nand U6766 (N_6766,N_5616,N_5301);
and U6767 (N_6767,N_5251,N_5270);
and U6768 (N_6768,N_5375,N_5037);
or U6769 (N_6769,N_5708,N_5488);
and U6770 (N_6770,N_5023,N_5590);
or U6771 (N_6771,N_5507,N_5801);
and U6772 (N_6772,N_5695,N_5998);
nand U6773 (N_6773,N_5321,N_5539);
and U6774 (N_6774,N_5959,N_5789);
nor U6775 (N_6775,N_5381,N_5031);
and U6776 (N_6776,N_5684,N_5027);
nor U6777 (N_6777,N_5381,N_5494);
and U6778 (N_6778,N_5738,N_5575);
nor U6779 (N_6779,N_5213,N_5543);
nor U6780 (N_6780,N_5536,N_5839);
or U6781 (N_6781,N_5357,N_5602);
and U6782 (N_6782,N_5599,N_5335);
nor U6783 (N_6783,N_5996,N_5299);
or U6784 (N_6784,N_5569,N_5994);
or U6785 (N_6785,N_5182,N_5043);
nor U6786 (N_6786,N_5827,N_5560);
nand U6787 (N_6787,N_5754,N_5929);
xnor U6788 (N_6788,N_5993,N_5536);
nor U6789 (N_6789,N_5995,N_5417);
and U6790 (N_6790,N_5719,N_5437);
or U6791 (N_6791,N_5199,N_5264);
nand U6792 (N_6792,N_5374,N_5326);
nand U6793 (N_6793,N_5328,N_5204);
nand U6794 (N_6794,N_5567,N_5497);
nand U6795 (N_6795,N_5115,N_5901);
and U6796 (N_6796,N_5771,N_5352);
nor U6797 (N_6797,N_5351,N_5285);
and U6798 (N_6798,N_5648,N_5426);
nand U6799 (N_6799,N_5676,N_5531);
and U6800 (N_6800,N_5674,N_5632);
and U6801 (N_6801,N_5877,N_5077);
or U6802 (N_6802,N_5082,N_5681);
nand U6803 (N_6803,N_5590,N_5307);
nor U6804 (N_6804,N_5520,N_5080);
and U6805 (N_6805,N_5231,N_5788);
or U6806 (N_6806,N_5353,N_5753);
nand U6807 (N_6807,N_5241,N_5505);
or U6808 (N_6808,N_5889,N_5587);
and U6809 (N_6809,N_5016,N_5563);
nor U6810 (N_6810,N_5018,N_5621);
nand U6811 (N_6811,N_5229,N_5258);
nand U6812 (N_6812,N_5796,N_5422);
and U6813 (N_6813,N_5536,N_5905);
and U6814 (N_6814,N_5167,N_5865);
xor U6815 (N_6815,N_5416,N_5364);
nand U6816 (N_6816,N_5237,N_5920);
xor U6817 (N_6817,N_5401,N_5342);
xor U6818 (N_6818,N_5447,N_5419);
and U6819 (N_6819,N_5044,N_5991);
and U6820 (N_6820,N_5422,N_5401);
or U6821 (N_6821,N_5894,N_5208);
nor U6822 (N_6822,N_5241,N_5948);
nor U6823 (N_6823,N_5853,N_5778);
nand U6824 (N_6824,N_5167,N_5308);
and U6825 (N_6825,N_5120,N_5449);
nor U6826 (N_6826,N_5988,N_5325);
nor U6827 (N_6827,N_5895,N_5520);
nand U6828 (N_6828,N_5499,N_5677);
nor U6829 (N_6829,N_5858,N_5908);
and U6830 (N_6830,N_5662,N_5660);
and U6831 (N_6831,N_5324,N_5013);
xor U6832 (N_6832,N_5809,N_5091);
and U6833 (N_6833,N_5873,N_5615);
and U6834 (N_6834,N_5270,N_5739);
or U6835 (N_6835,N_5754,N_5383);
nor U6836 (N_6836,N_5073,N_5493);
xnor U6837 (N_6837,N_5113,N_5170);
nor U6838 (N_6838,N_5015,N_5420);
nor U6839 (N_6839,N_5708,N_5521);
nor U6840 (N_6840,N_5214,N_5272);
nor U6841 (N_6841,N_5115,N_5890);
nand U6842 (N_6842,N_5042,N_5737);
nor U6843 (N_6843,N_5330,N_5946);
nor U6844 (N_6844,N_5224,N_5262);
and U6845 (N_6845,N_5726,N_5429);
nor U6846 (N_6846,N_5159,N_5615);
or U6847 (N_6847,N_5622,N_5207);
nand U6848 (N_6848,N_5186,N_5598);
and U6849 (N_6849,N_5285,N_5676);
or U6850 (N_6850,N_5924,N_5627);
nand U6851 (N_6851,N_5687,N_5594);
xnor U6852 (N_6852,N_5061,N_5027);
xor U6853 (N_6853,N_5468,N_5136);
and U6854 (N_6854,N_5917,N_5939);
and U6855 (N_6855,N_5437,N_5559);
xor U6856 (N_6856,N_5273,N_5104);
xnor U6857 (N_6857,N_5311,N_5957);
nor U6858 (N_6858,N_5819,N_5266);
nor U6859 (N_6859,N_5181,N_5878);
or U6860 (N_6860,N_5560,N_5372);
nor U6861 (N_6861,N_5233,N_5250);
and U6862 (N_6862,N_5416,N_5264);
nand U6863 (N_6863,N_5861,N_5727);
or U6864 (N_6864,N_5379,N_5173);
nor U6865 (N_6865,N_5806,N_5232);
nand U6866 (N_6866,N_5382,N_5643);
nor U6867 (N_6867,N_5492,N_5832);
and U6868 (N_6868,N_5946,N_5986);
nor U6869 (N_6869,N_5409,N_5485);
and U6870 (N_6870,N_5563,N_5195);
or U6871 (N_6871,N_5160,N_5465);
nand U6872 (N_6872,N_5738,N_5555);
nand U6873 (N_6873,N_5090,N_5813);
and U6874 (N_6874,N_5876,N_5225);
nand U6875 (N_6875,N_5722,N_5236);
nand U6876 (N_6876,N_5642,N_5909);
nand U6877 (N_6877,N_5041,N_5967);
nand U6878 (N_6878,N_5603,N_5438);
nor U6879 (N_6879,N_5137,N_5965);
or U6880 (N_6880,N_5557,N_5231);
nand U6881 (N_6881,N_5062,N_5830);
and U6882 (N_6882,N_5789,N_5322);
or U6883 (N_6883,N_5698,N_5415);
nand U6884 (N_6884,N_5503,N_5496);
nand U6885 (N_6885,N_5089,N_5696);
nor U6886 (N_6886,N_5743,N_5860);
or U6887 (N_6887,N_5649,N_5490);
nand U6888 (N_6888,N_5401,N_5692);
xnor U6889 (N_6889,N_5992,N_5808);
or U6890 (N_6890,N_5926,N_5999);
nor U6891 (N_6891,N_5330,N_5770);
and U6892 (N_6892,N_5767,N_5797);
nor U6893 (N_6893,N_5831,N_5013);
nand U6894 (N_6894,N_5085,N_5103);
and U6895 (N_6895,N_5281,N_5850);
and U6896 (N_6896,N_5238,N_5906);
nor U6897 (N_6897,N_5072,N_5991);
nand U6898 (N_6898,N_5047,N_5162);
and U6899 (N_6899,N_5928,N_5573);
nand U6900 (N_6900,N_5188,N_5619);
nand U6901 (N_6901,N_5483,N_5069);
nand U6902 (N_6902,N_5833,N_5294);
and U6903 (N_6903,N_5140,N_5784);
or U6904 (N_6904,N_5171,N_5007);
nand U6905 (N_6905,N_5556,N_5330);
nor U6906 (N_6906,N_5398,N_5426);
and U6907 (N_6907,N_5113,N_5674);
and U6908 (N_6908,N_5489,N_5380);
nor U6909 (N_6909,N_5972,N_5238);
and U6910 (N_6910,N_5290,N_5883);
and U6911 (N_6911,N_5291,N_5381);
nand U6912 (N_6912,N_5149,N_5702);
nor U6913 (N_6913,N_5178,N_5629);
and U6914 (N_6914,N_5697,N_5430);
nand U6915 (N_6915,N_5975,N_5988);
nor U6916 (N_6916,N_5501,N_5245);
nor U6917 (N_6917,N_5954,N_5522);
nor U6918 (N_6918,N_5233,N_5876);
nor U6919 (N_6919,N_5686,N_5812);
nand U6920 (N_6920,N_5475,N_5262);
nand U6921 (N_6921,N_5250,N_5871);
and U6922 (N_6922,N_5309,N_5498);
and U6923 (N_6923,N_5214,N_5930);
nand U6924 (N_6924,N_5023,N_5355);
nor U6925 (N_6925,N_5700,N_5488);
and U6926 (N_6926,N_5140,N_5616);
or U6927 (N_6927,N_5835,N_5034);
nor U6928 (N_6928,N_5109,N_5936);
nor U6929 (N_6929,N_5137,N_5222);
nor U6930 (N_6930,N_5696,N_5455);
nor U6931 (N_6931,N_5036,N_5823);
or U6932 (N_6932,N_5524,N_5123);
nor U6933 (N_6933,N_5317,N_5464);
or U6934 (N_6934,N_5562,N_5011);
nand U6935 (N_6935,N_5799,N_5576);
and U6936 (N_6936,N_5956,N_5756);
xnor U6937 (N_6937,N_5614,N_5101);
nor U6938 (N_6938,N_5907,N_5500);
nand U6939 (N_6939,N_5608,N_5147);
nand U6940 (N_6940,N_5684,N_5790);
xor U6941 (N_6941,N_5188,N_5825);
nand U6942 (N_6942,N_5571,N_5438);
or U6943 (N_6943,N_5170,N_5261);
xnor U6944 (N_6944,N_5446,N_5891);
nand U6945 (N_6945,N_5595,N_5287);
or U6946 (N_6946,N_5556,N_5042);
nor U6947 (N_6947,N_5565,N_5139);
nor U6948 (N_6948,N_5203,N_5325);
and U6949 (N_6949,N_5782,N_5851);
or U6950 (N_6950,N_5210,N_5257);
nand U6951 (N_6951,N_5550,N_5058);
nor U6952 (N_6952,N_5415,N_5217);
nand U6953 (N_6953,N_5691,N_5868);
or U6954 (N_6954,N_5049,N_5261);
or U6955 (N_6955,N_5065,N_5774);
or U6956 (N_6956,N_5154,N_5173);
nor U6957 (N_6957,N_5347,N_5394);
or U6958 (N_6958,N_5744,N_5239);
xnor U6959 (N_6959,N_5084,N_5998);
nand U6960 (N_6960,N_5420,N_5718);
or U6961 (N_6961,N_5894,N_5361);
nand U6962 (N_6962,N_5062,N_5561);
nor U6963 (N_6963,N_5891,N_5987);
nand U6964 (N_6964,N_5392,N_5721);
nor U6965 (N_6965,N_5399,N_5138);
nor U6966 (N_6966,N_5500,N_5190);
nand U6967 (N_6967,N_5898,N_5877);
nand U6968 (N_6968,N_5132,N_5422);
nand U6969 (N_6969,N_5824,N_5636);
xnor U6970 (N_6970,N_5380,N_5247);
and U6971 (N_6971,N_5422,N_5895);
xnor U6972 (N_6972,N_5116,N_5044);
nand U6973 (N_6973,N_5676,N_5624);
and U6974 (N_6974,N_5681,N_5034);
xor U6975 (N_6975,N_5094,N_5510);
nand U6976 (N_6976,N_5089,N_5629);
xor U6977 (N_6977,N_5888,N_5008);
or U6978 (N_6978,N_5824,N_5609);
and U6979 (N_6979,N_5559,N_5905);
or U6980 (N_6980,N_5187,N_5466);
nand U6981 (N_6981,N_5996,N_5831);
nor U6982 (N_6982,N_5963,N_5523);
nor U6983 (N_6983,N_5519,N_5669);
and U6984 (N_6984,N_5467,N_5268);
nor U6985 (N_6985,N_5525,N_5609);
nor U6986 (N_6986,N_5908,N_5817);
and U6987 (N_6987,N_5648,N_5817);
nand U6988 (N_6988,N_5521,N_5116);
and U6989 (N_6989,N_5654,N_5008);
or U6990 (N_6990,N_5548,N_5417);
nand U6991 (N_6991,N_5869,N_5962);
xor U6992 (N_6992,N_5861,N_5500);
nor U6993 (N_6993,N_5756,N_5460);
nor U6994 (N_6994,N_5260,N_5942);
or U6995 (N_6995,N_5203,N_5511);
and U6996 (N_6996,N_5271,N_5591);
nand U6997 (N_6997,N_5206,N_5749);
or U6998 (N_6998,N_5375,N_5268);
nand U6999 (N_6999,N_5576,N_5827);
nor U7000 (N_7000,N_6555,N_6194);
nor U7001 (N_7001,N_6997,N_6825);
or U7002 (N_7002,N_6607,N_6633);
nor U7003 (N_7003,N_6466,N_6850);
or U7004 (N_7004,N_6550,N_6819);
nor U7005 (N_7005,N_6108,N_6130);
nor U7006 (N_7006,N_6144,N_6580);
nor U7007 (N_7007,N_6849,N_6690);
nand U7008 (N_7008,N_6400,N_6349);
xnor U7009 (N_7009,N_6116,N_6360);
or U7010 (N_7010,N_6622,N_6013);
and U7011 (N_7011,N_6554,N_6595);
and U7012 (N_7012,N_6242,N_6733);
or U7013 (N_7013,N_6228,N_6642);
and U7014 (N_7014,N_6816,N_6402);
xor U7015 (N_7015,N_6931,N_6484);
nor U7016 (N_7016,N_6190,N_6851);
nor U7017 (N_7017,N_6756,N_6391);
xor U7018 (N_7018,N_6051,N_6004);
nor U7019 (N_7019,N_6372,N_6781);
nand U7020 (N_7020,N_6262,N_6741);
nand U7021 (N_7021,N_6202,N_6635);
nor U7022 (N_7022,N_6670,N_6937);
nor U7023 (N_7023,N_6582,N_6500);
and U7024 (N_7024,N_6193,N_6674);
or U7025 (N_7025,N_6615,N_6824);
or U7026 (N_7026,N_6886,N_6659);
or U7027 (N_7027,N_6857,N_6137);
nand U7028 (N_7028,N_6316,N_6697);
nor U7029 (N_7029,N_6176,N_6217);
xnor U7030 (N_7030,N_6169,N_6146);
and U7031 (N_7031,N_6513,N_6074);
nand U7032 (N_7032,N_6737,N_6258);
nand U7033 (N_7033,N_6195,N_6265);
nor U7034 (N_7034,N_6029,N_6090);
or U7035 (N_7035,N_6437,N_6044);
or U7036 (N_7036,N_6596,N_6359);
and U7037 (N_7037,N_6318,N_6460);
or U7038 (N_7038,N_6968,N_6821);
nor U7039 (N_7039,N_6061,N_6052);
nand U7040 (N_7040,N_6462,N_6842);
nor U7041 (N_7041,N_6150,N_6661);
nand U7042 (N_7042,N_6219,N_6124);
xnor U7043 (N_7043,N_6080,N_6143);
nand U7044 (N_7044,N_6406,N_6245);
xor U7045 (N_7045,N_6485,N_6673);
and U7046 (N_7046,N_6616,N_6012);
and U7047 (N_7047,N_6896,N_6155);
nand U7048 (N_7048,N_6758,N_6542);
xnor U7049 (N_7049,N_6643,N_6083);
nor U7050 (N_7050,N_6275,N_6474);
and U7051 (N_7051,N_6109,N_6114);
and U7052 (N_7052,N_6105,N_6742);
or U7053 (N_7053,N_6652,N_6605);
and U7054 (N_7054,N_6235,N_6000);
or U7055 (N_7055,N_6971,N_6617);
nor U7056 (N_7056,N_6656,N_6805);
or U7057 (N_7057,N_6984,N_6443);
xnor U7058 (N_7058,N_6632,N_6711);
xor U7059 (N_7059,N_6764,N_6367);
and U7060 (N_7060,N_6363,N_6919);
nand U7061 (N_7061,N_6895,N_6836);
nor U7062 (N_7062,N_6230,N_6151);
or U7063 (N_7063,N_6158,N_6054);
nor U7064 (N_7064,N_6645,N_6060);
nor U7065 (N_7065,N_6777,N_6592);
xor U7066 (N_7066,N_6410,N_6947);
nor U7067 (N_7067,N_6006,N_6983);
xor U7068 (N_7068,N_6153,N_6848);
and U7069 (N_7069,N_6878,N_6558);
xnor U7070 (N_7070,N_6695,N_6309);
or U7071 (N_7071,N_6820,N_6979);
and U7072 (N_7072,N_6089,N_6864);
nand U7073 (N_7073,N_6521,N_6148);
or U7074 (N_7074,N_6862,N_6476);
nand U7075 (N_7075,N_6099,N_6334);
nor U7076 (N_7076,N_6956,N_6749);
or U7077 (N_7077,N_6268,N_6882);
or U7078 (N_7078,N_6122,N_6998);
and U7079 (N_7079,N_6530,N_6488);
or U7080 (N_7080,N_6253,N_6822);
nand U7081 (N_7081,N_6952,N_6813);
and U7082 (N_7082,N_6017,N_6776);
or U7083 (N_7083,N_6573,N_6837);
nor U7084 (N_7084,N_6671,N_6240);
nor U7085 (N_7085,N_6694,N_6536);
nand U7086 (N_7086,N_6430,N_6803);
nand U7087 (N_7087,N_6755,N_6375);
and U7088 (N_7088,N_6570,N_6250);
or U7089 (N_7089,N_6270,N_6233);
nor U7090 (N_7090,N_6691,N_6753);
and U7091 (N_7091,N_6067,N_6765);
or U7092 (N_7092,N_6724,N_6746);
or U7093 (N_7093,N_6221,N_6809);
and U7094 (N_7094,N_6967,N_6501);
and U7095 (N_7095,N_6175,N_6823);
or U7096 (N_7096,N_6593,N_6413);
and U7097 (N_7097,N_6728,N_6881);
or U7098 (N_7098,N_6818,N_6496);
or U7099 (N_7099,N_6440,N_6664);
xnor U7100 (N_7100,N_6037,N_6342);
nor U7101 (N_7101,N_6871,N_6296);
nor U7102 (N_7102,N_6668,N_6735);
and U7103 (N_7103,N_6658,N_6913);
xor U7104 (N_7104,N_6393,N_6731);
and U7105 (N_7105,N_6395,N_6002);
or U7106 (N_7106,N_6241,N_6970);
nand U7107 (N_7107,N_6608,N_6348);
or U7108 (N_7108,N_6503,N_6401);
and U7109 (N_7109,N_6154,N_6302);
or U7110 (N_7110,N_6743,N_6778);
nor U7111 (N_7111,N_6291,N_6933);
nand U7112 (N_7112,N_6586,N_6773);
nor U7113 (N_7113,N_6720,N_6900);
and U7114 (N_7114,N_6251,N_6768);
nand U7115 (N_7115,N_6034,N_6444);
nand U7116 (N_7116,N_6185,N_6843);
nor U7117 (N_7117,N_6222,N_6508);
nand U7118 (N_7118,N_6775,N_6954);
and U7119 (N_7119,N_6799,N_6252);
and U7120 (N_7120,N_6304,N_6800);
or U7121 (N_7121,N_6057,N_6201);
xor U7122 (N_7122,N_6610,N_6650);
xor U7123 (N_7123,N_6127,N_6058);
or U7124 (N_7124,N_6714,N_6392);
nor U7125 (N_7125,N_6133,N_6667);
nor U7126 (N_7126,N_6449,N_6928);
or U7127 (N_7127,N_6338,N_6976);
nor U7128 (N_7128,N_6161,N_6293);
nor U7129 (N_7129,N_6020,N_6512);
nand U7130 (N_7130,N_6894,N_6552);
nor U7131 (N_7131,N_6079,N_6834);
nor U7132 (N_7132,N_6023,N_6914);
or U7133 (N_7133,N_6386,N_6638);
nand U7134 (N_7134,N_6523,N_6789);
and U7135 (N_7135,N_6906,N_6428);
nor U7136 (N_7136,N_6620,N_6340);
or U7137 (N_7137,N_6792,N_6634);
or U7138 (N_7138,N_6289,N_6015);
nor U7139 (N_7139,N_6588,N_6166);
and U7140 (N_7140,N_6766,N_6149);
nand U7141 (N_7141,N_6011,N_6647);
nand U7142 (N_7142,N_6483,N_6688);
xor U7143 (N_7143,N_6021,N_6292);
nor U7144 (N_7144,N_6300,N_6666);
xnor U7145 (N_7145,N_6996,N_6055);
and U7146 (N_7146,N_6008,N_6978);
or U7147 (N_7147,N_6517,N_6341);
nand U7148 (N_7148,N_6625,N_6899);
or U7149 (N_7149,N_6653,N_6738);
nor U7150 (N_7150,N_6925,N_6793);
or U7151 (N_7151,N_6452,N_6326);
or U7152 (N_7152,N_6702,N_6641);
nand U7153 (N_7153,N_6467,N_6762);
nand U7154 (N_7154,N_6703,N_6085);
and U7155 (N_7155,N_6721,N_6510);
or U7156 (N_7156,N_6352,N_6473);
nor U7157 (N_7157,N_6128,N_6716);
nor U7158 (N_7158,N_6432,N_6243);
or U7159 (N_7159,N_6328,N_6854);
nand U7160 (N_7160,N_6421,N_6584);
nand U7161 (N_7161,N_6880,N_6319);
and U7162 (N_7162,N_6237,N_6490);
nor U7163 (N_7163,N_6889,N_6547);
and U7164 (N_7164,N_6959,N_6752);
or U7165 (N_7165,N_6147,N_6431);
or U7166 (N_7166,N_6434,N_6929);
or U7167 (N_7167,N_6684,N_6170);
or U7168 (N_7168,N_6229,N_6179);
and U7169 (N_7169,N_6331,N_6827);
or U7170 (N_7170,N_6212,N_6323);
nand U7171 (N_7171,N_6718,N_6639);
nand U7172 (N_7172,N_6110,N_6298);
nand U7173 (N_7173,N_6208,N_6748);
nor U7174 (N_7174,N_6927,N_6187);
and U7175 (N_7175,N_6747,N_6022);
and U7176 (N_7176,N_6203,N_6942);
nand U7177 (N_7177,N_6327,N_6140);
and U7178 (N_7178,N_6086,N_6374);
nor U7179 (N_7179,N_6009,N_6081);
and U7180 (N_7180,N_6723,N_6760);
nor U7181 (N_7181,N_6516,N_6415);
nor U7182 (N_7182,N_6409,N_6761);
and U7183 (N_7183,N_6692,N_6568);
or U7184 (N_7184,N_6569,N_6985);
or U7185 (N_7185,N_6199,N_6627);
nor U7186 (N_7186,N_6729,N_6172);
nor U7187 (N_7187,N_6091,N_6590);
nand U7188 (N_7188,N_6311,N_6301);
nand U7189 (N_7189,N_6279,N_6047);
or U7190 (N_7190,N_6031,N_6288);
nor U7191 (N_7191,N_6908,N_6059);
and U7192 (N_7192,N_6946,N_6307);
and U7193 (N_7193,N_6427,N_6003);
and U7194 (N_7194,N_6405,N_6356);
nand U7195 (N_7195,N_6975,N_6637);
nand U7196 (N_7196,N_6280,N_6982);
nor U7197 (N_7197,N_6907,N_6884);
xnor U7198 (N_7198,N_6024,N_6377);
or U7199 (N_7199,N_6494,N_6062);
or U7200 (N_7200,N_6990,N_6248);
nor U7201 (N_7201,N_6887,N_6142);
xnor U7202 (N_7202,N_6365,N_6010);
and U7203 (N_7203,N_6551,N_6068);
nor U7204 (N_7204,N_6225,N_6489);
or U7205 (N_7205,N_6274,N_6699);
xor U7206 (N_7206,N_6897,N_6845);
nand U7207 (N_7207,N_6657,N_6713);
or U7208 (N_7208,N_6538,N_6422);
nand U7209 (N_7209,N_6041,N_6308);
nand U7210 (N_7210,N_6770,N_6621);
nor U7211 (N_7211,N_6868,N_6254);
or U7212 (N_7212,N_6838,N_6438);
nand U7213 (N_7213,N_6585,N_6103);
or U7214 (N_7214,N_6999,N_6577);
nor U7215 (N_7215,N_6672,N_6345);
nor U7216 (N_7216,N_6373,N_6915);
nor U7217 (N_7217,N_6120,N_6772);
nand U7218 (N_7218,N_6705,N_6314);
or U7219 (N_7219,N_6710,N_6532);
xnor U7220 (N_7220,N_6704,N_6094);
or U7221 (N_7221,N_6941,N_6325);
and U7222 (N_7222,N_6157,N_6491);
nand U7223 (N_7223,N_6507,N_6918);
nand U7224 (N_7224,N_6994,N_6101);
nor U7225 (N_7225,N_6665,N_6788);
nand U7226 (N_7226,N_6313,N_6763);
xnor U7227 (N_7227,N_6812,N_6287);
nor U7228 (N_7228,N_6972,N_6877);
or U7229 (N_7229,N_6576,N_6830);
or U7230 (N_7230,N_6113,N_6425);
and U7231 (N_7231,N_6197,N_6414);
and U7232 (N_7232,N_6016,N_6981);
nor U7233 (N_7233,N_6324,N_6563);
nand U7234 (N_7234,N_6992,N_6932);
and U7235 (N_7235,N_6064,N_6571);
or U7236 (N_7236,N_6701,N_6549);
and U7237 (N_7237,N_6249,N_6644);
or U7238 (N_7238,N_6888,N_6506);
nand U7239 (N_7239,N_6403,N_6599);
and U7240 (N_7240,N_6329,N_6798);
nor U7241 (N_7241,N_6231,N_6548);
and U7242 (N_7242,N_6511,N_6767);
nand U7243 (N_7243,N_6682,N_6239);
nor U7244 (N_7244,N_6935,N_6260);
nand U7245 (N_7245,N_6346,N_6870);
nor U7246 (N_7246,N_6531,N_6750);
and U7247 (N_7247,N_6030,N_6278);
nand U7248 (N_7248,N_6626,N_6567);
xor U7249 (N_7249,N_6852,N_6285);
and U7250 (N_7250,N_6910,N_6174);
and U7251 (N_7251,N_6078,N_6457);
and U7252 (N_7252,N_6214,N_6387);
and U7253 (N_7253,N_6236,N_6361);
nand U7254 (N_7254,N_6336,N_6383);
nand U7255 (N_7255,N_6829,N_6192);
nand U7256 (N_7256,N_6924,N_6802);
or U7257 (N_7257,N_6299,N_6435);
and U7258 (N_7258,N_6290,N_6305);
xor U7259 (N_7259,N_6930,N_6223);
and U7260 (N_7260,N_6358,N_6537);
and U7261 (N_7261,N_6541,N_6869);
nand U7262 (N_7262,N_6459,N_6875);
or U7263 (N_7263,N_6038,N_6722);
nand U7264 (N_7264,N_6053,N_6337);
and U7265 (N_7265,N_6602,N_6132);
xnor U7266 (N_7266,N_6196,N_6418);
nor U7267 (N_7267,N_6589,N_6339);
and U7268 (N_7268,N_6712,N_6417);
nor U7269 (N_7269,N_6993,N_6272);
and U7270 (N_7270,N_6559,N_6732);
and U7271 (N_7271,N_6923,N_6479);
and U7272 (N_7272,N_6049,N_6583);
and U7273 (N_7273,N_6495,N_6446);
or U7274 (N_7274,N_6465,N_6315);
nand U7275 (N_7275,N_6651,N_6603);
nand U7276 (N_7276,N_6261,N_6715);
nor U7277 (N_7277,N_6893,N_6892);
nand U7278 (N_7278,N_6436,N_6575);
and U7279 (N_7279,N_6458,N_6412);
nand U7280 (N_7280,N_6283,N_6546);
nor U7281 (N_7281,N_6594,N_6681);
or U7282 (N_7282,N_6902,N_6696);
and U7283 (N_7283,N_6679,N_6138);
and U7284 (N_7284,N_6126,N_6087);
nand U7285 (N_7285,N_6963,N_6045);
or U7286 (N_7286,N_6282,N_6926);
or U7287 (N_7287,N_6032,N_6654);
nand U7288 (N_7288,N_6384,N_6450);
and U7289 (N_7289,N_6419,N_6950);
nand U7290 (N_7290,N_6744,N_6680);
nand U7291 (N_7291,N_6519,N_6844);
nand U7292 (N_7292,N_6007,N_6487);
and U7293 (N_7293,N_6039,N_6831);
nor U7294 (N_7294,N_6662,N_6543);
nand U7295 (N_7295,N_6791,N_6481);
nor U7296 (N_7296,N_6591,N_6163);
nor U7297 (N_7297,N_6276,N_6164);
and U7298 (N_7298,N_6046,N_6376);
xor U7299 (N_7299,N_6553,N_6957);
nor U7300 (N_7300,N_6439,N_6227);
nand U7301 (N_7301,N_6303,N_6183);
nor U7302 (N_7302,N_6306,N_6669);
or U7303 (N_7303,N_6475,N_6189);
and U7304 (N_7304,N_6574,N_6477);
nand U7305 (N_7305,N_6612,N_6787);
nand U7306 (N_7306,N_6611,N_6226);
xor U7307 (N_7307,N_6097,N_6948);
nor U7308 (N_7308,N_6587,N_6390);
and U7309 (N_7309,N_6357,N_6790);
nor U7310 (N_7310,N_6423,N_6808);
or U7311 (N_7311,N_6456,N_6973);
and U7312 (N_7312,N_6040,N_6861);
and U7313 (N_7313,N_6118,N_6560);
nand U7314 (N_7314,N_6911,N_6026);
nor U7315 (N_7315,N_6294,N_6332);
or U7316 (N_7316,N_6152,N_6297);
nor U7317 (N_7317,N_6841,N_6561);
nand U7318 (N_7318,N_6522,N_6786);
and U7319 (N_7319,N_6050,N_6186);
and U7320 (N_7320,N_6991,N_6131);
or U7321 (N_7321,N_6271,N_6112);
nand U7322 (N_7322,N_6833,N_6033);
nor U7323 (N_7323,N_6480,N_6092);
and U7324 (N_7324,N_6213,N_6404);
nor U7325 (N_7325,N_6156,N_6578);
or U7326 (N_7326,N_6826,N_6876);
and U7327 (N_7327,N_6613,N_6408);
and U7328 (N_7328,N_6106,N_6663);
nand U7329 (N_7329,N_6598,N_6835);
nand U7330 (N_7330,N_6920,N_6277);
or U7331 (N_7331,N_6872,N_6453);
and U7332 (N_7332,N_6362,N_6234);
nor U7333 (N_7333,N_6115,N_6505);
xor U7334 (N_7334,N_6267,N_6125);
or U7335 (N_7335,N_6069,N_6579);
nor U7336 (N_7336,N_6839,N_6028);
or U7337 (N_7337,N_6111,N_6018);
or U7338 (N_7338,N_6840,N_6366);
nand U7339 (N_7339,N_6461,N_6977);
nor U7340 (N_7340,N_6618,N_6389);
and U7341 (N_7341,N_6557,N_6205);
nand U7342 (N_7342,N_6454,N_6220);
nor U7343 (N_7343,N_6980,N_6725);
xnor U7344 (N_7344,N_6953,N_6853);
nand U7345 (N_7345,N_6098,N_6520);
or U7346 (N_7346,N_6545,N_6354);
nand U7347 (N_7347,N_6939,N_6206);
or U7348 (N_7348,N_6534,N_6685);
nor U7349 (N_7349,N_6076,N_6266);
and U7350 (N_7350,N_6198,N_6614);
nand U7351 (N_7351,N_6660,N_6909);
nor U7352 (N_7352,N_6916,N_6879);
nand U7353 (N_7353,N_6257,N_6121);
nand U7354 (N_7354,N_6426,N_6343);
and U7355 (N_7355,N_6082,N_6141);
or U7356 (N_7356,N_6965,N_6535);
and U7357 (N_7357,N_6486,N_6420);
xnor U7358 (N_7358,N_6273,N_6075);
nand U7359 (N_7359,N_6102,N_6188);
nor U7360 (N_7360,N_6215,N_6182);
and U7361 (N_7361,N_6247,N_6649);
or U7362 (N_7362,N_6264,N_6027);
and U7363 (N_7363,N_6811,N_6167);
or U7364 (N_7364,N_6529,N_6917);
nor U7365 (N_7365,N_6025,N_6416);
xor U7366 (N_7366,N_6785,N_6646);
nand U7367 (N_7367,N_6232,N_6177);
and U7368 (N_7368,N_6539,N_6771);
nor U7369 (N_7369,N_6631,N_6441);
nand U7370 (N_7370,N_6863,N_6335);
nor U7371 (N_7371,N_6514,N_6001);
nor U7372 (N_7372,N_6369,N_6810);
or U7373 (N_7373,N_6019,N_6989);
and U7374 (N_7374,N_6938,N_6779);
or U7375 (N_7375,N_6606,N_6609);
and U7376 (N_7376,N_6333,N_6399);
nor U7377 (N_7377,N_6209,N_6726);
or U7378 (N_7378,N_6502,N_6165);
nand U7379 (N_7379,N_6683,N_6944);
nor U7380 (N_7380,N_6686,N_6655);
nand U7381 (N_7381,N_6904,N_6244);
xnor U7382 (N_7382,N_6388,N_6256);
nand U7383 (N_7383,N_6740,N_6964);
nand U7384 (N_7384,N_6949,N_6093);
nor U7385 (N_7385,N_6936,N_6556);
nor U7386 (N_7386,N_6084,N_6312);
or U7387 (N_7387,N_6524,N_6730);
and U7388 (N_7388,N_6322,N_6499);
nand U7389 (N_7389,N_6969,N_6424);
nand U7390 (N_7390,N_6200,N_6509);
or U7391 (N_7391,N_6463,N_6317);
or U7392 (N_7392,N_6096,N_6648);
xor U7393 (N_7393,N_6210,N_6447);
or U7394 (N_7394,N_6544,N_6736);
or U7395 (N_7395,N_6675,N_6347);
xnor U7396 (N_7396,N_6478,N_6689);
nand U7397 (N_7397,N_6448,N_6619);
nor U7398 (N_7398,N_6707,N_6504);
and U7399 (N_7399,N_6471,N_6727);
nand U7400 (N_7400,N_6350,N_6498);
and U7401 (N_7401,N_6564,N_6987);
nand U7402 (N_7402,N_6072,N_6940);
or U7403 (N_7403,N_6005,N_6071);
and U7404 (N_7404,N_6890,N_6482);
and U7405 (N_7405,N_6739,N_6378);
and U7406 (N_7406,N_6717,N_6636);
nor U7407 (N_7407,N_6706,N_6988);
xnor U7408 (N_7408,N_6445,N_6429);
and U7409 (N_7409,N_6769,N_6100);
and U7410 (N_7410,N_6135,N_6922);
xnor U7411 (N_7411,N_6381,N_6451);
nand U7412 (N_7412,N_6180,N_6397);
or U7413 (N_7413,N_6754,N_6065);
or U7414 (N_7414,N_6411,N_6497);
nand U7415 (N_7415,N_6310,N_6396);
nand U7416 (N_7416,N_6832,N_6119);
nand U7417 (N_7417,N_6986,N_6604);
or U7418 (N_7418,N_6533,N_6263);
nand U7419 (N_7419,N_6943,N_6796);
nand U7420 (N_7420,N_6814,N_6070);
and U7421 (N_7421,N_6469,N_6709);
or U7422 (N_7422,N_6794,N_6597);
and U7423 (N_7423,N_6353,N_6912);
or U7424 (N_7424,N_6751,N_6623);
or U7425 (N_7425,N_6145,N_6160);
or U7426 (N_7426,N_6995,N_6398);
and U7427 (N_7427,N_6104,N_6281);
xnor U7428 (N_7428,N_6966,N_6470);
or U7429 (N_7429,N_6958,N_6382);
or U7430 (N_7430,N_6073,N_6173);
nand U7431 (N_7431,N_6204,N_6846);
nand U7432 (N_7432,N_6066,N_6783);
and U7433 (N_7433,N_6368,N_6858);
nand U7434 (N_7434,N_6181,N_6693);
nor U7435 (N_7435,N_6745,N_6216);
nand U7436 (N_7436,N_6734,N_6117);
nor U7437 (N_7437,N_6259,N_6286);
and U7438 (N_7438,N_6159,N_6860);
xor U7439 (N_7439,N_6905,N_6171);
nor U7440 (N_7440,N_6370,N_6921);
nand U7441 (N_7441,N_6866,N_6883);
nor U7442 (N_7442,N_6708,N_6628);
nor U7443 (N_7443,N_6218,N_6640);
and U7444 (N_7444,N_6063,N_6806);
or U7445 (N_7445,N_6255,N_6136);
nor U7446 (N_7446,N_6807,N_6036);
and U7447 (N_7447,N_6847,N_6855);
or U7448 (N_7448,N_6077,N_6817);
or U7449 (N_7449,N_6238,N_6795);
or U7450 (N_7450,N_6043,N_6364);
and U7451 (N_7451,N_6385,N_6295);
or U7452 (N_7452,N_6867,N_6859);
xor U7453 (N_7453,N_6442,N_6934);
nor U7454 (N_7454,N_6951,N_6962);
and U7455 (N_7455,N_6472,N_6492);
or U7456 (N_7456,N_6246,N_6759);
nor U7457 (N_7457,N_6874,N_6527);
and U7458 (N_7458,N_6945,N_6168);
or U7459 (N_7459,N_6873,N_6107);
and U7460 (N_7460,N_6455,N_6518);
and U7461 (N_7461,N_6464,N_6774);
nor U7462 (N_7462,N_6581,N_6433);
nor U7463 (N_7463,N_6139,N_6528);
nand U7464 (N_7464,N_6629,N_6901);
nand U7465 (N_7465,N_6284,N_6630);
nand U7466 (N_7466,N_6042,N_6572);
and U7467 (N_7467,N_6525,N_6678);
and U7468 (N_7468,N_6379,N_6700);
nand U7469 (N_7469,N_6355,N_6468);
nor U7470 (N_7470,N_6207,N_6955);
nand U7471 (N_7471,N_6601,N_6757);
nand U7472 (N_7472,N_6088,N_6123);
nand U7473 (N_7473,N_6960,N_6269);
and U7474 (N_7474,N_6780,N_6565);
nand U7475 (N_7475,N_6891,N_6698);
nor U7476 (N_7476,N_6394,N_6540);
or U7477 (N_7477,N_6865,N_6885);
or U7478 (N_7478,N_6380,N_6961);
nand U7479 (N_7479,N_6191,N_6797);
nand U7480 (N_7480,N_6224,N_6035);
nor U7481 (N_7481,N_6048,N_6493);
or U7482 (N_7482,N_6095,N_6624);
nand U7483 (N_7483,N_6211,N_6014);
nand U7484 (N_7484,N_6321,N_6526);
or U7485 (N_7485,N_6184,N_6178);
nor U7486 (N_7486,N_6562,N_6719);
nand U7487 (N_7487,N_6566,N_6515);
xnor U7488 (N_7488,N_6782,N_6677);
nor U7489 (N_7489,N_6407,N_6898);
nor U7490 (N_7490,N_6320,N_6828);
or U7491 (N_7491,N_6804,N_6600);
and U7492 (N_7492,N_6815,N_6371);
nor U7493 (N_7493,N_6676,N_6351);
xor U7494 (N_7494,N_6784,N_6330);
nor U7495 (N_7495,N_6344,N_6687);
nand U7496 (N_7496,N_6056,N_6134);
or U7497 (N_7497,N_6801,N_6903);
xnor U7498 (N_7498,N_6162,N_6129);
or U7499 (N_7499,N_6974,N_6856);
nand U7500 (N_7500,N_6931,N_6336);
nand U7501 (N_7501,N_6304,N_6097);
nor U7502 (N_7502,N_6411,N_6455);
and U7503 (N_7503,N_6738,N_6655);
nand U7504 (N_7504,N_6736,N_6959);
and U7505 (N_7505,N_6948,N_6135);
or U7506 (N_7506,N_6510,N_6228);
and U7507 (N_7507,N_6398,N_6545);
or U7508 (N_7508,N_6302,N_6784);
nand U7509 (N_7509,N_6888,N_6826);
nand U7510 (N_7510,N_6017,N_6111);
and U7511 (N_7511,N_6952,N_6343);
nand U7512 (N_7512,N_6071,N_6179);
and U7513 (N_7513,N_6068,N_6770);
or U7514 (N_7514,N_6920,N_6763);
or U7515 (N_7515,N_6522,N_6910);
or U7516 (N_7516,N_6155,N_6885);
xor U7517 (N_7517,N_6130,N_6895);
or U7518 (N_7518,N_6972,N_6553);
and U7519 (N_7519,N_6246,N_6109);
xor U7520 (N_7520,N_6847,N_6743);
and U7521 (N_7521,N_6489,N_6505);
xor U7522 (N_7522,N_6175,N_6830);
and U7523 (N_7523,N_6424,N_6200);
xor U7524 (N_7524,N_6716,N_6075);
nand U7525 (N_7525,N_6361,N_6624);
nor U7526 (N_7526,N_6137,N_6584);
or U7527 (N_7527,N_6920,N_6598);
and U7528 (N_7528,N_6298,N_6041);
or U7529 (N_7529,N_6979,N_6520);
or U7530 (N_7530,N_6940,N_6526);
or U7531 (N_7531,N_6646,N_6400);
and U7532 (N_7532,N_6688,N_6196);
and U7533 (N_7533,N_6577,N_6350);
and U7534 (N_7534,N_6549,N_6643);
nor U7535 (N_7535,N_6642,N_6672);
nand U7536 (N_7536,N_6465,N_6709);
nor U7537 (N_7537,N_6937,N_6791);
nand U7538 (N_7538,N_6882,N_6508);
or U7539 (N_7539,N_6150,N_6372);
nor U7540 (N_7540,N_6219,N_6658);
and U7541 (N_7541,N_6911,N_6355);
and U7542 (N_7542,N_6124,N_6305);
or U7543 (N_7543,N_6015,N_6184);
nand U7544 (N_7544,N_6599,N_6690);
or U7545 (N_7545,N_6091,N_6451);
nand U7546 (N_7546,N_6945,N_6026);
and U7547 (N_7547,N_6823,N_6898);
nand U7548 (N_7548,N_6927,N_6532);
nand U7549 (N_7549,N_6319,N_6264);
nor U7550 (N_7550,N_6343,N_6604);
nor U7551 (N_7551,N_6217,N_6572);
or U7552 (N_7552,N_6709,N_6380);
and U7553 (N_7553,N_6855,N_6761);
nor U7554 (N_7554,N_6591,N_6201);
nand U7555 (N_7555,N_6005,N_6377);
nand U7556 (N_7556,N_6606,N_6186);
nor U7557 (N_7557,N_6162,N_6395);
nand U7558 (N_7558,N_6310,N_6731);
xnor U7559 (N_7559,N_6274,N_6120);
nand U7560 (N_7560,N_6672,N_6150);
nand U7561 (N_7561,N_6353,N_6218);
and U7562 (N_7562,N_6637,N_6869);
or U7563 (N_7563,N_6148,N_6633);
nand U7564 (N_7564,N_6216,N_6241);
and U7565 (N_7565,N_6155,N_6645);
and U7566 (N_7566,N_6266,N_6710);
nor U7567 (N_7567,N_6842,N_6473);
xor U7568 (N_7568,N_6219,N_6359);
and U7569 (N_7569,N_6963,N_6485);
xnor U7570 (N_7570,N_6496,N_6522);
or U7571 (N_7571,N_6679,N_6185);
and U7572 (N_7572,N_6808,N_6524);
nand U7573 (N_7573,N_6374,N_6358);
nand U7574 (N_7574,N_6615,N_6280);
nor U7575 (N_7575,N_6463,N_6740);
or U7576 (N_7576,N_6859,N_6616);
nand U7577 (N_7577,N_6960,N_6501);
and U7578 (N_7578,N_6462,N_6472);
nand U7579 (N_7579,N_6400,N_6923);
nand U7580 (N_7580,N_6041,N_6979);
and U7581 (N_7581,N_6342,N_6878);
xnor U7582 (N_7582,N_6549,N_6490);
or U7583 (N_7583,N_6598,N_6063);
or U7584 (N_7584,N_6974,N_6729);
or U7585 (N_7585,N_6310,N_6531);
or U7586 (N_7586,N_6896,N_6494);
or U7587 (N_7587,N_6002,N_6473);
nand U7588 (N_7588,N_6098,N_6530);
nand U7589 (N_7589,N_6741,N_6278);
nand U7590 (N_7590,N_6165,N_6350);
and U7591 (N_7591,N_6960,N_6421);
nor U7592 (N_7592,N_6206,N_6720);
or U7593 (N_7593,N_6991,N_6320);
or U7594 (N_7594,N_6190,N_6848);
or U7595 (N_7595,N_6472,N_6920);
and U7596 (N_7596,N_6609,N_6061);
and U7597 (N_7597,N_6242,N_6011);
nor U7598 (N_7598,N_6341,N_6519);
nand U7599 (N_7599,N_6302,N_6726);
nor U7600 (N_7600,N_6089,N_6484);
or U7601 (N_7601,N_6363,N_6725);
nand U7602 (N_7602,N_6106,N_6728);
or U7603 (N_7603,N_6150,N_6570);
xor U7604 (N_7604,N_6198,N_6336);
xnor U7605 (N_7605,N_6772,N_6785);
or U7606 (N_7606,N_6213,N_6672);
xor U7607 (N_7607,N_6818,N_6552);
nor U7608 (N_7608,N_6077,N_6095);
and U7609 (N_7609,N_6555,N_6138);
xnor U7610 (N_7610,N_6703,N_6255);
nor U7611 (N_7611,N_6386,N_6565);
or U7612 (N_7612,N_6778,N_6260);
or U7613 (N_7613,N_6946,N_6434);
xnor U7614 (N_7614,N_6928,N_6494);
nand U7615 (N_7615,N_6988,N_6469);
xnor U7616 (N_7616,N_6294,N_6711);
and U7617 (N_7617,N_6173,N_6457);
and U7618 (N_7618,N_6369,N_6397);
nor U7619 (N_7619,N_6260,N_6424);
nand U7620 (N_7620,N_6241,N_6675);
nand U7621 (N_7621,N_6503,N_6565);
xnor U7622 (N_7622,N_6605,N_6472);
or U7623 (N_7623,N_6494,N_6297);
nand U7624 (N_7624,N_6860,N_6740);
nand U7625 (N_7625,N_6185,N_6624);
xnor U7626 (N_7626,N_6970,N_6406);
nand U7627 (N_7627,N_6924,N_6923);
and U7628 (N_7628,N_6788,N_6845);
nand U7629 (N_7629,N_6309,N_6605);
nor U7630 (N_7630,N_6740,N_6542);
and U7631 (N_7631,N_6250,N_6196);
and U7632 (N_7632,N_6648,N_6612);
or U7633 (N_7633,N_6086,N_6929);
or U7634 (N_7634,N_6916,N_6061);
or U7635 (N_7635,N_6885,N_6782);
and U7636 (N_7636,N_6439,N_6482);
nand U7637 (N_7637,N_6062,N_6947);
nand U7638 (N_7638,N_6370,N_6013);
and U7639 (N_7639,N_6380,N_6482);
and U7640 (N_7640,N_6799,N_6265);
nand U7641 (N_7641,N_6546,N_6354);
nor U7642 (N_7642,N_6912,N_6360);
nand U7643 (N_7643,N_6729,N_6900);
nor U7644 (N_7644,N_6972,N_6063);
and U7645 (N_7645,N_6108,N_6730);
or U7646 (N_7646,N_6796,N_6767);
nand U7647 (N_7647,N_6033,N_6989);
or U7648 (N_7648,N_6692,N_6854);
or U7649 (N_7649,N_6837,N_6245);
nand U7650 (N_7650,N_6615,N_6943);
and U7651 (N_7651,N_6319,N_6886);
or U7652 (N_7652,N_6724,N_6681);
nor U7653 (N_7653,N_6689,N_6429);
and U7654 (N_7654,N_6189,N_6226);
xnor U7655 (N_7655,N_6318,N_6062);
or U7656 (N_7656,N_6715,N_6807);
and U7657 (N_7657,N_6007,N_6950);
or U7658 (N_7658,N_6755,N_6769);
nor U7659 (N_7659,N_6512,N_6573);
nor U7660 (N_7660,N_6331,N_6617);
or U7661 (N_7661,N_6605,N_6008);
or U7662 (N_7662,N_6369,N_6691);
and U7663 (N_7663,N_6988,N_6897);
and U7664 (N_7664,N_6415,N_6234);
and U7665 (N_7665,N_6524,N_6476);
and U7666 (N_7666,N_6926,N_6567);
nand U7667 (N_7667,N_6330,N_6056);
xor U7668 (N_7668,N_6846,N_6956);
nand U7669 (N_7669,N_6989,N_6603);
nor U7670 (N_7670,N_6315,N_6852);
nor U7671 (N_7671,N_6009,N_6962);
and U7672 (N_7672,N_6893,N_6122);
or U7673 (N_7673,N_6570,N_6343);
nor U7674 (N_7674,N_6562,N_6994);
nand U7675 (N_7675,N_6523,N_6938);
xor U7676 (N_7676,N_6900,N_6533);
or U7677 (N_7677,N_6968,N_6970);
nor U7678 (N_7678,N_6360,N_6692);
or U7679 (N_7679,N_6992,N_6221);
and U7680 (N_7680,N_6419,N_6148);
nand U7681 (N_7681,N_6121,N_6710);
nand U7682 (N_7682,N_6007,N_6662);
and U7683 (N_7683,N_6221,N_6452);
or U7684 (N_7684,N_6866,N_6935);
or U7685 (N_7685,N_6827,N_6581);
and U7686 (N_7686,N_6016,N_6446);
and U7687 (N_7687,N_6062,N_6249);
nand U7688 (N_7688,N_6750,N_6087);
nor U7689 (N_7689,N_6190,N_6527);
or U7690 (N_7690,N_6519,N_6895);
nand U7691 (N_7691,N_6099,N_6184);
and U7692 (N_7692,N_6902,N_6962);
nand U7693 (N_7693,N_6129,N_6690);
and U7694 (N_7694,N_6147,N_6481);
or U7695 (N_7695,N_6273,N_6913);
or U7696 (N_7696,N_6989,N_6847);
and U7697 (N_7697,N_6233,N_6908);
or U7698 (N_7698,N_6283,N_6121);
or U7699 (N_7699,N_6648,N_6008);
or U7700 (N_7700,N_6201,N_6536);
or U7701 (N_7701,N_6162,N_6088);
nor U7702 (N_7702,N_6516,N_6736);
or U7703 (N_7703,N_6905,N_6963);
or U7704 (N_7704,N_6590,N_6036);
or U7705 (N_7705,N_6498,N_6060);
nand U7706 (N_7706,N_6798,N_6557);
and U7707 (N_7707,N_6244,N_6206);
nand U7708 (N_7708,N_6277,N_6278);
nor U7709 (N_7709,N_6672,N_6897);
or U7710 (N_7710,N_6392,N_6272);
xnor U7711 (N_7711,N_6622,N_6680);
and U7712 (N_7712,N_6799,N_6855);
nand U7713 (N_7713,N_6745,N_6936);
nor U7714 (N_7714,N_6784,N_6326);
or U7715 (N_7715,N_6361,N_6596);
and U7716 (N_7716,N_6320,N_6459);
nand U7717 (N_7717,N_6805,N_6437);
or U7718 (N_7718,N_6527,N_6086);
and U7719 (N_7719,N_6921,N_6115);
nor U7720 (N_7720,N_6273,N_6323);
nor U7721 (N_7721,N_6905,N_6517);
or U7722 (N_7722,N_6747,N_6722);
nor U7723 (N_7723,N_6416,N_6347);
and U7724 (N_7724,N_6238,N_6753);
or U7725 (N_7725,N_6742,N_6594);
and U7726 (N_7726,N_6547,N_6046);
nand U7727 (N_7727,N_6232,N_6466);
xor U7728 (N_7728,N_6098,N_6554);
nand U7729 (N_7729,N_6656,N_6618);
or U7730 (N_7730,N_6547,N_6782);
and U7731 (N_7731,N_6322,N_6104);
or U7732 (N_7732,N_6124,N_6785);
and U7733 (N_7733,N_6734,N_6850);
xnor U7734 (N_7734,N_6467,N_6064);
and U7735 (N_7735,N_6022,N_6230);
nand U7736 (N_7736,N_6083,N_6790);
xor U7737 (N_7737,N_6111,N_6325);
or U7738 (N_7738,N_6165,N_6616);
or U7739 (N_7739,N_6809,N_6385);
and U7740 (N_7740,N_6355,N_6543);
nor U7741 (N_7741,N_6822,N_6640);
nand U7742 (N_7742,N_6166,N_6109);
nand U7743 (N_7743,N_6654,N_6539);
and U7744 (N_7744,N_6174,N_6334);
xor U7745 (N_7745,N_6501,N_6846);
nor U7746 (N_7746,N_6806,N_6638);
nor U7747 (N_7747,N_6289,N_6381);
and U7748 (N_7748,N_6996,N_6954);
nor U7749 (N_7749,N_6369,N_6239);
or U7750 (N_7750,N_6374,N_6699);
nor U7751 (N_7751,N_6701,N_6501);
nor U7752 (N_7752,N_6431,N_6459);
and U7753 (N_7753,N_6898,N_6749);
or U7754 (N_7754,N_6240,N_6607);
nand U7755 (N_7755,N_6355,N_6168);
nor U7756 (N_7756,N_6304,N_6518);
nand U7757 (N_7757,N_6280,N_6105);
nor U7758 (N_7758,N_6339,N_6657);
nor U7759 (N_7759,N_6855,N_6688);
or U7760 (N_7760,N_6405,N_6671);
nor U7761 (N_7761,N_6238,N_6623);
nor U7762 (N_7762,N_6787,N_6487);
or U7763 (N_7763,N_6597,N_6363);
and U7764 (N_7764,N_6750,N_6918);
and U7765 (N_7765,N_6923,N_6339);
and U7766 (N_7766,N_6939,N_6763);
or U7767 (N_7767,N_6261,N_6755);
or U7768 (N_7768,N_6123,N_6207);
and U7769 (N_7769,N_6596,N_6979);
xor U7770 (N_7770,N_6253,N_6390);
nand U7771 (N_7771,N_6686,N_6636);
or U7772 (N_7772,N_6254,N_6805);
xor U7773 (N_7773,N_6919,N_6870);
or U7774 (N_7774,N_6212,N_6508);
nand U7775 (N_7775,N_6634,N_6105);
xor U7776 (N_7776,N_6028,N_6259);
nor U7777 (N_7777,N_6200,N_6960);
nor U7778 (N_7778,N_6898,N_6772);
and U7779 (N_7779,N_6002,N_6902);
and U7780 (N_7780,N_6811,N_6934);
or U7781 (N_7781,N_6606,N_6192);
nand U7782 (N_7782,N_6759,N_6921);
nand U7783 (N_7783,N_6608,N_6340);
nor U7784 (N_7784,N_6746,N_6658);
or U7785 (N_7785,N_6591,N_6813);
and U7786 (N_7786,N_6120,N_6327);
and U7787 (N_7787,N_6596,N_6968);
nand U7788 (N_7788,N_6233,N_6100);
and U7789 (N_7789,N_6058,N_6005);
nand U7790 (N_7790,N_6886,N_6162);
nand U7791 (N_7791,N_6057,N_6383);
nor U7792 (N_7792,N_6887,N_6542);
nand U7793 (N_7793,N_6463,N_6176);
nand U7794 (N_7794,N_6551,N_6809);
or U7795 (N_7795,N_6946,N_6480);
and U7796 (N_7796,N_6762,N_6461);
nor U7797 (N_7797,N_6284,N_6072);
or U7798 (N_7798,N_6520,N_6291);
xnor U7799 (N_7799,N_6567,N_6222);
nand U7800 (N_7800,N_6354,N_6385);
or U7801 (N_7801,N_6722,N_6356);
and U7802 (N_7802,N_6458,N_6599);
and U7803 (N_7803,N_6152,N_6184);
nand U7804 (N_7804,N_6556,N_6884);
or U7805 (N_7805,N_6151,N_6671);
nor U7806 (N_7806,N_6596,N_6495);
nor U7807 (N_7807,N_6401,N_6659);
nor U7808 (N_7808,N_6936,N_6510);
nor U7809 (N_7809,N_6887,N_6666);
nor U7810 (N_7810,N_6621,N_6802);
nor U7811 (N_7811,N_6127,N_6535);
nand U7812 (N_7812,N_6757,N_6477);
or U7813 (N_7813,N_6463,N_6578);
nor U7814 (N_7814,N_6225,N_6073);
and U7815 (N_7815,N_6487,N_6011);
and U7816 (N_7816,N_6615,N_6722);
and U7817 (N_7817,N_6242,N_6564);
nor U7818 (N_7818,N_6389,N_6073);
and U7819 (N_7819,N_6363,N_6214);
nor U7820 (N_7820,N_6207,N_6978);
and U7821 (N_7821,N_6715,N_6396);
xnor U7822 (N_7822,N_6597,N_6673);
or U7823 (N_7823,N_6895,N_6477);
nor U7824 (N_7824,N_6606,N_6764);
or U7825 (N_7825,N_6254,N_6270);
nand U7826 (N_7826,N_6240,N_6625);
xor U7827 (N_7827,N_6196,N_6800);
or U7828 (N_7828,N_6226,N_6077);
and U7829 (N_7829,N_6632,N_6362);
nor U7830 (N_7830,N_6508,N_6849);
and U7831 (N_7831,N_6083,N_6497);
nor U7832 (N_7832,N_6328,N_6520);
or U7833 (N_7833,N_6193,N_6910);
xor U7834 (N_7834,N_6620,N_6683);
nand U7835 (N_7835,N_6387,N_6110);
and U7836 (N_7836,N_6350,N_6976);
nand U7837 (N_7837,N_6264,N_6468);
or U7838 (N_7838,N_6014,N_6570);
nor U7839 (N_7839,N_6999,N_6197);
and U7840 (N_7840,N_6176,N_6802);
nand U7841 (N_7841,N_6860,N_6060);
and U7842 (N_7842,N_6229,N_6917);
and U7843 (N_7843,N_6693,N_6594);
nand U7844 (N_7844,N_6812,N_6831);
nor U7845 (N_7845,N_6078,N_6048);
nor U7846 (N_7846,N_6387,N_6945);
nor U7847 (N_7847,N_6530,N_6111);
and U7848 (N_7848,N_6649,N_6778);
and U7849 (N_7849,N_6554,N_6315);
xnor U7850 (N_7850,N_6841,N_6970);
nand U7851 (N_7851,N_6376,N_6111);
or U7852 (N_7852,N_6135,N_6994);
or U7853 (N_7853,N_6149,N_6848);
or U7854 (N_7854,N_6794,N_6377);
and U7855 (N_7855,N_6000,N_6613);
nand U7856 (N_7856,N_6801,N_6804);
nand U7857 (N_7857,N_6732,N_6337);
nor U7858 (N_7858,N_6167,N_6040);
or U7859 (N_7859,N_6919,N_6731);
xnor U7860 (N_7860,N_6015,N_6713);
xor U7861 (N_7861,N_6730,N_6774);
xnor U7862 (N_7862,N_6544,N_6026);
nand U7863 (N_7863,N_6913,N_6188);
nand U7864 (N_7864,N_6569,N_6721);
and U7865 (N_7865,N_6545,N_6026);
nand U7866 (N_7866,N_6311,N_6853);
nor U7867 (N_7867,N_6928,N_6680);
or U7868 (N_7868,N_6350,N_6245);
or U7869 (N_7869,N_6057,N_6811);
nand U7870 (N_7870,N_6802,N_6469);
nor U7871 (N_7871,N_6303,N_6222);
nor U7872 (N_7872,N_6506,N_6924);
nor U7873 (N_7873,N_6705,N_6528);
or U7874 (N_7874,N_6120,N_6864);
nand U7875 (N_7875,N_6867,N_6231);
and U7876 (N_7876,N_6241,N_6634);
nand U7877 (N_7877,N_6920,N_6686);
nand U7878 (N_7878,N_6504,N_6852);
and U7879 (N_7879,N_6895,N_6808);
xnor U7880 (N_7880,N_6764,N_6624);
nor U7881 (N_7881,N_6307,N_6566);
nor U7882 (N_7882,N_6572,N_6474);
and U7883 (N_7883,N_6231,N_6698);
and U7884 (N_7884,N_6056,N_6451);
nand U7885 (N_7885,N_6368,N_6859);
nor U7886 (N_7886,N_6319,N_6979);
and U7887 (N_7887,N_6899,N_6420);
nand U7888 (N_7888,N_6593,N_6006);
xor U7889 (N_7889,N_6075,N_6605);
or U7890 (N_7890,N_6147,N_6662);
nor U7891 (N_7891,N_6687,N_6456);
nand U7892 (N_7892,N_6266,N_6423);
nand U7893 (N_7893,N_6263,N_6987);
nor U7894 (N_7894,N_6941,N_6918);
nand U7895 (N_7895,N_6832,N_6925);
and U7896 (N_7896,N_6451,N_6110);
and U7897 (N_7897,N_6068,N_6930);
and U7898 (N_7898,N_6806,N_6017);
nand U7899 (N_7899,N_6708,N_6096);
and U7900 (N_7900,N_6926,N_6274);
nor U7901 (N_7901,N_6886,N_6133);
nand U7902 (N_7902,N_6806,N_6892);
and U7903 (N_7903,N_6565,N_6994);
or U7904 (N_7904,N_6796,N_6969);
and U7905 (N_7905,N_6278,N_6567);
and U7906 (N_7906,N_6259,N_6164);
or U7907 (N_7907,N_6113,N_6810);
nor U7908 (N_7908,N_6860,N_6707);
nand U7909 (N_7909,N_6200,N_6349);
nor U7910 (N_7910,N_6133,N_6606);
or U7911 (N_7911,N_6621,N_6893);
nor U7912 (N_7912,N_6860,N_6280);
and U7913 (N_7913,N_6316,N_6889);
or U7914 (N_7914,N_6789,N_6358);
or U7915 (N_7915,N_6419,N_6119);
nor U7916 (N_7916,N_6571,N_6848);
xnor U7917 (N_7917,N_6021,N_6024);
and U7918 (N_7918,N_6300,N_6354);
and U7919 (N_7919,N_6005,N_6268);
nor U7920 (N_7920,N_6992,N_6026);
nor U7921 (N_7921,N_6252,N_6516);
and U7922 (N_7922,N_6511,N_6084);
or U7923 (N_7923,N_6266,N_6153);
nor U7924 (N_7924,N_6793,N_6003);
nor U7925 (N_7925,N_6263,N_6285);
and U7926 (N_7926,N_6553,N_6873);
xnor U7927 (N_7927,N_6329,N_6473);
nor U7928 (N_7928,N_6791,N_6857);
nand U7929 (N_7929,N_6693,N_6000);
nand U7930 (N_7930,N_6549,N_6275);
or U7931 (N_7931,N_6327,N_6186);
nor U7932 (N_7932,N_6845,N_6532);
nand U7933 (N_7933,N_6263,N_6267);
or U7934 (N_7934,N_6477,N_6198);
nor U7935 (N_7935,N_6498,N_6504);
nand U7936 (N_7936,N_6109,N_6366);
xnor U7937 (N_7937,N_6918,N_6118);
nor U7938 (N_7938,N_6923,N_6219);
nand U7939 (N_7939,N_6149,N_6908);
and U7940 (N_7940,N_6946,N_6993);
nor U7941 (N_7941,N_6958,N_6488);
and U7942 (N_7942,N_6008,N_6160);
nand U7943 (N_7943,N_6635,N_6815);
or U7944 (N_7944,N_6158,N_6842);
nand U7945 (N_7945,N_6405,N_6048);
or U7946 (N_7946,N_6463,N_6576);
or U7947 (N_7947,N_6150,N_6653);
or U7948 (N_7948,N_6596,N_6029);
xnor U7949 (N_7949,N_6926,N_6035);
nor U7950 (N_7950,N_6667,N_6153);
xor U7951 (N_7951,N_6209,N_6486);
nor U7952 (N_7952,N_6545,N_6878);
or U7953 (N_7953,N_6804,N_6435);
nor U7954 (N_7954,N_6922,N_6707);
or U7955 (N_7955,N_6567,N_6002);
and U7956 (N_7956,N_6266,N_6567);
and U7957 (N_7957,N_6253,N_6028);
and U7958 (N_7958,N_6977,N_6103);
nand U7959 (N_7959,N_6495,N_6720);
nand U7960 (N_7960,N_6965,N_6569);
and U7961 (N_7961,N_6411,N_6950);
and U7962 (N_7962,N_6047,N_6554);
and U7963 (N_7963,N_6101,N_6495);
nand U7964 (N_7964,N_6799,N_6659);
nand U7965 (N_7965,N_6344,N_6066);
xor U7966 (N_7966,N_6053,N_6385);
nand U7967 (N_7967,N_6333,N_6881);
and U7968 (N_7968,N_6807,N_6013);
or U7969 (N_7969,N_6847,N_6128);
nand U7970 (N_7970,N_6485,N_6620);
nor U7971 (N_7971,N_6271,N_6240);
nand U7972 (N_7972,N_6550,N_6042);
xor U7973 (N_7973,N_6869,N_6167);
nand U7974 (N_7974,N_6209,N_6583);
nand U7975 (N_7975,N_6958,N_6345);
and U7976 (N_7976,N_6355,N_6055);
or U7977 (N_7977,N_6532,N_6450);
and U7978 (N_7978,N_6246,N_6515);
nand U7979 (N_7979,N_6917,N_6672);
or U7980 (N_7980,N_6199,N_6711);
nor U7981 (N_7981,N_6919,N_6020);
nor U7982 (N_7982,N_6113,N_6840);
nand U7983 (N_7983,N_6931,N_6399);
and U7984 (N_7984,N_6873,N_6316);
nand U7985 (N_7985,N_6427,N_6523);
nand U7986 (N_7986,N_6121,N_6497);
nor U7987 (N_7987,N_6159,N_6278);
xnor U7988 (N_7988,N_6369,N_6460);
nor U7989 (N_7989,N_6648,N_6843);
nand U7990 (N_7990,N_6018,N_6839);
nor U7991 (N_7991,N_6787,N_6575);
and U7992 (N_7992,N_6034,N_6751);
nand U7993 (N_7993,N_6260,N_6044);
nand U7994 (N_7994,N_6772,N_6635);
nand U7995 (N_7995,N_6109,N_6155);
nor U7996 (N_7996,N_6930,N_6369);
nand U7997 (N_7997,N_6935,N_6559);
and U7998 (N_7998,N_6049,N_6360);
nand U7999 (N_7999,N_6667,N_6291);
and U8000 (N_8000,N_7419,N_7480);
nand U8001 (N_8001,N_7500,N_7114);
nor U8002 (N_8002,N_7659,N_7612);
nor U8003 (N_8003,N_7970,N_7215);
or U8004 (N_8004,N_7524,N_7903);
nand U8005 (N_8005,N_7740,N_7210);
nor U8006 (N_8006,N_7607,N_7559);
nor U8007 (N_8007,N_7562,N_7532);
or U8008 (N_8008,N_7365,N_7546);
and U8009 (N_8009,N_7677,N_7466);
and U8010 (N_8010,N_7759,N_7953);
nor U8011 (N_8011,N_7795,N_7023);
nor U8012 (N_8012,N_7905,N_7248);
nor U8013 (N_8013,N_7827,N_7609);
and U8014 (N_8014,N_7338,N_7586);
or U8015 (N_8015,N_7197,N_7367);
and U8016 (N_8016,N_7025,N_7521);
and U8017 (N_8017,N_7582,N_7848);
and U8018 (N_8018,N_7307,N_7530);
or U8019 (N_8019,N_7988,N_7637);
and U8020 (N_8020,N_7671,N_7774);
nor U8021 (N_8021,N_7491,N_7969);
xnor U8022 (N_8022,N_7997,N_7817);
and U8023 (N_8023,N_7856,N_7601);
or U8024 (N_8024,N_7138,N_7155);
and U8025 (N_8025,N_7029,N_7372);
and U8026 (N_8026,N_7018,N_7212);
nor U8027 (N_8027,N_7523,N_7489);
or U8028 (N_8028,N_7353,N_7031);
and U8029 (N_8029,N_7900,N_7726);
or U8030 (N_8030,N_7450,N_7922);
nor U8031 (N_8031,N_7719,N_7065);
nand U8032 (N_8032,N_7995,N_7376);
and U8033 (N_8033,N_7460,N_7705);
or U8034 (N_8034,N_7429,N_7973);
and U8035 (N_8035,N_7946,N_7402);
or U8036 (N_8036,N_7454,N_7565);
or U8037 (N_8037,N_7685,N_7139);
nor U8038 (N_8038,N_7068,N_7805);
and U8039 (N_8039,N_7295,N_7779);
and U8040 (N_8040,N_7405,N_7787);
and U8041 (N_8041,N_7940,N_7157);
nand U8042 (N_8042,N_7002,N_7878);
or U8043 (N_8043,N_7588,N_7178);
or U8044 (N_8044,N_7301,N_7538);
nand U8045 (N_8045,N_7358,N_7391);
and U8046 (N_8046,N_7596,N_7886);
xor U8047 (N_8047,N_7704,N_7778);
or U8048 (N_8048,N_7964,N_7850);
or U8049 (N_8049,N_7716,N_7933);
and U8050 (N_8050,N_7238,N_7789);
or U8051 (N_8051,N_7870,N_7724);
nand U8052 (N_8052,N_7649,N_7552);
nand U8053 (N_8053,N_7600,N_7110);
nand U8054 (N_8054,N_7116,N_7161);
or U8055 (N_8055,N_7978,N_7881);
and U8056 (N_8056,N_7887,N_7478);
nand U8057 (N_8057,N_7822,N_7440);
xor U8058 (N_8058,N_7811,N_7245);
or U8059 (N_8059,N_7496,N_7807);
and U8060 (N_8060,N_7132,N_7578);
nor U8061 (N_8061,N_7217,N_7333);
and U8062 (N_8062,N_7776,N_7207);
xnor U8063 (N_8063,N_7050,N_7961);
or U8064 (N_8064,N_7173,N_7077);
and U8065 (N_8065,N_7738,N_7854);
and U8066 (N_8066,N_7912,N_7472);
or U8067 (N_8067,N_7640,N_7696);
nand U8068 (N_8068,N_7202,N_7182);
nor U8069 (N_8069,N_7543,N_7192);
nand U8070 (N_8070,N_7894,N_7263);
nor U8071 (N_8071,N_7209,N_7330);
xnor U8072 (N_8072,N_7525,N_7769);
xnor U8073 (N_8073,N_7898,N_7979);
nand U8074 (N_8074,N_7184,N_7583);
and U8075 (N_8075,N_7258,N_7698);
and U8076 (N_8076,N_7804,N_7166);
nand U8077 (N_8077,N_7022,N_7368);
or U8078 (N_8078,N_7336,N_7400);
and U8079 (N_8079,N_7357,N_7104);
and U8080 (N_8080,N_7843,N_7921);
or U8081 (N_8081,N_7679,N_7529);
xnor U8082 (N_8082,N_7066,N_7619);
nor U8083 (N_8083,N_7510,N_7722);
nor U8084 (N_8084,N_7329,N_7935);
nand U8085 (N_8085,N_7823,N_7259);
nor U8086 (N_8086,N_7063,N_7540);
and U8087 (N_8087,N_7305,N_7627);
and U8088 (N_8088,N_7061,N_7622);
or U8089 (N_8089,N_7183,N_7687);
nor U8090 (N_8090,N_7032,N_7320);
nand U8091 (N_8091,N_7651,N_7852);
or U8092 (N_8092,N_7474,N_7732);
nand U8093 (N_8093,N_7153,N_7008);
and U8094 (N_8094,N_7513,N_7845);
nor U8095 (N_8095,N_7869,N_7929);
nor U8096 (N_8096,N_7299,N_7322);
or U8097 (N_8097,N_7624,N_7415);
nor U8098 (N_8098,N_7163,N_7392);
nand U8099 (N_8099,N_7831,N_7051);
nor U8100 (N_8100,N_7941,N_7052);
or U8101 (N_8101,N_7060,N_7930);
and U8102 (N_8102,N_7587,N_7455);
xor U8103 (N_8103,N_7802,N_7545);
nand U8104 (N_8104,N_7526,N_7409);
and U8105 (N_8105,N_7420,N_7959);
or U8106 (N_8106,N_7119,N_7571);
xnor U8107 (N_8107,N_7319,N_7731);
or U8108 (N_8108,N_7105,N_7218);
and U8109 (N_8109,N_7663,N_7620);
and U8110 (N_8110,N_7554,N_7385);
or U8111 (N_8111,N_7047,N_7889);
and U8112 (N_8112,N_7884,N_7388);
or U8113 (N_8113,N_7511,N_7862);
nor U8114 (N_8114,N_7390,N_7252);
nor U8115 (N_8115,N_7021,N_7493);
xor U8116 (N_8116,N_7304,N_7230);
nor U8117 (N_8117,N_7610,N_7585);
nor U8118 (N_8118,N_7243,N_7851);
or U8119 (N_8119,N_7115,N_7377);
nor U8120 (N_8120,N_7593,N_7793);
xnor U8121 (N_8121,N_7767,N_7280);
nand U8122 (N_8122,N_7577,N_7459);
or U8123 (N_8123,N_7276,N_7556);
or U8124 (N_8124,N_7824,N_7707);
nor U8125 (N_8125,N_7384,N_7439);
and U8126 (N_8126,N_7356,N_7968);
nand U8127 (N_8127,N_7855,N_7414);
nand U8128 (N_8128,N_7026,N_7096);
xnor U8129 (N_8129,N_7818,N_7290);
and U8130 (N_8130,N_7312,N_7124);
nor U8131 (N_8131,N_7794,N_7902);
and U8132 (N_8132,N_7505,N_7058);
and U8133 (N_8133,N_7265,N_7531);
and U8134 (N_8134,N_7594,N_7380);
and U8135 (N_8135,N_7099,N_7249);
and U8136 (N_8136,N_7150,N_7581);
or U8137 (N_8137,N_7470,N_7433);
nand U8138 (N_8138,N_7448,N_7499);
nand U8139 (N_8139,N_7713,N_7048);
nor U8140 (N_8140,N_7362,N_7225);
nand U8141 (N_8141,N_7498,N_7275);
or U8142 (N_8142,N_7700,N_7798);
nand U8143 (N_8143,N_7131,N_7840);
nand U8144 (N_8144,N_7931,N_7465);
nor U8145 (N_8145,N_7289,N_7246);
or U8146 (N_8146,N_7378,N_7345);
or U8147 (N_8147,N_7014,N_7788);
nor U8148 (N_8148,N_7042,N_7867);
and U8149 (N_8149,N_7231,N_7681);
nand U8150 (N_8150,N_7170,N_7775);
or U8151 (N_8151,N_7591,N_7118);
nor U8152 (N_8152,N_7514,N_7974);
nand U8153 (N_8153,N_7736,N_7201);
or U8154 (N_8154,N_7062,N_7456);
xnor U8155 (N_8155,N_7885,N_7171);
nor U8156 (N_8156,N_7172,N_7605);
and U8157 (N_8157,N_7348,N_7294);
or U8158 (N_8158,N_7471,N_7355);
nand U8159 (N_8159,N_7085,N_7036);
nor U8160 (N_8160,N_7999,N_7741);
nor U8161 (N_8161,N_7200,N_7809);
and U8162 (N_8162,N_7302,N_7560);
nor U8163 (N_8163,N_7948,N_7866);
nor U8164 (N_8164,N_7650,N_7092);
nor U8165 (N_8165,N_7227,N_7684);
and U8166 (N_8166,N_7401,N_7914);
or U8167 (N_8167,N_7495,N_7223);
and U8168 (N_8168,N_7045,N_7241);
nand U8169 (N_8169,N_7670,N_7232);
and U8170 (N_8170,N_7516,N_7806);
nor U8171 (N_8171,N_7690,N_7396);
and U8172 (N_8172,N_7148,N_7069);
nor U8173 (N_8173,N_7725,N_7782);
nand U8174 (N_8174,N_7980,N_7261);
or U8175 (N_8175,N_7548,N_7688);
and U8176 (N_8176,N_7476,N_7342);
nand U8177 (N_8177,N_7557,N_7568);
and U8178 (N_8178,N_7360,N_7167);
or U8179 (N_8179,N_7379,N_7247);
nand U8180 (N_8180,N_7760,N_7418);
or U8181 (N_8181,N_7103,N_7177);
and U8182 (N_8182,N_7542,N_7638);
nor U8183 (N_8183,N_7134,N_7221);
nor U8184 (N_8184,N_7686,N_7094);
nor U8185 (N_8185,N_7438,N_7043);
and U8186 (N_8186,N_7120,N_7475);
nor U8187 (N_8187,N_7936,N_7947);
and U8188 (N_8188,N_7720,N_7692);
nand U8189 (N_8189,N_7175,N_7410);
xnor U8190 (N_8190,N_7044,N_7703);
nand U8191 (N_8191,N_7370,N_7332);
or U8192 (N_8192,N_7815,N_7626);
nand U8193 (N_8193,N_7925,N_7920);
and U8194 (N_8194,N_7313,N_7204);
nor U8195 (N_8195,N_7235,N_7539);
and U8196 (N_8196,N_7727,N_7352);
and U8197 (N_8197,N_7458,N_7484);
or U8198 (N_8198,N_7233,N_7211);
or U8199 (N_8199,N_7917,N_7697);
and U8200 (N_8200,N_7229,N_7615);
and U8201 (N_8201,N_7468,N_7250);
xor U8202 (N_8202,N_7563,N_7618);
nor U8203 (N_8203,N_7287,N_7897);
nor U8204 (N_8204,N_7162,N_7359);
or U8205 (N_8205,N_7363,N_7340);
nand U8206 (N_8206,N_7130,N_7187);
xor U8207 (N_8207,N_7133,N_7989);
or U8208 (N_8208,N_7269,N_7966);
xnor U8209 (N_8209,N_7317,N_7088);
nor U8210 (N_8210,N_7196,N_7706);
nor U8211 (N_8211,N_7151,N_7205);
nor U8212 (N_8212,N_7518,N_7399);
and U8213 (N_8213,N_7003,N_7676);
or U8214 (N_8214,N_7303,N_7464);
xor U8215 (N_8215,N_7708,N_7871);
nor U8216 (N_8216,N_7982,N_7279);
nand U8217 (N_8217,N_7469,N_7331);
nor U8218 (N_8218,N_7764,N_7642);
xnor U8219 (N_8219,N_7836,N_7857);
xnor U8220 (N_8220,N_7406,N_7631);
xnor U8221 (N_8221,N_7604,N_7617);
nand U8222 (N_8222,N_7628,N_7408);
or U8223 (N_8223,N_7254,N_7971);
and U8224 (N_8224,N_7260,N_7424);
nand U8225 (N_8225,N_7723,N_7423);
and U8226 (N_8226,N_7517,N_7444);
and U8227 (N_8227,N_7747,N_7387);
nor U8228 (N_8228,N_7452,N_7300);
xor U8229 (N_8229,N_7658,N_7037);
xor U8230 (N_8230,N_7007,N_7435);
xnor U8231 (N_8231,N_7100,N_7504);
xor U8232 (N_8232,N_7812,N_7841);
nor U8233 (N_8233,N_7195,N_7830);
nor U8234 (N_8234,N_7761,N_7743);
and U8235 (N_8235,N_7519,N_7821);
nand U8236 (N_8236,N_7951,N_7801);
nand U8237 (N_8237,N_7645,N_7421);
and U8238 (N_8238,N_7534,N_7797);
nand U8239 (N_8239,N_7570,N_7799);
nand U8240 (N_8240,N_7441,N_7773);
nand U8241 (N_8241,N_7004,N_7427);
nand U8242 (N_8242,N_7832,N_7189);
nand U8243 (N_8243,N_7506,N_7371);
nor U8244 (N_8244,N_7579,N_7009);
and U8245 (N_8245,N_7298,N_7580);
and U8246 (N_8246,N_7839,N_7567);
nor U8247 (N_8247,N_7373,N_7907);
nand U8248 (N_8248,N_7111,N_7286);
or U8249 (N_8249,N_7636,N_7820);
xor U8250 (N_8250,N_7006,N_7284);
xor U8251 (N_8251,N_7422,N_7923);
or U8252 (N_8252,N_7654,N_7070);
or U8253 (N_8253,N_7666,N_7086);
xnor U8254 (N_8254,N_7486,N_7220);
nand U8255 (N_8255,N_7792,N_7056);
nand U8256 (N_8256,N_7266,N_7990);
nor U8257 (N_8257,N_7149,N_7308);
nand U8258 (N_8258,N_7093,N_7785);
xor U8259 (N_8259,N_7592,N_7129);
nor U8260 (N_8260,N_7411,N_7730);
or U8261 (N_8261,N_7674,N_7143);
xor U8262 (N_8262,N_7208,N_7906);
nand U8263 (N_8263,N_7253,N_7739);
or U8264 (N_8264,N_7680,N_7262);
nand U8265 (N_8265,N_7672,N_7011);
or U8266 (N_8266,N_7347,N_7547);
nor U8267 (N_8267,N_7780,N_7492);
or U8268 (N_8268,N_7494,N_7842);
and U8269 (N_8269,N_7437,N_7828);
and U8270 (N_8270,N_7017,N_7950);
and U8271 (N_8271,N_7012,N_7657);
nand U8272 (N_8272,N_7430,N_7228);
nand U8273 (N_8273,N_7834,N_7122);
and U8274 (N_8274,N_7569,N_7899);
nor U8275 (N_8275,N_7351,N_7853);
nor U8276 (N_8276,N_7381,N_7847);
or U8277 (N_8277,N_7781,N_7436);
nor U8278 (N_8278,N_7996,N_7074);
xor U8279 (N_8279,N_7140,N_7135);
and U8280 (N_8280,N_7306,N_7669);
nand U8281 (N_8281,N_7644,N_7264);
nand U8282 (N_8282,N_7909,N_7758);
and U8283 (N_8283,N_7473,N_7763);
or U8284 (N_8284,N_7431,N_7354);
or U8285 (N_8285,N_7369,N_7653);
and U8286 (N_8286,N_7753,N_7236);
or U8287 (N_8287,N_7020,N_7323);
nand U8288 (N_8288,N_7908,N_7942);
nand U8289 (N_8289,N_7611,N_7891);
and U8290 (N_8290,N_7702,N_7179);
and U8291 (N_8291,N_7034,N_7710);
or U8292 (N_8292,N_7310,N_7326);
and U8293 (N_8293,N_7549,N_7112);
or U8294 (N_8294,N_7507,N_7107);
and U8295 (N_8295,N_7718,N_7937);
xnor U8296 (N_8296,N_7682,N_7589);
nand U8297 (N_8297,N_7616,N_7413);
or U8298 (N_8298,N_7904,N_7482);
nor U8299 (N_8299,N_7064,N_7483);
and U8300 (N_8300,N_7629,N_7488);
and U8301 (N_8301,N_7734,N_7271);
or U8302 (N_8302,N_7386,N_7960);
and U8303 (N_8303,N_7224,N_7939);
nand U8304 (N_8304,N_7084,N_7555);
nor U8305 (N_8305,N_7136,N_7872);
or U8306 (N_8306,N_7544,N_7407);
or U8307 (N_8307,N_7442,N_7079);
nand U8308 (N_8308,N_7695,N_7073);
nor U8309 (N_8309,N_7327,N_7206);
or U8310 (N_8310,N_7467,N_7987);
nor U8311 (N_8311,N_7274,N_7146);
and U8312 (N_8312,N_7551,N_7389);
nor U8313 (N_8313,N_7113,N_7394);
or U8314 (N_8314,N_7028,N_7334);
or U8315 (N_8315,N_7846,N_7984);
nand U8316 (N_8316,N_7145,N_7267);
and U8317 (N_8317,N_7943,N_7101);
xor U8318 (N_8318,N_7983,N_7533);
xnor U8319 (N_8319,N_7662,N_7076);
nor U8320 (N_8320,N_7621,N_7875);
xnor U8321 (N_8321,N_7463,N_7515);
or U8322 (N_8322,N_7282,N_7522);
or U8323 (N_8323,N_7457,N_7185);
or U8324 (N_8324,N_7121,N_7913);
nor U8325 (N_8325,N_7374,N_7054);
or U8326 (N_8326,N_7072,N_7558);
or U8327 (N_8327,N_7046,N_7152);
nand U8328 (N_8328,N_7098,N_7715);
or U8329 (N_8329,N_7655,N_7991);
nor U8330 (N_8330,N_7154,N_7451);
xor U8331 (N_8331,N_7337,N_7089);
or U8332 (N_8332,N_7998,N_7453);
nand U8333 (N_8333,N_7067,N_7016);
or U8334 (N_8334,N_7599,N_7994);
and U8335 (N_8335,N_7859,N_7417);
nor U8336 (N_8336,N_7024,N_7144);
xor U8337 (N_8337,N_7993,N_7520);
and U8338 (N_8338,N_7838,N_7826);
xor U8339 (N_8339,N_7075,N_7040);
xnor U8340 (N_8340,N_7892,N_7268);
and U8341 (N_8341,N_7646,N_7039);
or U8342 (N_8342,N_7382,N_7728);
or U8343 (N_8343,N_7364,N_7564);
nand U8344 (N_8344,N_7746,N_7479);
and U8345 (N_8345,N_7693,N_7485);
and U8346 (N_8346,N_7311,N_7639);
or U8347 (N_8347,N_7919,N_7770);
or U8348 (N_8348,N_7689,N_7019);
and U8349 (N_8349,N_7833,N_7446);
nor U8350 (N_8350,N_7501,N_7814);
nor U8351 (N_8351,N_7749,N_7010);
nand U8352 (N_8352,N_7324,N_7890);
and U8353 (N_8353,N_7273,N_7328);
or U8354 (N_8354,N_7709,N_7733);
and U8355 (N_8355,N_7508,N_7745);
nor U8356 (N_8356,N_7366,N_7927);
and U8357 (N_8357,N_7194,N_7729);
or U8358 (N_8358,N_7321,N_7712);
nor U8359 (N_8359,N_7606,N_7127);
or U8360 (N_8360,N_7952,N_7967);
nor U8361 (N_8361,N_7090,N_7277);
nor U8362 (N_8362,N_7945,N_7876);
nor U8363 (N_8363,N_7035,N_7608);
nand U8364 (N_8364,N_7240,N_7123);
nor U8365 (N_8365,N_7678,N_7791);
nor U8366 (N_8366,N_7222,N_7633);
nand U8367 (N_8367,N_7180,N_7675);
nand U8368 (N_8368,N_7958,N_7752);
and U8369 (N_8369,N_7916,N_7428);
or U8370 (N_8370,N_7445,N_7783);
or U8371 (N_8371,N_7575,N_7944);
or U8372 (N_8372,N_7270,N_7765);
nor U8373 (N_8373,N_7398,N_7449);
xor U8374 (N_8374,N_7176,N_7819);
nor U8375 (N_8375,N_7535,N_7314);
nor U8376 (N_8376,N_7393,N_7226);
nand U8377 (N_8377,N_7893,N_7203);
and U8378 (N_8378,N_7701,N_7160);
or U8379 (N_8379,N_7896,N_7717);
and U8380 (N_8380,N_7808,N_7986);
nand U8381 (N_8381,N_7137,N_7404);
xor U8382 (N_8382,N_7335,N_7158);
or U8383 (N_8383,N_7186,N_7080);
nand U8384 (N_8384,N_7087,N_7790);
nand U8385 (N_8385,N_7901,N_7873);
or U8386 (N_8386,N_7656,N_7613);
nand U8387 (N_8387,N_7647,N_7584);
nor U8388 (N_8388,N_7985,N_7648);
or U8389 (N_8389,N_7879,N_7497);
nand U8390 (N_8390,N_7877,N_7000);
and U8391 (N_8391,N_7863,N_7426);
nand U8392 (N_8392,N_7316,N_7188);
nor U8393 (N_8393,N_7572,N_7315);
nand U8394 (N_8394,N_7432,N_7512);
or U8395 (N_8395,N_7341,N_7256);
and U8396 (N_8396,N_7527,N_7038);
and U8397 (N_8397,N_7918,N_7053);
and U8398 (N_8398,N_7837,N_7574);
or U8399 (N_8399,N_7447,N_7934);
or U8400 (N_8400,N_7285,N_7748);
and U8401 (N_8401,N_7536,N_7796);
nand U8402 (N_8402,N_7962,N_7005);
xnor U8403 (N_8403,N_7643,N_7434);
or U8404 (N_8404,N_7566,N_7537);
and U8405 (N_8405,N_7383,N_7237);
or U8406 (N_8406,N_7425,N_7641);
nor U8407 (N_8407,N_7403,N_7234);
xor U8408 (N_8408,N_7976,N_7082);
or U8409 (N_8409,N_7754,N_7757);
and U8410 (N_8410,N_7296,N_7078);
nor U8411 (N_8411,N_7095,N_7281);
xor U8412 (N_8412,N_7255,N_7668);
and U8413 (N_8413,N_7813,N_7126);
nand U8414 (N_8414,N_7954,N_7128);
or U8415 (N_8415,N_7156,N_7766);
and U8416 (N_8416,N_7125,N_7168);
nor U8417 (N_8417,N_7957,N_7597);
nand U8418 (N_8418,N_7963,N_7926);
and U8419 (N_8419,N_7595,N_7142);
xnor U8420 (N_8420,N_7829,N_7242);
nand U8421 (N_8421,N_7932,N_7590);
nand U8422 (N_8422,N_7938,N_7015);
nor U8423 (N_8423,N_7652,N_7573);
and U8424 (N_8424,N_7291,N_7057);
and U8425 (N_8425,N_7239,N_7803);
xnor U8426 (N_8426,N_7744,N_7602);
nor U8427 (N_8427,N_7293,N_7667);
nor U8428 (N_8428,N_7816,N_7825);
nand U8429 (N_8429,N_7477,N_7462);
nand U8430 (N_8430,N_7750,N_7216);
xnor U8431 (N_8431,N_7159,N_7972);
or U8432 (N_8432,N_7771,N_7956);
nor U8433 (N_8433,N_7858,N_7198);
nand U8434 (N_8434,N_7349,N_7660);
or U8435 (N_8435,N_7001,N_7880);
xor U8436 (N_8436,N_7509,N_7768);
nor U8437 (N_8437,N_7059,N_7911);
or U8438 (N_8438,N_7083,N_7461);
nand U8439 (N_8439,N_7106,N_7292);
nand U8440 (N_8440,N_7055,N_7735);
nand U8441 (N_8441,N_7108,N_7257);
nor U8442 (N_8442,N_7861,N_7346);
nand U8443 (N_8443,N_7244,N_7283);
xnor U8444 (N_8444,N_7214,N_7071);
xor U8445 (N_8445,N_7416,N_7755);
nand U8446 (N_8446,N_7864,N_7190);
and U8447 (N_8447,N_7502,N_7213);
or U8448 (N_8448,N_7949,N_7109);
nor U8449 (N_8449,N_7910,N_7924);
or U8450 (N_8450,N_7251,N_7598);
nor U8451 (N_8451,N_7888,N_7165);
and U8452 (N_8452,N_7711,N_7772);
and U8453 (N_8453,N_7849,N_7343);
and U8454 (N_8454,N_7683,N_7030);
nand U8455 (N_8455,N_7883,N_7786);
or U8456 (N_8456,N_7141,N_7350);
and U8457 (N_8457,N_7977,N_7844);
xor U8458 (N_8458,N_7714,N_7091);
nand U8459 (N_8459,N_7375,N_7219);
nor U8460 (N_8460,N_7550,N_7955);
and U8461 (N_8461,N_7325,N_7117);
xnor U8462 (N_8462,N_7721,N_7528);
or U8463 (N_8463,N_7865,N_7634);
or U8464 (N_8464,N_7412,N_7835);
and U8465 (N_8465,N_7874,N_7868);
nor U8466 (N_8466,N_7756,N_7965);
nand U8467 (N_8467,N_7975,N_7481);
nand U8468 (N_8468,N_7751,N_7625);
or U8469 (N_8469,N_7742,N_7199);
and U8470 (N_8470,N_7603,N_7191);
or U8471 (N_8471,N_7033,N_7561);
nor U8472 (N_8472,N_7164,N_7297);
nor U8473 (N_8473,N_7981,N_7694);
nand U8474 (N_8474,N_7102,N_7027);
nand U8475 (N_8475,N_7288,N_7395);
nor U8476 (N_8476,N_7915,N_7699);
and U8477 (N_8477,N_7553,N_7800);
and U8478 (N_8478,N_7661,N_7397);
nand U8479 (N_8479,N_7673,N_7635);
or U8480 (N_8480,N_7193,N_7049);
nand U8481 (N_8481,N_7632,N_7097);
or U8482 (N_8482,N_7013,N_7503);
and U8483 (N_8483,N_7882,N_7777);
or U8484 (N_8484,N_7147,N_7169);
and U8485 (N_8485,N_7490,N_7762);
and U8486 (N_8486,N_7541,N_7344);
or U8487 (N_8487,N_7614,N_7928);
nor U8488 (N_8488,N_7623,N_7487);
nand U8489 (N_8489,N_7664,N_7041);
xor U8490 (N_8490,N_7318,N_7737);
or U8491 (N_8491,N_7576,N_7810);
nor U8492 (N_8492,N_7361,N_7443);
and U8493 (N_8493,N_7895,N_7278);
or U8494 (N_8494,N_7691,N_7174);
nor U8495 (N_8495,N_7339,N_7784);
or U8496 (N_8496,N_7630,N_7081);
nor U8497 (N_8497,N_7992,N_7665);
xnor U8498 (N_8498,N_7309,N_7272);
or U8499 (N_8499,N_7860,N_7181);
nor U8500 (N_8500,N_7267,N_7158);
nand U8501 (N_8501,N_7348,N_7610);
nor U8502 (N_8502,N_7940,N_7578);
nor U8503 (N_8503,N_7125,N_7193);
nand U8504 (N_8504,N_7603,N_7536);
nand U8505 (N_8505,N_7645,N_7128);
nand U8506 (N_8506,N_7175,N_7686);
nor U8507 (N_8507,N_7747,N_7263);
or U8508 (N_8508,N_7175,N_7440);
nor U8509 (N_8509,N_7443,N_7100);
and U8510 (N_8510,N_7321,N_7627);
xor U8511 (N_8511,N_7591,N_7560);
or U8512 (N_8512,N_7607,N_7360);
or U8513 (N_8513,N_7548,N_7571);
nand U8514 (N_8514,N_7094,N_7197);
nor U8515 (N_8515,N_7833,N_7307);
nand U8516 (N_8516,N_7463,N_7131);
and U8517 (N_8517,N_7981,N_7638);
nand U8518 (N_8518,N_7978,N_7747);
nand U8519 (N_8519,N_7981,N_7523);
and U8520 (N_8520,N_7325,N_7927);
or U8521 (N_8521,N_7233,N_7612);
nand U8522 (N_8522,N_7896,N_7194);
or U8523 (N_8523,N_7309,N_7490);
xnor U8524 (N_8524,N_7160,N_7128);
xnor U8525 (N_8525,N_7258,N_7780);
xnor U8526 (N_8526,N_7220,N_7494);
nor U8527 (N_8527,N_7634,N_7487);
nand U8528 (N_8528,N_7178,N_7076);
xor U8529 (N_8529,N_7098,N_7748);
xnor U8530 (N_8530,N_7055,N_7642);
nor U8531 (N_8531,N_7930,N_7996);
nor U8532 (N_8532,N_7172,N_7624);
nor U8533 (N_8533,N_7080,N_7899);
nand U8534 (N_8534,N_7389,N_7175);
and U8535 (N_8535,N_7195,N_7580);
nand U8536 (N_8536,N_7976,N_7477);
nand U8537 (N_8537,N_7053,N_7503);
or U8538 (N_8538,N_7169,N_7801);
xnor U8539 (N_8539,N_7880,N_7836);
xor U8540 (N_8540,N_7050,N_7421);
nand U8541 (N_8541,N_7520,N_7066);
nand U8542 (N_8542,N_7163,N_7580);
or U8543 (N_8543,N_7375,N_7228);
nor U8544 (N_8544,N_7654,N_7235);
or U8545 (N_8545,N_7914,N_7463);
nor U8546 (N_8546,N_7851,N_7983);
nand U8547 (N_8547,N_7775,N_7296);
and U8548 (N_8548,N_7121,N_7516);
and U8549 (N_8549,N_7603,N_7721);
and U8550 (N_8550,N_7947,N_7245);
nor U8551 (N_8551,N_7890,N_7646);
xor U8552 (N_8552,N_7172,N_7317);
nor U8553 (N_8553,N_7150,N_7246);
nor U8554 (N_8554,N_7546,N_7836);
and U8555 (N_8555,N_7493,N_7561);
nand U8556 (N_8556,N_7971,N_7190);
nor U8557 (N_8557,N_7590,N_7761);
or U8558 (N_8558,N_7853,N_7170);
nor U8559 (N_8559,N_7337,N_7064);
nor U8560 (N_8560,N_7724,N_7760);
nand U8561 (N_8561,N_7647,N_7883);
nand U8562 (N_8562,N_7430,N_7068);
nor U8563 (N_8563,N_7674,N_7453);
nand U8564 (N_8564,N_7536,N_7715);
xor U8565 (N_8565,N_7784,N_7566);
nor U8566 (N_8566,N_7355,N_7828);
xor U8567 (N_8567,N_7653,N_7742);
or U8568 (N_8568,N_7380,N_7708);
and U8569 (N_8569,N_7549,N_7150);
or U8570 (N_8570,N_7547,N_7241);
nand U8571 (N_8571,N_7618,N_7330);
nor U8572 (N_8572,N_7098,N_7019);
nor U8573 (N_8573,N_7969,N_7148);
nor U8574 (N_8574,N_7287,N_7856);
nand U8575 (N_8575,N_7359,N_7968);
and U8576 (N_8576,N_7198,N_7355);
nor U8577 (N_8577,N_7211,N_7950);
xor U8578 (N_8578,N_7611,N_7862);
and U8579 (N_8579,N_7817,N_7517);
or U8580 (N_8580,N_7941,N_7917);
or U8581 (N_8581,N_7172,N_7916);
nand U8582 (N_8582,N_7243,N_7899);
nor U8583 (N_8583,N_7789,N_7995);
nand U8584 (N_8584,N_7657,N_7156);
or U8585 (N_8585,N_7274,N_7604);
nand U8586 (N_8586,N_7837,N_7730);
and U8587 (N_8587,N_7890,N_7209);
or U8588 (N_8588,N_7710,N_7223);
nand U8589 (N_8589,N_7651,N_7321);
or U8590 (N_8590,N_7359,N_7453);
xnor U8591 (N_8591,N_7588,N_7563);
and U8592 (N_8592,N_7740,N_7509);
and U8593 (N_8593,N_7537,N_7036);
and U8594 (N_8594,N_7865,N_7388);
xnor U8595 (N_8595,N_7320,N_7955);
or U8596 (N_8596,N_7791,N_7367);
xor U8597 (N_8597,N_7009,N_7947);
nand U8598 (N_8598,N_7407,N_7760);
nand U8599 (N_8599,N_7596,N_7462);
nor U8600 (N_8600,N_7358,N_7436);
xor U8601 (N_8601,N_7657,N_7807);
and U8602 (N_8602,N_7820,N_7417);
and U8603 (N_8603,N_7217,N_7794);
xor U8604 (N_8604,N_7808,N_7165);
or U8605 (N_8605,N_7679,N_7418);
nand U8606 (N_8606,N_7459,N_7553);
or U8607 (N_8607,N_7399,N_7849);
or U8608 (N_8608,N_7411,N_7599);
or U8609 (N_8609,N_7680,N_7681);
xnor U8610 (N_8610,N_7527,N_7582);
or U8611 (N_8611,N_7468,N_7023);
and U8612 (N_8612,N_7423,N_7017);
nor U8613 (N_8613,N_7390,N_7547);
nand U8614 (N_8614,N_7829,N_7778);
or U8615 (N_8615,N_7745,N_7714);
xnor U8616 (N_8616,N_7943,N_7613);
nor U8617 (N_8617,N_7844,N_7981);
and U8618 (N_8618,N_7010,N_7878);
or U8619 (N_8619,N_7374,N_7905);
nor U8620 (N_8620,N_7801,N_7948);
and U8621 (N_8621,N_7847,N_7891);
or U8622 (N_8622,N_7971,N_7827);
xor U8623 (N_8623,N_7305,N_7889);
or U8624 (N_8624,N_7484,N_7841);
nand U8625 (N_8625,N_7485,N_7943);
and U8626 (N_8626,N_7362,N_7389);
nor U8627 (N_8627,N_7091,N_7049);
xor U8628 (N_8628,N_7141,N_7020);
or U8629 (N_8629,N_7630,N_7330);
nor U8630 (N_8630,N_7697,N_7483);
nand U8631 (N_8631,N_7612,N_7447);
and U8632 (N_8632,N_7026,N_7471);
and U8633 (N_8633,N_7421,N_7427);
and U8634 (N_8634,N_7552,N_7407);
nor U8635 (N_8635,N_7386,N_7967);
nor U8636 (N_8636,N_7008,N_7835);
nor U8637 (N_8637,N_7738,N_7188);
nor U8638 (N_8638,N_7625,N_7118);
nand U8639 (N_8639,N_7336,N_7031);
nand U8640 (N_8640,N_7507,N_7181);
nand U8641 (N_8641,N_7392,N_7040);
and U8642 (N_8642,N_7546,N_7308);
and U8643 (N_8643,N_7658,N_7484);
nand U8644 (N_8644,N_7428,N_7607);
and U8645 (N_8645,N_7303,N_7361);
and U8646 (N_8646,N_7779,N_7492);
or U8647 (N_8647,N_7459,N_7442);
and U8648 (N_8648,N_7403,N_7944);
nand U8649 (N_8649,N_7740,N_7114);
and U8650 (N_8650,N_7448,N_7888);
nor U8651 (N_8651,N_7865,N_7876);
or U8652 (N_8652,N_7794,N_7520);
or U8653 (N_8653,N_7354,N_7832);
and U8654 (N_8654,N_7214,N_7828);
nor U8655 (N_8655,N_7589,N_7433);
xor U8656 (N_8656,N_7660,N_7995);
and U8657 (N_8657,N_7247,N_7714);
nand U8658 (N_8658,N_7052,N_7362);
and U8659 (N_8659,N_7825,N_7892);
and U8660 (N_8660,N_7432,N_7453);
nor U8661 (N_8661,N_7608,N_7752);
nand U8662 (N_8662,N_7629,N_7102);
or U8663 (N_8663,N_7671,N_7422);
or U8664 (N_8664,N_7490,N_7255);
nand U8665 (N_8665,N_7783,N_7875);
nand U8666 (N_8666,N_7575,N_7675);
and U8667 (N_8667,N_7563,N_7407);
nand U8668 (N_8668,N_7896,N_7643);
nand U8669 (N_8669,N_7767,N_7048);
nor U8670 (N_8670,N_7986,N_7488);
nand U8671 (N_8671,N_7735,N_7831);
and U8672 (N_8672,N_7867,N_7342);
or U8673 (N_8673,N_7414,N_7636);
and U8674 (N_8674,N_7048,N_7610);
and U8675 (N_8675,N_7867,N_7156);
nor U8676 (N_8676,N_7496,N_7801);
or U8677 (N_8677,N_7302,N_7617);
or U8678 (N_8678,N_7760,N_7704);
or U8679 (N_8679,N_7521,N_7961);
nor U8680 (N_8680,N_7382,N_7014);
nand U8681 (N_8681,N_7171,N_7358);
nand U8682 (N_8682,N_7673,N_7384);
nor U8683 (N_8683,N_7227,N_7914);
and U8684 (N_8684,N_7390,N_7082);
and U8685 (N_8685,N_7313,N_7396);
nand U8686 (N_8686,N_7457,N_7288);
or U8687 (N_8687,N_7878,N_7172);
nor U8688 (N_8688,N_7703,N_7939);
and U8689 (N_8689,N_7846,N_7582);
nor U8690 (N_8690,N_7675,N_7317);
nor U8691 (N_8691,N_7031,N_7634);
xor U8692 (N_8692,N_7559,N_7720);
nor U8693 (N_8693,N_7784,N_7508);
or U8694 (N_8694,N_7091,N_7250);
xor U8695 (N_8695,N_7662,N_7156);
or U8696 (N_8696,N_7881,N_7392);
nor U8697 (N_8697,N_7550,N_7489);
and U8698 (N_8698,N_7967,N_7067);
or U8699 (N_8699,N_7620,N_7250);
nand U8700 (N_8700,N_7469,N_7441);
or U8701 (N_8701,N_7373,N_7490);
nor U8702 (N_8702,N_7775,N_7271);
and U8703 (N_8703,N_7593,N_7709);
or U8704 (N_8704,N_7806,N_7895);
or U8705 (N_8705,N_7369,N_7174);
and U8706 (N_8706,N_7895,N_7207);
and U8707 (N_8707,N_7450,N_7847);
nor U8708 (N_8708,N_7615,N_7951);
and U8709 (N_8709,N_7147,N_7267);
or U8710 (N_8710,N_7068,N_7564);
or U8711 (N_8711,N_7068,N_7094);
or U8712 (N_8712,N_7574,N_7558);
and U8713 (N_8713,N_7464,N_7478);
xnor U8714 (N_8714,N_7364,N_7164);
nand U8715 (N_8715,N_7541,N_7304);
xnor U8716 (N_8716,N_7510,N_7178);
or U8717 (N_8717,N_7461,N_7945);
or U8718 (N_8718,N_7746,N_7111);
and U8719 (N_8719,N_7624,N_7345);
and U8720 (N_8720,N_7447,N_7214);
nor U8721 (N_8721,N_7144,N_7915);
nor U8722 (N_8722,N_7883,N_7781);
or U8723 (N_8723,N_7720,N_7248);
or U8724 (N_8724,N_7260,N_7713);
nand U8725 (N_8725,N_7477,N_7331);
and U8726 (N_8726,N_7188,N_7293);
nor U8727 (N_8727,N_7066,N_7305);
nor U8728 (N_8728,N_7835,N_7342);
xor U8729 (N_8729,N_7889,N_7592);
or U8730 (N_8730,N_7392,N_7641);
and U8731 (N_8731,N_7244,N_7724);
or U8732 (N_8732,N_7446,N_7880);
or U8733 (N_8733,N_7832,N_7953);
nand U8734 (N_8734,N_7276,N_7831);
or U8735 (N_8735,N_7926,N_7855);
nor U8736 (N_8736,N_7169,N_7105);
xnor U8737 (N_8737,N_7874,N_7067);
nand U8738 (N_8738,N_7295,N_7946);
xnor U8739 (N_8739,N_7109,N_7323);
xor U8740 (N_8740,N_7575,N_7055);
nand U8741 (N_8741,N_7835,N_7214);
nor U8742 (N_8742,N_7163,N_7260);
nand U8743 (N_8743,N_7515,N_7718);
nand U8744 (N_8744,N_7066,N_7989);
or U8745 (N_8745,N_7291,N_7165);
nor U8746 (N_8746,N_7482,N_7496);
and U8747 (N_8747,N_7240,N_7592);
nor U8748 (N_8748,N_7809,N_7554);
or U8749 (N_8749,N_7834,N_7479);
nand U8750 (N_8750,N_7398,N_7516);
nand U8751 (N_8751,N_7976,N_7504);
nand U8752 (N_8752,N_7374,N_7215);
or U8753 (N_8753,N_7589,N_7163);
xnor U8754 (N_8754,N_7670,N_7668);
or U8755 (N_8755,N_7133,N_7680);
and U8756 (N_8756,N_7352,N_7818);
nor U8757 (N_8757,N_7457,N_7081);
or U8758 (N_8758,N_7696,N_7899);
or U8759 (N_8759,N_7894,N_7308);
nor U8760 (N_8760,N_7214,N_7877);
nand U8761 (N_8761,N_7944,N_7776);
or U8762 (N_8762,N_7747,N_7246);
nor U8763 (N_8763,N_7683,N_7967);
nor U8764 (N_8764,N_7370,N_7812);
and U8765 (N_8765,N_7298,N_7973);
and U8766 (N_8766,N_7523,N_7100);
nand U8767 (N_8767,N_7186,N_7135);
nor U8768 (N_8768,N_7917,N_7985);
nand U8769 (N_8769,N_7300,N_7460);
nor U8770 (N_8770,N_7187,N_7258);
nand U8771 (N_8771,N_7599,N_7701);
or U8772 (N_8772,N_7876,N_7059);
and U8773 (N_8773,N_7114,N_7615);
or U8774 (N_8774,N_7472,N_7933);
and U8775 (N_8775,N_7380,N_7000);
or U8776 (N_8776,N_7849,N_7971);
nor U8777 (N_8777,N_7919,N_7430);
and U8778 (N_8778,N_7742,N_7591);
and U8779 (N_8779,N_7276,N_7507);
nor U8780 (N_8780,N_7783,N_7384);
or U8781 (N_8781,N_7322,N_7627);
nand U8782 (N_8782,N_7167,N_7531);
or U8783 (N_8783,N_7373,N_7106);
and U8784 (N_8784,N_7674,N_7649);
and U8785 (N_8785,N_7690,N_7515);
and U8786 (N_8786,N_7166,N_7696);
nand U8787 (N_8787,N_7911,N_7800);
nand U8788 (N_8788,N_7362,N_7151);
nor U8789 (N_8789,N_7608,N_7150);
and U8790 (N_8790,N_7161,N_7811);
nand U8791 (N_8791,N_7216,N_7284);
and U8792 (N_8792,N_7269,N_7774);
or U8793 (N_8793,N_7074,N_7937);
and U8794 (N_8794,N_7147,N_7196);
nor U8795 (N_8795,N_7805,N_7263);
nor U8796 (N_8796,N_7915,N_7548);
nor U8797 (N_8797,N_7270,N_7945);
xnor U8798 (N_8798,N_7178,N_7668);
or U8799 (N_8799,N_7377,N_7436);
nor U8800 (N_8800,N_7174,N_7768);
nand U8801 (N_8801,N_7157,N_7948);
nand U8802 (N_8802,N_7598,N_7990);
nand U8803 (N_8803,N_7680,N_7710);
nand U8804 (N_8804,N_7884,N_7734);
and U8805 (N_8805,N_7479,N_7285);
or U8806 (N_8806,N_7821,N_7733);
nor U8807 (N_8807,N_7368,N_7561);
and U8808 (N_8808,N_7618,N_7216);
or U8809 (N_8809,N_7291,N_7585);
and U8810 (N_8810,N_7749,N_7260);
or U8811 (N_8811,N_7613,N_7734);
xor U8812 (N_8812,N_7874,N_7964);
xnor U8813 (N_8813,N_7453,N_7571);
nand U8814 (N_8814,N_7572,N_7778);
and U8815 (N_8815,N_7020,N_7994);
and U8816 (N_8816,N_7764,N_7110);
nand U8817 (N_8817,N_7814,N_7945);
nor U8818 (N_8818,N_7200,N_7051);
and U8819 (N_8819,N_7577,N_7063);
nand U8820 (N_8820,N_7883,N_7854);
and U8821 (N_8821,N_7242,N_7810);
or U8822 (N_8822,N_7626,N_7740);
xor U8823 (N_8823,N_7631,N_7255);
nor U8824 (N_8824,N_7302,N_7941);
xnor U8825 (N_8825,N_7703,N_7283);
nor U8826 (N_8826,N_7762,N_7886);
or U8827 (N_8827,N_7324,N_7169);
or U8828 (N_8828,N_7117,N_7651);
nand U8829 (N_8829,N_7013,N_7892);
nand U8830 (N_8830,N_7296,N_7890);
nor U8831 (N_8831,N_7739,N_7389);
nor U8832 (N_8832,N_7896,N_7703);
nand U8833 (N_8833,N_7305,N_7003);
or U8834 (N_8834,N_7909,N_7330);
and U8835 (N_8835,N_7559,N_7759);
nor U8836 (N_8836,N_7713,N_7641);
nand U8837 (N_8837,N_7587,N_7322);
and U8838 (N_8838,N_7490,N_7329);
xor U8839 (N_8839,N_7097,N_7588);
or U8840 (N_8840,N_7112,N_7144);
or U8841 (N_8841,N_7582,N_7418);
nand U8842 (N_8842,N_7726,N_7484);
nand U8843 (N_8843,N_7273,N_7817);
xnor U8844 (N_8844,N_7360,N_7029);
and U8845 (N_8845,N_7999,N_7132);
nand U8846 (N_8846,N_7660,N_7226);
and U8847 (N_8847,N_7009,N_7697);
nor U8848 (N_8848,N_7038,N_7452);
and U8849 (N_8849,N_7435,N_7092);
and U8850 (N_8850,N_7234,N_7577);
or U8851 (N_8851,N_7086,N_7113);
nand U8852 (N_8852,N_7404,N_7696);
nand U8853 (N_8853,N_7618,N_7589);
nor U8854 (N_8854,N_7373,N_7057);
or U8855 (N_8855,N_7687,N_7215);
or U8856 (N_8856,N_7236,N_7304);
nand U8857 (N_8857,N_7813,N_7599);
nor U8858 (N_8858,N_7577,N_7313);
nand U8859 (N_8859,N_7276,N_7614);
nand U8860 (N_8860,N_7069,N_7045);
xnor U8861 (N_8861,N_7889,N_7135);
nor U8862 (N_8862,N_7670,N_7675);
and U8863 (N_8863,N_7364,N_7618);
nor U8864 (N_8864,N_7528,N_7983);
and U8865 (N_8865,N_7555,N_7466);
and U8866 (N_8866,N_7542,N_7129);
and U8867 (N_8867,N_7975,N_7159);
and U8868 (N_8868,N_7767,N_7073);
xnor U8869 (N_8869,N_7921,N_7403);
or U8870 (N_8870,N_7778,N_7444);
or U8871 (N_8871,N_7978,N_7483);
or U8872 (N_8872,N_7405,N_7181);
nor U8873 (N_8873,N_7392,N_7528);
or U8874 (N_8874,N_7419,N_7071);
nand U8875 (N_8875,N_7939,N_7376);
nand U8876 (N_8876,N_7079,N_7378);
and U8877 (N_8877,N_7300,N_7418);
or U8878 (N_8878,N_7584,N_7132);
nor U8879 (N_8879,N_7738,N_7673);
and U8880 (N_8880,N_7820,N_7347);
nand U8881 (N_8881,N_7448,N_7973);
and U8882 (N_8882,N_7959,N_7220);
nand U8883 (N_8883,N_7831,N_7315);
or U8884 (N_8884,N_7025,N_7557);
xnor U8885 (N_8885,N_7129,N_7115);
and U8886 (N_8886,N_7032,N_7463);
xor U8887 (N_8887,N_7184,N_7595);
and U8888 (N_8888,N_7704,N_7674);
xor U8889 (N_8889,N_7838,N_7433);
nor U8890 (N_8890,N_7911,N_7656);
nand U8891 (N_8891,N_7176,N_7296);
and U8892 (N_8892,N_7700,N_7840);
nor U8893 (N_8893,N_7687,N_7719);
nand U8894 (N_8894,N_7566,N_7806);
nor U8895 (N_8895,N_7068,N_7997);
nor U8896 (N_8896,N_7630,N_7218);
and U8897 (N_8897,N_7164,N_7972);
nor U8898 (N_8898,N_7792,N_7091);
and U8899 (N_8899,N_7370,N_7201);
or U8900 (N_8900,N_7433,N_7101);
nand U8901 (N_8901,N_7153,N_7880);
nor U8902 (N_8902,N_7794,N_7298);
or U8903 (N_8903,N_7921,N_7586);
nor U8904 (N_8904,N_7621,N_7457);
and U8905 (N_8905,N_7788,N_7801);
nand U8906 (N_8906,N_7675,N_7020);
nand U8907 (N_8907,N_7763,N_7094);
nand U8908 (N_8908,N_7554,N_7807);
nand U8909 (N_8909,N_7015,N_7828);
nand U8910 (N_8910,N_7459,N_7894);
xor U8911 (N_8911,N_7149,N_7617);
nand U8912 (N_8912,N_7684,N_7349);
or U8913 (N_8913,N_7116,N_7760);
nand U8914 (N_8914,N_7529,N_7800);
nand U8915 (N_8915,N_7435,N_7114);
nand U8916 (N_8916,N_7644,N_7267);
or U8917 (N_8917,N_7094,N_7856);
nand U8918 (N_8918,N_7939,N_7778);
nor U8919 (N_8919,N_7449,N_7925);
or U8920 (N_8920,N_7528,N_7371);
nand U8921 (N_8921,N_7344,N_7319);
or U8922 (N_8922,N_7902,N_7810);
nor U8923 (N_8923,N_7379,N_7167);
xor U8924 (N_8924,N_7155,N_7147);
nand U8925 (N_8925,N_7292,N_7375);
nor U8926 (N_8926,N_7290,N_7302);
xnor U8927 (N_8927,N_7628,N_7486);
nand U8928 (N_8928,N_7652,N_7364);
and U8929 (N_8929,N_7512,N_7520);
nand U8930 (N_8930,N_7496,N_7634);
nor U8931 (N_8931,N_7965,N_7449);
xor U8932 (N_8932,N_7273,N_7214);
and U8933 (N_8933,N_7825,N_7833);
xor U8934 (N_8934,N_7644,N_7808);
nand U8935 (N_8935,N_7654,N_7001);
or U8936 (N_8936,N_7290,N_7991);
or U8937 (N_8937,N_7207,N_7492);
nor U8938 (N_8938,N_7207,N_7702);
nor U8939 (N_8939,N_7324,N_7099);
or U8940 (N_8940,N_7101,N_7043);
nand U8941 (N_8941,N_7951,N_7299);
nor U8942 (N_8942,N_7861,N_7146);
nand U8943 (N_8943,N_7114,N_7441);
or U8944 (N_8944,N_7617,N_7651);
nor U8945 (N_8945,N_7975,N_7970);
xnor U8946 (N_8946,N_7012,N_7789);
and U8947 (N_8947,N_7654,N_7718);
nor U8948 (N_8948,N_7294,N_7917);
nor U8949 (N_8949,N_7329,N_7204);
and U8950 (N_8950,N_7390,N_7825);
nand U8951 (N_8951,N_7107,N_7813);
nor U8952 (N_8952,N_7533,N_7969);
and U8953 (N_8953,N_7672,N_7141);
or U8954 (N_8954,N_7535,N_7186);
nand U8955 (N_8955,N_7931,N_7004);
or U8956 (N_8956,N_7131,N_7075);
nand U8957 (N_8957,N_7230,N_7551);
xnor U8958 (N_8958,N_7281,N_7759);
or U8959 (N_8959,N_7245,N_7130);
and U8960 (N_8960,N_7398,N_7411);
nand U8961 (N_8961,N_7927,N_7795);
nand U8962 (N_8962,N_7071,N_7837);
nor U8963 (N_8963,N_7835,N_7924);
and U8964 (N_8964,N_7059,N_7634);
or U8965 (N_8965,N_7622,N_7782);
nor U8966 (N_8966,N_7681,N_7815);
and U8967 (N_8967,N_7126,N_7179);
or U8968 (N_8968,N_7177,N_7970);
or U8969 (N_8969,N_7251,N_7374);
nor U8970 (N_8970,N_7493,N_7294);
and U8971 (N_8971,N_7360,N_7528);
nand U8972 (N_8972,N_7888,N_7864);
nor U8973 (N_8973,N_7509,N_7561);
nand U8974 (N_8974,N_7119,N_7618);
and U8975 (N_8975,N_7323,N_7419);
nor U8976 (N_8976,N_7756,N_7150);
and U8977 (N_8977,N_7227,N_7607);
nor U8978 (N_8978,N_7503,N_7840);
xnor U8979 (N_8979,N_7106,N_7482);
nand U8980 (N_8980,N_7088,N_7479);
or U8981 (N_8981,N_7764,N_7145);
xnor U8982 (N_8982,N_7677,N_7066);
nor U8983 (N_8983,N_7956,N_7338);
xnor U8984 (N_8984,N_7776,N_7117);
nand U8985 (N_8985,N_7482,N_7642);
or U8986 (N_8986,N_7095,N_7274);
xnor U8987 (N_8987,N_7328,N_7146);
or U8988 (N_8988,N_7335,N_7427);
nor U8989 (N_8989,N_7667,N_7873);
nor U8990 (N_8990,N_7741,N_7030);
and U8991 (N_8991,N_7473,N_7904);
and U8992 (N_8992,N_7839,N_7003);
nor U8993 (N_8993,N_7570,N_7635);
nor U8994 (N_8994,N_7018,N_7439);
or U8995 (N_8995,N_7290,N_7759);
or U8996 (N_8996,N_7988,N_7311);
and U8997 (N_8997,N_7592,N_7335);
nand U8998 (N_8998,N_7214,N_7610);
nand U8999 (N_8999,N_7115,N_7936);
nor U9000 (N_9000,N_8019,N_8529);
nand U9001 (N_9001,N_8482,N_8960);
or U9002 (N_9002,N_8064,N_8615);
nor U9003 (N_9003,N_8820,N_8479);
nand U9004 (N_9004,N_8503,N_8212);
nand U9005 (N_9005,N_8800,N_8806);
nand U9006 (N_9006,N_8886,N_8403);
and U9007 (N_9007,N_8786,N_8207);
or U9008 (N_9008,N_8317,N_8091);
nor U9009 (N_9009,N_8430,N_8802);
and U9010 (N_9010,N_8020,N_8156);
and U9011 (N_9011,N_8650,N_8547);
xor U9012 (N_9012,N_8137,N_8050);
nor U9013 (N_9013,N_8121,N_8285);
or U9014 (N_9014,N_8318,N_8898);
nand U9015 (N_9015,N_8413,N_8573);
nor U9016 (N_9016,N_8648,N_8556);
and U9017 (N_9017,N_8376,N_8441);
nor U9018 (N_9018,N_8001,N_8607);
xor U9019 (N_9019,N_8335,N_8257);
nand U9020 (N_9020,N_8688,N_8589);
nor U9021 (N_9021,N_8095,N_8080);
or U9022 (N_9022,N_8689,N_8011);
and U9023 (N_9023,N_8136,N_8971);
xor U9024 (N_9024,N_8400,N_8794);
and U9025 (N_9025,N_8878,N_8591);
and U9026 (N_9026,N_8465,N_8893);
or U9027 (N_9027,N_8172,N_8250);
nand U9028 (N_9028,N_8846,N_8978);
and U9029 (N_9029,N_8005,N_8338);
and U9030 (N_9030,N_8135,N_8296);
nand U9031 (N_9031,N_8033,N_8412);
nand U9032 (N_9032,N_8635,N_8309);
nand U9033 (N_9033,N_8795,N_8475);
and U9034 (N_9034,N_8674,N_8414);
or U9035 (N_9035,N_8041,N_8633);
and U9036 (N_9036,N_8944,N_8558);
and U9037 (N_9037,N_8476,N_8670);
nor U9038 (N_9038,N_8518,N_8507);
or U9039 (N_9039,N_8961,N_8662);
xnor U9040 (N_9040,N_8779,N_8983);
and U9041 (N_9041,N_8949,N_8423);
nor U9042 (N_9042,N_8473,N_8532);
nand U9043 (N_9043,N_8625,N_8941);
and U9044 (N_9044,N_8762,N_8667);
or U9045 (N_9045,N_8323,N_8066);
nand U9046 (N_9046,N_8189,N_8557);
nand U9047 (N_9047,N_8551,N_8147);
and U9048 (N_9048,N_8138,N_8994);
nor U9049 (N_9049,N_8314,N_8459);
nand U9050 (N_9050,N_8218,N_8866);
nand U9051 (N_9051,N_8942,N_8491);
and U9052 (N_9052,N_8478,N_8108);
or U9053 (N_9053,N_8014,N_8924);
nor U9054 (N_9054,N_8833,N_8882);
nand U9055 (N_9055,N_8930,N_8153);
or U9056 (N_9056,N_8398,N_8406);
nand U9057 (N_9057,N_8493,N_8322);
nand U9058 (N_9058,N_8399,N_8577);
nand U9059 (N_9059,N_8624,N_8150);
nor U9060 (N_9060,N_8817,N_8467);
or U9061 (N_9061,N_8791,N_8756);
or U9062 (N_9062,N_8197,N_8186);
xnor U9063 (N_9063,N_8010,N_8916);
and U9064 (N_9064,N_8098,N_8954);
xor U9065 (N_9065,N_8517,N_8977);
nand U9066 (N_9066,N_8142,N_8238);
xnor U9067 (N_9067,N_8454,N_8235);
and U9068 (N_9068,N_8416,N_8282);
or U9069 (N_9069,N_8899,N_8021);
and U9070 (N_9070,N_8735,N_8139);
or U9071 (N_9071,N_8696,N_8592);
and U9072 (N_9072,N_8443,N_8658);
and U9073 (N_9073,N_8720,N_8274);
nor U9074 (N_9074,N_8373,N_8939);
nand U9075 (N_9075,N_8222,N_8788);
nand U9076 (N_9076,N_8940,N_8120);
nor U9077 (N_9077,N_8361,N_8740);
nand U9078 (N_9078,N_8643,N_8051);
nand U9079 (N_9079,N_8700,N_8495);
nor U9080 (N_9080,N_8884,N_8769);
nor U9081 (N_9081,N_8901,N_8713);
or U9082 (N_9082,N_8703,N_8328);
nand U9083 (N_9083,N_8126,N_8140);
nor U9084 (N_9084,N_8370,N_8075);
nand U9085 (N_9085,N_8260,N_8044);
or U9086 (N_9086,N_8289,N_8492);
and U9087 (N_9087,N_8654,N_8773);
or U9088 (N_9088,N_8436,N_8783);
nand U9089 (N_9089,N_8819,N_8524);
nand U9090 (N_9090,N_8921,N_8669);
nor U9091 (N_9091,N_8234,N_8319);
and U9092 (N_9092,N_8141,N_8683);
or U9093 (N_9093,N_8923,N_8796);
or U9094 (N_9094,N_8502,N_8391);
and U9095 (N_9095,N_8256,N_8526);
or U9096 (N_9096,N_8588,N_8000);
nor U9097 (N_9097,N_8022,N_8247);
xor U9098 (N_9098,N_8426,N_8088);
and U9099 (N_9099,N_8745,N_8811);
and U9100 (N_9100,N_8619,N_8856);
and U9101 (N_9101,N_8191,N_8099);
or U9102 (N_9102,N_8841,N_8448);
or U9103 (N_9103,N_8341,N_8251);
and U9104 (N_9104,N_8254,N_8867);
or U9105 (N_9105,N_8934,N_8550);
or U9106 (N_9106,N_8455,N_8178);
nor U9107 (N_9107,N_8089,N_8754);
nor U9108 (N_9108,N_8849,N_8008);
nor U9109 (N_9109,N_8598,N_8936);
nand U9110 (N_9110,N_8312,N_8621);
and U9111 (N_9111,N_8082,N_8638);
xnor U9112 (N_9112,N_8776,N_8928);
or U9113 (N_9113,N_8931,N_8876);
or U9114 (N_9114,N_8175,N_8986);
nand U9115 (N_9115,N_8634,N_8469);
and U9116 (N_9116,N_8881,N_8687);
nor U9117 (N_9117,N_8673,N_8110);
nand U9118 (N_9118,N_8836,N_8225);
xnor U9119 (N_9119,N_8699,N_8292);
and U9120 (N_9120,N_8221,N_8715);
nor U9121 (N_9121,N_8750,N_8723);
and U9122 (N_9122,N_8027,N_8204);
nor U9123 (N_9123,N_8891,N_8678);
nand U9124 (N_9124,N_8324,N_8626);
nand U9125 (N_9125,N_8728,N_8821);
xor U9126 (N_9126,N_8716,N_8685);
nand U9127 (N_9127,N_8052,N_8964);
and U9128 (N_9128,N_8917,N_8585);
nand U9129 (N_9129,N_8780,N_8616);
or U9130 (N_9130,N_8872,N_8451);
and U9131 (N_9131,N_8976,N_8392);
or U9132 (N_9132,N_8599,N_8636);
nand U9133 (N_9133,N_8239,N_8329);
or U9134 (N_9134,N_8970,N_8693);
nand U9135 (N_9135,N_8261,N_8902);
nor U9136 (N_9136,N_8013,N_8540);
and U9137 (N_9137,N_8536,N_8488);
and U9138 (N_9138,N_8060,N_8367);
or U9139 (N_9139,N_8885,N_8539);
and U9140 (N_9140,N_8736,N_8071);
and U9141 (N_9141,N_8704,N_8632);
xnor U9142 (N_9142,N_8365,N_8957);
xor U9143 (N_9143,N_8049,N_8107);
xnor U9144 (N_9144,N_8070,N_8613);
nand U9145 (N_9145,N_8900,N_8490);
nand U9146 (N_9146,N_8321,N_8462);
xor U9147 (N_9147,N_8340,N_8894);
and U9148 (N_9148,N_8439,N_8216);
xor U9149 (N_9149,N_8345,N_8926);
and U9150 (N_9150,N_8533,N_8920);
nor U9151 (N_9151,N_8999,N_8727);
and U9152 (N_9152,N_8384,N_8982);
or U9153 (N_9153,N_8183,N_8032);
nor U9154 (N_9154,N_8283,N_8313);
nand U9155 (N_9155,N_8004,N_8838);
or U9156 (N_9156,N_8668,N_8804);
and U9157 (N_9157,N_8170,N_8009);
or U9158 (N_9158,N_8372,N_8036);
nor U9159 (N_9159,N_8094,N_8530);
xnor U9160 (N_9160,N_8695,N_8602);
nand U9161 (N_9161,N_8415,N_8908);
nor U9162 (N_9162,N_8404,N_8103);
nand U9163 (N_9163,N_8694,N_8143);
or U9164 (N_9164,N_8746,N_8336);
nor U9165 (N_9165,N_8311,N_8040);
or U9166 (N_9166,N_8741,N_8357);
and U9167 (N_9167,N_8584,N_8061);
xnor U9168 (N_9168,N_8243,N_8093);
xor U9169 (N_9169,N_8481,N_8790);
nand U9170 (N_9170,N_8664,N_8100);
and U9171 (N_9171,N_8927,N_8549);
and U9172 (N_9172,N_8435,N_8951);
and U9173 (N_9173,N_8355,N_8277);
nand U9174 (N_9174,N_8732,N_8755);
and U9175 (N_9175,N_8179,N_8586);
nand U9176 (N_9176,N_8768,N_8701);
nor U9177 (N_9177,N_8113,N_8686);
and U9178 (N_9178,N_8035,N_8055);
or U9179 (N_9179,N_8171,N_8677);
or U9180 (N_9180,N_8752,N_8822);
and U9181 (N_9181,N_8571,N_8155);
nand U9182 (N_9182,N_8937,N_8209);
or U9183 (N_9183,N_8269,N_8470);
nor U9184 (N_9184,N_8028,N_8538);
and U9185 (N_9185,N_8227,N_8631);
nand U9186 (N_9186,N_8220,N_8965);
nor U9187 (N_9187,N_8839,N_8609);
nand U9188 (N_9188,N_8590,N_8639);
xnor U9189 (N_9189,N_8241,N_8017);
nor U9190 (N_9190,N_8883,N_8386);
nand U9191 (N_9191,N_8515,N_8346);
or U9192 (N_9192,N_8874,N_8935);
nor U9193 (N_9193,N_8118,N_8682);
xnor U9194 (N_9194,N_8764,N_8763);
nand U9195 (N_9195,N_8180,N_8500);
or U9196 (N_9196,N_8114,N_8188);
xor U9197 (N_9197,N_8237,N_8904);
nor U9198 (N_9198,N_8043,N_8684);
xnor U9199 (N_9199,N_8047,N_8166);
and U9200 (N_9200,N_8045,N_8531);
or U9201 (N_9201,N_8486,N_8730);
and U9202 (N_9202,N_8992,N_8984);
nand U9203 (N_9203,N_8460,N_8434);
nand U9204 (N_9204,N_8306,N_8279);
nor U9205 (N_9205,N_8829,N_8054);
nand U9206 (N_9206,N_8496,N_8554);
nand U9207 (N_9207,N_8661,N_8985);
and U9208 (N_9208,N_8056,N_8253);
nor U9209 (N_9209,N_8919,N_8331);
xor U9210 (N_9210,N_8561,N_8205);
or U9211 (N_9211,N_8182,N_8038);
xor U9212 (N_9212,N_8844,N_8990);
nor U9213 (N_9213,N_8302,N_8339);
and U9214 (N_9214,N_8078,N_8840);
and U9215 (N_9215,N_8947,N_8544);
and U9216 (N_9216,N_8378,N_8215);
and U9217 (N_9217,N_8692,N_8062);
xor U9218 (N_9218,N_8363,N_8437);
or U9219 (N_9219,N_8697,N_8226);
nand U9220 (N_9220,N_8420,N_8909);
or U9221 (N_9221,N_8086,N_8158);
xor U9222 (N_9222,N_8721,N_8981);
xnor U9223 (N_9223,N_8417,N_8897);
nand U9224 (N_9224,N_8382,N_8498);
xnor U9225 (N_9225,N_8301,N_8287);
and U9226 (N_9226,N_8512,N_8154);
or U9227 (N_9227,N_8611,N_8514);
nor U9228 (N_9228,N_8691,N_8905);
and U9229 (N_9229,N_8641,N_8761);
xnor U9230 (N_9230,N_8812,N_8711);
nand U9231 (N_9231,N_8003,N_8758);
or U9232 (N_9232,N_8578,N_8456);
nor U9233 (N_9233,N_8039,N_8892);
or U9234 (N_9234,N_8548,N_8831);
xnor U9235 (N_9235,N_8782,N_8474);
xnor U9236 (N_9236,N_8160,N_8480);
and U9237 (N_9237,N_8722,N_8652);
nor U9238 (N_9238,N_8268,N_8115);
or U9239 (N_9239,N_8858,N_8046);
nor U9240 (N_9240,N_8411,N_8079);
nor U9241 (N_9241,N_8824,N_8332);
or U9242 (N_9242,N_8063,N_8431);
and U9243 (N_9243,N_8195,N_8489);
nand U9244 (N_9244,N_8427,N_8042);
or U9245 (N_9245,N_8472,N_8593);
nor U9246 (N_9246,N_8162,N_8265);
or U9247 (N_9247,N_8570,N_8203);
or U9248 (N_9248,N_8401,N_8208);
xor U9249 (N_9249,N_8127,N_8012);
nand U9250 (N_9250,N_8176,N_8288);
and U9251 (N_9251,N_8354,N_8105);
nor U9252 (N_9252,N_8211,N_8381);
nor U9253 (N_9253,N_8871,N_8968);
nor U9254 (N_9254,N_8785,N_8863);
nand U9255 (N_9255,N_8709,N_8825);
nor U9256 (N_9256,N_8604,N_8334);
and U9257 (N_9257,N_8527,N_8869);
or U9258 (N_9258,N_8830,N_8672);
or U9259 (N_9259,N_8383,N_8255);
nor U9260 (N_9260,N_8397,N_8092);
and U9261 (N_9261,N_8083,N_8865);
nand U9262 (N_9262,N_8366,N_8574);
nand U9263 (N_9263,N_8537,N_8975);
or U9264 (N_9264,N_8501,N_8772);
or U9265 (N_9265,N_8666,N_8980);
xnor U9266 (N_9266,N_8177,N_8903);
and U9267 (N_9267,N_8958,N_8076);
nor U9268 (N_9268,N_8375,N_8006);
or U9269 (N_9269,N_8352,N_8133);
nor U9270 (N_9270,N_8655,N_8167);
nor U9271 (N_9271,N_8124,N_8390);
xnor U9272 (N_9272,N_8729,N_8873);
or U9273 (N_9273,N_8326,N_8181);
nand U9274 (N_9274,N_8813,N_8997);
or U9275 (N_9275,N_8775,N_8291);
nand U9276 (N_9276,N_8304,N_8974);
and U9277 (N_9277,N_8660,N_8955);
xor U9278 (N_9278,N_8199,N_8396);
or U9279 (N_9279,N_8766,N_8647);
or U9280 (N_9280,N_8466,N_8429);
nor U9281 (N_9281,N_8708,N_8680);
nand U9282 (N_9282,N_8037,N_8534);
nand U9283 (N_9283,N_8031,N_8349);
and U9284 (N_9284,N_8284,N_8030);
or U9285 (N_9285,N_8966,N_8827);
nor U9286 (N_9286,N_8351,N_8065);
nand U9287 (N_9287,N_8552,N_8575);
nand U9288 (N_9288,N_8316,N_8508);
nand U9289 (N_9289,N_8911,N_8485);
or U9290 (N_9290,N_8676,N_8567);
nand U9291 (N_9291,N_8294,N_8069);
nor U9292 (N_9292,N_8198,N_8712);
and U9293 (N_9293,N_8048,N_8690);
xnor U9294 (N_9294,N_8330,N_8275);
or U9295 (N_9295,N_8249,N_8428);
or U9296 (N_9296,N_8244,N_8146);
and U9297 (N_9297,N_8950,N_8477);
or U9298 (N_9298,N_8808,N_8151);
or U9299 (N_9299,N_8228,N_8096);
nor U9300 (N_9300,N_8513,N_8369);
or U9301 (N_9301,N_8068,N_8998);
nor U9302 (N_9302,N_8337,N_8025);
and U9303 (N_9303,N_8077,N_8603);
or U9304 (N_9304,N_8963,N_8327);
or U9305 (N_9305,N_8353,N_8224);
and U9306 (N_9306,N_8023,N_8267);
nor U9307 (N_9307,N_8714,N_8572);
nor U9308 (N_9308,N_8457,N_8608);
xnor U9309 (N_9309,N_8281,N_8810);
xnor U9310 (N_9310,N_8751,N_8938);
xnor U9311 (N_9311,N_8545,N_8563);
and U9312 (N_9312,N_8286,N_8645);
or U9313 (N_9313,N_8315,N_8956);
nor U9314 (N_9314,N_8174,N_8418);
and U9315 (N_9315,N_8343,N_8348);
nand U9316 (N_9316,N_8159,N_8018);
nand U9317 (N_9317,N_8620,N_8972);
and U9318 (N_9318,N_8850,N_8359);
nor U9319 (N_9319,N_8895,N_8471);
xor U9320 (N_9320,N_8259,N_8333);
and U9321 (N_9321,N_8562,N_8360);
nor U9322 (N_9322,N_8217,N_8959);
nor U9323 (N_9323,N_8059,N_8236);
nor U9324 (N_9324,N_8628,N_8067);
or U9325 (N_9325,N_8444,N_8681);
and U9326 (N_9326,N_8637,N_8523);
nor U9327 (N_9327,N_8272,N_8362);
and U9328 (N_9328,N_8263,N_8432);
nand U9329 (N_9329,N_8494,N_8717);
or U9330 (N_9330,N_8053,N_8163);
nor U9331 (N_9331,N_8854,N_8101);
and U9332 (N_9332,N_8542,N_8646);
xnor U9333 (N_9333,N_8541,N_8425);
nand U9334 (N_9334,N_8803,N_8629);
xor U9335 (N_9335,N_8969,N_8622);
nor U9336 (N_9336,N_8487,N_8525);
nor U9337 (N_9337,N_8845,N_8387);
or U9338 (N_9338,N_8057,N_8072);
xnor U9339 (N_9339,N_8298,N_8168);
or U9340 (N_9340,N_8879,N_8112);
xor U9341 (N_9341,N_8600,N_8553);
or U9342 (N_9342,N_8568,N_8748);
nor U9343 (N_9343,N_8910,N_8857);
nor U9344 (N_9344,N_8152,N_8605);
and U9345 (N_9345,N_8380,N_8617);
xor U9346 (N_9346,N_8771,N_8521);
nor U9347 (N_9347,N_8266,N_8297);
and U9348 (N_9348,N_8202,N_8358);
nand U9349 (N_9349,N_8623,N_8445);
or U9350 (N_9350,N_8388,N_8371);
or U9351 (N_9351,N_8122,N_8698);
nor U9352 (N_9352,N_8596,N_8555);
nand U9353 (N_9353,N_8506,N_8516);
nor U9354 (N_9354,N_8424,N_8979);
nand U9355 (N_9355,N_8201,N_8580);
nor U9356 (N_9356,N_8194,N_8085);
xnor U9357 (N_9357,N_8601,N_8024);
nor U9358 (N_9358,N_8084,N_8889);
nor U9359 (N_9359,N_8913,N_8410);
or U9360 (N_9360,N_8859,N_8393);
nand U9361 (N_9361,N_8461,N_8757);
nor U9362 (N_9362,N_8509,N_8657);
xor U9363 (N_9363,N_8438,N_8325);
and U9364 (N_9364,N_8743,N_8111);
and U9365 (N_9365,N_8952,N_8246);
nor U9366 (N_9366,N_8742,N_8123);
xnor U9367 (N_9367,N_8356,N_8058);
and U9368 (N_9368,N_8912,N_8861);
nand U9369 (N_9369,N_8193,N_8967);
and U9370 (N_9370,N_8777,N_8187);
nor U9371 (N_9371,N_8446,N_8814);
and U9372 (N_9372,N_8102,N_8864);
nor U9373 (N_9373,N_8546,N_8770);
nand U9374 (N_9374,N_8165,N_8164);
nor U9375 (N_9375,N_8468,N_8271);
nor U9376 (N_9376,N_8733,N_8922);
xnor U9377 (N_9377,N_8875,N_8989);
nor U9378 (N_9378,N_8344,N_8258);
xnor U9379 (N_9379,N_8368,N_8364);
nand U9380 (N_9380,N_8774,N_8656);
nand U9381 (N_9381,N_8851,N_8389);
nand U9382 (N_9382,N_8737,N_8834);
or U9383 (N_9383,N_8200,N_8242);
nand U9384 (N_9384,N_8823,N_8993);
nand U9385 (N_9385,N_8131,N_8528);
nand U9386 (N_9386,N_8350,N_8097);
or U9387 (N_9387,N_8767,N_8706);
and U9388 (N_9388,N_8837,N_8948);
and U9389 (N_9389,N_8996,N_8644);
nor U9390 (N_9390,N_8106,N_8442);
nor U9391 (N_9391,N_8447,N_8962);
or U9392 (N_9392,N_8034,N_8248);
and U9393 (N_9393,N_8073,N_8002);
nand U9394 (N_9394,N_8015,N_8125);
xor U9395 (N_9395,N_8305,N_8781);
and U9396 (N_9396,N_8145,N_8738);
and U9397 (N_9397,N_8579,N_8792);
or U9398 (N_9398,N_8347,N_8449);
and U9399 (N_9399,N_8233,N_8510);
nor U9400 (N_9400,N_8918,N_8805);
and U9401 (N_9401,N_8848,N_8231);
nand U9402 (N_9402,N_8230,N_8262);
nor U9403 (N_9403,N_8214,N_8877);
nand U9404 (N_9404,N_8801,N_8835);
or U9405 (N_9405,N_8219,N_8890);
nor U9406 (N_9406,N_8651,N_8206);
nand U9407 (N_9407,N_8973,N_8725);
xor U9408 (N_9408,N_8295,N_8280);
nor U9409 (N_9409,N_8169,N_8148);
and U9410 (N_9410,N_8119,N_8760);
and U9411 (N_9411,N_8270,N_8724);
nor U9412 (N_9412,N_8659,N_8653);
and U9413 (N_9413,N_8310,N_8734);
and U9414 (N_9414,N_8559,N_8594);
and U9415 (N_9415,N_8987,N_8753);
nor U9416 (N_9416,N_8452,N_8190);
or U9417 (N_9417,N_8988,N_8818);
nand U9418 (N_9418,N_8229,N_8192);
or U9419 (N_9419,N_8815,N_8026);
nand U9420 (N_9420,N_8303,N_8320);
xnor U9421 (N_9421,N_8842,N_8421);
and U9422 (N_9422,N_8852,N_8293);
or U9423 (N_9423,N_8299,N_8870);
and U9424 (N_9424,N_8793,N_8029);
and U9425 (N_9425,N_8484,N_8679);
and U9426 (N_9426,N_8290,N_8116);
nand U9427 (N_9427,N_8453,N_8543);
nor U9428 (N_9428,N_8307,N_8915);
and U9429 (N_9429,N_8535,N_8587);
and U9430 (N_9430,N_8196,N_8744);
or U9431 (N_9431,N_8618,N_8953);
and U9432 (N_9432,N_8374,N_8847);
nor U9433 (N_9433,N_8185,N_8377);
nor U9434 (N_9434,N_8798,N_8109);
and U9435 (N_9435,N_8896,N_8497);
or U9436 (N_9436,N_8583,N_8522);
or U9437 (N_9437,N_8627,N_8419);
nand U9438 (N_9438,N_8173,N_8184);
nand U9439 (N_9439,N_8134,N_8104);
nor U9440 (N_9440,N_8929,N_8278);
or U9441 (N_9441,N_8395,N_8519);
and U9442 (N_9442,N_8862,N_8582);
nand U9443 (N_9443,N_8614,N_8925);
xnor U9444 (N_9444,N_8799,N_8499);
nand U9445 (N_9445,N_8880,N_8422);
and U9446 (N_9446,N_8707,N_8149);
nor U9447 (N_9447,N_8843,N_8807);
or U9448 (N_9448,N_8932,N_8906);
nand U9449 (N_9449,N_8232,N_8264);
nor U9450 (N_9450,N_8784,N_8665);
or U9451 (N_9451,N_8749,N_8649);
or U9452 (N_9452,N_8759,N_8907);
nor U9453 (N_9453,N_8560,N_8300);
or U9454 (N_9454,N_8765,N_8464);
or U9455 (N_9455,N_8450,N_8081);
nor U9456 (N_9456,N_8565,N_8705);
nor U9457 (N_9457,N_8308,N_8245);
nor U9458 (N_9458,N_8710,N_8797);
nor U9459 (N_9459,N_8273,N_8610);
or U9460 (N_9460,N_8853,N_8074);
or U9461 (N_9461,N_8157,N_8210);
and U9462 (N_9462,N_8991,N_8569);
nor U9463 (N_9463,N_8402,N_8809);
and U9464 (N_9464,N_8630,N_8566);
nor U9465 (N_9465,N_8828,N_8252);
nor U9466 (N_9466,N_8995,N_8090);
and U9467 (N_9467,N_8161,N_8379);
and U9468 (N_9468,N_8511,N_8888);
nor U9469 (N_9469,N_8789,N_8130);
or U9470 (N_9470,N_8826,N_8606);
or U9471 (N_9471,N_8597,N_8887);
and U9472 (N_9472,N_8117,N_8576);
nand U9473 (N_9473,N_8394,N_8946);
and U9474 (N_9474,N_8144,N_8440);
nand U9475 (N_9475,N_8458,N_8855);
or U9476 (N_9476,N_8213,N_8671);
and U9477 (N_9477,N_8816,N_8612);
and U9478 (N_9478,N_8832,N_8505);
and U9479 (N_9479,N_8016,N_8719);
nor U9480 (N_9480,N_8385,N_8408);
xor U9481 (N_9481,N_8778,N_8132);
or U9482 (N_9482,N_8087,N_8520);
nand U9483 (N_9483,N_8914,N_8564);
nand U9484 (N_9484,N_8702,N_8483);
xnor U9485 (N_9485,N_8433,N_8675);
or U9486 (N_9486,N_8581,N_8128);
and U9487 (N_9487,N_8739,N_8595);
nand U9488 (N_9488,N_8407,N_8731);
and U9489 (N_9489,N_8463,N_8933);
or U9490 (N_9490,N_8409,N_8342);
or U9491 (N_9491,N_8747,N_8642);
nor U9492 (N_9492,N_8276,N_8663);
xor U9493 (N_9493,N_8405,N_8223);
nand U9494 (N_9494,N_8007,N_8945);
or U9495 (N_9495,N_8129,N_8860);
and U9496 (N_9496,N_8240,N_8943);
nand U9497 (N_9497,N_8868,N_8504);
and U9498 (N_9498,N_8718,N_8726);
nand U9499 (N_9499,N_8640,N_8787);
nor U9500 (N_9500,N_8532,N_8054);
xor U9501 (N_9501,N_8555,N_8449);
nand U9502 (N_9502,N_8041,N_8947);
or U9503 (N_9503,N_8659,N_8853);
nor U9504 (N_9504,N_8489,N_8290);
or U9505 (N_9505,N_8245,N_8942);
xor U9506 (N_9506,N_8795,N_8768);
nor U9507 (N_9507,N_8300,N_8524);
nand U9508 (N_9508,N_8440,N_8497);
nand U9509 (N_9509,N_8379,N_8144);
xnor U9510 (N_9510,N_8897,N_8081);
nor U9511 (N_9511,N_8262,N_8987);
xor U9512 (N_9512,N_8255,N_8826);
and U9513 (N_9513,N_8371,N_8348);
xnor U9514 (N_9514,N_8323,N_8727);
and U9515 (N_9515,N_8875,N_8502);
nor U9516 (N_9516,N_8852,N_8742);
or U9517 (N_9517,N_8362,N_8202);
and U9518 (N_9518,N_8009,N_8094);
and U9519 (N_9519,N_8590,N_8043);
xor U9520 (N_9520,N_8218,N_8432);
or U9521 (N_9521,N_8819,N_8966);
and U9522 (N_9522,N_8734,N_8989);
or U9523 (N_9523,N_8926,N_8061);
nand U9524 (N_9524,N_8730,N_8562);
and U9525 (N_9525,N_8600,N_8706);
nor U9526 (N_9526,N_8552,N_8120);
nor U9527 (N_9527,N_8396,N_8561);
nor U9528 (N_9528,N_8694,N_8991);
nor U9529 (N_9529,N_8182,N_8841);
nand U9530 (N_9530,N_8596,N_8072);
xnor U9531 (N_9531,N_8481,N_8467);
nor U9532 (N_9532,N_8832,N_8303);
xor U9533 (N_9533,N_8264,N_8273);
xor U9534 (N_9534,N_8705,N_8804);
nand U9535 (N_9535,N_8189,N_8593);
nor U9536 (N_9536,N_8545,N_8189);
nand U9537 (N_9537,N_8296,N_8551);
nand U9538 (N_9538,N_8527,N_8107);
nand U9539 (N_9539,N_8269,N_8790);
or U9540 (N_9540,N_8931,N_8151);
or U9541 (N_9541,N_8930,N_8514);
and U9542 (N_9542,N_8519,N_8405);
and U9543 (N_9543,N_8540,N_8364);
or U9544 (N_9544,N_8467,N_8538);
or U9545 (N_9545,N_8576,N_8839);
and U9546 (N_9546,N_8111,N_8079);
and U9547 (N_9547,N_8498,N_8288);
or U9548 (N_9548,N_8517,N_8542);
nor U9549 (N_9549,N_8873,N_8695);
nor U9550 (N_9550,N_8918,N_8887);
nand U9551 (N_9551,N_8010,N_8432);
or U9552 (N_9552,N_8367,N_8477);
xor U9553 (N_9553,N_8447,N_8021);
nor U9554 (N_9554,N_8025,N_8047);
nand U9555 (N_9555,N_8757,N_8391);
nand U9556 (N_9556,N_8115,N_8087);
nand U9557 (N_9557,N_8861,N_8092);
and U9558 (N_9558,N_8996,N_8435);
nand U9559 (N_9559,N_8869,N_8716);
and U9560 (N_9560,N_8358,N_8551);
or U9561 (N_9561,N_8441,N_8189);
nand U9562 (N_9562,N_8341,N_8169);
nand U9563 (N_9563,N_8128,N_8882);
nand U9564 (N_9564,N_8784,N_8371);
nand U9565 (N_9565,N_8398,N_8413);
or U9566 (N_9566,N_8951,N_8753);
and U9567 (N_9567,N_8581,N_8272);
or U9568 (N_9568,N_8060,N_8752);
and U9569 (N_9569,N_8393,N_8778);
nand U9570 (N_9570,N_8997,N_8539);
nand U9571 (N_9571,N_8166,N_8652);
and U9572 (N_9572,N_8630,N_8308);
nor U9573 (N_9573,N_8698,N_8085);
nor U9574 (N_9574,N_8965,N_8448);
nor U9575 (N_9575,N_8349,N_8678);
or U9576 (N_9576,N_8723,N_8565);
or U9577 (N_9577,N_8632,N_8582);
nor U9578 (N_9578,N_8464,N_8239);
nand U9579 (N_9579,N_8900,N_8269);
and U9580 (N_9580,N_8831,N_8476);
nand U9581 (N_9581,N_8048,N_8161);
or U9582 (N_9582,N_8054,N_8994);
and U9583 (N_9583,N_8358,N_8641);
nand U9584 (N_9584,N_8794,N_8192);
or U9585 (N_9585,N_8466,N_8628);
or U9586 (N_9586,N_8816,N_8362);
nor U9587 (N_9587,N_8222,N_8595);
or U9588 (N_9588,N_8941,N_8305);
nor U9589 (N_9589,N_8767,N_8268);
nor U9590 (N_9590,N_8119,N_8187);
or U9591 (N_9591,N_8606,N_8994);
nand U9592 (N_9592,N_8955,N_8399);
nand U9593 (N_9593,N_8817,N_8524);
nor U9594 (N_9594,N_8821,N_8855);
and U9595 (N_9595,N_8670,N_8776);
and U9596 (N_9596,N_8796,N_8222);
nand U9597 (N_9597,N_8715,N_8311);
nor U9598 (N_9598,N_8759,N_8929);
nand U9599 (N_9599,N_8299,N_8408);
nand U9600 (N_9600,N_8030,N_8820);
or U9601 (N_9601,N_8063,N_8041);
nand U9602 (N_9602,N_8774,N_8000);
or U9603 (N_9603,N_8041,N_8339);
xor U9604 (N_9604,N_8541,N_8505);
nor U9605 (N_9605,N_8763,N_8819);
nor U9606 (N_9606,N_8422,N_8556);
or U9607 (N_9607,N_8312,N_8981);
xor U9608 (N_9608,N_8582,N_8677);
nand U9609 (N_9609,N_8221,N_8296);
or U9610 (N_9610,N_8075,N_8419);
nand U9611 (N_9611,N_8554,N_8548);
nor U9612 (N_9612,N_8301,N_8764);
and U9613 (N_9613,N_8882,N_8395);
nand U9614 (N_9614,N_8093,N_8088);
nand U9615 (N_9615,N_8667,N_8334);
and U9616 (N_9616,N_8040,N_8854);
or U9617 (N_9617,N_8911,N_8747);
or U9618 (N_9618,N_8426,N_8841);
nor U9619 (N_9619,N_8130,N_8007);
xnor U9620 (N_9620,N_8187,N_8799);
nor U9621 (N_9621,N_8433,N_8019);
nand U9622 (N_9622,N_8209,N_8135);
nor U9623 (N_9623,N_8733,N_8845);
and U9624 (N_9624,N_8742,N_8146);
nand U9625 (N_9625,N_8540,N_8733);
xor U9626 (N_9626,N_8691,N_8997);
xor U9627 (N_9627,N_8226,N_8571);
nand U9628 (N_9628,N_8213,N_8720);
and U9629 (N_9629,N_8775,N_8278);
nor U9630 (N_9630,N_8579,N_8933);
or U9631 (N_9631,N_8749,N_8385);
nor U9632 (N_9632,N_8078,N_8097);
nor U9633 (N_9633,N_8474,N_8625);
and U9634 (N_9634,N_8829,N_8718);
xor U9635 (N_9635,N_8645,N_8031);
or U9636 (N_9636,N_8303,N_8300);
and U9637 (N_9637,N_8679,N_8526);
nor U9638 (N_9638,N_8731,N_8061);
or U9639 (N_9639,N_8232,N_8996);
nand U9640 (N_9640,N_8616,N_8276);
nor U9641 (N_9641,N_8216,N_8501);
or U9642 (N_9642,N_8420,N_8426);
nor U9643 (N_9643,N_8292,N_8294);
or U9644 (N_9644,N_8290,N_8009);
or U9645 (N_9645,N_8212,N_8857);
and U9646 (N_9646,N_8019,N_8637);
nor U9647 (N_9647,N_8905,N_8741);
or U9648 (N_9648,N_8312,N_8278);
or U9649 (N_9649,N_8671,N_8312);
nand U9650 (N_9650,N_8182,N_8142);
or U9651 (N_9651,N_8298,N_8807);
and U9652 (N_9652,N_8451,N_8121);
nand U9653 (N_9653,N_8310,N_8809);
xnor U9654 (N_9654,N_8377,N_8407);
nand U9655 (N_9655,N_8638,N_8646);
xnor U9656 (N_9656,N_8004,N_8902);
nor U9657 (N_9657,N_8202,N_8218);
xor U9658 (N_9658,N_8357,N_8185);
nand U9659 (N_9659,N_8711,N_8488);
and U9660 (N_9660,N_8110,N_8722);
nor U9661 (N_9661,N_8698,N_8096);
or U9662 (N_9662,N_8538,N_8939);
and U9663 (N_9663,N_8737,N_8170);
nor U9664 (N_9664,N_8965,N_8841);
xor U9665 (N_9665,N_8706,N_8918);
nor U9666 (N_9666,N_8469,N_8446);
xor U9667 (N_9667,N_8777,N_8516);
or U9668 (N_9668,N_8677,N_8727);
or U9669 (N_9669,N_8528,N_8288);
xor U9670 (N_9670,N_8354,N_8441);
or U9671 (N_9671,N_8261,N_8155);
and U9672 (N_9672,N_8183,N_8760);
and U9673 (N_9673,N_8594,N_8097);
nor U9674 (N_9674,N_8945,N_8002);
nor U9675 (N_9675,N_8285,N_8314);
nor U9676 (N_9676,N_8298,N_8082);
nand U9677 (N_9677,N_8523,N_8562);
or U9678 (N_9678,N_8944,N_8648);
and U9679 (N_9679,N_8933,N_8960);
or U9680 (N_9680,N_8504,N_8677);
and U9681 (N_9681,N_8259,N_8664);
nand U9682 (N_9682,N_8510,N_8609);
and U9683 (N_9683,N_8072,N_8310);
xor U9684 (N_9684,N_8317,N_8786);
and U9685 (N_9685,N_8067,N_8941);
nor U9686 (N_9686,N_8662,N_8256);
nor U9687 (N_9687,N_8617,N_8051);
nor U9688 (N_9688,N_8489,N_8331);
nand U9689 (N_9689,N_8665,N_8835);
nand U9690 (N_9690,N_8923,N_8385);
nor U9691 (N_9691,N_8413,N_8016);
nor U9692 (N_9692,N_8619,N_8532);
nor U9693 (N_9693,N_8671,N_8519);
or U9694 (N_9694,N_8931,N_8464);
or U9695 (N_9695,N_8020,N_8959);
or U9696 (N_9696,N_8305,N_8554);
and U9697 (N_9697,N_8691,N_8990);
nand U9698 (N_9698,N_8153,N_8716);
or U9699 (N_9699,N_8969,N_8252);
and U9700 (N_9700,N_8932,N_8184);
nand U9701 (N_9701,N_8427,N_8132);
or U9702 (N_9702,N_8813,N_8633);
xnor U9703 (N_9703,N_8985,N_8660);
nand U9704 (N_9704,N_8714,N_8877);
and U9705 (N_9705,N_8050,N_8284);
xor U9706 (N_9706,N_8065,N_8511);
or U9707 (N_9707,N_8122,N_8383);
or U9708 (N_9708,N_8820,N_8316);
and U9709 (N_9709,N_8412,N_8732);
nand U9710 (N_9710,N_8686,N_8653);
nor U9711 (N_9711,N_8810,N_8009);
and U9712 (N_9712,N_8040,N_8304);
or U9713 (N_9713,N_8220,N_8425);
and U9714 (N_9714,N_8492,N_8615);
nand U9715 (N_9715,N_8245,N_8885);
xnor U9716 (N_9716,N_8530,N_8021);
or U9717 (N_9717,N_8625,N_8003);
nor U9718 (N_9718,N_8286,N_8707);
or U9719 (N_9719,N_8205,N_8946);
or U9720 (N_9720,N_8650,N_8173);
or U9721 (N_9721,N_8870,N_8425);
nor U9722 (N_9722,N_8267,N_8426);
and U9723 (N_9723,N_8328,N_8476);
nor U9724 (N_9724,N_8190,N_8922);
nor U9725 (N_9725,N_8822,N_8887);
nor U9726 (N_9726,N_8542,N_8957);
and U9727 (N_9727,N_8267,N_8255);
nand U9728 (N_9728,N_8055,N_8437);
nor U9729 (N_9729,N_8227,N_8616);
or U9730 (N_9730,N_8200,N_8784);
and U9731 (N_9731,N_8422,N_8686);
and U9732 (N_9732,N_8475,N_8534);
and U9733 (N_9733,N_8601,N_8847);
nand U9734 (N_9734,N_8920,N_8857);
nand U9735 (N_9735,N_8626,N_8188);
and U9736 (N_9736,N_8510,N_8664);
and U9737 (N_9737,N_8716,N_8868);
nor U9738 (N_9738,N_8373,N_8298);
or U9739 (N_9739,N_8542,N_8827);
or U9740 (N_9740,N_8365,N_8504);
nand U9741 (N_9741,N_8307,N_8009);
or U9742 (N_9742,N_8878,N_8165);
nor U9743 (N_9743,N_8087,N_8186);
and U9744 (N_9744,N_8485,N_8962);
nand U9745 (N_9745,N_8758,N_8806);
nand U9746 (N_9746,N_8385,N_8168);
nand U9747 (N_9747,N_8417,N_8597);
xnor U9748 (N_9748,N_8254,N_8156);
nand U9749 (N_9749,N_8245,N_8898);
and U9750 (N_9750,N_8085,N_8887);
xnor U9751 (N_9751,N_8485,N_8619);
nand U9752 (N_9752,N_8350,N_8175);
nor U9753 (N_9753,N_8529,N_8776);
or U9754 (N_9754,N_8047,N_8887);
and U9755 (N_9755,N_8993,N_8898);
or U9756 (N_9756,N_8386,N_8541);
nor U9757 (N_9757,N_8467,N_8271);
nor U9758 (N_9758,N_8134,N_8426);
or U9759 (N_9759,N_8888,N_8972);
nand U9760 (N_9760,N_8593,N_8469);
or U9761 (N_9761,N_8563,N_8822);
nand U9762 (N_9762,N_8649,N_8082);
xor U9763 (N_9763,N_8462,N_8487);
nand U9764 (N_9764,N_8359,N_8507);
and U9765 (N_9765,N_8857,N_8144);
or U9766 (N_9766,N_8355,N_8463);
nor U9767 (N_9767,N_8679,N_8778);
nor U9768 (N_9768,N_8600,N_8444);
or U9769 (N_9769,N_8813,N_8949);
and U9770 (N_9770,N_8790,N_8864);
nand U9771 (N_9771,N_8739,N_8072);
and U9772 (N_9772,N_8938,N_8143);
and U9773 (N_9773,N_8740,N_8878);
nand U9774 (N_9774,N_8443,N_8253);
or U9775 (N_9775,N_8635,N_8729);
nand U9776 (N_9776,N_8053,N_8983);
or U9777 (N_9777,N_8432,N_8574);
and U9778 (N_9778,N_8158,N_8073);
xnor U9779 (N_9779,N_8459,N_8681);
or U9780 (N_9780,N_8085,N_8693);
nand U9781 (N_9781,N_8659,N_8254);
xor U9782 (N_9782,N_8134,N_8421);
or U9783 (N_9783,N_8610,N_8544);
nor U9784 (N_9784,N_8347,N_8606);
nand U9785 (N_9785,N_8302,N_8009);
xor U9786 (N_9786,N_8994,N_8508);
or U9787 (N_9787,N_8915,N_8191);
and U9788 (N_9788,N_8788,N_8420);
or U9789 (N_9789,N_8957,N_8033);
nor U9790 (N_9790,N_8121,N_8800);
nor U9791 (N_9791,N_8864,N_8974);
nand U9792 (N_9792,N_8964,N_8333);
nor U9793 (N_9793,N_8156,N_8792);
and U9794 (N_9794,N_8309,N_8454);
or U9795 (N_9795,N_8219,N_8593);
nor U9796 (N_9796,N_8676,N_8987);
xor U9797 (N_9797,N_8538,N_8938);
xnor U9798 (N_9798,N_8912,N_8031);
or U9799 (N_9799,N_8899,N_8104);
or U9800 (N_9800,N_8148,N_8323);
and U9801 (N_9801,N_8542,N_8679);
and U9802 (N_9802,N_8526,N_8769);
or U9803 (N_9803,N_8732,N_8016);
nand U9804 (N_9804,N_8928,N_8620);
and U9805 (N_9805,N_8998,N_8915);
nand U9806 (N_9806,N_8207,N_8052);
nor U9807 (N_9807,N_8766,N_8073);
or U9808 (N_9808,N_8884,N_8989);
nand U9809 (N_9809,N_8303,N_8520);
nor U9810 (N_9810,N_8886,N_8594);
nor U9811 (N_9811,N_8421,N_8259);
nand U9812 (N_9812,N_8925,N_8569);
nand U9813 (N_9813,N_8862,N_8710);
and U9814 (N_9814,N_8789,N_8262);
and U9815 (N_9815,N_8790,N_8341);
nand U9816 (N_9816,N_8200,N_8155);
nor U9817 (N_9817,N_8454,N_8853);
nand U9818 (N_9818,N_8167,N_8230);
nor U9819 (N_9819,N_8278,N_8758);
nor U9820 (N_9820,N_8736,N_8423);
nor U9821 (N_9821,N_8066,N_8232);
or U9822 (N_9822,N_8258,N_8406);
nand U9823 (N_9823,N_8572,N_8822);
nor U9824 (N_9824,N_8479,N_8500);
nor U9825 (N_9825,N_8666,N_8957);
nor U9826 (N_9826,N_8538,N_8555);
nand U9827 (N_9827,N_8258,N_8670);
nand U9828 (N_9828,N_8500,N_8496);
and U9829 (N_9829,N_8245,N_8051);
xor U9830 (N_9830,N_8245,N_8279);
or U9831 (N_9831,N_8706,N_8789);
nand U9832 (N_9832,N_8600,N_8802);
nor U9833 (N_9833,N_8497,N_8790);
nand U9834 (N_9834,N_8248,N_8455);
nand U9835 (N_9835,N_8572,N_8203);
or U9836 (N_9836,N_8934,N_8085);
xor U9837 (N_9837,N_8712,N_8600);
xnor U9838 (N_9838,N_8324,N_8474);
or U9839 (N_9839,N_8694,N_8175);
or U9840 (N_9840,N_8721,N_8136);
nor U9841 (N_9841,N_8027,N_8308);
xnor U9842 (N_9842,N_8085,N_8691);
nor U9843 (N_9843,N_8344,N_8899);
nand U9844 (N_9844,N_8357,N_8178);
or U9845 (N_9845,N_8211,N_8744);
and U9846 (N_9846,N_8924,N_8816);
nor U9847 (N_9847,N_8686,N_8590);
nand U9848 (N_9848,N_8917,N_8408);
nand U9849 (N_9849,N_8964,N_8193);
nor U9850 (N_9850,N_8968,N_8808);
nand U9851 (N_9851,N_8422,N_8833);
and U9852 (N_9852,N_8862,N_8324);
and U9853 (N_9853,N_8634,N_8854);
or U9854 (N_9854,N_8466,N_8331);
nor U9855 (N_9855,N_8487,N_8139);
or U9856 (N_9856,N_8227,N_8619);
or U9857 (N_9857,N_8051,N_8995);
nor U9858 (N_9858,N_8621,N_8718);
and U9859 (N_9859,N_8635,N_8186);
nor U9860 (N_9860,N_8044,N_8182);
xor U9861 (N_9861,N_8306,N_8405);
xnor U9862 (N_9862,N_8739,N_8413);
nor U9863 (N_9863,N_8657,N_8908);
and U9864 (N_9864,N_8810,N_8263);
nor U9865 (N_9865,N_8934,N_8235);
nor U9866 (N_9866,N_8821,N_8163);
and U9867 (N_9867,N_8828,N_8234);
and U9868 (N_9868,N_8447,N_8634);
nand U9869 (N_9869,N_8879,N_8454);
xnor U9870 (N_9870,N_8861,N_8116);
and U9871 (N_9871,N_8767,N_8341);
nand U9872 (N_9872,N_8991,N_8821);
and U9873 (N_9873,N_8950,N_8545);
or U9874 (N_9874,N_8477,N_8880);
and U9875 (N_9875,N_8272,N_8242);
nor U9876 (N_9876,N_8539,N_8754);
xnor U9877 (N_9877,N_8845,N_8818);
nand U9878 (N_9878,N_8006,N_8662);
nand U9879 (N_9879,N_8938,N_8185);
and U9880 (N_9880,N_8295,N_8266);
and U9881 (N_9881,N_8500,N_8466);
nand U9882 (N_9882,N_8489,N_8842);
nor U9883 (N_9883,N_8865,N_8743);
nand U9884 (N_9884,N_8110,N_8178);
nor U9885 (N_9885,N_8343,N_8958);
and U9886 (N_9886,N_8932,N_8923);
nand U9887 (N_9887,N_8908,N_8038);
nand U9888 (N_9888,N_8385,N_8498);
or U9889 (N_9889,N_8457,N_8672);
nand U9890 (N_9890,N_8600,N_8271);
and U9891 (N_9891,N_8443,N_8563);
and U9892 (N_9892,N_8791,N_8579);
nand U9893 (N_9893,N_8325,N_8951);
nor U9894 (N_9894,N_8797,N_8047);
and U9895 (N_9895,N_8602,N_8983);
xnor U9896 (N_9896,N_8171,N_8221);
nor U9897 (N_9897,N_8997,N_8746);
xor U9898 (N_9898,N_8872,N_8212);
and U9899 (N_9899,N_8602,N_8863);
xnor U9900 (N_9900,N_8950,N_8461);
or U9901 (N_9901,N_8465,N_8243);
nor U9902 (N_9902,N_8288,N_8243);
nor U9903 (N_9903,N_8635,N_8806);
or U9904 (N_9904,N_8155,N_8685);
nor U9905 (N_9905,N_8341,N_8126);
and U9906 (N_9906,N_8297,N_8851);
nor U9907 (N_9907,N_8420,N_8720);
and U9908 (N_9908,N_8565,N_8015);
or U9909 (N_9909,N_8654,N_8350);
and U9910 (N_9910,N_8013,N_8394);
nand U9911 (N_9911,N_8472,N_8389);
nand U9912 (N_9912,N_8605,N_8974);
and U9913 (N_9913,N_8998,N_8184);
and U9914 (N_9914,N_8804,N_8606);
nand U9915 (N_9915,N_8926,N_8483);
nor U9916 (N_9916,N_8854,N_8425);
xnor U9917 (N_9917,N_8805,N_8630);
nand U9918 (N_9918,N_8683,N_8433);
or U9919 (N_9919,N_8341,N_8082);
or U9920 (N_9920,N_8020,N_8483);
nor U9921 (N_9921,N_8298,N_8771);
and U9922 (N_9922,N_8936,N_8811);
xor U9923 (N_9923,N_8255,N_8678);
xor U9924 (N_9924,N_8991,N_8421);
nor U9925 (N_9925,N_8078,N_8559);
xor U9926 (N_9926,N_8272,N_8724);
or U9927 (N_9927,N_8267,N_8167);
and U9928 (N_9928,N_8276,N_8334);
nor U9929 (N_9929,N_8192,N_8133);
nor U9930 (N_9930,N_8379,N_8961);
nand U9931 (N_9931,N_8505,N_8579);
nor U9932 (N_9932,N_8072,N_8295);
nor U9933 (N_9933,N_8144,N_8980);
and U9934 (N_9934,N_8740,N_8083);
and U9935 (N_9935,N_8560,N_8104);
and U9936 (N_9936,N_8254,N_8035);
nand U9937 (N_9937,N_8936,N_8248);
nand U9938 (N_9938,N_8932,N_8381);
nor U9939 (N_9939,N_8996,N_8451);
xor U9940 (N_9940,N_8969,N_8687);
nor U9941 (N_9941,N_8527,N_8483);
or U9942 (N_9942,N_8641,N_8594);
or U9943 (N_9943,N_8899,N_8931);
or U9944 (N_9944,N_8557,N_8796);
or U9945 (N_9945,N_8124,N_8820);
or U9946 (N_9946,N_8763,N_8725);
or U9947 (N_9947,N_8412,N_8278);
nand U9948 (N_9948,N_8115,N_8263);
and U9949 (N_9949,N_8411,N_8296);
nor U9950 (N_9950,N_8884,N_8038);
and U9951 (N_9951,N_8480,N_8627);
or U9952 (N_9952,N_8005,N_8551);
nand U9953 (N_9953,N_8340,N_8309);
nor U9954 (N_9954,N_8147,N_8951);
or U9955 (N_9955,N_8061,N_8012);
or U9956 (N_9956,N_8347,N_8894);
and U9957 (N_9957,N_8305,N_8511);
nor U9958 (N_9958,N_8685,N_8858);
or U9959 (N_9959,N_8238,N_8086);
nor U9960 (N_9960,N_8441,N_8332);
and U9961 (N_9961,N_8159,N_8624);
or U9962 (N_9962,N_8207,N_8854);
nor U9963 (N_9963,N_8255,N_8704);
or U9964 (N_9964,N_8919,N_8058);
or U9965 (N_9965,N_8309,N_8271);
nand U9966 (N_9966,N_8787,N_8978);
nor U9967 (N_9967,N_8550,N_8974);
or U9968 (N_9968,N_8555,N_8261);
or U9969 (N_9969,N_8956,N_8210);
and U9970 (N_9970,N_8301,N_8194);
and U9971 (N_9971,N_8767,N_8112);
or U9972 (N_9972,N_8507,N_8488);
or U9973 (N_9973,N_8522,N_8035);
and U9974 (N_9974,N_8469,N_8026);
or U9975 (N_9975,N_8978,N_8795);
and U9976 (N_9976,N_8271,N_8540);
or U9977 (N_9977,N_8701,N_8259);
or U9978 (N_9978,N_8925,N_8626);
nor U9979 (N_9979,N_8188,N_8962);
nor U9980 (N_9980,N_8744,N_8392);
nor U9981 (N_9981,N_8452,N_8164);
nor U9982 (N_9982,N_8081,N_8041);
nand U9983 (N_9983,N_8274,N_8365);
xnor U9984 (N_9984,N_8162,N_8418);
or U9985 (N_9985,N_8257,N_8253);
nand U9986 (N_9986,N_8418,N_8597);
and U9987 (N_9987,N_8206,N_8051);
nand U9988 (N_9988,N_8684,N_8185);
xnor U9989 (N_9989,N_8303,N_8110);
and U9990 (N_9990,N_8987,N_8164);
nand U9991 (N_9991,N_8749,N_8716);
nor U9992 (N_9992,N_8304,N_8349);
and U9993 (N_9993,N_8979,N_8555);
nor U9994 (N_9994,N_8483,N_8899);
or U9995 (N_9995,N_8291,N_8235);
nor U9996 (N_9996,N_8752,N_8045);
nor U9997 (N_9997,N_8460,N_8414);
and U9998 (N_9998,N_8642,N_8623);
or U9999 (N_9999,N_8234,N_8442);
nand UO_0 (O_0,N_9956,N_9471);
nor UO_1 (O_1,N_9394,N_9981);
and UO_2 (O_2,N_9553,N_9266);
xor UO_3 (O_3,N_9004,N_9835);
and UO_4 (O_4,N_9057,N_9098);
xor UO_5 (O_5,N_9872,N_9606);
and UO_6 (O_6,N_9194,N_9491);
nand UO_7 (O_7,N_9311,N_9242);
nand UO_8 (O_8,N_9556,N_9416);
xnor UO_9 (O_9,N_9882,N_9966);
or UO_10 (O_10,N_9274,N_9030);
or UO_11 (O_11,N_9457,N_9347);
and UO_12 (O_12,N_9975,N_9176);
and UO_13 (O_13,N_9875,N_9074);
and UO_14 (O_14,N_9636,N_9614);
nand UO_15 (O_15,N_9657,N_9760);
nor UO_16 (O_16,N_9679,N_9929);
or UO_17 (O_17,N_9714,N_9314);
and UO_18 (O_18,N_9191,N_9379);
and UO_19 (O_19,N_9385,N_9174);
nor UO_20 (O_20,N_9041,N_9490);
or UO_21 (O_21,N_9122,N_9091);
nor UO_22 (O_22,N_9983,N_9251);
or UO_23 (O_23,N_9617,N_9392);
and UO_24 (O_24,N_9009,N_9878);
nor UO_25 (O_25,N_9737,N_9149);
nor UO_26 (O_26,N_9367,N_9836);
and UO_27 (O_27,N_9500,N_9934);
or UO_28 (O_28,N_9376,N_9622);
or UO_29 (O_29,N_9293,N_9791);
and UO_30 (O_30,N_9087,N_9248);
and UO_31 (O_31,N_9106,N_9017);
nor UO_32 (O_32,N_9543,N_9620);
nand UO_33 (O_33,N_9339,N_9300);
xor UO_34 (O_34,N_9955,N_9774);
or UO_35 (O_35,N_9072,N_9838);
nor UO_36 (O_36,N_9233,N_9272);
xor UO_37 (O_37,N_9834,N_9375);
or UO_38 (O_38,N_9532,N_9582);
xnor UO_39 (O_39,N_9720,N_9800);
nor UO_40 (O_40,N_9255,N_9103);
or UO_41 (O_41,N_9434,N_9411);
and UO_42 (O_42,N_9298,N_9031);
xnor UO_43 (O_43,N_9913,N_9662);
and UO_44 (O_44,N_9018,N_9277);
nand UO_45 (O_45,N_9598,N_9978);
and UO_46 (O_46,N_9717,N_9597);
or UO_47 (O_47,N_9499,N_9778);
nor UO_48 (O_48,N_9509,N_9159);
nor UO_49 (O_49,N_9039,N_9084);
nor UO_50 (O_50,N_9750,N_9768);
and UO_51 (O_51,N_9855,N_9535);
nor UO_52 (O_52,N_9050,N_9328);
and UO_53 (O_53,N_9080,N_9549);
nand UO_54 (O_54,N_9708,N_9295);
or UO_55 (O_55,N_9204,N_9974);
and UO_56 (O_56,N_9970,N_9584);
or UO_57 (O_57,N_9056,N_9216);
nand UO_58 (O_58,N_9296,N_9938);
nor UO_59 (O_59,N_9349,N_9062);
and UO_60 (O_60,N_9630,N_9104);
and UO_61 (O_61,N_9828,N_9188);
nor UO_62 (O_62,N_9023,N_9670);
or UO_63 (O_63,N_9944,N_9270);
or UO_64 (O_64,N_9051,N_9797);
nor UO_65 (O_65,N_9503,N_9766);
and UO_66 (O_66,N_9664,N_9195);
nor UO_67 (O_67,N_9355,N_9868);
and UO_68 (O_68,N_9169,N_9583);
and UO_69 (O_69,N_9267,N_9345);
nor UO_70 (O_70,N_9782,N_9640);
and UO_71 (O_71,N_9603,N_9982);
or UO_72 (O_72,N_9458,N_9015);
nand UO_73 (O_73,N_9097,N_9819);
nor UO_74 (O_74,N_9923,N_9413);
or UO_75 (O_75,N_9523,N_9891);
or UO_76 (O_76,N_9324,N_9439);
and UO_77 (O_77,N_9874,N_9867);
and UO_78 (O_78,N_9447,N_9014);
nor UO_79 (O_79,N_9764,N_9109);
or UO_80 (O_80,N_9455,N_9035);
nand UO_81 (O_81,N_9526,N_9680);
nand UO_82 (O_82,N_9564,N_9541);
and UO_83 (O_83,N_9420,N_9772);
nand UO_84 (O_84,N_9817,N_9605);
or UO_85 (O_85,N_9646,N_9137);
xnor UO_86 (O_86,N_9613,N_9007);
or UO_87 (O_87,N_9907,N_9390);
and UO_88 (O_88,N_9610,N_9108);
and UO_89 (O_89,N_9842,N_9733);
nor UO_90 (O_90,N_9847,N_9093);
nand UO_91 (O_91,N_9673,N_9016);
nand UO_92 (O_92,N_9719,N_9412);
nand UO_93 (O_93,N_9914,N_9644);
xnor UO_94 (O_94,N_9684,N_9825);
or UO_95 (O_95,N_9323,N_9130);
or UO_96 (O_96,N_9936,N_9950);
or UO_97 (O_97,N_9542,N_9378);
nor UO_98 (O_98,N_9048,N_9538);
nand UO_99 (O_99,N_9182,N_9550);
nor UO_100 (O_100,N_9384,N_9453);
and UO_101 (O_101,N_9609,N_9281);
nor UO_102 (O_102,N_9568,N_9168);
and UO_103 (O_103,N_9735,N_9705);
nand UO_104 (O_104,N_9128,N_9706);
or UO_105 (O_105,N_9659,N_9818);
and UO_106 (O_106,N_9200,N_9724);
nor UO_107 (O_107,N_9107,N_9886);
nand UO_108 (O_108,N_9520,N_9813);
xor UO_109 (O_109,N_9952,N_9132);
xnor UO_110 (O_110,N_9902,N_9309);
or UO_111 (O_111,N_9743,N_9124);
nor UO_112 (O_112,N_9740,N_9739);
nand UO_113 (O_113,N_9313,N_9892);
or UO_114 (O_114,N_9231,N_9859);
and UO_115 (O_115,N_9076,N_9029);
nor UO_116 (O_116,N_9082,N_9258);
or UO_117 (O_117,N_9885,N_9780);
nand UO_118 (O_118,N_9770,N_9444);
and UO_119 (O_119,N_9883,N_9346);
nor UO_120 (O_120,N_9158,N_9424);
xnor UO_121 (O_121,N_9754,N_9781);
nand UO_122 (O_122,N_9320,N_9228);
or UO_123 (O_123,N_9700,N_9359);
or UO_124 (O_124,N_9213,N_9683);
nand UO_125 (O_125,N_9887,N_9333);
or UO_126 (O_126,N_9515,N_9466);
nand UO_127 (O_127,N_9984,N_9371);
nand UO_128 (O_128,N_9064,N_9665);
or UO_129 (O_129,N_9473,N_9111);
nor UO_130 (O_130,N_9101,N_9634);
nor UO_131 (O_131,N_9330,N_9381);
and UO_132 (O_132,N_9910,N_9729);
xor UO_133 (O_133,N_9462,N_9113);
nand UO_134 (O_134,N_9297,N_9736);
or UO_135 (O_135,N_9331,N_9723);
and UO_136 (O_136,N_9954,N_9011);
and UO_137 (O_137,N_9933,N_9927);
nand UO_138 (O_138,N_9506,N_9884);
or UO_139 (O_139,N_9587,N_9998);
nor UO_140 (O_140,N_9329,N_9181);
and UO_141 (O_141,N_9960,N_9157);
or UO_142 (O_142,N_9555,N_9962);
nor UO_143 (O_143,N_9534,N_9469);
nor UO_144 (O_144,N_9880,N_9881);
nor UO_145 (O_145,N_9059,N_9682);
or UO_146 (O_146,N_9055,N_9493);
nor UO_147 (O_147,N_9687,N_9257);
or UO_148 (O_148,N_9627,N_9635);
and UO_149 (O_149,N_9177,N_9341);
nor UO_150 (O_150,N_9900,N_9336);
or UO_151 (O_151,N_9917,N_9437);
or UO_152 (O_152,N_9649,N_9979);
or UO_153 (O_153,N_9372,N_9840);
and UO_154 (O_154,N_9839,N_9226);
or UO_155 (O_155,N_9273,N_9013);
nor UO_156 (O_156,N_9429,N_9691);
or UO_157 (O_157,N_9285,N_9941);
nand UO_158 (O_158,N_9809,N_9485);
or UO_159 (O_159,N_9096,N_9256);
and UO_160 (O_160,N_9987,N_9578);
and UO_161 (O_161,N_9557,N_9012);
nor UO_162 (O_162,N_9033,N_9655);
and UO_163 (O_163,N_9088,N_9170);
nor UO_164 (O_164,N_9856,N_9230);
xor UO_165 (O_165,N_9316,N_9484);
nand UO_166 (O_166,N_9653,N_9734);
and UO_167 (O_167,N_9721,N_9036);
nor UO_168 (O_168,N_9574,N_9260);
and UO_169 (O_169,N_9674,N_9593);
nor UO_170 (O_170,N_9661,N_9548);
nand UO_171 (O_171,N_9250,N_9776);
or UO_172 (O_172,N_9395,N_9504);
or UO_173 (O_173,N_9896,N_9607);
nor UO_174 (O_174,N_9862,N_9284);
and UO_175 (O_175,N_9689,N_9214);
and UO_176 (O_176,N_9786,N_9784);
nand UO_177 (O_177,N_9652,N_9792);
and UO_178 (O_178,N_9483,N_9702);
nand UO_179 (O_179,N_9287,N_9428);
and UO_180 (O_180,N_9816,N_9077);
nor UO_181 (O_181,N_9079,N_9432);
xor UO_182 (O_182,N_9890,N_9858);
xor UO_183 (O_183,N_9445,N_9299);
and UO_184 (O_184,N_9322,N_9259);
or UO_185 (O_185,N_9581,N_9380);
and UO_186 (O_186,N_9579,N_9854);
or UO_187 (O_187,N_9748,N_9730);
xor UO_188 (O_188,N_9366,N_9871);
or UO_189 (O_189,N_9183,N_9551);
nand UO_190 (O_190,N_9105,N_9671);
xnor UO_191 (O_191,N_9946,N_9305);
nand UO_192 (O_192,N_9086,N_9419);
xor UO_193 (O_193,N_9830,N_9407);
nand UO_194 (O_194,N_9722,N_9775);
nand UO_195 (O_195,N_9901,N_9222);
nor UO_196 (O_196,N_9224,N_9431);
nor UO_197 (O_197,N_9192,N_9758);
or UO_198 (O_198,N_9089,N_9461);
and UO_199 (O_199,N_9522,N_9771);
or UO_200 (O_200,N_9712,N_9544);
nor UO_201 (O_201,N_9387,N_9127);
nor UO_202 (O_202,N_9291,N_9211);
nand UO_203 (O_203,N_9247,N_9894);
nor UO_204 (O_204,N_9262,N_9190);
or UO_205 (O_205,N_9136,N_9761);
xnor UO_206 (O_206,N_9377,N_9915);
and UO_207 (O_207,N_9241,N_9547);
nor UO_208 (O_208,N_9102,N_9586);
and UO_209 (O_209,N_9186,N_9650);
and UO_210 (O_210,N_9278,N_9117);
nand UO_211 (O_211,N_9645,N_9417);
nor UO_212 (O_212,N_9678,N_9232);
nor UO_213 (O_213,N_9773,N_9427);
and UO_214 (O_214,N_9423,N_9566);
and UO_215 (O_215,N_9326,N_9308);
nand UO_216 (O_216,N_9713,N_9477);
nor UO_217 (O_217,N_9386,N_9133);
or UO_218 (O_218,N_9873,N_9121);
nor UO_219 (O_219,N_9225,N_9140);
nand UO_220 (O_220,N_9363,N_9595);
xor UO_221 (O_221,N_9741,N_9876);
nand UO_222 (O_222,N_9561,N_9513);
xor UO_223 (O_223,N_9686,N_9451);
or UO_224 (O_224,N_9340,N_9234);
nand UO_225 (O_225,N_9788,N_9067);
or UO_226 (O_226,N_9560,N_9221);
nand UO_227 (O_227,N_9253,N_9034);
nand UO_228 (O_228,N_9647,N_9348);
nor UO_229 (O_229,N_9604,N_9038);
or UO_230 (O_230,N_9977,N_9053);
xnor UO_231 (O_231,N_9958,N_9027);
nand UO_232 (O_232,N_9718,N_9154);
or UO_233 (O_233,N_9342,N_9530);
nand UO_234 (O_234,N_9318,N_9135);
xnor UO_235 (O_235,N_9672,N_9658);
nor UO_236 (O_236,N_9220,N_9252);
nand UO_237 (O_237,N_9510,N_9205);
or UO_238 (O_238,N_9354,N_9060);
nand UO_239 (O_239,N_9529,N_9010);
xnor UO_240 (O_240,N_9276,N_9812);
or UO_241 (O_241,N_9238,N_9539);
and UO_242 (O_242,N_9288,N_9237);
or UO_243 (O_243,N_9498,N_9994);
or UO_244 (O_244,N_9254,N_9826);
and UO_245 (O_245,N_9454,N_9594);
xnor UO_246 (O_246,N_9943,N_9240);
nor UO_247 (O_247,N_9474,N_9843);
nand UO_248 (O_248,N_9338,N_9271);
nand UO_249 (O_249,N_9217,N_9352);
nor UO_250 (O_250,N_9728,N_9081);
and UO_251 (O_251,N_9279,N_9175);
nor UO_252 (O_252,N_9755,N_9196);
nor UO_253 (O_253,N_9621,N_9959);
nand UO_254 (O_254,N_9212,N_9094);
and UO_255 (O_255,N_9688,N_9747);
or UO_256 (O_256,N_9099,N_9292);
or UO_257 (O_257,N_9919,N_9951);
and UO_258 (O_258,N_9567,N_9866);
or UO_259 (O_259,N_9798,N_9861);
or UO_260 (O_260,N_9832,N_9391);
nor UO_261 (O_261,N_9058,N_9964);
nand UO_262 (O_262,N_9920,N_9388);
and UO_263 (O_263,N_9619,N_9853);
and UO_264 (O_264,N_9189,N_9845);
and UO_265 (O_265,N_9403,N_9463);
nor UO_266 (O_266,N_9236,N_9945);
nor UO_267 (O_267,N_9280,N_9289);
nand UO_268 (O_268,N_9996,N_9042);
nand UO_269 (O_269,N_9024,N_9531);
or UO_270 (O_270,N_9801,N_9441);
or UO_271 (O_271,N_9559,N_9043);
nand UO_272 (O_272,N_9249,N_9973);
nor UO_273 (O_273,N_9732,N_9536);
and UO_274 (O_274,N_9187,N_9160);
or UO_275 (O_275,N_9501,N_9435);
nand UO_276 (O_276,N_9208,N_9779);
xor UO_277 (O_277,N_9667,N_9669);
and UO_278 (O_278,N_9494,N_9351);
and UO_279 (O_279,N_9756,N_9590);
nor UO_280 (O_280,N_9065,N_9406);
or UO_281 (O_281,N_9690,N_9898);
nor UO_282 (O_282,N_9472,N_9668);
and UO_283 (O_283,N_9931,N_9997);
nand UO_284 (O_284,N_9525,N_9275);
and UO_285 (O_285,N_9162,N_9628);
nor UO_286 (O_286,N_9841,N_9511);
or UO_287 (O_287,N_9942,N_9283);
nand UO_288 (O_288,N_9641,N_9215);
nor UO_289 (O_289,N_9971,N_9731);
and UO_290 (O_290,N_9408,N_9460);
nor UO_291 (O_291,N_9602,N_9999);
and UO_292 (O_292,N_9167,N_9393);
nand UO_293 (O_293,N_9165,N_9244);
xnor UO_294 (O_294,N_9134,N_9580);
nand UO_295 (O_295,N_9025,N_9206);
or UO_296 (O_296,N_9002,N_9294);
and UO_297 (O_297,N_9040,N_9235);
and UO_298 (O_298,N_9245,N_9546);
nand UO_299 (O_299,N_9161,N_9193);
and UO_300 (O_300,N_9178,N_9207);
and UO_301 (O_301,N_9304,N_9047);
or UO_302 (O_302,N_9637,N_9571);
or UO_303 (O_303,N_9343,N_9846);
or UO_304 (O_304,N_9396,N_9696);
or UO_305 (O_305,N_9803,N_9143);
and UO_306 (O_306,N_9948,N_9849);
nand UO_307 (O_307,N_9957,N_9239);
nor UO_308 (O_308,N_9261,N_9425);
or UO_309 (O_309,N_9001,N_9918);
nor UO_310 (O_310,N_9608,N_9155);
xnor UO_311 (O_311,N_9577,N_9402);
or UO_312 (O_312,N_9935,N_9654);
or UO_313 (O_313,N_9022,N_9726);
or UO_314 (O_314,N_9600,N_9796);
xor UO_315 (O_315,N_9020,N_9071);
or UO_316 (O_316,N_9335,N_9704);
or UO_317 (O_317,N_9418,N_9307);
and UO_318 (O_318,N_9599,N_9401);
and UO_319 (O_319,N_9448,N_9626);
nand UO_320 (O_320,N_9479,N_9616);
and UO_321 (O_321,N_9759,N_9456);
and UO_322 (O_322,N_9459,N_9404);
and UO_323 (O_323,N_9497,N_9889);
xor UO_324 (O_324,N_9110,N_9694);
nor UO_325 (O_325,N_9464,N_9037);
nand UO_326 (O_326,N_9449,N_9837);
and UO_327 (O_327,N_9831,N_9061);
or UO_328 (O_328,N_9166,N_9519);
and UO_329 (O_329,N_9752,N_9442);
nor UO_330 (O_330,N_9633,N_9601);
or UO_331 (O_331,N_9656,N_9681);
or UO_332 (O_332,N_9319,N_9487);
or UO_333 (O_333,N_9807,N_9793);
nand UO_334 (O_334,N_9045,N_9073);
and UO_335 (O_335,N_9138,N_9725);
and UO_336 (O_336,N_9869,N_9742);
and UO_337 (O_337,N_9209,N_9976);
and UO_338 (O_338,N_9783,N_9325);
or UO_339 (O_339,N_9930,N_9492);
nor UO_340 (O_340,N_9481,N_9199);
nor UO_341 (O_341,N_9480,N_9524);
nand UO_342 (O_342,N_9624,N_9749);
or UO_343 (O_343,N_9436,N_9374);
nand UO_344 (O_344,N_9360,N_9625);
or UO_345 (O_345,N_9185,N_9877);
nand UO_346 (O_346,N_9075,N_9623);
nor UO_347 (O_347,N_9769,N_9400);
nor UO_348 (O_348,N_9450,N_9833);
xnor UO_349 (O_349,N_9937,N_9692);
and UO_350 (O_350,N_9083,N_9710);
nor UO_351 (O_351,N_9715,N_9264);
nand UO_352 (O_352,N_9171,N_9677);
nand UO_353 (O_353,N_9787,N_9963);
and UO_354 (O_354,N_9006,N_9701);
nand UO_355 (O_355,N_9821,N_9814);
and UO_356 (O_356,N_9201,N_9358);
nor UO_357 (O_357,N_9008,N_9932);
and UO_358 (O_358,N_9939,N_9049);
xnor UO_359 (O_359,N_9990,N_9585);
xnor UO_360 (O_360,N_9085,N_9306);
or UO_361 (O_361,N_9021,N_9589);
nand UO_362 (O_362,N_9414,N_9409);
nor UO_363 (O_363,N_9844,N_9507);
or UO_364 (O_364,N_9227,N_9762);
and UO_365 (O_365,N_9899,N_9139);
and UO_366 (O_366,N_9823,N_9642);
or UO_367 (O_367,N_9468,N_9790);
and UO_368 (O_368,N_9829,N_9476);
nor UO_369 (O_369,N_9146,N_9246);
or UO_370 (O_370,N_9452,N_9757);
and UO_371 (O_371,N_9369,N_9398);
xor UO_372 (O_372,N_9815,N_9632);
or UO_373 (O_373,N_9986,N_9703);
nor UO_374 (O_374,N_9985,N_9044);
nor UO_375 (O_375,N_9365,N_9916);
or UO_376 (O_376,N_9903,N_9820);
and UO_377 (O_377,N_9765,N_9286);
and UO_378 (O_378,N_9777,N_9897);
xor UO_379 (O_379,N_9851,N_9618);
and UO_380 (O_380,N_9475,N_9651);
and UO_381 (O_381,N_9119,N_9095);
nor UO_382 (O_382,N_9940,N_9070);
xnor UO_383 (O_383,N_9810,N_9905);
and UO_384 (O_384,N_9827,N_9282);
nor UO_385 (O_385,N_9972,N_9421);
or UO_386 (O_386,N_9612,N_9019);
xor UO_387 (O_387,N_9357,N_9993);
and UO_388 (O_388,N_9895,N_9502);
nand UO_389 (O_389,N_9629,N_9745);
nor UO_390 (O_390,N_9980,N_9799);
and UO_391 (O_391,N_9518,N_9115);
nand UO_392 (O_392,N_9806,N_9558);
xnor UO_393 (O_393,N_9334,N_9879);
nand UO_394 (O_394,N_9505,N_9908);
or UO_395 (O_395,N_9751,N_9638);
nand UO_396 (O_396,N_9268,N_9969);
and UO_397 (O_397,N_9909,N_9926);
nand UO_398 (O_398,N_9126,N_9517);
nor UO_399 (O_399,N_9588,N_9203);
and UO_400 (O_400,N_9151,N_9353);
nor UO_401 (O_401,N_9685,N_9516);
or UO_402 (O_402,N_9397,N_9545);
nand UO_403 (O_403,N_9290,N_9310);
nor UO_404 (O_404,N_9148,N_9695);
and UO_405 (O_405,N_9860,N_9848);
nand UO_406 (O_406,N_9364,N_9697);
or UO_407 (O_407,N_9123,N_9991);
xnor UO_408 (O_408,N_9144,N_9968);
or UO_409 (O_409,N_9922,N_9301);
or UO_410 (O_410,N_9120,N_9912);
xor UO_411 (O_411,N_9857,N_9785);
nand UO_412 (O_412,N_9763,N_9949);
nand UO_413 (O_413,N_9573,N_9592);
nand UO_414 (O_414,N_9467,N_9906);
and UO_415 (O_415,N_9727,N_9052);
nor UO_416 (O_416,N_9389,N_9537);
nand UO_417 (O_417,N_9716,N_9631);
nand UO_418 (O_418,N_9361,N_9967);
nor UO_419 (O_419,N_9443,N_9184);
or UO_420 (O_420,N_9422,N_9953);
and UO_421 (O_421,N_9527,N_9565);
or UO_422 (O_422,N_9989,N_9362);
and UO_423 (O_423,N_9643,N_9554);
nand UO_424 (O_424,N_9303,N_9486);
or UO_425 (O_425,N_9805,N_9399);
or UO_426 (O_426,N_9965,N_9410);
nor UO_427 (O_427,N_9069,N_9753);
nand UO_428 (O_428,N_9470,N_9988);
and UO_429 (O_429,N_9430,N_9032);
nand UO_430 (O_430,N_9767,N_9570);
nor UO_431 (O_431,N_9824,N_9489);
and UO_432 (O_432,N_9648,N_9163);
nor UO_433 (O_433,N_9063,N_9663);
or UO_434 (O_434,N_9066,N_9321);
nor UO_435 (O_435,N_9028,N_9210);
or UO_436 (O_436,N_9415,N_9533);
nor UO_437 (O_437,N_9446,N_9512);
nand UO_438 (O_438,N_9738,N_9078);
and UO_439 (O_439,N_9591,N_9693);
nor UO_440 (O_440,N_9003,N_9100);
or UO_441 (O_441,N_9269,N_9344);
and UO_442 (O_442,N_9572,N_9676);
nor UO_443 (O_443,N_9569,N_9433);
nor UO_444 (O_444,N_9698,N_9666);
nor UO_445 (O_445,N_9528,N_9150);
nand UO_446 (O_446,N_9576,N_9928);
nand UO_447 (O_447,N_9197,N_9675);
or UO_448 (O_448,N_9164,N_9145);
nand UO_449 (O_449,N_9005,N_9317);
or UO_450 (O_450,N_9921,N_9804);
or UO_451 (O_451,N_9888,N_9552);
nor UO_452 (O_452,N_9229,N_9370);
nand UO_453 (O_453,N_9495,N_9173);
nand UO_454 (O_454,N_9852,N_9440);
nand UO_455 (O_455,N_9660,N_9611);
nor UO_456 (O_456,N_9961,N_9924);
nand UO_457 (O_457,N_9789,N_9865);
xor UO_458 (O_458,N_9118,N_9046);
nand UO_459 (O_459,N_9356,N_9350);
nor UO_460 (O_460,N_9925,N_9219);
xor UO_461 (O_461,N_9180,N_9090);
and UO_462 (O_462,N_9092,N_9265);
and UO_463 (O_463,N_9327,N_9699);
nand UO_464 (O_464,N_9744,N_9794);
xnor UO_465 (O_465,N_9054,N_9540);
nand UO_466 (O_466,N_9368,N_9026);
or UO_467 (O_467,N_9114,N_9141);
and UO_468 (O_468,N_9373,N_9172);
nor UO_469 (O_469,N_9129,N_9382);
and UO_470 (O_470,N_9563,N_9802);
or UO_471 (O_471,N_9383,N_9000);
nor UO_472 (O_472,N_9863,N_9153);
xor UO_473 (O_473,N_9112,N_9864);
or UO_474 (O_474,N_9131,N_9332);
nor UO_475 (O_475,N_9746,N_9795);
nor UO_476 (O_476,N_9514,N_9575);
and UO_477 (O_477,N_9179,N_9808);
and UO_478 (O_478,N_9156,N_9904);
nand UO_479 (O_479,N_9995,N_9707);
nor UO_480 (O_480,N_9562,N_9615);
xor UO_481 (O_481,N_9521,N_9125);
nor UO_482 (O_482,N_9709,N_9711);
or UO_483 (O_483,N_9508,N_9302);
or UO_484 (O_484,N_9947,N_9152);
and UO_485 (O_485,N_9312,N_9405);
nand UO_486 (O_486,N_9596,N_9992);
and UO_487 (O_487,N_9263,N_9147);
xor UO_488 (O_488,N_9202,N_9911);
and UO_489 (O_489,N_9822,N_9068);
nand UO_490 (O_490,N_9850,N_9893);
xor UO_491 (O_491,N_9478,N_9870);
nor UO_492 (O_492,N_9218,N_9496);
or UO_493 (O_493,N_9142,N_9223);
nand UO_494 (O_494,N_9482,N_9465);
nand UO_495 (O_495,N_9426,N_9315);
nand UO_496 (O_496,N_9488,N_9243);
nor UO_497 (O_497,N_9639,N_9116);
nor UO_498 (O_498,N_9198,N_9811);
or UO_499 (O_499,N_9337,N_9438);
nor UO_500 (O_500,N_9213,N_9697);
or UO_501 (O_501,N_9887,N_9337);
nand UO_502 (O_502,N_9423,N_9281);
or UO_503 (O_503,N_9189,N_9144);
nor UO_504 (O_504,N_9707,N_9229);
xnor UO_505 (O_505,N_9126,N_9712);
or UO_506 (O_506,N_9560,N_9789);
nor UO_507 (O_507,N_9367,N_9393);
or UO_508 (O_508,N_9781,N_9766);
nor UO_509 (O_509,N_9297,N_9695);
nor UO_510 (O_510,N_9374,N_9271);
nand UO_511 (O_511,N_9901,N_9039);
or UO_512 (O_512,N_9137,N_9621);
and UO_513 (O_513,N_9765,N_9736);
and UO_514 (O_514,N_9733,N_9674);
nand UO_515 (O_515,N_9496,N_9368);
or UO_516 (O_516,N_9096,N_9764);
nor UO_517 (O_517,N_9434,N_9449);
nand UO_518 (O_518,N_9726,N_9669);
nor UO_519 (O_519,N_9157,N_9271);
or UO_520 (O_520,N_9644,N_9657);
xnor UO_521 (O_521,N_9981,N_9406);
nand UO_522 (O_522,N_9169,N_9072);
or UO_523 (O_523,N_9198,N_9145);
nor UO_524 (O_524,N_9014,N_9534);
xor UO_525 (O_525,N_9915,N_9494);
xnor UO_526 (O_526,N_9443,N_9404);
nor UO_527 (O_527,N_9039,N_9756);
and UO_528 (O_528,N_9906,N_9815);
or UO_529 (O_529,N_9963,N_9223);
nand UO_530 (O_530,N_9080,N_9222);
and UO_531 (O_531,N_9576,N_9382);
nand UO_532 (O_532,N_9934,N_9631);
or UO_533 (O_533,N_9087,N_9439);
or UO_534 (O_534,N_9700,N_9449);
nand UO_535 (O_535,N_9933,N_9845);
or UO_536 (O_536,N_9302,N_9503);
or UO_537 (O_537,N_9827,N_9566);
nand UO_538 (O_538,N_9827,N_9190);
nand UO_539 (O_539,N_9186,N_9913);
and UO_540 (O_540,N_9638,N_9290);
nand UO_541 (O_541,N_9040,N_9742);
and UO_542 (O_542,N_9459,N_9882);
nand UO_543 (O_543,N_9451,N_9866);
or UO_544 (O_544,N_9401,N_9998);
and UO_545 (O_545,N_9084,N_9058);
nor UO_546 (O_546,N_9342,N_9089);
and UO_547 (O_547,N_9378,N_9795);
nor UO_548 (O_548,N_9889,N_9302);
and UO_549 (O_549,N_9171,N_9013);
nand UO_550 (O_550,N_9541,N_9441);
nand UO_551 (O_551,N_9339,N_9188);
or UO_552 (O_552,N_9952,N_9149);
nand UO_553 (O_553,N_9289,N_9510);
nand UO_554 (O_554,N_9120,N_9717);
or UO_555 (O_555,N_9248,N_9143);
nor UO_556 (O_556,N_9663,N_9139);
nor UO_557 (O_557,N_9348,N_9512);
nand UO_558 (O_558,N_9796,N_9846);
or UO_559 (O_559,N_9891,N_9892);
or UO_560 (O_560,N_9404,N_9723);
and UO_561 (O_561,N_9054,N_9541);
xnor UO_562 (O_562,N_9899,N_9953);
nand UO_563 (O_563,N_9407,N_9372);
nor UO_564 (O_564,N_9518,N_9725);
nand UO_565 (O_565,N_9699,N_9519);
nand UO_566 (O_566,N_9304,N_9061);
or UO_567 (O_567,N_9017,N_9118);
nand UO_568 (O_568,N_9720,N_9077);
nor UO_569 (O_569,N_9347,N_9514);
nor UO_570 (O_570,N_9844,N_9177);
nor UO_571 (O_571,N_9127,N_9561);
nor UO_572 (O_572,N_9238,N_9326);
and UO_573 (O_573,N_9064,N_9800);
or UO_574 (O_574,N_9108,N_9368);
and UO_575 (O_575,N_9984,N_9652);
and UO_576 (O_576,N_9601,N_9117);
or UO_577 (O_577,N_9700,N_9035);
or UO_578 (O_578,N_9949,N_9598);
nor UO_579 (O_579,N_9298,N_9304);
nand UO_580 (O_580,N_9574,N_9586);
or UO_581 (O_581,N_9167,N_9596);
or UO_582 (O_582,N_9454,N_9234);
nor UO_583 (O_583,N_9035,N_9114);
nor UO_584 (O_584,N_9819,N_9969);
nand UO_585 (O_585,N_9240,N_9458);
nor UO_586 (O_586,N_9401,N_9535);
and UO_587 (O_587,N_9514,N_9130);
nand UO_588 (O_588,N_9787,N_9558);
and UO_589 (O_589,N_9378,N_9160);
or UO_590 (O_590,N_9818,N_9552);
and UO_591 (O_591,N_9972,N_9594);
or UO_592 (O_592,N_9254,N_9332);
nand UO_593 (O_593,N_9722,N_9000);
nor UO_594 (O_594,N_9617,N_9088);
and UO_595 (O_595,N_9506,N_9992);
nand UO_596 (O_596,N_9242,N_9504);
nand UO_597 (O_597,N_9880,N_9096);
xor UO_598 (O_598,N_9963,N_9632);
or UO_599 (O_599,N_9274,N_9742);
xnor UO_600 (O_600,N_9595,N_9531);
and UO_601 (O_601,N_9857,N_9698);
nor UO_602 (O_602,N_9955,N_9141);
and UO_603 (O_603,N_9038,N_9772);
nand UO_604 (O_604,N_9161,N_9396);
xnor UO_605 (O_605,N_9833,N_9092);
or UO_606 (O_606,N_9078,N_9562);
nand UO_607 (O_607,N_9124,N_9437);
and UO_608 (O_608,N_9072,N_9155);
and UO_609 (O_609,N_9765,N_9010);
nor UO_610 (O_610,N_9657,N_9021);
and UO_611 (O_611,N_9319,N_9147);
nand UO_612 (O_612,N_9317,N_9368);
nand UO_613 (O_613,N_9837,N_9980);
or UO_614 (O_614,N_9080,N_9174);
and UO_615 (O_615,N_9676,N_9877);
or UO_616 (O_616,N_9865,N_9055);
and UO_617 (O_617,N_9362,N_9972);
or UO_618 (O_618,N_9284,N_9233);
nor UO_619 (O_619,N_9516,N_9404);
nor UO_620 (O_620,N_9891,N_9870);
or UO_621 (O_621,N_9492,N_9246);
and UO_622 (O_622,N_9093,N_9906);
and UO_623 (O_623,N_9651,N_9615);
and UO_624 (O_624,N_9766,N_9916);
xor UO_625 (O_625,N_9030,N_9070);
nand UO_626 (O_626,N_9450,N_9733);
and UO_627 (O_627,N_9362,N_9789);
xor UO_628 (O_628,N_9214,N_9070);
nand UO_629 (O_629,N_9702,N_9783);
or UO_630 (O_630,N_9771,N_9837);
nor UO_631 (O_631,N_9384,N_9250);
xor UO_632 (O_632,N_9631,N_9559);
nor UO_633 (O_633,N_9144,N_9389);
nor UO_634 (O_634,N_9090,N_9751);
or UO_635 (O_635,N_9308,N_9653);
nand UO_636 (O_636,N_9822,N_9898);
or UO_637 (O_637,N_9305,N_9029);
or UO_638 (O_638,N_9033,N_9025);
and UO_639 (O_639,N_9292,N_9984);
nor UO_640 (O_640,N_9354,N_9795);
and UO_641 (O_641,N_9366,N_9462);
nor UO_642 (O_642,N_9075,N_9654);
nand UO_643 (O_643,N_9817,N_9735);
nand UO_644 (O_644,N_9784,N_9026);
nor UO_645 (O_645,N_9992,N_9675);
and UO_646 (O_646,N_9385,N_9795);
nand UO_647 (O_647,N_9395,N_9884);
or UO_648 (O_648,N_9492,N_9793);
nand UO_649 (O_649,N_9550,N_9833);
and UO_650 (O_650,N_9927,N_9059);
nand UO_651 (O_651,N_9470,N_9361);
nand UO_652 (O_652,N_9430,N_9193);
xor UO_653 (O_653,N_9597,N_9482);
or UO_654 (O_654,N_9046,N_9006);
nand UO_655 (O_655,N_9007,N_9715);
and UO_656 (O_656,N_9530,N_9156);
or UO_657 (O_657,N_9761,N_9438);
and UO_658 (O_658,N_9726,N_9970);
nor UO_659 (O_659,N_9287,N_9527);
nand UO_660 (O_660,N_9046,N_9773);
nand UO_661 (O_661,N_9632,N_9004);
or UO_662 (O_662,N_9112,N_9322);
or UO_663 (O_663,N_9068,N_9597);
nand UO_664 (O_664,N_9724,N_9900);
nor UO_665 (O_665,N_9240,N_9223);
nor UO_666 (O_666,N_9655,N_9308);
xor UO_667 (O_667,N_9963,N_9381);
nor UO_668 (O_668,N_9644,N_9819);
nor UO_669 (O_669,N_9292,N_9051);
and UO_670 (O_670,N_9546,N_9174);
or UO_671 (O_671,N_9293,N_9591);
nand UO_672 (O_672,N_9021,N_9212);
nand UO_673 (O_673,N_9330,N_9100);
nor UO_674 (O_674,N_9238,N_9749);
nand UO_675 (O_675,N_9994,N_9618);
xnor UO_676 (O_676,N_9782,N_9994);
nand UO_677 (O_677,N_9505,N_9360);
or UO_678 (O_678,N_9889,N_9615);
and UO_679 (O_679,N_9637,N_9985);
nor UO_680 (O_680,N_9634,N_9994);
or UO_681 (O_681,N_9395,N_9455);
and UO_682 (O_682,N_9581,N_9520);
nor UO_683 (O_683,N_9876,N_9329);
and UO_684 (O_684,N_9378,N_9427);
or UO_685 (O_685,N_9073,N_9822);
and UO_686 (O_686,N_9505,N_9772);
or UO_687 (O_687,N_9748,N_9420);
nor UO_688 (O_688,N_9505,N_9316);
and UO_689 (O_689,N_9483,N_9883);
nand UO_690 (O_690,N_9223,N_9781);
nand UO_691 (O_691,N_9086,N_9942);
nor UO_692 (O_692,N_9826,N_9349);
or UO_693 (O_693,N_9784,N_9898);
or UO_694 (O_694,N_9498,N_9285);
or UO_695 (O_695,N_9022,N_9531);
and UO_696 (O_696,N_9756,N_9506);
and UO_697 (O_697,N_9084,N_9739);
nor UO_698 (O_698,N_9408,N_9422);
xnor UO_699 (O_699,N_9847,N_9078);
or UO_700 (O_700,N_9113,N_9400);
and UO_701 (O_701,N_9633,N_9967);
nor UO_702 (O_702,N_9373,N_9924);
nor UO_703 (O_703,N_9835,N_9526);
or UO_704 (O_704,N_9187,N_9004);
nand UO_705 (O_705,N_9074,N_9436);
nand UO_706 (O_706,N_9389,N_9838);
nand UO_707 (O_707,N_9082,N_9375);
nand UO_708 (O_708,N_9887,N_9661);
and UO_709 (O_709,N_9821,N_9311);
nor UO_710 (O_710,N_9100,N_9496);
and UO_711 (O_711,N_9635,N_9545);
or UO_712 (O_712,N_9621,N_9208);
or UO_713 (O_713,N_9582,N_9553);
nor UO_714 (O_714,N_9418,N_9902);
and UO_715 (O_715,N_9677,N_9859);
and UO_716 (O_716,N_9818,N_9588);
nor UO_717 (O_717,N_9593,N_9562);
nor UO_718 (O_718,N_9784,N_9302);
nor UO_719 (O_719,N_9657,N_9987);
or UO_720 (O_720,N_9545,N_9463);
nand UO_721 (O_721,N_9570,N_9576);
or UO_722 (O_722,N_9223,N_9713);
nor UO_723 (O_723,N_9976,N_9741);
nor UO_724 (O_724,N_9390,N_9167);
nand UO_725 (O_725,N_9434,N_9007);
xnor UO_726 (O_726,N_9261,N_9638);
nor UO_727 (O_727,N_9702,N_9564);
and UO_728 (O_728,N_9465,N_9605);
and UO_729 (O_729,N_9508,N_9117);
nand UO_730 (O_730,N_9186,N_9975);
nand UO_731 (O_731,N_9564,N_9338);
nor UO_732 (O_732,N_9037,N_9146);
or UO_733 (O_733,N_9081,N_9046);
nor UO_734 (O_734,N_9080,N_9685);
or UO_735 (O_735,N_9810,N_9438);
or UO_736 (O_736,N_9395,N_9177);
and UO_737 (O_737,N_9400,N_9365);
nand UO_738 (O_738,N_9646,N_9923);
nand UO_739 (O_739,N_9668,N_9515);
or UO_740 (O_740,N_9925,N_9793);
and UO_741 (O_741,N_9615,N_9351);
nand UO_742 (O_742,N_9023,N_9053);
xnor UO_743 (O_743,N_9488,N_9418);
or UO_744 (O_744,N_9332,N_9695);
nor UO_745 (O_745,N_9957,N_9168);
nor UO_746 (O_746,N_9653,N_9807);
nor UO_747 (O_747,N_9578,N_9604);
nand UO_748 (O_748,N_9747,N_9985);
nor UO_749 (O_749,N_9245,N_9204);
nor UO_750 (O_750,N_9002,N_9443);
or UO_751 (O_751,N_9594,N_9249);
nor UO_752 (O_752,N_9134,N_9570);
and UO_753 (O_753,N_9698,N_9069);
nor UO_754 (O_754,N_9312,N_9289);
and UO_755 (O_755,N_9356,N_9832);
and UO_756 (O_756,N_9336,N_9123);
or UO_757 (O_757,N_9914,N_9787);
and UO_758 (O_758,N_9328,N_9230);
nand UO_759 (O_759,N_9246,N_9330);
or UO_760 (O_760,N_9564,N_9907);
and UO_761 (O_761,N_9628,N_9457);
nand UO_762 (O_762,N_9962,N_9320);
and UO_763 (O_763,N_9637,N_9148);
xor UO_764 (O_764,N_9517,N_9080);
xor UO_765 (O_765,N_9265,N_9585);
or UO_766 (O_766,N_9701,N_9583);
nor UO_767 (O_767,N_9982,N_9121);
nand UO_768 (O_768,N_9955,N_9900);
nor UO_769 (O_769,N_9869,N_9181);
nand UO_770 (O_770,N_9461,N_9408);
and UO_771 (O_771,N_9796,N_9791);
nor UO_772 (O_772,N_9685,N_9970);
or UO_773 (O_773,N_9654,N_9061);
nand UO_774 (O_774,N_9825,N_9303);
nand UO_775 (O_775,N_9599,N_9411);
nand UO_776 (O_776,N_9436,N_9607);
nand UO_777 (O_777,N_9057,N_9989);
and UO_778 (O_778,N_9312,N_9937);
and UO_779 (O_779,N_9596,N_9036);
and UO_780 (O_780,N_9835,N_9698);
and UO_781 (O_781,N_9453,N_9248);
or UO_782 (O_782,N_9514,N_9450);
or UO_783 (O_783,N_9187,N_9032);
nand UO_784 (O_784,N_9297,N_9667);
or UO_785 (O_785,N_9392,N_9796);
nor UO_786 (O_786,N_9578,N_9688);
nand UO_787 (O_787,N_9624,N_9655);
nand UO_788 (O_788,N_9397,N_9042);
nand UO_789 (O_789,N_9022,N_9521);
nor UO_790 (O_790,N_9342,N_9926);
xnor UO_791 (O_791,N_9753,N_9260);
or UO_792 (O_792,N_9173,N_9658);
nor UO_793 (O_793,N_9737,N_9921);
or UO_794 (O_794,N_9686,N_9621);
nand UO_795 (O_795,N_9471,N_9627);
nand UO_796 (O_796,N_9593,N_9183);
nand UO_797 (O_797,N_9289,N_9593);
nand UO_798 (O_798,N_9778,N_9393);
or UO_799 (O_799,N_9573,N_9177);
nor UO_800 (O_800,N_9797,N_9795);
or UO_801 (O_801,N_9349,N_9521);
xnor UO_802 (O_802,N_9247,N_9942);
or UO_803 (O_803,N_9927,N_9287);
nor UO_804 (O_804,N_9810,N_9012);
nor UO_805 (O_805,N_9125,N_9163);
and UO_806 (O_806,N_9984,N_9790);
or UO_807 (O_807,N_9361,N_9618);
or UO_808 (O_808,N_9554,N_9836);
nor UO_809 (O_809,N_9033,N_9708);
or UO_810 (O_810,N_9195,N_9885);
nor UO_811 (O_811,N_9550,N_9463);
or UO_812 (O_812,N_9926,N_9222);
and UO_813 (O_813,N_9138,N_9219);
nand UO_814 (O_814,N_9964,N_9550);
nor UO_815 (O_815,N_9869,N_9117);
or UO_816 (O_816,N_9298,N_9641);
and UO_817 (O_817,N_9181,N_9687);
or UO_818 (O_818,N_9450,N_9776);
xor UO_819 (O_819,N_9617,N_9198);
and UO_820 (O_820,N_9615,N_9913);
and UO_821 (O_821,N_9100,N_9365);
and UO_822 (O_822,N_9686,N_9850);
nor UO_823 (O_823,N_9564,N_9132);
and UO_824 (O_824,N_9642,N_9179);
or UO_825 (O_825,N_9480,N_9503);
or UO_826 (O_826,N_9199,N_9503);
and UO_827 (O_827,N_9568,N_9441);
nor UO_828 (O_828,N_9718,N_9214);
or UO_829 (O_829,N_9359,N_9658);
nor UO_830 (O_830,N_9780,N_9442);
nand UO_831 (O_831,N_9946,N_9427);
and UO_832 (O_832,N_9179,N_9875);
and UO_833 (O_833,N_9121,N_9136);
and UO_834 (O_834,N_9420,N_9118);
nor UO_835 (O_835,N_9950,N_9432);
xor UO_836 (O_836,N_9739,N_9949);
and UO_837 (O_837,N_9447,N_9985);
nor UO_838 (O_838,N_9240,N_9442);
nor UO_839 (O_839,N_9717,N_9234);
and UO_840 (O_840,N_9315,N_9807);
and UO_841 (O_841,N_9794,N_9252);
and UO_842 (O_842,N_9307,N_9111);
or UO_843 (O_843,N_9077,N_9536);
nor UO_844 (O_844,N_9513,N_9546);
or UO_845 (O_845,N_9036,N_9225);
nand UO_846 (O_846,N_9232,N_9817);
nor UO_847 (O_847,N_9450,N_9503);
nand UO_848 (O_848,N_9425,N_9621);
or UO_849 (O_849,N_9940,N_9239);
nor UO_850 (O_850,N_9689,N_9987);
and UO_851 (O_851,N_9150,N_9341);
nand UO_852 (O_852,N_9276,N_9534);
and UO_853 (O_853,N_9229,N_9443);
xnor UO_854 (O_854,N_9237,N_9111);
and UO_855 (O_855,N_9335,N_9064);
or UO_856 (O_856,N_9171,N_9968);
and UO_857 (O_857,N_9645,N_9310);
and UO_858 (O_858,N_9609,N_9931);
nand UO_859 (O_859,N_9916,N_9420);
or UO_860 (O_860,N_9518,N_9361);
and UO_861 (O_861,N_9177,N_9569);
and UO_862 (O_862,N_9757,N_9040);
or UO_863 (O_863,N_9904,N_9778);
nor UO_864 (O_864,N_9609,N_9870);
nor UO_865 (O_865,N_9437,N_9647);
nand UO_866 (O_866,N_9828,N_9648);
nor UO_867 (O_867,N_9697,N_9899);
or UO_868 (O_868,N_9868,N_9758);
or UO_869 (O_869,N_9319,N_9194);
nand UO_870 (O_870,N_9953,N_9312);
xor UO_871 (O_871,N_9160,N_9383);
or UO_872 (O_872,N_9533,N_9404);
nor UO_873 (O_873,N_9566,N_9706);
nand UO_874 (O_874,N_9689,N_9118);
nand UO_875 (O_875,N_9887,N_9790);
or UO_876 (O_876,N_9555,N_9104);
or UO_877 (O_877,N_9616,N_9588);
and UO_878 (O_878,N_9475,N_9786);
or UO_879 (O_879,N_9573,N_9679);
nand UO_880 (O_880,N_9195,N_9732);
nand UO_881 (O_881,N_9345,N_9944);
nor UO_882 (O_882,N_9267,N_9696);
nor UO_883 (O_883,N_9391,N_9785);
nor UO_884 (O_884,N_9431,N_9264);
and UO_885 (O_885,N_9093,N_9844);
and UO_886 (O_886,N_9124,N_9995);
nand UO_887 (O_887,N_9433,N_9773);
and UO_888 (O_888,N_9512,N_9608);
nand UO_889 (O_889,N_9055,N_9848);
and UO_890 (O_890,N_9642,N_9180);
nor UO_891 (O_891,N_9843,N_9209);
or UO_892 (O_892,N_9560,N_9376);
nor UO_893 (O_893,N_9787,N_9337);
nand UO_894 (O_894,N_9622,N_9310);
or UO_895 (O_895,N_9184,N_9053);
nor UO_896 (O_896,N_9294,N_9219);
xor UO_897 (O_897,N_9899,N_9489);
or UO_898 (O_898,N_9448,N_9332);
nor UO_899 (O_899,N_9681,N_9367);
nor UO_900 (O_900,N_9367,N_9747);
and UO_901 (O_901,N_9094,N_9873);
nand UO_902 (O_902,N_9880,N_9343);
and UO_903 (O_903,N_9119,N_9155);
nand UO_904 (O_904,N_9255,N_9868);
or UO_905 (O_905,N_9975,N_9507);
nand UO_906 (O_906,N_9420,N_9357);
or UO_907 (O_907,N_9592,N_9468);
or UO_908 (O_908,N_9373,N_9647);
and UO_909 (O_909,N_9070,N_9052);
nand UO_910 (O_910,N_9949,N_9110);
xor UO_911 (O_911,N_9386,N_9680);
nand UO_912 (O_912,N_9764,N_9780);
nand UO_913 (O_913,N_9738,N_9113);
nor UO_914 (O_914,N_9561,N_9210);
nor UO_915 (O_915,N_9344,N_9780);
nor UO_916 (O_916,N_9185,N_9251);
nor UO_917 (O_917,N_9854,N_9939);
or UO_918 (O_918,N_9384,N_9287);
nor UO_919 (O_919,N_9593,N_9150);
nor UO_920 (O_920,N_9302,N_9125);
nor UO_921 (O_921,N_9587,N_9058);
nand UO_922 (O_922,N_9815,N_9788);
and UO_923 (O_923,N_9258,N_9454);
and UO_924 (O_924,N_9887,N_9928);
xor UO_925 (O_925,N_9105,N_9209);
nand UO_926 (O_926,N_9066,N_9340);
and UO_927 (O_927,N_9650,N_9785);
and UO_928 (O_928,N_9868,N_9192);
nand UO_929 (O_929,N_9761,N_9129);
nand UO_930 (O_930,N_9924,N_9655);
or UO_931 (O_931,N_9850,N_9960);
or UO_932 (O_932,N_9829,N_9624);
xor UO_933 (O_933,N_9501,N_9999);
or UO_934 (O_934,N_9614,N_9491);
and UO_935 (O_935,N_9303,N_9380);
nand UO_936 (O_936,N_9978,N_9910);
and UO_937 (O_937,N_9975,N_9287);
and UO_938 (O_938,N_9394,N_9880);
nand UO_939 (O_939,N_9738,N_9262);
nor UO_940 (O_940,N_9479,N_9014);
nor UO_941 (O_941,N_9530,N_9034);
xor UO_942 (O_942,N_9539,N_9361);
or UO_943 (O_943,N_9036,N_9818);
nor UO_944 (O_944,N_9498,N_9316);
or UO_945 (O_945,N_9850,N_9093);
nor UO_946 (O_946,N_9423,N_9927);
and UO_947 (O_947,N_9006,N_9099);
and UO_948 (O_948,N_9188,N_9669);
or UO_949 (O_949,N_9651,N_9652);
and UO_950 (O_950,N_9633,N_9712);
or UO_951 (O_951,N_9070,N_9432);
and UO_952 (O_952,N_9812,N_9095);
or UO_953 (O_953,N_9125,N_9516);
and UO_954 (O_954,N_9243,N_9180);
nand UO_955 (O_955,N_9295,N_9975);
nand UO_956 (O_956,N_9248,N_9819);
nor UO_957 (O_957,N_9748,N_9229);
nor UO_958 (O_958,N_9674,N_9256);
nand UO_959 (O_959,N_9549,N_9685);
or UO_960 (O_960,N_9600,N_9725);
and UO_961 (O_961,N_9520,N_9745);
nand UO_962 (O_962,N_9003,N_9878);
or UO_963 (O_963,N_9206,N_9150);
xor UO_964 (O_964,N_9846,N_9608);
nor UO_965 (O_965,N_9313,N_9248);
and UO_966 (O_966,N_9885,N_9201);
or UO_967 (O_967,N_9876,N_9755);
or UO_968 (O_968,N_9381,N_9733);
and UO_969 (O_969,N_9670,N_9754);
or UO_970 (O_970,N_9126,N_9216);
xor UO_971 (O_971,N_9166,N_9417);
nand UO_972 (O_972,N_9710,N_9957);
nor UO_973 (O_973,N_9380,N_9699);
xor UO_974 (O_974,N_9866,N_9502);
nor UO_975 (O_975,N_9463,N_9899);
nor UO_976 (O_976,N_9845,N_9888);
or UO_977 (O_977,N_9262,N_9765);
or UO_978 (O_978,N_9373,N_9709);
or UO_979 (O_979,N_9863,N_9129);
nand UO_980 (O_980,N_9587,N_9803);
nand UO_981 (O_981,N_9414,N_9860);
and UO_982 (O_982,N_9917,N_9110);
nor UO_983 (O_983,N_9570,N_9122);
nand UO_984 (O_984,N_9627,N_9070);
nand UO_985 (O_985,N_9483,N_9157);
or UO_986 (O_986,N_9822,N_9612);
and UO_987 (O_987,N_9325,N_9293);
and UO_988 (O_988,N_9179,N_9323);
and UO_989 (O_989,N_9872,N_9587);
and UO_990 (O_990,N_9103,N_9813);
or UO_991 (O_991,N_9106,N_9343);
or UO_992 (O_992,N_9756,N_9326);
or UO_993 (O_993,N_9053,N_9827);
nor UO_994 (O_994,N_9124,N_9071);
nor UO_995 (O_995,N_9036,N_9455);
nor UO_996 (O_996,N_9790,N_9612);
nor UO_997 (O_997,N_9467,N_9542);
nor UO_998 (O_998,N_9461,N_9468);
nand UO_999 (O_999,N_9585,N_9097);
or UO_1000 (O_1000,N_9185,N_9002);
nand UO_1001 (O_1001,N_9691,N_9160);
nor UO_1002 (O_1002,N_9187,N_9503);
or UO_1003 (O_1003,N_9010,N_9549);
xor UO_1004 (O_1004,N_9628,N_9796);
nor UO_1005 (O_1005,N_9020,N_9782);
nand UO_1006 (O_1006,N_9934,N_9738);
and UO_1007 (O_1007,N_9926,N_9106);
and UO_1008 (O_1008,N_9987,N_9207);
or UO_1009 (O_1009,N_9859,N_9897);
nor UO_1010 (O_1010,N_9730,N_9052);
nor UO_1011 (O_1011,N_9962,N_9707);
nor UO_1012 (O_1012,N_9062,N_9633);
nor UO_1013 (O_1013,N_9046,N_9542);
nor UO_1014 (O_1014,N_9943,N_9790);
or UO_1015 (O_1015,N_9127,N_9215);
xor UO_1016 (O_1016,N_9777,N_9539);
or UO_1017 (O_1017,N_9442,N_9956);
and UO_1018 (O_1018,N_9862,N_9774);
or UO_1019 (O_1019,N_9529,N_9886);
xor UO_1020 (O_1020,N_9521,N_9498);
xor UO_1021 (O_1021,N_9973,N_9996);
nand UO_1022 (O_1022,N_9193,N_9711);
nand UO_1023 (O_1023,N_9520,N_9733);
nor UO_1024 (O_1024,N_9481,N_9320);
xnor UO_1025 (O_1025,N_9185,N_9149);
nor UO_1026 (O_1026,N_9624,N_9694);
or UO_1027 (O_1027,N_9011,N_9155);
or UO_1028 (O_1028,N_9955,N_9083);
nand UO_1029 (O_1029,N_9966,N_9888);
nor UO_1030 (O_1030,N_9664,N_9212);
nand UO_1031 (O_1031,N_9888,N_9682);
xor UO_1032 (O_1032,N_9368,N_9330);
and UO_1033 (O_1033,N_9295,N_9312);
nand UO_1034 (O_1034,N_9438,N_9898);
nor UO_1035 (O_1035,N_9151,N_9431);
nand UO_1036 (O_1036,N_9415,N_9535);
or UO_1037 (O_1037,N_9646,N_9491);
nor UO_1038 (O_1038,N_9885,N_9712);
nand UO_1039 (O_1039,N_9912,N_9954);
and UO_1040 (O_1040,N_9775,N_9336);
xor UO_1041 (O_1041,N_9324,N_9909);
nor UO_1042 (O_1042,N_9875,N_9378);
and UO_1043 (O_1043,N_9110,N_9029);
and UO_1044 (O_1044,N_9835,N_9192);
xnor UO_1045 (O_1045,N_9162,N_9420);
or UO_1046 (O_1046,N_9206,N_9371);
xor UO_1047 (O_1047,N_9856,N_9402);
and UO_1048 (O_1048,N_9588,N_9934);
nand UO_1049 (O_1049,N_9835,N_9535);
nor UO_1050 (O_1050,N_9655,N_9047);
nand UO_1051 (O_1051,N_9558,N_9104);
nor UO_1052 (O_1052,N_9297,N_9859);
nand UO_1053 (O_1053,N_9289,N_9223);
nand UO_1054 (O_1054,N_9571,N_9203);
and UO_1055 (O_1055,N_9691,N_9366);
and UO_1056 (O_1056,N_9701,N_9014);
nand UO_1057 (O_1057,N_9009,N_9340);
nand UO_1058 (O_1058,N_9152,N_9124);
or UO_1059 (O_1059,N_9162,N_9025);
xnor UO_1060 (O_1060,N_9788,N_9399);
or UO_1061 (O_1061,N_9726,N_9047);
xor UO_1062 (O_1062,N_9017,N_9719);
or UO_1063 (O_1063,N_9507,N_9576);
nand UO_1064 (O_1064,N_9311,N_9009);
xnor UO_1065 (O_1065,N_9678,N_9372);
nor UO_1066 (O_1066,N_9555,N_9546);
or UO_1067 (O_1067,N_9838,N_9539);
nor UO_1068 (O_1068,N_9040,N_9722);
or UO_1069 (O_1069,N_9993,N_9060);
or UO_1070 (O_1070,N_9935,N_9662);
nor UO_1071 (O_1071,N_9288,N_9399);
and UO_1072 (O_1072,N_9177,N_9830);
or UO_1073 (O_1073,N_9400,N_9441);
or UO_1074 (O_1074,N_9295,N_9062);
or UO_1075 (O_1075,N_9558,N_9460);
xnor UO_1076 (O_1076,N_9839,N_9364);
and UO_1077 (O_1077,N_9200,N_9334);
nor UO_1078 (O_1078,N_9589,N_9598);
nor UO_1079 (O_1079,N_9971,N_9207);
and UO_1080 (O_1080,N_9698,N_9553);
and UO_1081 (O_1081,N_9157,N_9041);
and UO_1082 (O_1082,N_9620,N_9786);
and UO_1083 (O_1083,N_9537,N_9303);
and UO_1084 (O_1084,N_9888,N_9000);
or UO_1085 (O_1085,N_9394,N_9574);
nor UO_1086 (O_1086,N_9323,N_9638);
or UO_1087 (O_1087,N_9913,N_9434);
nand UO_1088 (O_1088,N_9253,N_9340);
and UO_1089 (O_1089,N_9224,N_9391);
and UO_1090 (O_1090,N_9931,N_9451);
nand UO_1091 (O_1091,N_9700,N_9213);
xor UO_1092 (O_1092,N_9506,N_9005);
nand UO_1093 (O_1093,N_9648,N_9484);
nor UO_1094 (O_1094,N_9371,N_9897);
nand UO_1095 (O_1095,N_9341,N_9745);
nand UO_1096 (O_1096,N_9583,N_9087);
and UO_1097 (O_1097,N_9823,N_9214);
nor UO_1098 (O_1098,N_9259,N_9147);
nor UO_1099 (O_1099,N_9197,N_9083);
nor UO_1100 (O_1100,N_9049,N_9686);
nand UO_1101 (O_1101,N_9846,N_9823);
and UO_1102 (O_1102,N_9688,N_9450);
nand UO_1103 (O_1103,N_9353,N_9599);
and UO_1104 (O_1104,N_9261,N_9180);
and UO_1105 (O_1105,N_9606,N_9546);
and UO_1106 (O_1106,N_9438,N_9411);
or UO_1107 (O_1107,N_9173,N_9693);
or UO_1108 (O_1108,N_9948,N_9900);
and UO_1109 (O_1109,N_9359,N_9862);
or UO_1110 (O_1110,N_9926,N_9068);
or UO_1111 (O_1111,N_9398,N_9533);
nand UO_1112 (O_1112,N_9268,N_9494);
and UO_1113 (O_1113,N_9017,N_9728);
nor UO_1114 (O_1114,N_9454,N_9715);
nand UO_1115 (O_1115,N_9236,N_9524);
or UO_1116 (O_1116,N_9481,N_9689);
or UO_1117 (O_1117,N_9554,N_9197);
and UO_1118 (O_1118,N_9143,N_9915);
and UO_1119 (O_1119,N_9231,N_9499);
nor UO_1120 (O_1120,N_9430,N_9971);
nor UO_1121 (O_1121,N_9496,N_9065);
or UO_1122 (O_1122,N_9470,N_9721);
and UO_1123 (O_1123,N_9280,N_9019);
or UO_1124 (O_1124,N_9784,N_9021);
nor UO_1125 (O_1125,N_9545,N_9882);
or UO_1126 (O_1126,N_9096,N_9433);
nand UO_1127 (O_1127,N_9516,N_9259);
nor UO_1128 (O_1128,N_9833,N_9515);
and UO_1129 (O_1129,N_9259,N_9012);
or UO_1130 (O_1130,N_9666,N_9234);
nand UO_1131 (O_1131,N_9288,N_9081);
nor UO_1132 (O_1132,N_9947,N_9884);
xor UO_1133 (O_1133,N_9084,N_9805);
nor UO_1134 (O_1134,N_9457,N_9046);
nor UO_1135 (O_1135,N_9034,N_9438);
nor UO_1136 (O_1136,N_9494,N_9872);
nand UO_1137 (O_1137,N_9171,N_9262);
or UO_1138 (O_1138,N_9583,N_9838);
nand UO_1139 (O_1139,N_9222,N_9212);
xnor UO_1140 (O_1140,N_9019,N_9693);
nand UO_1141 (O_1141,N_9453,N_9204);
xor UO_1142 (O_1142,N_9167,N_9770);
nor UO_1143 (O_1143,N_9579,N_9597);
or UO_1144 (O_1144,N_9777,N_9933);
nor UO_1145 (O_1145,N_9436,N_9537);
and UO_1146 (O_1146,N_9880,N_9243);
nand UO_1147 (O_1147,N_9154,N_9549);
nand UO_1148 (O_1148,N_9020,N_9378);
and UO_1149 (O_1149,N_9650,N_9763);
or UO_1150 (O_1150,N_9268,N_9255);
or UO_1151 (O_1151,N_9860,N_9133);
nand UO_1152 (O_1152,N_9788,N_9373);
nand UO_1153 (O_1153,N_9071,N_9097);
nor UO_1154 (O_1154,N_9629,N_9216);
xnor UO_1155 (O_1155,N_9265,N_9244);
or UO_1156 (O_1156,N_9833,N_9038);
nand UO_1157 (O_1157,N_9622,N_9484);
or UO_1158 (O_1158,N_9001,N_9174);
and UO_1159 (O_1159,N_9789,N_9925);
or UO_1160 (O_1160,N_9610,N_9825);
or UO_1161 (O_1161,N_9199,N_9352);
or UO_1162 (O_1162,N_9406,N_9476);
and UO_1163 (O_1163,N_9007,N_9625);
nand UO_1164 (O_1164,N_9634,N_9301);
nor UO_1165 (O_1165,N_9319,N_9610);
or UO_1166 (O_1166,N_9736,N_9063);
nor UO_1167 (O_1167,N_9451,N_9513);
nand UO_1168 (O_1168,N_9194,N_9076);
xnor UO_1169 (O_1169,N_9278,N_9968);
nor UO_1170 (O_1170,N_9188,N_9981);
nand UO_1171 (O_1171,N_9841,N_9475);
nand UO_1172 (O_1172,N_9765,N_9543);
nand UO_1173 (O_1173,N_9805,N_9401);
and UO_1174 (O_1174,N_9333,N_9695);
and UO_1175 (O_1175,N_9377,N_9755);
nand UO_1176 (O_1176,N_9643,N_9772);
nor UO_1177 (O_1177,N_9493,N_9719);
xor UO_1178 (O_1178,N_9430,N_9195);
nand UO_1179 (O_1179,N_9058,N_9929);
nor UO_1180 (O_1180,N_9683,N_9135);
nor UO_1181 (O_1181,N_9529,N_9057);
or UO_1182 (O_1182,N_9959,N_9215);
xnor UO_1183 (O_1183,N_9034,N_9620);
or UO_1184 (O_1184,N_9917,N_9130);
nor UO_1185 (O_1185,N_9150,N_9735);
nor UO_1186 (O_1186,N_9854,N_9922);
nand UO_1187 (O_1187,N_9263,N_9856);
nand UO_1188 (O_1188,N_9249,N_9206);
nand UO_1189 (O_1189,N_9979,N_9975);
xnor UO_1190 (O_1190,N_9445,N_9563);
or UO_1191 (O_1191,N_9333,N_9322);
and UO_1192 (O_1192,N_9863,N_9577);
and UO_1193 (O_1193,N_9211,N_9802);
and UO_1194 (O_1194,N_9908,N_9565);
nor UO_1195 (O_1195,N_9977,N_9906);
or UO_1196 (O_1196,N_9382,N_9330);
nand UO_1197 (O_1197,N_9721,N_9118);
nor UO_1198 (O_1198,N_9784,N_9043);
nand UO_1199 (O_1199,N_9435,N_9395);
xor UO_1200 (O_1200,N_9198,N_9291);
nand UO_1201 (O_1201,N_9791,N_9448);
or UO_1202 (O_1202,N_9719,N_9413);
nand UO_1203 (O_1203,N_9554,N_9546);
or UO_1204 (O_1204,N_9755,N_9523);
nand UO_1205 (O_1205,N_9956,N_9495);
and UO_1206 (O_1206,N_9672,N_9580);
and UO_1207 (O_1207,N_9131,N_9015);
or UO_1208 (O_1208,N_9370,N_9735);
nor UO_1209 (O_1209,N_9665,N_9350);
and UO_1210 (O_1210,N_9887,N_9938);
or UO_1211 (O_1211,N_9538,N_9450);
nor UO_1212 (O_1212,N_9344,N_9100);
and UO_1213 (O_1213,N_9140,N_9864);
nor UO_1214 (O_1214,N_9390,N_9059);
xnor UO_1215 (O_1215,N_9693,N_9034);
xnor UO_1216 (O_1216,N_9606,N_9422);
nand UO_1217 (O_1217,N_9046,N_9328);
xnor UO_1218 (O_1218,N_9383,N_9422);
nand UO_1219 (O_1219,N_9459,N_9796);
or UO_1220 (O_1220,N_9129,N_9843);
and UO_1221 (O_1221,N_9071,N_9301);
nand UO_1222 (O_1222,N_9260,N_9987);
nand UO_1223 (O_1223,N_9367,N_9305);
xor UO_1224 (O_1224,N_9177,N_9201);
and UO_1225 (O_1225,N_9438,N_9177);
and UO_1226 (O_1226,N_9055,N_9408);
and UO_1227 (O_1227,N_9577,N_9327);
or UO_1228 (O_1228,N_9274,N_9366);
nor UO_1229 (O_1229,N_9545,N_9809);
nor UO_1230 (O_1230,N_9127,N_9196);
and UO_1231 (O_1231,N_9173,N_9366);
nor UO_1232 (O_1232,N_9993,N_9957);
nand UO_1233 (O_1233,N_9134,N_9319);
nand UO_1234 (O_1234,N_9163,N_9208);
nor UO_1235 (O_1235,N_9762,N_9600);
nand UO_1236 (O_1236,N_9670,N_9024);
nor UO_1237 (O_1237,N_9721,N_9269);
nand UO_1238 (O_1238,N_9514,N_9905);
nor UO_1239 (O_1239,N_9197,N_9143);
nand UO_1240 (O_1240,N_9402,N_9918);
nand UO_1241 (O_1241,N_9124,N_9135);
nand UO_1242 (O_1242,N_9564,N_9806);
nand UO_1243 (O_1243,N_9471,N_9429);
or UO_1244 (O_1244,N_9056,N_9405);
xnor UO_1245 (O_1245,N_9521,N_9839);
nand UO_1246 (O_1246,N_9998,N_9694);
nor UO_1247 (O_1247,N_9816,N_9812);
nor UO_1248 (O_1248,N_9472,N_9083);
nor UO_1249 (O_1249,N_9704,N_9326);
xor UO_1250 (O_1250,N_9487,N_9438);
or UO_1251 (O_1251,N_9439,N_9263);
nor UO_1252 (O_1252,N_9434,N_9879);
and UO_1253 (O_1253,N_9651,N_9650);
nand UO_1254 (O_1254,N_9161,N_9587);
or UO_1255 (O_1255,N_9869,N_9248);
nand UO_1256 (O_1256,N_9459,N_9083);
nor UO_1257 (O_1257,N_9353,N_9192);
nor UO_1258 (O_1258,N_9371,N_9308);
nand UO_1259 (O_1259,N_9551,N_9554);
nor UO_1260 (O_1260,N_9337,N_9388);
nand UO_1261 (O_1261,N_9138,N_9465);
nor UO_1262 (O_1262,N_9668,N_9519);
or UO_1263 (O_1263,N_9957,N_9144);
nor UO_1264 (O_1264,N_9134,N_9840);
and UO_1265 (O_1265,N_9416,N_9114);
nor UO_1266 (O_1266,N_9078,N_9689);
or UO_1267 (O_1267,N_9537,N_9736);
and UO_1268 (O_1268,N_9721,N_9354);
xnor UO_1269 (O_1269,N_9515,N_9719);
and UO_1270 (O_1270,N_9260,N_9150);
nor UO_1271 (O_1271,N_9577,N_9872);
or UO_1272 (O_1272,N_9473,N_9949);
or UO_1273 (O_1273,N_9799,N_9390);
and UO_1274 (O_1274,N_9193,N_9318);
and UO_1275 (O_1275,N_9033,N_9895);
and UO_1276 (O_1276,N_9098,N_9853);
or UO_1277 (O_1277,N_9190,N_9185);
or UO_1278 (O_1278,N_9260,N_9879);
nand UO_1279 (O_1279,N_9561,N_9346);
nor UO_1280 (O_1280,N_9709,N_9358);
and UO_1281 (O_1281,N_9196,N_9986);
nand UO_1282 (O_1282,N_9611,N_9985);
xor UO_1283 (O_1283,N_9700,N_9143);
or UO_1284 (O_1284,N_9414,N_9153);
nor UO_1285 (O_1285,N_9007,N_9486);
or UO_1286 (O_1286,N_9823,N_9830);
nor UO_1287 (O_1287,N_9119,N_9495);
or UO_1288 (O_1288,N_9550,N_9946);
nor UO_1289 (O_1289,N_9923,N_9354);
and UO_1290 (O_1290,N_9732,N_9706);
or UO_1291 (O_1291,N_9121,N_9741);
nand UO_1292 (O_1292,N_9076,N_9538);
or UO_1293 (O_1293,N_9779,N_9215);
and UO_1294 (O_1294,N_9269,N_9038);
nand UO_1295 (O_1295,N_9166,N_9334);
and UO_1296 (O_1296,N_9595,N_9599);
nand UO_1297 (O_1297,N_9138,N_9867);
nand UO_1298 (O_1298,N_9320,N_9570);
and UO_1299 (O_1299,N_9623,N_9182);
and UO_1300 (O_1300,N_9413,N_9621);
and UO_1301 (O_1301,N_9854,N_9034);
and UO_1302 (O_1302,N_9927,N_9436);
xor UO_1303 (O_1303,N_9852,N_9054);
or UO_1304 (O_1304,N_9253,N_9348);
xnor UO_1305 (O_1305,N_9338,N_9950);
nand UO_1306 (O_1306,N_9529,N_9449);
nor UO_1307 (O_1307,N_9118,N_9629);
xnor UO_1308 (O_1308,N_9597,N_9743);
or UO_1309 (O_1309,N_9091,N_9480);
or UO_1310 (O_1310,N_9869,N_9936);
nand UO_1311 (O_1311,N_9147,N_9320);
nand UO_1312 (O_1312,N_9054,N_9166);
nand UO_1313 (O_1313,N_9603,N_9878);
or UO_1314 (O_1314,N_9650,N_9331);
nand UO_1315 (O_1315,N_9175,N_9099);
nand UO_1316 (O_1316,N_9220,N_9263);
and UO_1317 (O_1317,N_9481,N_9026);
or UO_1318 (O_1318,N_9733,N_9134);
and UO_1319 (O_1319,N_9153,N_9445);
or UO_1320 (O_1320,N_9143,N_9032);
nor UO_1321 (O_1321,N_9392,N_9565);
nand UO_1322 (O_1322,N_9114,N_9748);
and UO_1323 (O_1323,N_9901,N_9023);
nand UO_1324 (O_1324,N_9383,N_9135);
nand UO_1325 (O_1325,N_9169,N_9757);
nor UO_1326 (O_1326,N_9381,N_9309);
nor UO_1327 (O_1327,N_9307,N_9515);
nand UO_1328 (O_1328,N_9025,N_9827);
and UO_1329 (O_1329,N_9086,N_9481);
and UO_1330 (O_1330,N_9013,N_9756);
nor UO_1331 (O_1331,N_9662,N_9495);
and UO_1332 (O_1332,N_9491,N_9851);
nand UO_1333 (O_1333,N_9370,N_9900);
or UO_1334 (O_1334,N_9122,N_9168);
or UO_1335 (O_1335,N_9648,N_9145);
and UO_1336 (O_1336,N_9386,N_9067);
xnor UO_1337 (O_1337,N_9859,N_9023);
nor UO_1338 (O_1338,N_9852,N_9769);
nand UO_1339 (O_1339,N_9947,N_9151);
and UO_1340 (O_1340,N_9717,N_9347);
or UO_1341 (O_1341,N_9992,N_9946);
nor UO_1342 (O_1342,N_9281,N_9884);
and UO_1343 (O_1343,N_9341,N_9076);
or UO_1344 (O_1344,N_9859,N_9902);
or UO_1345 (O_1345,N_9876,N_9368);
nand UO_1346 (O_1346,N_9297,N_9202);
xor UO_1347 (O_1347,N_9227,N_9149);
and UO_1348 (O_1348,N_9257,N_9064);
and UO_1349 (O_1349,N_9110,N_9107);
xnor UO_1350 (O_1350,N_9414,N_9960);
xor UO_1351 (O_1351,N_9658,N_9150);
xor UO_1352 (O_1352,N_9587,N_9723);
nand UO_1353 (O_1353,N_9172,N_9372);
and UO_1354 (O_1354,N_9613,N_9527);
or UO_1355 (O_1355,N_9227,N_9808);
xor UO_1356 (O_1356,N_9298,N_9741);
nor UO_1357 (O_1357,N_9212,N_9453);
nor UO_1358 (O_1358,N_9600,N_9929);
nor UO_1359 (O_1359,N_9098,N_9988);
nor UO_1360 (O_1360,N_9226,N_9456);
nand UO_1361 (O_1361,N_9201,N_9352);
xnor UO_1362 (O_1362,N_9220,N_9920);
and UO_1363 (O_1363,N_9292,N_9764);
nand UO_1364 (O_1364,N_9330,N_9788);
or UO_1365 (O_1365,N_9065,N_9302);
nor UO_1366 (O_1366,N_9268,N_9057);
nand UO_1367 (O_1367,N_9334,N_9412);
and UO_1368 (O_1368,N_9332,N_9781);
and UO_1369 (O_1369,N_9347,N_9707);
or UO_1370 (O_1370,N_9729,N_9954);
and UO_1371 (O_1371,N_9462,N_9182);
or UO_1372 (O_1372,N_9085,N_9816);
and UO_1373 (O_1373,N_9714,N_9526);
and UO_1374 (O_1374,N_9619,N_9247);
xnor UO_1375 (O_1375,N_9906,N_9214);
nand UO_1376 (O_1376,N_9215,N_9375);
or UO_1377 (O_1377,N_9172,N_9249);
nor UO_1378 (O_1378,N_9562,N_9335);
nand UO_1379 (O_1379,N_9610,N_9591);
or UO_1380 (O_1380,N_9069,N_9411);
nand UO_1381 (O_1381,N_9277,N_9819);
nand UO_1382 (O_1382,N_9319,N_9582);
nor UO_1383 (O_1383,N_9219,N_9119);
nand UO_1384 (O_1384,N_9584,N_9656);
nand UO_1385 (O_1385,N_9771,N_9586);
and UO_1386 (O_1386,N_9468,N_9664);
nor UO_1387 (O_1387,N_9752,N_9109);
and UO_1388 (O_1388,N_9891,N_9211);
and UO_1389 (O_1389,N_9455,N_9938);
nand UO_1390 (O_1390,N_9918,N_9878);
and UO_1391 (O_1391,N_9695,N_9014);
or UO_1392 (O_1392,N_9045,N_9292);
nand UO_1393 (O_1393,N_9083,N_9828);
and UO_1394 (O_1394,N_9020,N_9139);
xnor UO_1395 (O_1395,N_9448,N_9973);
and UO_1396 (O_1396,N_9422,N_9823);
nor UO_1397 (O_1397,N_9548,N_9227);
nor UO_1398 (O_1398,N_9433,N_9589);
nor UO_1399 (O_1399,N_9910,N_9368);
nor UO_1400 (O_1400,N_9142,N_9772);
and UO_1401 (O_1401,N_9798,N_9467);
and UO_1402 (O_1402,N_9734,N_9146);
nand UO_1403 (O_1403,N_9181,N_9325);
nor UO_1404 (O_1404,N_9645,N_9603);
or UO_1405 (O_1405,N_9669,N_9216);
and UO_1406 (O_1406,N_9930,N_9641);
nand UO_1407 (O_1407,N_9042,N_9524);
or UO_1408 (O_1408,N_9177,N_9687);
nand UO_1409 (O_1409,N_9478,N_9211);
or UO_1410 (O_1410,N_9989,N_9378);
nor UO_1411 (O_1411,N_9887,N_9179);
or UO_1412 (O_1412,N_9109,N_9117);
or UO_1413 (O_1413,N_9533,N_9282);
nand UO_1414 (O_1414,N_9599,N_9102);
and UO_1415 (O_1415,N_9518,N_9306);
and UO_1416 (O_1416,N_9881,N_9400);
and UO_1417 (O_1417,N_9072,N_9783);
or UO_1418 (O_1418,N_9371,N_9105);
nor UO_1419 (O_1419,N_9174,N_9102);
nand UO_1420 (O_1420,N_9924,N_9200);
or UO_1421 (O_1421,N_9530,N_9322);
and UO_1422 (O_1422,N_9552,N_9431);
nand UO_1423 (O_1423,N_9839,N_9005);
nor UO_1424 (O_1424,N_9324,N_9639);
or UO_1425 (O_1425,N_9659,N_9896);
xor UO_1426 (O_1426,N_9597,N_9165);
and UO_1427 (O_1427,N_9763,N_9986);
or UO_1428 (O_1428,N_9759,N_9651);
nand UO_1429 (O_1429,N_9344,N_9238);
nand UO_1430 (O_1430,N_9704,N_9153);
or UO_1431 (O_1431,N_9089,N_9743);
xnor UO_1432 (O_1432,N_9661,N_9545);
nand UO_1433 (O_1433,N_9910,N_9843);
nand UO_1434 (O_1434,N_9683,N_9100);
nor UO_1435 (O_1435,N_9704,N_9206);
or UO_1436 (O_1436,N_9972,N_9479);
nor UO_1437 (O_1437,N_9789,N_9609);
or UO_1438 (O_1438,N_9911,N_9060);
or UO_1439 (O_1439,N_9619,N_9928);
or UO_1440 (O_1440,N_9425,N_9106);
and UO_1441 (O_1441,N_9319,N_9960);
nor UO_1442 (O_1442,N_9630,N_9543);
or UO_1443 (O_1443,N_9640,N_9508);
xor UO_1444 (O_1444,N_9109,N_9530);
nand UO_1445 (O_1445,N_9661,N_9152);
nor UO_1446 (O_1446,N_9457,N_9434);
nor UO_1447 (O_1447,N_9223,N_9771);
and UO_1448 (O_1448,N_9931,N_9919);
nand UO_1449 (O_1449,N_9128,N_9411);
and UO_1450 (O_1450,N_9380,N_9873);
or UO_1451 (O_1451,N_9680,N_9561);
nor UO_1452 (O_1452,N_9993,N_9151);
and UO_1453 (O_1453,N_9255,N_9433);
and UO_1454 (O_1454,N_9335,N_9100);
and UO_1455 (O_1455,N_9147,N_9537);
nor UO_1456 (O_1456,N_9431,N_9256);
or UO_1457 (O_1457,N_9614,N_9527);
nor UO_1458 (O_1458,N_9939,N_9442);
nand UO_1459 (O_1459,N_9892,N_9836);
and UO_1460 (O_1460,N_9489,N_9507);
nor UO_1461 (O_1461,N_9711,N_9393);
and UO_1462 (O_1462,N_9937,N_9975);
nand UO_1463 (O_1463,N_9153,N_9459);
nand UO_1464 (O_1464,N_9579,N_9199);
and UO_1465 (O_1465,N_9849,N_9636);
nand UO_1466 (O_1466,N_9178,N_9838);
nand UO_1467 (O_1467,N_9344,N_9579);
and UO_1468 (O_1468,N_9082,N_9098);
nor UO_1469 (O_1469,N_9713,N_9676);
nand UO_1470 (O_1470,N_9200,N_9263);
xor UO_1471 (O_1471,N_9992,N_9184);
and UO_1472 (O_1472,N_9330,N_9622);
nand UO_1473 (O_1473,N_9271,N_9954);
nand UO_1474 (O_1474,N_9274,N_9976);
nor UO_1475 (O_1475,N_9793,N_9478);
nand UO_1476 (O_1476,N_9054,N_9010);
nor UO_1477 (O_1477,N_9751,N_9025);
nor UO_1478 (O_1478,N_9222,N_9410);
and UO_1479 (O_1479,N_9758,N_9336);
xor UO_1480 (O_1480,N_9452,N_9308);
nor UO_1481 (O_1481,N_9475,N_9090);
nor UO_1482 (O_1482,N_9578,N_9133);
nor UO_1483 (O_1483,N_9446,N_9229);
and UO_1484 (O_1484,N_9994,N_9936);
and UO_1485 (O_1485,N_9136,N_9883);
or UO_1486 (O_1486,N_9207,N_9703);
or UO_1487 (O_1487,N_9041,N_9090);
nor UO_1488 (O_1488,N_9621,N_9054);
and UO_1489 (O_1489,N_9401,N_9784);
nand UO_1490 (O_1490,N_9428,N_9095);
nand UO_1491 (O_1491,N_9195,N_9691);
nor UO_1492 (O_1492,N_9631,N_9693);
or UO_1493 (O_1493,N_9869,N_9487);
xor UO_1494 (O_1494,N_9738,N_9897);
or UO_1495 (O_1495,N_9161,N_9680);
nand UO_1496 (O_1496,N_9703,N_9276);
and UO_1497 (O_1497,N_9335,N_9363);
or UO_1498 (O_1498,N_9010,N_9808);
or UO_1499 (O_1499,N_9416,N_9407);
endmodule