module basic_500_3000_500_5_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_288,In_184);
or U1 (N_1,In_214,In_438);
and U2 (N_2,In_328,In_194);
nor U3 (N_3,In_443,In_414);
or U4 (N_4,In_499,In_221);
nand U5 (N_5,In_108,In_485);
or U6 (N_6,In_199,In_121);
nor U7 (N_7,In_62,In_31);
and U8 (N_8,In_212,In_81);
nor U9 (N_9,In_493,In_316);
or U10 (N_10,In_147,In_332);
or U11 (N_11,In_222,In_357);
and U12 (N_12,In_96,In_181);
nand U13 (N_13,In_176,In_336);
and U14 (N_14,In_454,In_489);
or U15 (N_15,In_282,In_14);
and U16 (N_16,In_123,In_48);
nand U17 (N_17,In_384,In_177);
nand U18 (N_18,In_143,In_205);
or U19 (N_19,In_124,In_141);
or U20 (N_20,In_428,In_75);
xor U21 (N_21,In_186,In_308);
or U22 (N_22,In_231,In_439);
and U23 (N_23,In_87,In_202);
and U24 (N_24,In_68,In_317);
nand U25 (N_25,In_174,In_497);
nand U26 (N_26,In_410,In_241);
nor U27 (N_27,In_109,In_498);
and U28 (N_28,In_496,In_269);
nor U29 (N_29,In_382,In_34);
nor U30 (N_30,In_298,In_99);
and U31 (N_31,In_237,In_460);
or U32 (N_32,In_230,In_245);
nand U33 (N_33,In_260,In_18);
nand U34 (N_34,In_315,In_37);
nor U35 (N_35,In_66,In_465);
and U36 (N_36,In_26,In_393);
or U37 (N_37,In_236,In_133);
or U38 (N_38,In_254,In_126);
nand U39 (N_39,In_4,In_193);
or U40 (N_40,In_275,In_165);
and U41 (N_41,In_9,In_69);
and U42 (N_42,In_183,In_197);
or U43 (N_43,In_94,In_137);
or U44 (N_44,In_268,In_156);
nor U45 (N_45,In_425,In_235);
nor U46 (N_46,In_159,In_368);
or U47 (N_47,In_430,In_115);
nor U48 (N_48,In_453,In_10);
or U49 (N_49,In_82,In_135);
nor U50 (N_50,In_243,In_29);
and U51 (N_51,In_385,In_50);
and U52 (N_52,In_293,In_93);
or U53 (N_53,In_35,In_140);
or U54 (N_54,In_11,In_191);
or U55 (N_55,In_257,In_487);
nor U56 (N_56,In_389,In_234);
nor U57 (N_57,In_111,In_103);
and U58 (N_58,In_210,In_355);
and U59 (N_59,In_219,In_118);
nor U60 (N_60,In_359,In_290);
nor U61 (N_61,In_432,In_74);
nor U62 (N_62,In_362,In_60);
nand U63 (N_63,In_131,In_461);
nor U64 (N_64,In_417,In_415);
nor U65 (N_65,In_155,In_311);
nor U66 (N_66,In_40,In_3);
nand U67 (N_67,In_217,In_195);
or U68 (N_68,In_441,In_449);
or U69 (N_69,In_23,In_365);
nor U70 (N_70,In_407,In_426);
nand U71 (N_71,In_240,In_46);
and U72 (N_72,In_476,In_271);
nor U73 (N_73,In_451,In_470);
or U74 (N_74,In_166,In_139);
and U75 (N_75,In_30,In_39);
or U76 (N_76,In_480,In_247);
and U77 (N_77,In_347,In_89);
or U78 (N_78,In_100,In_434);
and U79 (N_79,In_397,In_161);
nand U80 (N_80,In_283,In_180);
nor U81 (N_81,In_264,In_302);
or U82 (N_82,In_279,In_483);
nand U83 (N_83,In_20,In_276);
nor U84 (N_84,In_286,In_80);
and U85 (N_85,In_261,In_253);
nand U86 (N_86,In_297,In_255);
and U87 (N_87,In_0,In_95);
nand U88 (N_88,In_200,In_277);
nor U89 (N_89,In_201,In_471);
nor U90 (N_90,In_128,In_420);
or U91 (N_91,In_112,In_452);
or U92 (N_92,In_361,In_378);
and U93 (N_93,In_296,In_19);
and U94 (N_94,In_381,In_63);
or U95 (N_95,In_320,In_303);
and U96 (N_96,In_479,In_204);
or U97 (N_97,In_113,In_185);
and U98 (N_98,In_446,In_252);
nor U99 (N_99,In_206,In_188);
and U100 (N_100,In_49,In_73);
nor U101 (N_101,In_345,In_179);
nor U102 (N_102,In_225,In_85);
nor U103 (N_103,In_72,In_43);
and U104 (N_104,In_450,In_468);
nand U105 (N_105,In_292,In_91);
nor U106 (N_106,In_70,In_334);
nand U107 (N_107,In_348,In_171);
nor U108 (N_108,In_423,In_431);
nand U109 (N_109,In_102,In_250);
nand U110 (N_110,In_114,In_307);
nand U111 (N_111,In_396,In_411);
nor U112 (N_112,In_215,In_32);
or U113 (N_113,In_58,In_169);
nand U114 (N_114,In_106,In_481);
and U115 (N_115,In_309,In_65);
or U116 (N_116,In_55,In_101);
and U117 (N_117,In_251,In_474);
nor U118 (N_118,In_208,In_1);
and U119 (N_119,In_274,In_76);
or U120 (N_120,In_173,In_149);
and U121 (N_121,In_36,In_249);
nor U122 (N_122,In_145,In_41);
nor U123 (N_123,In_322,In_178);
nand U124 (N_124,In_246,In_248);
nand U125 (N_125,In_78,In_401);
nor U126 (N_126,In_482,In_67);
or U127 (N_127,In_233,In_459);
or U128 (N_128,In_291,In_61);
nor U129 (N_129,In_373,In_64);
nor U130 (N_130,In_144,In_228);
and U131 (N_131,In_192,In_151);
or U132 (N_132,In_437,In_472);
or U133 (N_133,In_340,In_270);
or U134 (N_134,In_2,In_213);
or U135 (N_135,In_182,In_464);
nand U136 (N_136,In_339,In_418);
nor U137 (N_137,In_372,In_278);
and U138 (N_138,In_491,In_444);
and U139 (N_139,In_7,In_272);
nand U140 (N_140,In_440,In_59);
nor U141 (N_141,In_462,In_370);
nand U142 (N_142,In_330,In_21);
or U143 (N_143,In_299,In_218);
nand U144 (N_144,In_338,In_343);
nand U145 (N_145,In_318,In_331);
or U146 (N_146,In_142,In_447);
nand U147 (N_147,In_400,In_337);
and U148 (N_148,In_342,In_266);
nand U149 (N_149,In_54,In_130);
and U150 (N_150,In_312,In_77);
nand U151 (N_151,In_374,In_267);
or U152 (N_152,In_492,In_15);
and U153 (N_153,In_146,In_168);
or U154 (N_154,In_388,In_242);
and U155 (N_155,In_198,In_424);
nand U156 (N_156,In_490,In_189);
or U157 (N_157,In_287,In_477);
or U158 (N_158,In_120,In_148);
nor U159 (N_159,In_326,In_445);
nor U160 (N_160,In_92,In_310);
nand U161 (N_161,In_304,In_203);
and U162 (N_162,In_314,In_8);
nor U163 (N_163,In_402,In_116);
nor U164 (N_164,In_38,In_398);
and U165 (N_165,In_392,In_256);
and U166 (N_166,In_375,In_97);
or U167 (N_167,In_335,In_220);
nor U168 (N_168,In_448,In_456);
nor U169 (N_169,In_224,In_44);
nor U170 (N_170,In_353,In_387);
nor U171 (N_171,In_239,In_466);
and U172 (N_172,In_281,In_419);
nor U173 (N_173,In_371,In_478);
and U174 (N_174,In_416,In_294);
nand U175 (N_175,In_346,In_170);
nand U176 (N_176,In_494,In_263);
nor U177 (N_177,In_356,In_232);
and U178 (N_178,In_51,In_160);
or U179 (N_179,In_408,In_52);
or U180 (N_180,In_258,In_24);
nand U181 (N_181,In_421,In_129);
nand U182 (N_182,In_262,In_344);
and U183 (N_183,In_358,In_17);
nor U184 (N_184,In_226,In_354);
nor U185 (N_185,In_158,In_57);
nand U186 (N_186,In_469,In_300);
or U187 (N_187,In_280,In_190);
and U188 (N_188,In_350,In_45);
nor U189 (N_189,In_98,In_285);
nor U190 (N_190,In_412,In_399);
or U191 (N_191,In_488,In_33);
and U192 (N_192,In_229,In_404);
and U193 (N_193,In_227,In_379);
nor U194 (N_194,In_157,In_265);
nand U195 (N_195,In_88,In_83);
nand U196 (N_196,In_409,In_117);
and U197 (N_197,In_138,In_323);
and U198 (N_198,In_403,In_325);
nor U199 (N_199,In_284,In_422);
nand U200 (N_200,In_244,In_390);
nand U201 (N_201,In_136,In_163);
or U202 (N_202,In_386,In_167);
and U203 (N_203,In_367,In_321);
nand U204 (N_204,In_329,In_84);
and U205 (N_205,In_305,In_162);
nor U206 (N_206,In_28,In_383);
and U207 (N_207,In_259,In_495);
and U208 (N_208,In_333,In_196);
and U209 (N_209,In_363,In_486);
nand U210 (N_210,In_132,In_164);
nor U211 (N_211,In_207,In_442);
and U212 (N_212,In_306,In_458);
nand U213 (N_213,In_413,In_13);
and U214 (N_214,In_104,In_435);
nor U215 (N_215,In_127,In_25);
nand U216 (N_216,In_436,In_238);
nor U217 (N_217,In_289,In_90);
nor U218 (N_218,In_71,In_223);
nand U219 (N_219,In_6,In_364);
nand U220 (N_220,In_406,In_79);
nand U221 (N_221,In_53,In_154);
nand U222 (N_222,In_324,In_27);
nand U223 (N_223,In_394,In_216);
nand U224 (N_224,In_273,In_405);
nor U225 (N_225,In_427,In_319);
and U226 (N_226,In_391,In_301);
nand U227 (N_227,In_463,In_47);
or U228 (N_228,In_125,In_313);
nor U229 (N_229,In_110,In_175);
or U230 (N_230,In_150,In_376);
nor U231 (N_231,In_395,In_16);
nand U232 (N_232,In_467,In_475);
nand U233 (N_233,In_369,In_352);
and U234 (N_234,In_429,In_457);
or U235 (N_235,In_152,In_211);
nand U236 (N_236,In_380,In_327);
nand U237 (N_237,In_209,In_56);
or U238 (N_238,In_473,In_341);
nor U239 (N_239,In_134,In_5);
nor U240 (N_240,In_122,In_42);
nand U241 (N_241,In_484,In_105);
nand U242 (N_242,In_351,In_107);
nand U243 (N_243,In_366,In_187);
and U244 (N_244,In_433,In_86);
nand U245 (N_245,In_172,In_349);
or U246 (N_246,In_360,In_295);
and U247 (N_247,In_12,In_455);
nand U248 (N_248,In_377,In_22);
nand U249 (N_249,In_119,In_153);
nor U250 (N_250,In_433,In_225);
nand U251 (N_251,In_318,In_309);
nor U252 (N_252,In_86,In_65);
nor U253 (N_253,In_395,In_101);
nor U254 (N_254,In_96,In_147);
or U255 (N_255,In_480,In_86);
nand U256 (N_256,In_0,In_243);
nand U257 (N_257,In_162,In_237);
or U258 (N_258,In_219,In_270);
or U259 (N_259,In_175,In_497);
nand U260 (N_260,In_215,In_327);
nand U261 (N_261,In_52,In_92);
nand U262 (N_262,In_80,In_82);
or U263 (N_263,In_82,In_322);
or U264 (N_264,In_173,In_108);
and U265 (N_265,In_87,In_491);
or U266 (N_266,In_477,In_295);
and U267 (N_267,In_468,In_53);
xor U268 (N_268,In_2,In_307);
nor U269 (N_269,In_399,In_241);
nor U270 (N_270,In_199,In_401);
and U271 (N_271,In_233,In_346);
nand U272 (N_272,In_474,In_365);
or U273 (N_273,In_12,In_424);
and U274 (N_274,In_55,In_306);
or U275 (N_275,In_262,In_308);
and U276 (N_276,In_235,In_342);
nor U277 (N_277,In_66,In_228);
or U278 (N_278,In_222,In_426);
and U279 (N_279,In_311,In_347);
nor U280 (N_280,In_174,In_65);
or U281 (N_281,In_187,In_76);
nand U282 (N_282,In_336,In_46);
or U283 (N_283,In_324,In_200);
xnor U284 (N_284,In_420,In_75);
nor U285 (N_285,In_176,In_364);
or U286 (N_286,In_227,In_47);
and U287 (N_287,In_49,In_166);
or U288 (N_288,In_347,In_294);
nand U289 (N_289,In_491,In_426);
nor U290 (N_290,In_110,In_132);
or U291 (N_291,In_294,In_202);
or U292 (N_292,In_28,In_248);
nor U293 (N_293,In_490,In_52);
nor U294 (N_294,In_477,In_404);
nor U295 (N_295,In_347,In_303);
or U296 (N_296,In_394,In_240);
or U297 (N_297,In_138,In_454);
and U298 (N_298,In_277,In_445);
and U299 (N_299,In_446,In_136);
nor U300 (N_300,In_395,In_109);
nor U301 (N_301,In_300,In_297);
and U302 (N_302,In_378,In_437);
and U303 (N_303,In_250,In_378);
nor U304 (N_304,In_170,In_219);
or U305 (N_305,In_396,In_78);
and U306 (N_306,In_249,In_86);
or U307 (N_307,In_478,In_355);
or U308 (N_308,In_285,In_55);
nand U309 (N_309,In_325,In_405);
and U310 (N_310,In_76,In_111);
or U311 (N_311,In_205,In_438);
nor U312 (N_312,In_128,In_404);
nor U313 (N_313,In_186,In_74);
nand U314 (N_314,In_154,In_379);
nor U315 (N_315,In_204,In_246);
or U316 (N_316,In_112,In_464);
nor U317 (N_317,In_409,In_348);
nor U318 (N_318,In_303,In_287);
nor U319 (N_319,In_455,In_330);
and U320 (N_320,In_130,In_352);
or U321 (N_321,In_360,In_336);
or U322 (N_322,In_191,In_484);
nor U323 (N_323,In_376,In_317);
and U324 (N_324,In_261,In_174);
and U325 (N_325,In_377,In_404);
nor U326 (N_326,In_22,In_446);
nand U327 (N_327,In_305,In_56);
nor U328 (N_328,In_409,In_264);
and U329 (N_329,In_65,In_2);
nor U330 (N_330,In_45,In_139);
and U331 (N_331,In_8,In_278);
and U332 (N_332,In_132,In_392);
nand U333 (N_333,In_174,In_414);
nand U334 (N_334,In_306,In_394);
and U335 (N_335,In_234,In_213);
or U336 (N_336,In_205,In_121);
nor U337 (N_337,In_40,In_452);
or U338 (N_338,In_340,In_295);
nand U339 (N_339,In_26,In_150);
and U340 (N_340,In_318,In_354);
and U341 (N_341,In_112,In_22);
nand U342 (N_342,In_472,In_125);
nand U343 (N_343,In_324,In_125);
and U344 (N_344,In_12,In_414);
or U345 (N_345,In_57,In_41);
nor U346 (N_346,In_309,In_66);
and U347 (N_347,In_125,In_286);
and U348 (N_348,In_106,In_269);
nand U349 (N_349,In_114,In_485);
or U350 (N_350,In_192,In_488);
nor U351 (N_351,In_421,In_9);
nor U352 (N_352,In_445,In_110);
nand U353 (N_353,In_129,In_381);
and U354 (N_354,In_379,In_373);
nand U355 (N_355,In_333,In_16);
nand U356 (N_356,In_486,In_1);
or U357 (N_357,In_470,In_377);
or U358 (N_358,In_123,In_169);
or U359 (N_359,In_469,In_238);
or U360 (N_360,In_364,In_463);
nor U361 (N_361,In_261,In_431);
nand U362 (N_362,In_140,In_243);
nand U363 (N_363,In_324,In_53);
nand U364 (N_364,In_79,In_234);
or U365 (N_365,In_264,In_397);
nand U366 (N_366,In_350,In_292);
or U367 (N_367,In_68,In_85);
or U368 (N_368,In_99,In_199);
or U369 (N_369,In_109,In_12);
nor U370 (N_370,In_294,In_55);
or U371 (N_371,In_172,In_162);
and U372 (N_372,In_81,In_228);
nor U373 (N_373,In_305,In_28);
or U374 (N_374,In_139,In_386);
and U375 (N_375,In_132,In_322);
and U376 (N_376,In_170,In_285);
or U377 (N_377,In_479,In_434);
nand U378 (N_378,In_83,In_391);
and U379 (N_379,In_362,In_22);
nor U380 (N_380,In_450,In_66);
and U381 (N_381,In_408,In_152);
nor U382 (N_382,In_202,In_478);
nor U383 (N_383,In_100,In_300);
or U384 (N_384,In_229,In_89);
or U385 (N_385,In_431,In_312);
nand U386 (N_386,In_152,In_123);
nor U387 (N_387,In_412,In_290);
nor U388 (N_388,In_44,In_328);
nor U389 (N_389,In_487,In_230);
nor U390 (N_390,In_440,In_54);
or U391 (N_391,In_219,In_455);
or U392 (N_392,In_202,In_307);
nand U393 (N_393,In_152,In_247);
nor U394 (N_394,In_90,In_244);
nor U395 (N_395,In_405,In_4);
or U396 (N_396,In_187,In_136);
nand U397 (N_397,In_369,In_173);
nand U398 (N_398,In_492,In_297);
or U399 (N_399,In_248,In_175);
nor U400 (N_400,In_355,In_75);
nand U401 (N_401,In_337,In_362);
nand U402 (N_402,In_486,In_293);
and U403 (N_403,In_433,In_11);
or U404 (N_404,In_36,In_465);
or U405 (N_405,In_41,In_26);
and U406 (N_406,In_365,In_251);
and U407 (N_407,In_215,In_304);
nand U408 (N_408,In_397,In_62);
nor U409 (N_409,In_268,In_451);
nor U410 (N_410,In_464,In_208);
and U411 (N_411,In_95,In_429);
nand U412 (N_412,In_435,In_162);
nand U413 (N_413,In_16,In_38);
nor U414 (N_414,In_311,In_473);
or U415 (N_415,In_73,In_231);
and U416 (N_416,In_47,In_264);
or U417 (N_417,In_313,In_233);
and U418 (N_418,In_448,In_152);
nand U419 (N_419,In_101,In_334);
or U420 (N_420,In_325,In_473);
and U421 (N_421,In_222,In_60);
nand U422 (N_422,In_441,In_476);
and U423 (N_423,In_338,In_220);
or U424 (N_424,In_355,In_2);
nand U425 (N_425,In_379,In_84);
and U426 (N_426,In_412,In_199);
or U427 (N_427,In_445,In_387);
nand U428 (N_428,In_56,In_311);
nand U429 (N_429,In_38,In_45);
nand U430 (N_430,In_137,In_318);
and U431 (N_431,In_1,In_249);
nand U432 (N_432,In_350,In_105);
or U433 (N_433,In_51,In_216);
nor U434 (N_434,In_321,In_1);
nand U435 (N_435,In_438,In_399);
or U436 (N_436,In_55,In_207);
nor U437 (N_437,In_230,In_356);
or U438 (N_438,In_266,In_255);
nor U439 (N_439,In_341,In_302);
nor U440 (N_440,In_62,In_30);
and U441 (N_441,In_462,In_403);
or U442 (N_442,In_316,In_179);
and U443 (N_443,In_316,In_242);
xor U444 (N_444,In_495,In_485);
nor U445 (N_445,In_423,In_348);
and U446 (N_446,In_435,In_406);
nand U447 (N_447,In_200,In_316);
nand U448 (N_448,In_285,In_267);
and U449 (N_449,In_294,In_32);
nor U450 (N_450,In_225,In_406);
nor U451 (N_451,In_211,In_71);
or U452 (N_452,In_183,In_75);
or U453 (N_453,In_435,In_182);
or U454 (N_454,In_411,In_237);
or U455 (N_455,In_144,In_7);
nor U456 (N_456,In_453,In_343);
or U457 (N_457,In_428,In_326);
or U458 (N_458,In_207,In_409);
or U459 (N_459,In_210,In_233);
or U460 (N_460,In_127,In_499);
and U461 (N_461,In_125,In_261);
or U462 (N_462,In_251,In_379);
and U463 (N_463,In_274,In_102);
and U464 (N_464,In_138,In_341);
or U465 (N_465,In_356,In_186);
nand U466 (N_466,In_38,In_407);
and U467 (N_467,In_497,In_165);
nand U468 (N_468,In_163,In_457);
xor U469 (N_469,In_474,In_434);
nor U470 (N_470,In_497,In_19);
nand U471 (N_471,In_288,In_495);
and U472 (N_472,In_202,In_58);
and U473 (N_473,In_413,In_345);
or U474 (N_474,In_205,In_490);
nor U475 (N_475,In_9,In_102);
or U476 (N_476,In_75,In_490);
and U477 (N_477,In_262,In_153);
or U478 (N_478,In_452,In_234);
and U479 (N_479,In_401,In_327);
nor U480 (N_480,In_237,In_222);
or U481 (N_481,In_242,In_62);
nand U482 (N_482,In_62,In_82);
and U483 (N_483,In_418,In_386);
and U484 (N_484,In_31,In_492);
nor U485 (N_485,In_314,In_222);
nand U486 (N_486,In_309,In_0);
nand U487 (N_487,In_335,In_69);
nand U488 (N_488,In_165,In_349);
nand U489 (N_489,In_102,In_476);
and U490 (N_490,In_69,In_419);
nor U491 (N_491,In_220,In_193);
xnor U492 (N_492,In_498,In_433);
or U493 (N_493,In_353,In_194);
and U494 (N_494,In_68,In_473);
or U495 (N_495,In_164,In_363);
or U496 (N_496,In_363,In_448);
nand U497 (N_497,In_56,In_324);
nand U498 (N_498,In_372,In_170);
and U499 (N_499,In_278,In_409);
nand U500 (N_500,In_375,In_452);
or U501 (N_501,In_314,In_109);
or U502 (N_502,In_422,In_447);
and U503 (N_503,In_145,In_315);
or U504 (N_504,In_213,In_128);
and U505 (N_505,In_256,In_309);
nand U506 (N_506,In_142,In_402);
or U507 (N_507,In_45,In_260);
or U508 (N_508,In_482,In_366);
and U509 (N_509,In_424,In_415);
xnor U510 (N_510,In_287,In_37);
nand U511 (N_511,In_109,In_141);
and U512 (N_512,In_12,In_244);
and U513 (N_513,In_389,In_269);
nand U514 (N_514,In_334,In_207);
nor U515 (N_515,In_172,In_20);
nor U516 (N_516,In_42,In_423);
or U517 (N_517,In_353,In_158);
xnor U518 (N_518,In_221,In_397);
and U519 (N_519,In_159,In_149);
nor U520 (N_520,In_204,In_114);
nor U521 (N_521,In_78,In_253);
or U522 (N_522,In_55,In_128);
nand U523 (N_523,In_479,In_350);
nor U524 (N_524,In_164,In_311);
nor U525 (N_525,In_93,In_118);
nor U526 (N_526,In_158,In_274);
and U527 (N_527,In_421,In_22);
nor U528 (N_528,In_486,In_496);
and U529 (N_529,In_234,In_119);
nor U530 (N_530,In_393,In_168);
and U531 (N_531,In_483,In_448);
and U532 (N_532,In_178,In_460);
or U533 (N_533,In_336,In_154);
nand U534 (N_534,In_105,In_353);
and U535 (N_535,In_8,In_169);
nor U536 (N_536,In_193,In_421);
nand U537 (N_537,In_391,In_305);
nand U538 (N_538,In_388,In_188);
and U539 (N_539,In_236,In_459);
nand U540 (N_540,In_491,In_236);
nor U541 (N_541,In_136,In_457);
or U542 (N_542,In_206,In_349);
nor U543 (N_543,In_289,In_248);
nand U544 (N_544,In_78,In_135);
or U545 (N_545,In_131,In_353);
and U546 (N_546,In_121,In_259);
nor U547 (N_547,In_243,In_3);
nand U548 (N_548,In_240,In_342);
nand U549 (N_549,In_123,In_362);
nor U550 (N_550,In_23,In_418);
nand U551 (N_551,In_217,In_15);
or U552 (N_552,In_132,In_131);
nor U553 (N_553,In_33,In_218);
or U554 (N_554,In_329,In_152);
or U555 (N_555,In_81,In_278);
or U556 (N_556,In_407,In_434);
nor U557 (N_557,In_309,In_391);
and U558 (N_558,In_201,In_49);
nand U559 (N_559,In_253,In_324);
nor U560 (N_560,In_417,In_420);
nor U561 (N_561,In_345,In_245);
or U562 (N_562,In_262,In_252);
nor U563 (N_563,In_455,In_132);
nand U564 (N_564,In_120,In_47);
nor U565 (N_565,In_297,In_277);
nand U566 (N_566,In_385,In_309);
and U567 (N_567,In_28,In_58);
nor U568 (N_568,In_82,In_412);
and U569 (N_569,In_93,In_476);
nand U570 (N_570,In_108,In_435);
and U571 (N_571,In_479,In_220);
and U572 (N_572,In_308,In_356);
nor U573 (N_573,In_241,In_337);
nor U574 (N_574,In_116,In_95);
or U575 (N_575,In_104,In_345);
nand U576 (N_576,In_273,In_339);
or U577 (N_577,In_245,In_74);
nand U578 (N_578,In_432,In_401);
nand U579 (N_579,In_266,In_376);
and U580 (N_580,In_151,In_112);
and U581 (N_581,In_16,In_256);
or U582 (N_582,In_31,In_269);
or U583 (N_583,In_76,In_322);
or U584 (N_584,In_368,In_249);
and U585 (N_585,In_389,In_79);
nor U586 (N_586,In_42,In_260);
nand U587 (N_587,In_72,In_16);
nor U588 (N_588,In_231,In_379);
nand U589 (N_589,In_132,In_220);
nand U590 (N_590,In_417,In_480);
and U591 (N_591,In_201,In_453);
or U592 (N_592,In_284,In_40);
nand U593 (N_593,In_293,In_170);
or U594 (N_594,In_123,In_322);
or U595 (N_595,In_174,In_365);
nand U596 (N_596,In_261,In_423);
nand U597 (N_597,In_404,In_46);
nor U598 (N_598,In_278,In_379);
or U599 (N_599,In_43,In_96);
or U600 (N_600,N_436,N_342);
nor U601 (N_601,N_419,N_9);
and U602 (N_602,N_253,N_180);
or U603 (N_603,N_562,N_329);
nor U604 (N_604,N_501,N_414);
and U605 (N_605,N_413,N_529);
nand U606 (N_606,N_429,N_24);
nor U607 (N_607,N_498,N_406);
xor U608 (N_608,N_264,N_170);
nor U609 (N_609,N_62,N_547);
or U610 (N_610,N_208,N_460);
nor U611 (N_611,N_12,N_548);
nand U612 (N_612,N_257,N_488);
and U613 (N_613,N_124,N_151);
nand U614 (N_614,N_318,N_55);
xnor U615 (N_615,N_68,N_287);
or U616 (N_616,N_493,N_274);
nand U617 (N_617,N_63,N_566);
nand U618 (N_618,N_204,N_374);
nor U619 (N_619,N_381,N_120);
and U620 (N_620,N_317,N_80);
and U621 (N_621,N_357,N_355);
nand U622 (N_622,N_17,N_399);
nand U623 (N_623,N_393,N_74);
and U624 (N_624,N_153,N_331);
nand U625 (N_625,N_451,N_137);
or U626 (N_626,N_30,N_244);
and U627 (N_627,N_16,N_134);
nand U628 (N_628,N_513,N_554);
and U629 (N_629,N_28,N_416);
and U630 (N_630,N_135,N_76);
or U631 (N_631,N_471,N_371);
or U632 (N_632,N_226,N_360);
and U633 (N_633,N_2,N_586);
nor U634 (N_634,N_64,N_350);
and U635 (N_635,N_510,N_567);
or U636 (N_636,N_33,N_127);
nor U637 (N_637,N_237,N_370);
nor U638 (N_638,N_428,N_211);
or U639 (N_639,N_277,N_125);
nor U640 (N_640,N_197,N_387);
nand U641 (N_641,N_71,N_402);
and U642 (N_642,N_221,N_549);
nor U643 (N_643,N_40,N_546);
or U644 (N_644,N_243,N_66);
or U645 (N_645,N_553,N_580);
and U646 (N_646,N_223,N_213);
nand U647 (N_647,N_344,N_299);
nor U648 (N_648,N_111,N_190);
and U649 (N_649,N_316,N_266);
or U650 (N_650,N_236,N_434);
or U651 (N_651,N_288,N_570);
nand U652 (N_652,N_397,N_443);
or U653 (N_653,N_311,N_385);
nand U654 (N_654,N_322,N_272);
or U655 (N_655,N_14,N_439);
xor U656 (N_656,N_340,N_198);
nor U657 (N_657,N_54,N_352);
or U658 (N_658,N_537,N_115);
or U659 (N_659,N_533,N_247);
nor U660 (N_660,N_392,N_260);
nand U661 (N_661,N_194,N_530);
or U662 (N_662,N_305,N_19);
nor U663 (N_663,N_467,N_187);
nand U664 (N_664,N_246,N_379);
or U665 (N_665,N_309,N_522);
or U666 (N_666,N_104,N_384);
and U667 (N_667,N_368,N_256);
and U668 (N_668,N_388,N_312);
nand U669 (N_669,N_118,N_278);
or U670 (N_670,N_26,N_596);
nand U671 (N_671,N_251,N_425);
nand U672 (N_672,N_473,N_22);
nor U673 (N_673,N_382,N_32);
or U674 (N_674,N_486,N_235);
and U675 (N_675,N_84,N_349);
and U676 (N_676,N_590,N_283);
and U677 (N_677,N_248,N_446);
nor U678 (N_678,N_81,N_10);
or U679 (N_679,N_395,N_75);
nor U680 (N_680,N_107,N_521);
nand U681 (N_681,N_82,N_39);
nand U682 (N_682,N_571,N_8);
nand U683 (N_683,N_441,N_5);
nand U684 (N_684,N_177,N_293);
nor U685 (N_685,N_575,N_377);
nand U686 (N_686,N_527,N_52);
and U687 (N_687,N_503,N_430);
nand U688 (N_688,N_363,N_262);
and U689 (N_689,N_336,N_528);
nor U690 (N_690,N_232,N_573);
nand U691 (N_691,N_523,N_65);
nor U692 (N_692,N_176,N_324);
nor U693 (N_693,N_435,N_507);
and U694 (N_694,N_505,N_119);
or U695 (N_695,N_43,N_483);
or U696 (N_696,N_106,N_588);
nor U697 (N_697,N_462,N_415);
and U698 (N_698,N_544,N_512);
nor U699 (N_699,N_178,N_156);
nor U700 (N_700,N_200,N_576);
or U701 (N_701,N_550,N_275);
and U702 (N_702,N_18,N_240);
nor U703 (N_703,N_144,N_188);
nor U704 (N_704,N_96,N_300);
and U705 (N_705,N_270,N_207);
nand U706 (N_706,N_389,N_356);
nand U707 (N_707,N_372,N_79);
or U708 (N_708,N_591,N_339);
and U709 (N_709,N_87,N_564);
nor U710 (N_710,N_585,N_476);
or U711 (N_711,N_38,N_481);
nor U712 (N_712,N_23,N_140);
and U713 (N_713,N_408,N_319);
nor U714 (N_714,N_122,N_132);
and U715 (N_715,N_390,N_252);
nand U716 (N_716,N_296,N_0);
and U717 (N_717,N_404,N_323);
nand U718 (N_718,N_193,N_411);
or U719 (N_719,N_220,N_268);
nand U720 (N_720,N_407,N_485);
and U721 (N_721,N_496,N_574);
and U722 (N_722,N_378,N_472);
and U723 (N_723,N_44,N_139);
nand U724 (N_724,N_540,N_103);
nor U725 (N_725,N_165,N_263);
nor U726 (N_726,N_155,N_47);
nand U727 (N_727,N_508,N_149);
or U728 (N_728,N_346,N_138);
nand U729 (N_729,N_45,N_94);
xor U730 (N_730,N_233,N_3);
or U731 (N_731,N_347,N_449);
nor U732 (N_732,N_444,N_37);
and U733 (N_733,N_225,N_11);
and U734 (N_734,N_215,N_185);
or U735 (N_735,N_560,N_558);
nand U736 (N_736,N_228,N_326);
nor U737 (N_737,N_181,N_465);
nor U738 (N_738,N_280,N_520);
or U739 (N_739,N_427,N_433);
and U740 (N_740,N_209,N_453);
nand U741 (N_741,N_499,N_83);
and U742 (N_742,N_231,N_468);
nand U743 (N_743,N_517,N_142);
and U744 (N_744,N_121,N_217);
or U745 (N_745,N_196,N_95);
and U746 (N_746,N_51,N_391);
or U747 (N_747,N_568,N_164);
nand U748 (N_748,N_146,N_29);
nor U749 (N_749,N_302,N_531);
and U750 (N_750,N_375,N_285);
nor U751 (N_751,N_269,N_361);
nand U752 (N_752,N_304,N_182);
nor U753 (N_753,N_61,N_48);
nor U754 (N_754,N_158,N_310);
nand U755 (N_755,N_369,N_561);
nor U756 (N_756,N_380,N_131);
nand U757 (N_757,N_201,N_186);
nand U758 (N_758,N_458,N_545);
nand U759 (N_759,N_241,N_482);
nor U760 (N_760,N_337,N_86);
or U761 (N_761,N_437,N_136);
nand U762 (N_762,N_234,N_25);
nand U763 (N_763,N_58,N_455);
nor U764 (N_764,N_452,N_290);
or U765 (N_765,N_117,N_294);
and U766 (N_766,N_261,N_218);
or U767 (N_767,N_516,N_480);
nor U768 (N_768,N_298,N_525);
nand U769 (N_769,N_592,N_184);
nor U770 (N_770,N_597,N_163);
or U771 (N_771,N_333,N_418);
or U772 (N_772,N_1,N_69);
nor U773 (N_773,N_157,N_175);
nand U774 (N_774,N_598,N_569);
and U775 (N_775,N_143,N_367);
nand U776 (N_776,N_89,N_490);
and U777 (N_777,N_171,N_365);
nor U778 (N_778,N_551,N_500);
nor U779 (N_779,N_239,N_470);
nor U780 (N_780,N_572,N_72);
nor U781 (N_781,N_191,N_448);
nand U782 (N_782,N_109,N_295);
nor U783 (N_783,N_478,N_174);
and U784 (N_784,N_447,N_396);
or U785 (N_785,N_254,N_281);
and U786 (N_786,N_212,N_42);
or U787 (N_787,N_276,N_487);
nor U788 (N_788,N_210,N_330);
or U789 (N_789,N_412,N_250);
nand U790 (N_790,N_35,N_366);
or U791 (N_791,N_21,N_474);
or U792 (N_792,N_199,N_582);
or U793 (N_793,N_179,N_489);
and U794 (N_794,N_594,N_341);
and U795 (N_795,N_327,N_362);
nand U796 (N_796,N_282,N_354);
nand U797 (N_797,N_168,N_314);
nor U798 (N_798,N_67,N_494);
or U799 (N_799,N_373,N_114);
nand U800 (N_800,N_129,N_315);
or U801 (N_801,N_543,N_166);
and U802 (N_802,N_90,N_41);
or U803 (N_803,N_581,N_53);
nand U804 (N_804,N_353,N_587);
and U805 (N_805,N_279,N_159);
or U806 (N_806,N_148,N_538);
nand U807 (N_807,N_405,N_245);
or U808 (N_808,N_93,N_286);
nor U809 (N_809,N_161,N_559);
and U810 (N_810,N_464,N_578);
or U811 (N_811,N_255,N_113);
and U812 (N_812,N_227,N_292);
nand U813 (N_813,N_101,N_518);
nor U814 (N_814,N_536,N_141);
or U815 (N_815,N_459,N_92);
nor U816 (N_816,N_15,N_535);
nor U817 (N_817,N_289,N_440);
nand U818 (N_818,N_31,N_565);
nor U819 (N_819,N_504,N_555);
and U820 (N_820,N_541,N_152);
nand U821 (N_821,N_422,N_308);
nand U822 (N_822,N_50,N_20);
and U823 (N_823,N_205,N_307);
and U824 (N_824,N_526,N_303);
and U825 (N_825,N_57,N_130);
or U826 (N_826,N_206,N_258);
and U827 (N_827,N_154,N_259);
or U828 (N_828,N_334,N_173);
nand U829 (N_829,N_423,N_162);
nand U830 (N_830,N_400,N_583);
or U831 (N_831,N_328,N_306);
and U832 (N_832,N_438,N_599);
nor U833 (N_833,N_338,N_249);
nand U834 (N_834,N_99,N_313);
or U835 (N_835,N_105,N_497);
and U836 (N_836,N_359,N_123);
nand U837 (N_837,N_203,N_450);
nor U838 (N_838,N_557,N_454);
nor U839 (N_839,N_579,N_466);
nor U840 (N_840,N_189,N_475);
nor U841 (N_841,N_301,N_383);
or U842 (N_842,N_514,N_70);
nand U843 (N_843,N_60,N_358);
nand U844 (N_844,N_195,N_49);
or U845 (N_845,N_126,N_167);
or U846 (N_846,N_59,N_445);
nand U847 (N_847,N_267,N_577);
nor U848 (N_848,N_364,N_348);
nand U849 (N_849,N_202,N_116);
and U850 (N_850,N_78,N_511);
nor U851 (N_851,N_563,N_556);
nor U852 (N_852,N_265,N_584);
nand U853 (N_853,N_401,N_133);
or U854 (N_854,N_56,N_424);
or U855 (N_855,N_542,N_36);
nand U856 (N_856,N_442,N_102);
nand U857 (N_857,N_456,N_420);
and U858 (N_858,N_160,N_110);
and U859 (N_859,N_230,N_595);
and U860 (N_860,N_183,N_552);
nand U861 (N_861,N_457,N_351);
nor U862 (N_862,N_491,N_219);
and U863 (N_863,N_495,N_417);
nand U864 (N_864,N_432,N_284);
nor U865 (N_865,N_273,N_145);
nand U866 (N_866,N_150,N_539);
or U867 (N_867,N_73,N_325);
or U868 (N_868,N_484,N_222);
nand U869 (N_869,N_98,N_403);
and U870 (N_870,N_410,N_593);
nor U871 (N_871,N_534,N_27);
and U872 (N_872,N_398,N_477);
nand U873 (N_873,N_6,N_409);
nand U874 (N_874,N_4,N_519);
nand U875 (N_875,N_214,N_46);
or U876 (N_876,N_297,N_112);
nand U877 (N_877,N_502,N_506);
or U878 (N_878,N_291,N_376);
nand U879 (N_879,N_431,N_461);
nor U880 (N_880,N_321,N_229);
and U881 (N_881,N_386,N_509);
and U882 (N_882,N_13,N_394);
and U883 (N_883,N_172,N_426);
and U884 (N_884,N_343,N_100);
nor U885 (N_885,N_97,N_332);
nand U886 (N_886,N_169,N_238);
nor U887 (N_887,N_77,N_108);
nor U888 (N_888,N_88,N_463);
and U889 (N_889,N_147,N_216);
nand U890 (N_890,N_515,N_532);
nor U891 (N_891,N_224,N_320);
and U892 (N_892,N_524,N_421);
and U893 (N_893,N_242,N_192);
nand U894 (N_894,N_589,N_128);
and U895 (N_895,N_271,N_7);
and U896 (N_896,N_469,N_335);
nor U897 (N_897,N_85,N_492);
nor U898 (N_898,N_34,N_479);
or U899 (N_899,N_91,N_345);
nand U900 (N_900,N_368,N_366);
and U901 (N_901,N_54,N_304);
nor U902 (N_902,N_165,N_316);
or U903 (N_903,N_226,N_212);
nor U904 (N_904,N_582,N_226);
nand U905 (N_905,N_387,N_368);
or U906 (N_906,N_305,N_522);
and U907 (N_907,N_537,N_201);
nand U908 (N_908,N_262,N_171);
and U909 (N_909,N_202,N_281);
or U910 (N_910,N_224,N_201);
and U911 (N_911,N_64,N_37);
nor U912 (N_912,N_590,N_216);
and U913 (N_913,N_345,N_527);
or U914 (N_914,N_357,N_303);
and U915 (N_915,N_12,N_556);
nor U916 (N_916,N_551,N_284);
nor U917 (N_917,N_139,N_230);
nand U918 (N_918,N_115,N_330);
or U919 (N_919,N_322,N_307);
or U920 (N_920,N_432,N_531);
nor U921 (N_921,N_489,N_38);
or U922 (N_922,N_514,N_510);
nand U923 (N_923,N_431,N_464);
nand U924 (N_924,N_322,N_86);
nor U925 (N_925,N_453,N_119);
and U926 (N_926,N_403,N_563);
and U927 (N_927,N_569,N_322);
nor U928 (N_928,N_224,N_435);
and U929 (N_929,N_267,N_441);
nand U930 (N_930,N_11,N_36);
nand U931 (N_931,N_544,N_408);
and U932 (N_932,N_495,N_227);
or U933 (N_933,N_42,N_454);
nand U934 (N_934,N_213,N_459);
nand U935 (N_935,N_511,N_243);
nand U936 (N_936,N_538,N_206);
xnor U937 (N_937,N_561,N_297);
and U938 (N_938,N_221,N_72);
and U939 (N_939,N_110,N_257);
or U940 (N_940,N_526,N_358);
or U941 (N_941,N_2,N_216);
nor U942 (N_942,N_97,N_305);
or U943 (N_943,N_24,N_7);
and U944 (N_944,N_311,N_153);
and U945 (N_945,N_485,N_189);
or U946 (N_946,N_418,N_317);
nand U947 (N_947,N_526,N_310);
or U948 (N_948,N_481,N_229);
and U949 (N_949,N_164,N_371);
nand U950 (N_950,N_81,N_317);
or U951 (N_951,N_234,N_20);
nor U952 (N_952,N_33,N_296);
or U953 (N_953,N_565,N_116);
nand U954 (N_954,N_545,N_32);
nand U955 (N_955,N_89,N_421);
and U956 (N_956,N_335,N_284);
or U957 (N_957,N_219,N_265);
or U958 (N_958,N_206,N_191);
and U959 (N_959,N_257,N_203);
nor U960 (N_960,N_311,N_464);
and U961 (N_961,N_93,N_189);
and U962 (N_962,N_28,N_305);
nor U963 (N_963,N_339,N_483);
nor U964 (N_964,N_71,N_316);
and U965 (N_965,N_94,N_464);
nor U966 (N_966,N_511,N_429);
or U967 (N_967,N_303,N_519);
nand U968 (N_968,N_423,N_196);
nand U969 (N_969,N_438,N_538);
or U970 (N_970,N_537,N_295);
nor U971 (N_971,N_34,N_372);
nand U972 (N_972,N_107,N_262);
nand U973 (N_973,N_574,N_437);
nor U974 (N_974,N_464,N_228);
or U975 (N_975,N_273,N_376);
xor U976 (N_976,N_131,N_544);
and U977 (N_977,N_30,N_529);
or U978 (N_978,N_138,N_421);
or U979 (N_979,N_439,N_72);
and U980 (N_980,N_569,N_445);
and U981 (N_981,N_413,N_528);
nor U982 (N_982,N_431,N_69);
or U983 (N_983,N_322,N_381);
or U984 (N_984,N_185,N_392);
or U985 (N_985,N_329,N_381);
nor U986 (N_986,N_97,N_160);
xnor U987 (N_987,N_14,N_234);
nand U988 (N_988,N_160,N_245);
or U989 (N_989,N_464,N_424);
nor U990 (N_990,N_268,N_205);
or U991 (N_991,N_274,N_445);
nand U992 (N_992,N_551,N_315);
nand U993 (N_993,N_571,N_249);
nand U994 (N_994,N_478,N_239);
xor U995 (N_995,N_329,N_207);
and U996 (N_996,N_383,N_63);
nand U997 (N_997,N_490,N_323);
nand U998 (N_998,N_476,N_318);
and U999 (N_999,N_11,N_91);
nand U1000 (N_1000,N_514,N_84);
and U1001 (N_1001,N_197,N_469);
nand U1002 (N_1002,N_339,N_340);
and U1003 (N_1003,N_25,N_204);
nand U1004 (N_1004,N_289,N_85);
nor U1005 (N_1005,N_110,N_130);
and U1006 (N_1006,N_412,N_498);
nand U1007 (N_1007,N_559,N_61);
or U1008 (N_1008,N_388,N_533);
nor U1009 (N_1009,N_503,N_31);
and U1010 (N_1010,N_571,N_388);
or U1011 (N_1011,N_251,N_420);
xnor U1012 (N_1012,N_263,N_496);
nand U1013 (N_1013,N_273,N_32);
and U1014 (N_1014,N_231,N_54);
nor U1015 (N_1015,N_193,N_524);
nor U1016 (N_1016,N_527,N_176);
and U1017 (N_1017,N_384,N_242);
and U1018 (N_1018,N_306,N_596);
and U1019 (N_1019,N_595,N_142);
or U1020 (N_1020,N_494,N_318);
nand U1021 (N_1021,N_237,N_401);
or U1022 (N_1022,N_211,N_124);
and U1023 (N_1023,N_148,N_95);
and U1024 (N_1024,N_567,N_241);
nor U1025 (N_1025,N_185,N_240);
or U1026 (N_1026,N_545,N_134);
or U1027 (N_1027,N_29,N_98);
nor U1028 (N_1028,N_71,N_480);
nand U1029 (N_1029,N_431,N_59);
nor U1030 (N_1030,N_157,N_547);
nand U1031 (N_1031,N_445,N_465);
or U1032 (N_1032,N_104,N_75);
or U1033 (N_1033,N_459,N_35);
nor U1034 (N_1034,N_357,N_37);
and U1035 (N_1035,N_480,N_554);
and U1036 (N_1036,N_377,N_583);
and U1037 (N_1037,N_407,N_497);
or U1038 (N_1038,N_42,N_441);
nor U1039 (N_1039,N_11,N_408);
nand U1040 (N_1040,N_228,N_412);
nand U1041 (N_1041,N_197,N_424);
and U1042 (N_1042,N_47,N_254);
nor U1043 (N_1043,N_473,N_398);
nor U1044 (N_1044,N_450,N_95);
or U1045 (N_1045,N_43,N_120);
nor U1046 (N_1046,N_323,N_313);
and U1047 (N_1047,N_101,N_243);
or U1048 (N_1048,N_172,N_9);
and U1049 (N_1049,N_22,N_453);
nor U1050 (N_1050,N_592,N_580);
nor U1051 (N_1051,N_303,N_256);
nand U1052 (N_1052,N_210,N_90);
nand U1053 (N_1053,N_350,N_212);
nand U1054 (N_1054,N_129,N_237);
and U1055 (N_1055,N_559,N_27);
or U1056 (N_1056,N_143,N_407);
or U1057 (N_1057,N_596,N_380);
nor U1058 (N_1058,N_279,N_503);
nand U1059 (N_1059,N_343,N_326);
xor U1060 (N_1060,N_597,N_272);
nand U1061 (N_1061,N_266,N_322);
and U1062 (N_1062,N_213,N_375);
and U1063 (N_1063,N_260,N_445);
nor U1064 (N_1064,N_413,N_79);
nor U1065 (N_1065,N_186,N_557);
nor U1066 (N_1066,N_77,N_575);
or U1067 (N_1067,N_366,N_456);
nor U1068 (N_1068,N_103,N_194);
nand U1069 (N_1069,N_256,N_75);
or U1070 (N_1070,N_353,N_39);
and U1071 (N_1071,N_95,N_164);
or U1072 (N_1072,N_470,N_586);
nand U1073 (N_1073,N_481,N_292);
nor U1074 (N_1074,N_541,N_553);
nor U1075 (N_1075,N_541,N_378);
nor U1076 (N_1076,N_22,N_326);
and U1077 (N_1077,N_330,N_572);
or U1078 (N_1078,N_315,N_148);
and U1079 (N_1079,N_275,N_549);
and U1080 (N_1080,N_551,N_380);
or U1081 (N_1081,N_429,N_349);
nor U1082 (N_1082,N_573,N_90);
nand U1083 (N_1083,N_196,N_145);
and U1084 (N_1084,N_371,N_301);
nand U1085 (N_1085,N_537,N_495);
nand U1086 (N_1086,N_544,N_465);
or U1087 (N_1087,N_126,N_284);
nor U1088 (N_1088,N_545,N_228);
and U1089 (N_1089,N_345,N_88);
nand U1090 (N_1090,N_389,N_207);
nor U1091 (N_1091,N_165,N_315);
nand U1092 (N_1092,N_299,N_10);
nor U1093 (N_1093,N_105,N_220);
nor U1094 (N_1094,N_425,N_484);
and U1095 (N_1095,N_218,N_499);
and U1096 (N_1096,N_192,N_477);
nor U1097 (N_1097,N_51,N_530);
and U1098 (N_1098,N_297,N_430);
nand U1099 (N_1099,N_445,N_188);
nor U1100 (N_1100,N_351,N_577);
and U1101 (N_1101,N_175,N_0);
nand U1102 (N_1102,N_566,N_517);
and U1103 (N_1103,N_118,N_299);
and U1104 (N_1104,N_33,N_423);
nor U1105 (N_1105,N_311,N_250);
or U1106 (N_1106,N_156,N_448);
nor U1107 (N_1107,N_453,N_598);
nor U1108 (N_1108,N_403,N_82);
nor U1109 (N_1109,N_516,N_94);
or U1110 (N_1110,N_171,N_134);
and U1111 (N_1111,N_56,N_226);
nand U1112 (N_1112,N_103,N_365);
nor U1113 (N_1113,N_3,N_121);
and U1114 (N_1114,N_171,N_67);
nand U1115 (N_1115,N_540,N_349);
nand U1116 (N_1116,N_336,N_511);
nand U1117 (N_1117,N_260,N_353);
nor U1118 (N_1118,N_365,N_81);
or U1119 (N_1119,N_229,N_42);
or U1120 (N_1120,N_588,N_442);
nand U1121 (N_1121,N_89,N_195);
or U1122 (N_1122,N_332,N_352);
or U1123 (N_1123,N_177,N_136);
nor U1124 (N_1124,N_352,N_365);
nand U1125 (N_1125,N_221,N_60);
and U1126 (N_1126,N_591,N_418);
or U1127 (N_1127,N_267,N_283);
and U1128 (N_1128,N_42,N_532);
nor U1129 (N_1129,N_210,N_427);
and U1130 (N_1130,N_66,N_0);
nand U1131 (N_1131,N_93,N_296);
and U1132 (N_1132,N_78,N_532);
or U1133 (N_1133,N_568,N_566);
and U1134 (N_1134,N_584,N_293);
nor U1135 (N_1135,N_578,N_576);
xnor U1136 (N_1136,N_31,N_392);
nand U1137 (N_1137,N_443,N_312);
nor U1138 (N_1138,N_429,N_353);
nor U1139 (N_1139,N_502,N_521);
nand U1140 (N_1140,N_132,N_69);
nor U1141 (N_1141,N_474,N_372);
nand U1142 (N_1142,N_139,N_509);
or U1143 (N_1143,N_351,N_78);
nand U1144 (N_1144,N_503,N_254);
and U1145 (N_1145,N_12,N_404);
or U1146 (N_1146,N_301,N_112);
nand U1147 (N_1147,N_94,N_126);
nand U1148 (N_1148,N_570,N_497);
or U1149 (N_1149,N_566,N_96);
nand U1150 (N_1150,N_571,N_309);
nand U1151 (N_1151,N_532,N_349);
nor U1152 (N_1152,N_467,N_70);
and U1153 (N_1153,N_324,N_318);
nor U1154 (N_1154,N_558,N_315);
nor U1155 (N_1155,N_183,N_34);
and U1156 (N_1156,N_478,N_519);
or U1157 (N_1157,N_68,N_572);
or U1158 (N_1158,N_496,N_532);
nor U1159 (N_1159,N_448,N_385);
nand U1160 (N_1160,N_188,N_593);
and U1161 (N_1161,N_94,N_386);
nand U1162 (N_1162,N_394,N_277);
nand U1163 (N_1163,N_440,N_290);
or U1164 (N_1164,N_395,N_447);
nor U1165 (N_1165,N_123,N_171);
nor U1166 (N_1166,N_303,N_297);
nor U1167 (N_1167,N_85,N_436);
and U1168 (N_1168,N_0,N_196);
and U1169 (N_1169,N_576,N_523);
nand U1170 (N_1170,N_466,N_469);
or U1171 (N_1171,N_533,N_417);
or U1172 (N_1172,N_204,N_464);
and U1173 (N_1173,N_590,N_548);
and U1174 (N_1174,N_111,N_82);
nor U1175 (N_1175,N_496,N_106);
nand U1176 (N_1176,N_68,N_258);
or U1177 (N_1177,N_140,N_235);
and U1178 (N_1178,N_374,N_102);
nand U1179 (N_1179,N_412,N_381);
and U1180 (N_1180,N_463,N_193);
or U1181 (N_1181,N_312,N_13);
nand U1182 (N_1182,N_276,N_251);
or U1183 (N_1183,N_3,N_383);
or U1184 (N_1184,N_576,N_106);
nor U1185 (N_1185,N_352,N_244);
and U1186 (N_1186,N_385,N_400);
nor U1187 (N_1187,N_293,N_295);
nand U1188 (N_1188,N_559,N_251);
or U1189 (N_1189,N_364,N_178);
nor U1190 (N_1190,N_281,N_390);
or U1191 (N_1191,N_71,N_529);
nor U1192 (N_1192,N_151,N_474);
nand U1193 (N_1193,N_397,N_579);
and U1194 (N_1194,N_101,N_485);
nand U1195 (N_1195,N_460,N_272);
nor U1196 (N_1196,N_44,N_449);
or U1197 (N_1197,N_7,N_500);
and U1198 (N_1198,N_452,N_480);
nand U1199 (N_1199,N_21,N_55);
nand U1200 (N_1200,N_712,N_830);
or U1201 (N_1201,N_984,N_1133);
or U1202 (N_1202,N_1113,N_1063);
or U1203 (N_1203,N_722,N_901);
nor U1204 (N_1204,N_1110,N_1155);
or U1205 (N_1205,N_1070,N_1045);
or U1206 (N_1206,N_1187,N_640);
and U1207 (N_1207,N_1067,N_920);
nand U1208 (N_1208,N_1088,N_1198);
and U1209 (N_1209,N_738,N_868);
and U1210 (N_1210,N_903,N_1081);
nor U1211 (N_1211,N_1091,N_894);
or U1212 (N_1212,N_658,N_662);
or U1213 (N_1213,N_758,N_888);
or U1214 (N_1214,N_1086,N_697);
or U1215 (N_1215,N_1159,N_1185);
nor U1216 (N_1216,N_1118,N_1020);
nand U1217 (N_1217,N_977,N_849);
xor U1218 (N_1218,N_689,N_1094);
nor U1219 (N_1219,N_1038,N_938);
and U1220 (N_1220,N_703,N_879);
or U1221 (N_1221,N_989,N_843);
nor U1222 (N_1222,N_800,N_1097);
nand U1223 (N_1223,N_926,N_605);
or U1224 (N_1224,N_1033,N_713);
nand U1225 (N_1225,N_826,N_1017);
nor U1226 (N_1226,N_1010,N_1095);
or U1227 (N_1227,N_1047,N_931);
nand U1228 (N_1228,N_771,N_1034);
nor U1229 (N_1229,N_996,N_1079);
nand U1230 (N_1230,N_660,N_808);
nor U1231 (N_1231,N_1180,N_925);
and U1232 (N_1232,N_1169,N_1144);
or U1233 (N_1233,N_795,N_1011);
nor U1234 (N_1234,N_778,N_786);
and U1235 (N_1235,N_1040,N_856);
nor U1236 (N_1236,N_957,N_1152);
or U1237 (N_1237,N_917,N_902);
or U1238 (N_1238,N_864,N_1083);
nand U1239 (N_1239,N_971,N_763);
or U1240 (N_1240,N_740,N_1009);
and U1241 (N_1241,N_846,N_878);
and U1242 (N_1242,N_1082,N_742);
and U1243 (N_1243,N_764,N_937);
nor U1244 (N_1244,N_645,N_743);
and U1245 (N_1245,N_986,N_1078);
and U1246 (N_1246,N_1109,N_1071);
or U1247 (N_1247,N_757,N_622);
nor U1248 (N_1248,N_992,N_892);
and U1249 (N_1249,N_1195,N_867);
or U1250 (N_1250,N_1062,N_760);
nor U1251 (N_1251,N_885,N_784);
and U1252 (N_1252,N_747,N_814);
xnor U1253 (N_1253,N_1131,N_1019);
nor U1254 (N_1254,N_644,N_1149);
nor U1255 (N_1255,N_792,N_750);
nor U1256 (N_1256,N_891,N_1182);
nand U1257 (N_1257,N_987,N_872);
nand U1258 (N_1258,N_816,N_1106);
nand U1259 (N_1259,N_839,N_613);
nor U1260 (N_1260,N_635,N_781);
or U1261 (N_1261,N_1005,N_1143);
and U1262 (N_1262,N_705,N_833);
nand U1263 (N_1263,N_769,N_1012);
and U1264 (N_1264,N_995,N_844);
and U1265 (N_1265,N_620,N_639);
nor U1266 (N_1266,N_935,N_1018);
nor U1267 (N_1267,N_845,N_788);
nor U1268 (N_1268,N_1055,N_944);
or U1269 (N_1269,N_921,N_875);
nand U1270 (N_1270,N_663,N_779);
nor U1271 (N_1271,N_1048,N_1080);
and U1272 (N_1272,N_1073,N_690);
nor U1273 (N_1273,N_765,N_924);
and U1274 (N_1274,N_665,N_678);
nand U1275 (N_1275,N_1192,N_909);
nor U1276 (N_1276,N_600,N_632);
or U1277 (N_1277,N_945,N_670);
nand U1278 (N_1278,N_1154,N_941);
or U1279 (N_1279,N_828,N_1189);
nor U1280 (N_1280,N_1117,N_1087);
and U1281 (N_1281,N_772,N_676);
and U1282 (N_1282,N_708,N_677);
nand U1283 (N_1283,N_861,N_842);
and U1284 (N_1284,N_966,N_1116);
or U1285 (N_1285,N_1075,N_1130);
or U1286 (N_1286,N_756,N_1061);
nand U1287 (N_1287,N_895,N_1049);
or U1288 (N_1288,N_853,N_1026);
nand U1289 (N_1289,N_854,N_1015);
or U1290 (N_1290,N_1132,N_954);
and U1291 (N_1291,N_739,N_978);
nand U1292 (N_1292,N_647,N_923);
nor U1293 (N_1293,N_1181,N_634);
or U1294 (N_1294,N_907,N_964);
nor U1295 (N_1295,N_871,N_865);
and U1296 (N_1296,N_649,N_696);
nand U1297 (N_1297,N_729,N_919);
or U1298 (N_1298,N_818,N_751);
and U1299 (N_1299,N_711,N_719);
nor U1300 (N_1300,N_768,N_942);
nor U1301 (N_1301,N_1129,N_684);
nor U1302 (N_1302,N_1092,N_1065);
or U1303 (N_1303,N_1003,N_787);
nor U1304 (N_1304,N_619,N_824);
and U1305 (N_1305,N_1165,N_603);
and U1306 (N_1306,N_1194,N_1004);
nand U1307 (N_1307,N_1183,N_1103);
nand U1308 (N_1308,N_852,N_1108);
or U1309 (N_1309,N_922,N_961);
nor U1310 (N_1310,N_982,N_1058);
nand U1311 (N_1311,N_1046,N_911);
and U1312 (N_1312,N_749,N_1059);
or U1313 (N_1313,N_654,N_767);
nor U1314 (N_1314,N_1127,N_761);
and U1315 (N_1315,N_1199,N_1153);
nand U1316 (N_1316,N_621,N_821);
or U1317 (N_1317,N_806,N_1123);
nand U1318 (N_1318,N_766,N_835);
nand U1319 (N_1319,N_686,N_1030);
nor U1320 (N_1320,N_914,N_896);
nor U1321 (N_1321,N_720,N_812);
or U1322 (N_1322,N_1021,N_1147);
nand U1323 (N_1323,N_688,N_789);
or U1324 (N_1324,N_681,N_623);
or U1325 (N_1325,N_626,N_685);
nand U1326 (N_1326,N_753,N_1124);
nor U1327 (N_1327,N_981,N_904);
and U1328 (N_1328,N_1054,N_841);
nand U1329 (N_1329,N_933,N_1188);
nor U1330 (N_1330,N_886,N_735);
nor U1331 (N_1331,N_797,N_837);
nor U1332 (N_1332,N_775,N_1115);
or U1333 (N_1333,N_625,N_616);
or U1334 (N_1334,N_609,N_918);
nand U1335 (N_1335,N_683,N_1037);
or U1336 (N_1336,N_707,N_962);
nand U1337 (N_1337,N_1024,N_1085);
nand U1338 (N_1338,N_618,N_1043);
and U1339 (N_1339,N_906,N_1051);
nand U1340 (N_1340,N_1077,N_850);
nor U1341 (N_1341,N_1042,N_956);
or U1342 (N_1342,N_699,N_770);
nand U1343 (N_1343,N_637,N_866);
nand U1344 (N_1344,N_791,N_659);
nor U1345 (N_1345,N_927,N_940);
nor U1346 (N_1346,N_1028,N_668);
nor U1347 (N_1347,N_946,N_951);
or U1348 (N_1348,N_710,N_724);
nand U1349 (N_1349,N_967,N_1179);
nand U1350 (N_1350,N_1006,N_1044);
nand U1351 (N_1351,N_667,N_793);
nor U1352 (N_1352,N_669,N_947);
nor U1353 (N_1353,N_1157,N_858);
xnor U1354 (N_1354,N_785,N_1068);
or U1355 (N_1355,N_717,N_936);
and U1356 (N_1356,N_733,N_959);
or U1357 (N_1357,N_796,N_1056);
nand U1358 (N_1358,N_1025,N_979);
and U1359 (N_1359,N_1138,N_973);
nand U1360 (N_1360,N_916,N_759);
and U1361 (N_1361,N_716,N_780);
nand U1362 (N_1362,N_704,N_810);
and U1363 (N_1363,N_1173,N_836);
and U1364 (N_1364,N_627,N_1136);
nor U1365 (N_1365,N_1142,N_990);
nand U1366 (N_1366,N_746,N_817);
nor U1367 (N_1367,N_1190,N_748);
nand U1368 (N_1368,N_1074,N_1193);
and U1369 (N_1369,N_737,N_1076);
or U1370 (N_1370,N_706,N_890);
and U1371 (N_1371,N_1102,N_1191);
and U1372 (N_1372,N_624,N_807);
and U1373 (N_1373,N_646,N_829);
nor U1374 (N_1374,N_1176,N_855);
and U1375 (N_1375,N_762,N_862);
nor U1376 (N_1376,N_949,N_955);
nand U1377 (N_1377,N_932,N_790);
or U1378 (N_1378,N_969,N_715);
nor U1379 (N_1379,N_840,N_1031);
nand U1380 (N_1380,N_638,N_897);
and U1381 (N_1381,N_1196,N_1148);
nand U1382 (N_1382,N_869,N_801);
nand U1383 (N_1383,N_687,N_825);
nor U1384 (N_1384,N_602,N_1139);
or U1385 (N_1385,N_1093,N_754);
nand U1386 (N_1386,N_1096,N_636);
nand U1387 (N_1387,N_631,N_666);
nand U1388 (N_1388,N_1066,N_611);
or U1389 (N_1389,N_1089,N_726);
and U1390 (N_1390,N_873,N_939);
or U1391 (N_1391,N_783,N_883);
or U1392 (N_1392,N_972,N_1072);
or U1393 (N_1393,N_1016,N_838);
or U1394 (N_1394,N_815,N_672);
or U1395 (N_1395,N_1053,N_680);
nor U1396 (N_1396,N_948,N_701);
nand U1397 (N_1397,N_900,N_884);
or U1398 (N_1398,N_700,N_694);
xnor U1399 (N_1399,N_952,N_993);
or U1400 (N_1400,N_1022,N_848);
nor U1401 (N_1401,N_1158,N_1162);
nor U1402 (N_1402,N_774,N_1121);
nor U1403 (N_1403,N_887,N_1057);
nand U1404 (N_1404,N_1126,N_698);
nor U1405 (N_1405,N_912,N_671);
and U1406 (N_1406,N_1141,N_1168);
nor U1407 (N_1407,N_820,N_943);
and U1408 (N_1408,N_803,N_915);
or U1409 (N_1409,N_615,N_1029);
nor U1410 (N_1410,N_965,N_1171);
nand U1411 (N_1411,N_1104,N_604);
nand U1412 (N_1412,N_1064,N_628);
xnor U1413 (N_1413,N_610,N_1175);
nand U1414 (N_1414,N_730,N_643);
and U1415 (N_1415,N_827,N_831);
and U1416 (N_1416,N_963,N_1140);
nand U1417 (N_1417,N_1111,N_1167);
nand U1418 (N_1418,N_1013,N_1084);
and U1419 (N_1419,N_692,N_1119);
and U1420 (N_1420,N_798,N_679);
nor U1421 (N_1421,N_1163,N_997);
xor U1422 (N_1422,N_653,N_881);
nor U1423 (N_1423,N_1100,N_709);
nor U1424 (N_1424,N_882,N_799);
nor U1425 (N_1425,N_736,N_607);
nor U1426 (N_1426,N_1000,N_674);
and U1427 (N_1427,N_606,N_953);
and U1428 (N_1428,N_975,N_1052);
and U1429 (N_1429,N_612,N_970);
nor U1430 (N_1430,N_804,N_1177);
nor U1431 (N_1431,N_1050,N_1174);
nand U1432 (N_1432,N_809,N_734);
nor U1433 (N_1433,N_1032,N_655);
nand U1434 (N_1434,N_1161,N_983);
nand U1435 (N_1435,N_899,N_1186);
nor U1436 (N_1436,N_1098,N_1069);
nand U1437 (N_1437,N_682,N_908);
and U1438 (N_1438,N_725,N_988);
nand U1439 (N_1439,N_1197,N_650);
or U1440 (N_1440,N_656,N_1008);
nor U1441 (N_1441,N_819,N_1023);
and U1442 (N_1442,N_1001,N_958);
and U1443 (N_1443,N_877,N_999);
and U1444 (N_1444,N_1151,N_1178);
nor U1445 (N_1445,N_675,N_1007);
and U1446 (N_1446,N_857,N_929);
nor U1447 (N_1447,N_641,N_1099);
nand U1448 (N_1448,N_893,N_876);
nand U1449 (N_1449,N_860,N_1107);
nand U1450 (N_1450,N_1027,N_998);
or U1451 (N_1451,N_1039,N_782);
or U1452 (N_1452,N_1150,N_928);
or U1453 (N_1453,N_823,N_617);
and U1454 (N_1454,N_630,N_1160);
nor U1455 (N_1455,N_1036,N_889);
and U1456 (N_1456,N_1122,N_728);
nor U1457 (N_1457,N_664,N_794);
and U1458 (N_1458,N_657,N_880);
and U1459 (N_1459,N_1134,N_991);
and U1460 (N_1460,N_1146,N_960);
or U1461 (N_1461,N_898,N_608);
or U1462 (N_1462,N_1170,N_752);
nor U1463 (N_1463,N_934,N_629);
and U1464 (N_1464,N_661,N_1128);
and U1465 (N_1465,N_985,N_1156);
nor U1466 (N_1466,N_1166,N_673);
or U1467 (N_1467,N_648,N_652);
and U1468 (N_1468,N_741,N_1145);
or U1469 (N_1469,N_731,N_1135);
or U1470 (N_1470,N_744,N_1184);
and U1471 (N_1471,N_1137,N_718);
nor U1472 (N_1472,N_1090,N_755);
or U1473 (N_1473,N_851,N_910);
and U1474 (N_1474,N_614,N_1112);
and U1475 (N_1475,N_702,N_976);
nand U1476 (N_1476,N_695,N_773);
or U1477 (N_1477,N_1041,N_822);
or U1478 (N_1478,N_601,N_693);
nand U1479 (N_1479,N_811,N_651);
and U1480 (N_1480,N_968,N_1164);
and U1481 (N_1481,N_721,N_974);
and U1482 (N_1482,N_776,N_1101);
nand U1483 (N_1483,N_727,N_802);
nand U1484 (N_1484,N_777,N_1014);
nor U1485 (N_1485,N_642,N_913);
or U1486 (N_1486,N_723,N_950);
and U1487 (N_1487,N_1105,N_1002);
nor U1488 (N_1488,N_1120,N_714);
nor U1489 (N_1489,N_1172,N_1114);
nand U1490 (N_1490,N_832,N_859);
or U1491 (N_1491,N_691,N_874);
nand U1492 (N_1492,N_834,N_1060);
nor U1493 (N_1493,N_1035,N_805);
nor U1494 (N_1494,N_863,N_870);
and U1495 (N_1495,N_813,N_633);
nor U1496 (N_1496,N_732,N_847);
nor U1497 (N_1497,N_980,N_1125);
and U1498 (N_1498,N_905,N_930);
or U1499 (N_1499,N_994,N_745);
nand U1500 (N_1500,N_864,N_681);
and U1501 (N_1501,N_885,N_758);
nor U1502 (N_1502,N_699,N_986);
nand U1503 (N_1503,N_961,N_657);
nor U1504 (N_1504,N_1124,N_1134);
and U1505 (N_1505,N_1037,N_697);
nand U1506 (N_1506,N_967,N_696);
nor U1507 (N_1507,N_859,N_976);
and U1508 (N_1508,N_628,N_1038);
and U1509 (N_1509,N_645,N_969);
and U1510 (N_1510,N_1055,N_1184);
nand U1511 (N_1511,N_998,N_805);
nor U1512 (N_1512,N_1178,N_871);
or U1513 (N_1513,N_615,N_705);
and U1514 (N_1514,N_869,N_784);
nand U1515 (N_1515,N_795,N_1102);
nor U1516 (N_1516,N_678,N_1181);
nor U1517 (N_1517,N_710,N_1001);
nand U1518 (N_1518,N_878,N_963);
or U1519 (N_1519,N_721,N_1191);
or U1520 (N_1520,N_955,N_764);
or U1521 (N_1521,N_774,N_1040);
nand U1522 (N_1522,N_886,N_1077);
and U1523 (N_1523,N_1191,N_1169);
nand U1524 (N_1524,N_1191,N_730);
and U1525 (N_1525,N_1132,N_607);
and U1526 (N_1526,N_903,N_658);
nand U1527 (N_1527,N_668,N_641);
nor U1528 (N_1528,N_866,N_918);
or U1529 (N_1529,N_602,N_1119);
or U1530 (N_1530,N_1196,N_958);
nand U1531 (N_1531,N_993,N_859);
nor U1532 (N_1532,N_664,N_1023);
nor U1533 (N_1533,N_676,N_1037);
or U1534 (N_1534,N_962,N_732);
or U1535 (N_1535,N_1104,N_636);
and U1536 (N_1536,N_605,N_1191);
and U1537 (N_1537,N_1087,N_957);
and U1538 (N_1538,N_977,N_855);
and U1539 (N_1539,N_1020,N_732);
and U1540 (N_1540,N_1099,N_636);
nand U1541 (N_1541,N_977,N_1024);
or U1542 (N_1542,N_662,N_961);
nor U1543 (N_1543,N_1098,N_624);
and U1544 (N_1544,N_1168,N_977);
or U1545 (N_1545,N_725,N_1124);
nor U1546 (N_1546,N_995,N_1185);
nor U1547 (N_1547,N_628,N_618);
or U1548 (N_1548,N_800,N_759);
xnor U1549 (N_1549,N_812,N_739);
or U1550 (N_1550,N_1133,N_1075);
nor U1551 (N_1551,N_1111,N_1006);
nand U1552 (N_1552,N_1035,N_1043);
nor U1553 (N_1553,N_780,N_766);
and U1554 (N_1554,N_1013,N_850);
and U1555 (N_1555,N_651,N_769);
and U1556 (N_1556,N_877,N_705);
and U1557 (N_1557,N_715,N_615);
and U1558 (N_1558,N_950,N_1180);
xnor U1559 (N_1559,N_741,N_947);
nor U1560 (N_1560,N_961,N_1117);
nor U1561 (N_1561,N_659,N_847);
and U1562 (N_1562,N_602,N_1047);
or U1563 (N_1563,N_1093,N_1092);
nand U1564 (N_1564,N_819,N_898);
nand U1565 (N_1565,N_911,N_953);
or U1566 (N_1566,N_674,N_875);
and U1567 (N_1567,N_984,N_720);
or U1568 (N_1568,N_1029,N_1142);
nor U1569 (N_1569,N_1041,N_1069);
or U1570 (N_1570,N_829,N_850);
nor U1571 (N_1571,N_966,N_665);
nand U1572 (N_1572,N_701,N_983);
nand U1573 (N_1573,N_1113,N_1194);
or U1574 (N_1574,N_751,N_1051);
or U1575 (N_1575,N_1028,N_871);
nand U1576 (N_1576,N_983,N_1059);
nor U1577 (N_1577,N_1190,N_818);
and U1578 (N_1578,N_759,N_785);
nand U1579 (N_1579,N_1043,N_778);
and U1580 (N_1580,N_675,N_1004);
and U1581 (N_1581,N_795,N_1139);
and U1582 (N_1582,N_767,N_731);
or U1583 (N_1583,N_904,N_790);
nand U1584 (N_1584,N_899,N_1016);
or U1585 (N_1585,N_671,N_895);
or U1586 (N_1586,N_1022,N_1199);
nor U1587 (N_1587,N_1121,N_1166);
nor U1588 (N_1588,N_853,N_835);
and U1589 (N_1589,N_1128,N_828);
and U1590 (N_1590,N_1029,N_677);
nand U1591 (N_1591,N_685,N_743);
and U1592 (N_1592,N_616,N_790);
and U1593 (N_1593,N_945,N_927);
nor U1594 (N_1594,N_624,N_1029);
nor U1595 (N_1595,N_766,N_1070);
or U1596 (N_1596,N_1090,N_1074);
or U1597 (N_1597,N_921,N_1065);
nand U1598 (N_1598,N_976,N_630);
nor U1599 (N_1599,N_635,N_633);
or U1600 (N_1600,N_676,N_905);
nor U1601 (N_1601,N_651,N_1047);
nor U1602 (N_1602,N_945,N_1038);
nor U1603 (N_1603,N_782,N_604);
or U1604 (N_1604,N_1122,N_1058);
or U1605 (N_1605,N_853,N_740);
nor U1606 (N_1606,N_1058,N_929);
or U1607 (N_1607,N_949,N_1111);
nor U1608 (N_1608,N_728,N_677);
nand U1609 (N_1609,N_857,N_767);
nor U1610 (N_1610,N_1179,N_701);
and U1611 (N_1611,N_1053,N_1076);
or U1612 (N_1612,N_662,N_907);
nor U1613 (N_1613,N_748,N_1064);
and U1614 (N_1614,N_876,N_680);
nor U1615 (N_1615,N_1195,N_831);
nor U1616 (N_1616,N_1136,N_1019);
or U1617 (N_1617,N_740,N_795);
nor U1618 (N_1618,N_1079,N_1120);
and U1619 (N_1619,N_803,N_1013);
or U1620 (N_1620,N_959,N_678);
or U1621 (N_1621,N_798,N_1088);
nor U1622 (N_1622,N_812,N_833);
and U1623 (N_1623,N_1136,N_1062);
nor U1624 (N_1624,N_818,N_1128);
or U1625 (N_1625,N_1114,N_823);
or U1626 (N_1626,N_821,N_1073);
nor U1627 (N_1627,N_938,N_746);
or U1628 (N_1628,N_778,N_859);
nor U1629 (N_1629,N_944,N_749);
nor U1630 (N_1630,N_1109,N_753);
or U1631 (N_1631,N_996,N_987);
or U1632 (N_1632,N_602,N_922);
and U1633 (N_1633,N_614,N_917);
or U1634 (N_1634,N_661,N_696);
nand U1635 (N_1635,N_708,N_998);
nand U1636 (N_1636,N_632,N_882);
and U1637 (N_1637,N_825,N_623);
and U1638 (N_1638,N_1118,N_925);
nand U1639 (N_1639,N_939,N_1035);
and U1640 (N_1640,N_859,N_1121);
and U1641 (N_1641,N_804,N_1025);
nand U1642 (N_1642,N_1050,N_785);
nor U1643 (N_1643,N_766,N_833);
nand U1644 (N_1644,N_737,N_1086);
nor U1645 (N_1645,N_778,N_1031);
nand U1646 (N_1646,N_649,N_1181);
or U1647 (N_1647,N_1097,N_891);
nand U1648 (N_1648,N_882,N_1000);
nand U1649 (N_1649,N_772,N_1033);
and U1650 (N_1650,N_1146,N_1135);
nand U1651 (N_1651,N_966,N_706);
nor U1652 (N_1652,N_621,N_1050);
or U1653 (N_1653,N_616,N_904);
nand U1654 (N_1654,N_775,N_1028);
and U1655 (N_1655,N_1084,N_644);
nor U1656 (N_1656,N_740,N_942);
nand U1657 (N_1657,N_1158,N_877);
nand U1658 (N_1658,N_824,N_605);
nor U1659 (N_1659,N_1000,N_981);
nor U1660 (N_1660,N_1193,N_887);
nand U1661 (N_1661,N_981,N_672);
and U1662 (N_1662,N_1030,N_1040);
xnor U1663 (N_1663,N_817,N_1103);
or U1664 (N_1664,N_923,N_932);
nand U1665 (N_1665,N_819,N_789);
nand U1666 (N_1666,N_1041,N_872);
nor U1667 (N_1667,N_866,N_987);
nor U1668 (N_1668,N_1047,N_705);
and U1669 (N_1669,N_906,N_682);
nor U1670 (N_1670,N_1097,N_978);
and U1671 (N_1671,N_1063,N_1197);
and U1672 (N_1672,N_909,N_731);
and U1673 (N_1673,N_1051,N_884);
and U1674 (N_1674,N_1036,N_854);
nor U1675 (N_1675,N_654,N_985);
or U1676 (N_1676,N_1034,N_759);
or U1677 (N_1677,N_855,N_710);
and U1678 (N_1678,N_1025,N_763);
nor U1679 (N_1679,N_663,N_1037);
nand U1680 (N_1680,N_1002,N_650);
and U1681 (N_1681,N_819,N_647);
and U1682 (N_1682,N_676,N_1049);
and U1683 (N_1683,N_606,N_818);
nor U1684 (N_1684,N_1146,N_788);
nand U1685 (N_1685,N_1058,N_994);
nor U1686 (N_1686,N_1028,N_629);
nand U1687 (N_1687,N_719,N_814);
nand U1688 (N_1688,N_602,N_800);
or U1689 (N_1689,N_610,N_792);
nand U1690 (N_1690,N_1070,N_621);
and U1691 (N_1691,N_782,N_1116);
nor U1692 (N_1692,N_928,N_629);
nand U1693 (N_1693,N_756,N_993);
nand U1694 (N_1694,N_1169,N_1015);
nor U1695 (N_1695,N_1176,N_764);
or U1696 (N_1696,N_627,N_615);
nor U1697 (N_1697,N_671,N_810);
and U1698 (N_1698,N_736,N_939);
nand U1699 (N_1699,N_1161,N_1136);
nand U1700 (N_1700,N_790,N_882);
or U1701 (N_1701,N_652,N_697);
nor U1702 (N_1702,N_1037,N_1058);
or U1703 (N_1703,N_1147,N_794);
nor U1704 (N_1704,N_1177,N_1040);
nand U1705 (N_1705,N_1199,N_822);
nand U1706 (N_1706,N_603,N_1102);
nor U1707 (N_1707,N_801,N_1108);
nor U1708 (N_1708,N_985,N_623);
nand U1709 (N_1709,N_834,N_646);
nor U1710 (N_1710,N_1054,N_1179);
nor U1711 (N_1711,N_1177,N_1069);
nor U1712 (N_1712,N_1158,N_1002);
or U1713 (N_1713,N_806,N_609);
nand U1714 (N_1714,N_1048,N_913);
or U1715 (N_1715,N_933,N_953);
and U1716 (N_1716,N_1152,N_1158);
and U1717 (N_1717,N_1065,N_908);
or U1718 (N_1718,N_751,N_681);
nor U1719 (N_1719,N_1055,N_973);
nor U1720 (N_1720,N_1018,N_717);
and U1721 (N_1721,N_1062,N_1018);
or U1722 (N_1722,N_622,N_866);
or U1723 (N_1723,N_1151,N_1086);
nand U1724 (N_1724,N_671,N_767);
nor U1725 (N_1725,N_875,N_1139);
or U1726 (N_1726,N_944,N_824);
or U1727 (N_1727,N_626,N_788);
nor U1728 (N_1728,N_858,N_1098);
or U1729 (N_1729,N_752,N_740);
nor U1730 (N_1730,N_937,N_734);
nand U1731 (N_1731,N_1143,N_1120);
nand U1732 (N_1732,N_956,N_1039);
or U1733 (N_1733,N_1099,N_869);
nor U1734 (N_1734,N_1076,N_891);
or U1735 (N_1735,N_651,N_1013);
nor U1736 (N_1736,N_826,N_604);
nand U1737 (N_1737,N_901,N_1009);
and U1738 (N_1738,N_833,N_999);
nor U1739 (N_1739,N_642,N_1071);
and U1740 (N_1740,N_824,N_668);
nor U1741 (N_1741,N_848,N_968);
and U1742 (N_1742,N_710,N_794);
or U1743 (N_1743,N_947,N_1010);
xor U1744 (N_1744,N_899,N_880);
and U1745 (N_1745,N_1093,N_875);
nor U1746 (N_1746,N_1186,N_847);
nor U1747 (N_1747,N_1131,N_888);
and U1748 (N_1748,N_747,N_680);
nor U1749 (N_1749,N_682,N_678);
nor U1750 (N_1750,N_1188,N_744);
nor U1751 (N_1751,N_600,N_1158);
or U1752 (N_1752,N_998,N_914);
nor U1753 (N_1753,N_1114,N_841);
and U1754 (N_1754,N_800,N_872);
and U1755 (N_1755,N_928,N_1017);
or U1756 (N_1756,N_679,N_724);
nor U1757 (N_1757,N_1055,N_988);
nand U1758 (N_1758,N_1073,N_689);
and U1759 (N_1759,N_1062,N_670);
nand U1760 (N_1760,N_723,N_1092);
and U1761 (N_1761,N_896,N_687);
and U1762 (N_1762,N_1032,N_986);
nand U1763 (N_1763,N_1096,N_751);
nor U1764 (N_1764,N_1167,N_941);
xor U1765 (N_1765,N_1096,N_949);
and U1766 (N_1766,N_1010,N_1018);
and U1767 (N_1767,N_887,N_940);
or U1768 (N_1768,N_1179,N_1041);
and U1769 (N_1769,N_813,N_981);
and U1770 (N_1770,N_697,N_931);
or U1771 (N_1771,N_933,N_1190);
and U1772 (N_1772,N_789,N_630);
and U1773 (N_1773,N_610,N_788);
nor U1774 (N_1774,N_848,N_839);
or U1775 (N_1775,N_634,N_613);
nand U1776 (N_1776,N_1030,N_1133);
or U1777 (N_1777,N_766,N_942);
or U1778 (N_1778,N_757,N_735);
xnor U1779 (N_1779,N_836,N_934);
or U1780 (N_1780,N_721,N_634);
nor U1781 (N_1781,N_1043,N_859);
or U1782 (N_1782,N_866,N_1170);
nor U1783 (N_1783,N_1115,N_697);
nor U1784 (N_1784,N_948,N_1143);
and U1785 (N_1785,N_804,N_724);
nor U1786 (N_1786,N_907,N_841);
or U1787 (N_1787,N_939,N_1024);
xnor U1788 (N_1788,N_932,N_885);
or U1789 (N_1789,N_967,N_1117);
or U1790 (N_1790,N_1047,N_887);
nand U1791 (N_1791,N_1061,N_1040);
nor U1792 (N_1792,N_895,N_686);
or U1793 (N_1793,N_715,N_885);
nand U1794 (N_1794,N_745,N_846);
nand U1795 (N_1795,N_684,N_777);
nand U1796 (N_1796,N_1007,N_854);
or U1797 (N_1797,N_1150,N_966);
and U1798 (N_1798,N_667,N_1171);
nand U1799 (N_1799,N_916,N_1126);
or U1800 (N_1800,N_1419,N_1558);
nor U1801 (N_1801,N_1719,N_1795);
or U1802 (N_1802,N_1573,N_1352);
and U1803 (N_1803,N_1268,N_1298);
nand U1804 (N_1804,N_1338,N_1582);
nor U1805 (N_1805,N_1653,N_1743);
or U1806 (N_1806,N_1637,N_1206);
or U1807 (N_1807,N_1715,N_1713);
or U1808 (N_1808,N_1797,N_1485);
or U1809 (N_1809,N_1351,N_1335);
and U1810 (N_1810,N_1496,N_1207);
or U1811 (N_1811,N_1742,N_1315);
nor U1812 (N_1812,N_1477,N_1424);
nand U1813 (N_1813,N_1394,N_1384);
nor U1814 (N_1814,N_1473,N_1413);
nor U1815 (N_1815,N_1468,N_1537);
or U1816 (N_1816,N_1617,N_1684);
and U1817 (N_1817,N_1492,N_1505);
nand U1818 (N_1818,N_1423,N_1318);
nor U1819 (N_1819,N_1527,N_1396);
nand U1820 (N_1820,N_1345,N_1217);
or U1821 (N_1821,N_1578,N_1604);
nor U1822 (N_1822,N_1766,N_1717);
or U1823 (N_1823,N_1470,N_1326);
and U1824 (N_1824,N_1436,N_1619);
and U1825 (N_1825,N_1567,N_1562);
and U1826 (N_1826,N_1263,N_1392);
or U1827 (N_1827,N_1373,N_1220);
and U1828 (N_1828,N_1618,N_1565);
or U1829 (N_1829,N_1260,N_1560);
and U1830 (N_1830,N_1610,N_1606);
and U1831 (N_1831,N_1669,N_1639);
or U1832 (N_1832,N_1257,N_1445);
nand U1833 (N_1833,N_1512,N_1698);
nand U1834 (N_1834,N_1301,N_1236);
nor U1835 (N_1835,N_1375,N_1239);
nand U1836 (N_1836,N_1313,N_1320);
nor U1837 (N_1837,N_1678,N_1358);
nor U1838 (N_1838,N_1353,N_1398);
and U1839 (N_1839,N_1299,N_1613);
nor U1840 (N_1840,N_1689,N_1407);
or U1841 (N_1841,N_1750,N_1533);
xor U1842 (N_1842,N_1446,N_1339);
and U1843 (N_1843,N_1574,N_1620);
or U1844 (N_1844,N_1550,N_1551);
nand U1845 (N_1845,N_1685,N_1723);
nor U1846 (N_1846,N_1223,N_1648);
and U1847 (N_1847,N_1579,N_1690);
or U1848 (N_1848,N_1705,N_1366);
and U1849 (N_1849,N_1623,N_1385);
or U1850 (N_1850,N_1201,N_1367);
or U1851 (N_1851,N_1788,N_1203);
or U1852 (N_1852,N_1777,N_1302);
and U1853 (N_1853,N_1547,N_1314);
nand U1854 (N_1854,N_1494,N_1770);
and U1855 (N_1855,N_1549,N_1234);
and U1856 (N_1856,N_1703,N_1218);
nor U1857 (N_1857,N_1586,N_1645);
and U1858 (N_1858,N_1691,N_1249);
nand U1859 (N_1859,N_1670,N_1590);
nor U1860 (N_1860,N_1452,N_1232);
nand U1861 (N_1861,N_1487,N_1341);
nor U1862 (N_1862,N_1509,N_1288);
and U1863 (N_1863,N_1484,N_1675);
and U1864 (N_1864,N_1513,N_1526);
nor U1865 (N_1865,N_1229,N_1405);
nand U1866 (N_1866,N_1228,N_1621);
nand U1867 (N_1867,N_1528,N_1532);
or U1868 (N_1868,N_1246,N_1332);
and U1869 (N_1869,N_1215,N_1486);
nor U1870 (N_1870,N_1605,N_1278);
nand U1871 (N_1871,N_1601,N_1216);
and U1872 (N_1872,N_1269,N_1430);
nor U1873 (N_1873,N_1401,N_1438);
nor U1874 (N_1874,N_1741,N_1603);
nor U1875 (N_1875,N_1383,N_1535);
nor U1876 (N_1876,N_1589,N_1235);
nor U1877 (N_1877,N_1754,N_1388);
and U1878 (N_1878,N_1292,N_1611);
nand U1879 (N_1879,N_1785,N_1327);
nor U1880 (N_1880,N_1700,N_1525);
or U1881 (N_1881,N_1672,N_1219);
nor U1882 (N_1882,N_1556,N_1790);
nand U1883 (N_1883,N_1270,N_1518);
nand U1884 (N_1884,N_1646,N_1224);
and U1885 (N_1885,N_1557,N_1540);
nor U1886 (N_1886,N_1647,N_1328);
nor U1887 (N_1887,N_1696,N_1765);
nand U1888 (N_1888,N_1248,N_1774);
nand U1889 (N_1889,N_1222,N_1382);
and U1890 (N_1890,N_1522,N_1546);
or U1891 (N_1891,N_1297,N_1478);
and U1892 (N_1892,N_1208,N_1410);
nor U1893 (N_1893,N_1364,N_1609);
nor U1894 (N_1894,N_1439,N_1480);
or U1895 (N_1895,N_1497,N_1592);
nand U1896 (N_1896,N_1399,N_1429);
or U1897 (N_1897,N_1584,N_1283);
and U1898 (N_1898,N_1440,N_1200);
nand U1899 (N_1899,N_1659,N_1416);
nor U1900 (N_1900,N_1306,N_1371);
and U1901 (N_1901,N_1390,N_1799);
and U1902 (N_1902,N_1671,N_1643);
nand U1903 (N_1903,N_1425,N_1250);
nor U1904 (N_1904,N_1724,N_1627);
nor U1905 (N_1905,N_1340,N_1657);
nor U1906 (N_1906,N_1679,N_1458);
and U1907 (N_1907,N_1251,N_1597);
nor U1908 (N_1908,N_1787,N_1444);
or U1909 (N_1909,N_1295,N_1233);
nor U1910 (N_1910,N_1760,N_1329);
and U1911 (N_1911,N_1707,N_1252);
nand U1912 (N_1912,N_1402,N_1644);
or U1913 (N_1913,N_1596,N_1662);
and U1914 (N_1914,N_1769,N_1291);
nor U1915 (N_1915,N_1581,N_1431);
and U1916 (N_1916,N_1726,N_1414);
or U1917 (N_1917,N_1706,N_1534);
and U1918 (N_1918,N_1368,N_1363);
nand U1919 (N_1919,N_1391,N_1650);
nor U1920 (N_1920,N_1334,N_1516);
nor U1921 (N_1921,N_1290,N_1608);
nand U1922 (N_1922,N_1677,N_1602);
or U1923 (N_1923,N_1658,N_1475);
or U1924 (N_1924,N_1781,N_1293);
and U1925 (N_1925,N_1759,N_1272);
and U1926 (N_1926,N_1721,N_1515);
nand U1927 (N_1927,N_1740,N_1361);
xnor U1928 (N_1928,N_1455,N_1273);
or U1929 (N_1929,N_1541,N_1791);
nand U1930 (N_1930,N_1792,N_1312);
and U1931 (N_1931,N_1214,N_1409);
nand U1932 (N_1932,N_1271,N_1593);
nand U1933 (N_1933,N_1519,N_1266);
and U1934 (N_1934,N_1555,N_1701);
and U1935 (N_1935,N_1728,N_1450);
and U1936 (N_1936,N_1751,N_1282);
nor U1937 (N_1937,N_1511,N_1393);
nor U1938 (N_1938,N_1433,N_1231);
nand U1939 (N_1939,N_1694,N_1674);
nor U1940 (N_1940,N_1735,N_1552);
or U1941 (N_1941,N_1680,N_1521);
xnor U1942 (N_1942,N_1316,N_1309);
or U1943 (N_1943,N_1712,N_1542);
and U1944 (N_1944,N_1607,N_1744);
and U1945 (N_1945,N_1568,N_1614);
nand U1946 (N_1946,N_1704,N_1622);
nor U1947 (N_1947,N_1506,N_1630);
xor U1948 (N_1948,N_1559,N_1422);
nor U1949 (N_1949,N_1481,N_1600);
nor U1950 (N_1950,N_1508,N_1255);
nand U1951 (N_1951,N_1336,N_1595);
and U1952 (N_1952,N_1262,N_1369);
or U1953 (N_1953,N_1441,N_1253);
and U1954 (N_1954,N_1380,N_1664);
nand U1955 (N_1955,N_1554,N_1775);
nor U1956 (N_1956,N_1773,N_1544);
nor U1957 (N_1957,N_1699,N_1665);
nand U1958 (N_1958,N_1654,N_1265);
and U1959 (N_1959,N_1274,N_1570);
nor U1960 (N_1960,N_1771,N_1448);
nor U1961 (N_1961,N_1462,N_1503);
nand U1962 (N_1962,N_1786,N_1676);
nand U1963 (N_1963,N_1756,N_1354);
or U1964 (N_1964,N_1330,N_1510);
or U1965 (N_1965,N_1612,N_1240);
and U1966 (N_1966,N_1548,N_1718);
nand U1967 (N_1967,N_1649,N_1632);
and U1968 (N_1968,N_1447,N_1634);
nand U1969 (N_1969,N_1247,N_1357);
nand U1970 (N_1970,N_1711,N_1243);
nand U1971 (N_1971,N_1668,N_1736);
or U1972 (N_1972,N_1378,N_1564);
nor U1973 (N_1973,N_1673,N_1545);
or U1974 (N_1974,N_1529,N_1794);
and U1975 (N_1975,N_1488,N_1709);
and U1976 (N_1976,N_1418,N_1764);
nor U1977 (N_1977,N_1594,N_1708);
or U1978 (N_1978,N_1289,N_1238);
nor U1979 (N_1979,N_1737,N_1780);
and U1980 (N_1980,N_1426,N_1501);
and U1981 (N_1981,N_1482,N_1403);
or U1982 (N_1982,N_1520,N_1379);
and U1983 (N_1983,N_1517,N_1267);
nand U1984 (N_1984,N_1507,N_1796);
nor U1985 (N_1985,N_1287,N_1575);
nand U1986 (N_1986,N_1286,N_1748);
and U1987 (N_1987,N_1308,N_1479);
nand U1988 (N_1988,N_1281,N_1307);
nand U1989 (N_1989,N_1702,N_1628);
or U1990 (N_1990,N_1538,N_1710);
or U1991 (N_1991,N_1204,N_1294);
nand U1992 (N_1992,N_1625,N_1317);
or U1993 (N_1993,N_1276,N_1230);
nand U1994 (N_1994,N_1638,N_1563);
and U1995 (N_1995,N_1395,N_1599);
nor U1996 (N_1996,N_1733,N_1310);
and U1997 (N_1997,N_1783,N_1355);
and U1998 (N_1998,N_1681,N_1370);
and U1999 (N_1999,N_1209,N_1725);
nor U2000 (N_2000,N_1322,N_1210);
or U2001 (N_2001,N_1303,N_1530);
nor U2002 (N_2002,N_1640,N_1453);
and U2003 (N_2003,N_1729,N_1536);
nor U2004 (N_2004,N_1569,N_1739);
or U2005 (N_2005,N_1738,N_1523);
or U2006 (N_2006,N_1432,N_1434);
nor U2007 (N_2007,N_1227,N_1779);
nand U2008 (N_2008,N_1465,N_1346);
and U2009 (N_2009,N_1793,N_1349);
or U2010 (N_2010,N_1212,N_1767);
nor U2011 (N_2011,N_1504,N_1254);
nand U2012 (N_2012,N_1311,N_1731);
and U2013 (N_2013,N_1763,N_1730);
nor U2014 (N_2014,N_1758,N_1456);
nand U2015 (N_2015,N_1258,N_1304);
and U2016 (N_2016,N_1615,N_1296);
and U2017 (N_2017,N_1397,N_1350);
and U2018 (N_2018,N_1524,N_1400);
nand U2019 (N_2019,N_1261,N_1587);
or U2020 (N_2020,N_1459,N_1588);
and U2021 (N_2021,N_1749,N_1531);
nand U2022 (N_2022,N_1333,N_1500);
nor U2023 (N_2023,N_1277,N_1359);
nand U2024 (N_2024,N_1577,N_1467);
nand U2025 (N_2025,N_1420,N_1585);
and U2026 (N_2026,N_1331,N_1376);
xnor U2027 (N_2027,N_1716,N_1490);
nor U2028 (N_2028,N_1275,N_1344);
xnor U2029 (N_2029,N_1761,N_1360);
or U2030 (N_2030,N_1469,N_1576);
nor U2031 (N_2031,N_1747,N_1571);
and U2032 (N_2032,N_1583,N_1714);
or U2033 (N_2033,N_1543,N_1415);
or U2034 (N_2034,N_1381,N_1451);
or U2035 (N_2035,N_1242,N_1221);
or U2036 (N_2036,N_1474,N_1687);
nor U2037 (N_2037,N_1553,N_1651);
and U2038 (N_2038,N_1461,N_1225);
or U2039 (N_2039,N_1305,N_1321);
nor U2040 (N_2040,N_1493,N_1652);
or U2041 (N_2041,N_1372,N_1778);
nor U2042 (N_2042,N_1237,N_1757);
nor U2043 (N_2043,N_1631,N_1566);
nand U2044 (N_2044,N_1411,N_1406);
and U2045 (N_2045,N_1755,N_1768);
and U2046 (N_2046,N_1449,N_1337);
and U2047 (N_2047,N_1663,N_1211);
nor U2048 (N_2048,N_1435,N_1661);
or U2049 (N_2049,N_1457,N_1324);
nand U2050 (N_2050,N_1417,N_1695);
nand U2051 (N_2051,N_1244,N_1580);
or U2052 (N_2052,N_1561,N_1362);
nand U2053 (N_2053,N_1682,N_1624);
xor U2054 (N_2054,N_1591,N_1259);
nand U2055 (N_2055,N_1202,N_1374);
or U2056 (N_2056,N_1464,N_1343);
nor U2057 (N_2057,N_1772,N_1629);
or U2058 (N_2058,N_1745,N_1746);
nand U2059 (N_2059,N_1514,N_1693);
or U2060 (N_2060,N_1720,N_1442);
nand U2061 (N_2061,N_1280,N_1734);
nor U2062 (N_2062,N_1683,N_1408);
nor U2063 (N_2063,N_1466,N_1776);
nand U2064 (N_2064,N_1598,N_1782);
nor U2065 (N_2065,N_1472,N_1427);
or U2066 (N_2066,N_1498,N_1688);
nor U2067 (N_2067,N_1641,N_1460);
nand U2068 (N_2068,N_1642,N_1489);
nand U2069 (N_2069,N_1471,N_1762);
or U2070 (N_2070,N_1437,N_1245);
nor U2071 (N_2071,N_1300,N_1491);
nor U2072 (N_2072,N_1365,N_1347);
or U2073 (N_2073,N_1404,N_1752);
and U2074 (N_2074,N_1722,N_1377);
nor U2075 (N_2075,N_1443,N_1284);
nor U2076 (N_2076,N_1463,N_1660);
and U2077 (N_2077,N_1572,N_1727);
nand U2078 (N_2078,N_1789,N_1213);
nor U2079 (N_2079,N_1784,N_1389);
nand U2080 (N_2080,N_1656,N_1256);
or U2081 (N_2081,N_1616,N_1692);
nand U2082 (N_2082,N_1636,N_1226);
nor U2083 (N_2083,N_1319,N_1666);
and U2084 (N_2084,N_1732,N_1483);
or U2085 (N_2085,N_1279,N_1633);
nand U2086 (N_2086,N_1476,N_1205);
or U2087 (N_2087,N_1241,N_1342);
and U2088 (N_2088,N_1798,N_1686);
and U2089 (N_2089,N_1495,N_1285);
or U2090 (N_2090,N_1356,N_1626);
and U2091 (N_2091,N_1323,N_1753);
or U2092 (N_2092,N_1539,N_1428);
and U2093 (N_2093,N_1454,N_1697);
and U2094 (N_2094,N_1386,N_1412);
or U2095 (N_2095,N_1387,N_1421);
nand U2096 (N_2096,N_1502,N_1655);
and U2097 (N_2097,N_1264,N_1325);
nor U2098 (N_2098,N_1635,N_1667);
and U2099 (N_2099,N_1348,N_1499);
nand U2100 (N_2100,N_1284,N_1231);
nand U2101 (N_2101,N_1244,N_1405);
nor U2102 (N_2102,N_1579,N_1506);
nand U2103 (N_2103,N_1282,N_1536);
nor U2104 (N_2104,N_1632,N_1719);
nor U2105 (N_2105,N_1429,N_1596);
and U2106 (N_2106,N_1608,N_1512);
nor U2107 (N_2107,N_1435,N_1769);
nor U2108 (N_2108,N_1214,N_1344);
nand U2109 (N_2109,N_1793,N_1553);
and U2110 (N_2110,N_1463,N_1340);
nand U2111 (N_2111,N_1418,N_1461);
nand U2112 (N_2112,N_1747,N_1333);
nor U2113 (N_2113,N_1483,N_1262);
and U2114 (N_2114,N_1469,N_1787);
or U2115 (N_2115,N_1352,N_1659);
or U2116 (N_2116,N_1439,N_1683);
or U2117 (N_2117,N_1701,N_1210);
or U2118 (N_2118,N_1766,N_1346);
nand U2119 (N_2119,N_1606,N_1762);
nor U2120 (N_2120,N_1243,N_1716);
or U2121 (N_2121,N_1282,N_1266);
and U2122 (N_2122,N_1490,N_1285);
nand U2123 (N_2123,N_1454,N_1247);
and U2124 (N_2124,N_1506,N_1237);
or U2125 (N_2125,N_1517,N_1792);
and U2126 (N_2126,N_1429,N_1371);
or U2127 (N_2127,N_1745,N_1753);
or U2128 (N_2128,N_1530,N_1766);
or U2129 (N_2129,N_1282,N_1264);
nand U2130 (N_2130,N_1554,N_1698);
or U2131 (N_2131,N_1302,N_1243);
and U2132 (N_2132,N_1622,N_1403);
nor U2133 (N_2133,N_1445,N_1289);
nand U2134 (N_2134,N_1757,N_1451);
nand U2135 (N_2135,N_1324,N_1637);
nor U2136 (N_2136,N_1335,N_1470);
nor U2137 (N_2137,N_1506,N_1536);
nor U2138 (N_2138,N_1452,N_1370);
nor U2139 (N_2139,N_1208,N_1358);
or U2140 (N_2140,N_1335,N_1635);
nor U2141 (N_2141,N_1584,N_1237);
nor U2142 (N_2142,N_1680,N_1221);
nor U2143 (N_2143,N_1422,N_1339);
nand U2144 (N_2144,N_1363,N_1596);
nor U2145 (N_2145,N_1582,N_1272);
or U2146 (N_2146,N_1316,N_1384);
or U2147 (N_2147,N_1527,N_1342);
nand U2148 (N_2148,N_1799,N_1678);
nor U2149 (N_2149,N_1489,N_1512);
nand U2150 (N_2150,N_1635,N_1701);
or U2151 (N_2151,N_1708,N_1299);
and U2152 (N_2152,N_1497,N_1279);
nor U2153 (N_2153,N_1609,N_1564);
or U2154 (N_2154,N_1612,N_1577);
or U2155 (N_2155,N_1361,N_1332);
and U2156 (N_2156,N_1567,N_1775);
or U2157 (N_2157,N_1231,N_1776);
and U2158 (N_2158,N_1793,N_1593);
or U2159 (N_2159,N_1759,N_1293);
or U2160 (N_2160,N_1676,N_1413);
and U2161 (N_2161,N_1727,N_1315);
nor U2162 (N_2162,N_1321,N_1625);
nand U2163 (N_2163,N_1622,N_1340);
nand U2164 (N_2164,N_1376,N_1701);
nor U2165 (N_2165,N_1682,N_1699);
nand U2166 (N_2166,N_1247,N_1390);
nand U2167 (N_2167,N_1787,N_1339);
nand U2168 (N_2168,N_1577,N_1466);
or U2169 (N_2169,N_1294,N_1725);
nor U2170 (N_2170,N_1331,N_1383);
nand U2171 (N_2171,N_1376,N_1223);
nand U2172 (N_2172,N_1544,N_1492);
and U2173 (N_2173,N_1460,N_1502);
and U2174 (N_2174,N_1497,N_1337);
or U2175 (N_2175,N_1564,N_1371);
nor U2176 (N_2176,N_1483,N_1637);
nor U2177 (N_2177,N_1474,N_1399);
nand U2178 (N_2178,N_1676,N_1444);
and U2179 (N_2179,N_1423,N_1616);
nand U2180 (N_2180,N_1767,N_1461);
nand U2181 (N_2181,N_1619,N_1569);
nand U2182 (N_2182,N_1608,N_1427);
nor U2183 (N_2183,N_1233,N_1694);
nand U2184 (N_2184,N_1254,N_1714);
and U2185 (N_2185,N_1297,N_1620);
nor U2186 (N_2186,N_1378,N_1682);
and U2187 (N_2187,N_1678,N_1632);
and U2188 (N_2188,N_1675,N_1754);
or U2189 (N_2189,N_1414,N_1442);
or U2190 (N_2190,N_1771,N_1514);
nor U2191 (N_2191,N_1741,N_1255);
or U2192 (N_2192,N_1399,N_1266);
nor U2193 (N_2193,N_1508,N_1246);
or U2194 (N_2194,N_1224,N_1520);
nor U2195 (N_2195,N_1685,N_1722);
nor U2196 (N_2196,N_1621,N_1738);
nand U2197 (N_2197,N_1235,N_1713);
or U2198 (N_2198,N_1299,N_1732);
nor U2199 (N_2199,N_1499,N_1554);
nand U2200 (N_2200,N_1251,N_1408);
and U2201 (N_2201,N_1444,N_1618);
or U2202 (N_2202,N_1314,N_1637);
and U2203 (N_2203,N_1670,N_1785);
and U2204 (N_2204,N_1506,N_1751);
and U2205 (N_2205,N_1557,N_1433);
or U2206 (N_2206,N_1572,N_1248);
or U2207 (N_2207,N_1495,N_1313);
and U2208 (N_2208,N_1684,N_1602);
or U2209 (N_2209,N_1694,N_1441);
nand U2210 (N_2210,N_1217,N_1225);
or U2211 (N_2211,N_1557,N_1214);
and U2212 (N_2212,N_1460,N_1377);
nor U2213 (N_2213,N_1237,N_1432);
nand U2214 (N_2214,N_1598,N_1574);
and U2215 (N_2215,N_1395,N_1709);
nor U2216 (N_2216,N_1607,N_1609);
nor U2217 (N_2217,N_1532,N_1208);
and U2218 (N_2218,N_1648,N_1799);
nand U2219 (N_2219,N_1390,N_1285);
nand U2220 (N_2220,N_1380,N_1597);
and U2221 (N_2221,N_1663,N_1670);
or U2222 (N_2222,N_1541,N_1790);
nor U2223 (N_2223,N_1303,N_1274);
or U2224 (N_2224,N_1523,N_1739);
and U2225 (N_2225,N_1273,N_1787);
nor U2226 (N_2226,N_1711,N_1521);
nor U2227 (N_2227,N_1434,N_1553);
or U2228 (N_2228,N_1723,N_1212);
nor U2229 (N_2229,N_1649,N_1593);
nand U2230 (N_2230,N_1438,N_1334);
nand U2231 (N_2231,N_1455,N_1333);
nor U2232 (N_2232,N_1578,N_1291);
nand U2233 (N_2233,N_1569,N_1433);
nor U2234 (N_2234,N_1232,N_1609);
nand U2235 (N_2235,N_1454,N_1359);
or U2236 (N_2236,N_1572,N_1216);
nor U2237 (N_2237,N_1791,N_1373);
nor U2238 (N_2238,N_1278,N_1478);
nor U2239 (N_2239,N_1350,N_1765);
nor U2240 (N_2240,N_1683,N_1412);
nor U2241 (N_2241,N_1243,N_1329);
or U2242 (N_2242,N_1271,N_1784);
nor U2243 (N_2243,N_1444,N_1620);
or U2244 (N_2244,N_1677,N_1657);
and U2245 (N_2245,N_1670,N_1233);
nand U2246 (N_2246,N_1353,N_1515);
and U2247 (N_2247,N_1650,N_1654);
nand U2248 (N_2248,N_1438,N_1253);
and U2249 (N_2249,N_1671,N_1673);
and U2250 (N_2250,N_1448,N_1341);
or U2251 (N_2251,N_1479,N_1222);
and U2252 (N_2252,N_1417,N_1722);
nor U2253 (N_2253,N_1226,N_1706);
or U2254 (N_2254,N_1732,N_1643);
or U2255 (N_2255,N_1655,N_1239);
and U2256 (N_2256,N_1367,N_1311);
and U2257 (N_2257,N_1391,N_1496);
and U2258 (N_2258,N_1428,N_1426);
nand U2259 (N_2259,N_1276,N_1583);
nand U2260 (N_2260,N_1416,N_1531);
nand U2261 (N_2261,N_1458,N_1682);
and U2262 (N_2262,N_1492,N_1488);
nor U2263 (N_2263,N_1350,N_1542);
nand U2264 (N_2264,N_1339,N_1492);
and U2265 (N_2265,N_1688,N_1462);
and U2266 (N_2266,N_1446,N_1777);
nand U2267 (N_2267,N_1654,N_1727);
and U2268 (N_2268,N_1683,N_1750);
nand U2269 (N_2269,N_1584,N_1481);
nand U2270 (N_2270,N_1757,N_1342);
or U2271 (N_2271,N_1650,N_1274);
or U2272 (N_2272,N_1362,N_1452);
or U2273 (N_2273,N_1706,N_1519);
nor U2274 (N_2274,N_1358,N_1530);
nand U2275 (N_2275,N_1310,N_1309);
and U2276 (N_2276,N_1552,N_1566);
xor U2277 (N_2277,N_1762,N_1795);
nand U2278 (N_2278,N_1293,N_1796);
and U2279 (N_2279,N_1536,N_1275);
nor U2280 (N_2280,N_1483,N_1770);
and U2281 (N_2281,N_1603,N_1406);
nor U2282 (N_2282,N_1360,N_1229);
or U2283 (N_2283,N_1305,N_1723);
or U2284 (N_2284,N_1318,N_1309);
and U2285 (N_2285,N_1337,N_1657);
and U2286 (N_2286,N_1736,N_1518);
and U2287 (N_2287,N_1423,N_1454);
and U2288 (N_2288,N_1789,N_1555);
nand U2289 (N_2289,N_1520,N_1357);
nand U2290 (N_2290,N_1526,N_1470);
or U2291 (N_2291,N_1703,N_1626);
or U2292 (N_2292,N_1799,N_1473);
or U2293 (N_2293,N_1687,N_1329);
or U2294 (N_2294,N_1619,N_1612);
or U2295 (N_2295,N_1338,N_1300);
or U2296 (N_2296,N_1287,N_1548);
nor U2297 (N_2297,N_1293,N_1787);
or U2298 (N_2298,N_1566,N_1577);
nand U2299 (N_2299,N_1684,N_1355);
and U2300 (N_2300,N_1361,N_1395);
or U2301 (N_2301,N_1332,N_1446);
nor U2302 (N_2302,N_1388,N_1444);
or U2303 (N_2303,N_1396,N_1570);
nand U2304 (N_2304,N_1616,N_1487);
and U2305 (N_2305,N_1606,N_1269);
or U2306 (N_2306,N_1205,N_1754);
xnor U2307 (N_2307,N_1386,N_1485);
nand U2308 (N_2308,N_1537,N_1755);
or U2309 (N_2309,N_1529,N_1678);
or U2310 (N_2310,N_1330,N_1354);
and U2311 (N_2311,N_1544,N_1508);
or U2312 (N_2312,N_1289,N_1438);
or U2313 (N_2313,N_1560,N_1653);
and U2314 (N_2314,N_1598,N_1491);
and U2315 (N_2315,N_1670,N_1758);
nor U2316 (N_2316,N_1377,N_1685);
nand U2317 (N_2317,N_1755,N_1610);
nand U2318 (N_2318,N_1341,N_1679);
and U2319 (N_2319,N_1562,N_1755);
or U2320 (N_2320,N_1385,N_1541);
and U2321 (N_2321,N_1530,N_1395);
and U2322 (N_2322,N_1666,N_1645);
nand U2323 (N_2323,N_1520,N_1333);
and U2324 (N_2324,N_1486,N_1225);
or U2325 (N_2325,N_1623,N_1231);
nand U2326 (N_2326,N_1422,N_1747);
nor U2327 (N_2327,N_1629,N_1765);
nand U2328 (N_2328,N_1645,N_1700);
nand U2329 (N_2329,N_1751,N_1232);
nor U2330 (N_2330,N_1316,N_1718);
nor U2331 (N_2331,N_1485,N_1694);
or U2332 (N_2332,N_1624,N_1793);
or U2333 (N_2333,N_1643,N_1438);
nor U2334 (N_2334,N_1796,N_1217);
nor U2335 (N_2335,N_1476,N_1316);
nand U2336 (N_2336,N_1610,N_1407);
or U2337 (N_2337,N_1218,N_1472);
or U2338 (N_2338,N_1355,N_1482);
or U2339 (N_2339,N_1689,N_1234);
nor U2340 (N_2340,N_1509,N_1710);
or U2341 (N_2341,N_1371,N_1666);
or U2342 (N_2342,N_1715,N_1310);
nor U2343 (N_2343,N_1447,N_1400);
and U2344 (N_2344,N_1539,N_1373);
or U2345 (N_2345,N_1392,N_1612);
and U2346 (N_2346,N_1331,N_1714);
and U2347 (N_2347,N_1471,N_1371);
or U2348 (N_2348,N_1222,N_1643);
nor U2349 (N_2349,N_1290,N_1607);
nand U2350 (N_2350,N_1377,N_1522);
nand U2351 (N_2351,N_1208,N_1708);
or U2352 (N_2352,N_1434,N_1746);
nand U2353 (N_2353,N_1344,N_1372);
and U2354 (N_2354,N_1744,N_1740);
and U2355 (N_2355,N_1755,N_1383);
and U2356 (N_2356,N_1738,N_1407);
and U2357 (N_2357,N_1568,N_1653);
or U2358 (N_2358,N_1443,N_1766);
or U2359 (N_2359,N_1489,N_1626);
or U2360 (N_2360,N_1649,N_1202);
or U2361 (N_2361,N_1335,N_1454);
and U2362 (N_2362,N_1758,N_1297);
nand U2363 (N_2363,N_1754,N_1597);
and U2364 (N_2364,N_1254,N_1382);
and U2365 (N_2365,N_1553,N_1420);
and U2366 (N_2366,N_1368,N_1319);
nor U2367 (N_2367,N_1355,N_1753);
and U2368 (N_2368,N_1751,N_1794);
and U2369 (N_2369,N_1219,N_1692);
or U2370 (N_2370,N_1614,N_1278);
nand U2371 (N_2371,N_1421,N_1239);
or U2372 (N_2372,N_1248,N_1725);
and U2373 (N_2373,N_1624,N_1791);
nand U2374 (N_2374,N_1422,N_1239);
or U2375 (N_2375,N_1671,N_1749);
nand U2376 (N_2376,N_1490,N_1245);
or U2377 (N_2377,N_1662,N_1337);
nor U2378 (N_2378,N_1692,N_1552);
and U2379 (N_2379,N_1418,N_1717);
or U2380 (N_2380,N_1275,N_1753);
and U2381 (N_2381,N_1630,N_1395);
nor U2382 (N_2382,N_1483,N_1436);
nor U2383 (N_2383,N_1695,N_1250);
or U2384 (N_2384,N_1234,N_1573);
and U2385 (N_2385,N_1533,N_1285);
nor U2386 (N_2386,N_1713,N_1456);
or U2387 (N_2387,N_1744,N_1757);
nor U2388 (N_2388,N_1740,N_1261);
nor U2389 (N_2389,N_1585,N_1436);
or U2390 (N_2390,N_1455,N_1374);
nor U2391 (N_2391,N_1404,N_1205);
and U2392 (N_2392,N_1504,N_1263);
nand U2393 (N_2393,N_1334,N_1539);
and U2394 (N_2394,N_1730,N_1555);
nor U2395 (N_2395,N_1560,N_1686);
and U2396 (N_2396,N_1567,N_1402);
nand U2397 (N_2397,N_1667,N_1770);
or U2398 (N_2398,N_1272,N_1409);
nand U2399 (N_2399,N_1719,N_1336);
nor U2400 (N_2400,N_2185,N_2017);
nand U2401 (N_2401,N_1868,N_1912);
or U2402 (N_2402,N_2339,N_2225);
nor U2403 (N_2403,N_1892,N_2381);
nor U2404 (N_2404,N_1884,N_2087);
nand U2405 (N_2405,N_2078,N_2263);
nor U2406 (N_2406,N_2049,N_2242);
nand U2407 (N_2407,N_2142,N_1921);
nor U2408 (N_2408,N_2134,N_2260);
nor U2409 (N_2409,N_2300,N_2039);
nand U2410 (N_2410,N_1925,N_1904);
and U2411 (N_2411,N_2181,N_2131);
or U2412 (N_2412,N_1991,N_1990);
nand U2413 (N_2413,N_2344,N_1929);
nand U2414 (N_2414,N_2203,N_2050);
or U2415 (N_2415,N_2084,N_2335);
and U2416 (N_2416,N_2325,N_2223);
or U2417 (N_2417,N_1997,N_1807);
or U2418 (N_2418,N_2005,N_2371);
nand U2419 (N_2419,N_2199,N_2194);
nand U2420 (N_2420,N_2146,N_1926);
or U2421 (N_2421,N_1900,N_2316);
and U2422 (N_2422,N_1969,N_2154);
and U2423 (N_2423,N_2130,N_2269);
nor U2424 (N_2424,N_2220,N_2137);
or U2425 (N_2425,N_2274,N_1810);
nand U2426 (N_2426,N_2243,N_1883);
and U2427 (N_2427,N_2168,N_2148);
nand U2428 (N_2428,N_1945,N_2392);
or U2429 (N_2429,N_2279,N_1967);
and U2430 (N_2430,N_1861,N_1999);
nand U2431 (N_2431,N_2319,N_1872);
or U2432 (N_2432,N_2023,N_2202);
nand U2433 (N_2433,N_1869,N_2293);
and U2434 (N_2434,N_1911,N_1901);
or U2435 (N_2435,N_2015,N_2031);
nand U2436 (N_2436,N_2113,N_1812);
nor U2437 (N_2437,N_2310,N_2390);
and U2438 (N_2438,N_2121,N_2200);
nand U2439 (N_2439,N_1808,N_2327);
and U2440 (N_2440,N_1874,N_2110);
nand U2441 (N_2441,N_2256,N_1944);
and U2442 (N_2442,N_2287,N_2233);
and U2443 (N_2443,N_2045,N_2069);
nor U2444 (N_2444,N_2032,N_1855);
nor U2445 (N_2445,N_1870,N_2391);
nor U2446 (N_2446,N_1927,N_2071);
and U2447 (N_2447,N_1930,N_2103);
nand U2448 (N_2448,N_2350,N_1894);
and U2449 (N_2449,N_2234,N_2138);
and U2450 (N_2450,N_2075,N_2167);
or U2451 (N_2451,N_2240,N_2129);
nor U2452 (N_2452,N_2052,N_2324);
and U2453 (N_2453,N_2229,N_2334);
or U2454 (N_2454,N_1987,N_2021);
and U2455 (N_2455,N_1983,N_2333);
nor U2456 (N_2456,N_2192,N_2309);
and U2457 (N_2457,N_2359,N_2288);
or U2458 (N_2458,N_2383,N_2208);
nand U2459 (N_2459,N_2117,N_2216);
and U2460 (N_2460,N_1830,N_1994);
and U2461 (N_2461,N_2304,N_1972);
and U2462 (N_2462,N_1877,N_2248);
nand U2463 (N_2463,N_2090,N_2369);
nand U2464 (N_2464,N_2341,N_2160);
or U2465 (N_2465,N_1970,N_2043);
nor U2466 (N_2466,N_1956,N_2299);
nor U2467 (N_2467,N_2025,N_1837);
or U2468 (N_2468,N_1984,N_2282);
nor U2469 (N_2469,N_1862,N_2384);
or U2470 (N_2470,N_2176,N_1851);
nand U2471 (N_2471,N_2337,N_2246);
nand U2472 (N_2472,N_1922,N_2053);
nor U2473 (N_2473,N_1913,N_2056);
or U2474 (N_2474,N_2067,N_1839);
nor U2475 (N_2475,N_2089,N_1964);
or U2476 (N_2476,N_1893,N_1961);
and U2477 (N_2477,N_1801,N_2171);
nand U2478 (N_2478,N_2252,N_1988);
nand U2479 (N_2479,N_2387,N_2001);
nand U2480 (N_2480,N_2106,N_1903);
nand U2481 (N_2481,N_2258,N_1953);
and U2482 (N_2482,N_2317,N_2235);
and U2483 (N_2483,N_2169,N_2281);
and U2484 (N_2484,N_2395,N_2016);
and U2485 (N_2485,N_2128,N_1905);
nor U2486 (N_2486,N_1829,N_1958);
and U2487 (N_2487,N_1820,N_2211);
or U2488 (N_2488,N_2259,N_2266);
and U2489 (N_2489,N_2116,N_2284);
nor U2490 (N_2490,N_2152,N_1840);
nand U2491 (N_2491,N_1805,N_2217);
nand U2492 (N_2492,N_2082,N_2157);
and U2493 (N_2493,N_2012,N_1804);
nor U2494 (N_2494,N_2101,N_2081);
nor U2495 (N_2495,N_1955,N_1890);
nand U2496 (N_2496,N_1938,N_2115);
or U2497 (N_2497,N_2112,N_2096);
nand U2498 (N_2498,N_2238,N_1876);
and U2499 (N_2499,N_2253,N_2007);
nor U2500 (N_2500,N_2011,N_2014);
nand U2501 (N_2501,N_2175,N_1985);
nand U2502 (N_2502,N_2141,N_2353);
or U2503 (N_2503,N_2037,N_1935);
xor U2504 (N_2504,N_1885,N_1871);
nand U2505 (N_2505,N_1941,N_1813);
nor U2506 (N_2506,N_2074,N_2098);
nor U2507 (N_2507,N_2394,N_1942);
nor U2508 (N_2508,N_2026,N_2000);
xnor U2509 (N_2509,N_2298,N_2352);
and U2510 (N_2510,N_1924,N_2262);
nor U2511 (N_2511,N_1838,N_1828);
nor U2512 (N_2512,N_2318,N_1814);
nor U2513 (N_2513,N_2048,N_1850);
and U2514 (N_2514,N_2356,N_2190);
nand U2515 (N_2515,N_1873,N_2374);
nand U2516 (N_2516,N_2255,N_1859);
and U2517 (N_2517,N_2268,N_2330);
nor U2518 (N_2518,N_2212,N_2061);
and U2519 (N_2519,N_1986,N_1943);
or U2520 (N_2520,N_1880,N_2083);
nand U2521 (N_2521,N_2351,N_2094);
nor U2522 (N_2522,N_2024,N_2245);
and U2523 (N_2523,N_1923,N_2188);
nor U2524 (N_2524,N_2206,N_2241);
nand U2525 (N_2525,N_2177,N_2095);
nor U2526 (N_2526,N_2119,N_2178);
nor U2527 (N_2527,N_1879,N_2380);
and U2528 (N_2528,N_2354,N_1980);
nand U2529 (N_2529,N_1852,N_2349);
or U2530 (N_2530,N_1858,N_2251);
nor U2531 (N_2531,N_2174,N_2120);
or U2532 (N_2532,N_1906,N_1845);
nand U2533 (N_2533,N_1898,N_2261);
nand U2534 (N_2534,N_2063,N_2044);
and U2535 (N_2535,N_2099,N_2313);
and U2536 (N_2536,N_2280,N_1908);
nor U2537 (N_2537,N_2179,N_2046);
and U2538 (N_2538,N_1975,N_2204);
nand U2539 (N_2539,N_2301,N_2382);
and U2540 (N_2540,N_1878,N_2302);
nor U2541 (N_2541,N_2158,N_1976);
or U2542 (N_2542,N_1896,N_1940);
nand U2543 (N_2543,N_2197,N_2165);
nand U2544 (N_2544,N_1907,N_1881);
and U2545 (N_2545,N_1996,N_1952);
nand U2546 (N_2546,N_2150,N_1947);
or U2547 (N_2547,N_1819,N_2227);
and U2548 (N_2548,N_2038,N_2109);
nand U2549 (N_2549,N_1933,N_2355);
and U2550 (N_2550,N_1950,N_2265);
or U2551 (N_2551,N_1843,N_2172);
nor U2552 (N_2552,N_2385,N_1915);
nand U2553 (N_2553,N_2195,N_2221);
nor U2554 (N_2554,N_1959,N_2273);
nor U2555 (N_2555,N_1979,N_1914);
nor U2556 (N_2556,N_2164,N_2034);
nor U2557 (N_2557,N_2062,N_2140);
nor U2558 (N_2558,N_2139,N_1800);
and U2559 (N_2559,N_2186,N_1966);
or U2560 (N_2560,N_1854,N_2207);
or U2561 (N_2561,N_1836,N_2159);
nand U2562 (N_2562,N_2232,N_1887);
nor U2563 (N_2563,N_2022,N_2010);
or U2564 (N_2564,N_2149,N_2076);
nand U2565 (N_2565,N_2323,N_1974);
nand U2566 (N_2566,N_2289,N_2118);
nor U2567 (N_2567,N_1866,N_2272);
nand U2568 (N_2568,N_2342,N_2183);
nand U2569 (N_2569,N_2198,N_1889);
nand U2570 (N_2570,N_2064,N_2315);
or U2571 (N_2571,N_1834,N_2239);
nand U2572 (N_2572,N_1835,N_1897);
or U2573 (N_2573,N_2080,N_1960);
or U2574 (N_2574,N_2283,N_2060);
nor U2575 (N_2575,N_2013,N_1917);
nor U2576 (N_2576,N_1936,N_1957);
nand U2577 (N_2577,N_2018,N_1916);
nand U2578 (N_2578,N_2377,N_2123);
nand U2579 (N_2579,N_2393,N_2189);
nand U2580 (N_2580,N_1977,N_1848);
and U2581 (N_2581,N_2028,N_2147);
and U2582 (N_2582,N_2218,N_2182);
nand U2583 (N_2583,N_1846,N_2161);
nand U2584 (N_2584,N_2366,N_1995);
and U2585 (N_2585,N_1899,N_1932);
nor U2586 (N_2586,N_1882,N_1832);
nand U2587 (N_2587,N_2041,N_2294);
nor U2588 (N_2588,N_2143,N_2162);
and U2589 (N_2589,N_2378,N_2308);
and U2590 (N_2590,N_1891,N_2136);
and U2591 (N_2591,N_1920,N_2077);
and U2592 (N_2592,N_1946,N_2020);
nor U2593 (N_2593,N_1856,N_2357);
and U2594 (N_2594,N_2275,N_1816);
nor U2595 (N_2595,N_2321,N_2055);
and U2596 (N_2596,N_2320,N_1909);
or U2597 (N_2597,N_1827,N_2187);
and U2598 (N_2598,N_1824,N_1826);
or U2599 (N_2599,N_2073,N_1841);
nor U2600 (N_2600,N_2367,N_2271);
and U2601 (N_2601,N_2003,N_1817);
and U2602 (N_2602,N_1803,N_2388);
nand U2603 (N_2603,N_2244,N_1963);
nor U2604 (N_2604,N_2398,N_2085);
nor U2605 (N_2605,N_2004,N_1811);
or U2606 (N_2606,N_2155,N_2151);
or U2607 (N_2607,N_2270,N_2219);
and U2608 (N_2608,N_2305,N_2329);
or U2609 (N_2609,N_2311,N_2047);
or U2610 (N_2610,N_2086,N_2191);
and U2611 (N_2611,N_2336,N_2346);
nor U2612 (N_2612,N_2114,N_2322);
nor U2613 (N_2613,N_2250,N_2224);
nor U2614 (N_2614,N_1982,N_1981);
and U2615 (N_2615,N_2286,N_2009);
and U2616 (N_2616,N_2226,N_2370);
or U2617 (N_2617,N_2328,N_2209);
and U2618 (N_2618,N_2030,N_2331);
nand U2619 (N_2619,N_2205,N_2295);
xor U2620 (N_2620,N_2306,N_1934);
nand U2621 (N_2621,N_2111,N_1998);
nand U2622 (N_2622,N_1978,N_2173);
nand U2623 (N_2623,N_2042,N_2332);
nor U2624 (N_2624,N_2285,N_1989);
nor U2625 (N_2625,N_2264,N_1886);
nand U2626 (N_2626,N_2372,N_1919);
or U2627 (N_2627,N_2057,N_1949);
and U2628 (N_2628,N_2291,N_1962);
or U2629 (N_2629,N_2163,N_2122);
or U2630 (N_2630,N_2124,N_2035);
and U2631 (N_2631,N_1831,N_2375);
nand U2632 (N_2632,N_2249,N_2180);
and U2633 (N_2633,N_2133,N_2214);
or U2634 (N_2634,N_2326,N_2247);
nand U2635 (N_2635,N_2236,N_2365);
or U2636 (N_2636,N_2126,N_2303);
or U2637 (N_2637,N_2193,N_1888);
nor U2638 (N_2638,N_1895,N_2312);
nand U2639 (N_2639,N_2364,N_2125);
and U2640 (N_2640,N_2100,N_2058);
nand U2641 (N_2641,N_2093,N_1860);
nand U2642 (N_2642,N_2145,N_2362);
nand U2643 (N_2643,N_1993,N_2002);
or U2644 (N_2644,N_1928,N_2292);
nor U2645 (N_2645,N_2033,N_2215);
and U2646 (N_2646,N_2153,N_1954);
nand U2647 (N_2647,N_2059,N_2314);
and U2648 (N_2648,N_2396,N_2347);
nor U2649 (N_2649,N_1802,N_1821);
or U2650 (N_2650,N_2029,N_2278);
nor U2651 (N_2651,N_2104,N_1823);
nand U2652 (N_2652,N_2135,N_2105);
nand U2653 (N_2653,N_1809,N_2358);
and U2654 (N_2654,N_1931,N_1992);
or U2655 (N_2655,N_2257,N_2213);
nor U2656 (N_2656,N_1825,N_2231);
or U2657 (N_2657,N_1849,N_1973);
or U2658 (N_2658,N_1806,N_1937);
nand U2659 (N_2659,N_2373,N_2019);
nand U2660 (N_2660,N_2170,N_2222);
nor U2661 (N_2661,N_1865,N_2051);
or U2662 (N_2662,N_2210,N_1857);
and U2663 (N_2663,N_1853,N_2376);
or U2664 (N_2664,N_2127,N_1842);
and U2665 (N_2665,N_2184,N_1818);
nand U2666 (N_2666,N_2068,N_2360);
nor U2667 (N_2667,N_2348,N_2036);
and U2668 (N_2668,N_2361,N_2196);
nor U2669 (N_2669,N_2254,N_1918);
and U2670 (N_2670,N_2363,N_2072);
nand U2671 (N_2671,N_2054,N_1910);
nand U2672 (N_2672,N_1863,N_2144);
and U2673 (N_2673,N_2070,N_1951);
nand U2674 (N_2674,N_1965,N_2065);
or U2675 (N_2675,N_2040,N_2156);
and U2676 (N_2676,N_2267,N_2338);
xor U2677 (N_2677,N_1948,N_2340);
or U2678 (N_2678,N_2108,N_1968);
or U2679 (N_2679,N_2102,N_2296);
nand U2680 (N_2680,N_2088,N_2079);
nor U2681 (N_2681,N_2066,N_2343);
nor U2682 (N_2682,N_2091,N_2397);
or U2683 (N_2683,N_2201,N_1844);
nand U2684 (N_2684,N_2008,N_1822);
nand U2685 (N_2685,N_1864,N_2277);
and U2686 (N_2686,N_2092,N_1847);
and U2687 (N_2687,N_1902,N_2228);
xor U2688 (N_2688,N_2166,N_2386);
or U2689 (N_2689,N_2027,N_2389);
and U2690 (N_2690,N_2307,N_1833);
or U2691 (N_2691,N_1867,N_2368);
or U2692 (N_2692,N_2399,N_1939);
and U2693 (N_2693,N_2276,N_2297);
nor U2694 (N_2694,N_2132,N_2107);
and U2695 (N_2695,N_2237,N_1815);
nor U2696 (N_2696,N_2379,N_2230);
nand U2697 (N_2697,N_1875,N_2290);
or U2698 (N_2698,N_2097,N_2345);
nand U2699 (N_2699,N_2006,N_1971);
nor U2700 (N_2700,N_1830,N_2339);
nor U2701 (N_2701,N_1883,N_1888);
and U2702 (N_2702,N_1970,N_2321);
nor U2703 (N_2703,N_1836,N_2071);
and U2704 (N_2704,N_2075,N_2242);
or U2705 (N_2705,N_2353,N_2377);
and U2706 (N_2706,N_1831,N_2285);
or U2707 (N_2707,N_1953,N_2091);
or U2708 (N_2708,N_2238,N_1802);
or U2709 (N_2709,N_1947,N_1864);
and U2710 (N_2710,N_1968,N_1977);
and U2711 (N_2711,N_2285,N_1837);
nor U2712 (N_2712,N_2131,N_2387);
nor U2713 (N_2713,N_2372,N_2262);
nor U2714 (N_2714,N_2010,N_1938);
nor U2715 (N_2715,N_1940,N_2013);
nand U2716 (N_2716,N_1871,N_2254);
and U2717 (N_2717,N_2158,N_1830);
nor U2718 (N_2718,N_2215,N_1987);
and U2719 (N_2719,N_1897,N_1903);
or U2720 (N_2720,N_1947,N_1907);
nor U2721 (N_2721,N_1843,N_1845);
nand U2722 (N_2722,N_1840,N_2298);
nand U2723 (N_2723,N_2321,N_2389);
nor U2724 (N_2724,N_2335,N_2145);
and U2725 (N_2725,N_1952,N_2399);
nor U2726 (N_2726,N_1864,N_1921);
and U2727 (N_2727,N_2141,N_2181);
and U2728 (N_2728,N_1822,N_1990);
and U2729 (N_2729,N_2316,N_2399);
and U2730 (N_2730,N_1830,N_1923);
nor U2731 (N_2731,N_2000,N_2025);
or U2732 (N_2732,N_2274,N_2171);
nand U2733 (N_2733,N_1968,N_1903);
nor U2734 (N_2734,N_1958,N_2011);
or U2735 (N_2735,N_2384,N_2318);
or U2736 (N_2736,N_2066,N_1804);
or U2737 (N_2737,N_2314,N_2367);
or U2738 (N_2738,N_2017,N_2199);
nand U2739 (N_2739,N_2378,N_2342);
nor U2740 (N_2740,N_2217,N_2301);
nor U2741 (N_2741,N_2243,N_2035);
and U2742 (N_2742,N_2004,N_1933);
nand U2743 (N_2743,N_1949,N_2218);
and U2744 (N_2744,N_1869,N_1859);
nor U2745 (N_2745,N_2028,N_1912);
or U2746 (N_2746,N_2353,N_1964);
nor U2747 (N_2747,N_2286,N_2203);
nor U2748 (N_2748,N_2178,N_2325);
nor U2749 (N_2749,N_2140,N_2049);
nor U2750 (N_2750,N_2207,N_2225);
nand U2751 (N_2751,N_2081,N_1988);
or U2752 (N_2752,N_1896,N_1951);
and U2753 (N_2753,N_2162,N_2058);
nor U2754 (N_2754,N_2216,N_2037);
or U2755 (N_2755,N_2319,N_2147);
and U2756 (N_2756,N_2361,N_2044);
nor U2757 (N_2757,N_2284,N_2178);
nor U2758 (N_2758,N_1819,N_2279);
nand U2759 (N_2759,N_2108,N_1982);
nor U2760 (N_2760,N_2053,N_2327);
nor U2761 (N_2761,N_2303,N_2054);
and U2762 (N_2762,N_2151,N_1936);
nor U2763 (N_2763,N_2376,N_2185);
or U2764 (N_2764,N_1985,N_2361);
or U2765 (N_2765,N_2048,N_1976);
or U2766 (N_2766,N_2300,N_2383);
or U2767 (N_2767,N_2167,N_1989);
and U2768 (N_2768,N_2018,N_2171);
nand U2769 (N_2769,N_2033,N_1974);
nand U2770 (N_2770,N_2160,N_1933);
nand U2771 (N_2771,N_2240,N_2022);
nor U2772 (N_2772,N_1861,N_2382);
and U2773 (N_2773,N_2329,N_2010);
and U2774 (N_2774,N_1955,N_1814);
and U2775 (N_2775,N_1858,N_2344);
or U2776 (N_2776,N_1888,N_2072);
or U2777 (N_2777,N_2069,N_1948);
xor U2778 (N_2778,N_2228,N_1978);
nor U2779 (N_2779,N_2250,N_2168);
and U2780 (N_2780,N_1909,N_2273);
nand U2781 (N_2781,N_1830,N_1894);
nand U2782 (N_2782,N_2191,N_2231);
and U2783 (N_2783,N_2059,N_1984);
nor U2784 (N_2784,N_1968,N_2231);
or U2785 (N_2785,N_2207,N_1975);
or U2786 (N_2786,N_2311,N_2005);
or U2787 (N_2787,N_2338,N_2279);
nor U2788 (N_2788,N_2220,N_2148);
or U2789 (N_2789,N_2092,N_2234);
nand U2790 (N_2790,N_2389,N_1811);
nand U2791 (N_2791,N_2393,N_1928);
nor U2792 (N_2792,N_1853,N_2149);
nand U2793 (N_2793,N_2187,N_1872);
or U2794 (N_2794,N_2370,N_2297);
nor U2795 (N_2795,N_1816,N_2308);
and U2796 (N_2796,N_1985,N_2307);
nor U2797 (N_2797,N_1821,N_2068);
and U2798 (N_2798,N_2005,N_2054);
or U2799 (N_2799,N_1831,N_1869);
nand U2800 (N_2800,N_1853,N_2327);
nand U2801 (N_2801,N_2151,N_2042);
or U2802 (N_2802,N_1988,N_1962);
and U2803 (N_2803,N_2309,N_1801);
nand U2804 (N_2804,N_2273,N_2399);
or U2805 (N_2805,N_2006,N_1801);
and U2806 (N_2806,N_2034,N_2181);
or U2807 (N_2807,N_2203,N_2095);
nor U2808 (N_2808,N_1970,N_2085);
nand U2809 (N_2809,N_2163,N_2052);
and U2810 (N_2810,N_1828,N_2140);
nand U2811 (N_2811,N_2282,N_2369);
and U2812 (N_2812,N_2232,N_2292);
nand U2813 (N_2813,N_2241,N_2231);
nor U2814 (N_2814,N_2342,N_2217);
nand U2815 (N_2815,N_2315,N_1906);
and U2816 (N_2816,N_2180,N_2265);
nand U2817 (N_2817,N_1890,N_2349);
nor U2818 (N_2818,N_2177,N_1961);
and U2819 (N_2819,N_1804,N_1984);
and U2820 (N_2820,N_1822,N_1828);
and U2821 (N_2821,N_2010,N_2024);
or U2822 (N_2822,N_2055,N_1872);
and U2823 (N_2823,N_2318,N_2046);
nor U2824 (N_2824,N_2389,N_2170);
and U2825 (N_2825,N_1820,N_2147);
xor U2826 (N_2826,N_2263,N_2355);
nor U2827 (N_2827,N_2393,N_1939);
or U2828 (N_2828,N_1916,N_1910);
nand U2829 (N_2829,N_1940,N_2367);
nor U2830 (N_2830,N_1854,N_1877);
nor U2831 (N_2831,N_1929,N_2134);
nor U2832 (N_2832,N_2002,N_2017);
and U2833 (N_2833,N_2036,N_2137);
or U2834 (N_2834,N_1832,N_1939);
nand U2835 (N_2835,N_2100,N_2305);
or U2836 (N_2836,N_2376,N_2336);
and U2837 (N_2837,N_2071,N_2154);
or U2838 (N_2838,N_2324,N_2225);
nor U2839 (N_2839,N_2397,N_1819);
or U2840 (N_2840,N_1849,N_2082);
or U2841 (N_2841,N_1868,N_2304);
nand U2842 (N_2842,N_1809,N_2203);
or U2843 (N_2843,N_2170,N_1857);
nand U2844 (N_2844,N_2323,N_2191);
nand U2845 (N_2845,N_2220,N_2347);
and U2846 (N_2846,N_2269,N_1910);
or U2847 (N_2847,N_1894,N_2104);
and U2848 (N_2848,N_2135,N_1913);
nor U2849 (N_2849,N_1808,N_2310);
and U2850 (N_2850,N_2066,N_1972);
nor U2851 (N_2851,N_1956,N_2058);
or U2852 (N_2852,N_2021,N_2389);
or U2853 (N_2853,N_2146,N_2082);
nor U2854 (N_2854,N_2200,N_1808);
nor U2855 (N_2855,N_1943,N_2208);
and U2856 (N_2856,N_2227,N_1800);
nand U2857 (N_2857,N_2197,N_2110);
nand U2858 (N_2858,N_1896,N_2016);
and U2859 (N_2859,N_1995,N_2378);
nand U2860 (N_2860,N_2124,N_2020);
or U2861 (N_2861,N_2256,N_1883);
nor U2862 (N_2862,N_2321,N_1828);
and U2863 (N_2863,N_1930,N_2192);
and U2864 (N_2864,N_2176,N_2056);
nor U2865 (N_2865,N_2014,N_2007);
and U2866 (N_2866,N_2358,N_1831);
nand U2867 (N_2867,N_2327,N_2085);
nor U2868 (N_2868,N_2174,N_2329);
and U2869 (N_2869,N_2197,N_1844);
and U2870 (N_2870,N_2076,N_2374);
nor U2871 (N_2871,N_1901,N_2112);
or U2872 (N_2872,N_1998,N_2106);
nand U2873 (N_2873,N_2393,N_2138);
nor U2874 (N_2874,N_2121,N_2038);
or U2875 (N_2875,N_1814,N_2273);
and U2876 (N_2876,N_2095,N_1855);
and U2877 (N_2877,N_2044,N_1842);
nor U2878 (N_2878,N_2374,N_2274);
and U2879 (N_2879,N_2081,N_2231);
nor U2880 (N_2880,N_2042,N_2210);
or U2881 (N_2881,N_2115,N_2274);
and U2882 (N_2882,N_2075,N_2064);
nand U2883 (N_2883,N_2280,N_2059);
nand U2884 (N_2884,N_2238,N_2270);
and U2885 (N_2885,N_2042,N_2338);
nor U2886 (N_2886,N_2373,N_1909);
nor U2887 (N_2887,N_1941,N_1940);
or U2888 (N_2888,N_1810,N_2038);
or U2889 (N_2889,N_1935,N_2222);
or U2890 (N_2890,N_2102,N_2381);
or U2891 (N_2891,N_1999,N_2177);
nand U2892 (N_2892,N_2200,N_2244);
nand U2893 (N_2893,N_2279,N_1916);
nand U2894 (N_2894,N_1859,N_2307);
or U2895 (N_2895,N_2389,N_2248);
and U2896 (N_2896,N_1943,N_2355);
nand U2897 (N_2897,N_2061,N_2196);
and U2898 (N_2898,N_2331,N_1812);
and U2899 (N_2899,N_2173,N_2135);
or U2900 (N_2900,N_2360,N_2333);
and U2901 (N_2901,N_2160,N_2281);
and U2902 (N_2902,N_2374,N_2257);
and U2903 (N_2903,N_2291,N_1833);
nor U2904 (N_2904,N_2221,N_1962);
nand U2905 (N_2905,N_2130,N_2315);
or U2906 (N_2906,N_1850,N_1959);
and U2907 (N_2907,N_1968,N_2041);
nor U2908 (N_2908,N_1880,N_2362);
or U2909 (N_2909,N_2261,N_2024);
nor U2910 (N_2910,N_2114,N_1820);
nor U2911 (N_2911,N_2117,N_2222);
and U2912 (N_2912,N_1801,N_1901);
nand U2913 (N_2913,N_2324,N_2113);
or U2914 (N_2914,N_1883,N_1950);
nand U2915 (N_2915,N_2109,N_2209);
and U2916 (N_2916,N_2101,N_2148);
and U2917 (N_2917,N_2338,N_1895);
nand U2918 (N_2918,N_2073,N_2372);
nor U2919 (N_2919,N_2046,N_1908);
nand U2920 (N_2920,N_2236,N_2097);
or U2921 (N_2921,N_2017,N_2395);
nand U2922 (N_2922,N_1894,N_2089);
or U2923 (N_2923,N_1968,N_2110);
nand U2924 (N_2924,N_2266,N_2247);
or U2925 (N_2925,N_2067,N_2293);
xor U2926 (N_2926,N_1931,N_1814);
nor U2927 (N_2927,N_2335,N_1858);
nor U2928 (N_2928,N_1874,N_2104);
nor U2929 (N_2929,N_1898,N_1856);
and U2930 (N_2930,N_2187,N_1884);
or U2931 (N_2931,N_1994,N_1817);
or U2932 (N_2932,N_2020,N_2209);
nand U2933 (N_2933,N_2351,N_2286);
and U2934 (N_2934,N_2051,N_1936);
and U2935 (N_2935,N_1814,N_2101);
and U2936 (N_2936,N_2358,N_2269);
or U2937 (N_2937,N_2106,N_2381);
nor U2938 (N_2938,N_2253,N_2371);
and U2939 (N_2939,N_1904,N_2212);
nand U2940 (N_2940,N_1957,N_1926);
or U2941 (N_2941,N_2321,N_2379);
nand U2942 (N_2942,N_2318,N_1937);
nand U2943 (N_2943,N_2059,N_2271);
nand U2944 (N_2944,N_1990,N_1850);
xor U2945 (N_2945,N_2079,N_2159);
and U2946 (N_2946,N_2022,N_2069);
nand U2947 (N_2947,N_1852,N_2017);
nor U2948 (N_2948,N_2313,N_1967);
nor U2949 (N_2949,N_2138,N_2268);
nand U2950 (N_2950,N_2053,N_1960);
and U2951 (N_2951,N_1850,N_1885);
and U2952 (N_2952,N_2209,N_2063);
nand U2953 (N_2953,N_2168,N_2270);
nor U2954 (N_2954,N_1841,N_2048);
nor U2955 (N_2955,N_2396,N_2200);
nand U2956 (N_2956,N_2115,N_2081);
nand U2957 (N_2957,N_1958,N_2146);
or U2958 (N_2958,N_2012,N_2137);
or U2959 (N_2959,N_1887,N_2012);
and U2960 (N_2960,N_2225,N_2197);
or U2961 (N_2961,N_2271,N_2243);
or U2962 (N_2962,N_2104,N_1942);
nor U2963 (N_2963,N_2363,N_1865);
nor U2964 (N_2964,N_2349,N_1895);
or U2965 (N_2965,N_2223,N_2149);
nor U2966 (N_2966,N_2341,N_2233);
or U2967 (N_2967,N_1902,N_2317);
nand U2968 (N_2968,N_2379,N_1839);
nand U2969 (N_2969,N_2236,N_2132);
nand U2970 (N_2970,N_2284,N_2283);
nand U2971 (N_2971,N_2043,N_2037);
nand U2972 (N_2972,N_1871,N_2169);
and U2973 (N_2973,N_1839,N_2214);
or U2974 (N_2974,N_1808,N_2353);
nand U2975 (N_2975,N_1808,N_2140);
nor U2976 (N_2976,N_2293,N_2239);
or U2977 (N_2977,N_2229,N_2120);
or U2978 (N_2978,N_2211,N_2161);
nand U2979 (N_2979,N_1948,N_1855);
nor U2980 (N_2980,N_1981,N_2160);
or U2981 (N_2981,N_2276,N_1832);
nor U2982 (N_2982,N_1973,N_2017);
and U2983 (N_2983,N_2387,N_1802);
and U2984 (N_2984,N_2319,N_1830);
or U2985 (N_2985,N_2324,N_1821);
nor U2986 (N_2986,N_1964,N_1998);
nand U2987 (N_2987,N_2176,N_2154);
nor U2988 (N_2988,N_2100,N_2072);
and U2989 (N_2989,N_1837,N_2238);
nor U2990 (N_2990,N_2117,N_1849);
nor U2991 (N_2991,N_2318,N_1838);
and U2992 (N_2992,N_2375,N_1858);
xor U2993 (N_2993,N_2339,N_2236);
nand U2994 (N_2994,N_1991,N_2251);
nand U2995 (N_2995,N_2104,N_2050);
and U2996 (N_2996,N_2352,N_2388);
or U2997 (N_2997,N_2267,N_1832);
and U2998 (N_2998,N_1897,N_2389);
or U2999 (N_2999,N_2387,N_1845);
or UO_0 (O_0,N_2413,N_2704);
nand UO_1 (O_1,N_2626,N_2538);
nand UO_2 (O_2,N_2761,N_2541);
nor UO_3 (O_3,N_2673,N_2443);
and UO_4 (O_4,N_2890,N_2560);
nand UO_5 (O_5,N_2858,N_2803);
and UO_6 (O_6,N_2986,N_2598);
and UO_7 (O_7,N_2883,N_2435);
nand UO_8 (O_8,N_2765,N_2719);
and UO_9 (O_9,N_2874,N_2762);
nand UO_10 (O_10,N_2914,N_2663);
nand UO_11 (O_11,N_2679,N_2808);
and UO_12 (O_12,N_2984,N_2901);
nand UO_13 (O_13,N_2612,N_2463);
and UO_14 (O_14,N_2749,N_2603);
and UO_15 (O_15,N_2714,N_2742);
or UO_16 (O_16,N_2527,N_2817);
or UO_17 (O_17,N_2718,N_2850);
nand UO_18 (O_18,N_2716,N_2823);
nand UO_19 (O_19,N_2546,N_2720);
nor UO_20 (O_20,N_2552,N_2886);
nor UO_21 (O_21,N_2620,N_2834);
or UO_22 (O_22,N_2832,N_2793);
or UO_23 (O_23,N_2456,N_2508);
nor UO_24 (O_24,N_2977,N_2934);
nand UO_25 (O_25,N_2573,N_2558);
nand UO_26 (O_26,N_2807,N_2861);
or UO_27 (O_27,N_2630,N_2657);
and UO_28 (O_28,N_2494,N_2465);
nor UO_29 (O_29,N_2869,N_2493);
nor UO_30 (O_30,N_2650,N_2523);
and UO_31 (O_31,N_2550,N_2540);
nand UO_32 (O_32,N_2997,N_2422);
and UO_33 (O_33,N_2661,N_2894);
and UO_34 (O_34,N_2819,N_2577);
nand UO_35 (O_35,N_2642,N_2790);
nor UO_36 (O_36,N_2702,N_2649);
nor UO_37 (O_37,N_2458,N_2453);
nor UO_38 (O_38,N_2470,N_2543);
nand UO_39 (O_39,N_2654,N_2646);
or UO_40 (O_40,N_2431,N_2919);
nand UO_41 (O_41,N_2963,N_2755);
nand UO_42 (O_42,N_2833,N_2467);
nor UO_43 (O_43,N_2747,N_2684);
nor UO_44 (O_44,N_2644,N_2617);
nor UO_45 (O_45,N_2452,N_2896);
and UO_46 (O_46,N_2824,N_2722);
nand UO_47 (O_47,N_2578,N_2600);
or UO_48 (O_48,N_2821,N_2407);
nand UO_49 (O_49,N_2582,N_2961);
or UO_50 (O_50,N_2708,N_2763);
nand UO_51 (O_51,N_2619,N_2954);
nand UO_52 (O_52,N_2591,N_2444);
and UO_53 (O_53,N_2579,N_2802);
or UO_54 (O_54,N_2660,N_2903);
and UO_55 (O_55,N_2695,N_2962);
and UO_56 (O_56,N_2408,N_2696);
nand UO_57 (O_57,N_2733,N_2760);
xnor UO_58 (O_58,N_2454,N_2857);
nor UO_59 (O_59,N_2585,N_2417);
and UO_60 (O_60,N_2907,N_2884);
nor UO_61 (O_61,N_2736,N_2643);
or UO_62 (O_62,N_2952,N_2809);
nand UO_63 (O_63,N_2621,N_2932);
nand UO_64 (O_64,N_2451,N_2865);
nand UO_65 (O_65,N_2780,N_2420);
nand UO_66 (O_66,N_2876,N_2416);
nor UO_67 (O_67,N_2670,N_2516);
or UO_68 (O_68,N_2766,N_2640);
and UO_69 (O_69,N_2924,N_2918);
nand UO_70 (O_70,N_2521,N_2575);
or UO_71 (O_71,N_2860,N_2474);
and UO_72 (O_72,N_2949,N_2553);
and UO_73 (O_73,N_2625,N_2993);
nand UO_74 (O_74,N_2783,N_2814);
and UO_75 (O_75,N_2629,N_2837);
nor UO_76 (O_76,N_2647,N_2592);
nor UO_77 (O_77,N_2767,N_2801);
nor UO_78 (O_78,N_2912,N_2426);
or UO_79 (O_79,N_2948,N_2735);
nand UO_80 (O_80,N_2715,N_2922);
nor UO_81 (O_81,N_2485,N_2728);
nor UO_82 (O_82,N_2830,N_2496);
and UO_83 (O_83,N_2844,N_2539);
nor UO_84 (O_84,N_2439,N_2666);
or UO_85 (O_85,N_2622,N_2882);
nand UO_86 (O_86,N_2723,N_2786);
nor UO_87 (O_87,N_2991,N_2489);
and UO_88 (O_88,N_2522,N_2531);
or UO_89 (O_89,N_2935,N_2881);
nand UO_90 (O_90,N_2812,N_2528);
or UO_91 (O_91,N_2569,N_2771);
nor UO_92 (O_92,N_2532,N_2816);
or UO_93 (O_93,N_2820,N_2676);
nor UO_94 (O_94,N_2460,N_2423);
and UO_95 (O_95,N_2772,N_2965);
nor UO_96 (O_96,N_2587,N_2609);
or UO_97 (O_97,N_2478,N_2847);
nor UO_98 (O_98,N_2951,N_2811);
nand UO_99 (O_99,N_2871,N_2841);
and UO_100 (O_100,N_2893,N_2913);
nor UO_101 (O_101,N_2976,N_2504);
and UO_102 (O_102,N_2978,N_2506);
nor UO_103 (O_103,N_2971,N_2549);
nand UO_104 (O_104,N_2499,N_2992);
nor UO_105 (O_105,N_2983,N_2851);
and UO_106 (O_106,N_2655,N_2581);
or UO_107 (O_107,N_2799,N_2764);
xor UO_108 (O_108,N_2955,N_2511);
or UO_109 (O_109,N_2745,N_2729);
nor UO_110 (O_110,N_2623,N_2967);
or UO_111 (O_111,N_2905,N_2996);
nor UO_112 (O_112,N_2953,N_2939);
or UO_113 (O_113,N_2966,N_2678);
and UO_114 (O_114,N_2826,N_2639);
nor UO_115 (O_115,N_2503,N_2878);
or UO_116 (O_116,N_2746,N_2475);
and UO_117 (O_117,N_2594,N_2481);
and UO_118 (O_118,N_2477,N_2872);
and UO_119 (O_119,N_2942,N_2572);
and UO_120 (O_120,N_2839,N_2712);
nor UO_121 (O_121,N_2792,N_2958);
nor UO_122 (O_122,N_2611,N_2672);
nand UO_123 (O_123,N_2887,N_2694);
and UO_124 (O_124,N_2713,N_2662);
and UO_125 (O_125,N_2667,N_2936);
nand UO_126 (O_126,N_2748,N_2605);
nand UO_127 (O_127,N_2975,N_2599);
or UO_128 (O_128,N_2513,N_2469);
nor UO_129 (O_129,N_2681,N_2664);
and UO_130 (O_130,N_2900,N_2852);
and UO_131 (O_131,N_2525,N_2656);
nor UO_132 (O_132,N_2544,N_2437);
or UO_133 (O_133,N_2597,N_2788);
or UO_134 (O_134,N_2425,N_2777);
nor UO_135 (O_135,N_2491,N_2744);
or UO_136 (O_136,N_2999,N_2926);
nand UO_137 (O_137,N_2888,N_2947);
or UO_138 (O_138,N_2668,N_2682);
nor UO_139 (O_139,N_2979,N_2510);
or UO_140 (O_140,N_2449,N_2409);
nand UO_141 (O_141,N_2432,N_2574);
nand UO_142 (O_142,N_2536,N_2698);
nor UO_143 (O_143,N_2638,N_2968);
or UO_144 (O_144,N_2464,N_2957);
or UO_145 (O_145,N_2933,N_2985);
or UO_146 (O_146,N_2628,N_2879);
or UO_147 (O_147,N_2427,N_2904);
or UO_148 (O_148,N_2652,N_2709);
nor UO_149 (O_149,N_2806,N_2734);
or UO_150 (O_150,N_2800,N_2910);
nor UO_151 (O_151,N_2921,N_2773);
or UO_152 (O_152,N_2429,N_2956);
or UO_153 (O_153,N_2419,N_2756);
nor UO_154 (O_154,N_2457,N_2885);
xnor UO_155 (O_155,N_2778,N_2498);
and UO_156 (O_156,N_2891,N_2805);
or UO_157 (O_157,N_2862,N_2835);
nand UO_158 (O_158,N_2868,N_2653);
or UO_159 (O_159,N_2845,N_2468);
or UO_160 (O_160,N_2774,N_2683);
and UO_161 (O_161,N_2873,N_2534);
and UO_162 (O_162,N_2970,N_2787);
or UO_163 (O_163,N_2796,N_2563);
nand UO_164 (O_164,N_2405,N_2974);
and UO_165 (O_165,N_2758,N_2836);
or UO_166 (O_166,N_2909,N_2737);
and UO_167 (O_167,N_2524,N_2688);
nand UO_168 (O_168,N_2483,N_2512);
nor UO_169 (O_169,N_2410,N_2635);
nor UO_170 (O_170,N_2631,N_2404);
nor UO_171 (O_171,N_2440,N_2486);
or UO_172 (O_172,N_2789,N_2840);
nor UO_173 (O_173,N_2677,N_2559);
and UO_174 (O_174,N_2593,N_2495);
or UO_175 (O_175,N_2557,N_2665);
or UO_176 (O_176,N_2509,N_2445);
nor UO_177 (O_177,N_2870,N_2795);
nor UO_178 (O_178,N_2776,N_2717);
nor UO_179 (O_179,N_2810,N_2436);
nor UO_180 (O_180,N_2699,N_2990);
nor UO_181 (O_181,N_2945,N_2401);
nor UO_182 (O_182,N_2941,N_2438);
nand UO_183 (O_183,N_2691,N_2892);
and UO_184 (O_184,N_2447,N_2595);
nor UO_185 (O_185,N_2428,N_2406);
and UO_186 (O_186,N_2769,N_2658);
nor UO_187 (O_187,N_2705,N_2501);
and UO_188 (O_188,N_2565,N_2863);
nand UO_189 (O_189,N_2964,N_2446);
nor UO_190 (O_190,N_2606,N_2831);
xnor UO_191 (O_191,N_2785,N_2518);
nor UO_192 (O_192,N_2930,N_2994);
and UO_193 (O_193,N_2690,N_2915);
nand UO_194 (O_194,N_2645,N_2853);
and UO_195 (O_195,N_2759,N_2798);
and UO_196 (O_196,N_2537,N_2917);
nand UO_197 (O_197,N_2940,N_2507);
nand UO_198 (O_198,N_2727,N_2779);
nor UO_199 (O_199,N_2659,N_2487);
nor UO_200 (O_200,N_2981,N_2898);
nor UO_201 (O_201,N_2751,N_2757);
nor UO_202 (O_202,N_2421,N_2897);
and UO_203 (O_203,N_2929,N_2411);
nand UO_204 (O_204,N_2706,N_2472);
or UO_205 (O_205,N_2616,N_2430);
nand UO_206 (O_206,N_2584,N_2828);
nor UO_207 (O_207,N_2588,N_2680);
nand UO_208 (O_208,N_2944,N_2854);
nor UO_209 (O_209,N_2693,N_2782);
and UO_210 (O_210,N_2675,N_2741);
nor UO_211 (O_211,N_2490,N_2740);
nor UO_212 (O_212,N_2580,N_2995);
or UO_213 (O_213,N_2669,N_2482);
nand UO_214 (O_214,N_2959,N_2946);
nor UO_215 (O_215,N_2403,N_2542);
or UO_216 (O_216,N_2927,N_2931);
and UO_217 (O_217,N_2781,N_2842);
nand UO_218 (O_218,N_2916,N_2671);
nor UO_219 (O_219,N_2998,N_2730);
xnor UO_220 (O_220,N_2442,N_2415);
or UO_221 (O_221,N_2846,N_2479);
or UO_222 (O_222,N_2526,N_2721);
nand UO_223 (O_223,N_2768,N_2943);
nand UO_224 (O_224,N_2938,N_2637);
and UO_225 (O_225,N_2743,N_2618);
nand UO_226 (O_226,N_2641,N_2418);
or UO_227 (O_227,N_2908,N_2895);
or UO_228 (O_228,N_2554,N_2848);
and UO_229 (O_229,N_2703,N_2794);
and UO_230 (O_230,N_2545,N_2791);
and UO_231 (O_231,N_2980,N_2505);
nor UO_232 (O_232,N_2500,N_2697);
and UO_233 (O_233,N_2566,N_2583);
or UO_234 (O_234,N_2685,N_2412);
or UO_235 (O_235,N_2960,N_2448);
nor UO_236 (O_236,N_2610,N_2689);
and UO_237 (O_237,N_2866,N_2484);
and UO_238 (O_238,N_2920,N_2533);
nand UO_239 (O_239,N_2725,N_2636);
nand UO_240 (O_240,N_2987,N_2710);
and UO_241 (O_241,N_2434,N_2700);
nor UO_242 (O_242,N_2459,N_2450);
and UO_243 (O_243,N_2570,N_2515);
nand UO_244 (O_244,N_2535,N_2674);
or UO_245 (O_245,N_2613,N_2604);
and UO_246 (O_246,N_2775,N_2867);
or UO_247 (O_247,N_2731,N_2875);
and UO_248 (O_248,N_2520,N_2473);
and UO_249 (O_249,N_2989,N_2899);
nand UO_250 (O_250,N_2586,N_2530);
nand UO_251 (O_251,N_2590,N_2855);
and UO_252 (O_252,N_2471,N_2827);
and UO_253 (O_253,N_2973,N_2813);
and UO_254 (O_254,N_2634,N_2589);
or UO_255 (O_255,N_2923,N_2596);
or UO_256 (O_256,N_2750,N_2576);
and UO_257 (O_257,N_2608,N_2651);
or UO_258 (O_258,N_2497,N_2556);
nor UO_259 (O_259,N_2822,N_2455);
nand UO_260 (O_260,N_2732,N_2752);
and UO_261 (O_261,N_2849,N_2928);
nor UO_262 (O_262,N_2517,N_2562);
nand UO_263 (O_263,N_2476,N_2692);
nor UO_264 (O_264,N_2754,N_2462);
nand UO_265 (O_265,N_2902,N_2551);
and UO_266 (O_266,N_2466,N_2889);
nor UO_267 (O_267,N_2632,N_2753);
and UO_268 (O_268,N_2624,N_2564);
nand UO_269 (O_269,N_2433,N_2502);
nor UO_270 (O_270,N_2561,N_2950);
nand UO_271 (O_271,N_2770,N_2529);
or UO_272 (O_272,N_2461,N_2480);
or UO_273 (O_273,N_2982,N_2402);
xnor UO_274 (O_274,N_2711,N_2648);
nand UO_275 (O_275,N_2707,N_2969);
nand UO_276 (O_276,N_2519,N_2567);
nor UO_277 (O_277,N_2414,N_2627);
nand UO_278 (O_278,N_2701,N_2571);
and UO_279 (O_279,N_2818,N_2972);
nor UO_280 (O_280,N_2633,N_2687);
nor UO_281 (O_281,N_2607,N_2724);
or UO_282 (O_282,N_2686,N_2838);
and UO_283 (O_283,N_2784,N_2829);
nor UO_284 (O_284,N_2602,N_2856);
nand UO_285 (O_285,N_2739,N_2925);
nand UO_286 (O_286,N_2864,N_2441);
nor UO_287 (O_287,N_2906,N_2614);
nand UO_288 (O_288,N_2738,N_2880);
nor UO_289 (O_289,N_2615,N_2877);
and UO_290 (O_290,N_2815,N_2859);
nand UO_291 (O_291,N_2804,N_2843);
nand UO_292 (O_292,N_2988,N_2797);
nand UO_293 (O_293,N_2601,N_2568);
xnor UO_294 (O_294,N_2555,N_2911);
or UO_295 (O_295,N_2400,N_2547);
or UO_296 (O_296,N_2424,N_2488);
nand UO_297 (O_297,N_2492,N_2726);
and UO_298 (O_298,N_2514,N_2548);
and UO_299 (O_299,N_2937,N_2825);
and UO_300 (O_300,N_2439,N_2676);
and UO_301 (O_301,N_2966,N_2859);
and UO_302 (O_302,N_2934,N_2541);
or UO_303 (O_303,N_2891,N_2976);
nor UO_304 (O_304,N_2495,N_2826);
nor UO_305 (O_305,N_2474,N_2533);
and UO_306 (O_306,N_2870,N_2416);
or UO_307 (O_307,N_2930,N_2795);
or UO_308 (O_308,N_2439,N_2780);
and UO_309 (O_309,N_2912,N_2747);
and UO_310 (O_310,N_2499,N_2890);
nor UO_311 (O_311,N_2814,N_2584);
nor UO_312 (O_312,N_2635,N_2747);
and UO_313 (O_313,N_2837,N_2534);
or UO_314 (O_314,N_2646,N_2919);
nand UO_315 (O_315,N_2653,N_2778);
nand UO_316 (O_316,N_2807,N_2587);
nand UO_317 (O_317,N_2533,N_2817);
nor UO_318 (O_318,N_2874,N_2904);
nand UO_319 (O_319,N_2842,N_2594);
or UO_320 (O_320,N_2412,N_2802);
nor UO_321 (O_321,N_2466,N_2624);
nor UO_322 (O_322,N_2891,N_2826);
nand UO_323 (O_323,N_2603,N_2563);
nor UO_324 (O_324,N_2934,N_2984);
and UO_325 (O_325,N_2561,N_2982);
or UO_326 (O_326,N_2615,N_2601);
and UO_327 (O_327,N_2881,N_2575);
nor UO_328 (O_328,N_2507,N_2427);
nand UO_329 (O_329,N_2420,N_2509);
or UO_330 (O_330,N_2413,N_2736);
nor UO_331 (O_331,N_2711,N_2483);
and UO_332 (O_332,N_2930,N_2818);
nor UO_333 (O_333,N_2977,N_2762);
or UO_334 (O_334,N_2788,N_2562);
nor UO_335 (O_335,N_2804,N_2784);
or UO_336 (O_336,N_2491,N_2764);
nand UO_337 (O_337,N_2601,N_2838);
and UO_338 (O_338,N_2749,N_2978);
nor UO_339 (O_339,N_2561,N_2931);
and UO_340 (O_340,N_2521,N_2781);
and UO_341 (O_341,N_2763,N_2881);
and UO_342 (O_342,N_2733,N_2743);
nand UO_343 (O_343,N_2754,N_2463);
nand UO_344 (O_344,N_2972,N_2566);
or UO_345 (O_345,N_2584,N_2612);
nor UO_346 (O_346,N_2844,N_2856);
nor UO_347 (O_347,N_2468,N_2714);
nand UO_348 (O_348,N_2779,N_2485);
nor UO_349 (O_349,N_2447,N_2562);
nor UO_350 (O_350,N_2602,N_2432);
nor UO_351 (O_351,N_2660,N_2667);
nand UO_352 (O_352,N_2635,N_2798);
and UO_353 (O_353,N_2807,N_2456);
nand UO_354 (O_354,N_2919,N_2535);
nand UO_355 (O_355,N_2602,N_2409);
or UO_356 (O_356,N_2832,N_2747);
or UO_357 (O_357,N_2556,N_2798);
nand UO_358 (O_358,N_2404,N_2632);
nand UO_359 (O_359,N_2816,N_2618);
nor UO_360 (O_360,N_2431,N_2556);
or UO_361 (O_361,N_2469,N_2952);
nand UO_362 (O_362,N_2957,N_2918);
and UO_363 (O_363,N_2845,N_2640);
nor UO_364 (O_364,N_2900,N_2516);
nand UO_365 (O_365,N_2536,N_2946);
nor UO_366 (O_366,N_2841,N_2431);
nor UO_367 (O_367,N_2536,N_2829);
nor UO_368 (O_368,N_2960,N_2986);
and UO_369 (O_369,N_2986,N_2633);
or UO_370 (O_370,N_2842,N_2532);
and UO_371 (O_371,N_2604,N_2567);
or UO_372 (O_372,N_2754,N_2712);
nor UO_373 (O_373,N_2678,N_2615);
nand UO_374 (O_374,N_2540,N_2867);
nor UO_375 (O_375,N_2732,N_2902);
or UO_376 (O_376,N_2568,N_2726);
nor UO_377 (O_377,N_2551,N_2711);
or UO_378 (O_378,N_2844,N_2528);
nand UO_379 (O_379,N_2857,N_2912);
nor UO_380 (O_380,N_2580,N_2671);
and UO_381 (O_381,N_2725,N_2775);
and UO_382 (O_382,N_2496,N_2852);
or UO_383 (O_383,N_2412,N_2958);
and UO_384 (O_384,N_2891,N_2581);
nor UO_385 (O_385,N_2844,N_2923);
nor UO_386 (O_386,N_2706,N_2537);
or UO_387 (O_387,N_2944,N_2739);
or UO_388 (O_388,N_2881,N_2624);
nand UO_389 (O_389,N_2479,N_2754);
or UO_390 (O_390,N_2980,N_2836);
nor UO_391 (O_391,N_2916,N_2519);
nand UO_392 (O_392,N_2775,N_2439);
nor UO_393 (O_393,N_2886,N_2730);
nor UO_394 (O_394,N_2638,N_2449);
nand UO_395 (O_395,N_2844,N_2892);
and UO_396 (O_396,N_2754,N_2845);
nand UO_397 (O_397,N_2889,N_2947);
and UO_398 (O_398,N_2958,N_2732);
nor UO_399 (O_399,N_2525,N_2967);
and UO_400 (O_400,N_2440,N_2569);
nor UO_401 (O_401,N_2676,N_2865);
or UO_402 (O_402,N_2610,N_2528);
and UO_403 (O_403,N_2441,N_2996);
nor UO_404 (O_404,N_2778,N_2559);
and UO_405 (O_405,N_2892,N_2869);
xor UO_406 (O_406,N_2569,N_2467);
nand UO_407 (O_407,N_2518,N_2503);
nor UO_408 (O_408,N_2606,N_2905);
or UO_409 (O_409,N_2935,N_2561);
and UO_410 (O_410,N_2960,N_2736);
nand UO_411 (O_411,N_2548,N_2476);
and UO_412 (O_412,N_2752,N_2822);
and UO_413 (O_413,N_2872,N_2746);
nand UO_414 (O_414,N_2486,N_2805);
or UO_415 (O_415,N_2586,N_2993);
nor UO_416 (O_416,N_2490,N_2416);
and UO_417 (O_417,N_2610,N_2926);
and UO_418 (O_418,N_2562,N_2458);
nand UO_419 (O_419,N_2928,N_2990);
or UO_420 (O_420,N_2563,N_2902);
nor UO_421 (O_421,N_2446,N_2520);
nand UO_422 (O_422,N_2988,N_2753);
and UO_423 (O_423,N_2782,N_2445);
and UO_424 (O_424,N_2419,N_2603);
and UO_425 (O_425,N_2815,N_2426);
nand UO_426 (O_426,N_2981,N_2949);
and UO_427 (O_427,N_2619,N_2710);
nand UO_428 (O_428,N_2574,N_2747);
nor UO_429 (O_429,N_2917,N_2531);
nor UO_430 (O_430,N_2996,N_2754);
nor UO_431 (O_431,N_2545,N_2968);
nor UO_432 (O_432,N_2523,N_2721);
nor UO_433 (O_433,N_2813,N_2633);
nor UO_434 (O_434,N_2698,N_2761);
and UO_435 (O_435,N_2561,N_2576);
xnor UO_436 (O_436,N_2670,N_2493);
or UO_437 (O_437,N_2970,N_2614);
and UO_438 (O_438,N_2468,N_2910);
nor UO_439 (O_439,N_2746,N_2835);
or UO_440 (O_440,N_2670,N_2639);
nor UO_441 (O_441,N_2547,N_2874);
nor UO_442 (O_442,N_2884,N_2976);
and UO_443 (O_443,N_2675,N_2923);
nand UO_444 (O_444,N_2786,N_2572);
nor UO_445 (O_445,N_2813,N_2857);
nand UO_446 (O_446,N_2810,N_2709);
and UO_447 (O_447,N_2518,N_2909);
nand UO_448 (O_448,N_2930,N_2499);
nand UO_449 (O_449,N_2950,N_2968);
nor UO_450 (O_450,N_2499,N_2871);
nand UO_451 (O_451,N_2705,N_2746);
nand UO_452 (O_452,N_2484,N_2825);
and UO_453 (O_453,N_2538,N_2957);
and UO_454 (O_454,N_2404,N_2569);
or UO_455 (O_455,N_2837,N_2926);
nor UO_456 (O_456,N_2971,N_2418);
or UO_457 (O_457,N_2951,N_2575);
nand UO_458 (O_458,N_2416,N_2459);
and UO_459 (O_459,N_2771,N_2924);
nor UO_460 (O_460,N_2694,N_2970);
and UO_461 (O_461,N_2422,N_2497);
nor UO_462 (O_462,N_2573,N_2653);
and UO_463 (O_463,N_2875,N_2433);
or UO_464 (O_464,N_2556,N_2708);
nand UO_465 (O_465,N_2833,N_2489);
nand UO_466 (O_466,N_2753,N_2714);
and UO_467 (O_467,N_2682,N_2422);
nand UO_468 (O_468,N_2754,N_2649);
nand UO_469 (O_469,N_2804,N_2507);
nand UO_470 (O_470,N_2832,N_2548);
nor UO_471 (O_471,N_2900,N_2792);
nor UO_472 (O_472,N_2746,N_2518);
nor UO_473 (O_473,N_2440,N_2937);
or UO_474 (O_474,N_2798,N_2592);
or UO_475 (O_475,N_2796,N_2806);
or UO_476 (O_476,N_2656,N_2702);
and UO_477 (O_477,N_2451,N_2641);
nor UO_478 (O_478,N_2523,N_2694);
nor UO_479 (O_479,N_2880,N_2450);
nand UO_480 (O_480,N_2876,N_2667);
nand UO_481 (O_481,N_2809,N_2414);
or UO_482 (O_482,N_2412,N_2954);
or UO_483 (O_483,N_2446,N_2866);
and UO_484 (O_484,N_2559,N_2665);
and UO_485 (O_485,N_2554,N_2715);
nand UO_486 (O_486,N_2513,N_2493);
and UO_487 (O_487,N_2526,N_2651);
and UO_488 (O_488,N_2850,N_2976);
or UO_489 (O_489,N_2546,N_2963);
nor UO_490 (O_490,N_2444,N_2513);
nor UO_491 (O_491,N_2926,N_2510);
or UO_492 (O_492,N_2435,N_2696);
and UO_493 (O_493,N_2843,N_2668);
nor UO_494 (O_494,N_2758,N_2420);
nor UO_495 (O_495,N_2833,N_2908);
nor UO_496 (O_496,N_2931,N_2754);
nand UO_497 (O_497,N_2481,N_2682);
and UO_498 (O_498,N_2701,N_2507);
nand UO_499 (O_499,N_2702,N_2891);
endmodule