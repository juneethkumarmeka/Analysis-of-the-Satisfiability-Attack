module basic_500_3000_500_60_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_306,In_19);
and U1 (N_1,In_128,In_347);
and U2 (N_2,In_337,In_265);
nor U3 (N_3,In_326,In_407);
nand U4 (N_4,In_282,In_37);
nand U5 (N_5,In_115,In_158);
nand U6 (N_6,In_84,In_109);
and U7 (N_7,In_134,In_429);
nand U8 (N_8,In_452,In_386);
or U9 (N_9,In_194,In_174);
nor U10 (N_10,In_129,In_322);
nand U11 (N_11,In_215,In_271);
and U12 (N_12,In_332,In_400);
xnor U13 (N_13,In_434,In_11);
and U14 (N_14,In_153,In_177);
and U15 (N_15,In_225,In_187);
nor U16 (N_16,In_117,In_294);
nand U17 (N_17,In_184,In_431);
and U18 (N_18,In_28,In_139);
nor U19 (N_19,In_159,In_257);
or U20 (N_20,In_258,In_165);
or U21 (N_21,In_68,In_42);
nand U22 (N_22,In_412,In_395);
or U23 (N_23,In_490,In_104);
nor U24 (N_24,In_263,In_107);
nand U25 (N_25,In_405,In_100);
nor U26 (N_26,In_415,In_471);
or U27 (N_27,In_232,In_18);
nand U28 (N_28,In_53,In_195);
or U29 (N_29,In_192,In_460);
or U30 (N_30,In_489,In_176);
or U31 (N_31,In_166,In_150);
and U32 (N_32,In_61,In_143);
or U33 (N_33,In_323,In_410);
or U34 (N_34,In_210,In_457);
or U35 (N_35,In_438,In_356);
nand U36 (N_36,In_329,In_246);
or U37 (N_37,In_133,In_487);
or U38 (N_38,In_335,In_341);
and U39 (N_39,In_454,In_307);
and U40 (N_40,In_58,In_51);
and U41 (N_41,In_21,In_288);
or U42 (N_42,In_342,In_126);
and U43 (N_43,In_87,In_496);
nand U44 (N_44,In_334,In_259);
nand U45 (N_45,In_238,In_3);
nand U46 (N_46,In_64,In_339);
or U47 (N_47,In_445,In_488);
and U48 (N_48,In_244,In_144);
or U49 (N_49,In_388,In_82);
and U50 (N_50,In_469,In_237);
nand U51 (N_51,In_127,In_151);
nor U52 (N_52,In_125,In_304);
nand U53 (N_53,In_262,In_264);
or U54 (N_54,In_57,In_299);
nor U55 (N_55,In_131,In_396);
or U56 (N_56,In_448,In_92);
nor U57 (N_57,In_408,In_204);
nor U58 (N_58,In_80,In_170);
or U59 (N_59,N_44,In_212);
nand U60 (N_60,In_316,N_12);
nand U61 (N_61,In_274,In_137);
nand U62 (N_62,In_474,In_378);
xnor U63 (N_63,In_463,In_135);
nand U64 (N_64,In_498,N_48);
nand U65 (N_65,In_376,N_19);
nor U66 (N_66,In_494,In_152);
or U67 (N_67,In_77,In_56);
nand U68 (N_68,N_42,In_358);
and U69 (N_69,In_24,In_15);
or U70 (N_70,In_373,In_303);
or U71 (N_71,In_136,N_6);
nand U72 (N_72,N_30,In_312);
xnor U73 (N_73,In_313,In_71);
or U74 (N_74,In_449,In_470);
and U75 (N_75,N_38,In_97);
and U76 (N_76,In_462,In_252);
nand U77 (N_77,In_477,In_140);
nand U78 (N_78,In_466,In_267);
nand U79 (N_79,In_10,In_268);
nand U80 (N_80,N_11,In_359);
or U81 (N_81,In_285,In_355);
nor U82 (N_82,In_75,In_30);
and U83 (N_83,In_442,N_14);
nand U84 (N_84,In_66,In_230);
nor U85 (N_85,In_214,In_436);
or U86 (N_86,In_227,In_298);
or U87 (N_87,In_7,In_468);
nand U88 (N_88,N_49,N_35);
nand U89 (N_89,In_317,In_38);
nand U90 (N_90,In_2,In_86);
nand U91 (N_91,In_31,In_254);
or U92 (N_92,In_62,In_72);
nand U93 (N_93,In_450,In_451);
and U94 (N_94,In_394,In_392);
nand U95 (N_95,In_147,In_22);
or U96 (N_96,In_65,In_275);
and U97 (N_97,In_121,In_455);
and U98 (N_98,In_251,In_141);
nand U99 (N_99,In_497,N_7);
nand U100 (N_100,In_379,In_91);
nand U101 (N_101,In_132,In_340);
or U102 (N_102,In_495,In_52);
and U103 (N_103,In_371,In_499);
or U104 (N_104,In_309,In_280);
and U105 (N_105,In_154,In_33);
and U106 (N_106,In_404,In_467);
nor U107 (N_107,In_351,In_1);
or U108 (N_108,N_21,N_24);
nor U109 (N_109,In_12,In_302);
or U110 (N_110,N_63,In_433);
nor U111 (N_111,In_428,N_53);
or U112 (N_112,N_8,In_23);
and U113 (N_113,N_86,N_65);
or U114 (N_114,In_156,N_10);
and U115 (N_115,N_61,In_146);
or U116 (N_116,N_73,In_486);
nand U117 (N_117,N_68,In_180);
nor U118 (N_118,N_88,In_476);
nor U119 (N_119,In_363,In_325);
xor U120 (N_120,N_47,In_456);
or U121 (N_121,In_20,In_219);
nor U122 (N_122,In_34,In_14);
and U123 (N_123,N_50,N_37);
nor U124 (N_124,In_96,In_491);
or U125 (N_125,N_45,In_300);
nand U126 (N_126,In_393,N_74);
and U127 (N_127,In_402,In_48);
or U128 (N_128,In_223,In_206);
or U129 (N_129,In_441,In_324);
or U130 (N_130,In_191,In_105);
nand U131 (N_131,N_39,In_362);
nand U132 (N_132,In_493,N_58);
nor U133 (N_133,In_171,In_284);
nand U134 (N_134,In_399,In_220);
nand U135 (N_135,In_183,In_245);
nand U136 (N_136,In_295,In_122);
nand U137 (N_137,N_41,In_269);
or U138 (N_138,In_461,In_277);
or U139 (N_139,In_361,N_64);
nand U140 (N_140,N_20,In_99);
nand U141 (N_141,In_124,In_443);
and U142 (N_142,In_403,In_76);
xor U143 (N_143,In_293,In_439);
and U144 (N_144,In_243,In_397);
nand U145 (N_145,N_5,In_483);
or U146 (N_146,In_364,N_79);
or U147 (N_147,In_46,In_182);
or U148 (N_148,In_235,N_75);
nor U149 (N_149,In_482,In_167);
and U150 (N_150,In_387,In_5);
or U151 (N_151,N_56,N_101);
or U152 (N_152,In_207,In_173);
nor U153 (N_153,In_458,N_46);
nor U154 (N_154,N_40,In_198);
nand U155 (N_155,In_116,In_260);
or U156 (N_156,In_54,N_94);
nor U157 (N_157,In_286,N_2);
nand U158 (N_158,In_50,N_126);
nand U159 (N_159,N_22,In_163);
or U160 (N_160,In_473,In_222);
or U161 (N_161,N_108,In_142);
nor U162 (N_162,In_327,N_90);
nor U163 (N_163,In_377,N_25);
nor U164 (N_164,N_148,In_118);
and U165 (N_165,In_168,In_345);
or U166 (N_166,In_218,N_124);
or U167 (N_167,N_139,In_242);
or U168 (N_168,In_270,N_106);
nand U169 (N_169,In_8,In_465);
and U170 (N_170,In_103,In_343);
nor U171 (N_171,In_106,N_105);
and U172 (N_172,In_49,In_240);
and U173 (N_173,N_123,In_276);
and U174 (N_174,N_33,N_109);
or U175 (N_175,In_85,In_63);
nand U176 (N_176,In_0,In_432);
and U177 (N_177,In_74,N_0);
nor U178 (N_178,In_224,N_82);
nor U179 (N_179,In_190,N_83);
nand U180 (N_180,N_52,In_385);
or U181 (N_181,In_196,In_484);
nand U182 (N_182,N_60,In_374);
and U183 (N_183,In_89,In_338);
nor U184 (N_184,N_96,In_426);
or U185 (N_185,In_247,N_62);
nor U186 (N_186,In_81,In_289);
nand U187 (N_187,In_79,In_459);
nand U188 (N_188,In_199,In_60);
nand U189 (N_189,In_221,In_231);
nor U190 (N_190,In_348,In_211);
xnor U191 (N_191,In_205,In_305);
and U192 (N_192,In_301,In_380);
and U193 (N_193,In_279,N_112);
nor U194 (N_194,In_485,N_134);
nand U195 (N_195,In_93,In_73);
and U196 (N_196,In_90,In_440);
nor U197 (N_197,In_88,In_391);
or U198 (N_198,In_447,N_23);
or U199 (N_199,In_43,In_114);
or U200 (N_200,In_175,N_187);
nand U201 (N_201,N_197,In_47);
nor U202 (N_202,In_112,In_188);
and U203 (N_203,N_55,N_177);
nor U204 (N_204,N_164,In_41);
and U205 (N_205,N_17,In_197);
and U206 (N_206,In_398,N_51);
and U207 (N_207,In_383,N_180);
nand U208 (N_208,In_375,N_16);
nor U209 (N_209,In_353,In_266);
nor U210 (N_210,N_161,N_95);
or U211 (N_211,N_32,In_4);
or U212 (N_212,In_256,In_145);
or U213 (N_213,In_401,N_128);
nor U214 (N_214,In_370,In_427);
nand U215 (N_215,N_93,In_365);
nor U216 (N_216,In_44,N_115);
and U217 (N_217,In_318,In_311);
or U218 (N_218,In_281,In_480);
or U219 (N_219,In_354,In_113);
nand U220 (N_220,In_13,In_420);
xnor U221 (N_221,In_200,N_54);
nand U222 (N_222,N_72,In_320);
or U223 (N_223,In_255,In_9);
nor U224 (N_224,N_9,In_179);
nand U225 (N_225,In_226,N_129);
and U226 (N_226,In_148,N_162);
or U227 (N_227,In_384,In_59);
or U228 (N_228,N_70,In_185);
and U229 (N_229,In_169,N_150);
and U230 (N_230,N_184,In_352);
or U231 (N_231,In_366,N_188);
nand U232 (N_232,In_278,In_181);
nor U233 (N_233,In_328,In_344);
and U234 (N_234,In_213,In_349);
or U235 (N_235,N_183,In_250);
nor U236 (N_236,N_15,N_151);
and U237 (N_237,In_417,In_229);
nor U238 (N_238,N_172,In_389);
nand U239 (N_239,In_102,N_196);
nand U240 (N_240,In_418,In_413);
or U241 (N_241,N_97,In_228);
and U242 (N_242,In_216,N_157);
or U243 (N_243,N_149,N_78);
nand U244 (N_244,In_248,N_4);
and U245 (N_245,In_108,In_360);
or U246 (N_246,N_141,N_116);
nor U247 (N_247,In_162,N_171);
nand U248 (N_248,N_192,N_198);
or U249 (N_249,N_1,In_25);
and U250 (N_250,In_161,N_217);
and U251 (N_251,N_69,N_232);
or U252 (N_252,N_110,In_35);
or U253 (N_253,N_154,N_59);
nor U254 (N_254,In_425,In_390);
nor U255 (N_255,In_416,N_207);
nand U256 (N_256,In_32,In_287);
nor U257 (N_257,In_78,In_336);
nor U258 (N_258,In_16,N_137);
or U259 (N_259,N_221,N_166);
or U260 (N_260,N_200,In_291);
nor U261 (N_261,In_292,In_283);
or U262 (N_262,N_122,N_210);
or U263 (N_263,N_249,In_453);
and U264 (N_264,In_414,N_194);
nor U265 (N_265,In_430,In_155);
and U266 (N_266,N_237,N_155);
nor U267 (N_267,N_160,N_34);
or U268 (N_268,N_247,In_464);
and U269 (N_269,In_350,N_117);
nor U270 (N_270,In_249,In_193);
nor U271 (N_271,N_27,N_233);
and U272 (N_272,N_204,N_181);
or U273 (N_273,N_100,In_492);
nor U274 (N_274,N_231,N_211);
or U275 (N_275,In_164,N_118);
nor U276 (N_276,N_216,In_29);
nor U277 (N_277,In_120,N_223);
or U278 (N_278,N_173,N_111);
nor U279 (N_279,N_36,In_369);
nor U280 (N_280,In_296,In_479);
nor U281 (N_281,In_272,N_26);
nor U282 (N_282,N_175,N_229);
nor U283 (N_283,N_244,In_6);
nand U284 (N_284,N_145,In_321);
nand U285 (N_285,In_478,In_101);
or U286 (N_286,N_159,N_132);
xor U287 (N_287,N_167,N_222);
or U288 (N_288,N_104,N_178);
or U289 (N_289,N_18,In_419);
nor U290 (N_290,In_346,N_77);
or U291 (N_291,N_131,In_236);
or U292 (N_292,In_149,In_83);
nand U293 (N_293,In_472,In_424);
nor U294 (N_294,In_160,In_189);
nor U295 (N_295,N_67,In_69);
or U296 (N_296,In_310,N_127);
and U297 (N_297,In_382,N_133);
nor U298 (N_298,N_239,N_121);
nor U299 (N_299,In_422,N_80);
or U300 (N_300,N_273,N_257);
or U301 (N_301,N_213,N_290);
nor U302 (N_302,N_240,N_238);
nor U303 (N_303,N_297,In_290);
nor U304 (N_304,N_214,N_283);
and U305 (N_305,N_3,N_259);
and U306 (N_306,In_178,In_261);
and U307 (N_307,In_208,In_409);
nor U308 (N_308,In_331,N_219);
and U309 (N_309,In_315,N_103);
and U310 (N_310,In_157,N_203);
nor U311 (N_311,N_113,N_102);
and U312 (N_312,N_208,In_123);
nor U313 (N_313,N_242,In_319);
xnor U314 (N_314,N_255,N_13);
and U315 (N_315,N_142,N_268);
and U316 (N_316,N_182,N_272);
nor U317 (N_317,In_26,N_277);
nand U318 (N_318,N_28,N_264);
nand U319 (N_319,N_202,N_270);
nor U320 (N_320,N_84,N_119);
nor U321 (N_321,N_125,N_248);
or U322 (N_322,N_215,N_195);
and U323 (N_323,In_381,N_246);
xnor U324 (N_324,In_475,N_298);
nor U325 (N_325,In_172,In_297);
nor U326 (N_326,N_146,N_279);
xor U327 (N_327,In_119,In_233);
nand U328 (N_328,N_292,N_236);
nand U329 (N_329,In_111,N_92);
nor U330 (N_330,N_174,N_220);
xor U331 (N_331,N_165,In_45);
and U332 (N_332,N_269,N_99);
nor U333 (N_333,N_263,N_254);
or U334 (N_334,N_296,N_87);
nor U335 (N_335,N_286,In_202);
or U336 (N_336,In_357,N_241);
and U337 (N_337,N_287,N_107);
nor U338 (N_338,N_66,N_235);
and U339 (N_339,N_289,N_186);
nor U340 (N_340,In_273,In_241);
nor U341 (N_341,In_27,N_227);
nand U342 (N_342,In_130,N_156);
and U343 (N_343,N_299,In_437);
nand U344 (N_344,N_252,In_110);
nand U345 (N_345,N_201,N_230);
or U346 (N_346,N_114,In_368);
nor U347 (N_347,N_291,In_217);
and U348 (N_348,N_76,In_36);
nor U349 (N_349,N_275,N_85);
nor U350 (N_350,In_70,N_98);
or U351 (N_351,N_260,In_421);
nor U352 (N_352,In_67,N_176);
nand U353 (N_353,N_265,N_305);
or U354 (N_354,N_89,N_323);
and U355 (N_355,N_185,N_338);
or U356 (N_356,N_321,N_343);
and U357 (N_357,N_302,N_330);
nor U358 (N_358,N_193,In_234);
or U359 (N_359,N_303,N_271);
nor U360 (N_360,N_81,N_256);
nand U361 (N_361,N_312,In_446);
nand U362 (N_362,N_328,In_203);
and U363 (N_363,N_234,N_306);
nor U364 (N_364,In_411,N_301);
nor U365 (N_365,N_319,N_224);
or U366 (N_366,N_331,N_261);
or U367 (N_367,In_330,N_320);
and U368 (N_368,In_308,N_170);
nor U369 (N_369,N_327,N_288);
nand U370 (N_370,N_147,N_313);
or U371 (N_371,N_324,N_189);
nor U372 (N_372,N_158,In_17);
and U373 (N_373,N_31,N_136);
or U374 (N_374,N_317,N_43);
nand U375 (N_375,N_267,In_138);
or U376 (N_376,In_367,N_332);
nand U377 (N_377,N_294,In_314);
nand U378 (N_378,N_57,N_326);
xor U379 (N_379,N_339,N_334);
nand U380 (N_380,N_199,N_91);
or U381 (N_381,N_205,In_40);
and U382 (N_382,N_212,N_304);
nor U383 (N_383,In_372,N_266);
nor U384 (N_384,In_201,N_190);
nor U385 (N_385,N_143,N_163);
nor U386 (N_386,In_39,In_481);
nor U387 (N_387,N_168,In_423);
nor U388 (N_388,N_300,N_276);
nand U389 (N_389,N_348,N_285);
nor U390 (N_390,N_322,N_345);
nor U391 (N_391,N_310,N_329);
nand U392 (N_392,N_280,N_284);
nand U393 (N_393,N_340,In_435);
nand U394 (N_394,N_318,N_169);
nand U395 (N_395,N_314,In_94);
nand U396 (N_396,N_153,In_95);
and U397 (N_397,In_209,N_152);
nor U398 (N_398,N_140,N_253);
and U399 (N_399,N_251,N_342);
nand U400 (N_400,N_228,N_398);
or U401 (N_401,N_362,N_120);
xnor U402 (N_402,N_377,N_352);
nor U403 (N_403,N_308,N_144);
or U404 (N_404,N_378,N_381);
nand U405 (N_405,N_337,N_347);
nand U406 (N_406,N_179,N_335);
nand U407 (N_407,N_361,In_98);
or U408 (N_408,N_374,N_354);
nor U409 (N_409,N_364,N_386);
or U410 (N_410,N_389,N_357);
and U411 (N_411,N_359,N_243);
or U412 (N_412,N_226,N_367);
nor U413 (N_413,N_316,N_384);
and U414 (N_414,N_369,N_397);
nor U415 (N_415,N_293,N_346);
nor U416 (N_416,N_209,N_325);
or U417 (N_417,In_253,N_315);
or U418 (N_418,N_383,N_399);
or U419 (N_419,N_373,N_385);
nor U420 (N_420,In_333,N_71);
or U421 (N_421,N_375,N_295);
and U422 (N_422,N_358,N_135);
and U423 (N_423,N_388,In_239);
or U424 (N_424,N_382,N_387);
or U425 (N_425,N_396,N_282);
nor U426 (N_426,In_186,N_394);
nand U427 (N_427,N_371,N_218);
and U428 (N_428,In_444,N_353);
or U429 (N_429,N_258,N_191);
or U430 (N_430,N_130,N_307);
and U431 (N_431,In_55,N_250);
nor U432 (N_432,N_392,N_370);
nor U433 (N_433,N_336,N_225);
or U434 (N_434,N_390,N_262);
and U435 (N_435,N_341,N_356);
and U436 (N_436,N_372,N_278);
or U437 (N_437,N_350,N_380);
or U438 (N_438,N_355,N_395);
nand U439 (N_439,N_376,N_333);
nor U440 (N_440,N_365,N_349);
nor U441 (N_441,N_391,N_393);
nand U442 (N_442,N_363,N_281);
nand U443 (N_443,N_351,N_29);
nor U444 (N_444,N_379,In_406);
or U445 (N_445,N_344,N_309);
nor U446 (N_446,N_311,N_360);
and U447 (N_447,N_138,N_206);
and U448 (N_448,N_368,N_366);
nand U449 (N_449,N_274,N_245);
or U450 (N_450,N_448,N_440);
and U451 (N_451,N_435,N_412);
nor U452 (N_452,N_422,N_425);
or U453 (N_453,N_407,N_406);
nand U454 (N_454,N_414,N_447);
nor U455 (N_455,N_432,N_429);
or U456 (N_456,N_442,N_415);
nor U457 (N_457,N_426,N_402);
and U458 (N_458,N_437,N_404);
nor U459 (N_459,N_421,N_424);
or U460 (N_460,N_434,N_436);
nor U461 (N_461,N_431,N_427);
or U462 (N_462,N_443,N_441);
nor U463 (N_463,N_400,N_449);
nand U464 (N_464,N_444,N_419);
nand U465 (N_465,N_409,N_439);
nand U466 (N_466,N_423,N_410);
nor U467 (N_467,N_408,N_438);
nor U468 (N_468,N_433,N_411);
and U469 (N_469,N_405,N_430);
nor U470 (N_470,N_418,N_401);
and U471 (N_471,N_417,N_446);
nand U472 (N_472,N_413,N_416);
or U473 (N_473,N_428,N_445);
nand U474 (N_474,N_403,N_420);
or U475 (N_475,N_406,N_433);
and U476 (N_476,N_430,N_429);
nand U477 (N_477,N_419,N_430);
nor U478 (N_478,N_423,N_434);
or U479 (N_479,N_423,N_428);
nor U480 (N_480,N_436,N_442);
and U481 (N_481,N_421,N_404);
nor U482 (N_482,N_434,N_414);
xor U483 (N_483,N_449,N_422);
and U484 (N_484,N_445,N_442);
or U485 (N_485,N_410,N_402);
nor U486 (N_486,N_400,N_430);
nand U487 (N_487,N_441,N_409);
nor U488 (N_488,N_429,N_424);
nor U489 (N_489,N_404,N_420);
or U490 (N_490,N_411,N_437);
nand U491 (N_491,N_415,N_401);
and U492 (N_492,N_405,N_422);
nor U493 (N_493,N_415,N_424);
nand U494 (N_494,N_438,N_446);
nand U495 (N_495,N_419,N_423);
nand U496 (N_496,N_411,N_407);
nor U497 (N_497,N_410,N_403);
and U498 (N_498,N_446,N_402);
and U499 (N_499,N_409,N_424);
and U500 (N_500,N_483,N_494);
or U501 (N_501,N_481,N_477);
or U502 (N_502,N_465,N_475);
and U503 (N_503,N_487,N_478);
and U504 (N_504,N_496,N_463);
nand U505 (N_505,N_472,N_489);
nand U506 (N_506,N_466,N_462);
nor U507 (N_507,N_486,N_469);
nand U508 (N_508,N_476,N_479);
or U509 (N_509,N_474,N_464);
or U510 (N_510,N_467,N_473);
or U511 (N_511,N_454,N_495);
and U512 (N_512,N_459,N_482);
xor U513 (N_513,N_492,N_455);
or U514 (N_514,N_488,N_484);
xor U515 (N_515,N_460,N_468);
or U516 (N_516,N_485,N_480);
or U517 (N_517,N_497,N_456);
nand U518 (N_518,N_499,N_491);
and U519 (N_519,N_471,N_493);
or U520 (N_520,N_457,N_470);
nand U521 (N_521,N_450,N_490);
and U522 (N_522,N_458,N_452);
nor U523 (N_523,N_498,N_461);
or U524 (N_524,N_451,N_453);
xor U525 (N_525,N_475,N_467);
nand U526 (N_526,N_478,N_456);
nand U527 (N_527,N_450,N_470);
nand U528 (N_528,N_460,N_466);
nor U529 (N_529,N_459,N_456);
and U530 (N_530,N_489,N_473);
or U531 (N_531,N_460,N_485);
or U532 (N_532,N_454,N_467);
nor U533 (N_533,N_490,N_485);
and U534 (N_534,N_476,N_465);
or U535 (N_535,N_461,N_476);
or U536 (N_536,N_464,N_493);
nor U537 (N_537,N_460,N_474);
nor U538 (N_538,N_465,N_460);
and U539 (N_539,N_481,N_470);
nand U540 (N_540,N_489,N_469);
and U541 (N_541,N_496,N_487);
and U542 (N_542,N_484,N_494);
nand U543 (N_543,N_464,N_459);
or U544 (N_544,N_483,N_463);
or U545 (N_545,N_466,N_480);
or U546 (N_546,N_483,N_496);
and U547 (N_547,N_457,N_498);
nor U548 (N_548,N_469,N_471);
or U549 (N_549,N_466,N_463);
and U550 (N_550,N_501,N_507);
nor U551 (N_551,N_540,N_547);
nand U552 (N_552,N_518,N_534);
nor U553 (N_553,N_508,N_515);
nor U554 (N_554,N_509,N_532);
nand U555 (N_555,N_512,N_536);
nand U556 (N_556,N_514,N_513);
and U557 (N_557,N_535,N_504);
nor U558 (N_558,N_539,N_511);
xor U559 (N_559,N_503,N_546);
and U560 (N_560,N_520,N_533);
nand U561 (N_561,N_523,N_510);
nand U562 (N_562,N_506,N_538);
nor U563 (N_563,N_505,N_502);
nand U564 (N_564,N_500,N_524);
nor U565 (N_565,N_545,N_549);
or U566 (N_566,N_543,N_542);
and U567 (N_567,N_541,N_522);
or U568 (N_568,N_528,N_529);
xnor U569 (N_569,N_527,N_519);
or U570 (N_570,N_537,N_521);
nand U571 (N_571,N_530,N_526);
or U572 (N_572,N_531,N_525);
and U573 (N_573,N_517,N_548);
or U574 (N_574,N_544,N_516);
nor U575 (N_575,N_502,N_512);
xor U576 (N_576,N_545,N_532);
or U577 (N_577,N_539,N_540);
or U578 (N_578,N_529,N_502);
nor U579 (N_579,N_503,N_525);
nand U580 (N_580,N_511,N_528);
nand U581 (N_581,N_525,N_507);
nand U582 (N_582,N_535,N_529);
and U583 (N_583,N_507,N_545);
nor U584 (N_584,N_516,N_503);
nor U585 (N_585,N_544,N_525);
nand U586 (N_586,N_529,N_505);
nor U587 (N_587,N_510,N_517);
and U588 (N_588,N_524,N_531);
and U589 (N_589,N_504,N_528);
or U590 (N_590,N_540,N_515);
xnor U591 (N_591,N_543,N_506);
nor U592 (N_592,N_516,N_543);
and U593 (N_593,N_528,N_530);
and U594 (N_594,N_503,N_530);
nand U595 (N_595,N_500,N_521);
nor U596 (N_596,N_500,N_525);
or U597 (N_597,N_526,N_509);
and U598 (N_598,N_518,N_523);
or U599 (N_599,N_533,N_535);
or U600 (N_600,N_555,N_576);
and U601 (N_601,N_578,N_560);
and U602 (N_602,N_557,N_550);
and U603 (N_603,N_593,N_592);
nor U604 (N_604,N_583,N_579);
nand U605 (N_605,N_589,N_598);
nand U606 (N_606,N_552,N_595);
nand U607 (N_607,N_590,N_571);
nand U608 (N_608,N_597,N_556);
nor U609 (N_609,N_584,N_568);
and U610 (N_610,N_559,N_553);
xnor U611 (N_611,N_554,N_566);
or U612 (N_612,N_567,N_551);
and U613 (N_613,N_577,N_599);
or U614 (N_614,N_569,N_588);
nand U615 (N_615,N_591,N_572);
nand U616 (N_616,N_563,N_581);
nand U617 (N_617,N_565,N_585);
or U618 (N_618,N_582,N_573);
or U619 (N_619,N_570,N_575);
or U620 (N_620,N_580,N_561);
nand U621 (N_621,N_594,N_587);
and U622 (N_622,N_596,N_574);
and U623 (N_623,N_558,N_586);
nor U624 (N_624,N_564,N_562);
nand U625 (N_625,N_564,N_560);
and U626 (N_626,N_582,N_586);
nor U627 (N_627,N_551,N_590);
nand U628 (N_628,N_557,N_595);
and U629 (N_629,N_556,N_583);
or U630 (N_630,N_588,N_560);
and U631 (N_631,N_590,N_574);
nor U632 (N_632,N_552,N_555);
or U633 (N_633,N_590,N_588);
nor U634 (N_634,N_563,N_561);
nor U635 (N_635,N_599,N_552);
nor U636 (N_636,N_573,N_557);
nand U637 (N_637,N_594,N_599);
nor U638 (N_638,N_557,N_588);
or U639 (N_639,N_568,N_571);
and U640 (N_640,N_593,N_586);
or U641 (N_641,N_593,N_574);
nor U642 (N_642,N_595,N_567);
or U643 (N_643,N_587,N_555);
and U644 (N_644,N_582,N_579);
and U645 (N_645,N_567,N_593);
and U646 (N_646,N_567,N_599);
nand U647 (N_647,N_553,N_595);
or U648 (N_648,N_550,N_556);
or U649 (N_649,N_588,N_550);
or U650 (N_650,N_644,N_616);
and U651 (N_651,N_626,N_625);
nor U652 (N_652,N_622,N_606);
nor U653 (N_653,N_627,N_631);
xnor U654 (N_654,N_629,N_632);
and U655 (N_655,N_614,N_637);
nand U656 (N_656,N_618,N_628);
nand U657 (N_657,N_641,N_602);
nand U658 (N_658,N_630,N_612);
nor U659 (N_659,N_603,N_633);
nand U660 (N_660,N_607,N_611);
and U661 (N_661,N_624,N_640);
and U662 (N_662,N_609,N_636);
or U663 (N_663,N_642,N_615);
nand U664 (N_664,N_646,N_617);
nand U665 (N_665,N_610,N_621);
nand U666 (N_666,N_601,N_604);
or U667 (N_667,N_620,N_649);
nor U668 (N_668,N_635,N_639);
nand U669 (N_669,N_623,N_605);
nor U670 (N_670,N_608,N_645);
or U671 (N_671,N_613,N_638);
nor U672 (N_672,N_648,N_619);
nand U673 (N_673,N_634,N_647);
and U674 (N_674,N_600,N_643);
or U675 (N_675,N_609,N_646);
or U676 (N_676,N_633,N_639);
nor U677 (N_677,N_602,N_628);
and U678 (N_678,N_619,N_628);
and U679 (N_679,N_614,N_633);
nand U680 (N_680,N_647,N_639);
nor U681 (N_681,N_624,N_647);
and U682 (N_682,N_615,N_614);
or U683 (N_683,N_629,N_622);
nor U684 (N_684,N_608,N_646);
nor U685 (N_685,N_646,N_605);
and U686 (N_686,N_608,N_612);
nand U687 (N_687,N_603,N_626);
nand U688 (N_688,N_620,N_621);
nand U689 (N_689,N_638,N_617);
and U690 (N_690,N_648,N_649);
and U691 (N_691,N_607,N_614);
or U692 (N_692,N_636,N_608);
nor U693 (N_693,N_635,N_613);
and U694 (N_694,N_602,N_623);
nand U695 (N_695,N_643,N_648);
and U696 (N_696,N_615,N_616);
and U697 (N_697,N_610,N_648);
nand U698 (N_698,N_610,N_639);
nand U699 (N_699,N_647,N_621);
or U700 (N_700,N_667,N_695);
xnor U701 (N_701,N_657,N_674);
and U702 (N_702,N_686,N_671);
nand U703 (N_703,N_687,N_665);
or U704 (N_704,N_661,N_669);
or U705 (N_705,N_676,N_691);
nor U706 (N_706,N_696,N_681);
and U707 (N_707,N_652,N_677);
nor U708 (N_708,N_662,N_693);
nor U709 (N_709,N_694,N_670);
and U710 (N_710,N_688,N_650);
nand U711 (N_711,N_685,N_654);
or U712 (N_712,N_656,N_673);
xor U713 (N_713,N_697,N_660);
nor U714 (N_714,N_659,N_680);
or U715 (N_715,N_679,N_668);
or U716 (N_716,N_672,N_655);
nor U717 (N_717,N_698,N_683);
nand U718 (N_718,N_692,N_651);
nand U719 (N_719,N_666,N_699);
or U720 (N_720,N_678,N_675);
or U721 (N_721,N_653,N_690);
or U722 (N_722,N_658,N_689);
or U723 (N_723,N_663,N_664);
and U724 (N_724,N_682,N_684);
and U725 (N_725,N_656,N_660);
nand U726 (N_726,N_666,N_692);
nor U727 (N_727,N_659,N_652);
and U728 (N_728,N_667,N_662);
or U729 (N_729,N_699,N_697);
or U730 (N_730,N_692,N_680);
xnor U731 (N_731,N_650,N_673);
nor U732 (N_732,N_679,N_653);
and U733 (N_733,N_666,N_673);
and U734 (N_734,N_675,N_656);
and U735 (N_735,N_670,N_673);
nor U736 (N_736,N_650,N_679);
nor U737 (N_737,N_692,N_682);
and U738 (N_738,N_657,N_663);
nor U739 (N_739,N_677,N_692);
nand U740 (N_740,N_650,N_682);
and U741 (N_741,N_664,N_667);
or U742 (N_742,N_679,N_683);
nand U743 (N_743,N_686,N_658);
nand U744 (N_744,N_676,N_651);
or U745 (N_745,N_667,N_678);
or U746 (N_746,N_689,N_664);
or U747 (N_747,N_683,N_681);
nor U748 (N_748,N_680,N_662);
or U749 (N_749,N_688,N_678);
nand U750 (N_750,N_736,N_715);
nand U751 (N_751,N_739,N_747);
or U752 (N_752,N_746,N_731);
and U753 (N_753,N_738,N_730);
and U754 (N_754,N_732,N_700);
and U755 (N_755,N_724,N_745);
and U756 (N_756,N_734,N_733);
nand U757 (N_757,N_712,N_718);
or U758 (N_758,N_744,N_721);
or U759 (N_759,N_743,N_716);
and U760 (N_760,N_704,N_725);
or U761 (N_761,N_729,N_735);
xnor U762 (N_762,N_726,N_749);
or U763 (N_763,N_701,N_702);
and U764 (N_764,N_720,N_737);
nor U765 (N_765,N_741,N_706);
nor U766 (N_766,N_727,N_748);
nand U767 (N_767,N_728,N_722);
and U768 (N_768,N_719,N_740);
and U769 (N_769,N_723,N_714);
nand U770 (N_770,N_711,N_708);
nor U771 (N_771,N_742,N_703);
or U772 (N_772,N_717,N_707);
nand U773 (N_773,N_709,N_705);
and U774 (N_774,N_710,N_713);
and U775 (N_775,N_730,N_720);
nand U776 (N_776,N_738,N_711);
or U777 (N_777,N_742,N_706);
nand U778 (N_778,N_746,N_730);
and U779 (N_779,N_714,N_737);
nor U780 (N_780,N_716,N_700);
nor U781 (N_781,N_722,N_730);
nor U782 (N_782,N_745,N_719);
nand U783 (N_783,N_723,N_716);
nand U784 (N_784,N_728,N_734);
nand U785 (N_785,N_710,N_720);
and U786 (N_786,N_732,N_713);
and U787 (N_787,N_733,N_720);
and U788 (N_788,N_743,N_714);
or U789 (N_789,N_743,N_727);
or U790 (N_790,N_711,N_736);
nand U791 (N_791,N_716,N_718);
nor U792 (N_792,N_713,N_741);
or U793 (N_793,N_725,N_734);
nand U794 (N_794,N_744,N_708);
and U795 (N_795,N_731,N_719);
or U796 (N_796,N_744,N_731);
and U797 (N_797,N_717,N_706);
nand U798 (N_798,N_702,N_720);
or U799 (N_799,N_732,N_701);
and U800 (N_800,N_761,N_787);
nand U801 (N_801,N_796,N_755);
or U802 (N_802,N_751,N_782);
nand U803 (N_803,N_757,N_759);
nor U804 (N_804,N_766,N_786);
and U805 (N_805,N_793,N_775);
nor U806 (N_806,N_798,N_770);
or U807 (N_807,N_783,N_799);
nand U808 (N_808,N_771,N_765);
nand U809 (N_809,N_788,N_790);
and U810 (N_810,N_773,N_792);
or U811 (N_811,N_778,N_777);
and U812 (N_812,N_756,N_752);
or U813 (N_813,N_791,N_753);
or U814 (N_814,N_784,N_758);
and U815 (N_815,N_764,N_794);
nor U816 (N_816,N_750,N_780);
nor U817 (N_817,N_768,N_797);
or U818 (N_818,N_776,N_767);
xnor U819 (N_819,N_774,N_762);
and U820 (N_820,N_772,N_763);
nor U821 (N_821,N_785,N_789);
nand U822 (N_822,N_769,N_779);
and U823 (N_823,N_781,N_760);
or U824 (N_824,N_795,N_754);
and U825 (N_825,N_767,N_758);
nand U826 (N_826,N_783,N_772);
nor U827 (N_827,N_780,N_794);
and U828 (N_828,N_776,N_787);
or U829 (N_829,N_784,N_787);
nand U830 (N_830,N_769,N_789);
or U831 (N_831,N_798,N_780);
nand U832 (N_832,N_786,N_788);
and U833 (N_833,N_766,N_767);
and U834 (N_834,N_753,N_789);
or U835 (N_835,N_777,N_788);
and U836 (N_836,N_757,N_762);
or U837 (N_837,N_798,N_788);
and U838 (N_838,N_752,N_768);
or U839 (N_839,N_795,N_752);
or U840 (N_840,N_796,N_768);
or U841 (N_841,N_796,N_798);
or U842 (N_842,N_799,N_758);
nor U843 (N_843,N_769,N_751);
nand U844 (N_844,N_766,N_797);
or U845 (N_845,N_754,N_794);
nor U846 (N_846,N_770,N_788);
and U847 (N_847,N_777,N_759);
nor U848 (N_848,N_760,N_765);
xnor U849 (N_849,N_770,N_761);
nor U850 (N_850,N_845,N_823);
nor U851 (N_851,N_804,N_825);
nor U852 (N_852,N_835,N_829);
and U853 (N_853,N_808,N_830);
nand U854 (N_854,N_844,N_806);
or U855 (N_855,N_818,N_833);
and U856 (N_856,N_807,N_832);
or U857 (N_857,N_801,N_821);
nor U858 (N_858,N_816,N_838);
or U859 (N_859,N_809,N_817);
nor U860 (N_860,N_824,N_800);
nor U861 (N_861,N_805,N_813);
nor U862 (N_862,N_802,N_847);
nand U863 (N_863,N_827,N_837);
and U864 (N_864,N_820,N_803);
nand U865 (N_865,N_841,N_811);
and U866 (N_866,N_828,N_840);
or U867 (N_867,N_842,N_810);
nor U868 (N_868,N_819,N_839);
nand U869 (N_869,N_848,N_834);
and U870 (N_870,N_836,N_846);
nor U871 (N_871,N_815,N_849);
xor U872 (N_872,N_822,N_812);
and U873 (N_873,N_843,N_831);
nand U874 (N_874,N_826,N_814);
or U875 (N_875,N_845,N_803);
nand U876 (N_876,N_841,N_846);
nor U877 (N_877,N_837,N_823);
or U878 (N_878,N_819,N_815);
nor U879 (N_879,N_827,N_824);
nor U880 (N_880,N_838,N_811);
nand U881 (N_881,N_832,N_834);
or U882 (N_882,N_818,N_832);
or U883 (N_883,N_842,N_826);
nand U884 (N_884,N_826,N_802);
or U885 (N_885,N_809,N_818);
or U886 (N_886,N_844,N_818);
nor U887 (N_887,N_830,N_835);
nor U888 (N_888,N_827,N_814);
or U889 (N_889,N_847,N_822);
and U890 (N_890,N_802,N_808);
or U891 (N_891,N_810,N_822);
nor U892 (N_892,N_841,N_843);
nor U893 (N_893,N_842,N_849);
nand U894 (N_894,N_834,N_843);
or U895 (N_895,N_815,N_800);
or U896 (N_896,N_849,N_816);
nand U897 (N_897,N_812,N_827);
nand U898 (N_898,N_813,N_835);
or U899 (N_899,N_828,N_815);
nand U900 (N_900,N_860,N_855);
and U901 (N_901,N_890,N_861);
nand U902 (N_902,N_850,N_898);
or U903 (N_903,N_878,N_862);
and U904 (N_904,N_874,N_856);
nor U905 (N_905,N_859,N_864);
nand U906 (N_906,N_853,N_895);
and U907 (N_907,N_877,N_869);
nor U908 (N_908,N_894,N_893);
nand U909 (N_909,N_872,N_899);
and U910 (N_910,N_876,N_885);
nor U911 (N_911,N_863,N_880);
and U912 (N_912,N_854,N_897);
and U913 (N_913,N_851,N_867);
or U914 (N_914,N_857,N_875);
and U915 (N_915,N_881,N_888);
nor U916 (N_916,N_892,N_896);
xor U917 (N_917,N_873,N_889);
and U918 (N_918,N_891,N_870);
and U919 (N_919,N_886,N_868);
nor U920 (N_920,N_871,N_865);
and U921 (N_921,N_858,N_852);
and U922 (N_922,N_887,N_883);
nor U923 (N_923,N_879,N_884);
xnor U924 (N_924,N_866,N_882);
nand U925 (N_925,N_871,N_863);
and U926 (N_926,N_872,N_894);
nor U927 (N_927,N_857,N_853);
nor U928 (N_928,N_897,N_894);
xnor U929 (N_929,N_893,N_864);
and U930 (N_930,N_884,N_890);
or U931 (N_931,N_851,N_857);
and U932 (N_932,N_898,N_863);
nor U933 (N_933,N_890,N_898);
nor U934 (N_934,N_858,N_899);
and U935 (N_935,N_858,N_855);
nor U936 (N_936,N_885,N_896);
xor U937 (N_937,N_896,N_891);
and U938 (N_938,N_879,N_891);
and U939 (N_939,N_858,N_875);
and U940 (N_940,N_890,N_860);
nor U941 (N_941,N_880,N_874);
nor U942 (N_942,N_850,N_899);
nand U943 (N_943,N_877,N_863);
or U944 (N_944,N_893,N_853);
nand U945 (N_945,N_877,N_892);
nand U946 (N_946,N_885,N_861);
nand U947 (N_947,N_896,N_875);
nand U948 (N_948,N_862,N_853);
xnor U949 (N_949,N_889,N_862);
and U950 (N_950,N_913,N_939);
and U951 (N_951,N_934,N_942);
and U952 (N_952,N_938,N_925);
nor U953 (N_953,N_935,N_909);
nor U954 (N_954,N_923,N_941);
nand U955 (N_955,N_905,N_932);
xor U956 (N_956,N_922,N_904);
and U957 (N_957,N_949,N_928);
nor U958 (N_958,N_915,N_936);
nand U959 (N_959,N_926,N_927);
and U960 (N_960,N_947,N_900);
or U961 (N_961,N_920,N_914);
and U962 (N_962,N_911,N_921);
nor U963 (N_963,N_930,N_929);
and U964 (N_964,N_937,N_916);
nand U965 (N_965,N_901,N_948);
and U966 (N_966,N_931,N_918);
xnor U967 (N_967,N_912,N_903);
and U968 (N_968,N_919,N_924);
nor U969 (N_969,N_944,N_917);
nand U970 (N_970,N_945,N_933);
nor U971 (N_971,N_907,N_908);
nor U972 (N_972,N_943,N_902);
nor U973 (N_973,N_906,N_940);
and U974 (N_974,N_946,N_910);
nor U975 (N_975,N_906,N_913);
nor U976 (N_976,N_924,N_932);
nor U977 (N_977,N_927,N_908);
nand U978 (N_978,N_946,N_922);
nand U979 (N_979,N_942,N_936);
xor U980 (N_980,N_905,N_901);
and U981 (N_981,N_903,N_926);
xnor U982 (N_982,N_942,N_911);
or U983 (N_983,N_919,N_925);
nor U984 (N_984,N_914,N_911);
nor U985 (N_985,N_902,N_905);
and U986 (N_986,N_907,N_930);
nand U987 (N_987,N_944,N_948);
nor U988 (N_988,N_905,N_916);
or U989 (N_989,N_902,N_936);
nand U990 (N_990,N_922,N_915);
or U991 (N_991,N_931,N_949);
nand U992 (N_992,N_926,N_902);
nor U993 (N_993,N_902,N_928);
or U994 (N_994,N_914,N_902);
nand U995 (N_995,N_902,N_925);
and U996 (N_996,N_930,N_927);
nor U997 (N_997,N_945,N_928);
xor U998 (N_998,N_936,N_935);
and U999 (N_999,N_938,N_914);
and U1000 (N_1000,N_956,N_982);
or U1001 (N_1001,N_983,N_972);
and U1002 (N_1002,N_979,N_986);
nand U1003 (N_1003,N_955,N_962);
or U1004 (N_1004,N_976,N_954);
and U1005 (N_1005,N_988,N_980);
and U1006 (N_1006,N_987,N_951);
xnor U1007 (N_1007,N_991,N_993);
nand U1008 (N_1008,N_981,N_997);
and U1009 (N_1009,N_977,N_968);
nor U1010 (N_1010,N_999,N_966);
nand U1011 (N_1011,N_953,N_978);
and U1012 (N_1012,N_975,N_994);
nand U1013 (N_1013,N_958,N_952);
or U1014 (N_1014,N_974,N_961);
and U1015 (N_1015,N_965,N_989);
nand U1016 (N_1016,N_960,N_950);
nand U1017 (N_1017,N_971,N_990);
nand U1018 (N_1018,N_985,N_998);
nand U1019 (N_1019,N_957,N_967);
nor U1020 (N_1020,N_959,N_963);
nor U1021 (N_1021,N_973,N_969);
xor U1022 (N_1022,N_970,N_992);
nand U1023 (N_1023,N_964,N_984);
or U1024 (N_1024,N_995,N_996);
and U1025 (N_1025,N_955,N_977);
xnor U1026 (N_1026,N_979,N_970);
nand U1027 (N_1027,N_986,N_996);
and U1028 (N_1028,N_969,N_974);
xor U1029 (N_1029,N_994,N_954);
and U1030 (N_1030,N_998,N_999);
nand U1031 (N_1031,N_957,N_961);
and U1032 (N_1032,N_973,N_953);
or U1033 (N_1033,N_991,N_973);
or U1034 (N_1034,N_985,N_968);
or U1035 (N_1035,N_998,N_975);
and U1036 (N_1036,N_989,N_988);
or U1037 (N_1037,N_982,N_979);
or U1038 (N_1038,N_999,N_963);
and U1039 (N_1039,N_984,N_953);
or U1040 (N_1040,N_977,N_980);
or U1041 (N_1041,N_978,N_960);
nand U1042 (N_1042,N_995,N_971);
nand U1043 (N_1043,N_957,N_999);
nor U1044 (N_1044,N_991,N_954);
and U1045 (N_1045,N_955,N_985);
nand U1046 (N_1046,N_979,N_951);
nand U1047 (N_1047,N_950,N_989);
xor U1048 (N_1048,N_995,N_977);
nor U1049 (N_1049,N_991,N_979);
nor U1050 (N_1050,N_1015,N_1036);
or U1051 (N_1051,N_1049,N_1002);
and U1052 (N_1052,N_1018,N_1006);
nand U1053 (N_1053,N_1035,N_1027);
or U1054 (N_1054,N_1034,N_1009);
and U1055 (N_1055,N_1013,N_1022);
nor U1056 (N_1056,N_1019,N_1011);
nand U1057 (N_1057,N_1004,N_1029);
nor U1058 (N_1058,N_1014,N_1003);
or U1059 (N_1059,N_1039,N_1010);
and U1060 (N_1060,N_1020,N_1043);
and U1061 (N_1061,N_1024,N_1026);
and U1062 (N_1062,N_1048,N_1031);
nor U1063 (N_1063,N_1045,N_1028);
xor U1064 (N_1064,N_1000,N_1007);
nor U1065 (N_1065,N_1032,N_1030);
xor U1066 (N_1066,N_1041,N_1033);
nor U1067 (N_1067,N_1038,N_1025);
or U1068 (N_1068,N_1046,N_1037);
and U1069 (N_1069,N_1005,N_1021);
and U1070 (N_1070,N_1012,N_1023);
nor U1071 (N_1071,N_1042,N_1008);
or U1072 (N_1072,N_1047,N_1044);
or U1073 (N_1073,N_1001,N_1040);
xnor U1074 (N_1074,N_1016,N_1017);
or U1075 (N_1075,N_1005,N_1034);
xor U1076 (N_1076,N_1037,N_1032);
or U1077 (N_1077,N_1034,N_1001);
xor U1078 (N_1078,N_1016,N_1020);
nor U1079 (N_1079,N_1014,N_1007);
or U1080 (N_1080,N_1043,N_1038);
and U1081 (N_1081,N_1008,N_1013);
or U1082 (N_1082,N_1020,N_1046);
nor U1083 (N_1083,N_1046,N_1030);
nand U1084 (N_1084,N_1043,N_1039);
nor U1085 (N_1085,N_1027,N_1038);
nand U1086 (N_1086,N_1021,N_1001);
and U1087 (N_1087,N_1025,N_1026);
xnor U1088 (N_1088,N_1032,N_1009);
nor U1089 (N_1089,N_1022,N_1045);
xnor U1090 (N_1090,N_1038,N_1020);
nor U1091 (N_1091,N_1016,N_1022);
or U1092 (N_1092,N_1033,N_1017);
and U1093 (N_1093,N_1003,N_1024);
nor U1094 (N_1094,N_1037,N_1049);
nor U1095 (N_1095,N_1007,N_1011);
nor U1096 (N_1096,N_1001,N_1013);
nor U1097 (N_1097,N_1015,N_1017);
nor U1098 (N_1098,N_1000,N_1040);
nand U1099 (N_1099,N_1044,N_1038);
or U1100 (N_1100,N_1059,N_1068);
nor U1101 (N_1101,N_1088,N_1052);
or U1102 (N_1102,N_1074,N_1076);
nand U1103 (N_1103,N_1055,N_1053);
and U1104 (N_1104,N_1064,N_1083);
and U1105 (N_1105,N_1063,N_1072);
nor U1106 (N_1106,N_1082,N_1092);
xnor U1107 (N_1107,N_1073,N_1098);
or U1108 (N_1108,N_1070,N_1080);
nand U1109 (N_1109,N_1077,N_1084);
nand U1110 (N_1110,N_1051,N_1086);
and U1111 (N_1111,N_1060,N_1095);
nand U1112 (N_1112,N_1094,N_1079);
or U1113 (N_1113,N_1056,N_1099);
nand U1114 (N_1114,N_1057,N_1067);
nor U1115 (N_1115,N_1061,N_1058);
or U1116 (N_1116,N_1096,N_1085);
and U1117 (N_1117,N_1090,N_1071);
nand U1118 (N_1118,N_1087,N_1054);
and U1119 (N_1119,N_1069,N_1081);
nor U1120 (N_1120,N_1089,N_1097);
and U1121 (N_1121,N_1050,N_1091);
xnor U1122 (N_1122,N_1093,N_1066);
and U1123 (N_1123,N_1075,N_1078);
nor U1124 (N_1124,N_1065,N_1062);
nor U1125 (N_1125,N_1089,N_1067);
or U1126 (N_1126,N_1092,N_1095);
and U1127 (N_1127,N_1068,N_1052);
nor U1128 (N_1128,N_1061,N_1059);
nand U1129 (N_1129,N_1059,N_1071);
nand U1130 (N_1130,N_1084,N_1052);
or U1131 (N_1131,N_1078,N_1083);
and U1132 (N_1132,N_1054,N_1050);
nand U1133 (N_1133,N_1068,N_1085);
xor U1134 (N_1134,N_1057,N_1085);
nand U1135 (N_1135,N_1082,N_1095);
and U1136 (N_1136,N_1069,N_1091);
nor U1137 (N_1137,N_1079,N_1057);
nor U1138 (N_1138,N_1054,N_1056);
nor U1139 (N_1139,N_1050,N_1094);
nand U1140 (N_1140,N_1087,N_1083);
and U1141 (N_1141,N_1075,N_1096);
nor U1142 (N_1142,N_1074,N_1070);
nor U1143 (N_1143,N_1085,N_1072);
nand U1144 (N_1144,N_1097,N_1054);
nand U1145 (N_1145,N_1086,N_1066);
and U1146 (N_1146,N_1061,N_1091);
or U1147 (N_1147,N_1089,N_1075);
nor U1148 (N_1148,N_1097,N_1073);
nand U1149 (N_1149,N_1067,N_1087);
nand U1150 (N_1150,N_1132,N_1123);
or U1151 (N_1151,N_1142,N_1114);
nor U1152 (N_1152,N_1147,N_1116);
and U1153 (N_1153,N_1122,N_1148);
nor U1154 (N_1154,N_1135,N_1104);
or U1155 (N_1155,N_1115,N_1106);
or U1156 (N_1156,N_1102,N_1100);
and U1157 (N_1157,N_1144,N_1131);
or U1158 (N_1158,N_1141,N_1127);
or U1159 (N_1159,N_1140,N_1124);
and U1160 (N_1160,N_1105,N_1101);
nand U1161 (N_1161,N_1130,N_1121);
or U1162 (N_1162,N_1134,N_1129);
nand U1163 (N_1163,N_1109,N_1118);
nor U1164 (N_1164,N_1136,N_1128);
or U1165 (N_1165,N_1138,N_1125);
nand U1166 (N_1166,N_1137,N_1107);
xor U1167 (N_1167,N_1112,N_1146);
nor U1168 (N_1168,N_1139,N_1117);
xnor U1169 (N_1169,N_1145,N_1120);
or U1170 (N_1170,N_1143,N_1119);
or U1171 (N_1171,N_1126,N_1113);
nor U1172 (N_1172,N_1133,N_1110);
and U1173 (N_1173,N_1103,N_1149);
and U1174 (N_1174,N_1108,N_1111);
or U1175 (N_1175,N_1148,N_1112);
xnor U1176 (N_1176,N_1108,N_1146);
nand U1177 (N_1177,N_1111,N_1127);
nand U1178 (N_1178,N_1125,N_1136);
or U1179 (N_1179,N_1143,N_1142);
nor U1180 (N_1180,N_1122,N_1115);
nor U1181 (N_1181,N_1133,N_1100);
or U1182 (N_1182,N_1121,N_1142);
nand U1183 (N_1183,N_1142,N_1102);
nand U1184 (N_1184,N_1128,N_1110);
and U1185 (N_1185,N_1127,N_1122);
nor U1186 (N_1186,N_1130,N_1122);
and U1187 (N_1187,N_1147,N_1141);
or U1188 (N_1188,N_1142,N_1144);
and U1189 (N_1189,N_1139,N_1122);
nor U1190 (N_1190,N_1130,N_1125);
or U1191 (N_1191,N_1137,N_1119);
or U1192 (N_1192,N_1130,N_1111);
nand U1193 (N_1193,N_1103,N_1132);
and U1194 (N_1194,N_1130,N_1109);
nor U1195 (N_1195,N_1146,N_1113);
nand U1196 (N_1196,N_1133,N_1123);
nand U1197 (N_1197,N_1107,N_1123);
and U1198 (N_1198,N_1142,N_1148);
and U1199 (N_1199,N_1120,N_1122);
or U1200 (N_1200,N_1176,N_1168);
nand U1201 (N_1201,N_1165,N_1191);
and U1202 (N_1202,N_1167,N_1195);
nand U1203 (N_1203,N_1158,N_1186);
nand U1204 (N_1204,N_1190,N_1183);
or U1205 (N_1205,N_1198,N_1187);
xnor U1206 (N_1206,N_1179,N_1196);
and U1207 (N_1207,N_1159,N_1163);
or U1208 (N_1208,N_1197,N_1169);
and U1209 (N_1209,N_1175,N_1152);
or U1210 (N_1210,N_1178,N_1188);
xnor U1211 (N_1211,N_1173,N_1182);
nand U1212 (N_1212,N_1164,N_1151);
nor U1213 (N_1213,N_1166,N_1185);
xnor U1214 (N_1214,N_1153,N_1194);
or U1215 (N_1215,N_1199,N_1177);
nor U1216 (N_1216,N_1192,N_1150);
nand U1217 (N_1217,N_1189,N_1157);
nand U1218 (N_1218,N_1174,N_1193);
nand U1219 (N_1219,N_1154,N_1162);
nor U1220 (N_1220,N_1160,N_1161);
and U1221 (N_1221,N_1155,N_1171);
or U1222 (N_1222,N_1170,N_1172);
or U1223 (N_1223,N_1184,N_1180);
nand U1224 (N_1224,N_1181,N_1156);
and U1225 (N_1225,N_1163,N_1196);
and U1226 (N_1226,N_1175,N_1183);
nor U1227 (N_1227,N_1169,N_1153);
nor U1228 (N_1228,N_1181,N_1157);
and U1229 (N_1229,N_1197,N_1193);
nand U1230 (N_1230,N_1155,N_1188);
nor U1231 (N_1231,N_1155,N_1150);
nor U1232 (N_1232,N_1154,N_1152);
nor U1233 (N_1233,N_1186,N_1181);
or U1234 (N_1234,N_1183,N_1172);
or U1235 (N_1235,N_1185,N_1161);
or U1236 (N_1236,N_1150,N_1152);
or U1237 (N_1237,N_1154,N_1177);
and U1238 (N_1238,N_1172,N_1177);
nand U1239 (N_1239,N_1161,N_1150);
or U1240 (N_1240,N_1161,N_1194);
and U1241 (N_1241,N_1164,N_1193);
nor U1242 (N_1242,N_1192,N_1181);
nand U1243 (N_1243,N_1184,N_1156);
nand U1244 (N_1244,N_1161,N_1199);
nor U1245 (N_1245,N_1179,N_1156);
or U1246 (N_1246,N_1161,N_1152);
and U1247 (N_1247,N_1189,N_1193);
or U1248 (N_1248,N_1179,N_1189);
nor U1249 (N_1249,N_1160,N_1165);
and U1250 (N_1250,N_1218,N_1247);
nand U1251 (N_1251,N_1203,N_1242);
and U1252 (N_1252,N_1243,N_1220);
and U1253 (N_1253,N_1236,N_1231);
nor U1254 (N_1254,N_1208,N_1249);
nor U1255 (N_1255,N_1234,N_1221);
nor U1256 (N_1256,N_1230,N_1202);
and U1257 (N_1257,N_1211,N_1226);
and U1258 (N_1258,N_1240,N_1206);
xor U1259 (N_1259,N_1212,N_1214);
or U1260 (N_1260,N_1224,N_1229);
and U1261 (N_1261,N_1239,N_1235);
or U1262 (N_1262,N_1216,N_1225);
or U1263 (N_1263,N_1200,N_1210);
and U1264 (N_1264,N_1237,N_1248);
nand U1265 (N_1265,N_1215,N_1233);
nor U1266 (N_1266,N_1232,N_1209);
or U1267 (N_1267,N_1244,N_1219);
or U1268 (N_1268,N_1204,N_1213);
nor U1269 (N_1269,N_1227,N_1223);
xnor U1270 (N_1270,N_1245,N_1217);
xor U1271 (N_1271,N_1222,N_1207);
and U1272 (N_1272,N_1246,N_1238);
and U1273 (N_1273,N_1201,N_1205);
nand U1274 (N_1274,N_1228,N_1241);
and U1275 (N_1275,N_1201,N_1243);
nor U1276 (N_1276,N_1209,N_1249);
nor U1277 (N_1277,N_1248,N_1218);
nand U1278 (N_1278,N_1245,N_1220);
nand U1279 (N_1279,N_1244,N_1231);
or U1280 (N_1280,N_1236,N_1243);
nand U1281 (N_1281,N_1244,N_1226);
or U1282 (N_1282,N_1212,N_1243);
nor U1283 (N_1283,N_1222,N_1239);
nand U1284 (N_1284,N_1245,N_1209);
and U1285 (N_1285,N_1247,N_1221);
nor U1286 (N_1286,N_1239,N_1213);
and U1287 (N_1287,N_1224,N_1242);
nand U1288 (N_1288,N_1223,N_1213);
and U1289 (N_1289,N_1226,N_1213);
nor U1290 (N_1290,N_1234,N_1225);
and U1291 (N_1291,N_1247,N_1203);
and U1292 (N_1292,N_1229,N_1202);
or U1293 (N_1293,N_1243,N_1203);
nor U1294 (N_1294,N_1228,N_1210);
nor U1295 (N_1295,N_1210,N_1215);
or U1296 (N_1296,N_1241,N_1217);
or U1297 (N_1297,N_1214,N_1209);
nor U1298 (N_1298,N_1244,N_1245);
or U1299 (N_1299,N_1200,N_1228);
nor U1300 (N_1300,N_1285,N_1269);
and U1301 (N_1301,N_1298,N_1268);
and U1302 (N_1302,N_1291,N_1296);
and U1303 (N_1303,N_1282,N_1284);
and U1304 (N_1304,N_1265,N_1255);
nor U1305 (N_1305,N_1274,N_1290);
nor U1306 (N_1306,N_1256,N_1280);
nor U1307 (N_1307,N_1281,N_1266);
nor U1308 (N_1308,N_1275,N_1258);
and U1309 (N_1309,N_1287,N_1270);
nor U1310 (N_1310,N_1264,N_1279);
nor U1311 (N_1311,N_1289,N_1286);
and U1312 (N_1312,N_1261,N_1263);
nor U1313 (N_1313,N_1253,N_1283);
or U1314 (N_1314,N_1260,N_1250);
nor U1315 (N_1315,N_1251,N_1288);
nand U1316 (N_1316,N_1297,N_1267);
or U1317 (N_1317,N_1262,N_1278);
or U1318 (N_1318,N_1277,N_1257);
and U1319 (N_1319,N_1292,N_1272);
nor U1320 (N_1320,N_1252,N_1295);
or U1321 (N_1321,N_1276,N_1271);
and U1322 (N_1322,N_1293,N_1254);
or U1323 (N_1323,N_1273,N_1294);
nand U1324 (N_1324,N_1259,N_1299);
nor U1325 (N_1325,N_1274,N_1256);
or U1326 (N_1326,N_1254,N_1261);
and U1327 (N_1327,N_1296,N_1297);
and U1328 (N_1328,N_1296,N_1294);
nor U1329 (N_1329,N_1256,N_1258);
or U1330 (N_1330,N_1289,N_1282);
or U1331 (N_1331,N_1255,N_1271);
nand U1332 (N_1332,N_1278,N_1280);
nand U1333 (N_1333,N_1288,N_1267);
nor U1334 (N_1334,N_1284,N_1276);
or U1335 (N_1335,N_1283,N_1280);
nand U1336 (N_1336,N_1254,N_1250);
xor U1337 (N_1337,N_1284,N_1266);
and U1338 (N_1338,N_1284,N_1261);
or U1339 (N_1339,N_1290,N_1284);
nor U1340 (N_1340,N_1272,N_1282);
and U1341 (N_1341,N_1284,N_1299);
and U1342 (N_1342,N_1250,N_1278);
or U1343 (N_1343,N_1281,N_1299);
nor U1344 (N_1344,N_1271,N_1266);
xnor U1345 (N_1345,N_1277,N_1250);
nor U1346 (N_1346,N_1274,N_1270);
nor U1347 (N_1347,N_1288,N_1299);
and U1348 (N_1348,N_1257,N_1281);
nand U1349 (N_1349,N_1292,N_1297);
nor U1350 (N_1350,N_1341,N_1340);
or U1351 (N_1351,N_1301,N_1316);
nand U1352 (N_1352,N_1305,N_1300);
or U1353 (N_1353,N_1317,N_1331);
nor U1354 (N_1354,N_1324,N_1339);
and U1355 (N_1355,N_1335,N_1312);
or U1356 (N_1356,N_1322,N_1320);
nand U1357 (N_1357,N_1303,N_1309);
nor U1358 (N_1358,N_1310,N_1304);
and U1359 (N_1359,N_1315,N_1349);
nor U1360 (N_1360,N_1325,N_1342);
or U1361 (N_1361,N_1306,N_1323);
nor U1362 (N_1362,N_1314,N_1327);
nor U1363 (N_1363,N_1308,N_1336);
nand U1364 (N_1364,N_1347,N_1329);
nor U1365 (N_1365,N_1348,N_1345);
and U1366 (N_1366,N_1326,N_1346);
or U1367 (N_1367,N_1344,N_1328);
nand U1368 (N_1368,N_1319,N_1307);
and U1369 (N_1369,N_1313,N_1330);
and U1370 (N_1370,N_1318,N_1333);
or U1371 (N_1371,N_1338,N_1302);
and U1372 (N_1372,N_1337,N_1311);
nand U1373 (N_1373,N_1343,N_1321);
nand U1374 (N_1374,N_1332,N_1334);
nand U1375 (N_1375,N_1345,N_1325);
nor U1376 (N_1376,N_1341,N_1338);
nor U1377 (N_1377,N_1327,N_1300);
and U1378 (N_1378,N_1334,N_1339);
nand U1379 (N_1379,N_1313,N_1319);
nor U1380 (N_1380,N_1311,N_1313);
or U1381 (N_1381,N_1313,N_1340);
or U1382 (N_1382,N_1331,N_1332);
or U1383 (N_1383,N_1338,N_1330);
or U1384 (N_1384,N_1325,N_1347);
or U1385 (N_1385,N_1309,N_1324);
nand U1386 (N_1386,N_1344,N_1305);
nor U1387 (N_1387,N_1337,N_1345);
or U1388 (N_1388,N_1305,N_1313);
and U1389 (N_1389,N_1322,N_1332);
nor U1390 (N_1390,N_1337,N_1336);
and U1391 (N_1391,N_1345,N_1330);
nand U1392 (N_1392,N_1314,N_1336);
and U1393 (N_1393,N_1321,N_1310);
nor U1394 (N_1394,N_1328,N_1326);
nor U1395 (N_1395,N_1332,N_1314);
nor U1396 (N_1396,N_1304,N_1337);
nand U1397 (N_1397,N_1349,N_1328);
and U1398 (N_1398,N_1315,N_1335);
or U1399 (N_1399,N_1306,N_1301);
and U1400 (N_1400,N_1358,N_1350);
or U1401 (N_1401,N_1357,N_1370);
nor U1402 (N_1402,N_1353,N_1392);
or U1403 (N_1403,N_1371,N_1394);
and U1404 (N_1404,N_1379,N_1351);
nand U1405 (N_1405,N_1359,N_1352);
nand U1406 (N_1406,N_1363,N_1395);
nand U1407 (N_1407,N_1373,N_1377);
and U1408 (N_1408,N_1381,N_1388);
nor U1409 (N_1409,N_1393,N_1355);
or U1410 (N_1410,N_1367,N_1354);
or U1411 (N_1411,N_1383,N_1375);
nor U1412 (N_1412,N_1356,N_1368);
nor U1413 (N_1413,N_1399,N_1397);
and U1414 (N_1414,N_1387,N_1361);
nand U1415 (N_1415,N_1360,N_1366);
nand U1416 (N_1416,N_1398,N_1364);
nor U1417 (N_1417,N_1386,N_1396);
and U1418 (N_1418,N_1384,N_1385);
xnor U1419 (N_1419,N_1380,N_1374);
and U1420 (N_1420,N_1389,N_1365);
nor U1421 (N_1421,N_1369,N_1376);
or U1422 (N_1422,N_1378,N_1382);
and U1423 (N_1423,N_1362,N_1391);
or U1424 (N_1424,N_1390,N_1372);
and U1425 (N_1425,N_1354,N_1372);
and U1426 (N_1426,N_1399,N_1366);
nor U1427 (N_1427,N_1363,N_1364);
nand U1428 (N_1428,N_1381,N_1390);
and U1429 (N_1429,N_1395,N_1354);
nor U1430 (N_1430,N_1357,N_1358);
nand U1431 (N_1431,N_1396,N_1361);
nand U1432 (N_1432,N_1381,N_1395);
nor U1433 (N_1433,N_1387,N_1357);
and U1434 (N_1434,N_1363,N_1357);
nand U1435 (N_1435,N_1374,N_1369);
xnor U1436 (N_1436,N_1382,N_1386);
nand U1437 (N_1437,N_1376,N_1379);
nor U1438 (N_1438,N_1376,N_1362);
nor U1439 (N_1439,N_1360,N_1378);
and U1440 (N_1440,N_1396,N_1384);
nor U1441 (N_1441,N_1359,N_1371);
nand U1442 (N_1442,N_1379,N_1372);
nand U1443 (N_1443,N_1389,N_1394);
nand U1444 (N_1444,N_1387,N_1371);
or U1445 (N_1445,N_1381,N_1372);
and U1446 (N_1446,N_1363,N_1374);
nor U1447 (N_1447,N_1357,N_1374);
xor U1448 (N_1448,N_1372,N_1363);
nand U1449 (N_1449,N_1396,N_1390);
nand U1450 (N_1450,N_1413,N_1437);
and U1451 (N_1451,N_1444,N_1414);
nand U1452 (N_1452,N_1426,N_1425);
or U1453 (N_1453,N_1448,N_1420);
nand U1454 (N_1454,N_1441,N_1400);
xnor U1455 (N_1455,N_1438,N_1412);
or U1456 (N_1456,N_1443,N_1418);
or U1457 (N_1457,N_1449,N_1442);
or U1458 (N_1458,N_1405,N_1416);
nand U1459 (N_1459,N_1434,N_1432);
nand U1460 (N_1460,N_1430,N_1423);
or U1461 (N_1461,N_1403,N_1404);
and U1462 (N_1462,N_1415,N_1446);
nor U1463 (N_1463,N_1411,N_1427);
or U1464 (N_1464,N_1439,N_1440);
nor U1465 (N_1465,N_1424,N_1410);
nand U1466 (N_1466,N_1406,N_1436);
and U1467 (N_1467,N_1402,N_1429);
and U1468 (N_1468,N_1419,N_1428);
nand U1469 (N_1469,N_1431,N_1407);
or U1470 (N_1470,N_1447,N_1409);
or U1471 (N_1471,N_1421,N_1417);
nand U1472 (N_1472,N_1408,N_1433);
and U1473 (N_1473,N_1445,N_1422);
or U1474 (N_1474,N_1401,N_1435);
nand U1475 (N_1475,N_1425,N_1411);
or U1476 (N_1476,N_1435,N_1430);
nand U1477 (N_1477,N_1447,N_1421);
nor U1478 (N_1478,N_1412,N_1402);
nand U1479 (N_1479,N_1443,N_1429);
nand U1480 (N_1480,N_1435,N_1400);
and U1481 (N_1481,N_1403,N_1420);
or U1482 (N_1482,N_1410,N_1445);
nand U1483 (N_1483,N_1418,N_1411);
or U1484 (N_1484,N_1431,N_1418);
nor U1485 (N_1485,N_1446,N_1400);
nor U1486 (N_1486,N_1414,N_1436);
nor U1487 (N_1487,N_1406,N_1408);
nor U1488 (N_1488,N_1449,N_1445);
and U1489 (N_1489,N_1429,N_1415);
or U1490 (N_1490,N_1401,N_1426);
and U1491 (N_1491,N_1440,N_1442);
nand U1492 (N_1492,N_1404,N_1417);
nor U1493 (N_1493,N_1441,N_1424);
nor U1494 (N_1494,N_1403,N_1417);
and U1495 (N_1495,N_1403,N_1426);
nor U1496 (N_1496,N_1443,N_1407);
or U1497 (N_1497,N_1413,N_1424);
and U1498 (N_1498,N_1441,N_1447);
and U1499 (N_1499,N_1435,N_1415);
or U1500 (N_1500,N_1463,N_1462);
or U1501 (N_1501,N_1497,N_1473);
nand U1502 (N_1502,N_1478,N_1456);
or U1503 (N_1503,N_1458,N_1453);
nand U1504 (N_1504,N_1452,N_1476);
nand U1505 (N_1505,N_1469,N_1466);
or U1506 (N_1506,N_1494,N_1482);
and U1507 (N_1507,N_1459,N_1479);
nor U1508 (N_1508,N_1499,N_1495);
and U1509 (N_1509,N_1488,N_1471);
nand U1510 (N_1510,N_1496,N_1461);
or U1511 (N_1511,N_1490,N_1454);
nor U1512 (N_1512,N_1489,N_1485);
nor U1513 (N_1513,N_1470,N_1481);
and U1514 (N_1514,N_1468,N_1492);
or U1515 (N_1515,N_1451,N_1484);
or U1516 (N_1516,N_1493,N_1487);
and U1517 (N_1517,N_1460,N_1450);
nor U1518 (N_1518,N_1477,N_1498);
nor U1519 (N_1519,N_1486,N_1472);
nand U1520 (N_1520,N_1475,N_1465);
nand U1521 (N_1521,N_1491,N_1483);
or U1522 (N_1522,N_1474,N_1457);
nor U1523 (N_1523,N_1455,N_1464);
nor U1524 (N_1524,N_1480,N_1467);
or U1525 (N_1525,N_1463,N_1499);
nand U1526 (N_1526,N_1463,N_1497);
nor U1527 (N_1527,N_1488,N_1472);
and U1528 (N_1528,N_1467,N_1455);
nand U1529 (N_1529,N_1489,N_1450);
and U1530 (N_1530,N_1454,N_1477);
and U1531 (N_1531,N_1469,N_1475);
nand U1532 (N_1532,N_1452,N_1472);
and U1533 (N_1533,N_1488,N_1459);
nor U1534 (N_1534,N_1464,N_1493);
or U1535 (N_1535,N_1482,N_1455);
and U1536 (N_1536,N_1464,N_1477);
nor U1537 (N_1537,N_1485,N_1477);
nor U1538 (N_1538,N_1474,N_1493);
xor U1539 (N_1539,N_1455,N_1468);
and U1540 (N_1540,N_1499,N_1469);
nor U1541 (N_1541,N_1456,N_1467);
xnor U1542 (N_1542,N_1458,N_1482);
or U1543 (N_1543,N_1490,N_1462);
xnor U1544 (N_1544,N_1494,N_1471);
nand U1545 (N_1545,N_1495,N_1456);
nor U1546 (N_1546,N_1463,N_1468);
or U1547 (N_1547,N_1465,N_1488);
and U1548 (N_1548,N_1468,N_1458);
and U1549 (N_1549,N_1458,N_1465);
nand U1550 (N_1550,N_1534,N_1517);
and U1551 (N_1551,N_1537,N_1535);
nor U1552 (N_1552,N_1541,N_1549);
or U1553 (N_1553,N_1547,N_1533);
nand U1554 (N_1554,N_1536,N_1505);
or U1555 (N_1555,N_1512,N_1542);
nor U1556 (N_1556,N_1546,N_1519);
or U1557 (N_1557,N_1529,N_1525);
xor U1558 (N_1558,N_1510,N_1509);
nor U1559 (N_1559,N_1518,N_1545);
xnor U1560 (N_1560,N_1520,N_1524);
and U1561 (N_1561,N_1504,N_1530);
and U1562 (N_1562,N_1526,N_1539);
nor U1563 (N_1563,N_1513,N_1528);
nand U1564 (N_1564,N_1506,N_1523);
nor U1565 (N_1565,N_1516,N_1515);
nand U1566 (N_1566,N_1521,N_1527);
nand U1567 (N_1567,N_1532,N_1538);
xor U1568 (N_1568,N_1500,N_1544);
or U1569 (N_1569,N_1540,N_1501);
and U1570 (N_1570,N_1548,N_1511);
and U1571 (N_1571,N_1522,N_1507);
nor U1572 (N_1572,N_1508,N_1503);
nand U1573 (N_1573,N_1543,N_1514);
and U1574 (N_1574,N_1502,N_1531);
and U1575 (N_1575,N_1518,N_1515);
nand U1576 (N_1576,N_1506,N_1546);
or U1577 (N_1577,N_1505,N_1525);
or U1578 (N_1578,N_1519,N_1525);
xor U1579 (N_1579,N_1549,N_1525);
or U1580 (N_1580,N_1517,N_1525);
or U1581 (N_1581,N_1503,N_1509);
and U1582 (N_1582,N_1516,N_1527);
nand U1583 (N_1583,N_1529,N_1534);
and U1584 (N_1584,N_1516,N_1528);
and U1585 (N_1585,N_1546,N_1537);
nor U1586 (N_1586,N_1531,N_1549);
nor U1587 (N_1587,N_1527,N_1512);
or U1588 (N_1588,N_1549,N_1527);
and U1589 (N_1589,N_1531,N_1527);
or U1590 (N_1590,N_1509,N_1508);
or U1591 (N_1591,N_1528,N_1514);
or U1592 (N_1592,N_1538,N_1529);
or U1593 (N_1593,N_1525,N_1544);
nor U1594 (N_1594,N_1501,N_1549);
nand U1595 (N_1595,N_1520,N_1531);
or U1596 (N_1596,N_1519,N_1528);
nand U1597 (N_1597,N_1512,N_1546);
nand U1598 (N_1598,N_1523,N_1516);
nor U1599 (N_1599,N_1500,N_1530);
nor U1600 (N_1600,N_1557,N_1595);
nand U1601 (N_1601,N_1562,N_1575);
and U1602 (N_1602,N_1580,N_1555);
nor U1603 (N_1603,N_1553,N_1570);
nand U1604 (N_1604,N_1567,N_1589);
nand U1605 (N_1605,N_1594,N_1585);
and U1606 (N_1606,N_1566,N_1591);
nand U1607 (N_1607,N_1552,N_1560);
or U1608 (N_1608,N_1583,N_1597);
and U1609 (N_1609,N_1590,N_1568);
nor U1610 (N_1610,N_1587,N_1579);
nor U1611 (N_1611,N_1573,N_1565);
nand U1612 (N_1612,N_1550,N_1584);
or U1613 (N_1613,N_1569,N_1564);
xnor U1614 (N_1614,N_1588,N_1551);
nand U1615 (N_1615,N_1581,N_1558);
or U1616 (N_1616,N_1582,N_1593);
nor U1617 (N_1617,N_1554,N_1559);
nor U1618 (N_1618,N_1596,N_1592);
or U1619 (N_1619,N_1576,N_1586);
xor U1620 (N_1620,N_1599,N_1574);
nor U1621 (N_1621,N_1556,N_1561);
nor U1622 (N_1622,N_1578,N_1563);
nor U1623 (N_1623,N_1571,N_1598);
nand U1624 (N_1624,N_1577,N_1572);
or U1625 (N_1625,N_1578,N_1587);
or U1626 (N_1626,N_1596,N_1590);
xor U1627 (N_1627,N_1567,N_1598);
nand U1628 (N_1628,N_1586,N_1562);
nand U1629 (N_1629,N_1589,N_1571);
or U1630 (N_1630,N_1599,N_1552);
nand U1631 (N_1631,N_1569,N_1559);
nor U1632 (N_1632,N_1578,N_1571);
or U1633 (N_1633,N_1595,N_1575);
and U1634 (N_1634,N_1571,N_1588);
nor U1635 (N_1635,N_1571,N_1590);
nor U1636 (N_1636,N_1570,N_1575);
nand U1637 (N_1637,N_1554,N_1596);
xnor U1638 (N_1638,N_1576,N_1594);
nand U1639 (N_1639,N_1580,N_1581);
and U1640 (N_1640,N_1579,N_1580);
and U1641 (N_1641,N_1599,N_1567);
or U1642 (N_1642,N_1587,N_1591);
nand U1643 (N_1643,N_1581,N_1575);
and U1644 (N_1644,N_1553,N_1579);
or U1645 (N_1645,N_1561,N_1562);
or U1646 (N_1646,N_1595,N_1587);
or U1647 (N_1647,N_1580,N_1589);
nor U1648 (N_1648,N_1571,N_1567);
nand U1649 (N_1649,N_1550,N_1594);
nand U1650 (N_1650,N_1610,N_1613);
nand U1651 (N_1651,N_1606,N_1620);
nand U1652 (N_1652,N_1635,N_1623);
or U1653 (N_1653,N_1619,N_1636);
and U1654 (N_1654,N_1642,N_1605);
nand U1655 (N_1655,N_1624,N_1645);
or U1656 (N_1656,N_1600,N_1646);
nand U1657 (N_1657,N_1633,N_1618);
nor U1658 (N_1658,N_1641,N_1629);
and U1659 (N_1659,N_1615,N_1612);
or U1660 (N_1660,N_1643,N_1617);
nand U1661 (N_1661,N_1637,N_1627);
nor U1662 (N_1662,N_1634,N_1622);
or U1663 (N_1663,N_1602,N_1614);
or U1664 (N_1664,N_1631,N_1647);
xor U1665 (N_1665,N_1603,N_1604);
or U1666 (N_1666,N_1607,N_1601);
and U1667 (N_1667,N_1628,N_1649);
or U1668 (N_1668,N_1639,N_1638);
or U1669 (N_1669,N_1640,N_1648);
and U1670 (N_1670,N_1616,N_1630);
nand U1671 (N_1671,N_1608,N_1611);
nor U1672 (N_1672,N_1621,N_1609);
xnor U1673 (N_1673,N_1644,N_1625);
nor U1674 (N_1674,N_1626,N_1632);
and U1675 (N_1675,N_1606,N_1633);
nor U1676 (N_1676,N_1625,N_1619);
and U1677 (N_1677,N_1614,N_1629);
nor U1678 (N_1678,N_1608,N_1621);
nor U1679 (N_1679,N_1633,N_1644);
nor U1680 (N_1680,N_1616,N_1643);
or U1681 (N_1681,N_1607,N_1600);
or U1682 (N_1682,N_1618,N_1606);
nor U1683 (N_1683,N_1637,N_1602);
nand U1684 (N_1684,N_1600,N_1635);
nor U1685 (N_1685,N_1600,N_1632);
nor U1686 (N_1686,N_1606,N_1643);
nor U1687 (N_1687,N_1636,N_1649);
and U1688 (N_1688,N_1629,N_1600);
nand U1689 (N_1689,N_1636,N_1633);
or U1690 (N_1690,N_1608,N_1648);
or U1691 (N_1691,N_1613,N_1627);
or U1692 (N_1692,N_1644,N_1616);
or U1693 (N_1693,N_1628,N_1626);
nand U1694 (N_1694,N_1641,N_1624);
and U1695 (N_1695,N_1600,N_1638);
nor U1696 (N_1696,N_1624,N_1633);
or U1697 (N_1697,N_1615,N_1622);
nand U1698 (N_1698,N_1632,N_1641);
and U1699 (N_1699,N_1638,N_1629);
and U1700 (N_1700,N_1688,N_1663);
and U1701 (N_1701,N_1676,N_1695);
or U1702 (N_1702,N_1696,N_1698);
or U1703 (N_1703,N_1658,N_1683);
or U1704 (N_1704,N_1678,N_1664);
nor U1705 (N_1705,N_1662,N_1684);
nand U1706 (N_1706,N_1656,N_1655);
and U1707 (N_1707,N_1668,N_1677);
nand U1708 (N_1708,N_1650,N_1682);
or U1709 (N_1709,N_1681,N_1653);
and U1710 (N_1710,N_1675,N_1661);
or U1711 (N_1711,N_1657,N_1651);
or U1712 (N_1712,N_1665,N_1692);
and U1713 (N_1713,N_1679,N_1667);
nor U1714 (N_1714,N_1686,N_1659);
and U1715 (N_1715,N_1671,N_1673);
or U1716 (N_1716,N_1690,N_1687);
nand U1717 (N_1717,N_1652,N_1654);
or U1718 (N_1718,N_1685,N_1699);
nand U1719 (N_1719,N_1666,N_1680);
or U1720 (N_1720,N_1672,N_1694);
nand U1721 (N_1721,N_1693,N_1674);
nor U1722 (N_1722,N_1669,N_1670);
or U1723 (N_1723,N_1697,N_1691);
or U1724 (N_1724,N_1689,N_1660);
or U1725 (N_1725,N_1671,N_1653);
nand U1726 (N_1726,N_1681,N_1684);
or U1727 (N_1727,N_1683,N_1676);
nand U1728 (N_1728,N_1657,N_1655);
and U1729 (N_1729,N_1668,N_1689);
nor U1730 (N_1730,N_1694,N_1654);
xnor U1731 (N_1731,N_1657,N_1698);
or U1732 (N_1732,N_1696,N_1656);
and U1733 (N_1733,N_1653,N_1650);
and U1734 (N_1734,N_1675,N_1668);
nor U1735 (N_1735,N_1663,N_1665);
nor U1736 (N_1736,N_1675,N_1695);
nor U1737 (N_1737,N_1664,N_1690);
nand U1738 (N_1738,N_1680,N_1667);
and U1739 (N_1739,N_1657,N_1690);
nor U1740 (N_1740,N_1672,N_1688);
nor U1741 (N_1741,N_1677,N_1698);
nand U1742 (N_1742,N_1664,N_1697);
nand U1743 (N_1743,N_1665,N_1662);
xor U1744 (N_1744,N_1651,N_1671);
nand U1745 (N_1745,N_1665,N_1688);
nand U1746 (N_1746,N_1694,N_1660);
or U1747 (N_1747,N_1687,N_1673);
nor U1748 (N_1748,N_1664,N_1652);
or U1749 (N_1749,N_1673,N_1664);
and U1750 (N_1750,N_1729,N_1738);
and U1751 (N_1751,N_1706,N_1742);
and U1752 (N_1752,N_1704,N_1703);
or U1753 (N_1753,N_1721,N_1712);
and U1754 (N_1754,N_1701,N_1745);
and U1755 (N_1755,N_1710,N_1705);
or U1756 (N_1756,N_1727,N_1714);
or U1757 (N_1757,N_1717,N_1700);
and U1758 (N_1758,N_1725,N_1747);
and U1759 (N_1759,N_1722,N_1743);
nor U1760 (N_1760,N_1741,N_1728);
nor U1761 (N_1761,N_1736,N_1740);
nor U1762 (N_1762,N_1735,N_1730);
and U1763 (N_1763,N_1702,N_1719);
nor U1764 (N_1764,N_1724,N_1720);
nand U1765 (N_1765,N_1707,N_1746);
or U1766 (N_1766,N_1718,N_1708);
and U1767 (N_1767,N_1739,N_1744);
nor U1768 (N_1768,N_1716,N_1734);
nor U1769 (N_1769,N_1711,N_1726);
and U1770 (N_1770,N_1733,N_1748);
nand U1771 (N_1771,N_1749,N_1715);
nor U1772 (N_1772,N_1713,N_1737);
nand U1773 (N_1773,N_1731,N_1732);
or U1774 (N_1774,N_1709,N_1723);
nand U1775 (N_1775,N_1732,N_1742);
and U1776 (N_1776,N_1739,N_1745);
nand U1777 (N_1777,N_1746,N_1740);
nor U1778 (N_1778,N_1708,N_1734);
nor U1779 (N_1779,N_1735,N_1728);
nand U1780 (N_1780,N_1722,N_1734);
nand U1781 (N_1781,N_1730,N_1738);
or U1782 (N_1782,N_1743,N_1702);
nand U1783 (N_1783,N_1706,N_1702);
nand U1784 (N_1784,N_1706,N_1714);
nand U1785 (N_1785,N_1719,N_1714);
or U1786 (N_1786,N_1708,N_1725);
or U1787 (N_1787,N_1724,N_1721);
and U1788 (N_1788,N_1744,N_1730);
and U1789 (N_1789,N_1726,N_1713);
and U1790 (N_1790,N_1720,N_1747);
or U1791 (N_1791,N_1742,N_1737);
nor U1792 (N_1792,N_1704,N_1722);
or U1793 (N_1793,N_1719,N_1746);
or U1794 (N_1794,N_1729,N_1733);
or U1795 (N_1795,N_1716,N_1737);
nand U1796 (N_1796,N_1712,N_1746);
or U1797 (N_1797,N_1720,N_1738);
nand U1798 (N_1798,N_1706,N_1700);
and U1799 (N_1799,N_1736,N_1707);
or U1800 (N_1800,N_1778,N_1758);
nor U1801 (N_1801,N_1791,N_1750);
nand U1802 (N_1802,N_1799,N_1771);
and U1803 (N_1803,N_1786,N_1754);
or U1804 (N_1804,N_1780,N_1798);
or U1805 (N_1805,N_1766,N_1761);
nand U1806 (N_1806,N_1763,N_1769);
nor U1807 (N_1807,N_1775,N_1762);
and U1808 (N_1808,N_1782,N_1764);
and U1809 (N_1809,N_1792,N_1788);
nand U1810 (N_1810,N_1777,N_1774);
or U1811 (N_1811,N_1772,N_1783);
and U1812 (N_1812,N_1773,N_1755);
and U1813 (N_1813,N_1776,N_1759);
and U1814 (N_1814,N_1753,N_1794);
xnor U1815 (N_1815,N_1784,N_1787);
and U1816 (N_1816,N_1785,N_1795);
nand U1817 (N_1817,N_1767,N_1752);
xor U1818 (N_1818,N_1770,N_1760);
or U1819 (N_1819,N_1790,N_1779);
or U1820 (N_1820,N_1751,N_1789);
or U1821 (N_1821,N_1797,N_1756);
nand U1822 (N_1822,N_1765,N_1757);
and U1823 (N_1823,N_1768,N_1796);
nor U1824 (N_1824,N_1793,N_1781);
and U1825 (N_1825,N_1786,N_1797);
or U1826 (N_1826,N_1789,N_1783);
and U1827 (N_1827,N_1778,N_1788);
nand U1828 (N_1828,N_1772,N_1779);
nand U1829 (N_1829,N_1774,N_1795);
and U1830 (N_1830,N_1760,N_1762);
and U1831 (N_1831,N_1778,N_1759);
nor U1832 (N_1832,N_1776,N_1756);
nor U1833 (N_1833,N_1767,N_1777);
nor U1834 (N_1834,N_1786,N_1783);
and U1835 (N_1835,N_1753,N_1795);
nor U1836 (N_1836,N_1783,N_1787);
or U1837 (N_1837,N_1793,N_1765);
nor U1838 (N_1838,N_1762,N_1763);
nor U1839 (N_1839,N_1770,N_1780);
nor U1840 (N_1840,N_1791,N_1798);
and U1841 (N_1841,N_1790,N_1767);
nand U1842 (N_1842,N_1780,N_1762);
nand U1843 (N_1843,N_1788,N_1785);
nand U1844 (N_1844,N_1767,N_1796);
and U1845 (N_1845,N_1795,N_1767);
nand U1846 (N_1846,N_1799,N_1768);
or U1847 (N_1847,N_1793,N_1755);
or U1848 (N_1848,N_1798,N_1776);
and U1849 (N_1849,N_1777,N_1781);
xor U1850 (N_1850,N_1807,N_1816);
and U1851 (N_1851,N_1806,N_1828);
nand U1852 (N_1852,N_1824,N_1829);
or U1853 (N_1853,N_1804,N_1842);
and U1854 (N_1854,N_1810,N_1837);
or U1855 (N_1855,N_1835,N_1843);
or U1856 (N_1856,N_1848,N_1827);
nor U1857 (N_1857,N_1820,N_1805);
nor U1858 (N_1858,N_1847,N_1832);
and U1859 (N_1859,N_1808,N_1844);
and U1860 (N_1860,N_1826,N_1801);
or U1861 (N_1861,N_1817,N_1822);
and U1862 (N_1862,N_1830,N_1825);
nor U1863 (N_1863,N_1846,N_1812);
nor U1864 (N_1864,N_1819,N_1800);
and U1865 (N_1865,N_1809,N_1838);
nand U1866 (N_1866,N_1834,N_1823);
nand U1867 (N_1867,N_1803,N_1836);
and U1868 (N_1868,N_1814,N_1849);
nor U1869 (N_1869,N_1802,N_1845);
and U1870 (N_1870,N_1840,N_1811);
nor U1871 (N_1871,N_1839,N_1841);
and U1872 (N_1872,N_1831,N_1818);
and U1873 (N_1873,N_1815,N_1833);
nand U1874 (N_1874,N_1821,N_1813);
nor U1875 (N_1875,N_1818,N_1846);
xor U1876 (N_1876,N_1819,N_1820);
nor U1877 (N_1877,N_1842,N_1814);
or U1878 (N_1878,N_1824,N_1811);
xnor U1879 (N_1879,N_1824,N_1817);
nor U1880 (N_1880,N_1838,N_1805);
nand U1881 (N_1881,N_1834,N_1838);
and U1882 (N_1882,N_1825,N_1811);
or U1883 (N_1883,N_1802,N_1815);
xor U1884 (N_1884,N_1809,N_1800);
or U1885 (N_1885,N_1830,N_1829);
nand U1886 (N_1886,N_1828,N_1827);
xnor U1887 (N_1887,N_1812,N_1813);
and U1888 (N_1888,N_1813,N_1800);
nand U1889 (N_1889,N_1820,N_1833);
and U1890 (N_1890,N_1847,N_1804);
or U1891 (N_1891,N_1848,N_1812);
and U1892 (N_1892,N_1847,N_1833);
and U1893 (N_1893,N_1848,N_1810);
and U1894 (N_1894,N_1840,N_1819);
nand U1895 (N_1895,N_1813,N_1832);
and U1896 (N_1896,N_1810,N_1841);
nand U1897 (N_1897,N_1849,N_1811);
nand U1898 (N_1898,N_1844,N_1835);
or U1899 (N_1899,N_1846,N_1842);
nor U1900 (N_1900,N_1881,N_1850);
or U1901 (N_1901,N_1897,N_1861);
nor U1902 (N_1902,N_1896,N_1890);
nand U1903 (N_1903,N_1882,N_1854);
and U1904 (N_1904,N_1866,N_1886);
nand U1905 (N_1905,N_1871,N_1879);
and U1906 (N_1906,N_1892,N_1883);
or U1907 (N_1907,N_1863,N_1872);
and U1908 (N_1908,N_1891,N_1889);
nor U1909 (N_1909,N_1894,N_1877);
nor U1910 (N_1910,N_1874,N_1864);
and U1911 (N_1911,N_1899,N_1868);
nor U1912 (N_1912,N_1855,N_1862);
and U1913 (N_1913,N_1876,N_1870);
and U1914 (N_1914,N_1852,N_1853);
and U1915 (N_1915,N_1851,N_1893);
nand U1916 (N_1916,N_1859,N_1888);
or U1917 (N_1917,N_1878,N_1884);
nand U1918 (N_1918,N_1873,N_1856);
nand U1919 (N_1919,N_1865,N_1887);
or U1920 (N_1920,N_1869,N_1895);
nor U1921 (N_1921,N_1857,N_1875);
and U1922 (N_1922,N_1898,N_1867);
or U1923 (N_1923,N_1860,N_1858);
nand U1924 (N_1924,N_1880,N_1885);
xnor U1925 (N_1925,N_1880,N_1853);
nand U1926 (N_1926,N_1888,N_1877);
nor U1927 (N_1927,N_1895,N_1873);
nand U1928 (N_1928,N_1899,N_1878);
and U1929 (N_1929,N_1856,N_1893);
nand U1930 (N_1930,N_1876,N_1857);
nand U1931 (N_1931,N_1892,N_1868);
nor U1932 (N_1932,N_1874,N_1853);
and U1933 (N_1933,N_1899,N_1858);
nor U1934 (N_1934,N_1853,N_1865);
nor U1935 (N_1935,N_1896,N_1877);
or U1936 (N_1936,N_1899,N_1867);
and U1937 (N_1937,N_1863,N_1859);
nor U1938 (N_1938,N_1891,N_1893);
and U1939 (N_1939,N_1860,N_1895);
and U1940 (N_1940,N_1879,N_1882);
or U1941 (N_1941,N_1853,N_1871);
nor U1942 (N_1942,N_1857,N_1898);
nor U1943 (N_1943,N_1877,N_1858);
and U1944 (N_1944,N_1875,N_1891);
nand U1945 (N_1945,N_1855,N_1878);
or U1946 (N_1946,N_1897,N_1855);
and U1947 (N_1947,N_1882,N_1864);
or U1948 (N_1948,N_1883,N_1879);
nor U1949 (N_1949,N_1853,N_1877);
nor U1950 (N_1950,N_1939,N_1921);
nand U1951 (N_1951,N_1917,N_1919);
nor U1952 (N_1952,N_1915,N_1931);
or U1953 (N_1953,N_1918,N_1946);
or U1954 (N_1954,N_1900,N_1901);
and U1955 (N_1955,N_1932,N_1914);
nand U1956 (N_1956,N_1934,N_1911);
or U1957 (N_1957,N_1916,N_1936);
or U1958 (N_1958,N_1906,N_1920);
nand U1959 (N_1959,N_1940,N_1948);
and U1960 (N_1960,N_1908,N_1907);
or U1961 (N_1961,N_1937,N_1929);
xor U1962 (N_1962,N_1923,N_1903);
and U1963 (N_1963,N_1938,N_1928);
nor U1964 (N_1964,N_1930,N_1904);
or U1965 (N_1965,N_1924,N_1922);
or U1966 (N_1966,N_1945,N_1926);
or U1967 (N_1967,N_1947,N_1949);
or U1968 (N_1968,N_1910,N_1942);
nand U1969 (N_1969,N_1905,N_1944);
or U1970 (N_1970,N_1909,N_1943);
nand U1971 (N_1971,N_1912,N_1913);
or U1972 (N_1972,N_1902,N_1927);
or U1973 (N_1973,N_1935,N_1933);
nand U1974 (N_1974,N_1941,N_1925);
and U1975 (N_1975,N_1904,N_1929);
nand U1976 (N_1976,N_1914,N_1942);
nor U1977 (N_1977,N_1921,N_1920);
or U1978 (N_1978,N_1931,N_1912);
and U1979 (N_1979,N_1924,N_1927);
or U1980 (N_1980,N_1932,N_1903);
and U1981 (N_1981,N_1938,N_1946);
nor U1982 (N_1982,N_1912,N_1927);
nor U1983 (N_1983,N_1937,N_1939);
and U1984 (N_1984,N_1907,N_1923);
nand U1985 (N_1985,N_1940,N_1936);
and U1986 (N_1986,N_1939,N_1933);
or U1987 (N_1987,N_1937,N_1900);
and U1988 (N_1988,N_1931,N_1901);
or U1989 (N_1989,N_1941,N_1930);
nand U1990 (N_1990,N_1907,N_1904);
and U1991 (N_1991,N_1917,N_1924);
nand U1992 (N_1992,N_1939,N_1924);
nand U1993 (N_1993,N_1913,N_1911);
and U1994 (N_1994,N_1947,N_1938);
nand U1995 (N_1995,N_1918,N_1942);
nand U1996 (N_1996,N_1917,N_1926);
or U1997 (N_1997,N_1903,N_1907);
nor U1998 (N_1998,N_1943,N_1932);
and U1999 (N_1999,N_1932,N_1902);
nor U2000 (N_2000,N_1983,N_1957);
and U2001 (N_2001,N_1999,N_1955);
nor U2002 (N_2002,N_1994,N_1975);
or U2003 (N_2003,N_1973,N_1969);
nor U2004 (N_2004,N_1974,N_1967);
or U2005 (N_2005,N_1995,N_1986);
and U2006 (N_2006,N_1988,N_1978);
or U2007 (N_2007,N_1956,N_1993);
nand U2008 (N_2008,N_1959,N_1977);
xnor U2009 (N_2009,N_1952,N_1985);
nor U2010 (N_2010,N_1982,N_1968);
xor U2011 (N_2011,N_1960,N_1950);
nand U2012 (N_2012,N_1979,N_1984);
or U2013 (N_2013,N_1966,N_1963);
nor U2014 (N_2014,N_1965,N_1958);
nand U2015 (N_2015,N_1980,N_1953);
and U2016 (N_2016,N_1990,N_1998);
and U2017 (N_2017,N_1964,N_1976);
or U2018 (N_2018,N_1971,N_1997);
nand U2019 (N_2019,N_1970,N_1991);
and U2020 (N_2020,N_1989,N_1951);
and U2021 (N_2021,N_1961,N_1992);
nor U2022 (N_2022,N_1996,N_1954);
or U2023 (N_2023,N_1981,N_1972);
or U2024 (N_2024,N_1962,N_1987);
nor U2025 (N_2025,N_1978,N_1994);
and U2026 (N_2026,N_1968,N_1991);
nor U2027 (N_2027,N_1953,N_1970);
or U2028 (N_2028,N_1973,N_1957);
and U2029 (N_2029,N_1972,N_1984);
nor U2030 (N_2030,N_1996,N_1952);
nand U2031 (N_2031,N_1969,N_1994);
nor U2032 (N_2032,N_1972,N_1979);
nand U2033 (N_2033,N_1993,N_1992);
nand U2034 (N_2034,N_1961,N_1990);
and U2035 (N_2035,N_1969,N_1968);
nand U2036 (N_2036,N_1990,N_1955);
or U2037 (N_2037,N_1960,N_1986);
or U2038 (N_2038,N_1959,N_1978);
nor U2039 (N_2039,N_1970,N_1987);
and U2040 (N_2040,N_1968,N_1966);
or U2041 (N_2041,N_1953,N_1978);
nor U2042 (N_2042,N_1988,N_1951);
nor U2043 (N_2043,N_1999,N_1978);
xnor U2044 (N_2044,N_1991,N_1957);
nor U2045 (N_2045,N_1983,N_1987);
nand U2046 (N_2046,N_1961,N_1973);
xor U2047 (N_2047,N_1962,N_1973);
nand U2048 (N_2048,N_1970,N_1977);
or U2049 (N_2049,N_1981,N_1977);
nand U2050 (N_2050,N_2018,N_2005);
and U2051 (N_2051,N_2019,N_2045);
xor U2052 (N_2052,N_2002,N_2004);
and U2053 (N_2053,N_2016,N_2031);
or U2054 (N_2054,N_2020,N_2043);
nor U2055 (N_2055,N_2006,N_2032);
nor U2056 (N_2056,N_2044,N_2022);
and U2057 (N_2057,N_2026,N_2033);
nor U2058 (N_2058,N_2003,N_2012);
nand U2059 (N_2059,N_2046,N_2042);
nor U2060 (N_2060,N_2009,N_2040);
nand U2061 (N_2061,N_2011,N_2028);
nor U2062 (N_2062,N_2036,N_2048);
or U2063 (N_2063,N_2001,N_2030);
or U2064 (N_2064,N_2034,N_2023);
nand U2065 (N_2065,N_2047,N_2015);
nor U2066 (N_2066,N_2038,N_2029);
xor U2067 (N_2067,N_2000,N_2049);
and U2068 (N_2068,N_2010,N_2024);
and U2069 (N_2069,N_2021,N_2041);
nor U2070 (N_2070,N_2027,N_2008);
and U2071 (N_2071,N_2017,N_2014);
and U2072 (N_2072,N_2013,N_2039);
or U2073 (N_2073,N_2025,N_2007);
or U2074 (N_2074,N_2037,N_2035);
or U2075 (N_2075,N_2014,N_2010);
nand U2076 (N_2076,N_2035,N_2012);
nand U2077 (N_2077,N_2022,N_2003);
or U2078 (N_2078,N_2046,N_2017);
or U2079 (N_2079,N_2007,N_2026);
and U2080 (N_2080,N_2020,N_2028);
nor U2081 (N_2081,N_2027,N_2001);
nor U2082 (N_2082,N_2010,N_2021);
and U2083 (N_2083,N_2028,N_2004);
nor U2084 (N_2084,N_2011,N_2036);
nand U2085 (N_2085,N_2043,N_2040);
xnor U2086 (N_2086,N_2023,N_2045);
or U2087 (N_2087,N_2002,N_2015);
xor U2088 (N_2088,N_2010,N_2007);
xor U2089 (N_2089,N_2000,N_2040);
nor U2090 (N_2090,N_2049,N_2017);
nor U2091 (N_2091,N_2038,N_2019);
or U2092 (N_2092,N_2007,N_2039);
nor U2093 (N_2093,N_2005,N_2026);
nand U2094 (N_2094,N_2031,N_2018);
and U2095 (N_2095,N_2036,N_2013);
and U2096 (N_2096,N_2038,N_2017);
nand U2097 (N_2097,N_2043,N_2022);
nand U2098 (N_2098,N_2011,N_2027);
and U2099 (N_2099,N_2017,N_2009);
and U2100 (N_2100,N_2072,N_2062);
or U2101 (N_2101,N_2097,N_2091);
and U2102 (N_2102,N_2054,N_2078);
nor U2103 (N_2103,N_2094,N_2099);
and U2104 (N_2104,N_2098,N_2084);
nor U2105 (N_2105,N_2092,N_2066);
nand U2106 (N_2106,N_2064,N_2074);
or U2107 (N_2107,N_2093,N_2071);
nor U2108 (N_2108,N_2087,N_2075);
nor U2109 (N_2109,N_2083,N_2096);
or U2110 (N_2110,N_2090,N_2089);
nand U2111 (N_2111,N_2086,N_2058);
or U2112 (N_2112,N_2077,N_2067);
and U2113 (N_2113,N_2061,N_2080);
nor U2114 (N_2114,N_2057,N_2082);
and U2115 (N_2115,N_2050,N_2051);
nand U2116 (N_2116,N_2065,N_2079);
or U2117 (N_2117,N_2069,N_2055);
and U2118 (N_2118,N_2076,N_2095);
xnor U2119 (N_2119,N_2052,N_2088);
and U2120 (N_2120,N_2060,N_2073);
and U2121 (N_2121,N_2059,N_2070);
or U2122 (N_2122,N_2056,N_2085);
and U2123 (N_2123,N_2068,N_2063);
nand U2124 (N_2124,N_2081,N_2053);
and U2125 (N_2125,N_2079,N_2060);
nand U2126 (N_2126,N_2098,N_2066);
nor U2127 (N_2127,N_2054,N_2086);
nor U2128 (N_2128,N_2057,N_2079);
and U2129 (N_2129,N_2064,N_2088);
and U2130 (N_2130,N_2085,N_2074);
or U2131 (N_2131,N_2057,N_2052);
or U2132 (N_2132,N_2062,N_2096);
nand U2133 (N_2133,N_2099,N_2061);
nor U2134 (N_2134,N_2055,N_2063);
nand U2135 (N_2135,N_2068,N_2062);
or U2136 (N_2136,N_2063,N_2052);
or U2137 (N_2137,N_2084,N_2067);
and U2138 (N_2138,N_2091,N_2054);
nand U2139 (N_2139,N_2086,N_2074);
and U2140 (N_2140,N_2089,N_2074);
or U2141 (N_2141,N_2092,N_2078);
xor U2142 (N_2142,N_2050,N_2066);
or U2143 (N_2143,N_2070,N_2063);
nand U2144 (N_2144,N_2070,N_2055);
or U2145 (N_2145,N_2070,N_2050);
and U2146 (N_2146,N_2055,N_2072);
nand U2147 (N_2147,N_2051,N_2064);
nand U2148 (N_2148,N_2070,N_2071);
or U2149 (N_2149,N_2091,N_2082);
nor U2150 (N_2150,N_2122,N_2113);
or U2151 (N_2151,N_2117,N_2144);
and U2152 (N_2152,N_2101,N_2136);
or U2153 (N_2153,N_2125,N_2134);
and U2154 (N_2154,N_2133,N_2109);
nand U2155 (N_2155,N_2105,N_2141);
and U2156 (N_2156,N_2148,N_2126);
or U2157 (N_2157,N_2138,N_2146);
nor U2158 (N_2158,N_2102,N_2108);
or U2159 (N_2159,N_2110,N_2121);
or U2160 (N_2160,N_2135,N_2107);
nand U2161 (N_2161,N_2149,N_2119);
or U2162 (N_2162,N_2103,N_2123);
xor U2163 (N_2163,N_2128,N_2124);
xor U2164 (N_2164,N_2116,N_2137);
and U2165 (N_2165,N_2100,N_2120);
nand U2166 (N_2166,N_2132,N_2114);
or U2167 (N_2167,N_2118,N_2112);
xor U2168 (N_2168,N_2111,N_2142);
nand U2169 (N_2169,N_2145,N_2131);
nor U2170 (N_2170,N_2115,N_2130);
and U2171 (N_2171,N_2104,N_2147);
and U2172 (N_2172,N_2139,N_2127);
nand U2173 (N_2173,N_2129,N_2106);
and U2174 (N_2174,N_2143,N_2140);
and U2175 (N_2175,N_2139,N_2106);
nor U2176 (N_2176,N_2122,N_2104);
nand U2177 (N_2177,N_2111,N_2118);
xor U2178 (N_2178,N_2127,N_2105);
and U2179 (N_2179,N_2112,N_2123);
nand U2180 (N_2180,N_2143,N_2115);
nor U2181 (N_2181,N_2111,N_2144);
and U2182 (N_2182,N_2105,N_2121);
or U2183 (N_2183,N_2121,N_2141);
and U2184 (N_2184,N_2143,N_2114);
and U2185 (N_2185,N_2140,N_2109);
nand U2186 (N_2186,N_2109,N_2125);
or U2187 (N_2187,N_2147,N_2141);
nor U2188 (N_2188,N_2118,N_2133);
nor U2189 (N_2189,N_2144,N_2112);
nor U2190 (N_2190,N_2128,N_2118);
and U2191 (N_2191,N_2135,N_2139);
nand U2192 (N_2192,N_2142,N_2143);
xor U2193 (N_2193,N_2123,N_2102);
and U2194 (N_2194,N_2143,N_2124);
nor U2195 (N_2195,N_2110,N_2123);
nand U2196 (N_2196,N_2115,N_2107);
or U2197 (N_2197,N_2141,N_2113);
nor U2198 (N_2198,N_2113,N_2101);
nor U2199 (N_2199,N_2143,N_2130);
xnor U2200 (N_2200,N_2195,N_2174);
nand U2201 (N_2201,N_2154,N_2176);
and U2202 (N_2202,N_2162,N_2193);
nand U2203 (N_2203,N_2186,N_2169);
nor U2204 (N_2204,N_2151,N_2172);
or U2205 (N_2205,N_2170,N_2191);
and U2206 (N_2206,N_2177,N_2184);
and U2207 (N_2207,N_2171,N_2163);
or U2208 (N_2208,N_2152,N_2157);
and U2209 (N_2209,N_2190,N_2156);
nor U2210 (N_2210,N_2173,N_2165);
xor U2211 (N_2211,N_2189,N_2194);
nor U2212 (N_2212,N_2166,N_2196);
and U2213 (N_2213,N_2182,N_2187);
or U2214 (N_2214,N_2167,N_2159);
and U2215 (N_2215,N_2197,N_2181);
and U2216 (N_2216,N_2179,N_2150);
or U2217 (N_2217,N_2161,N_2199);
or U2218 (N_2218,N_2188,N_2192);
and U2219 (N_2219,N_2164,N_2155);
nand U2220 (N_2220,N_2198,N_2168);
and U2221 (N_2221,N_2185,N_2183);
nor U2222 (N_2222,N_2153,N_2178);
nand U2223 (N_2223,N_2175,N_2158);
or U2224 (N_2224,N_2180,N_2160);
and U2225 (N_2225,N_2154,N_2168);
nor U2226 (N_2226,N_2164,N_2162);
and U2227 (N_2227,N_2154,N_2159);
or U2228 (N_2228,N_2191,N_2183);
or U2229 (N_2229,N_2154,N_2180);
or U2230 (N_2230,N_2152,N_2163);
or U2231 (N_2231,N_2164,N_2177);
nand U2232 (N_2232,N_2196,N_2169);
and U2233 (N_2233,N_2197,N_2166);
and U2234 (N_2234,N_2151,N_2196);
and U2235 (N_2235,N_2173,N_2152);
nand U2236 (N_2236,N_2195,N_2171);
nand U2237 (N_2237,N_2161,N_2175);
or U2238 (N_2238,N_2194,N_2185);
or U2239 (N_2239,N_2175,N_2167);
or U2240 (N_2240,N_2174,N_2168);
and U2241 (N_2241,N_2179,N_2196);
nor U2242 (N_2242,N_2187,N_2194);
nand U2243 (N_2243,N_2163,N_2178);
nand U2244 (N_2244,N_2164,N_2194);
or U2245 (N_2245,N_2168,N_2191);
nand U2246 (N_2246,N_2179,N_2158);
nand U2247 (N_2247,N_2155,N_2183);
and U2248 (N_2248,N_2169,N_2198);
or U2249 (N_2249,N_2185,N_2191);
nand U2250 (N_2250,N_2223,N_2221);
nor U2251 (N_2251,N_2211,N_2219);
nand U2252 (N_2252,N_2209,N_2210);
or U2253 (N_2253,N_2202,N_2249);
xnor U2254 (N_2254,N_2200,N_2217);
or U2255 (N_2255,N_2233,N_2204);
nand U2256 (N_2256,N_2236,N_2234);
nand U2257 (N_2257,N_2215,N_2244);
or U2258 (N_2258,N_2240,N_2246);
or U2259 (N_2259,N_2226,N_2214);
or U2260 (N_2260,N_2206,N_2237);
nor U2261 (N_2261,N_2220,N_2227);
and U2262 (N_2262,N_2208,N_2212);
nand U2263 (N_2263,N_2207,N_2205);
nand U2264 (N_2264,N_2247,N_2229);
and U2265 (N_2265,N_2238,N_2235);
or U2266 (N_2266,N_2218,N_2230);
nor U2267 (N_2267,N_2241,N_2231);
and U2268 (N_2268,N_2232,N_2239);
nor U2269 (N_2269,N_2213,N_2248);
xor U2270 (N_2270,N_2224,N_2245);
nor U2271 (N_2271,N_2222,N_2228);
and U2272 (N_2272,N_2216,N_2201);
nand U2273 (N_2273,N_2243,N_2203);
nand U2274 (N_2274,N_2242,N_2225);
nand U2275 (N_2275,N_2217,N_2236);
and U2276 (N_2276,N_2208,N_2239);
nand U2277 (N_2277,N_2236,N_2230);
nand U2278 (N_2278,N_2206,N_2249);
and U2279 (N_2279,N_2207,N_2241);
or U2280 (N_2280,N_2216,N_2234);
or U2281 (N_2281,N_2242,N_2206);
or U2282 (N_2282,N_2232,N_2237);
nand U2283 (N_2283,N_2200,N_2226);
and U2284 (N_2284,N_2219,N_2228);
nand U2285 (N_2285,N_2241,N_2213);
and U2286 (N_2286,N_2245,N_2217);
and U2287 (N_2287,N_2221,N_2214);
nand U2288 (N_2288,N_2228,N_2238);
and U2289 (N_2289,N_2212,N_2200);
nand U2290 (N_2290,N_2219,N_2209);
xor U2291 (N_2291,N_2235,N_2237);
nor U2292 (N_2292,N_2233,N_2239);
nand U2293 (N_2293,N_2211,N_2212);
and U2294 (N_2294,N_2201,N_2241);
and U2295 (N_2295,N_2205,N_2208);
or U2296 (N_2296,N_2208,N_2202);
and U2297 (N_2297,N_2234,N_2219);
nand U2298 (N_2298,N_2240,N_2247);
or U2299 (N_2299,N_2228,N_2236);
nor U2300 (N_2300,N_2252,N_2254);
or U2301 (N_2301,N_2285,N_2286);
or U2302 (N_2302,N_2263,N_2272);
nor U2303 (N_2303,N_2294,N_2256);
or U2304 (N_2304,N_2280,N_2274);
and U2305 (N_2305,N_2267,N_2282);
and U2306 (N_2306,N_2262,N_2293);
xnor U2307 (N_2307,N_2296,N_2257);
or U2308 (N_2308,N_2265,N_2259);
nor U2309 (N_2309,N_2260,N_2291);
nand U2310 (N_2310,N_2289,N_2268);
and U2311 (N_2311,N_2251,N_2271);
nand U2312 (N_2312,N_2255,N_2287);
or U2313 (N_2313,N_2295,N_2269);
and U2314 (N_2314,N_2253,N_2284);
nand U2315 (N_2315,N_2275,N_2258);
nand U2316 (N_2316,N_2276,N_2281);
and U2317 (N_2317,N_2250,N_2283);
and U2318 (N_2318,N_2279,N_2264);
nor U2319 (N_2319,N_2278,N_2297);
nor U2320 (N_2320,N_2298,N_2292);
and U2321 (N_2321,N_2261,N_2299);
nor U2322 (N_2322,N_2273,N_2270);
nor U2323 (N_2323,N_2288,N_2266);
nand U2324 (N_2324,N_2290,N_2277);
or U2325 (N_2325,N_2296,N_2276);
nor U2326 (N_2326,N_2284,N_2252);
nor U2327 (N_2327,N_2296,N_2261);
nor U2328 (N_2328,N_2287,N_2266);
nor U2329 (N_2329,N_2269,N_2257);
nand U2330 (N_2330,N_2286,N_2271);
or U2331 (N_2331,N_2296,N_2286);
nor U2332 (N_2332,N_2276,N_2265);
xnor U2333 (N_2333,N_2289,N_2266);
or U2334 (N_2334,N_2274,N_2250);
nor U2335 (N_2335,N_2295,N_2293);
and U2336 (N_2336,N_2290,N_2267);
nor U2337 (N_2337,N_2264,N_2268);
or U2338 (N_2338,N_2288,N_2286);
and U2339 (N_2339,N_2291,N_2258);
or U2340 (N_2340,N_2286,N_2275);
nand U2341 (N_2341,N_2268,N_2294);
nand U2342 (N_2342,N_2287,N_2259);
and U2343 (N_2343,N_2277,N_2286);
and U2344 (N_2344,N_2275,N_2278);
nand U2345 (N_2345,N_2260,N_2252);
nand U2346 (N_2346,N_2271,N_2289);
nor U2347 (N_2347,N_2278,N_2258);
nand U2348 (N_2348,N_2280,N_2279);
xor U2349 (N_2349,N_2276,N_2268);
nor U2350 (N_2350,N_2307,N_2308);
nand U2351 (N_2351,N_2319,N_2311);
or U2352 (N_2352,N_2333,N_2325);
nor U2353 (N_2353,N_2344,N_2340);
nor U2354 (N_2354,N_2317,N_2330);
and U2355 (N_2355,N_2315,N_2303);
or U2356 (N_2356,N_2323,N_2334);
and U2357 (N_2357,N_2316,N_2312);
or U2358 (N_2358,N_2320,N_2347);
nor U2359 (N_2359,N_2343,N_2314);
nor U2360 (N_2360,N_2313,N_2305);
or U2361 (N_2361,N_2348,N_2306);
and U2362 (N_2362,N_2329,N_2338);
or U2363 (N_2363,N_2328,N_2349);
or U2364 (N_2364,N_2327,N_2302);
or U2365 (N_2365,N_2304,N_2301);
nor U2366 (N_2366,N_2322,N_2345);
and U2367 (N_2367,N_2335,N_2339);
and U2368 (N_2368,N_2341,N_2326);
and U2369 (N_2369,N_2300,N_2337);
nor U2370 (N_2370,N_2324,N_2331);
or U2371 (N_2371,N_2318,N_2310);
or U2372 (N_2372,N_2332,N_2346);
and U2373 (N_2373,N_2309,N_2336);
and U2374 (N_2374,N_2342,N_2321);
and U2375 (N_2375,N_2323,N_2322);
nor U2376 (N_2376,N_2311,N_2345);
nor U2377 (N_2377,N_2304,N_2335);
and U2378 (N_2378,N_2329,N_2324);
and U2379 (N_2379,N_2311,N_2316);
nor U2380 (N_2380,N_2311,N_2339);
nor U2381 (N_2381,N_2320,N_2318);
nand U2382 (N_2382,N_2332,N_2309);
nor U2383 (N_2383,N_2333,N_2336);
or U2384 (N_2384,N_2340,N_2312);
nor U2385 (N_2385,N_2311,N_2336);
nor U2386 (N_2386,N_2326,N_2307);
and U2387 (N_2387,N_2313,N_2344);
or U2388 (N_2388,N_2315,N_2347);
nand U2389 (N_2389,N_2301,N_2324);
nor U2390 (N_2390,N_2341,N_2343);
or U2391 (N_2391,N_2302,N_2313);
nand U2392 (N_2392,N_2326,N_2310);
nor U2393 (N_2393,N_2313,N_2338);
nand U2394 (N_2394,N_2308,N_2334);
and U2395 (N_2395,N_2339,N_2325);
or U2396 (N_2396,N_2333,N_2341);
xor U2397 (N_2397,N_2320,N_2312);
nor U2398 (N_2398,N_2348,N_2337);
and U2399 (N_2399,N_2340,N_2305);
or U2400 (N_2400,N_2383,N_2358);
and U2401 (N_2401,N_2390,N_2387);
and U2402 (N_2402,N_2397,N_2363);
or U2403 (N_2403,N_2380,N_2351);
or U2404 (N_2404,N_2381,N_2368);
or U2405 (N_2405,N_2364,N_2379);
nand U2406 (N_2406,N_2370,N_2361);
nand U2407 (N_2407,N_2374,N_2399);
or U2408 (N_2408,N_2388,N_2371);
nand U2409 (N_2409,N_2398,N_2373);
or U2410 (N_2410,N_2392,N_2359);
and U2411 (N_2411,N_2352,N_2378);
nand U2412 (N_2412,N_2360,N_2372);
and U2413 (N_2413,N_2353,N_2385);
or U2414 (N_2414,N_2394,N_2366);
or U2415 (N_2415,N_2354,N_2362);
nand U2416 (N_2416,N_2367,N_2395);
nor U2417 (N_2417,N_2382,N_2375);
nand U2418 (N_2418,N_2384,N_2377);
or U2419 (N_2419,N_2350,N_2391);
xnor U2420 (N_2420,N_2396,N_2389);
nor U2421 (N_2421,N_2365,N_2355);
and U2422 (N_2422,N_2393,N_2356);
or U2423 (N_2423,N_2357,N_2376);
nand U2424 (N_2424,N_2369,N_2386);
nand U2425 (N_2425,N_2387,N_2371);
nor U2426 (N_2426,N_2374,N_2381);
nand U2427 (N_2427,N_2395,N_2366);
xor U2428 (N_2428,N_2368,N_2358);
or U2429 (N_2429,N_2364,N_2395);
or U2430 (N_2430,N_2357,N_2395);
nand U2431 (N_2431,N_2361,N_2380);
nand U2432 (N_2432,N_2357,N_2390);
nor U2433 (N_2433,N_2353,N_2381);
and U2434 (N_2434,N_2378,N_2377);
and U2435 (N_2435,N_2367,N_2392);
or U2436 (N_2436,N_2382,N_2394);
nand U2437 (N_2437,N_2395,N_2380);
nor U2438 (N_2438,N_2398,N_2355);
nand U2439 (N_2439,N_2384,N_2359);
and U2440 (N_2440,N_2376,N_2381);
or U2441 (N_2441,N_2398,N_2392);
nor U2442 (N_2442,N_2386,N_2391);
nand U2443 (N_2443,N_2367,N_2373);
nand U2444 (N_2444,N_2398,N_2387);
nor U2445 (N_2445,N_2386,N_2368);
nand U2446 (N_2446,N_2353,N_2380);
and U2447 (N_2447,N_2381,N_2379);
or U2448 (N_2448,N_2384,N_2355);
and U2449 (N_2449,N_2367,N_2363);
or U2450 (N_2450,N_2427,N_2413);
or U2451 (N_2451,N_2411,N_2401);
nor U2452 (N_2452,N_2449,N_2443);
nor U2453 (N_2453,N_2424,N_2448);
nand U2454 (N_2454,N_2420,N_2439);
nand U2455 (N_2455,N_2408,N_2436);
and U2456 (N_2456,N_2426,N_2418);
nand U2457 (N_2457,N_2414,N_2441);
nand U2458 (N_2458,N_2438,N_2433);
xnor U2459 (N_2459,N_2404,N_2440);
and U2460 (N_2460,N_2429,N_2445);
nand U2461 (N_2461,N_2406,N_2415);
nand U2462 (N_2462,N_2446,N_2409);
nor U2463 (N_2463,N_2444,N_2403);
and U2464 (N_2464,N_2431,N_2419);
nand U2465 (N_2465,N_2407,N_2437);
or U2466 (N_2466,N_2435,N_2400);
nor U2467 (N_2467,N_2432,N_2417);
or U2468 (N_2468,N_2442,N_2422);
nor U2469 (N_2469,N_2428,N_2423);
or U2470 (N_2470,N_2447,N_2416);
nor U2471 (N_2471,N_2434,N_2430);
xnor U2472 (N_2472,N_2425,N_2412);
and U2473 (N_2473,N_2410,N_2421);
and U2474 (N_2474,N_2402,N_2405);
nand U2475 (N_2475,N_2423,N_2433);
nor U2476 (N_2476,N_2418,N_2443);
and U2477 (N_2477,N_2404,N_2424);
and U2478 (N_2478,N_2413,N_2423);
and U2479 (N_2479,N_2432,N_2412);
nor U2480 (N_2480,N_2414,N_2403);
nand U2481 (N_2481,N_2434,N_2417);
nor U2482 (N_2482,N_2423,N_2407);
or U2483 (N_2483,N_2417,N_2436);
or U2484 (N_2484,N_2410,N_2411);
nand U2485 (N_2485,N_2414,N_2409);
nor U2486 (N_2486,N_2432,N_2404);
nor U2487 (N_2487,N_2414,N_2400);
nor U2488 (N_2488,N_2402,N_2425);
or U2489 (N_2489,N_2434,N_2441);
nor U2490 (N_2490,N_2406,N_2423);
nor U2491 (N_2491,N_2416,N_2414);
and U2492 (N_2492,N_2439,N_2414);
nand U2493 (N_2493,N_2430,N_2405);
and U2494 (N_2494,N_2433,N_2416);
or U2495 (N_2495,N_2426,N_2434);
or U2496 (N_2496,N_2447,N_2439);
nand U2497 (N_2497,N_2423,N_2441);
nand U2498 (N_2498,N_2411,N_2408);
nand U2499 (N_2499,N_2402,N_2403);
or U2500 (N_2500,N_2498,N_2470);
or U2501 (N_2501,N_2469,N_2485);
and U2502 (N_2502,N_2473,N_2493);
or U2503 (N_2503,N_2487,N_2491);
and U2504 (N_2504,N_2472,N_2483);
or U2505 (N_2505,N_2495,N_2456);
and U2506 (N_2506,N_2496,N_2478);
and U2507 (N_2507,N_2474,N_2492);
and U2508 (N_2508,N_2460,N_2464);
nor U2509 (N_2509,N_2458,N_2457);
nor U2510 (N_2510,N_2462,N_2484);
nor U2511 (N_2511,N_2489,N_2486);
or U2512 (N_2512,N_2453,N_2479);
and U2513 (N_2513,N_2477,N_2463);
and U2514 (N_2514,N_2467,N_2471);
or U2515 (N_2515,N_2454,N_2466);
nand U2516 (N_2516,N_2450,N_2499);
nand U2517 (N_2517,N_2452,N_2475);
nor U2518 (N_2518,N_2482,N_2465);
or U2519 (N_2519,N_2476,N_2490);
and U2520 (N_2520,N_2480,N_2494);
nor U2521 (N_2521,N_2455,N_2459);
and U2522 (N_2522,N_2468,N_2497);
or U2523 (N_2523,N_2461,N_2488);
or U2524 (N_2524,N_2481,N_2451);
or U2525 (N_2525,N_2458,N_2474);
nand U2526 (N_2526,N_2482,N_2475);
nand U2527 (N_2527,N_2495,N_2453);
nand U2528 (N_2528,N_2497,N_2487);
or U2529 (N_2529,N_2490,N_2458);
or U2530 (N_2530,N_2451,N_2479);
or U2531 (N_2531,N_2484,N_2497);
or U2532 (N_2532,N_2485,N_2496);
nor U2533 (N_2533,N_2472,N_2497);
nand U2534 (N_2534,N_2451,N_2496);
or U2535 (N_2535,N_2473,N_2474);
or U2536 (N_2536,N_2481,N_2485);
or U2537 (N_2537,N_2451,N_2454);
or U2538 (N_2538,N_2480,N_2459);
nor U2539 (N_2539,N_2485,N_2498);
nor U2540 (N_2540,N_2480,N_2470);
or U2541 (N_2541,N_2474,N_2452);
nand U2542 (N_2542,N_2458,N_2492);
or U2543 (N_2543,N_2463,N_2481);
xnor U2544 (N_2544,N_2465,N_2479);
or U2545 (N_2545,N_2479,N_2498);
or U2546 (N_2546,N_2456,N_2467);
nor U2547 (N_2547,N_2474,N_2499);
or U2548 (N_2548,N_2457,N_2484);
and U2549 (N_2549,N_2496,N_2484);
nand U2550 (N_2550,N_2525,N_2524);
nor U2551 (N_2551,N_2533,N_2512);
or U2552 (N_2552,N_2538,N_2505);
nand U2553 (N_2553,N_2509,N_2542);
nand U2554 (N_2554,N_2511,N_2518);
nand U2555 (N_2555,N_2528,N_2548);
nand U2556 (N_2556,N_2536,N_2537);
nor U2557 (N_2557,N_2540,N_2510);
and U2558 (N_2558,N_2513,N_2543);
and U2559 (N_2559,N_2539,N_2502);
nand U2560 (N_2560,N_2503,N_2549);
nor U2561 (N_2561,N_2535,N_2547);
nor U2562 (N_2562,N_2519,N_2500);
nor U2563 (N_2563,N_2523,N_2521);
and U2564 (N_2564,N_2516,N_2506);
nor U2565 (N_2565,N_2531,N_2530);
or U2566 (N_2566,N_2541,N_2504);
nand U2567 (N_2567,N_2515,N_2514);
nor U2568 (N_2568,N_2527,N_2546);
and U2569 (N_2569,N_2520,N_2507);
nor U2570 (N_2570,N_2529,N_2544);
or U2571 (N_2571,N_2532,N_2534);
nor U2572 (N_2572,N_2526,N_2545);
nand U2573 (N_2573,N_2522,N_2517);
nand U2574 (N_2574,N_2501,N_2508);
and U2575 (N_2575,N_2512,N_2537);
and U2576 (N_2576,N_2502,N_2525);
nand U2577 (N_2577,N_2534,N_2519);
or U2578 (N_2578,N_2517,N_2508);
and U2579 (N_2579,N_2502,N_2531);
nand U2580 (N_2580,N_2518,N_2526);
or U2581 (N_2581,N_2506,N_2539);
or U2582 (N_2582,N_2512,N_2505);
and U2583 (N_2583,N_2536,N_2542);
or U2584 (N_2584,N_2544,N_2525);
nand U2585 (N_2585,N_2546,N_2504);
or U2586 (N_2586,N_2527,N_2502);
or U2587 (N_2587,N_2513,N_2541);
xor U2588 (N_2588,N_2536,N_2529);
and U2589 (N_2589,N_2502,N_2547);
or U2590 (N_2590,N_2513,N_2523);
nand U2591 (N_2591,N_2530,N_2541);
or U2592 (N_2592,N_2519,N_2528);
nor U2593 (N_2593,N_2501,N_2510);
nand U2594 (N_2594,N_2500,N_2547);
xor U2595 (N_2595,N_2532,N_2501);
nor U2596 (N_2596,N_2519,N_2525);
and U2597 (N_2597,N_2506,N_2528);
nor U2598 (N_2598,N_2511,N_2506);
nor U2599 (N_2599,N_2502,N_2509);
or U2600 (N_2600,N_2561,N_2574);
xnor U2601 (N_2601,N_2580,N_2579);
nand U2602 (N_2602,N_2592,N_2581);
nand U2603 (N_2603,N_2563,N_2567);
and U2604 (N_2604,N_2564,N_2572);
and U2605 (N_2605,N_2560,N_2593);
nand U2606 (N_2606,N_2556,N_2568);
and U2607 (N_2607,N_2566,N_2562);
nand U2608 (N_2608,N_2578,N_2598);
nor U2609 (N_2609,N_2554,N_2551);
and U2610 (N_2610,N_2590,N_2575);
nor U2611 (N_2611,N_2582,N_2586);
nor U2612 (N_2612,N_2550,N_2553);
nor U2613 (N_2613,N_2594,N_2597);
or U2614 (N_2614,N_2571,N_2570);
or U2615 (N_2615,N_2588,N_2555);
or U2616 (N_2616,N_2583,N_2565);
or U2617 (N_2617,N_2576,N_2599);
and U2618 (N_2618,N_2577,N_2557);
or U2619 (N_2619,N_2552,N_2585);
or U2620 (N_2620,N_2587,N_2595);
nor U2621 (N_2621,N_2558,N_2589);
nand U2622 (N_2622,N_2573,N_2596);
or U2623 (N_2623,N_2584,N_2559);
nand U2624 (N_2624,N_2569,N_2591);
nor U2625 (N_2625,N_2597,N_2584);
nand U2626 (N_2626,N_2589,N_2576);
and U2627 (N_2627,N_2561,N_2585);
nand U2628 (N_2628,N_2571,N_2559);
nand U2629 (N_2629,N_2599,N_2583);
and U2630 (N_2630,N_2561,N_2581);
and U2631 (N_2631,N_2561,N_2599);
or U2632 (N_2632,N_2560,N_2582);
and U2633 (N_2633,N_2553,N_2596);
or U2634 (N_2634,N_2566,N_2580);
nor U2635 (N_2635,N_2571,N_2582);
or U2636 (N_2636,N_2597,N_2578);
and U2637 (N_2637,N_2587,N_2598);
nand U2638 (N_2638,N_2557,N_2572);
or U2639 (N_2639,N_2580,N_2581);
nor U2640 (N_2640,N_2576,N_2583);
xor U2641 (N_2641,N_2589,N_2591);
and U2642 (N_2642,N_2559,N_2585);
nor U2643 (N_2643,N_2572,N_2592);
and U2644 (N_2644,N_2578,N_2582);
or U2645 (N_2645,N_2597,N_2563);
nand U2646 (N_2646,N_2556,N_2587);
nand U2647 (N_2647,N_2581,N_2587);
or U2648 (N_2648,N_2592,N_2577);
and U2649 (N_2649,N_2564,N_2556);
or U2650 (N_2650,N_2634,N_2620);
nor U2651 (N_2651,N_2643,N_2636);
nand U2652 (N_2652,N_2633,N_2602);
and U2653 (N_2653,N_2600,N_2612);
nand U2654 (N_2654,N_2623,N_2647);
nand U2655 (N_2655,N_2625,N_2622);
or U2656 (N_2656,N_2648,N_2615);
nor U2657 (N_2657,N_2619,N_2641);
and U2658 (N_2658,N_2624,N_2630);
and U2659 (N_2659,N_2611,N_2635);
and U2660 (N_2660,N_2629,N_2610);
nand U2661 (N_2661,N_2632,N_2603);
nor U2662 (N_2662,N_2621,N_2640);
nor U2663 (N_2663,N_2608,N_2642);
or U2664 (N_2664,N_2637,N_2639);
or U2665 (N_2665,N_2617,N_2606);
nand U2666 (N_2666,N_2631,N_2638);
and U2667 (N_2667,N_2616,N_2649);
or U2668 (N_2668,N_2618,N_2605);
xnor U2669 (N_2669,N_2609,N_2604);
nor U2670 (N_2670,N_2644,N_2613);
and U2671 (N_2671,N_2601,N_2626);
nor U2672 (N_2672,N_2645,N_2607);
and U2673 (N_2673,N_2614,N_2627);
nor U2674 (N_2674,N_2628,N_2646);
nor U2675 (N_2675,N_2608,N_2643);
nand U2676 (N_2676,N_2611,N_2629);
nand U2677 (N_2677,N_2602,N_2644);
nand U2678 (N_2678,N_2605,N_2609);
nor U2679 (N_2679,N_2627,N_2626);
nand U2680 (N_2680,N_2602,N_2641);
or U2681 (N_2681,N_2618,N_2607);
nand U2682 (N_2682,N_2605,N_2617);
nand U2683 (N_2683,N_2632,N_2608);
nor U2684 (N_2684,N_2625,N_2619);
and U2685 (N_2685,N_2629,N_2601);
nor U2686 (N_2686,N_2631,N_2633);
nand U2687 (N_2687,N_2616,N_2627);
and U2688 (N_2688,N_2625,N_2629);
or U2689 (N_2689,N_2622,N_2623);
nand U2690 (N_2690,N_2625,N_2607);
or U2691 (N_2691,N_2649,N_2639);
and U2692 (N_2692,N_2626,N_2621);
nor U2693 (N_2693,N_2617,N_2601);
and U2694 (N_2694,N_2619,N_2637);
nand U2695 (N_2695,N_2633,N_2645);
and U2696 (N_2696,N_2646,N_2620);
nand U2697 (N_2697,N_2622,N_2621);
or U2698 (N_2698,N_2648,N_2620);
nor U2699 (N_2699,N_2613,N_2627);
or U2700 (N_2700,N_2687,N_2699);
xor U2701 (N_2701,N_2698,N_2681);
and U2702 (N_2702,N_2668,N_2659);
nand U2703 (N_2703,N_2665,N_2666);
or U2704 (N_2704,N_2661,N_2679);
and U2705 (N_2705,N_2684,N_2695);
nor U2706 (N_2706,N_2653,N_2656);
or U2707 (N_2707,N_2658,N_2669);
nand U2708 (N_2708,N_2670,N_2693);
and U2709 (N_2709,N_2674,N_2676);
and U2710 (N_2710,N_2650,N_2697);
or U2711 (N_2711,N_2677,N_2694);
or U2712 (N_2712,N_2682,N_2696);
or U2713 (N_2713,N_2673,N_2692);
nor U2714 (N_2714,N_2683,N_2685);
or U2715 (N_2715,N_2675,N_2662);
nor U2716 (N_2716,N_2686,N_2678);
nand U2717 (N_2717,N_2672,N_2651);
or U2718 (N_2718,N_2671,N_2690);
nand U2719 (N_2719,N_2691,N_2660);
nor U2720 (N_2720,N_2652,N_2664);
nor U2721 (N_2721,N_2657,N_2688);
nor U2722 (N_2722,N_2654,N_2689);
nor U2723 (N_2723,N_2663,N_2680);
nand U2724 (N_2724,N_2667,N_2655);
or U2725 (N_2725,N_2690,N_2650);
or U2726 (N_2726,N_2691,N_2651);
and U2727 (N_2727,N_2656,N_2695);
nand U2728 (N_2728,N_2651,N_2668);
or U2729 (N_2729,N_2685,N_2650);
nand U2730 (N_2730,N_2680,N_2677);
nor U2731 (N_2731,N_2652,N_2687);
and U2732 (N_2732,N_2692,N_2699);
nand U2733 (N_2733,N_2673,N_2682);
or U2734 (N_2734,N_2659,N_2660);
nand U2735 (N_2735,N_2654,N_2671);
nand U2736 (N_2736,N_2694,N_2675);
nor U2737 (N_2737,N_2660,N_2674);
or U2738 (N_2738,N_2669,N_2676);
nor U2739 (N_2739,N_2691,N_2659);
nor U2740 (N_2740,N_2676,N_2681);
or U2741 (N_2741,N_2674,N_2657);
or U2742 (N_2742,N_2683,N_2671);
nor U2743 (N_2743,N_2676,N_2687);
or U2744 (N_2744,N_2657,N_2656);
and U2745 (N_2745,N_2670,N_2672);
xor U2746 (N_2746,N_2654,N_2656);
nor U2747 (N_2747,N_2689,N_2661);
and U2748 (N_2748,N_2679,N_2699);
and U2749 (N_2749,N_2691,N_2679);
nand U2750 (N_2750,N_2710,N_2738);
and U2751 (N_2751,N_2718,N_2725);
nand U2752 (N_2752,N_2715,N_2717);
or U2753 (N_2753,N_2722,N_2709);
or U2754 (N_2754,N_2740,N_2716);
or U2755 (N_2755,N_2735,N_2745);
or U2756 (N_2756,N_2731,N_2742);
nand U2757 (N_2757,N_2700,N_2706);
nand U2758 (N_2758,N_2732,N_2712);
nor U2759 (N_2759,N_2734,N_2723);
or U2760 (N_2760,N_2728,N_2721);
or U2761 (N_2761,N_2747,N_2737);
or U2762 (N_2762,N_2705,N_2730);
xor U2763 (N_2763,N_2741,N_2749);
or U2764 (N_2764,N_2746,N_2720);
and U2765 (N_2765,N_2701,N_2704);
and U2766 (N_2766,N_2729,N_2733);
and U2767 (N_2767,N_2714,N_2703);
nand U2768 (N_2768,N_2719,N_2707);
nand U2769 (N_2769,N_2739,N_2736);
or U2770 (N_2770,N_2726,N_2708);
and U2771 (N_2771,N_2724,N_2727);
nor U2772 (N_2772,N_2711,N_2713);
or U2773 (N_2773,N_2744,N_2743);
nor U2774 (N_2774,N_2702,N_2748);
xnor U2775 (N_2775,N_2714,N_2739);
and U2776 (N_2776,N_2732,N_2739);
nor U2777 (N_2777,N_2741,N_2705);
or U2778 (N_2778,N_2734,N_2741);
and U2779 (N_2779,N_2735,N_2714);
nor U2780 (N_2780,N_2729,N_2705);
or U2781 (N_2781,N_2708,N_2714);
or U2782 (N_2782,N_2700,N_2740);
or U2783 (N_2783,N_2743,N_2701);
nor U2784 (N_2784,N_2734,N_2731);
nand U2785 (N_2785,N_2737,N_2728);
nor U2786 (N_2786,N_2732,N_2734);
and U2787 (N_2787,N_2730,N_2737);
nand U2788 (N_2788,N_2742,N_2747);
nand U2789 (N_2789,N_2735,N_2701);
or U2790 (N_2790,N_2700,N_2732);
or U2791 (N_2791,N_2741,N_2738);
nand U2792 (N_2792,N_2734,N_2701);
and U2793 (N_2793,N_2704,N_2702);
or U2794 (N_2794,N_2707,N_2734);
nor U2795 (N_2795,N_2722,N_2717);
nand U2796 (N_2796,N_2744,N_2706);
or U2797 (N_2797,N_2725,N_2744);
nand U2798 (N_2798,N_2720,N_2741);
nand U2799 (N_2799,N_2725,N_2741);
nor U2800 (N_2800,N_2793,N_2751);
or U2801 (N_2801,N_2755,N_2765);
or U2802 (N_2802,N_2778,N_2776);
nor U2803 (N_2803,N_2753,N_2762);
and U2804 (N_2804,N_2750,N_2754);
nor U2805 (N_2805,N_2756,N_2795);
or U2806 (N_2806,N_2771,N_2773);
nor U2807 (N_2807,N_2763,N_2781);
and U2808 (N_2808,N_2766,N_2777);
nor U2809 (N_2809,N_2758,N_2790);
nand U2810 (N_2810,N_2775,N_2782);
and U2811 (N_2811,N_2799,N_2768);
and U2812 (N_2812,N_2764,N_2787);
or U2813 (N_2813,N_2784,N_2767);
or U2814 (N_2814,N_2779,N_2770);
nand U2815 (N_2815,N_2794,N_2797);
nand U2816 (N_2816,N_2774,N_2798);
nand U2817 (N_2817,N_2761,N_2791);
and U2818 (N_2818,N_2785,N_2789);
and U2819 (N_2819,N_2769,N_2783);
and U2820 (N_2820,N_2772,N_2788);
nand U2821 (N_2821,N_2786,N_2757);
nand U2822 (N_2822,N_2760,N_2752);
and U2823 (N_2823,N_2792,N_2780);
or U2824 (N_2824,N_2796,N_2759);
nand U2825 (N_2825,N_2772,N_2790);
or U2826 (N_2826,N_2764,N_2783);
nor U2827 (N_2827,N_2792,N_2794);
or U2828 (N_2828,N_2791,N_2790);
and U2829 (N_2829,N_2779,N_2769);
nor U2830 (N_2830,N_2779,N_2773);
and U2831 (N_2831,N_2777,N_2797);
or U2832 (N_2832,N_2776,N_2755);
nand U2833 (N_2833,N_2773,N_2788);
nor U2834 (N_2834,N_2779,N_2767);
and U2835 (N_2835,N_2751,N_2753);
and U2836 (N_2836,N_2758,N_2769);
or U2837 (N_2837,N_2771,N_2761);
or U2838 (N_2838,N_2792,N_2793);
or U2839 (N_2839,N_2761,N_2768);
or U2840 (N_2840,N_2777,N_2782);
and U2841 (N_2841,N_2761,N_2794);
nor U2842 (N_2842,N_2778,N_2759);
and U2843 (N_2843,N_2778,N_2762);
nor U2844 (N_2844,N_2753,N_2787);
nand U2845 (N_2845,N_2795,N_2781);
or U2846 (N_2846,N_2781,N_2771);
nand U2847 (N_2847,N_2760,N_2775);
nand U2848 (N_2848,N_2776,N_2797);
or U2849 (N_2849,N_2782,N_2761);
nand U2850 (N_2850,N_2833,N_2846);
xnor U2851 (N_2851,N_2807,N_2818);
nor U2852 (N_2852,N_2813,N_2805);
or U2853 (N_2853,N_2838,N_2801);
nand U2854 (N_2854,N_2803,N_2848);
nand U2855 (N_2855,N_2817,N_2820);
nor U2856 (N_2856,N_2829,N_2847);
nor U2857 (N_2857,N_2842,N_2836);
nor U2858 (N_2858,N_2808,N_2823);
or U2859 (N_2859,N_2824,N_2834);
nor U2860 (N_2860,N_2821,N_2816);
or U2861 (N_2861,N_2840,N_2845);
nand U2862 (N_2862,N_2809,N_2812);
nand U2863 (N_2863,N_2828,N_2826);
and U2864 (N_2864,N_2819,N_2802);
nand U2865 (N_2865,N_2839,N_2825);
or U2866 (N_2866,N_2811,N_2810);
and U2867 (N_2867,N_2822,N_2806);
and U2868 (N_2868,N_2837,N_2814);
nand U2869 (N_2869,N_2832,N_2835);
and U2870 (N_2870,N_2800,N_2830);
nor U2871 (N_2871,N_2844,N_2849);
nand U2872 (N_2872,N_2815,N_2841);
nor U2873 (N_2873,N_2827,N_2831);
nor U2874 (N_2874,N_2804,N_2843);
nor U2875 (N_2875,N_2811,N_2828);
nor U2876 (N_2876,N_2806,N_2825);
or U2877 (N_2877,N_2811,N_2838);
nand U2878 (N_2878,N_2815,N_2820);
nor U2879 (N_2879,N_2841,N_2809);
or U2880 (N_2880,N_2818,N_2814);
nor U2881 (N_2881,N_2837,N_2809);
or U2882 (N_2882,N_2804,N_2834);
xnor U2883 (N_2883,N_2805,N_2834);
or U2884 (N_2884,N_2820,N_2833);
and U2885 (N_2885,N_2839,N_2803);
nand U2886 (N_2886,N_2844,N_2840);
and U2887 (N_2887,N_2820,N_2843);
and U2888 (N_2888,N_2834,N_2825);
nand U2889 (N_2889,N_2837,N_2822);
nor U2890 (N_2890,N_2827,N_2816);
nor U2891 (N_2891,N_2815,N_2835);
or U2892 (N_2892,N_2808,N_2803);
or U2893 (N_2893,N_2819,N_2838);
nor U2894 (N_2894,N_2801,N_2810);
nor U2895 (N_2895,N_2824,N_2846);
nor U2896 (N_2896,N_2847,N_2806);
or U2897 (N_2897,N_2822,N_2803);
xnor U2898 (N_2898,N_2802,N_2817);
nor U2899 (N_2899,N_2805,N_2803);
nand U2900 (N_2900,N_2869,N_2855);
nand U2901 (N_2901,N_2888,N_2876);
or U2902 (N_2902,N_2875,N_2885);
xor U2903 (N_2903,N_2854,N_2853);
or U2904 (N_2904,N_2879,N_2893);
xor U2905 (N_2905,N_2873,N_2858);
or U2906 (N_2906,N_2857,N_2897);
and U2907 (N_2907,N_2881,N_2871);
or U2908 (N_2908,N_2895,N_2878);
and U2909 (N_2909,N_2863,N_2862);
nand U2910 (N_2910,N_2896,N_2872);
nor U2911 (N_2911,N_2887,N_2864);
and U2912 (N_2912,N_2892,N_2851);
nand U2913 (N_2913,N_2856,N_2891);
or U2914 (N_2914,N_2890,N_2883);
nand U2915 (N_2915,N_2850,N_2889);
xor U2916 (N_2916,N_2861,N_2859);
or U2917 (N_2917,N_2898,N_2882);
nand U2918 (N_2918,N_2860,N_2880);
or U2919 (N_2919,N_2894,N_2867);
and U2920 (N_2920,N_2877,N_2868);
and U2921 (N_2921,N_2866,N_2886);
xor U2922 (N_2922,N_2870,N_2865);
or U2923 (N_2923,N_2852,N_2874);
or U2924 (N_2924,N_2899,N_2884);
or U2925 (N_2925,N_2871,N_2891);
nor U2926 (N_2926,N_2863,N_2867);
nand U2927 (N_2927,N_2865,N_2881);
nor U2928 (N_2928,N_2879,N_2880);
and U2929 (N_2929,N_2855,N_2889);
and U2930 (N_2930,N_2858,N_2872);
and U2931 (N_2931,N_2852,N_2864);
nor U2932 (N_2932,N_2858,N_2864);
or U2933 (N_2933,N_2865,N_2895);
or U2934 (N_2934,N_2891,N_2879);
nand U2935 (N_2935,N_2860,N_2857);
nor U2936 (N_2936,N_2867,N_2862);
and U2937 (N_2937,N_2875,N_2878);
and U2938 (N_2938,N_2871,N_2853);
nand U2939 (N_2939,N_2896,N_2867);
nor U2940 (N_2940,N_2889,N_2877);
nand U2941 (N_2941,N_2850,N_2859);
or U2942 (N_2942,N_2880,N_2876);
nor U2943 (N_2943,N_2860,N_2889);
nor U2944 (N_2944,N_2860,N_2874);
or U2945 (N_2945,N_2878,N_2877);
or U2946 (N_2946,N_2896,N_2861);
and U2947 (N_2947,N_2853,N_2898);
nor U2948 (N_2948,N_2865,N_2886);
nand U2949 (N_2949,N_2886,N_2898);
nor U2950 (N_2950,N_2902,N_2914);
nand U2951 (N_2951,N_2918,N_2915);
and U2952 (N_2952,N_2909,N_2939);
nand U2953 (N_2953,N_2947,N_2924);
nor U2954 (N_2954,N_2936,N_2912);
nor U2955 (N_2955,N_2943,N_2913);
nor U2956 (N_2956,N_2934,N_2908);
nor U2957 (N_2957,N_2921,N_2919);
nand U2958 (N_2958,N_2927,N_2905);
nand U2959 (N_2959,N_2904,N_2933);
nand U2960 (N_2960,N_2911,N_2942);
nor U2961 (N_2961,N_2935,N_2945);
and U2962 (N_2962,N_2946,N_2925);
nand U2963 (N_2963,N_2920,N_2926);
or U2964 (N_2964,N_2929,N_2930);
and U2965 (N_2965,N_2903,N_2900);
nor U2966 (N_2966,N_2907,N_2931);
and U2967 (N_2967,N_2901,N_2938);
nand U2968 (N_2968,N_2928,N_2949);
and U2969 (N_2969,N_2916,N_2948);
and U2970 (N_2970,N_2923,N_2932);
and U2971 (N_2971,N_2906,N_2944);
or U2972 (N_2972,N_2940,N_2941);
nand U2973 (N_2973,N_2937,N_2917);
nor U2974 (N_2974,N_2910,N_2922);
and U2975 (N_2975,N_2928,N_2906);
nor U2976 (N_2976,N_2928,N_2902);
and U2977 (N_2977,N_2940,N_2919);
or U2978 (N_2978,N_2934,N_2917);
or U2979 (N_2979,N_2901,N_2928);
nor U2980 (N_2980,N_2946,N_2941);
nor U2981 (N_2981,N_2929,N_2912);
nor U2982 (N_2982,N_2947,N_2945);
or U2983 (N_2983,N_2940,N_2937);
and U2984 (N_2984,N_2903,N_2927);
nand U2985 (N_2985,N_2940,N_2948);
nor U2986 (N_2986,N_2933,N_2915);
and U2987 (N_2987,N_2902,N_2934);
nand U2988 (N_2988,N_2942,N_2923);
and U2989 (N_2989,N_2918,N_2946);
nor U2990 (N_2990,N_2917,N_2949);
nor U2991 (N_2991,N_2909,N_2940);
and U2992 (N_2992,N_2940,N_2928);
nor U2993 (N_2993,N_2945,N_2922);
or U2994 (N_2994,N_2920,N_2909);
nor U2995 (N_2995,N_2938,N_2900);
nor U2996 (N_2996,N_2925,N_2941);
and U2997 (N_2997,N_2903,N_2924);
nor U2998 (N_2998,N_2938,N_2936);
and U2999 (N_2999,N_2915,N_2941);
or UO_0 (O_0,N_2970,N_2966);
nor UO_1 (O_1,N_2998,N_2991);
or UO_2 (O_2,N_2973,N_2994);
nand UO_3 (O_3,N_2963,N_2996);
nor UO_4 (O_4,N_2968,N_2989);
or UO_5 (O_5,N_2964,N_2974);
or UO_6 (O_6,N_2981,N_2987);
nand UO_7 (O_7,N_2960,N_2986);
or UO_8 (O_8,N_2953,N_2961);
nand UO_9 (O_9,N_2959,N_2979);
or UO_10 (O_10,N_2997,N_2983);
or UO_11 (O_11,N_2969,N_2993);
nor UO_12 (O_12,N_2956,N_2952);
nor UO_13 (O_13,N_2980,N_2978);
nand UO_14 (O_14,N_2984,N_2972);
nor UO_15 (O_15,N_2950,N_2975);
or UO_16 (O_16,N_2992,N_2965);
or UO_17 (O_17,N_2976,N_2988);
or UO_18 (O_18,N_2962,N_2990);
and UO_19 (O_19,N_2954,N_2995);
nand UO_20 (O_20,N_2999,N_2957);
nand UO_21 (O_21,N_2977,N_2967);
or UO_22 (O_22,N_2985,N_2958);
nor UO_23 (O_23,N_2951,N_2955);
nor UO_24 (O_24,N_2971,N_2982);
and UO_25 (O_25,N_2967,N_2987);
xor UO_26 (O_26,N_2973,N_2955);
or UO_27 (O_27,N_2982,N_2996);
or UO_28 (O_28,N_2970,N_2963);
nor UO_29 (O_29,N_2987,N_2955);
and UO_30 (O_30,N_2989,N_2994);
and UO_31 (O_31,N_2961,N_2962);
nand UO_32 (O_32,N_2979,N_2974);
nor UO_33 (O_33,N_2999,N_2953);
nor UO_34 (O_34,N_2985,N_2956);
nand UO_35 (O_35,N_2988,N_2987);
nand UO_36 (O_36,N_2967,N_2999);
nor UO_37 (O_37,N_2960,N_2965);
nor UO_38 (O_38,N_2951,N_2974);
xnor UO_39 (O_39,N_2968,N_2964);
nand UO_40 (O_40,N_2971,N_2983);
or UO_41 (O_41,N_2995,N_2972);
nand UO_42 (O_42,N_2994,N_2979);
or UO_43 (O_43,N_2972,N_2964);
and UO_44 (O_44,N_2952,N_2997);
and UO_45 (O_45,N_2979,N_2952);
and UO_46 (O_46,N_2993,N_2971);
nor UO_47 (O_47,N_2989,N_2996);
or UO_48 (O_48,N_2970,N_2995);
and UO_49 (O_49,N_2988,N_2980);
nor UO_50 (O_50,N_2989,N_2956);
nor UO_51 (O_51,N_2967,N_2953);
and UO_52 (O_52,N_2970,N_2958);
and UO_53 (O_53,N_2954,N_2956);
nor UO_54 (O_54,N_2951,N_2959);
nand UO_55 (O_55,N_2964,N_2954);
or UO_56 (O_56,N_2995,N_2973);
or UO_57 (O_57,N_2957,N_2968);
or UO_58 (O_58,N_2991,N_2959);
and UO_59 (O_59,N_2978,N_2986);
nor UO_60 (O_60,N_2959,N_2997);
nor UO_61 (O_61,N_2968,N_2986);
nor UO_62 (O_62,N_2997,N_2998);
or UO_63 (O_63,N_2961,N_2973);
nand UO_64 (O_64,N_2950,N_2984);
or UO_65 (O_65,N_2988,N_2971);
nand UO_66 (O_66,N_2991,N_2967);
or UO_67 (O_67,N_2960,N_2988);
nor UO_68 (O_68,N_2962,N_2986);
nand UO_69 (O_69,N_2981,N_2959);
nand UO_70 (O_70,N_2977,N_2964);
or UO_71 (O_71,N_2952,N_2991);
nand UO_72 (O_72,N_2950,N_2964);
nor UO_73 (O_73,N_2987,N_2985);
or UO_74 (O_74,N_2958,N_2995);
or UO_75 (O_75,N_2985,N_2976);
or UO_76 (O_76,N_2979,N_2961);
or UO_77 (O_77,N_2964,N_2987);
xor UO_78 (O_78,N_2995,N_2951);
or UO_79 (O_79,N_2981,N_2961);
or UO_80 (O_80,N_2999,N_2965);
or UO_81 (O_81,N_2972,N_2985);
nand UO_82 (O_82,N_2958,N_2978);
and UO_83 (O_83,N_2980,N_2983);
nand UO_84 (O_84,N_2998,N_2958);
nand UO_85 (O_85,N_2991,N_2989);
or UO_86 (O_86,N_2990,N_2967);
or UO_87 (O_87,N_2977,N_2963);
nand UO_88 (O_88,N_2975,N_2978);
nand UO_89 (O_89,N_2977,N_2992);
and UO_90 (O_90,N_2968,N_2999);
and UO_91 (O_91,N_2967,N_2969);
nand UO_92 (O_92,N_2967,N_2984);
and UO_93 (O_93,N_2959,N_2965);
nand UO_94 (O_94,N_2982,N_2992);
and UO_95 (O_95,N_2966,N_2977);
nand UO_96 (O_96,N_2998,N_2995);
or UO_97 (O_97,N_2978,N_2962);
or UO_98 (O_98,N_2963,N_2967);
nand UO_99 (O_99,N_2981,N_2988);
nand UO_100 (O_100,N_2987,N_2997);
and UO_101 (O_101,N_2996,N_2991);
nand UO_102 (O_102,N_2986,N_2995);
xor UO_103 (O_103,N_2957,N_2996);
nand UO_104 (O_104,N_2969,N_2954);
and UO_105 (O_105,N_2982,N_2997);
nand UO_106 (O_106,N_2973,N_2977);
or UO_107 (O_107,N_2950,N_2992);
and UO_108 (O_108,N_2963,N_2954);
nand UO_109 (O_109,N_2961,N_2959);
nor UO_110 (O_110,N_2993,N_2970);
nor UO_111 (O_111,N_2980,N_2961);
and UO_112 (O_112,N_2969,N_2960);
nand UO_113 (O_113,N_2979,N_2989);
nand UO_114 (O_114,N_2982,N_2990);
or UO_115 (O_115,N_2975,N_2963);
and UO_116 (O_116,N_2955,N_2970);
nor UO_117 (O_117,N_2968,N_2977);
nor UO_118 (O_118,N_2983,N_2987);
and UO_119 (O_119,N_2969,N_2972);
or UO_120 (O_120,N_2971,N_2998);
nor UO_121 (O_121,N_2955,N_2974);
or UO_122 (O_122,N_2983,N_2990);
nor UO_123 (O_123,N_2982,N_2999);
nor UO_124 (O_124,N_2996,N_2998);
or UO_125 (O_125,N_2960,N_2964);
or UO_126 (O_126,N_2962,N_2968);
nor UO_127 (O_127,N_2959,N_2964);
nand UO_128 (O_128,N_2995,N_2980);
nand UO_129 (O_129,N_2985,N_2982);
or UO_130 (O_130,N_2966,N_2984);
and UO_131 (O_131,N_2960,N_2962);
and UO_132 (O_132,N_2980,N_2987);
nand UO_133 (O_133,N_2999,N_2990);
nor UO_134 (O_134,N_2956,N_2990);
or UO_135 (O_135,N_2982,N_2978);
nor UO_136 (O_136,N_2996,N_2992);
nor UO_137 (O_137,N_2996,N_2999);
nand UO_138 (O_138,N_2995,N_2965);
and UO_139 (O_139,N_2984,N_2991);
and UO_140 (O_140,N_2969,N_2997);
nand UO_141 (O_141,N_2973,N_2965);
and UO_142 (O_142,N_2971,N_2985);
nand UO_143 (O_143,N_2952,N_2981);
nor UO_144 (O_144,N_2961,N_2970);
and UO_145 (O_145,N_2977,N_2959);
nor UO_146 (O_146,N_2990,N_2970);
nand UO_147 (O_147,N_2959,N_2952);
or UO_148 (O_148,N_2978,N_2996);
nand UO_149 (O_149,N_2986,N_2961);
or UO_150 (O_150,N_2968,N_2958);
or UO_151 (O_151,N_2980,N_2989);
or UO_152 (O_152,N_2979,N_2978);
nor UO_153 (O_153,N_2952,N_2993);
and UO_154 (O_154,N_2997,N_2984);
nand UO_155 (O_155,N_2957,N_2955);
and UO_156 (O_156,N_2970,N_2952);
xnor UO_157 (O_157,N_2980,N_2957);
nor UO_158 (O_158,N_2994,N_2950);
or UO_159 (O_159,N_2997,N_2967);
and UO_160 (O_160,N_2952,N_2969);
and UO_161 (O_161,N_2982,N_2959);
nand UO_162 (O_162,N_2954,N_2994);
nor UO_163 (O_163,N_2966,N_2981);
nor UO_164 (O_164,N_2970,N_2971);
and UO_165 (O_165,N_2970,N_2973);
nor UO_166 (O_166,N_2969,N_2994);
nand UO_167 (O_167,N_2973,N_2957);
or UO_168 (O_168,N_2965,N_2981);
nand UO_169 (O_169,N_2953,N_2970);
or UO_170 (O_170,N_2972,N_2961);
or UO_171 (O_171,N_2964,N_2961);
nor UO_172 (O_172,N_2986,N_2956);
nand UO_173 (O_173,N_2978,N_2961);
and UO_174 (O_174,N_2973,N_2989);
or UO_175 (O_175,N_2955,N_2961);
nor UO_176 (O_176,N_2969,N_2984);
nor UO_177 (O_177,N_2955,N_2976);
or UO_178 (O_178,N_2960,N_2989);
nor UO_179 (O_179,N_2990,N_2975);
and UO_180 (O_180,N_2986,N_2969);
and UO_181 (O_181,N_2989,N_2988);
or UO_182 (O_182,N_2952,N_2988);
nor UO_183 (O_183,N_2975,N_2966);
nor UO_184 (O_184,N_2950,N_2974);
and UO_185 (O_185,N_2980,N_2954);
and UO_186 (O_186,N_2978,N_2992);
xnor UO_187 (O_187,N_2969,N_2980);
nand UO_188 (O_188,N_2956,N_2993);
and UO_189 (O_189,N_2956,N_2975);
or UO_190 (O_190,N_2954,N_2992);
xor UO_191 (O_191,N_2963,N_2950);
or UO_192 (O_192,N_2964,N_2984);
and UO_193 (O_193,N_2987,N_2972);
nor UO_194 (O_194,N_2957,N_2985);
and UO_195 (O_195,N_2957,N_2989);
nor UO_196 (O_196,N_2993,N_2972);
nand UO_197 (O_197,N_2987,N_2979);
and UO_198 (O_198,N_2951,N_2998);
and UO_199 (O_199,N_2975,N_2985);
nor UO_200 (O_200,N_2952,N_2975);
nor UO_201 (O_201,N_2958,N_2997);
and UO_202 (O_202,N_2965,N_2969);
nor UO_203 (O_203,N_2972,N_2974);
nor UO_204 (O_204,N_2983,N_2986);
and UO_205 (O_205,N_2956,N_2962);
and UO_206 (O_206,N_2973,N_2985);
and UO_207 (O_207,N_2985,N_2950);
and UO_208 (O_208,N_2955,N_2972);
or UO_209 (O_209,N_2993,N_2992);
nand UO_210 (O_210,N_2967,N_2964);
nor UO_211 (O_211,N_2992,N_2958);
nor UO_212 (O_212,N_2962,N_2972);
nand UO_213 (O_213,N_2950,N_2991);
or UO_214 (O_214,N_2957,N_2998);
nor UO_215 (O_215,N_2962,N_2995);
nand UO_216 (O_216,N_2966,N_2957);
nor UO_217 (O_217,N_2986,N_2970);
nand UO_218 (O_218,N_2999,N_2960);
nand UO_219 (O_219,N_2987,N_2998);
nor UO_220 (O_220,N_2999,N_2983);
or UO_221 (O_221,N_2988,N_2970);
nand UO_222 (O_222,N_2984,N_2998);
xnor UO_223 (O_223,N_2973,N_2956);
nand UO_224 (O_224,N_2979,N_2992);
and UO_225 (O_225,N_2994,N_2982);
and UO_226 (O_226,N_2952,N_2982);
and UO_227 (O_227,N_2998,N_2983);
and UO_228 (O_228,N_2966,N_2958);
nor UO_229 (O_229,N_2984,N_2992);
xnor UO_230 (O_230,N_2992,N_2986);
and UO_231 (O_231,N_2958,N_2962);
nor UO_232 (O_232,N_2979,N_2951);
nor UO_233 (O_233,N_2992,N_2995);
nand UO_234 (O_234,N_2950,N_2959);
or UO_235 (O_235,N_2983,N_2982);
or UO_236 (O_236,N_2975,N_2993);
nand UO_237 (O_237,N_2983,N_2955);
nand UO_238 (O_238,N_2957,N_2993);
nor UO_239 (O_239,N_2954,N_2959);
nand UO_240 (O_240,N_2990,N_2998);
and UO_241 (O_241,N_2983,N_2989);
nor UO_242 (O_242,N_2970,N_2974);
nor UO_243 (O_243,N_2990,N_2977);
nand UO_244 (O_244,N_2964,N_2998);
or UO_245 (O_245,N_2977,N_2987);
nor UO_246 (O_246,N_2955,N_2954);
nand UO_247 (O_247,N_2960,N_2998);
nand UO_248 (O_248,N_2956,N_2995);
or UO_249 (O_249,N_2980,N_2955);
nand UO_250 (O_250,N_2976,N_2956);
nor UO_251 (O_251,N_2994,N_2984);
or UO_252 (O_252,N_2983,N_2984);
and UO_253 (O_253,N_2995,N_2950);
or UO_254 (O_254,N_2985,N_2979);
nor UO_255 (O_255,N_2951,N_2953);
nor UO_256 (O_256,N_2988,N_2993);
nand UO_257 (O_257,N_2978,N_2995);
or UO_258 (O_258,N_2974,N_2980);
and UO_259 (O_259,N_2973,N_2963);
or UO_260 (O_260,N_2985,N_2955);
nor UO_261 (O_261,N_2953,N_2996);
nand UO_262 (O_262,N_2986,N_2988);
nand UO_263 (O_263,N_2966,N_2972);
nor UO_264 (O_264,N_2952,N_2998);
and UO_265 (O_265,N_2962,N_2985);
or UO_266 (O_266,N_2975,N_2969);
nor UO_267 (O_267,N_2966,N_2997);
nor UO_268 (O_268,N_2993,N_2962);
or UO_269 (O_269,N_2991,N_2981);
or UO_270 (O_270,N_2966,N_2992);
nand UO_271 (O_271,N_2967,N_2976);
or UO_272 (O_272,N_2961,N_2985);
or UO_273 (O_273,N_2986,N_2989);
or UO_274 (O_274,N_2993,N_2994);
or UO_275 (O_275,N_2962,N_2969);
nor UO_276 (O_276,N_2977,N_2981);
or UO_277 (O_277,N_2964,N_2952);
nand UO_278 (O_278,N_2992,N_2989);
nor UO_279 (O_279,N_2966,N_2973);
nand UO_280 (O_280,N_2983,N_2963);
nor UO_281 (O_281,N_2967,N_2973);
xnor UO_282 (O_282,N_2959,N_2960);
or UO_283 (O_283,N_2981,N_2956);
nand UO_284 (O_284,N_2959,N_2984);
nand UO_285 (O_285,N_2985,N_2954);
and UO_286 (O_286,N_2961,N_2994);
nand UO_287 (O_287,N_2989,N_2987);
xnor UO_288 (O_288,N_2978,N_2989);
or UO_289 (O_289,N_2994,N_2995);
and UO_290 (O_290,N_2997,N_2971);
and UO_291 (O_291,N_2990,N_2986);
and UO_292 (O_292,N_2970,N_2996);
nand UO_293 (O_293,N_2987,N_2959);
nand UO_294 (O_294,N_2973,N_2993);
nor UO_295 (O_295,N_2992,N_2952);
nand UO_296 (O_296,N_2974,N_2960);
and UO_297 (O_297,N_2951,N_2977);
and UO_298 (O_298,N_2977,N_2979);
nor UO_299 (O_299,N_2959,N_2962);
nand UO_300 (O_300,N_2973,N_2998);
nor UO_301 (O_301,N_2954,N_2991);
nand UO_302 (O_302,N_2964,N_2956);
and UO_303 (O_303,N_2974,N_2985);
and UO_304 (O_304,N_2998,N_2978);
or UO_305 (O_305,N_2965,N_2982);
nand UO_306 (O_306,N_2954,N_2988);
and UO_307 (O_307,N_2959,N_2998);
nand UO_308 (O_308,N_2957,N_2965);
nand UO_309 (O_309,N_2957,N_2956);
or UO_310 (O_310,N_2965,N_2962);
and UO_311 (O_311,N_2951,N_2989);
or UO_312 (O_312,N_2953,N_2973);
nand UO_313 (O_313,N_2996,N_2990);
nand UO_314 (O_314,N_2982,N_2955);
and UO_315 (O_315,N_2964,N_2991);
nor UO_316 (O_316,N_2994,N_2990);
nor UO_317 (O_317,N_2981,N_2950);
or UO_318 (O_318,N_2953,N_2960);
nor UO_319 (O_319,N_2988,N_2995);
and UO_320 (O_320,N_2985,N_2959);
nand UO_321 (O_321,N_2998,N_2963);
and UO_322 (O_322,N_2956,N_2996);
nand UO_323 (O_323,N_2974,N_2973);
nor UO_324 (O_324,N_2995,N_2957);
nand UO_325 (O_325,N_2980,N_2985);
nor UO_326 (O_326,N_2960,N_2968);
nor UO_327 (O_327,N_2974,N_2969);
nand UO_328 (O_328,N_2955,N_2952);
nor UO_329 (O_329,N_2976,N_2974);
or UO_330 (O_330,N_2998,N_2950);
xor UO_331 (O_331,N_2959,N_2967);
nand UO_332 (O_332,N_2997,N_2962);
or UO_333 (O_333,N_2965,N_2993);
or UO_334 (O_334,N_2988,N_2953);
or UO_335 (O_335,N_2965,N_2980);
nor UO_336 (O_336,N_2958,N_2961);
xnor UO_337 (O_337,N_2978,N_2977);
or UO_338 (O_338,N_2978,N_2956);
nor UO_339 (O_339,N_2979,N_2969);
nand UO_340 (O_340,N_2962,N_2982);
nand UO_341 (O_341,N_2973,N_2975);
or UO_342 (O_342,N_2994,N_2957);
nor UO_343 (O_343,N_2979,N_2960);
or UO_344 (O_344,N_2976,N_2964);
or UO_345 (O_345,N_2956,N_2979);
or UO_346 (O_346,N_2968,N_2954);
or UO_347 (O_347,N_2989,N_2982);
xor UO_348 (O_348,N_2991,N_2995);
and UO_349 (O_349,N_2959,N_2955);
nand UO_350 (O_350,N_2965,N_2953);
or UO_351 (O_351,N_2977,N_2988);
nand UO_352 (O_352,N_2990,N_2979);
nand UO_353 (O_353,N_2969,N_2966);
nand UO_354 (O_354,N_2968,N_2963);
nand UO_355 (O_355,N_2954,N_2976);
nor UO_356 (O_356,N_2958,N_2976);
and UO_357 (O_357,N_2981,N_2970);
nor UO_358 (O_358,N_2994,N_2955);
nor UO_359 (O_359,N_2990,N_2959);
nor UO_360 (O_360,N_2990,N_2953);
and UO_361 (O_361,N_2974,N_2989);
nand UO_362 (O_362,N_2983,N_2951);
and UO_363 (O_363,N_2991,N_2977);
or UO_364 (O_364,N_2993,N_2961);
xnor UO_365 (O_365,N_2978,N_2966);
nor UO_366 (O_366,N_2990,N_2997);
and UO_367 (O_367,N_2950,N_2996);
or UO_368 (O_368,N_2957,N_2953);
and UO_369 (O_369,N_2953,N_2978);
or UO_370 (O_370,N_2988,N_2972);
nand UO_371 (O_371,N_2952,N_2986);
nand UO_372 (O_372,N_2986,N_2958);
and UO_373 (O_373,N_2957,N_2991);
and UO_374 (O_374,N_2978,N_2997);
nand UO_375 (O_375,N_2966,N_2990);
xor UO_376 (O_376,N_2955,N_2991);
nand UO_377 (O_377,N_2976,N_2981);
nor UO_378 (O_378,N_2972,N_2994);
nand UO_379 (O_379,N_2995,N_2959);
nand UO_380 (O_380,N_2953,N_2958);
nor UO_381 (O_381,N_2971,N_2952);
nand UO_382 (O_382,N_2994,N_2977);
and UO_383 (O_383,N_2992,N_2988);
nand UO_384 (O_384,N_2983,N_2960);
nand UO_385 (O_385,N_2995,N_2999);
or UO_386 (O_386,N_2997,N_2979);
nand UO_387 (O_387,N_2953,N_2989);
and UO_388 (O_388,N_2971,N_2959);
and UO_389 (O_389,N_2981,N_2962);
nor UO_390 (O_390,N_2986,N_2950);
and UO_391 (O_391,N_2968,N_2972);
or UO_392 (O_392,N_2974,N_2997);
nand UO_393 (O_393,N_2994,N_2981);
nor UO_394 (O_394,N_2959,N_2996);
and UO_395 (O_395,N_2986,N_2971);
and UO_396 (O_396,N_2994,N_2966);
nor UO_397 (O_397,N_2956,N_2999);
nor UO_398 (O_398,N_2998,N_2974);
nand UO_399 (O_399,N_2962,N_2953);
or UO_400 (O_400,N_2964,N_2955);
and UO_401 (O_401,N_2967,N_2955);
or UO_402 (O_402,N_2950,N_2988);
or UO_403 (O_403,N_2998,N_2967);
or UO_404 (O_404,N_2972,N_2986);
nor UO_405 (O_405,N_2982,N_2966);
or UO_406 (O_406,N_2992,N_2975);
nand UO_407 (O_407,N_2975,N_2988);
nor UO_408 (O_408,N_2984,N_2990);
and UO_409 (O_409,N_2950,N_2954);
and UO_410 (O_410,N_2999,N_2987);
nor UO_411 (O_411,N_2961,N_2957);
nor UO_412 (O_412,N_2951,N_2991);
nand UO_413 (O_413,N_2980,N_2953);
nor UO_414 (O_414,N_2983,N_2976);
and UO_415 (O_415,N_2971,N_2980);
or UO_416 (O_416,N_2975,N_2983);
and UO_417 (O_417,N_2969,N_2971);
nor UO_418 (O_418,N_2960,N_2966);
xor UO_419 (O_419,N_2954,N_2981);
xnor UO_420 (O_420,N_2974,N_2952);
nor UO_421 (O_421,N_2961,N_2998);
nor UO_422 (O_422,N_2959,N_2986);
nand UO_423 (O_423,N_2981,N_2999);
and UO_424 (O_424,N_2976,N_2984);
nand UO_425 (O_425,N_2960,N_2972);
or UO_426 (O_426,N_2965,N_2975);
nor UO_427 (O_427,N_2999,N_2992);
and UO_428 (O_428,N_2951,N_2994);
and UO_429 (O_429,N_2969,N_2978);
and UO_430 (O_430,N_2991,N_2963);
or UO_431 (O_431,N_2976,N_2973);
xnor UO_432 (O_432,N_2994,N_2988);
nand UO_433 (O_433,N_2991,N_2997);
nand UO_434 (O_434,N_2972,N_2992);
nand UO_435 (O_435,N_2958,N_2957);
nand UO_436 (O_436,N_2965,N_2961);
or UO_437 (O_437,N_2980,N_2981);
and UO_438 (O_438,N_2990,N_2991);
nor UO_439 (O_439,N_2984,N_2978);
or UO_440 (O_440,N_2963,N_2979);
nand UO_441 (O_441,N_2960,N_2967);
nor UO_442 (O_442,N_2984,N_2981);
or UO_443 (O_443,N_2965,N_2984);
nor UO_444 (O_444,N_2951,N_2964);
nor UO_445 (O_445,N_2976,N_2972);
or UO_446 (O_446,N_2972,N_2982);
or UO_447 (O_447,N_2999,N_2989);
xnor UO_448 (O_448,N_2999,N_2998);
or UO_449 (O_449,N_2958,N_2983);
and UO_450 (O_450,N_2989,N_2961);
nor UO_451 (O_451,N_2958,N_2954);
and UO_452 (O_452,N_2988,N_2991);
nor UO_453 (O_453,N_2950,N_2987);
nand UO_454 (O_454,N_2979,N_2972);
nand UO_455 (O_455,N_2981,N_2964);
nand UO_456 (O_456,N_2962,N_2963);
and UO_457 (O_457,N_2997,N_2973);
nand UO_458 (O_458,N_2969,N_2990);
nand UO_459 (O_459,N_2966,N_2983);
or UO_460 (O_460,N_2993,N_2976);
xnor UO_461 (O_461,N_2979,N_2998);
and UO_462 (O_462,N_2999,N_2975);
and UO_463 (O_463,N_2986,N_2975);
or UO_464 (O_464,N_2980,N_2975);
nand UO_465 (O_465,N_2978,N_2960);
and UO_466 (O_466,N_2958,N_2964);
or UO_467 (O_467,N_2986,N_2974);
or UO_468 (O_468,N_2950,N_2993);
or UO_469 (O_469,N_2965,N_2956);
and UO_470 (O_470,N_2992,N_2990);
nand UO_471 (O_471,N_2995,N_2974);
nor UO_472 (O_472,N_2992,N_2963);
or UO_473 (O_473,N_2989,N_2958);
nand UO_474 (O_474,N_2990,N_2972);
or UO_475 (O_475,N_2985,N_2998);
and UO_476 (O_476,N_2987,N_2956);
or UO_477 (O_477,N_2977,N_2972);
nor UO_478 (O_478,N_2981,N_2960);
nand UO_479 (O_479,N_2970,N_2987);
and UO_480 (O_480,N_2951,N_2950);
nand UO_481 (O_481,N_2954,N_2970);
nand UO_482 (O_482,N_2986,N_2979);
nand UO_483 (O_483,N_2971,N_2990);
or UO_484 (O_484,N_2986,N_2964);
and UO_485 (O_485,N_2997,N_2988);
and UO_486 (O_486,N_2989,N_2950);
nor UO_487 (O_487,N_2967,N_2988);
or UO_488 (O_488,N_2983,N_2952);
nor UO_489 (O_489,N_2968,N_2980);
nand UO_490 (O_490,N_2951,N_2973);
nand UO_491 (O_491,N_2998,N_2981);
nand UO_492 (O_492,N_2971,N_2966);
nor UO_493 (O_493,N_2995,N_2975);
or UO_494 (O_494,N_2977,N_2961);
nor UO_495 (O_495,N_2950,N_2958);
nor UO_496 (O_496,N_2971,N_2958);
nor UO_497 (O_497,N_2982,N_2987);
and UO_498 (O_498,N_2994,N_2968);
nor UO_499 (O_499,N_2976,N_2953);
endmodule