module basic_3000_30000_3500_3_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20001,N_20005,N_20006,N_20007,N_20008,N_20009,N_20012,N_20013,N_20014,N_20017,N_20018,N_20020,N_20021,N_20024,N_20025,N_20026,N_20028,N_20030,N_20032,N_20033,N_20034,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20060,N_20061,N_20063,N_20064,N_20066,N_20067,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20078,N_20080,N_20082,N_20083,N_20084,N_20086,N_20087,N_20089,N_20090,N_20092,N_20094,N_20095,N_20096,N_20100,N_20101,N_20102,N_20104,N_20105,N_20106,N_20107,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20119,N_20120,N_20121,N_20122,N_20123,N_20125,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20136,N_20137,N_20138,N_20139,N_20140,N_20143,N_20145,N_20146,N_20150,N_20151,N_20152,N_20154,N_20155,N_20157,N_20158,N_20159,N_20160,N_20162,N_20164,N_20165,N_20166,N_20167,N_20169,N_20170,N_20172,N_20173,N_20174,N_20178,N_20179,N_20183,N_20184,N_20185,N_20186,N_20187,N_20190,N_20192,N_20193,N_20194,N_20195,N_20199,N_20200,N_20201,N_20202,N_20203,N_20206,N_20207,N_20208,N_20212,N_20215,N_20216,N_20219,N_20220,N_20222,N_20224,N_20225,N_20227,N_20228,N_20229,N_20231,N_20232,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20244,N_20248,N_20249,N_20250,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20259,N_20260,N_20261,N_20262,N_20263,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20286,N_20288,N_20290,N_20291,N_20292,N_20293,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20305,N_20306,N_20308,N_20309,N_20310,N_20312,N_20313,N_20314,N_20316,N_20318,N_20319,N_20320,N_20322,N_20323,N_20324,N_20327,N_20328,N_20330,N_20331,N_20332,N_20334,N_20335,N_20337,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20364,N_20367,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20379,N_20380,N_20382,N_20383,N_20384,N_20385,N_20386,N_20388,N_20389,N_20391,N_20394,N_20395,N_20396,N_20397,N_20399,N_20400,N_20402,N_20404,N_20406,N_20407,N_20409,N_20411,N_20412,N_20414,N_20415,N_20417,N_20418,N_20419,N_20420,N_20421,N_20424,N_20426,N_20427,N_20428,N_20429,N_20430,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20442,N_20444,N_20445,N_20448,N_20450,N_20451,N_20452,N_20455,N_20456,N_20457,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20472,N_20474,N_20475,N_20476,N_20477,N_20478,N_20480,N_20482,N_20483,N_20484,N_20485,N_20486,N_20488,N_20490,N_20491,N_20492,N_20495,N_20496,N_20497,N_20498,N_20500,N_20501,N_20502,N_20503,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20517,N_20519,N_20520,N_20522,N_20527,N_20528,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20537,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20547,N_20550,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20566,N_20567,N_20568,N_20570,N_20571,N_20572,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20587,N_20588,N_20590,N_20592,N_20594,N_20595,N_20597,N_20598,N_20600,N_20601,N_20603,N_20604,N_20605,N_20607,N_20609,N_20611,N_20612,N_20614,N_20616,N_20617,N_20618,N_20620,N_20621,N_20622,N_20624,N_20625,N_20626,N_20627,N_20628,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20638,N_20644,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20656,N_20657,N_20658,N_20659,N_20660,N_20662,N_20663,N_20664,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20676,N_20678,N_20679,N_20681,N_20682,N_20686,N_20687,N_20689,N_20692,N_20693,N_20696,N_20698,N_20700,N_20701,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20712,N_20717,N_20718,N_20720,N_20722,N_20723,N_20724,N_20726,N_20727,N_20730,N_20733,N_20735,N_20737,N_20739,N_20740,N_20741,N_20742,N_20745,N_20746,N_20748,N_20749,N_20750,N_20752,N_20753,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20762,N_20764,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20777,N_20778,N_20779,N_20780,N_20782,N_20784,N_20785,N_20789,N_20792,N_20793,N_20794,N_20795,N_20796,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20817,N_20819,N_20820,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20857,N_20858,N_20859,N_20862,N_20864,N_20865,N_20866,N_20867,N_20870,N_20871,N_20874,N_20876,N_20877,N_20878,N_20880,N_20881,N_20882,N_20883,N_20884,N_20886,N_20887,N_20888,N_20889,N_20890,N_20892,N_20893,N_20894,N_20899,N_20900,N_20901,N_20905,N_20906,N_20907,N_20909,N_20910,N_20911,N_20913,N_20914,N_20915,N_20916,N_20917,N_20919,N_20920,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20931,N_20933,N_20934,N_20935,N_20937,N_20938,N_20939,N_20940,N_20943,N_20944,N_20945,N_20946,N_20947,N_20949,N_20950,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20970,N_20971,N_20972,N_20973,N_20976,N_20978,N_20979,N_20981,N_20982,N_20983,N_20985,N_20986,N_20987,N_20988,N_20989,N_20991,N_20992,N_20994,N_20995,N_20996,N_20997,N_20999,N_21001,N_21004,N_21005,N_21006,N_21007,N_21008,N_21012,N_21013,N_21014,N_21015,N_21016,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21032,N_21034,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21046,N_21047,N_21048,N_21049,N_21050,N_21052,N_21054,N_21055,N_21058,N_21060,N_21061,N_21062,N_21063,N_21064,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21076,N_21078,N_21079,N_21080,N_21081,N_21084,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21104,N_21105,N_21106,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21115,N_21116,N_21121,N_21122,N_21123,N_21125,N_21126,N_21127,N_21129,N_21132,N_21133,N_21135,N_21138,N_21139,N_21140,N_21141,N_21143,N_21144,N_21145,N_21148,N_21149,N_21150,N_21151,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21183,N_21184,N_21185,N_21186,N_21188,N_21189,N_21192,N_21193,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21206,N_21208,N_21211,N_21212,N_21214,N_21216,N_21217,N_21218,N_21219,N_21220,N_21223,N_21224,N_21225,N_21228,N_21229,N_21231,N_21233,N_21234,N_21235,N_21237,N_21239,N_21240,N_21241,N_21242,N_21243,N_21246,N_21247,N_21248,N_21250,N_21251,N_21253,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21269,N_21270,N_21271,N_21272,N_21275,N_21276,N_21277,N_21278,N_21279,N_21281,N_21282,N_21283,N_21284,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21295,N_21296,N_21297,N_21300,N_21302,N_21303,N_21304,N_21306,N_21307,N_21308,N_21309,N_21311,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21322,N_21323,N_21324,N_21325,N_21327,N_21328,N_21332,N_21333,N_21334,N_21335,N_21338,N_21339,N_21340,N_21341,N_21343,N_21344,N_21345,N_21346,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21362,N_21364,N_21366,N_21368,N_21369,N_21370,N_21372,N_21374,N_21376,N_21377,N_21378,N_21379,N_21381,N_21384,N_21385,N_21387,N_21388,N_21390,N_21392,N_21393,N_21394,N_21398,N_21401,N_21402,N_21403,N_21404,N_21405,N_21408,N_21410,N_21411,N_21412,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21425,N_21426,N_21427,N_21428,N_21429,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21441,N_21444,N_21445,N_21446,N_21447,N_21450,N_21451,N_21453,N_21454,N_21456,N_21458,N_21462,N_21463,N_21466,N_21467,N_21468,N_21470,N_21471,N_21473,N_21474,N_21475,N_21477,N_21478,N_21480,N_21481,N_21483,N_21484,N_21485,N_21486,N_21489,N_21492,N_21494,N_21495,N_21497,N_21498,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21521,N_21523,N_21524,N_21528,N_21529,N_21530,N_21532,N_21534,N_21535,N_21536,N_21538,N_21540,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21550,N_21552,N_21553,N_21555,N_21556,N_21558,N_21559,N_21561,N_21562,N_21563,N_21564,N_21566,N_21567,N_21568,N_21569,N_21571,N_21573,N_21574,N_21575,N_21576,N_21577,N_21580,N_21581,N_21582,N_21583,N_21584,N_21586,N_21589,N_21590,N_21591,N_21592,N_21593,N_21595,N_21596,N_21597,N_21598,N_21599,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21611,N_21612,N_21613,N_21614,N_21615,N_21617,N_21618,N_21621,N_21622,N_21624,N_21626,N_21628,N_21629,N_21630,N_21631,N_21635,N_21636,N_21637,N_21638,N_21640,N_21643,N_21645,N_21646,N_21647,N_21649,N_21650,N_21651,N_21653,N_21655,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21664,N_21665,N_21666,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21686,N_21688,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21709,N_21710,N_21711,N_21712,N_21713,N_21715,N_21716,N_21717,N_21719,N_21722,N_21725,N_21728,N_21729,N_21730,N_21731,N_21732,N_21735,N_21736,N_21737,N_21738,N_21740,N_21741,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21754,N_21755,N_21756,N_21757,N_21759,N_21760,N_21761,N_21762,N_21764,N_21768,N_21770,N_21772,N_21774,N_21777,N_21778,N_21780,N_21781,N_21783,N_21788,N_21790,N_21791,N_21793,N_21794,N_21795,N_21796,N_21797,N_21800,N_21802,N_21803,N_21806,N_21807,N_21808,N_21809,N_21811,N_21812,N_21813,N_21814,N_21815,N_21817,N_21818,N_21819,N_21822,N_21823,N_21826,N_21827,N_21828,N_21830,N_21831,N_21832,N_21834,N_21835,N_21836,N_21838,N_21839,N_21842,N_21843,N_21844,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21853,N_21855,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21865,N_21866,N_21867,N_21868,N_21869,N_21871,N_21875,N_21877,N_21878,N_21880,N_21881,N_21882,N_21883,N_21884,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21894,N_21895,N_21896,N_21897,N_21898,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21915,N_21917,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21928,N_21929,N_21930,N_21931,N_21932,N_21934,N_21938,N_21940,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21952,N_21953,N_21954,N_21957,N_21958,N_21959,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21971,N_21972,N_21974,N_21975,N_21976,N_21977,N_21978,N_21982,N_21983,N_21984,N_21985,N_21986,N_21988,N_21989,N_21991,N_21993,N_21994,N_21995,N_21997,N_21998,N_22000,N_22001,N_22002,N_22007,N_22008,N_22011,N_22012,N_22014,N_22015,N_22017,N_22022,N_22023,N_22024,N_22026,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22049,N_22053,N_22054,N_22057,N_22058,N_22060,N_22061,N_22063,N_22064,N_22065,N_22066,N_22068,N_22069,N_22070,N_22071,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22090,N_22092,N_22093,N_22094,N_22095,N_22097,N_22098,N_22100,N_22102,N_22103,N_22104,N_22105,N_22106,N_22108,N_22109,N_22111,N_22113,N_22114,N_22115,N_22118,N_22119,N_22120,N_22122,N_22123,N_22124,N_22125,N_22126,N_22129,N_22130,N_22131,N_22133,N_22136,N_22137,N_22138,N_22140,N_22141,N_22143,N_22144,N_22145,N_22146,N_22148,N_22149,N_22150,N_22151,N_22153,N_22155,N_22159,N_22160,N_22162,N_22163,N_22164,N_22166,N_22167,N_22168,N_22169,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22180,N_22182,N_22183,N_22184,N_22185,N_22188,N_22189,N_22194,N_22196,N_22197,N_22198,N_22199,N_22200,N_22202,N_22204,N_22205,N_22206,N_22207,N_22210,N_22211,N_22212,N_22213,N_22214,N_22216,N_22217,N_22219,N_22220,N_22221,N_22227,N_22229,N_22230,N_22236,N_22237,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22249,N_22252,N_22253,N_22255,N_22256,N_22258,N_22259,N_22260,N_22262,N_22263,N_22265,N_22267,N_22268,N_22269,N_22271,N_22275,N_22277,N_22278,N_22279,N_22280,N_22283,N_22284,N_22285,N_22286,N_22290,N_22291,N_22292,N_22294,N_22295,N_22296,N_22298,N_22299,N_22301,N_22302,N_22305,N_22306,N_22307,N_22309,N_22311,N_22313,N_22314,N_22315,N_22316,N_22317,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22327,N_22330,N_22331,N_22333,N_22334,N_22335,N_22336,N_22340,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22351,N_22352,N_22353,N_22354,N_22356,N_22357,N_22359,N_22361,N_22362,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22372,N_22373,N_22375,N_22376,N_22378,N_22379,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22388,N_22389,N_22390,N_22391,N_22392,N_22395,N_22396,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22411,N_22414,N_22416,N_22417,N_22421,N_22423,N_22424,N_22425,N_22427,N_22428,N_22429,N_22432,N_22433,N_22434,N_22435,N_22437,N_22438,N_22440,N_22443,N_22444,N_22446,N_22447,N_22449,N_22451,N_22452,N_22453,N_22454,N_22455,N_22457,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22468,N_22469,N_22471,N_22474,N_22475,N_22476,N_22478,N_22479,N_22480,N_22483,N_22485,N_22486,N_22488,N_22491,N_22492,N_22493,N_22495,N_22497,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22506,N_22508,N_22510,N_22511,N_22512,N_22513,N_22514,N_22516,N_22517,N_22518,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22528,N_22529,N_22533,N_22534,N_22535,N_22536,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22549,N_22550,N_22552,N_22553,N_22555,N_22556,N_22558,N_22559,N_22560,N_22562,N_22565,N_22566,N_22568,N_22569,N_22571,N_22572,N_22573,N_22574,N_22575,N_22577,N_22578,N_22580,N_22581,N_22582,N_22584,N_22585,N_22586,N_22589,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22611,N_22615,N_22616,N_22617,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22634,N_22636,N_22639,N_22641,N_22643,N_22644,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22653,N_22654,N_22656,N_22657,N_22658,N_22659,N_22660,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22678,N_22679,N_22680,N_22682,N_22683,N_22684,N_22685,N_22687,N_22688,N_22689,N_22690,N_22692,N_22694,N_22695,N_22697,N_22700,N_22701,N_22704,N_22707,N_22709,N_22711,N_22712,N_22713,N_22714,N_22715,N_22718,N_22719,N_22720,N_22721,N_22722,N_22724,N_22725,N_22726,N_22728,N_22729,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22739,N_22740,N_22741,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22758,N_22761,N_22762,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22772,N_22773,N_22775,N_22777,N_22779,N_22781,N_22782,N_22783,N_22784,N_22786,N_22787,N_22788,N_22789,N_22790,N_22792,N_22795,N_22796,N_22797,N_22799,N_22800,N_22801,N_22803,N_22805,N_22807,N_22808,N_22809,N_22810,N_22812,N_22813,N_22814,N_22816,N_22817,N_22819,N_22820,N_22824,N_22826,N_22827,N_22829,N_22832,N_22834,N_22835,N_22837,N_22838,N_22839,N_22842,N_22843,N_22844,N_22846,N_22848,N_22849,N_22850,N_22851,N_22852,N_22854,N_22855,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22865,N_22866,N_22867,N_22869,N_22870,N_22872,N_22873,N_22874,N_22875,N_22877,N_22878,N_22879,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22888,N_22890,N_22891,N_22892,N_22893,N_22894,N_22896,N_22897,N_22898,N_22900,N_22901,N_22902,N_22903,N_22905,N_22906,N_22909,N_22910,N_22911,N_22912,N_22913,N_22915,N_22917,N_22918,N_22919,N_22920,N_22921,N_22923,N_22924,N_22926,N_22927,N_22928,N_22930,N_22931,N_22932,N_22934,N_22936,N_22938,N_22939,N_22940,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22951,N_22952,N_22955,N_22957,N_22958,N_22959,N_22960,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22971,N_22972,N_22975,N_22977,N_22979,N_22981,N_22982,N_22984,N_22986,N_22990,N_22991,N_22992,N_22993,N_22995,N_22996,N_22997,N_22998,N_22999,N_23001,N_23002,N_23003,N_23004,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23016,N_23017,N_23019,N_23020,N_23022,N_23024,N_23025,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23043,N_23050,N_23051,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23070,N_23071,N_23073,N_23075,N_23076,N_23077,N_23079,N_23080,N_23081,N_23082,N_23083,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23097,N_23098,N_23101,N_23102,N_23103,N_23104,N_23107,N_23108,N_23109,N_23111,N_23113,N_23114,N_23115,N_23117,N_23118,N_23119,N_23121,N_23122,N_23126,N_23128,N_23130,N_23132,N_23133,N_23134,N_23135,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23147,N_23148,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23157,N_23158,N_23161,N_23162,N_23164,N_23165,N_23166,N_23169,N_23170,N_23173,N_23174,N_23175,N_23177,N_23179,N_23180,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23191,N_23192,N_23193,N_23195,N_23197,N_23198,N_23199,N_23200,N_23203,N_23205,N_23207,N_23208,N_23210,N_23211,N_23212,N_23213,N_23214,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23224,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23237,N_23238,N_23239,N_23240,N_23241,N_23244,N_23245,N_23248,N_23250,N_23251,N_23253,N_23254,N_23255,N_23256,N_23259,N_23260,N_23262,N_23264,N_23265,N_23266,N_23268,N_23271,N_23273,N_23275,N_23276,N_23277,N_23278,N_23280,N_23282,N_23286,N_23287,N_23288,N_23289,N_23290,N_23292,N_23293,N_23294,N_23295,N_23297,N_23298,N_23299,N_23300,N_23302,N_23303,N_23304,N_23305,N_23308,N_23309,N_23310,N_23311,N_23313,N_23315,N_23316,N_23317,N_23320,N_23321,N_23322,N_23323,N_23325,N_23326,N_23327,N_23330,N_23331,N_23334,N_23335,N_23338,N_23339,N_23340,N_23341,N_23342,N_23344,N_23345,N_23346,N_23347,N_23349,N_23350,N_23352,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23369,N_23371,N_23372,N_23374,N_23375,N_23376,N_23377,N_23378,N_23381,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23391,N_23393,N_23397,N_23398,N_23399,N_23400,N_23401,N_23403,N_23404,N_23406,N_23408,N_23409,N_23410,N_23411,N_23412,N_23415,N_23416,N_23418,N_23419,N_23421,N_23423,N_23424,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23448,N_23449,N_23450,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23460,N_23461,N_23465,N_23466,N_23467,N_23468,N_23470,N_23472,N_23473,N_23477,N_23478,N_23480,N_23481,N_23483,N_23484,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23496,N_23497,N_23499,N_23501,N_23502,N_23503,N_23506,N_23508,N_23509,N_23510,N_23512,N_23513,N_23514,N_23517,N_23518,N_23519,N_23520,N_23522,N_23523,N_23525,N_23526,N_23529,N_23530,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23540,N_23541,N_23542,N_23543,N_23545,N_23546,N_23547,N_23548,N_23549,N_23551,N_23553,N_23554,N_23555,N_23556,N_23558,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23568,N_23570,N_23571,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23582,N_23583,N_23584,N_23585,N_23586,N_23588,N_23589,N_23590,N_23591,N_23593,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23602,N_23603,N_23604,N_23606,N_23609,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23619,N_23621,N_23623,N_23624,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23635,N_23636,N_23640,N_23642,N_23644,N_23646,N_23647,N_23648,N_23649,N_23652,N_23654,N_23655,N_23656,N_23658,N_23659,N_23660,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23683,N_23684,N_23685,N_23687,N_23691,N_23692,N_23695,N_23696,N_23697,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23706,N_23707,N_23708,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23726,N_23727,N_23732,N_23737,N_23738,N_23739,N_23740,N_23741,N_23743,N_23744,N_23746,N_23747,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23756,N_23757,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23767,N_23768,N_23770,N_23772,N_23773,N_23774,N_23776,N_23777,N_23778,N_23780,N_23784,N_23786,N_23787,N_23788,N_23789,N_23791,N_23793,N_23794,N_23796,N_23797,N_23798,N_23800,N_23801,N_23803,N_23809,N_23811,N_23812,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23822,N_23823,N_23826,N_23827,N_23828,N_23829,N_23831,N_23833,N_23834,N_23836,N_23837,N_23838,N_23840,N_23842,N_23844,N_23847,N_23848,N_23850,N_23851,N_23852,N_23853,N_23855,N_23856,N_23858,N_23860,N_23861,N_23862,N_23863,N_23866,N_23867,N_23868,N_23870,N_23872,N_23875,N_23877,N_23878,N_23881,N_23883,N_23884,N_23886,N_23887,N_23888,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23921,N_23922,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23948,N_23950,N_23951,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23961,N_23962,N_23967,N_23968,N_23969,N_23972,N_23973,N_23975,N_23977,N_23978,N_23980,N_23981,N_23983,N_23985,N_23988,N_23989,N_23992,N_23993,N_23995,N_23996,N_23999,N_24000,N_24001,N_24004,N_24005,N_24007,N_24008,N_24013,N_24014,N_24015,N_24016,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24027,N_24028,N_24031,N_24035,N_24036,N_24038,N_24039,N_24041,N_24042,N_24043,N_24044,N_24045,N_24047,N_24048,N_24049,N_24050,N_24052,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24063,N_24065,N_24067,N_24068,N_24070,N_24071,N_24072,N_24073,N_24075,N_24076,N_24077,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24087,N_24088,N_24089,N_24091,N_24092,N_24094,N_24095,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24107,N_24109,N_24110,N_24111,N_24112,N_24115,N_24116,N_24117,N_24121,N_24123,N_24125,N_24126,N_24127,N_24128,N_24130,N_24131,N_24132,N_24133,N_24134,N_24136,N_24137,N_24138,N_24140,N_24141,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24152,N_24153,N_24154,N_24155,N_24156,N_24158,N_24159,N_24162,N_24163,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24174,N_24175,N_24176,N_24178,N_24179,N_24180,N_24182,N_24183,N_24186,N_24187,N_24190,N_24191,N_24192,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24202,N_24205,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24218,N_24220,N_24221,N_24222,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24232,N_24234,N_24236,N_24237,N_24238,N_24239,N_24241,N_24244,N_24246,N_24247,N_24248,N_24249,N_24251,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24262,N_24263,N_24265,N_24266,N_24269,N_24270,N_24271,N_24272,N_24273,N_24275,N_24276,N_24277,N_24278,N_24279,N_24281,N_24285,N_24286,N_24287,N_24288,N_24290,N_24291,N_24292,N_24294,N_24295,N_24296,N_24297,N_24299,N_24301,N_24302,N_24303,N_24304,N_24306,N_24307,N_24308,N_24309,N_24313,N_24314,N_24315,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24326,N_24328,N_24330,N_24332,N_24333,N_24334,N_24336,N_24337,N_24339,N_24340,N_24342,N_24343,N_24344,N_24350,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24368,N_24372,N_24373,N_24374,N_24378,N_24379,N_24380,N_24382,N_24383,N_24385,N_24386,N_24390,N_24391,N_24392,N_24395,N_24396,N_24399,N_24401,N_24402,N_24403,N_24404,N_24405,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24414,N_24415,N_24417,N_24418,N_24419,N_24420,N_24422,N_24425,N_24426,N_24427,N_24428,N_24431,N_24433,N_24434,N_24436,N_24438,N_24443,N_24444,N_24445,N_24446,N_24447,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24460,N_24461,N_24463,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24489,N_24490,N_24491,N_24493,N_24495,N_24496,N_24498,N_24499,N_24501,N_24502,N_24503,N_24505,N_24507,N_24508,N_24510,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24519,N_24520,N_24521,N_24523,N_24524,N_24525,N_24526,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24554,N_24555,N_24557,N_24559,N_24560,N_24562,N_24565,N_24567,N_24569,N_24570,N_24571,N_24572,N_24576,N_24579,N_24580,N_24581,N_24582,N_24583,N_24586,N_24587,N_24588,N_24589,N_24590,N_24592,N_24593,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24614,N_24617,N_24618,N_24619,N_24621,N_24623,N_24627,N_24629,N_24631,N_24634,N_24635,N_24636,N_24638,N_24639,N_24641,N_24642,N_24643,N_24644,N_24646,N_24648,N_24652,N_24654,N_24655,N_24656,N_24658,N_24659,N_24660,N_24663,N_24664,N_24665,N_24667,N_24669,N_24671,N_24672,N_24674,N_24677,N_24679,N_24680,N_24681,N_24683,N_24685,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24705,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24733,N_24735,N_24736,N_24740,N_24741,N_24743,N_24744,N_24745,N_24749,N_24750,N_24753,N_24754,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24766,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24776,N_24777,N_24778,N_24781,N_24782,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24803,N_24804,N_24805,N_24807,N_24808,N_24809,N_24811,N_24813,N_24817,N_24818,N_24819,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24832,N_24833,N_24834,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24846,N_24847,N_24848,N_24849,N_24851,N_24852,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24862,N_24863,N_24865,N_24867,N_24869,N_24871,N_24873,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24890,N_24891,N_24894,N_24895,N_24896,N_24898,N_24901,N_24902,N_24905,N_24907,N_24908,N_24909,N_24910,N_24911,N_24913,N_24914,N_24915,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24929,N_24932,N_24933,N_24935,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24950,N_24951,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24964,N_24965,N_24967,N_24968,N_24969,N_24970,N_24973,N_24975,N_24976,N_24977,N_24979,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24991,N_24992,N_24993,N_24995,N_24996,N_24998,N_24999,N_25000,N_25003,N_25004,N_25005,N_25007,N_25008,N_25009,N_25010,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25028,N_25029,N_25030,N_25031,N_25032,N_25034,N_25035,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25046,N_25047,N_25048,N_25049,N_25050,N_25053,N_25055,N_25056,N_25058,N_25059,N_25061,N_25062,N_25065,N_25066,N_25067,N_25069,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25080,N_25082,N_25084,N_25085,N_25087,N_25088,N_25089,N_25090,N_25092,N_25093,N_25094,N_25095,N_25096,N_25098,N_25099,N_25100,N_25102,N_25103,N_25107,N_25108,N_25109,N_25110,N_25111,N_25113,N_25114,N_25116,N_25117,N_25118,N_25119,N_25120,N_25122,N_25123,N_25124,N_25125,N_25126,N_25128,N_25129,N_25130,N_25131,N_25132,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25166,N_25167,N_25168,N_25170,N_25171,N_25172,N_25174,N_25175,N_25176,N_25178,N_25179,N_25182,N_25183,N_25184,N_25185,N_25187,N_25188,N_25189,N_25190,N_25192,N_25194,N_25195,N_25196,N_25197,N_25199,N_25200,N_25201,N_25204,N_25205,N_25206,N_25212,N_25214,N_25215,N_25217,N_25218,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25230,N_25231,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25241,N_25242,N_25244,N_25245,N_25246,N_25248,N_25249,N_25250,N_25252,N_25253,N_25255,N_25256,N_25257,N_25259,N_25260,N_25262,N_25263,N_25265,N_25267,N_25269,N_25270,N_25271,N_25272,N_25274,N_25277,N_25279,N_25280,N_25281,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25293,N_25294,N_25296,N_25297,N_25298,N_25300,N_25302,N_25303,N_25304,N_25306,N_25308,N_25309,N_25312,N_25313,N_25315,N_25316,N_25317,N_25320,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25330,N_25331,N_25332,N_25333,N_25334,N_25337,N_25338,N_25339,N_25341,N_25342,N_25343,N_25344,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25355,N_25356,N_25358,N_25359,N_25360,N_25361,N_25363,N_25364,N_25365,N_25366,N_25367,N_25369,N_25370,N_25371,N_25373,N_25374,N_25376,N_25377,N_25378,N_25379,N_25380,N_25382,N_25385,N_25386,N_25388,N_25389,N_25391,N_25392,N_25393,N_25394,N_25396,N_25397,N_25398,N_25399,N_25402,N_25403,N_25406,N_25407,N_25408,N_25409,N_25410,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25419,N_25420,N_25423,N_25424,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25436,N_25437,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25448,N_25449,N_25450,N_25451,N_25452,N_25454,N_25456,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25470,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25481,N_25483,N_25485,N_25486,N_25489,N_25493,N_25495,N_25496,N_25497,N_25498,N_25500,N_25503,N_25505,N_25508,N_25511,N_25512,N_25515,N_25516,N_25517,N_25518,N_25520,N_25521,N_25522,N_25523,N_25526,N_25528,N_25530,N_25531,N_25533,N_25536,N_25537,N_25538,N_25540,N_25544,N_25545,N_25547,N_25548,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25567,N_25569,N_25570,N_25571,N_25573,N_25575,N_25576,N_25577,N_25579,N_25581,N_25583,N_25584,N_25585,N_25586,N_25589,N_25590,N_25591,N_25592,N_25594,N_25595,N_25596,N_25597,N_25599,N_25601,N_25602,N_25603,N_25604,N_25605,N_25608,N_25610,N_25611,N_25612,N_25613,N_25615,N_25617,N_25618,N_25619,N_25620,N_25621,N_25623,N_25625,N_25626,N_25627,N_25629,N_25630,N_25631,N_25632,N_25635,N_25636,N_25640,N_25641,N_25642,N_25645,N_25646,N_25647,N_25651,N_25652,N_25653,N_25654,N_25655,N_25658,N_25659,N_25660,N_25663,N_25664,N_25665,N_25666,N_25668,N_25669,N_25670,N_25671,N_25674,N_25675,N_25676,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25687,N_25689,N_25691,N_25693,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25707,N_25710,N_25713,N_25714,N_25715,N_25716,N_25718,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25735,N_25741,N_25742,N_25744,N_25746,N_25747,N_25750,N_25751,N_25752,N_25755,N_25756,N_25758,N_25759,N_25760,N_25762,N_25764,N_25765,N_25767,N_25768,N_25769,N_25770,N_25772,N_25773,N_25775,N_25776,N_25777,N_25778,N_25779,N_25781,N_25782,N_25783,N_25784,N_25785,N_25788,N_25789,N_25790,N_25791,N_25793,N_25794,N_25795,N_25796,N_25797,N_25799,N_25800,N_25801,N_25802,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25812,N_25813,N_25814,N_25816,N_25817,N_25818,N_25819,N_25821,N_25822,N_25823,N_25825,N_25827,N_25828,N_25829,N_25830,N_25831,N_25833,N_25836,N_25837,N_25838,N_25840,N_25841,N_25844,N_25846,N_25847,N_25851,N_25852,N_25853,N_25855,N_25856,N_25858,N_25859,N_25860,N_25862,N_25863,N_25864,N_25866,N_25867,N_25868,N_25869,N_25871,N_25872,N_25876,N_25877,N_25878,N_25880,N_25881,N_25882,N_25885,N_25886,N_25889,N_25890,N_25891,N_25892,N_25893,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25910,N_25912,N_25915,N_25916,N_25917,N_25919,N_25921,N_25922,N_25924,N_25926,N_25929,N_25932,N_25933,N_25934,N_25935,N_25937,N_25939,N_25941,N_25942,N_25945,N_25946,N_25947,N_25948,N_25949,N_25951,N_25952,N_25953,N_25954,N_25957,N_25958,N_25959,N_25960,N_25961,N_25963,N_25964,N_25965,N_25966,N_25967,N_25970,N_25972,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25985,N_25986,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25999,N_26000,N_26001,N_26003,N_26005,N_26006,N_26007,N_26009,N_26010,N_26011,N_26013,N_26014,N_26015,N_26017,N_26020,N_26022,N_26023,N_26024,N_26025,N_26028,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26038,N_26039,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26051,N_26052,N_26053,N_26054,N_26056,N_26058,N_26061,N_26062,N_26063,N_26065,N_26066,N_26069,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26080,N_26081,N_26082,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26092,N_26093,N_26094,N_26096,N_26097,N_26100,N_26103,N_26104,N_26106,N_26107,N_26108,N_26109,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26124,N_26128,N_26129,N_26131,N_26132,N_26133,N_26134,N_26135,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26147,N_26149,N_26151,N_26152,N_26153,N_26155,N_26156,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26166,N_26167,N_26169,N_26170,N_26171,N_26173,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26187,N_26188,N_26189,N_26190,N_26191,N_26193,N_26194,N_26195,N_26197,N_26198,N_26199,N_26200,N_26201,N_26203,N_26204,N_26206,N_26207,N_26209,N_26210,N_26212,N_26213,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26225,N_26226,N_26229,N_26230,N_26232,N_26234,N_26237,N_26239,N_26241,N_26242,N_26243,N_26244,N_26246,N_26247,N_26248,N_26249,N_26250,N_26252,N_26253,N_26254,N_26255,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26266,N_26267,N_26268,N_26269,N_26271,N_26272,N_26273,N_26274,N_26275,N_26277,N_26279,N_26281,N_26282,N_26284,N_26286,N_26290,N_26291,N_26292,N_26293,N_26295,N_26297,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26310,N_26311,N_26312,N_26315,N_26317,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26331,N_26333,N_26334,N_26336,N_26341,N_26342,N_26345,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26355,N_26358,N_26359,N_26361,N_26362,N_26363,N_26364,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26377,N_26379,N_26380,N_26382,N_26383,N_26385,N_26386,N_26388,N_26389,N_26390,N_26391,N_26394,N_26395,N_26396,N_26400,N_26401,N_26402,N_26405,N_26407,N_26409,N_26410,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26420,N_26421,N_26423,N_26425,N_26427,N_26429,N_26430,N_26431,N_26432,N_26434,N_26436,N_26437,N_26438,N_26439,N_26440,N_26442,N_26444,N_26445,N_26447,N_26450,N_26451,N_26452,N_26455,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26465,N_26466,N_26467,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26478,N_26479,N_26480,N_26481,N_26482,N_26485,N_26487,N_26488,N_26490,N_26491,N_26492,N_26493,N_26498,N_26499,N_26500,N_26501,N_26503,N_26504,N_26505,N_26506,N_26508,N_26509,N_26511,N_26512,N_26513,N_26516,N_26517,N_26518,N_26520,N_26521,N_26522,N_26524,N_26526,N_26529,N_26532,N_26533,N_26535,N_26536,N_26537,N_26538,N_26539,N_26541,N_26542,N_26543,N_26545,N_26546,N_26548,N_26553,N_26555,N_26557,N_26558,N_26560,N_26562,N_26567,N_26569,N_26570,N_26572,N_26573,N_26576,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26603,N_26604,N_26605,N_26606,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26622,N_26624,N_26625,N_26628,N_26629,N_26630,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26641,N_26642,N_26643,N_26645,N_26646,N_26647,N_26648,N_26649,N_26651,N_26653,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26664,N_26665,N_26666,N_26667,N_26669,N_26670,N_26671,N_26673,N_26674,N_26676,N_26678,N_26680,N_26681,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26695,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26704,N_26706,N_26707,N_26709,N_26710,N_26711,N_26713,N_26714,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26733,N_26734,N_26735,N_26736,N_26738,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26748,N_26749,N_26750,N_26751,N_26753,N_26757,N_26759,N_26760,N_26761,N_26763,N_26764,N_26765,N_26766,N_26768,N_26769,N_26770,N_26772,N_26776,N_26779,N_26780,N_26781,N_26782,N_26784,N_26785,N_26786,N_26788,N_26791,N_26794,N_26795,N_26796,N_26797,N_26800,N_26801,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26824,N_26825,N_26826,N_26828,N_26829,N_26830,N_26831,N_26834,N_26836,N_26837,N_26838,N_26839,N_26841,N_26843,N_26845,N_26846,N_26847,N_26848,N_26851,N_26852,N_26853,N_26854,N_26856,N_26857,N_26858,N_26860,N_26861,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26877,N_26879,N_26880,N_26881,N_26882,N_26883,N_26885,N_26890,N_26891,N_26894,N_26897,N_26898,N_26899,N_26900,N_26902,N_26903,N_26904,N_26910,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26920,N_26921,N_26924,N_26925,N_26927,N_26928,N_26930,N_26931,N_26932,N_26933,N_26934,N_26936,N_26938,N_26939,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26955,N_26956,N_26958,N_26960,N_26961,N_26962,N_26965,N_26966,N_26967,N_26968,N_26971,N_26974,N_26975,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26985,N_26986,N_26987,N_26990,N_26991,N_26992,N_26996,N_26997,N_26998,N_26999,N_27000,N_27003,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27021,N_27022,N_27023,N_27024,N_27026,N_27029,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27048,N_27049,N_27050,N_27051,N_27052,N_27055,N_27056,N_27057,N_27060,N_27062,N_27063,N_27064,N_27066,N_27067,N_27069,N_27071,N_27072,N_27073,N_27074,N_27076,N_27078,N_27079,N_27080,N_27082,N_27083,N_27086,N_27087,N_27088,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27097,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27118,N_27119,N_27120,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27130,N_27132,N_27133,N_27134,N_27135,N_27136,N_27138,N_27140,N_27141,N_27145,N_27146,N_27147,N_27149,N_27151,N_27153,N_27156,N_27157,N_27158,N_27160,N_27162,N_27165,N_27167,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27177,N_27178,N_27180,N_27181,N_27182,N_27183,N_27185,N_27186,N_27187,N_27189,N_27190,N_27193,N_27194,N_27196,N_27199,N_27200,N_27201,N_27203,N_27204,N_27205,N_27207,N_27209,N_27210,N_27211,N_27212,N_27213,N_27215,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27224,N_27225,N_27226,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27236,N_27237,N_27243,N_27245,N_27246,N_27247,N_27248,N_27250,N_27252,N_27254,N_27255,N_27256,N_27257,N_27259,N_27260,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27272,N_27275,N_27277,N_27278,N_27280,N_27281,N_27283,N_27284,N_27285,N_27287,N_27288,N_27291,N_27292,N_27293,N_27295,N_27298,N_27299,N_27300,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27310,N_27312,N_27314,N_27315,N_27318,N_27320,N_27321,N_27322,N_27323,N_27325,N_27326,N_27328,N_27329,N_27331,N_27332,N_27333,N_27335,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27346,N_27347,N_27350,N_27351,N_27353,N_27355,N_27357,N_27359,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27368,N_27370,N_27372,N_27373,N_27375,N_27376,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27398,N_27402,N_27403,N_27405,N_27406,N_27408,N_27409,N_27413,N_27414,N_27415,N_27416,N_27419,N_27421,N_27422,N_27423,N_27425,N_27426,N_27427,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27438,N_27440,N_27443,N_27444,N_27447,N_27448,N_27449,N_27452,N_27453,N_27454,N_27455,N_27456,N_27458,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27474,N_27475,N_27476,N_27478,N_27480,N_27483,N_27484,N_27486,N_27487,N_27488,N_27489,N_27494,N_27495,N_27496,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27514,N_27517,N_27518,N_27519,N_27520,N_27521,N_27525,N_27526,N_27527,N_27528,N_27529,N_27531,N_27533,N_27534,N_27535,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27545,N_27546,N_27547,N_27549,N_27553,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27591,N_27592,N_27593,N_27594,N_27596,N_27597,N_27599,N_27600,N_27601,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27612,N_27613,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27631,N_27632,N_27633,N_27634,N_27637,N_27638,N_27639,N_27640,N_27642,N_27643,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27657,N_27658,N_27659,N_27660,N_27661,N_27663,N_27664,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27685,N_27686,N_27687,N_27691,N_27692,N_27693,N_27697,N_27700,N_27701,N_27702,N_27703,N_27704,N_27706,N_27708,N_27710,N_27711,N_27713,N_27714,N_27716,N_27718,N_27719,N_27720,N_27721,N_27722,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27735,N_27736,N_27737,N_27739,N_27740,N_27741,N_27742,N_27745,N_27747,N_27748,N_27749,N_27752,N_27753,N_27754,N_27759,N_27760,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27779,N_27781,N_27782,N_27785,N_27786,N_27788,N_27792,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27802,N_27803,N_27804,N_27806,N_27807,N_27809,N_27812,N_27814,N_27815,N_27816,N_27818,N_27820,N_27821,N_27824,N_27826,N_27827,N_27828,N_27830,N_27831,N_27832,N_27833,N_27835,N_27836,N_27837,N_27838,N_27839,N_27841,N_27842,N_27843,N_27845,N_27846,N_27847,N_27850,N_27851,N_27852,N_27853,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27867,N_27869,N_27871,N_27872,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27882,N_27883,N_27885,N_27889,N_27890,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27901,N_27902,N_27903,N_27905,N_27906,N_27907,N_27909,N_27910,N_27911,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27951,N_27952,N_27954,N_27955,N_27957,N_27959,N_27960,N_27961,N_27962,N_27964,N_27966,N_27969,N_27970,N_27972,N_27973,N_27974,N_27975,N_27977,N_27978,N_27979,N_27980,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27991,N_27992,N_27993,N_27994,N_27996,N_27998,N_27999,N_28000,N_28003,N_28004,N_28007,N_28009,N_28010,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28020,N_28021,N_28022,N_28023,N_28024,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28036,N_28037,N_28038,N_28039,N_28040,N_28042,N_28043,N_28044,N_28045,N_28046,N_28048,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28059,N_28060,N_28061,N_28062,N_28064,N_28067,N_28070,N_28071,N_28072,N_28075,N_28076,N_28078,N_28080,N_28081,N_28083,N_28084,N_28086,N_28087,N_28088,N_28090,N_28091,N_28093,N_28094,N_28095,N_28096,N_28100,N_28101,N_28102,N_28105,N_28106,N_28107,N_28110,N_28111,N_28112,N_28113,N_28115,N_28116,N_28117,N_28118,N_28120,N_28121,N_28123,N_28125,N_28126,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28143,N_28144,N_28149,N_28150,N_28152,N_28153,N_28154,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28171,N_28172,N_28173,N_28175,N_28176,N_28178,N_28179,N_28180,N_28181,N_28182,N_28184,N_28187,N_28188,N_28189,N_28190,N_28191,N_28193,N_28194,N_28196,N_28197,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28213,N_28214,N_28215,N_28216,N_28222,N_28224,N_28225,N_28226,N_28227,N_28229,N_28230,N_28232,N_28233,N_28234,N_28235,N_28238,N_28239,N_28240,N_28241,N_28242,N_28245,N_28247,N_28249,N_28251,N_28252,N_28253,N_28255,N_28256,N_28257,N_28258,N_28261,N_28263,N_28265,N_28266,N_28267,N_28268,N_28269,N_28271,N_28272,N_28273,N_28275,N_28276,N_28277,N_28278,N_28280,N_28282,N_28283,N_28284,N_28285,N_28291,N_28292,N_28293,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28306,N_28307,N_28308,N_28310,N_28314,N_28316,N_28317,N_28319,N_28320,N_28322,N_28324,N_28325,N_28327,N_28328,N_28330,N_28332,N_28333,N_28334,N_28335,N_28336,N_28338,N_28340,N_28341,N_28342,N_28343,N_28344,N_28346,N_28347,N_28348,N_28349,N_28350,N_28355,N_28356,N_28357,N_28358,N_28359,N_28362,N_28364,N_28366,N_28367,N_28368,N_28369,N_28373,N_28375,N_28376,N_28377,N_28378,N_28379,N_28381,N_28383,N_28384,N_28386,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28397,N_28398,N_28399,N_28400,N_28402,N_28403,N_28405,N_28406,N_28408,N_28409,N_28410,N_28411,N_28412,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28427,N_28429,N_28431,N_28432,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28461,N_28462,N_28463,N_28464,N_28467,N_28468,N_28470,N_28471,N_28474,N_28476,N_28477,N_28479,N_28482,N_28483,N_28485,N_28488,N_28490,N_28491,N_28492,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28502,N_28503,N_28504,N_28506,N_28507,N_28508,N_28509,N_28510,N_28512,N_28514,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28533,N_28534,N_28537,N_28538,N_28539,N_28540,N_28541,N_28543,N_28545,N_28546,N_28549,N_28551,N_28552,N_28554,N_28555,N_28556,N_28560,N_28561,N_28562,N_28564,N_28565,N_28566,N_28567,N_28568,N_28570,N_28572,N_28573,N_28574,N_28575,N_28577,N_28578,N_28580,N_28581,N_28583,N_28584,N_28585,N_28587,N_28588,N_28589,N_28590,N_28591,N_28593,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28605,N_28606,N_28607,N_28608,N_28611,N_28613,N_28614,N_28615,N_28618,N_28619,N_28626,N_28627,N_28629,N_28630,N_28632,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28652,N_28655,N_28656,N_28657,N_28659,N_28660,N_28661,N_28663,N_28665,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28674,N_28676,N_28679,N_28680,N_28681,N_28682,N_28684,N_28686,N_28687,N_28688,N_28690,N_28691,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28704,N_28705,N_28706,N_28708,N_28709,N_28710,N_28712,N_28714,N_28715,N_28717,N_28719,N_28720,N_28721,N_28722,N_28723,N_28725,N_28726,N_28727,N_28728,N_28731,N_28732,N_28733,N_28734,N_28735,N_28737,N_28738,N_28739,N_28740,N_28741,N_28743,N_28744,N_28747,N_28748,N_28749,N_28751,N_28753,N_28754,N_28755,N_28756,N_28757,N_28759,N_28760,N_28761,N_28762,N_28763,N_28766,N_28767,N_28768,N_28770,N_28771,N_28773,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28796,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28814,N_28816,N_28819,N_28821,N_28824,N_28825,N_28827,N_28828,N_28829,N_28830,N_28831,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28848,N_28849,N_28851,N_28852,N_28854,N_28855,N_28857,N_28858,N_28859,N_28862,N_28863,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28873,N_28874,N_28875,N_28876,N_28878,N_28879,N_28882,N_28883,N_28885,N_28887,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28915,N_28916,N_28918,N_28919,N_28920,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28938,N_28939,N_28940,N_28943,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28953,N_28954,N_28955,N_28956,N_28958,N_28960,N_28963,N_28965,N_28966,N_28967,N_28969,N_28970,N_28972,N_28973,N_28974,N_28975,N_28976,N_28978,N_28982,N_28984,N_28985,N_28986,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28997,N_28998,N_28999,N_29000,N_29002,N_29003,N_29006,N_29007,N_29009,N_29010,N_29011,N_29012,N_29014,N_29015,N_29016,N_29018,N_29023,N_29024,N_29026,N_29028,N_29029,N_29030,N_29031,N_29033,N_29035,N_29037,N_29038,N_29040,N_29041,N_29043,N_29045,N_29047,N_29048,N_29049,N_29051,N_29052,N_29053,N_29054,N_29056,N_29057,N_29059,N_29060,N_29062,N_29063,N_29066,N_29069,N_29070,N_29071,N_29073,N_29074,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29084,N_29085,N_29086,N_29087,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29098,N_29099,N_29102,N_29103,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29112,N_29114,N_29115,N_29116,N_29118,N_29119,N_29121,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29131,N_29134,N_29135,N_29136,N_29138,N_29143,N_29144,N_29145,N_29146,N_29147,N_29149,N_29152,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29174,N_29175,N_29176,N_29177,N_29178,N_29180,N_29183,N_29184,N_29185,N_29186,N_29188,N_29190,N_29191,N_29193,N_29194,N_29196,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29211,N_29212,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29228,N_29229,N_29230,N_29231,N_29233,N_29235,N_29236,N_29238,N_29239,N_29240,N_29243,N_29244,N_29245,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29256,N_29257,N_29258,N_29260,N_29262,N_29263,N_29264,N_29266,N_29269,N_29270,N_29272,N_29273,N_29275,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29285,N_29286,N_29287,N_29288,N_29290,N_29291,N_29292,N_29293,N_29294,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29305,N_29307,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29321,N_29323,N_29324,N_29326,N_29327,N_29328,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29340,N_29341,N_29343,N_29345,N_29347,N_29349,N_29350,N_29351,N_29352,N_29353,N_29355,N_29357,N_29358,N_29359,N_29360,N_29362,N_29364,N_29366,N_29367,N_29369,N_29370,N_29371,N_29372,N_29373,N_29375,N_29376,N_29377,N_29378,N_29382,N_29384,N_29385,N_29387,N_29388,N_29389,N_29390,N_29391,N_29393,N_29394,N_29396,N_29397,N_29399,N_29400,N_29401,N_29403,N_29404,N_29405,N_29406,N_29410,N_29411,N_29412,N_29413,N_29418,N_29419,N_29420,N_29421,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29432,N_29434,N_29436,N_29438,N_29439,N_29440,N_29442,N_29443,N_29444,N_29445,N_29448,N_29449,N_29450,N_29451,N_29453,N_29454,N_29455,N_29457,N_29458,N_29459,N_29460,N_29462,N_29464,N_29465,N_29466,N_29467,N_29469,N_29470,N_29471,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29485,N_29487,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29508,N_29510,N_29511,N_29513,N_29514,N_29516,N_29518,N_29519,N_29521,N_29522,N_29526,N_29528,N_29529,N_29532,N_29533,N_29536,N_29537,N_29539,N_29542,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29552,N_29553,N_29554,N_29555,N_29558,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29568,N_29570,N_29571,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29588,N_29589,N_29591,N_29592,N_29593,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29612,N_29613,N_29615,N_29616,N_29617,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29633,N_29634,N_29635,N_29636,N_29637,N_29639,N_29640,N_29641,N_29645,N_29646,N_29647,N_29650,N_29651,N_29654,N_29655,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29666,N_29667,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29685,N_29686,N_29689,N_29690,N_29691,N_29693,N_29695,N_29696,N_29697,N_29698,N_29700,N_29702,N_29703,N_29704,N_29706,N_29707,N_29712,N_29713,N_29714,N_29715,N_29716,N_29719,N_29721,N_29722,N_29725,N_29727,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29736,N_29737,N_29739,N_29742,N_29743,N_29744,N_29745,N_29747,N_29748,N_29750,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29766,N_29767,N_29768,N_29769,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29780,N_29781,N_29783,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29803,N_29805,N_29806,N_29807,N_29808,N_29810,N_29811,N_29820,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29840,N_29843,N_29844,N_29845,N_29847,N_29848,N_29849,N_29851,N_29852,N_29853,N_29856,N_29857,N_29858,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29872,N_29873,N_29874,N_29875,N_29877,N_29878,N_29879,N_29883,N_29885,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29898,N_29900,N_29901,N_29903,N_29904,N_29907,N_29909,N_29910,N_29912,N_29913,N_29920,N_29924,N_29930,N_29932,N_29933,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29945,N_29946,N_29947,N_29948,N_29950,N_29952,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29962,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998;
nand U0 (N_0,In_1514,In_1119);
xnor U1 (N_1,In_1229,In_1991);
nand U2 (N_2,In_1547,In_546);
and U3 (N_3,In_2287,In_1426);
nor U4 (N_4,In_791,In_1651);
or U5 (N_5,In_805,In_621);
or U6 (N_6,In_1139,In_877);
nor U7 (N_7,In_211,In_1901);
nand U8 (N_8,In_258,In_2965);
nor U9 (N_9,In_2262,In_39);
or U10 (N_10,In_1491,In_1376);
nor U11 (N_11,In_1503,In_583);
and U12 (N_12,In_229,In_2486);
nand U13 (N_13,In_1753,In_2442);
xor U14 (N_14,In_861,In_1921);
or U15 (N_15,In_1087,In_2997);
nor U16 (N_16,In_1019,In_1409);
nor U17 (N_17,In_2377,In_2110);
or U18 (N_18,In_2653,In_1294);
or U19 (N_19,In_112,In_578);
xor U20 (N_20,In_2853,In_2117);
nand U21 (N_21,In_1973,In_1007);
nand U22 (N_22,In_1918,In_1322);
nor U23 (N_23,In_858,In_1723);
nor U24 (N_24,In_1355,In_306);
or U25 (N_25,In_427,In_2251);
nor U26 (N_26,In_301,In_167);
xnor U27 (N_27,In_2699,In_2522);
nor U28 (N_28,In_1300,In_942);
nor U29 (N_29,In_815,In_2984);
and U30 (N_30,In_976,In_1198);
xnor U31 (N_31,In_2602,In_1914);
or U32 (N_32,In_788,In_2747);
xor U33 (N_33,In_1864,In_1689);
xnor U34 (N_34,In_909,In_1564);
or U35 (N_35,In_2426,In_2875);
and U36 (N_36,In_2375,In_1774);
nor U37 (N_37,In_1989,In_2986);
or U38 (N_38,In_2448,In_2970);
nand U39 (N_39,In_1776,In_2423);
and U40 (N_40,In_2983,In_263);
nor U41 (N_41,In_2750,In_1047);
nand U42 (N_42,In_118,In_224);
or U43 (N_43,In_2160,In_2381);
nand U44 (N_44,In_73,In_2643);
nor U45 (N_45,In_1385,In_448);
or U46 (N_46,In_987,In_2506);
or U47 (N_47,In_42,In_2547);
nand U48 (N_48,In_1907,In_1266);
nand U49 (N_49,In_2717,In_2291);
or U50 (N_50,In_985,In_1246);
and U51 (N_51,In_2848,In_2576);
and U52 (N_52,In_1234,In_1667);
xnor U53 (N_53,In_558,In_998);
nand U54 (N_54,In_1482,In_2277);
and U55 (N_55,In_144,In_435);
nor U56 (N_56,In_2850,In_626);
or U57 (N_57,In_924,In_62);
nand U58 (N_58,In_447,In_1185);
xnor U59 (N_59,In_2139,In_2860);
or U60 (N_60,In_2464,In_2684);
xor U61 (N_61,In_1625,In_1810);
nor U62 (N_62,In_2271,In_1736);
xor U63 (N_63,In_2795,In_2258);
nand U64 (N_64,In_430,In_542);
and U65 (N_65,In_504,In_659);
nor U66 (N_66,In_2912,In_2134);
or U67 (N_67,In_291,In_2951);
or U68 (N_68,In_947,In_613);
nor U69 (N_69,In_531,In_1944);
xor U70 (N_70,In_1572,In_309);
xor U71 (N_71,In_2922,In_846);
nand U72 (N_72,In_2072,In_2254);
and U73 (N_73,In_276,In_1100);
nor U74 (N_74,In_2786,In_2085);
xnor U75 (N_75,In_378,In_1039);
and U76 (N_76,In_2525,In_2639);
nor U77 (N_77,In_1211,In_1730);
nor U78 (N_78,In_168,In_1197);
xor U79 (N_79,In_191,In_783);
xor U80 (N_80,In_714,In_237);
nand U81 (N_81,In_1035,In_1721);
nor U82 (N_82,In_1069,In_1452);
or U83 (N_83,In_1546,In_2482);
and U84 (N_84,In_2540,In_2940);
xor U85 (N_85,In_687,In_2297);
xor U86 (N_86,In_1854,In_1113);
or U87 (N_87,In_1421,In_2052);
and U88 (N_88,In_2490,In_2273);
nor U89 (N_89,In_33,In_763);
nand U90 (N_90,In_1791,In_2167);
nor U91 (N_91,In_2820,In_1799);
and U92 (N_92,In_753,In_179);
xnor U93 (N_93,In_460,In_2348);
nor U94 (N_94,In_875,In_131);
or U95 (N_95,In_1362,In_2116);
or U96 (N_96,In_2059,In_2956);
or U97 (N_97,In_2510,In_2255);
nand U98 (N_98,In_2462,In_1390);
nor U99 (N_99,In_590,In_629);
xor U100 (N_100,In_2011,In_2051);
xnor U101 (N_101,In_1570,In_1559);
nor U102 (N_102,In_1557,In_601);
nand U103 (N_103,In_834,In_2946);
and U104 (N_104,In_2321,In_215);
and U105 (N_105,In_2125,In_2213);
xnor U106 (N_106,In_2972,In_2228);
nor U107 (N_107,In_2298,In_2189);
and U108 (N_108,In_1057,In_640);
xor U109 (N_109,In_157,In_2048);
xor U110 (N_110,In_103,In_1273);
or U111 (N_111,In_1207,In_1013);
nand U112 (N_112,In_2020,In_1126);
xor U113 (N_113,In_588,In_884);
nor U114 (N_114,In_287,In_737);
nor U115 (N_115,In_1205,In_2872);
nand U116 (N_116,In_1397,In_1088);
and U117 (N_117,In_598,In_2234);
xnor U118 (N_118,In_2264,In_953);
and U119 (N_119,In_1440,In_1147);
or U120 (N_120,In_1360,In_434);
and U121 (N_121,In_487,In_2557);
nand U122 (N_122,In_1208,In_64);
or U123 (N_123,In_1484,In_1314);
xor U124 (N_124,In_2887,In_1489);
or U125 (N_125,In_1654,In_1321);
or U126 (N_126,In_2917,In_1908);
nand U127 (N_127,In_307,In_1369);
and U128 (N_128,In_2526,In_226);
xnor U129 (N_129,In_381,In_2190);
xor U130 (N_130,In_717,In_1955);
and U131 (N_131,In_2199,In_397);
and U132 (N_132,In_1371,In_1105);
nand U133 (N_133,In_682,In_2045);
or U134 (N_134,In_1781,In_392);
nor U135 (N_135,In_1889,In_1716);
nand U136 (N_136,In_2855,In_2644);
nor U137 (N_137,In_555,In_244);
nor U138 (N_138,In_1109,In_1856);
and U139 (N_139,In_894,In_2885);
xnor U140 (N_140,In_2065,In_120);
nor U141 (N_141,In_2027,In_278);
nor U142 (N_142,In_2220,In_1662);
and U143 (N_143,In_320,In_1943);
xor U144 (N_144,In_384,In_1021);
xor U145 (N_145,In_2401,In_599);
nand U146 (N_146,In_711,In_1875);
and U147 (N_147,In_2186,In_2935);
nor U148 (N_148,In_2575,In_2837);
nand U149 (N_149,In_907,In_657);
nand U150 (N_150,In_926,In_1264);
or U151 (N_151,In_472,In_1950);
nand U152 (N_152,In_2856,In_614);
or U153 (N_153,In_1215,In_2934);
nand U154 (N_154,In_165,In_428);
nor U155 (N_155,In_2142,In_344);
or U156 (N_156,In_2242,In_477);
nor U157 (N_157,In_859,In_1978);
nor U158 (N_158,In_198,In_2500);
or U159 (N_159,In_256,In_1183);
xnor U160 (N_160,In_416,In_1518);
or U161 (N_161,In_2570,In_1699);
nand U162 (N_162,In_299,In_740);
nor U163 (N_163,In_194,In_2604);
nor U164 (N_164,In_2392,In_535);
xor U165 (N_165,In_1836,In_968);
nand U166 (N_166,In_718,In_2752);
nand U167 (N_167,In_2225,In_1114);
nand U168 (N_168,In_2589,In_681);
nand U169 (N_169,In_756,In_2936);
nor U170 (N_170,In_2324,In_1777);
and U171 (N_171,In_2122,In_1089);
and U172 (N_172,In_2430,In_510);
nor U173 (N_173,In_525,In_133);
xor U174 (N_174,In_2404,In_2531);
nand U175 (N_175,In_2610,In_1529);
nor U176 (N_176,In_1276,In_2283);
nor U177 (N_177,In_2474,In_679);
xor U178 (N_178,In_691,In_1511);
nor U179 (N_179,In_1399,In_620);
xor U180 (N_180,In_648,In_764);
xor U181 (N_181,In_349,In_1417);
nand U182 (N_182,In_917,In_1408);
nand U183 (N_183,In_1775,In_2006);
xor U184 (N_184,In_2802,In_8);
nand U185 (N_185,In_2074,In_1922);
nand U186 (N_186,In_914,In_1590);
nand U187 (N_187,In_1841,In_650);
nor U188 (N_188,In_1381,In_2996);
xor U189 (N_189,In_1219,In_2976);
nor U190 (N_190,In_656,In_409);
nor U191 (N_191,In_2230,In_2660);
xnor U192 (N_192,In_994,In_1182);
or U193 (N_193,In_1186,In_2680);
nand U194 (N_194,In_109,In_1439);
xor U195 (N_195,In_2374,In_1363);
nand U196 (N_196,In_45,In_160);
xnor U197 (N_197,In_2720,In_1884);
nand U198 (N_198,In_1940,In_2580);
nor U199 (N_199,In_592,In_1647);
xnor U200 (N_200,In_63,In_2345);
nand U201 (N_201,In_2094,In_2200);
nor U202 (N_202,In_537,In_2642);
xnor U203 (N_203,In_2670,In_2656);
or U204 (N_204,In_1562,In_1504);
nand U205 (N_205,In_2909,In_2154);
or U206 (N_206,In_853,In_28);
nand U207 (N_207,In_2330,In_2755);
nor U208 (N_208,In_530,In_1539);
nand U209 (N_209,In_483,In_2364);
nor U210 (N_210,In_2034,In_2807);
or U211 (N_211,In_1123,In_2729);
xnor U212 (N_212,In_334,In_2318);
and U213 (N_213,In_672,In_528);
nor U214 (N_214,In_1095,In_2708);
and U215 (N_215,In_1538,In_55);
nor U216 (N_216,In_943,In_1151);
and U217 (N_217,In_406,In_2621);
or U218 (N_218,In_2662,In_1458);
nor U219 (N_219,In_2967,In_2615);
nor U220 (N_220,In_1878,In_2465);
and U221 (N_221,In_2980,In_1118);
xnor U222 (N_222,In_1571,In_319);
or U223 (N_223,In_2443,In_91);
or U224 (N_224,In_390,In_628);
and U225 (N_225,In_1495,In_444);
nor U226 (N_226,In_1278,In_1610);
nand U227 (N_227,In_1804,In_1038);
or U228 (N_228,In_403,In_2767);
or U229 (N_229,In_2798,In_2455);
or U230 (N_230,In_1240,In_2647);
and U231 (N_231,In_1947,In_1949);
xnor U232 (N_232,In_2745,In_2892);
nand U233 (N_233,In_2864,In_1044);
nor U234 (N_234,In_2239,In_2947);
nor U235 (N_235,In_1096,In_16);
nor U236 (N_236,In_864,In_2961);
nand U237 (N_237,In_2873,In_2175);
xor U238 (N_238,In_1283,In_2520);
nand U239 (N_239,In_2565,In_2485);
or U240 (N_240,In_1618,In_354);
nor U241 (N_241,In_1206,In_2077);
nor U242 (N_242,In_2813,In_786);
nand U243 (N_243,In_2685,In_31);
and U244 (N_244,In_2757,In_2832);
or U245 (N_245,In_2379,In_841);
and U246 (N_246,In_2995,In_333);
nand U247 (N_247,In_1176,In_2247);
nor U248 (N_248,In_556,In_984);
and U249 (N_249,In_1823,In_2236);
nand U250 (N_250,In_485,In_832);
or U251 (N_251,In_2327,In_1137);
nor U252 (N_252,In_2418,In_2707);
and U253 (N_253,In_2666,In_1463);
nor U254 (N_254,In_1782,In_1257);
nand U255 (N_255,In_2484,In_2447);
nor U256 (N_256,In_1429,In_2834);
nand U257 (N_257,In_2742,In_1905);
and U258 (N_258,In_1432,In_1698);
or U259 (N_259,In_840,In_2756);
or U260 (N_260,In_56,In_1261);
or U261 (N_261,In_1814,In_275);
nor U262 (N_262,In_164,In_1772);
nand U263 (N_263,In_281,In_2126);
and U264 (N_264,In_895,In_716);
or U265 (N_265,In_1602,In_1064);
xnor U266 (N_266,In_1962,In_2775);
nor U267 (N_267,In_346,In_2928);
and U268 (N_268,In_2169,In_752);
or U269 (N_269,In_2545,In_443);
or U270 (N_270,In_499,In_2870);
and U271 (N_271,In_1419,In_1356);
nand U272 (N_272,In_1425,In_1926);
nor U273 (N_273,In_1838,In_1387);
or U274 (N_274,In_2269,In_413);
and U275 (N_275,In_2563,In_1595);
nor U276 (N_276,In_2607,In_342);
nand U277 (N_277,In_2638,In_1859);
and U278 (N_278,In_1085,In_2854);
nand U279 (N_279,In_1128,In_2672);
and U280 (N_280,In_1587,In_2257);
nor U281 (N_281,In_1980,In_410);
or U282 (N_282,In_101,In_2180);
or U283 (N_283,In_2050,In_990);
nand U284 (N_284,In_1826,In_2215);
or U285 (N_285,In_1427,In_660);
and U286 (N_286,In_65,In_1702);
nand U287 (N_287,In_2128,In_878);
and U288 (N_288,In_908,In_2926);
nand U289 (N_289,In_2688,In_902);
nor U290 (N_290,In_442,In_2876);
nand U291 (N_291,In_2583,In_273);
xor U292 (N_292,In_1820,In_105);
nand U293 (N_293,In_1325,In_111);
xnor U294 (N_294,In_1204,In_2552);
and U295 (N_295,In_1305,In_2036);
nand U296 (N_296,In_2212,In_200);
xor U297 (N_297,In_158,In_1338);
xnor U298 (N_298,In_1936,In_2938);
nor U299 (N_299,In_1402,In_2323);
and U300 (N_300,In_919,In_1701);
nor U301 (N_301,In_2655,In_844);
and U302 (N_302,In_2825,In_1522);
nand U303 (N_303,In_1500,In_84);
and U304 (N_304,In_89,In_50);
nor U305 (N_305,In_1401,In_2260);
xor U306 (N_306,In_954,In_1811);
or U307 (N_307,In_769,In_511);
or U308 (N_308,In_1135,In_1160);
nor U309 (N_309,In_95,In_2840);
nor U310 (N_310,In_2047,In_1302);
and U311 (N_311,In_295,In_1175);
nand U312 (N_312,In_1093,In_1307);
nand U313 (N_313,In_2715,In_2461);
or U314 (N_314,In_938,In_1184);
nand U315 (N_315,In_1014,In_5);
nand U316 (N_316,In_1284,In_1049);
nand U317 (N_317,In_773,In_2394);
and U318 (N_318,In_2746,In_2003);
xor U319 (N_319,In_2140,In_13);
or U320 (N_320,In_2793,In_731);
nand U321 (N_321,In_2070,In_1643);
and U322 (N_322,In_591,In_2356);
nor U323 (N_323,In_1188,In_549);
and U324 (N_324,In_2342,In_79);
nor U325 (N_325,In_1548,In_214);
nand U326 (N_326,In_2100,In_1468);
or U327 (N_327,In_1745,In_1833);
or U328 (N_328,In_2700,In_2410);
nand U329 (N_329,In_1200,In_609);
and U330 (N_330,In_494,In_1824);
or U331 (N_331,In_2705,In_122);
nand U332 (N_332,In_2818,In_2347);
nor U333 (N_333,In_813,In_205);
nand U334 (N_334,In_863,In_855);
xnor U335 (N_335,In_2411,In_280);
or U336 (N_336,In_514,In_389);
nand U337 (N_337,In_890,In_1343);
nand U338 (N_338,In_1853,In_2037);
nand U339 (N_339,In_2363,In_1703);
or U340 (N_340,In_2076,In_1247);
xor U341 (N_341,In_1451,In_1871);
nor U342 (N_342,In_1398,In_848);
xor U343 (N_343,In_776,In_2902);
or U344 (N_344,In_874,In_1022);
and U345 (N_345,In_2712,In_1976);
xnor U346 (N_346,In_1545,In_2451);
nor U347 (N_347,In_1683,In_75);
xor U348 (N_348,In_1645,In_187);
and U349 (N_349,In_1048,In_2982);
nor U350 (N_350,In_1011,In_2827);
xnor U351 (N_351,In_1964,In_2436);
or U352 (N_352,In_2509,In_2325);
nor U353 (N_353,In_166,In_1586);
or U354 (N_354,In_1675,In_1924);
xor U355 (N_355,In_2859,In_2454);
nand U356 (N_356,In_2626,In_358);
and U357 (N_357,In_2952,In_2916);
nor U358 (N_358,In_2337,In_870);
nor U359 (N_359,In_2222,In_2479);
xor U360 (N_360,In_595,In_2578);
nand U361 (N_361,In_977,In_305);
and U362 (N_362,In_2367,In_1852);
nand U363 (N_363,In_2343,In_2202);
and U364 (N_364,In_1560,In_1850);
nand U365 (N_365,In_1090,In_677);
or U366 (N_366,In_482,In_24);
or U367 (N_367,In_2237,In_666);
nor U368 (N_368,In_1469,In_931);
and U369 (N_369,In_2358,In_712);
and U370 (N_370,In_2906,In_170);
and U371 (N_371,In_429,In_1644);
and U372 (N_372,In_1435,In_2438);
nor U373 (N_373,In_1265,In_1711);
xor U374 (N_374,In_2868,In_2898);
or U375 (N_375,In_210,In_1285);
nand U376 (N_376,In_155,In_450);
and U377 (N_377,In_2599,In_387);
nand U378 (N_378,In_1187,In_2253);
or U379 (N_379,In_1552,In_2640);
nand U380 (N_380,In_2785,In_2921);
nor U381 (N_381,In_2810,In_1316);
xnor U382 (N_382,In_639,In_453);
and U383 (N_383,In_2311,In_2611);
or U384 (N_384,In_577,In_2651);
nor U385 (N_385,In_126,In_1301);
and U386 (N_386,In_1658,In_1475);
xor U387 (N_387,In_218,In_359);
nand U388 (N_388,In_2673,In_1712);
and U389 (N_389,In_2930,In_911);
xnor U390 (N_390,In_1462,In_2333);
and U391 (N_391,In_1555,In_2880);
nand U392 (N_392,In_982,In_1543);
or U393 (N_393,In_2749,In_1700);
xnor U394 (N_394,In_2409,In_1769);
or U395 (N_395,In_2130,In_1756);
xnor U396 (N_396,In_2722,In_634);
nor U397 (N_397,In_54,In_1152);
and U398 (N_398,In_2551,In_1512);
or U399 (N_399,In_2978,In_2267);
and U400 (N_400,In_2335,In_2194);
or U401 (N_401,In_2843,In_90);
nor U402 (N_402,In_1233,In_452);
and U403 (N_403,In_2014,In_996);
and U404 (N_404,In_2370,In_2429);
xnor U405 (N_405,In_2021,In_1874);
or U406 (N_406,In_270,In_582);
xnor U407 (N_407,In_2709,In_2847);
and U408 (N_408,In_6,In_1957);
or U409 (N_409,In_1173,In_2618);
and U410 (N_410,In_2698,In_2450);
and U411 (N_411,In_1212,In_1687);
and U412 (N_412,In_1953,In_701);
xor U413 (N_413,In_2731,In_2592);
xnor U414 (N_414,In_208,In_1194);
nor U415 (N_415,In_2549,In_329);
xnor U416 (N_416,In_608,In_439);
and U417 (N_417,In_2559,In_1330);
nor U418 (N_418,In_2596,In_322);
xnor U419 (N_419,In_847,In_2227);
or U420 (N_420,In_67,In_1816);
and U421 (N_421,In_469,In_2595);
nor U422 (N_422,In_1834,In_2999);
nor U423 (N_423,In_1225,In_1765);
nor U424 (N_424,In_2693,In_1568);
or U425 (N_425,In_1840,In_808);
nor U426 (N_426,In_825,In_1635);
nand U427 (N_427,In_2605,In_751);
xnor U428 (N_428,In_2679,In_1352);
nand U429 (N_429,In_554,In_1713);
nand U430 (N_430,In_2893,In_1785);
xnor U431 (N_431,In_552,In_513);
nand U432 (N_432,In_259,In_1773);
nand U433 (N_433,In_419,In_106);
and U434 (N_434,In_180,In_1849);
nor U435 (N_435,In_2771,In_2514);
or U436 (N_436,In_147,In_1719);
xor U437 (N_437,In_2470,In_1665);
and U438 (N_438,In_2453,In_2900);
nor U439 (N_439,In_1164,In_1954);
and U440 (N_440,In_476,In_2044);
nor U441 (N_441,In_850,In_1997);
nor U442 (N_442,In_1830,In_705);
nor U443 (N_443,In_2519,In_454);
nor U444 (N_444,In_1866,In_779);
nand U445 (N_445,In_2397,In_2606);
or U446 (N_446,In_2541,In_2765);
nand U447 (N_447,In_2445,In_2091);
xor U448 (N_448,In_1251,In_213);
and U449 (N_449,In_2838,In_2378);
and U450 (N_450,In_252,In_18);
or U451 (N_451,In_324,In_2718);
nor U452 (N_452,In_2248,In_221);
nor U453 (N_453,In_2646,In_314);
nor U454 (N_454,In_2294,In_2308);
nor U455 (N_455,In_1601,In_1697);
nor U456 (N_456,In_264,In_2663);
or U457 (N_457,In_683,In_26);
and U458 (N_458,In_1478,In_1910);
nand U459 (N_459,In_2261,In_741);
nor U460 (N_460,In_2622,In_2532);
or U461 (N_461,In_1574,In_283);
xor U462 (N_462,In_564,In_440);
nand U463 (N_463,In_2039,In_1430);
and U464 (N_464,In_1809,In_1904);
nor U465 (N_465,In_293,In_1592);
or U466 (N_466,In_1083,In_2152);
nor U467 (N_467,In_2413,In_644);
nor U468 (N_468,In_665,In_1970);
nand U469 (N_469,In_2508,In_2654);
or U470 (N_470,In_532,In_637);
xnor U471 (N_471,In_2488,In_647);
and U472 (N_472,In_449,In_29);
xor U473 (N_473,In_612,In_915);
and U474 (N_474,In_1827,In_780);
xor U475 (N_475,In_1348,In_2915);
xnor U476 (N_476,In_2881,In_353);
and U477 (N_477,In_2304,In_2503);
nor U478 (N_478,In_474,In_1112);
or U479 (N_479,In_2371,In_2328);
nand U480 (N_480,In_1082,In_1839);
xor U481 (N_481,In_1023,In_1192);
nor U482 (N_482,In_1053,In_2341);
and U483 (N_483,In_2962,In_2950);
and U484 (N_484,In_2010,In_1900);
and U485 (N_485,In_2231,In_2690);
or U486 (N_486,In_2704,In_1120);
or U487 (N_487,In_1883,In_2533);
nand U488 (N_488,In_2295,In_1043);
nand U489 (N_489,In_1920,In_1259);
or U490 (N_490,In_395,In_14);
and U491 (N_491,In_765,In_1414);
or U492 (N_492,In_1741,In_1752);
and U493 (N_493,In_1310,In_506);
nand U494 (N_494,In_851,In_2603);
and U495 (N_495,In_1861,In_1735);
and U496 (N_496,In_117,In_1540);
and U497 (N_497,In_394,In_2188);
or U498 (N_498,In_2161,In_518);
and U499 (N_499,In_1797,In_2351);
and U500 (N_500,In_1528,In_2046);
or U501 (N_501,In_2209,In_1664);
xor U502 (N_502,In_1056,In_725);
xnor U503 (N_503,In_2518,In_1030);
nand U504 (N_504,In_527,In_761);
or U505 (N_505,In_1818,In_573);
nand U506 (N_506,In_2732,In_1648);
xor U507 (N_507,In_2092,In_979);
and U508 (N_508,In_2082,In_1382);
nor U509 (N_509,In_1018,In_836);
xor U510 (N_510,In_2368,In_2831);
nand U511 (N_511,In_1933,In_1174);
nor U512 (N_512,In_2960,In_2015);
nand U513 (N_513,In_2290,In_536);
or U514 (N_514,In_99,In_2049);
xnor U515 (N_515,In_1923,In_2975);
nor U516 (N_516,In_1631,In_2990);
and U517 (N_517,In_2387,In_2030);
xnor U518 (N_518,In_680,In_2733);
and U519 (N_519,In_2927,In_2025);
or U520 (N_520,In_2417,In_2521);
xor U521 (N_521,In_922,In_662);
nand U522 (N_522,In_2738,In_1127);
or U523 (N_523,In_557,In_978);
or U524 (N_524,In_1705,In_2512);
or U525 (N_525,In_1029,In_2659);
and U526 (N_526,In_1274,In_104);
and U527 (N_527,In_2925,In_219);
xor U528 (N_528,In_336,In_1894);
nor U529 (N_529,In_2084,In_2883);
xnor U530 (N_530,In_1802,In_2103);
xnor U531 (N_531,In_604,In_1190);
xor U532 (N_532,In_617,In_367);
nor U533 (N_533,In_363,In_747);
nor U534 (N_534,In_945,In_2405);
xnor U535 (N_535,In_1391,In_2060);
and U536 (N_536,In_1146,In_829);
xor U537 (N_537,In_2494,In_2772);
nor U538 (N_538,In_1829,In_2625);
and U539 (N_539,In_1107,In_420);
xnor U540 (N_540,In_2195,In_1383);
nand U541 (N_541,In_1124,In_2104);
nor U542 (N_542,In_1649,In_197);
or U543 (N_543,In_2740,In_606);
and U544 (N_544,In_94,In_1692);
and U545 (N_545,In_2944,In_227);
and U546 (N_546,In_1751,In_2406);
and U547 (N_547,In_702,In_2609);
and U548 (N_548,In_951,In_1319);
nor U549 (N_549,In_1860,In_1966);
nand U550 (N_550,In_1457,In_2493);
or U551 (N_551,In_2109,In_937);
nor U552 (N_552,In_1315,In_2256);
and U553 (N_553,In_311,In_44);
xor U554 (N_554,In_432,In_901);
xor U555 (N_555,In_2937,In_1690);
or U556 (N_556,In_2312,In_889);
nand U557 (N_557,In_1282,In_1579);
xnor U558 (N_558,In_940,In_567);
nand U559 (N_559,In_383,In_941);
nor U560 (N_560,In_1862,In_2744);
xnor U561 (N_561,In_267,In_1652);
nand U562 (N_562,In_548,In_2858);
nand U563 (N_563,In_337,In_1454);
xor U564 (N_564,In_248,In_1759);
nand U565 (N_565,In_2851,In_2383);
nor U566 (N_566,In_17,In_1523);
and U567 (N_567,In_950,In_1031);
nor U568 (N_568,In_326,In_2682);
xnor U569 (N_569,In_4,In_2388);
nor U570 (N_570,In_300,In_1569);
or U571 (N_571,In_1524,In_2163);
and U572 (N_572,In_2400,In_1170);
nor U573 (N_573,In_619,In_2539);
nor U574 (N_574,In_642,In_1122);
xnor U575 (N_575,In_587,In_1906);
nor U576 (N_576,In_1235,In_2469);
xnor U577 (N_577,In_623,In_1242);
nor U578 (N_578,In_407,In_2302);
nor U579 (N_579,In_2845,In_2761);
nor U580 (N_580,In_2546,In_1106);
or U581 (N_581,In_399,In_192);
nor U582 (N_582,In_1263,In_1413);
xnor U583 (N_583,In_2939,In_674);
or U584 (N_584,In_470,In_2491);
nor U585 (N_585,In_1004,In_492);
or U586 (N_586,In_1734,In_876);
and U587 (N_587,In_1930,In_2382);
or U588 (N_588,In_2040,In_988);
or U589 (N_589,In_2101,In_1680);
or U590 (N_590,In_2790,In_1236);
nand U591 (N_591,In_107,In_2507);
and U592 (N_592,In_97,In_1344);
nand U593 (N_593,In_1999,In_2309);
xnor U594 (N_594,In_653,In_2770);
and U595 (N_595,In_562,In_586);
nor U596 (N_596,In_1868,In_920);
or U597 (N_597,In_486,In_2460);
nor U598 (N_598,In_1101,In_1727);
xnor U599 (N_599,In_1311,In_722);
xnor U600 (N_600,In_2111,In_975);
xnor U601 (N_601,In_2788,In_1159);
xnor U602 (N_602,In_733,In_2637);
nand U603 (N_603,In_1213,In_2584);
and U604 (N_604,In_2544,In_2805);
and U605 (N_605,In_2762,In_1858);
nor U606 (N_606,In_411,In_2568);
nand U607 (N_607,In_739,In_2017);
xnor U608 (N_608,In_1679,In_1230);
or U609 (N_609,In_114,In_2706);
or U610 (N_610,In_1060,In_957);
nand U611 (N_611,In_129,In_930);
or U612 (N_612,In_2734,In_775);
or U613 (N_613,In_1244,In_445);
or U614 (N_614,In_1193,In_2992);
xor U615 (N_615,In_1593,In_76);
nor U616 (N_616,In_1611,In_1453);
xnor U617 (N_617,In_2778,In_142);
nand U618 (N_618,In_1982,In_2696);
nand U619 (N_619,In_1725,In_421);
nand U620 (N_620,In_243,In_1405);
or U621 (N_621,In_508,In_607);
xnor U622 (N_622,In_770,In_139);
xor U623 (N_623,In_2701,In_1676);
nand U624 (N_624,In_997,In_2779);
or U625 (N_625,In_589,In_2723);
nand U626 (N_626,In_2069,In_1481);
nand U627 (N_627,In_41,In_1554);
nand U628 (N_628,In_1945,In_966);
nor U629 (N_629,In_1619,In_1133);
nand U630 (N_630,In_159,In_1917);
xor U631 (N_631,In_576,In_2487);
and U632 (N_632,In_819,In_480);
and U633 (N_633,In_302,In_921);
nand U634 (N_634,In_1641,In_1140);
xnor U635 (N_635,In_2288,In_93);
or U636 (N_636,In_1486,In_2424);
nand U637 (N_637,In_2086,In_708);
nor U638 (N_638,In_318,In_1749);
nand U639 (N_639,In_366,In_2613);
xnor U640 (N_640,In_2739,In_2808);
xor U641 (N_641,In_2434,In_2619);
nor U642 (N_642,In_1415,In_1821);
nor U643 (N_643,In_1354,In_1393);
or U644 (N_644,In_1070,In_1846);
and U645 (N_645,In_2991,In_490);
nor U646 (N_646,In_2329,In_2459);
nand U647 (N_647,In_1708,In_478);
xor U648 (N_648,In_1306,In_2768);
and U649 (N_649,In_343,In_539);
xnor U650 (N_650,In_1162,In_1012);
and U651 (N_651,In_1981,In_1042);
and U652 (N_652,In_35,In_1386);
xor U653 (N_653,In_1267,In_1795);
nand U654 (N_654,In_1886,In_575);
xor U655 (N_655,In_935,In_1279);
nand U656 (N_656,In_2674,In_1660);
xnor U657 (N_657,In_962,In_1709);
xnor U658 (N_658,In_1498,In_209);
xor U659 (N_659,In_1627,In_2617);
xnor U660 (N_660,In_1580,In_675);
or U661 (N_661,In_1466,In_206);
nand U662 (N_662,In_22,In_1798);
and U663 (N_663,In_3,In_260);
or U664 (N_664,In_2941,In_1145);
xnor U665 (N_665,In_355,In_970);
nand U666 (N_666,In_2179,In_1094);
xor U667 (N_667,In_458,In_2891);
and U668 (N_668,In_70,In_2658);
nand U669 (N_669,In_1888,In_1117);
or U670 (N_670,In_2007,In_1361);
and U671 (N_671,In_2197,In_869);
nor U672 (N_672,In_265,In_1882);
or U673 (N_673,In_1501,In_2033);
and U674 (N_674,In_1682,In_2665);
or U675 (N_675,In_2801,In_787);
or U676 (N_676,In_251,In_830);
or U677 (N_677,In_1624,In_2703);
nand U678 (N_678,In_1887,In_903);
nand U679 (N_679,In_456,In_298);
or U680 (N_680,In_1722,In_102);
xnor U681 (N_681,In_2569,In_1987);
nor U682 (N_682,In_1422,In_2355);
nand U683 (N_683,In_1526,In_727);
xnor U684 (N_684,In_1086,In_1142);
or U685 (N_685,In_382,In_1985);
or U686 (N_686,In_2736,In_2608);
and U687 (N_687,In_2948,In_2632);
or U688 (N_688,In_240,In_2001);
nand U689 (N_689,In_625,In_87);
nand U690 (N_690,In_1715,In_2884);
nand U691 (N_691,In_325,In_2737);
or U692 (N_692,In_331,In_2068);
xor U693 (N_693,In_2444,In_1743);
nand U694 (N_694,In_2135,In_52);
xor U695 (N_695,In_2959,In_2396);
nand U696 (N_696,In_2120,In_1783);
or U697 (N_697,In_1948,In_550);
nand U698 (N_698,In_2346,In_1801);
nor U699 (N_699,In_2386,In_2031);
nand U700 (N_700,In_1141,In_1958);
nor U701 (N_701,In_83,In_2143);
xnor U702 (N_702,In_2118,In_1891);
nand U703 (N_703,In_526,In_1003);
or U704 (N_704,In_279,In_736);
or U705 (N_705,In_2784,In_2313);
nand U706 (N_706,In_2555,In_467);
or U707 (N_707,In_2080,In_288);
nand U708 (N_708,In_964,In_615);
nand U709 (N_709,In_2064,In_1913);
nor U710 (N_710,In_2028,In_1959);
xnor U711 (N_711,In_364,In_2572);
nand U712 (N_712,In_2968,In_239);
or U713 (N_713,In_1217,In_2336);
nor U714 (N_714,In_53,In_1180);
xnor U715 (N_715,In_2556,In_1615);
xor U716 (N_716,In_1629,In_269);
nor U717 (N_717,In_2542,In_845);
or U718 (N_718,In_1806,In_2133);
or U719 (N_719,In_2942,In_605);
and U720 (N_720,In_1384,In_734);
nor U721 (N_721,In_2558,In_2158);
xor U722 (N_722,In_2502,In_594);
nand U723 (N_723,In_2276,In_2395);
or U724 (N_724,In_2402,In_865);
xor U725 (N_725,In_1465,In_1786);
xnor U726 (N_726,In_1561,In_882);
nand U727 (N_727,In_995,In_1467);
xnor U728 (N_728,In_2953,In_2949);
and U729 (N_729,In_983,In_1502);
or U730 (N_730,In_1111,In_1766);
or U731 (N_731,In_137,In_255);
nand U732 (N_732,In_2252,In_1015);
and U733 (N_733,In_1819,In_2758);
nand U734 (N_734,In_1392,In_2588);
nand U735 (N_735,In_422,In_2857);
or U736 (N_736,In_1613,In_228);
nor U737 (N_737,In_471,In_1375);
or U738 (N_738,In_735,In_404);
nand U739 (N_739,In_1626,In_831);
or U740 (N_740,In_1448,In_2232);
nor U741 (N_741,In_918,In_1253);
and U742 (N_742,In_2905,In_1521);
and U743 (N_743,In_934,In_2170);
xor U744 (N_744,In_323,In_868);
or U745 (N_745,In_2789,In_823);
xor U746 (N_746,In_1851,In_560);
nand U747 (N_747,In_854,In_565);
nor U748 (N_748,In_340,In_2867);
nor U749 (N_749,In_2352,In_1326);
and U750 (N_750,In_1650,In_610);
or U751 (N_751,In_1576,In_520);
nor U752 (N_752,In_928,In_38);
or U753 (N_753,In_2635,In_1460);
and U754 (N_754,In_1080,In_2792);
nand U755 (N_755,In_1499,In_2537);
nand U756 (N_756,In_1181,In_455);
and U757 (N_757,In_1815,In_2636);
and U758 (N_758,In_989,In_2344);
xnor U759 (N_759,In_2587,In_816);
nand U760 (N_760,In_1974,In_2914);
nor U761 (N_761,In_1755,In_247);
nor U762 (N_762,In_321,In_1671);
xor U763 (N_763,In_1956,In_1642);
xor U764 (N_764,In_1623,In_2166);
and U765 (N_765,In_2888,In_2);
xor U766 (N_766,In_1566,In_2694);
nor U767 (N_767,In_2721,In_1472);
and U768 (N_768,In_838,In_597);
xnor U769 (N_769,In_1380,In_1990);
nor U770 (N_770,In_986,In_1534);
nor U771 (N_771,In_2543,In_347);
nand U772 (N_772,In_2229,In_1178);
xnor U773 (N_773,In_1704,In_385);
nor U774 (N_774,In_459,In_46);
and U775 (N_775,In_23,In_2138);
xor U776 (N_776,In_15,In_1516);
nor U777 (N_777,In_618,In_2407);
nand U778 (N_778,In_1074,In_1050);
nand U779 (N_779,In_551,In_1364);
nor U780 (N_780,In_1617,In_203);
or U781 (N_781,In_670,In_1510);
xnor U782 (N_782,In_2185,In_491);
xnor U783 (N_783,In_1121,In_488);
nand U784 (N_784,In_2284,In_784);
nand U785 (N_785,In_115,In_1058);
or U786 (N_786,In_1598,In_1345);
or U787 (N_787,In_1323,In_785);
xor U788 (N_788,In_955,In_463);
xnor U789 (N_789,In_1313,In_1406);
xnor U790 (N_790,In_2814,In_524);
and U791 (N_791,In_2472,In_835);
nor U792 (N_792,In_559,In_2661);
nand U793 (N_793,In_2013,In_2299);
and U794 (N_794,In_568,In_412);
or U795 (N_795,In_1599,In_1277);
or U796 (N_796,In_2751,In_2811);
nor U797 (N_797,In_141,In_1269);
xnor U798 (N_798,In_468,In_1927);
nor U799 (N_799,In_1796,In_2691);
nor U800 (N_800,In_2282,In_2184);
nor U801 (N_801,In_2293,In_1591);
and U802 (N_802,In_2217,In_912);
and U803 (N_803,In_402,In_1196);
xor U804 (N_804,In_1104,In_697);
xor U805 (N_805,In_1909,In_116);
or U806 (N_806,In_534,In_2828);
xor U807 (N_807,In_1351,In_2319);
nor U808 (N_808,In_1803,In_78);
or U809 (N_809,In_2697,In_2797);
or U810 (N_810,In_1750,In_1983);
nand U811 (N_811,In_1445,In_2305);
nor U812 (N_812,In_190,In_584);
nand U813 (N_813,In_2393,In_1710);
or U814 (N_814,In_57,In_2527);
and U815 (N_815,In_2969,In_2794);
nand U816 (N_816,In_1033,In_266);
nand U817 (N_817,In_2886,In_496);
or U818 (N_818,In_2285,In_2144);
nor U819 (N_819,In_246,In_2441);
and U820 (N_820,In_1984,In_2279);
nor U821 (N_821,In_2681,In_272);
xor U822 (N_822,In_2719,In_1673);
and U823 (N_823,In_317,In_1436);
nand U824 (N_824,In_1129,In_1149);
nor U825 (N_825,In_580,In_2203);
nor U826 (N_826,In_1103,In_1622);
or U827 (N_827,In_2799,In_2224);
or U828 (N_828,In_960,In_1222);
or U829 (N_829,In_959,In_405);
nand U830 (N_830,In_1492,In_803);
nand U831 (N_831,In_473,In_1400);
and U832 (N_832,In_1286,In_2480);
and U833 (N_833,In_2063,In_1807);
nor U834 (N_834,In_505,In_1720);
nor U835 (N_835,In_1020,In_1694);
nor U836 (N_836,In_516,In_2427);
nand U837 (N_837,In_1932,In_2176);
and U838 (N_838,In_585,In_2743);
nor U839 (N_839,In_1317,In_1437);
nand U840 (N_840,In_1358,In_1477);
or U841 (N_841,In_2861,In_622);
or U842 (N_842,In_59,In_566);
and U843 (N_843,In_2773,In_1788);
and U844 (N_844,In_2038,In_2066);
xnor U845 (N_845,In_2903,In_2780);
and U846 (N_846,In_1365,In_1333);
nand U847 (N_847,In_797,In_1258);
nand U848 (N_848,In_2988,In_744);
nor U849 (N_849,In_1808,In_726);
xor U850 (N_850,In_1612,In_437);
or U851 (N_851,In_760,In_2300);
nor U852 (N_852,In_1972,In_2403);
or U853 (N_853,In_1768,In_1575);
nand U854 (N_854,In_2106,In_1255);
xnor U855 (N_855,In_212,In_2145);
and U856 (N_856,In_2265,In_2373);
and U857 (N_857,In_2511,In_2042);
xor U858 (N_858,In_2107,In_2650);
nor U859 (N_859,In_881,In_2032);
nor U860 (N_860,In_1081,In_1091);
or U861 (N_861,In_616,In_1337);
or U862 (N_862,In_2146,In_153);
nand U863 (N_863,In_61,In_1280);
nand U864 (N_864,In_789,In_2806);
or U865 (N_865,In_696,In_1359);
nor U866 (N_866,In_1125,In_757);
nor U867 (N_867,In_1068,In_1865);
xor U868 (N_868,In_543,In_2929);
nor U869 (N_869,In_1845,In_631);
nor U870 (N_870,In_1509,In_2073);
and U871 (N_871,In_689,In_361);
nor U872 (N_872,In_238,In_1728);
nand U873 (N_873,In_632,In_1449);
and U874 (N_874,In_790,In_1828);
nor U875 (N_875,In_1223,In_671);
xnor U876 (N_876,In_1525,In_2174);
nand U877 (N_877,In_2800,In_2754);
or U878 (N_878,In_939,In_1027);
and U879 (N_879,In_1108,In_721);
xor U880 (N_880,In_904,In_981);
xor U881 (N_881,In_809,In_967);
xor U882 (N_882,In_1747,In_1295);
or U883 (N_883,In_1331,In_603);
xor U884 (N_884,In_2191,In_285);
and U885 (N_885,In_1714,In_2878);
or U886 (N_886,In_652,In_66);
nand U887 (N_887,In_2955,In_2183);
nand U888 (N_888,In_2208,In_802);
and U889 (N_889,In_1066,In_386);
nor U890 (N_890,In_899,In_368);
xor U891 (N_891,In_339,In_130);
xor U892 (N_892,In_1771,In_2097);
nand U893 (N_893,In_1292,In_2561);
nand U894 (N_894,In_673,In_888);
nand U895 (N_895,In_1424,In_2416);
xor U896 (N_896,In_1742,In_732);
nand U897 (N_897,In_866,In_1842);
and U898 (N_898,In_910,In_1608);
or U899 (N_899,In_335,In_1075);
or U900 (N_900,In_2159,In_1199);
and U901 (N_901,In_993,In_1340);
or U902 (N_902,In_540,In_897);
xor U903 (N_903,In_2095,In_500);
or U904 (N_904,In_2399,In_1444);
and U905 (N_905,In_862,In_1844);
nand U906 (N_906,In_2204,In_2178);
nor U907 (N_907,In_426,In_161);
nand U908 (N_908,In_201,In_2766);
and U909 (N_909,In_2631,In_2597);
and U910 (N_910,In_242,In_2274);
nor U911 (N_911,In_2782,In_2233);
nand U912 (N_912,In_1672,In_1328);
and U913 (N_913,In_1433,In_1724);
nor U914 (N_914,In_2822,In_173);
and U915 (N_915,In_2538,In_2296);
nand U916 (N_916,In_154,In_27);
nor U917 (N_917,In_713,In_1494);
xor U918 (N_918,In_1604,In_2431);
and U919 (N_919,In_2809,In_1006);
xor U920 (N_920,In_1967,In_971);
or U921 (N_921,In_1009,In_684);
and U922 (N_922,In_1241,In_96);
xor U923 (N_923,In_316,In_310);
nand U924 (N_924,In_1729,In_1606);
and U925 (N_925,In_1471,In_872);
nor U926 (N_926,In_799,In_1026);
nand U927 (N_927,In_1036,In_1778);
nor U928 (N_928,In_1441,In_2777);
nand U929 (N_929,In_1837,In_522);
nor U930 (N_930,In_19,In_2678);
nor U931 (N_931,In_479,In_2280);
nor U932 (N_932,In_1998,In_2759);
xor U933 (N_933,In_110,In_1770);
or U934 (N_934,In_692,In_651);
nor U935 (N_935,In_1536,In_1939);
nor U936 (N_936,In_1434,In_303);
and U937 (N_937,In_1171,In_2322);
or U938 (N_938,In_2593,In_1296);
nor U939 (N_939,In_2895,In_1165);
nand U940 (N_940,In_2366,In_833);
and U941 (N_941,In_1737,In_2102);
and U942 (N_942,In_1892,In_742);
or U943 (N_943,In_1942,In_2332);
xor U944 (N_944,In_2457,In_1621);
xor U945 (N_945,In_1541,In_661);
nand U946 (N_946,In_1046,In_572);
xor U947 (N_947,In_2026,In_569);
and U948 (N_948,In_818,In_2842);
and U949 (N_949,In_1857,In_1628);
and U950 (N_950,In_1496,In_1731);
and U951 (N_951,In_2633,In_2966);
nand U952 (N_952,In_2998,In_1262);
and U953 (N_953,In_1054,In_2098);
or U954 (N_954,In_1377,In_1116);
or U955 (N_955,In_1556,In_1863);
nand U956 (N_956,In_2339,In_1443);
and U957 (N_957,In_2193,In_2369);
and U958 (N_958,In_184,In_145);
nor U959 (N_959,In_2354,In_2326);
nor U960 (N_960,In_2513,In_2499);
nand U961 (N_961,In_581,In_2024);
nand U962 (N_962,In_128,In_1298);
and U963 (N_963,In_2904,In_1992);
xnor U964 (N_964,In_2517,In_2005);
or U965 (N_965,In_1065,In_380);
nor U966 (N_966,In_156,In_730);
nor U967 (N_967,In_745,In_1479);
nand U968 (N_968,In_1825,In_1061);
or U969 (N_969,In_1166,In_1339);
nor U970 (N_970,In_1946,In_501);
nand U971 (N_971,In_1161,In_21);
xnor U972 (N_972,In_1873,In_1937);
nand U973 (N_973,In_1596,In_1527);
or U974 (N_974,In_2933,In_304);
and U975 (N_975,In_1226,In_388);
nor U976 (N_976,In_1835,In_2432);
or U977 (N_977,In_2989,In_2221);
and U978 (N_978,In_2687,In_2119);
or U979 (N_979,In_2035,In_177);
or U980 (N_980,In_1832,In_1138);
and U981 (N_981,In_2716,In_2560);
and U982 (N_982,In_2571,In_2869);
xnor U983 (N_983,In_963,In_669);
and U984 (N_984,In_332,In_493);
nor U985 (N_985,In_1916,In_466);
nand U986 (N_986,In_2422,In_2667);
and U987 (N_987,In_600,In_843);
or U988 (N_988,In_1335,In_451);
nor U989 (N_989,In_2958,In_217);
nand U990 (N_990,In_2839,In_1092);
and U991 (N_991,In_1893,In_414);
xor U992 (N_992,In_1519,In_1136);
nand U993 (N_993,In_1633,In_1485);
xnor U994 (N_994,In_1040,In_1637);
nand U995 (N_995,In_2331,In_1614);
and U996 (N_996,In_2245,In_2871);
or U997 (N_997,In_2115,In_2150);
and U998 (N_998,In_1620,In_1686);
xnor U999 (N_999,In_2973,In_2168);
nand U1000 (N_1000,In_86,In_391);
nor U1001 (N_1001,In_2550,In_1324);
and U1002 (N_1002,In_892,In_796);
xor U1003 (N_1003,In_290,In_638);
nor U1004 (N_1004,In_1169,In_2349);
and U1005 (N_1005,In_1202,In_1656);
xor U1006 (N_1006,In_2981,In_1684);
nand U1007 (N_1007,In_738,In_2496);
nor U1008 (N_1008,In_136,In_1706);
and U1009 (N_1009,In_1655,In_2630);
or U1010 (N_1010,In_2616,In_71);
xor U1011 (N_1011,In_913,In_1707);
xor U1012 (N_1012,In_484,In_124);
and U1013 (N_1013,In_596,In_1931);
nand U1014 (N_1014,In_119,In_2890);
nand U1015 (N_1015,In_1717,In_778);
nor U1016 (N_1016,In_464,In_2804);
and U1017 (N_1017,In_1961,In_148);
or U1018 (N_1018,In_1870,In_1549);
or U1019 (N_1019,In_2620,In_1346);
nor U1020 (N_1020,In_1394,In_593);
and U1021 (N_1021,In_826,In_1297);
xor U1022 (N_1022,In_519,In_1051);
or U1023 (N_1023,In_2415,In_185);
and U1024 (N_1024,In_1431,In_2882);
nand U1025 (N_1025,In_2760,In_1532);
and U1026 (N_1026,In_250,In_1657);
and U1027 (N_1027,In_991,In_232);
nor U1028 (N_1028,In_793,In_2523);
nand U1029 (N_1029,In_1189,In_2446);
nor U1030 (N_1030,In_360,In_1005);
nand U1031 (N_1031,In_2201,In_1156);
and U1032 (N_1032,In_1661,In_824);
or U1033 (N_1033,In_2471,In_85);
xor U1034 (N_1034,In_74,In_2817);
nand U1035 (N_1035,In_1531,In_1669);
nor U1036 (N_1036,In_1260,In_125);
and U1037 (N_1037,In_900,In_1497);
or U1038 (N_1038,In_2971,In_2149);
nand U1039 (N_1039,In_351,In_1977);
and U1040 (N_1040,In_30,In_956);
and U1041 (N_1041,In_2317,In_207);
xnor U1042 (N_1042,In_743,In_249);
xnor U1043 (N_1043,In_1372,In_1353);
and U1044 (N_1044,In_150,In_663);
or U1045 (N_1045,In_762,In_814);
and U1046 (N_1046,In_2206,In_2440);
xnor U1047 (N_1047,In_2414,In_312);
nand U1048 (N_1048,In_1659,In_1017);
or U1049 (N_1049,In_1636,In_801);
and U1050 (N_1050,In_1403,In_707);
nor U1051 (N_1051,In_417,In_1780);
nor U1052 (N_1052,In_2164,In_1968);
nand U1053 (N_1053,In_1670,In_457);
nor U1054 (N_1054,In_1303,In_1238);
nand U1055 (N_1055,In_1632,In_879);
or U1056 (N_1056,In_1969,In_1474);
xor U1057 (N_1057,In_2862,In_1334);
nor U1058 (N_1058,In_630,In_627);
or U1059 (N_1059,In_1455,In_1578);
xor U1060 (N_1060,In_1553,In_837);
nand U1061 (N_1061,In_1028,In_1373);
nand U1062 (N_1062,In_952,In_1925);
xnor U1063 (N_1063,In_512,In_507);
nor U1064 (N_1064,In_1563,In_2468);
or U1065 (N_1065,In_2826,In_1476);
and U1066 (N_1066,In_1903,In_2019);
or U1067 (N_1067,In_222,In_1446);
nand U1068 (N_1068,In_1537,In_1254);
and U1069 (N_1069,In_1368,In_234);
or U1070 (N_1070,In_1986,In_772);
xor U1071 (N_1071,In_1214,In_2724);
or U1072 (N_1072,In_1744,In_481);
xor U1073 (N_1073,In_767,In_1847);
or U1074 (N_1074,In_2477,In_2263);
nor U1075 (N_1075,In_2357,In_2918);
or U1076 (N_1076,In_2908,In_2889);
xnor U1077 (N_1077,In_2985,In_905);
nor U1078 (N_1078,In_2210,In_646);
nor U1079 (N_1079,In_2943,In_883);
nor U1080 (N_1080,In_1411,In_2504);
and U1081 (N_1081,In_169,In_2452);
xnor U1082 (N_1082,In_2974,In_2219);
and U1083 (N_1083,In_2141,In_2365);
or U1084 (N_1084,In_82,In_1084);
and U1085 (N_1085,In_2218,In_1055);
nor U1086 (N_1086,In_2078,In_424);
nand U1087 (N_1087,In_2919,In_2863);
xnor U1088 (N_1088,In_2105,In_719);
or U1089 (N_1089,In_1388,In_188);
xor U1090 (N_1090,In_755,In_1507);
and U1091 (N_1091,In_220,In_2753);
xor U1092 (N_1092,In_2894,In_2211);
nor U1093 (N_1093,In_2564,In_2096);
nor U1094 (N_1094,In_2901,In_1520);
nor U1095 (N_1095,In_274,In_2664);
or U1096 (N_1096,In_1605,In_400);
and U1097 (N_1097,In_1493,In_1450);
nor U1098 (N_1098,In_1203,In_149);
or U1099 (N_1099,In_393,In_2516);
xnor U1100 (N_1100,In_2054,In_2259);
nor U1101 (N_1101,In_887,In_40);
nor U1102 (N_1102,In_69,In_1473);
and U1103 (N_1103,In_81,In_1281);
and U1104 (N_1104,In_1063,In_2769);
or U1105 (N_1105,In_2334,In_2023);
nand U1106 (N_1106,In_961,In_2695);
nor U1107 (N_1107,In_1880,In_1872);
nand U1108 (N_1108,In_171,In_1374);
nand U1109 (N_1109,In_699,In_1634);
and U1110 (N_1110,In_341,In_1594);
xor U1111 (N_1111,In_2524,In_233);
and U1112 (N_1112,In_2376,In_372);
and U1113 (N_1113,In_2123,In_1256);
xnor U1114 (N_1114,In_1245,In_1290);
xor U1115 (N_1115,In_533,In_2677);
nand U1116 (N_1116,In_574,In_1988);
and U1117 (N_1117,In_538,In_2932);
xor U1118 (N_1118,In_1996,In_2022);
nand U1119 (N_1119,In_1567,In_2803);
or U1120 (N_1120,In_749,In_11);
nor U1121 (N_1121,In_1110,In_1396);
and U1122 (N_1122,In_860,In_1130);
or U1123 (N_1123,In_2079,In_330);
and U1124 (N_1124,In_2131,In_230);
or U1125 (N_1125,In_2505,In_235);
or U1126 (N_1126,In_134,In_1691);
nand U1127 (N_1127,In_1163,In_2846);
nor U1128 (N_1128,In_2475,In_771);
nand U1129 (N_1129,In_441,In_2243);
or U1130 (N_1130,In_1220,In_695);
and U1131 (N_1131,In_2071,In_462);
and U1132 (N_1132,In_2866,In_2979);
nor U1133 (N_1133,In_1530,In_1008);
nand U1134 (N_1134,In_2360,In_1157);
and U1135 (N_1135,In_1685,In_873);
xor U1136 (N_1136,In_2481,In_2675);
and U1137 (N_1137,In_1428,In_795);
nor U1138 (N_1138,In_327,In_1681);
nand U1139 (N_1139,In_645,In_1895);
and U1140 (N_1140,In_923,In_2844);
and U1141 (N_1141,In_123,In_1079);
or U1142 (N_1142,In_2815,In_1890);
or U1143 (N_1143,In_1201,In_654);
and U1144 (N_1144,In_1639,In_2012);
nand U1145 (N_1145,In_2272,In_1395);
xnor U1146 (N_1146,In_2275,In_1542);
xor U1147 (N_1147,In_1461,In_495);
or U1148 (N_1148,In_241,In_2235);
xor U1149 (N_1149,In_973,In_415);
xor U1150 (N_1150,In_2420,In_1447);
and U1151 (N_1151,In_563,In_268);
and U1152 (N_1152,In_1389,In_2108);
xor U1153 (N_1153,In_1309,In_676);
nand U1154 (N_1154,In_1971,In_2421);
nand U1155 (N_1155,In_1762,In_2478);
nor U1156 (N_1156,In_649,In_254);
and U1157 (N_1157,In_1600,In_365);
nor U1158 (N_1158,In_2562,In_1897);
nand U1159 (N_1159,In_204,In_371);
and U1160 (N_1160,In_1696,In_1154);
nand U1161 (N_1161,In_2586,In_925);
nor U1162 (N_1162,In_2187,In_135);
xnor U1163 (N_1163,In_1349,In_1653);
or U1164 (N_1164,In_2090,In_509);
xnor U1165 (N_1165,In_1965,In_1616);
and U1166 (N_1166,In_1350,In_1800);
xor U1167 (N_1167,In_2361,In_1416);
nand U1168 (N_1168,In_2389,In_1289);
or U1169 (N_1169,In_1928,In_1993);
or U1170 (N_1170,In_2362,In_315);
or U1171 (N_1171,In_1739,In_1144);
or U1172 (N_1172,In_2132,In_2591);
or U1173 (N_1173,In_2171,In_1688);
or U1174 (N_1174,In_2652,In_1740);
nor U1175 (N_1175,In_2896,In_2833);
and U1176 (N_1176,In_1533,In_624);
nor U1177 (N_1177,In_2634,In_2196);
and U1178 (N_1178,In_2735,In_1506);
or U1179 (N_1179,In_720,In_1573);
xnor U1180 (N_1180,In_2099,In_885);
nor U1181 (N_1181,In_1960,In_916);
nand U1182 (N_1182,In_2214,In_794);
or U1183 (N_1183,In_2075,In_2338);
nand U1184 (N_1184,In_1879,In_965);
or U1185 (N_1185,In_1442,In_1327);
or U1186 (N_1186,In_502,In_1902);
nand U1187 (N_1187,In_643,In_2489);
xor U1188 (N_1188,In_1638,In_1228);
nand U1189 (N_1189,In_2340,In_1848);
nor U1190 (N_1190,In_633,In_2008);
nor U1191 (N_1191,In_43,In_2865);
xnor U1192 (N_1192,In_1299,In_571);
and U1193 (N_1193,In_503,In_1733);
and U1194 (N_1194,In_2977,In_369);
nor U1195 (N_1195,In_357,In_842);
and U1196 (N_1196,In_1678,In_2310);
and U1197 (N_1197,In_2062,In_1738);
or U1198 (N_1198,In_936,In_1210);
xnor U1199 (N_1199,In_2162,In_2567);
and U1200 (N_1200,In_1216,In_2498);
or U1201 (N_1201,In_2649,In_1508);
and U1202 (N_1202,In_373,In_189);
or U1203 (N_1203,In_1589,In_658);
or U1204 (N_1204,In_2437,In_1221);
nand U1205 (N_1205,In_2671,In_1812);
xnor U1206 (N_1206,In_1831,In_2623);
xor U1207 (N_1207,In_1535,In_7);
and U1208 (N_1208,In_2686,In_1150);
or U1209 (N_1209,In_2964,In_2515);
xor U1210 (N_1210,In_2791,In_2648);
or U1211 (N_1211,In_1793,In_1045);
nand U1212 (N_1212,In_906,In_1412);
nand U1213 (N_1213,In_2497,In_2307);
or U1214 (N_1214,In_1912,In_2385);
or U1215 (N_1215,In_1581,In_162);
nand U1216 (N_1216,In_398,In_1607);
xnor U1217 (N_1217,In_113,In_529);
or U1218 (N_1218,In_1179,In_709);
nor U1219 (N_1219,In_2391,In_1726);
nor U1220 (N_1220,In_2067,In_2548);
nand U1221 (N_1221,In_2741,In_2136);
nor U1222 (N_1222,In_2821,In_182);
xor U1223 (N_1223,In_49,In_1763);
or U1224 (N_1224,In_1155,In_1078);
or U1225 (N_1225,In_515,In_2463);
nor U1226 (N_1226,In_261,In_282);
nand U1227 (N_1227,In_1794,In_1312);
nor U1228 (N_1228,In_461,In_138);
or U1229 (N_1229,In_774,In_700);
and U1230 (N_1230,In_1817,In_140);
xnor U1231 (N_1231,In_2913,In_2689);
nand U1232 (N_1232,In_2390,In_1076);
nand U1233 (N_1233,In_2029,In_446);
or U1234 (N_1234,In_1480,In_2412);
nand U1235 (N_1235,In_1357,In_183);
nor U1236 (N_1236,In_2910,In_2726);
and U1237 (N_1237,In_2877,In_1191);
or U1238 (N_1238,In_820,In_216);
and U1239 (N_1239,In_1250,In_1767);
nor U1240 (N_1240,In_1951,In_1764);
nor U1241 (N_1241,In_2439,In_2473);
xor U1242 (N_1242,In_51,In_2879);
or U1243 (N_1243,In_1758,In_2268);
or U1244 (N_1244,In_2018,In_1470);
xnor U1245 (N_1245,In_1732,In_1148);
xor U1246 (N_1246,In_1754,In_308);
nand U1247 (N_1247,In_1271,In_2093);
or U1248 (N_1248,In_1168,In_423);
or U1249 (N_1249,In_2812,In_1143);
xnor U1250 (N_1250,In_1919,In_2172);
or U1251 (N_1251,In_2841,In_1790);
xor U1252 (N_1252,In_2897,In_2121);
nor U1253 (N_1253,In_828,In_294);
xor U1254 (N_1254,In_313,In_2692);
nor U1255 (N_1255,In_2041,In_418);
and U1256 (N_1256,In_2153,In_2428);
nand U1257 (N_1257,In_1792,In_1167);
and U1258 (N_1258,In_929,In_2466);
or U1259 (N_1259,In_2165,In_849);
nand U1260 (N_1260,In_1748,In_408);
nor U1261 (N_1261,In_1410,In_34);
nand U1262 (N_1262,In_2816,In_1630);
and U1263 (N_1263,In_1195,In_1666);
nand U1264 (N_1264,In_2683,In_2192);
xor U1265 (N_1265,In_2714,In_710);
nor U1266 (N_1266,In_946,In_1668);
nor U1267 (N_1267,In_143,In_2585);
and U1268 (N_1268,In_1584,In_2907);
xnor U1269 (N_1269,In_2088,In_1544);
nand U1270 (N_1270,In_2316,In_152);
nand U1271 (N_1271,In_1784,In_2645);
or U1272 (N_1272,In_20,In_2433);
or U1273 (N_1273,In_1288,In_2147);
nand U1274 (N_1274,In_927,In_2823);
or U1275 (N_1275,In_1097,In_2058);
or U1276 (N_1276,In_2156,In_297);
nor U1277 (N_1277,In_80,In_225);
nor U1278 (N_1278,In_2353,In_58);
xnor U1279 (N_1279,In_1366,In_1098);
nand U1280 (N_1280,In_2320,In_748);
nor U1281 (N_1281,In_2612,In_348);
xor U1282 (N_1282,In_782,In_668);
nand U1283 (N_1283,In_2114,In_2710);
or U1284 (N_1284,In_10,In_690);
nand U1285 (N_1285,In_1332,In_2501);
or U1286 (N_1286,In_1609,In_2835);
or U1287 (N_1287,In_2713,In_2148);
nor U1288 (N_1288,In_2266,In_2931);
nor U1289 (N_1289,In_1318,In_1342);
nand U1290 (N_1290,In_374,In_2456);
nand U1291 (N_1291,In_694,In_47);
and U1292 (N_1292,In_1016,In_1224);
nor U1293 (N_1293,In_9,In_812);
or U1294 (N_1294,In_1515,In_108);
xor U1295 (N_1295,In_438,In_2774);
nor U1296 (N_1296,In_754,In_2787);
or U1297 (N_1297,In_2566,In_2994);
and U1298 (N_1298,In_1855,In_777);
and U1299 (N_1299,In_602,In_2601);
nand U1300 (N_1300,In_1952,In_2238);
nand U1301 (N_1301,In_1218,In_2993);
xnor U1302 (N_1302,In_2554,In_1979);
nor U1303 (N_1303,In_1585,In_867);
nor U1304 (N_1304,In_2641,In_2763);
nor U1305 (N_1305,In_2181,In_1231);
xnor U1306 (N_1306,In_2899,In_1347);
nor U1307 (N_1307,In_174,In_2205);
nor U1308 (N_1308,In_2582,In_781);
nor U1309 (N_1309,In_1746,In_328);
nor U1310 (N_1310,In_2476,In_0);
nand U1311 (N_1311,In_1024,In_2836);
or U1312 (N_1312,In_1,In_72);
and U1313 (N_1313,In_2627,In_759);
or U1314 (N_1314,In_1488,In_891);
nand U1315 (N_1315,In_2127,In_289);
xnor U1316 (N_1316,In_2924,In_685);
nand U1317 (N_1317,In_2350,In_1881);
nor U1318 (N_1318,In_1177,In_350);
and U1319 (N_1319,In_1239,In_1270);
or U1320 (N_1320,In_2764,In_2628);
or U1321 (N_1321,In_724,In_1935);
and U1322 (N_1322,In_2286,In_2281);
or U1323 (N_1323,In_2711,In_1899);
and U1324 (N_1324,In_1071,In_1010);
xnor U1325 (N_1325,In_1000,In_667);
or U1326 (N_1326,In_2945,In_804);
nand U1327 (N_1327,In_277,In_974);
and U1328 (N_1328,In_2016,In_886);
nand U1329 (N_1329,In_2874,In_2173);
and U1330 (N_1330,In_827,In_1367);
nor U1331 (N_1331,In_2536,In_1464);
nor U1332 (N_1332,In_2449,In_1813);
xor U1333 (N_1333,In_1287,In_2435);
nor U1334 (N_1334,In_641,In_1787);
xor U1335 (N_1335,In_2920,In_544);
or U1336 (N_1336,In_1423,In_338);
xor U1337 (N_1337,In_2301,In_852);
nor U1338 (N_1338,In_1115,In_1695);
or U1339 (N_1339,In_1308,In_686);
and U1340 (N_1340,In_2730,In_1072);
nor U1341 (N_1341,In_688,In_375);
xnor U1342 (N_1342,In_1153,In_1779);
and U1343 (N_1343,In_678,In_1073);
or U1344 (N_1344,In_2492,In_768);
xor U1345 (N_1345,In_2728,In_1252);
and U1346 (N_1346,In_2113,In_100);
xnor U1347 (N_1347,In_1336,In_1407);
or U1348 (N_1348,In_2987,In_800);
nor U1349 (N_1349,In_611,In_2963);
xnor U1350 (N_1350,In_497,In_433);
or U1351 (N_1351,In_1041,In_2081);
nand U1352 (N_1352,In_271,In_758);
and U1353 (N_1353,In_181,In_223);
nor U1354 (N_1354,In_32,In_2314);
xnor U1355 (N_1355,In_127,In_635);
nand U1356 (N_1356,In_807,In_517);
nand U1357 (N_1357,In_2590,In_2270);
xor U1358 (N_1358,In_992,In_60);
nand U1359 (N_1359,In_146,In_766);
or U1360 (N_1360,In_932,In_68);
nor U1361 (N_1361,In_356,In_262);
xnor U1362 (N_1362,In_202,In_1663);
and U1363 (N_1363,In_933,In_2250);
and U1364 (N_1364,In_1249,In_1757);
and U1365 (N_1365,In_553,In_2124);
or U1366 (N_1366,In_2129,In_1067);
nor U1367 (N_1367,In_12,In_1268);
xnor U1368 (N_1368,In_1404,In_1420);
xor U1369 (N_1369,In_2289,In_880);
xnor U1370 (N_1370,In_1677,In_1761);
and U1371 (N_1371,In_2783,In_541);
nand U1372 (N_1372,In_2089,In_1320);
or U1373 (N_1373,In_2727,In_1822);
xor U1374 (N_1374,In_2372,In_1718);
nor U1375 (N_1375,In_2573,In_98);
xnor U1376 (N_1376,In_948,In_132);
and U1377 (N_1377,In_2852,In_2824);
nand U1378 (N_1378,In_2598,In_1370);
nor U1379 (N_1379,In_2241,In_2182);
nand U1380 (N_1380,In_284,In_898);
and U1381 (N_1381,In_1934,In_2600);
and U1382 (N_1382,In_257,In_2581);
or U1383 (N_1383,In_2359,In_792);
xor U1384 (N_1384,In_199,In_2614);
nand U1385 (N_1385,In_2177,In_636);
or U1386 (N_1386,In_1032,In_2055);
xnor U1387 (N_1387,In_172,In_236);
and U1388 (N_1388,In_1938,In_1760);
nand U1389 (N_1389,In_1062,In_362);
xnor U1390 (N_1390,In_1582,In_698);
or U1391 (N_1391,In_811,In_2000);
xor U1392 (N_1392,In_521,In_1805);
or U1393 (N_1393,In_186,In_377);
nor U1394 (N_1394,In_2528,In_2408);
and U1395 (N_1395,In_2776,In_475);
or U1396 (N_1396,In_1025,In_1134);
nor U1397 (N_1397,In_1293,In_193);
xnor U1398 (N_1398,In_655,In_2425);
or U1399 (N_1399,In_1232,In_1646);
xnor U1400 (N_1400,In_1789,In_2380);
nand U1401 (N_1401,In_1291,In_1640);
or U1402 (N_1402,In_1341,In_2849);
nand U1403 (N_1403,In_746,In_999);
xnor U1404 (N_1404,In_1995,In_2535);
or U1405 (N_1405,In_498,In_1558);
or U1406 (N_1406,In_1172,In_1456);
and U1407 (N_1407,In_817,In_1077);
xnor U1408 (N_1408,In_579,In_1438);
nor U1409 (N_1409,In_704,In_370);
nor U1410 (N_1410,In_396,In_839);
and U1411 (N_1411,In_1248,In_1483);
and U1412 (N_1412,In_36,In_1487);
and U1413 (N_1413,In_2151,In_896);
or U1414 (N_1414,In_2594,In_822);
nand U1415 (N_1415,In_1304,In_2398);
nor U1416 (N_1416,In_2083,In_2574);
and U1417 (N_1417,In_723,In_706);
and U1418 (N_1418,In_1583,In_2384);
xor U1419 (N_1419,In_2002,In_1896);
or U1420 (N_1420,In_1059,In_561);
nand U1421 (N_1421,In_2303,In_1001);
nand U1422 (N_1422,In_1941,In_1603);
nand U1423 (N_1423,In_2043,In_1513);
xor U1424 (N_1424,In_1418,In_944);
xnor U1425 (N_1425,In_2198,In_1565);
and U1426 (N_1426,In_1915,In_1597);
or U1427 (N_1427,In_1869,In_523);
nor U1428 (N_1428,In_1002,In_2553);
and U1429 (N_1429,In_1898,In_2781);
nand U1430 (N_1430,In_2458,In_1877);
or U1431 (N_1431,In_1158,In_2829);
and U1432 (N_1432,In_2057,In_1551);
and U1433 (N_1433,In_2244,In_1975);
and U1434 (N_1434,In_2669,In_2306);
nor U1435 (N_1435,In_2911,In_810);
and U1436 (N_1436,In_1911,In_1132);
and U1437 (N_1437,In_2155,In_2292);
nand U1438 (N_1438,In_2246,In_806);
nor U1439 (N_1439,In_151,In_196);
nor U1440 (N_1440,In_750,In_2923);
nor U1441 (N_1441,In_1099,In_980);
nand U1442 (N_1442,In_92,In_2087);
xnor U1443 (N_1443,In_195,In_547);
nand U1444 (N_1444,In_2009,In_1243);
nor U1445 (N_1445,In_1102,In_231);
or U1446 (N_1446,In_1505,In_436);
or U1447 (N_1447,In_1227,In_2137);
or U1448 (N_1448,In_728,In_2216);
nor U1449 (N_1449,In_893,In_2467);
xnor U1450 (N_1450,In_401,In_2624);
nand U1451 (N_1451,In_48,In_949);
or U1452 (N_1452,In_1209,In_2577);
and U1453 (N_1453,In_376,In_1034);
nand U1454 (N_1454,In_2056,In_798);
and U1455 (N_1455,In_1693,In_1674);
and U1456 (N_1456,In_958,In_969);
and U1457 (N_1457,In_2061,In_296);
and U1458 (N_1458,In_664,In_425);
xor U1459 (N_1459,In_245,In_2419);
xnor U1460 (N_1460,In_2226,In_1885);
nor U1461 (N_1461,In_871,In_379);
or U1462 (N_1462,In_2954,In_1272);
and U1463 (N_1463,In_2207,In_1131);
and U1464 (N_1464,In_703,In_1843);
nand U1465 (N_1465,In_2249,In_2053);
xnor U1466 (N_1466,In_1994,In_1379);
nor U1467 (N_1467,In_1378,In_2819);
nand U1468 (N_1468,In_715,In_176);
and U1469 (N_1469,In_2957,In_1577);
nor U1470 (N_1470,In_2223,In_857);
or U1471 (N_1471,In_2668,In_545);
nand U1472 (N_1472,In_729,In_2534);
and U1473 (N_1473,In_1929,In_1517);
xor U1474 (N_1474,In_1867,In_1329);
nor U1475 (N_1475,In_2157,In_2676);
xnor U1476 (N_1476,In_1459,In_2657);
and U1477 (N_1477,In_465,In_1550);
nor U1478 (N_1478,In_2629,In_88);
or U1479 (N_1479,In_286,In_2315);
or U1480 (N_1480,In_175,In_2495);
or U1481 (N_1481,In_693,In_1490);
nor U1482 (N_1482,In_489,In_345);
or U1483 (N_1483,In_1275,In_972);
and U1484 (N_1484,In_2702,In_292);
or U1485 (N_1485,In_2483,In_431);
and U1486 (N_1486,In_163,In_37);
and U1487 (N_1487,In_121,In_2529);
or U1488 (N_1488,In_2725,In_2579);
or U1489 (N_1489,In_2240,In_2530);
or U1490 (N_1490,In_352,In_2796);
nand U1491 (N_1491,In_1052,In_2830);
nand U1492 (N_1492,In_2112,In_178);
and U1493 (N_1493,In_570,In_253);
nor U1494 (N_1494,In_77,In_1588);
or U1495 (N_1495,In_1963,In_2748);
and U1496 (N_1496,In_2004,In_2278);
xnor U1497 (N_1497,In_1237,In_1037);
nand U1498 (N_1498,In_856,In_821);
nor U1499 (N_1499,In_25,In_1876);
nor U1500 (N_1500,In_1772,In_455);
nand U1501 (N_1501,In_132,In_2280);
nor U1502 (N_1502,In_2528,In_423);
xor U1503 (N_1503,In_713,In_2440);
and U1504 (N_1504,In_452,In_1757);
xnor U1505 (N_1505,In_750,In_2613);
xnor U1506 (N_1506,In_1271,In_2965);
and U1507 (N_1507,In_1999,In_2627);
nand U1508 (N_1508,In_1618,In_1603);
and U1509 (N_1509,In_2931,In_1018);
and U1510 (N_1510,In_900,In_2025);
nand U1511 (N_1511,In_575,In_2939);
nor U1512 (N_1512,In_2588,In_2008);
nor U1513 (N_1513,In_514,In_1957);
xnor U1514 (N_1514,In_1430,In_1712);
xnor U1515 (N_1515,In_458,In_717);
nand U1516 (N_1516,In_697,In_1863);
or U1517 (N_1517,In_2036,In_1296);
nand U1518 (N_1518,In_1846,In_1826);
nor U1519 (N_1519,In_489,In_2430);
and U1520 (N_1520,In_612,In_769);
or U1521 (N_1521,In_807,In_1948);
xnor U1522 (N_1522,In_981,In_1165);
nor U1523 (N_1523,In_2763,In_2638);
nand U1524 (N_1524,In_747,In_2900);
nand U1525 (N_1525,In_975,In_1059);
xor U1526 (N_1526,In_2570,In_926);
or U1527 (N_1527,In_1212,In_1678);
nand U1528 (N_1528,In_1216,In_470);
nor U1529 (N_1529,In_1584,In_1120);
xnor U1530 (N_1530,In_862,In_1181);
and U1531 (N_1531,In_344,In_74);
nand U1532 (N_1532,In_797,In_2746);
nor U1533 (N_1533,In_1732,In_921);
nor U1534 (N_1534,In_2273,In_1884);
and U1535 (N_1535,In_2334,In_806);
and U1536 (N_1536,In_2614,In_253);
nor U1537 (N_1537,In_1054,In_1392);
xor U1538 (N_1538,In_513,In_1876);
xor U1539 (N_1539,In_262,In_2316);
and U1540 (N_1540,In_1330,In_753);
nor U1541 (N_1541,In_2477,In_1524);
nor U1542 (N_1542,In_2538,In_77);
xnor U1543 (N_1543,In_1228,In_2081);
nand U1544 (N_1544,In_1350,In_4);
xnor U1545 (N_1545,In_647,In_909);
nor U1546 (N_1546,In_1891,In_2926);
or U1547 (N_1547,In_2107,In_99);
xor U1548 (N_1548,In_1268,In_1569);
nand U1549 (N_1549,In_1239,In_1572);
and U1550 (N_1550,In_2280,In_1481);
or U1551 (N_1551,In_1992,In_1423);
nor U1552 (N_1552,In_1963,In_1923);
xor U1553 (N_1553,In_1673,In_1950);
nand U1554 (N_1554,In_137,In_703);
or U1555 (N_1555,In_2719,In_1791);
nor U1556 (N_1556,In_2666,In_126);
or U1557 (N_1557,In_2510,In_2050);
nand U1558 (N_1558,In_2485,In_2891);
xor U1559 (N_1559,In_2475,In_124);
or U1560 (N_1560,In_1324,In_2578);
xor U1561 (N_1561,In_2138,In_170);
nand U1562 (N_1562,In_2437,In_1015);
nand U1563 (N_1563,In_915,In_756);
or U1564 (N_1564,In_1384,In_821);
and U1565 (N_1565,In_2263,In_931);
xor U1566 (N_1566,In_923,In_1172);
or U1567 (N_1567,In_1062,In_277);
or U1568 (N_1568,In_877,In_1483);
nor U1569 (N_1569,In_1451,In_244);
nor U1570 (N_1570,In_2968,In_1614);
or U1571 (N_1571,In_2942,In_67);
or U1572 (N_1572,In_2393,In_1041);
or U1573 (N_1573,In_1304,In_2483);
nand U1574 (N_1574,In_1425,In_476);
nand U1575 (N_1575,In_576,In_1957);
xnor U1576 (N_1576,In_494,In_1899);
and U1577 (N_1577,In_336,In_1437);
and U1578 (N_1578,In_2913,In_2662);
nand U1579 (N_1579,In_2518,In_1092);
and U1580 (N_1580,In_849,In_2098);
or U1581 (N_1581,In_1529,In_1488);
nor U1582 (N_1582,In_2208,In_96);
or U1583 (N_1583,In_1099,In_2860);
or U1584 (N_1584,In_1734,In_2878);
and U1585 (N_1585,In_2970,In_1861);
or U1586 (N_1586,In_2578,In_885);
xor U1587 (N_1587,In_277,In_459);
nand U1588 (N_1588,In_1246,In_2240);
xnor U1589 (N_1589,In_1554,In_502);
xor U1590 (N_1590,In_35,In_2510);
nand U1591 (N_1591,In_197,In_2851);
nor U1592 (N_1592,In_2838,In_84);
nand U1593 (N_1593,In_133,In_1320);
nor U1594 (N_1594,In_1283,In_2756);
nand U1595 (N_1595,In_1867,In_331);
and U1596 (N_1596,In_2043,In_2084);
or U1597 (N_1597,In_2154,In_228);
nand U1598 (N_1598,In_2936,In_1249);
or U1599 (N_1599,In_1040,In_230);
nor U1600 (N_1600,In_2211,In_903);
nand U1601 (N_1601,In_1564,In_1414);
nor U1602 (N_1602,In_612,In_837);
or U1603 (N_1603,In_1995,In_597);
xnor U1604 (N_1604,In_56,In_695);
and U1605 (N_1605,In_1180,In_558);
and U1606 (N_1606,In_1699,In_2952);
xor U1607 (N_1607,In_2689,In_340);
and U1608 (N_1608,In_2720,In_1287);
or U1609 (N_1609,In_2974,In_1190);
or U1610 (N_1610,In_212,In_546);
nor U1611 (N_1611,In_710,In_911);
and U1612 (N_1612,In_1924,In_561);
nor U1613 (N_1613,In_1414,In_2652);
or U1614 (N_1614,In_430,In_2347);
or U1615 (N_1615,In_54,In_2140);
nor U1616 (N_1616,In_516,In_1667);
xor U1617 (N_1617,In_839,In_2357);
xor U1618 (N_1618,In_1346,In_672);
or U1619 (N_1619,In_2621,In_2722);
nor U1620 (N_1620,In_1962,In_1650);
nand U1621 (N_1621,In_587,In_2805);
and U1622 (N_1622,In_2387,In_750);
and U1623 (N_1623,In_1496,In_1268);
nor U1624 (N_1624,In_890,In_459);
and U1625 (N_1625,In_370,In_1792);
nand U1626 (N_1626,In_2083,In_1264);
nor U1627 (N_1627,In_1202,In_226);
and U1628 (N_1628,In_2046,In_856);
nor U1629 (N_1629,In_169,In_800);
nand U1630 (N_1630,In_1993,In_2576);
xor U1631 (N_1631,In_1579,In_2325);
nand U1632 (N_1632,In_1888,In_1620);
nor U1633 (N_1633,In_1668,In_833);
and U1634 (N_1634,In_2360,In_1390);
or U1635 (N_1635,In_2869,In_2350);
and U1636 (N_1636,In_1449,In_1210);
nor U1637 (N_1637,In_1928,In_2022);
nand U1638 (N_1638,In_1368,In_2970);
and U1639 (N_1639,In_745,In_394);
nor U1640 (N_1640,In_327,In_268);
nor U1641 (N_1641,In_2493,In_1968);
nand U1642 (N_1642,In_1391,In_493);
nor U1643 (N_1643,In_541,In_2237);
nand U1644 (N_1644,In_1732,In_293);
xnor U1645 (N_1645,In_1807,In_1860);
or U1646 (N_1646,In_1696,In_322);
and U1647 (N_1647,In_2365,In_2873);
or U1648 (N_1648,In_1564,In_165);
or U1649 (N_1649,In_584,In_1476);
and U1650 (N_1650,In_2793,In_1458);
nand U1651 (N_1651,In_2426,In_160);
nor U1652 (N_1652,In_1030,In_1903);
and U1653 (N_1653,In_1120,In_855);
or U1654 (N_1654,In_1976,In_2840);
nor U1655 (N_1655,In_949,In_380);
and U1656 (N_1656,In_132,In_262);
nor U1657 (N_1657,In_105,In_1736);
xnor U1658 (N_1658,In_44,In_925);
xnor U1659 (N_1659,In_412,In_1552);
xor U1660 (N_1660,In_2621,In_1217);
xnor U1661 (N_1661,In_1436,In_2375);
nor U1662 (N_1662,In_2852,In_425);
xor U1663 (N_1663,In_2201,In_1258);
nor U1664 (N_1664,In_1460,In_1257);
or U1665 (N_1665,In_69,In_2455);
xor U1666 (N_1666,In_231,In_2932);
or U1667 (N_1667,In_2282,In_2201);
or U1668 (N_1668,In_212,In_2901);
and U1669 (N_1669,In_384,In_1770);
nor U1670 (N_1670,In_1845,In_114);
or U1671 (N_1671,In_2798,In_502);
nand U1672 (N_1672,In_721,In_1531);
xnor U1673 (N_1673,In_2214,In_1843);
nand U1674 (N_1674,In_2938,In_1047);
or U1675 (N_1675,In_2174,In_731);
nor U1676 (N_1676,In_545,In_2125);
xor U1677 (N_1677,In_389,In_211);
and U1678 (N_1678,In_622,In_2914);
and U1679 (N_1679,In_74,In_621);
and U1680 (N_1680,In_2756,In_2725);
xnor U1681 (N_1681,In_2925,In_344);
nor U1682 (N_1682,In_401,In_2488);
nor U1683 (N_1683,In_1324,In_1552);
or U1684 (N_1684,In_521,In_1421);
xor U1685 (N_1685,In_2127,In_1356);
and U1686 (N_1686,In_394,In_1011);
xnor U1687 (N_1687,In_169,In_2770);
xor U1688 (N_1688,In_2139,In_879);
xor U1689 (N_1689,In_2006,In_1289);
xnor U1690 (N_1690,In_2116,In_1456);
nand U1691 (N_1691,In_959,In_1262);
nor U1692 (N_1692,In_716,In_2215);
nor U1693 (N_1693,In_667,In_1902);
xor U1694 (N_1694,In_2711,In_1384);
nand U1695 (N_1695,In_827,In_491);
xnor U1696 (N_1696,In_1077,In_1662);
nor U1697 (N_1697,In_518,In_632);
or U1698 (N_1698,In_1771,In_1491);
and U1699 (N_1699,In_1094,In_30);
nand U1700 (N_1700,In_94,In_1755);
nand U1701 (N_1701,In_1481,In_1517);
nor U1702 (N_1702,In_839,In_2094);
nor U1703 (N_1703,In_923,In_193);
nor U1704 (N_1704,In_1836,In_141);
or U1705 (N_1705,In_1871,In_2082);
or U1706 (N_1706,In_2702,In_1062);
nor U1707 (N_1707,In_717,In_1481);
or U1708 (N_1708,In_1551,In_875);
or U1709 (N_1709,In_270,In_2196);
or U1710 (N_1710,In_1882,In_87);
nand U1711 (N_1711,In_838,In_120);
and U1712 (N_1712,In_1804,In_2880);
xnor U1713 (N_1713,In_2055,In_1759);
and U1714 (N_1714,In_1826,In_1507);
xnor U1715 (N_1715,In_1860,In_2782);
nor U1716 (N_1716,In_746,In_473);
or U1717 (N_1717,In_916,In_1706);
or U1718 (N_1718,In_2189,In_2299);
xnor U1719 (N_1719,In_2045,In_2508);
and U1720 (N_1720,In_1034,In_2619);
and U1721 (N_1721,In_2548,In_2883);
xor U1722 (N_1722,In_862,In_887);
xnor U1723 (N_1723,In_2463,In_1099);
xor U1724 (N_1724,In_841,In_1137);
and U1725 (N_1725,In_1510,In_1692);
nand U1726 (N_1726,In_1807,In_2418);
nor U1727 (N_1727,In_490,In_1679);
nor U1728 (N_1728,In_2656,In_918);
nor U1729 (N_1729,In_907,In_614);
nor U1730 (N_1730,In_889,In_2249);
xnor U1731 (N_1731,In_165,In_2330);
nor U1732 (N_1732,In_1962,In_1010);
nor U1733 (N_1733,In_2603,In_2825);
or U1734 (N_1734,In_2175,In_1195);
and U1735 (N_1735,In_745,In_2094);
nor U1736 (N_1736,In_2450,In_1756);
and U1737 (N_1737,In_1992,In_2066);
or U1738 (N_1738,In_1465,In_1423);
or U1739 (N_1739,In_710,In_1190);
and U1740 (N_1740,In_695,In_1036);
nor U1741 (N_1741,In_380,In_2515);
nand U1742 (N_1742,In_2989,In_2233);
nand U1743 (N_1743,In_1646,In_1575);
nor U1744 (N_1744,In_2636,In_2621);
and U1745 (N_1745,In_1233,In_887);
and U1746 (N_1746,In_779,In_2256);
and U1747 (N_1747,In_1815,In_1267);
xnor U1748 (N_1748,In_2626,In_1206);
xor U1749 (N_1749,In_2422,In_2802);
and U1750 (N_1750,In_2497,In_2335);
and U1751 (N_1751,In_575,In_1841);
and U1752 (N_1752,In_1924,In_2984);
nand U1753 (N_1753,In_75,In_1848);
nor U1754 (N_1754,In_2823,In_2662);
or U1755 (N_1755,In_891,In_2755);
xnor U1756 (N_1756,In_2458,In_1522);
nor U1757 (N_1757,In_200,In_153);
nand U1758 (N_1758,In_252,In_774);
or U1759 (N_1759,In_922,In_583);
and U1760 (N_1760,In_2131,In_1460);
or U1761 (N_1761,In_371,In_2580);
and U1762 (N_1762,In_2550,In_540);
and U1763 (N_1763,In_2624,In_1349);
xnor U1764 (N_1764,In_2433,In_1433);
xor U1765 (N_1765,In_701,In_2810);
or U1766 (N_1766,In_325,In_564);
or U1767 (N_1767,In_1387,In_1469);
nor U1768 (N_1768,In_2920,In_1119);
and U1769 (N_1769,In_599,In_2487);
nor U1770 (N_1770,In_439,In_480);
nand U1771 (N_1771,In_636,In_1389);
and U1772 (N_1772,In_762,In_1781);
nand U1773 (N_1773,In_2884,In_2501);
nor U1774 (N_1774,In_1873,In_2632);
or U1775 (N_1775,In_255,In_2341);
and U1776 (N_1776,In_1672,In_2243);
nor U1777 (N_1777,In_670,In_2909);
xor U1778 (N_1778,In_2974,In_1840);
xnor U1779 (N_1779,In_1208,In_1407);
xor U1780 (N_1780,In_826,In_1965);
or U1781 (N_1781,In_625,In_379);
nor U1782 (N_1782,In_3,In_2285);
nand U1783 (N_1783,In_615,In_1962);
nor U1784 (N_1784,In_2947,In_2989);
or U1785 (N_1785,In_1668,In_954);
nand U1786 (N_1786,In_375,In_1258);
and U1787 (N_1787,In_2824,In_2837);
nand U1788 (N_1788,In_1149,In_2599);
nand U1789 (N_1789,In_2089,In_1572);
xnor U1790 (N_1790,In_20,In_1170);
and U1791 (N_1791,In_2997,In_1667);
nand U1792 (N_1792,In_253,In_2199);
or U1793 (N_1793,In_2594,In_2772);
and U1794 (N_1794,In_557,In_174);
xor U1795 (N_1795,In_2032,In_1060);
nor U1796 (N_1796,In_233,In_2711);
and U1797 (N_1797,In_103,In_1709);
nor U1798 (N_1798,In_743,In_2529);
and U1799 (N_1799,In_1212,In_1239);
and U1800 (N_1800,In_2801,In_138);
xnor U1801 (N_1801,In_2831,In_1447);
and U1802 (N_1802,In_2293,In_2182);
and U1803 (N_1803,In_2583,In_2170);
and U1804 (N_1804,In_2867,In_2865);
nor U1805 (N_1805,In_391,In_2299);
xnor U1806 (N_1806,In_1057,In_2057);
nand U1807 (N_1807,In_1246,In_2586);
or U1808 (N_1808,In_1399,In_34);
and U1809 (N_1809,In_304,In_2388);
nand U1810 (N_1810,In_1737,In_2849);
nor U1811 (N_1811,In_1346,In_920);
and U1812 (N_1812,In_390,In_260);
and U1813 (N_1813,In_2972,In_777);
nand U1814 (N_1814,In_2109,In_926);
nand U1815 (N_1815,In_46,In_391);
xnor U1816 (N_1816,In_1764,In_2288);
nor U1817 (N_1817,In_15,In_2356);
and U1818 (N_1818,In_1812,In_520);
nand U1819 (N_1819,In_895,In_2678);
nor U1820 (N_1820,In_2902,In_2820);
xnor U1821 (N_1821,In_1113,In_2958);
and U1822 (N_1822,In_2704,In_2453);
and U1823 (N_1823,In_2043,In_622);
and U1824 (N_1824,In_540,In_142);
xnor U1825 (N_1825,In_2112,In_2264);
xor U1826 (N_1826,In_1169,In_143);
nor U1827 (N_1827,In_1540,In_1947);
xnor U1828 (N_1828,In_1870,In_2339);
or U1829 (N_1829,In_2905,In_2065);
nor U1830 (N_1830,In_1565,In_1180);
xnor U1831 (N_1831,In_2403,In_806);
nand U1832 (N_1832,In_2479,In_794);
or U1833 (N_1833,In_2723,In_1960);
xnor U1834 (N_1834,In_625,In_439);
or U1835 (N_1835,In_1420,In_2563);
nand U1836 (N_1836,In_2052,In_2965);
nor U1837 (N_1837,In_1851,In_591);
nand U1838 (N_1838,In_2916,In_623);
nor U1839 (N_1839,In_376,In_2309);
xnor U1840 (N_1840,In_504,In_1068);
xnor U1841 (N_1841,In_2197,In_2203);
nor U1842 (N_1842,In_2338,In_2473);
or U1843 (N_1843,In_1354,In_268);
nor U1844 (N_1844,In_2935,In_1992);
nor U1845 (N_1845,In_1886,In_1729);
or U1846 (N_1846,In_2325,In_191);
nor U1847 (N_1847,In_1621,In_2897);
and U1848 (N_1848,In_322,In_2532);
nor U1849 (N_1849,In_987,In_2306);
and U1850 (N_1850,In_1380,In_1610);
xnor U1851 (N_1851,In_2821,In_1927);
nor U1852 (N_1852,In_899,In_2440);
nand U1853 (N_1853,In_356,In_344);
nor U1854 (N_1854,In_1960,In_649);
and U1855 (N_1855,In_604,In_123);
or U1856 (N_1856,In_522,In_1746);
xnor U1857 (N_1857,In_1444,In_2955);
or U1858 (N_1858,In_1116,In_771);
xor U1859 (N_1859,In_883,In_1200);
nand U1860 (N_1860,In_1692,In_2766);
nand U1861 (N_1861,In_1292,In_1379);
xor U1862 (N_1862,In_1582,In_2991);
and U1863 (N_1863,In_2815,In_1773);
or U1864 (N_1864,In_2383,In_459);
and U1865 (N_1865,In_2181,In_721);
nand U1866 (N_1866,In_2357,In_788);
nand U1867 (N_1867,In_1287,In_2127);
nand U1868 (N_1868,In_1265,In_477);
and U1869 (N_1869,In_1545,In_801);
xor U1870 (N_1870,In_2552,In_2206);
or U1871 (N_1871,In_1899,In_481);
nand U1872 (N_1872,In_2675,In_2967);
xnor U1873 (N_1873,In_2124,In_984);
nand U1874 (N_1874,In_760,In_1593);
nand U1875 (N_1875,In_758,In_2777);
nor U1876 (N_1876,In_610,In_457);
and U1877 (N_1877,In_646,In_1113);
nand U1878 (N_1878,In_2887,In_488);
xnor U1879 (N_1879,In_2003,In_2190);
or U1880 (N_1880,In_1772,In_2759);
xnor U1881 (N_1881,In_2543,In_2729);
or U1882 (N_1882,In_2345,In_2118);
or U1883 (N_1883,In_1160,In_2129);
or U1884 (N_1884,In_323,In_727);
or U1885 (N_1885,In_681,In_1904);
nand U1886 (N_1886,In_487,In_1543);
nor U1887 (N_1887,In_2484,In_2165);
nor U1888 (N_1888,In_934,In_793);
and U1889 (N_1889,In_2738,In_1546);
or U1890 (N_1890,In_661,In_1807);
xor U1891 (N_1891,In_160,In_197);
nor U1892 (N_1892,In_222,In_1042);
nand U1893 (N_1893,In_1946,In_2677);
nand U1894 (N_1894,In_1902,In_297);
xnor U1895 (N_1895,In_1283,In_2966);
nand U1896 (N_1896,In_2474,In_1766);
xnor U1897 (N_1897,In_1715,In_645);
xor U1898 (N_1898,In_1834,In_1398);
nor U1899 (N_1899,In_2762,In_1688);
xor U1900 (N_1900,In_493,In_187);
and U1901 (N_1901,In_2238,In_83);
nand U1902 (N_1902,In_1222,In_1587);
nand U1903 (N_1903,In_2005,In_1718);
and U1904 (N_1904,In_855,In_752);
nand U1905 (N_1905,In_2801,In_376);
or U1906 (N_1906,In_635,In_2585);
and U1907 (N_1907,In_2634,In_1949);
and U1908 (N_1908,In_2924,In_1443);
and U1909 (N_1909,In_647,In_126);
nand U1910 (N_1910,In_966,In_746);
xor U1911 (N_1911,In_73,In_233);
xor U1912 (N_1912,In_540,In_377);
nand U1913 (N_1913,In_549,In_989);
and U1914 (N_1914,In_1937,In_997);
or U1915 (N_1915,In_1784,In_652);
xor U1916 (N_1916,In_482,In_2769);
xnor U1917 (N_1917,In_2069,In_1636);
nor U1918 (N_1918,In_2495,In_2300);
nor U1919 (N_1919,In_354,In_2757);
xnor U1920 (N_1920,In_2440,In_2863);
xnor U1921 (N_1921,In_785,In_1906);
nand U1922 (N_1922,In_813,In_2340);
nand U1923 (N_1923,In_811,In_1171);
nor U1924 (N_1924,In_2346,In_305);
nand U1925 (N_1925,In_1904,In_2007);
or U1926 (N_1926,In_1633,In_1197);
and U1927 (N_1927,In_1282,In_1344);
nor U1928 (N_1928,In_1150,In_2216);
nand U1929 (N_1929,In_747,In_1413);
and U1930 (N_1930,In_760,In_1219);
and U1931 (N_1931,In_2893,In_1396);
or U1932 (N_1932,In_2111,In_1900);
or U1933 (N_1933,In_2755,In_1819);
nor U1934 (N_1934,In_446,In_2600);
xor U1935 (N_1935,In_2606,In_1072);
nor U1936 (N_1936,In_2909,In_348);
nor U1937 (N_1937,In_2792,In_1820);
and U1938 (N_1938,In_1925,In_1860);
and U1939 (N_1939,In_522,In_2247);
nor U1940 (N_1940,In_2911,In_896);
nor U1941 (N_1941,In_1408,In_1802);
and U1942 (N_1942,In_2478,In_1946);
nand U1943 (N_1943,In_2558,In_1516);
nand U1944 (N_1944,In_2227,In_2583);
xor U1945 (N_1945,In_238,In_2606);
xnor U1946 (N_1946,In_2194,In_202);
nand U1947 (N_1947,In_1723,In_923);
and U1948 (N_1948,In_150,In_2169);
and U1949 (N_1949,In_1711,In_643);
or U1950 (N_1950,In_2240,In_238);
nand U1951 (N_1951,In_1435,In_2935);
and U1952 (N_1952,In_2922,In_1057);
nand U1953 (N_1953,In_1893,In_762);
and U1954 (N_1954,In_1613,In_981);
nor U1955 (N_1955,In_1322,In_2691);
or U1956 (N_1956,In_884,In_1216);
and U1957 (N_1957,In_2450,In_538);
xnor U1958 (N_1958,In_685,In_2745);
or U1959 (N_1959,In_1847,In_1823);
or U1960 (N_1960,In_2277,In_226);
nor U1961 (N_1961,In_2798,In_2556);
nand U1962 (N_1962,In_2510,In_699);
or U1963 (N_1963,In_2979,In_495);
or U1964 (N_1964,In_2121,In_2241);
xnor U1965 (N_1965,In_981,In_1248);
or U1966 (N_1966,In_2411,In_1322);
or U1967 (N_1967,In_563,In_2600);
or U1968 (N_1968,In_1874,In_1127);
nand U1969 (N_1969,In_879,In_35);
nor U1970 (N_1970,In_2316,In_1141);
xor U1971 (N_1971,In_930,In_2680);
xnor U1972 (N_1972,In_2489,In_381);
and U1973 (N_1973,In_676,In_1737);
or U1974 (N_1974,In_1454,In_2242);
and U1975 (N_1975,In_174,In_1155);
xnor U1976 (N_1976,In_2774,In_565);
and U1977 (N_1977,In_297,In_2443);
and U1978 (N_1978,In_2297,In_1349);
or U1979 (N_1979,In_1313,In_1098);
nand U1980 (N_1980,In_1546,In_1857);
or U1981 (N_1981,In_852,In_993);
nand U1982 (N_1982,In_1678,In_287);
xor U1983 (N_1983,In_209,In_2609);
or U1984 (N_1984,In_2423,In_984);
xor U1985 (N_1985,In_183,In_1262);
or U1986 (N_1986,In_594,In_1433);
nand U1987 (N_1987,In_1915,In_1438);
nand U1988 (N_1988,In_235,In_708);
and U1989 (N_1989,In_186,In_65);
nand U1990 (N_1990,In_385,In_1867);
xor U1991 (N_1991,In_1788,In_1276);
nor U1992 (N_1992,In_727,In_2950);
nand U1993 (N_1993,In_399,In_1544);
nand U1994 (N_1994,In_1964,In_1374);
nand U1995 (N_1995,In_2687,In_1032);
or U1996 (N_1996,In_87,In_2826);
xnor U1997 (N_1997,In_1786,In_556);
and U1998 (N_1998,In_567,In_2754);
nor U1999 (N_1999,In_651,In_2361);
or U2000 (N_2000,In_1320,In_1646);
or U2001 (N_2001,In_995,In_169);
xnor U2002 (N_2002,In_1935,In_416);
xnor U2003 (N_2003,In_2000,In_116);
or U2004 (N_2004,In_1319,In_49);
nor U2005 (N_2005,In_800,In_807);
xor U2006 (N_2006,In_1129,In_2678);
xnor U2007 (N_2007,In_2316,In_2611);
or U2008 (N_2008,In_1679,In_19);
nand U2009 (N_2009,In_487,In_2448);
xor U2010 (N_2010,In_1613,In_4);
nand U2011 (N_2011,In_1936,In_2159);
nor U2012 (N_2012,In_1907,In_1318);
nand U2013 (N_2013,In_2020,In_1632);
nor U2014 (N_2014,In_1757,In_654);
nor U2015 (N_2015,In_874,In_1848);
nor U2016 (N_2016,In_247,In_1683);
nor U2017 (N_2017,In_1195,In_469);
xnor U2018 (N_2018,In_2413,In_675);
or U2019 (N_2019,In_2740,In_1336);
nor U2020 (N_2020,In_2062,In_1504);
nor U2021 (N_2021,In_528,In_1336);
nand U2022 (N_2022,In_1537,In_808);
nor U2023 (N_2023,In_2065,In_188);
nor U2024 (N_2024,In_1983,In_1485);
nand U2025 (N_2025,In_1800,In_1941);
nand U2026 (N_2026,In_801,In_1666);
nand U2027 (N_2027,In_1337,In_1300);
xor U2028 (N_2028,In_195,In_1694);
and U2029 (N_2029,In_1632,In_97);
nand U2030 (N_2030,In_903,In_1481);
or U2031 (N_2031,In_2341,In_612);
and U2032 (N_2032,In_1647,In_261);
nand U2033 (N_2033,In_2148,In_418);
or U2034 (N_2034,In_1419,In_2111);
or U2035 (N_2035,In_1217,In_1700);
nand U2036 (N_2036,In_1139,In_1187);
nand U2037 (N_2037,In_2876,In_1621);
or U2038 (N_2038,In_935,In_772);
or U2039 (N_2039,In_839,In_758);
nand U2040 (N_2040,In_480,In_1118);
nand U2041 (N_2041,In_2269,In_293);
nand U2042 (N_2042,In_1758,In_546);
xnor U2043 (N_2043,In_38,In_2460);
or U2044 (N_2044,In_1114,In_1262);
xor U2045 (N_2045,In_1542,In_1799);
nand U2046 (N_2046,In_2537,In_2714);
or U2047 (N_2047,In_2236,In_1444);
and U2048 (N_2048,In_2105,In_2806);
xnor U2049 (N_2049,In_2416,In_916);
nand U2050 (N_2050,In_1339,In_819);
xnor U2051 (N_2051,In_1945,In_2706);
and U2052 (N_2052,In_1721,In_2595);
nor U2053 (N_2053,In_620,In_1401);
or U2054 (N_2054,In_2137,In_2098);
or U2055 (N_2055,In_1420,In_2921);
nor U2056 (N_2056,In_469,In_1566);
xor U2057 (N_2057,In_1653,In_1655);
nor U2058 (N_2058,In_1907,In_2339);
nor U2059 (N_2059,In_1346,In_1224);
xor U2060 (N_2060,In_400,In_1742);
nand U2061 (N_2061,In_2521,In_1572);
nor U2062 (N_2062,In_803,In_46);
nor U2063 (N_2063,In_2912,In_2612);
or U2064 (N_2064,In_1101,In_552);
xnor U2065 (N_2065,In_1410,In_381);
or U2066 (N_2066,In_1130,In_1465);
or U2067 (N_2067,In_2716,In_1576);
xor U2068 (N_2068,In_1538,In_327);
or U2069 (N_2069,In_2394,In_1702);
nand U2070 (N_2070,In_1903,In_1227);
xor U2071 (N_2071,In_2324,In_2801);
or U2072 (N_2072,In_655,In_2823);
or U2073 (N_2073,In_2691,In_945);
nand U2074 (N_2074,In_643,In_1622);
xnor U2075 (N_2075,In_2688,In_106);
and U2076 (N_2076,In_2055,In_261);
nand U2077 (N_2077,In_1476,In_2024);
nand U2078 (N_2078,In_1808,In_2154);
nand U2079 (N_2079,In_1354,In_2634);
nor U2080 (N_2080,In_2974,In_1476);
nor U2081 (N_2081,In_1146,In_1240);
nor U2082 (N_2082,In_1225,In_2578);
or U2083 (N_2083,In_217,In_62);
xnor U2084 (N_2084,In_83,In_1424);
and U2085 (N_2085,In_1964,In_1404);
nor U2086 (N_2086,In_1367,In_964);
xor U2087 (N_2087,In_2224,In_85);
xor U2088 (N_2088,In_1880,In_2872);
or U2089 (N_2089,In_570,In_1457);
and U2090 (N_2090,In_2966,In_1211);
nand U2091 (N_2091,In_1636,In_2993);
xor U2092 (N_2092,In_1599,In_1585);
and U2093 (N_2093,In_2294,In_778);
or U2094 (N_2094,In_788,In_1769);
xnor U2095 (N_2095,In_742,In_905);
nand U2096 (N_2096,In_1518,In_55);
nor U2097 (N_2097,In_2952,In_2261);
xnor U2098 (N_2098,In_2506,In_1105);
xnor U2099 (N_2099,In_32,In_1086);
and U2100 (N_2100,In_553,In_1834);
nor U2101 (N_2101,In_1685,In_335);
nor U2102 (N_2102,In_1493,In_2189);
nand U2103 (N_2103,In_2658,In_2933);
or U2104 (N_2104,In_1817,In_976);
and U2105 (N_2105,In_422,In_932);
or U2106 (N_2106,In_1978,In_639);
xnor U2107 (N_2107,In_908,In_1165);
and U2108 (N_2108,In_1287,In_1580);
or U2109 (N_2109,In_756,In_2499);
nor U2110 (N_2110,In_1100,In_1308);
or U2111 (N_2111,In_1095,In_2546);
nand U2112 (N_2112,In_100,In_1778);
nor U2113 (N_2113,In_224,In_2684);
or U2114 (N_2114,In_2272,In_2365);
nand U2115 (N_2115,In_383,In_1594);
and U2116 (N_2116,In_2655,In_2783);
nor U2117 (N_2117,In_961,In_2668);
and U2118 (N_2118,In_1029,In_2495);
nand U2119 (N_2119,In_801,In_115);
nor U2120 (N_2120,In_2723,In_1155);
and U2121 (N_2121,In_2328,In_512);
nand U2122 (N_2122,In_1246,In_1200);
and U2123 (N_2123,In_1019,In_479);
and U2124 (N_2124,In_593,In_26);
and U2125 (N_2125,In_2984,In_2192);
nor U2126 (N_2126,In_568,In_227);
or U2127 (N_2127,In_574,In_2269);
nand U2128 (N_2128,In_1137,In_169);
nor U2129 (N_2129,In_1668,In_398);
nand U2130 (N_2130,In_1264,In_2758);
or U2131 (N_2131,In_2115,In_2853);
or U2132 (N_2132,In_1583,In_259);
and U2133 (N_2133,In_390,In_2608);
xor U2134 (N_2134,In_336,In_1351);
or U2135 (N_2135,In_32,In_1149);
and U2136 (N_2136,In_56,In_864);
nor U2137 (N_2137,In_2732,In_2575);
or U2138 (N_2138,In_2278,In_1291);
xor U2139 (N_2139,In_2624,In_1231);
xnor U2140 (N_2140,In_1233,In_1683);
or U2141 (N_2141,In_1947,In_489);
nand U2142 (N_2142,In_1178,In_2391);
nor U2143 (N_2143,In_224,In_1059);
xor U2144 (N_2144,In_1723,In_523);
nand U2145 (N_2145,In_2116,In_2931);
xnor U2146 (N_2146,In_418,In_2767);
nor U2147 (N_2147,In_2095,In_1572);
nand U2148 (N_2148,In_2709,In_39);
xor U2149 (N_2149,In_2338,In_1466);
nand U2150 (N_2150,In_2192,In_538);
nor U2151 (N_2151,In_214,In_961);
nand U2152 (N_2152,In_1789,In_2388);
nand U2153 (N_2153,In_726,In_860);
or U2154 (N_2154,In_1477,In_2549);
and U2155 (N_2155,In_2895,In_575);
nor U2156 (N_2156,In_669,In_1834);
nor U2157 (N_2157,In_2738,In_1830);
xor U2158 (N_2158,In_591,In_2436);
and U2159 (N_2159,In_2884,In_1180);
and U2160 (N_2160,In_105,In_626);
nor U2161 (N_2161,In_160,In_1732);
xor U2162 (N_2162,In_1198,In_441);
or U2163 (N_2163,In_281,In_1101);
or U2164 (N_2164,In_2294,In_678);
or U2165 (N_2165,In_1943,In_2379);
nand U2166 (N_2166,In_1120,In_1030);
and U2167 (N_2167,In_2969,In_2213);
nor U2168 (N_2168,In_2871,In_945);
nor U2169 (N_2169,In_2386,In_2073);
and U2170 (N_2170,In_1196,In_1020);
nor U2171 (N_2171,In_2945,In_983);
and U2172 (N_2172,In_1408,In_1661);
nor U2173 (N_2173,In_2465,In_1232);
xor U2174 (N_2174,In_839,In_7);
nor U2175 (N_2175,In_1758,In_1305);
nor U2176 (N_2176,In_2394,In_913);
nand U2177 (N_2177,In_2029,In_233);
nand U2178 (N_2178,In_1278,In_96);
nor U2179 (N_2179,In_2525,In_1204);
and U2180 (N_2180,In_641,In_1245);
nand U2181 (N_2181,In_1553,In_2493);
and U2182 (N_2182,In_1004,In_137);
and U2183 (N_2183,In_1719,In_1619);
and U2184 (N_2184,In_244,In_1113);
xnor U2185 (N_2185,In_2113,In_491);
and U2186 (N_2186,In_615,In_1003);
and U2187 (N_2187,In_185,In_790);
and U2188 (N_2188,In_1546,In_1338);
or U2189 (N_2189,In_495,In_75);
and U2190 (N_2190,In_1708,In_2569);
xor U2191 (N_2191,In_2764,In_1207);
xor U2192 (N_2192,In_432,In_967);
xnor U2193 (N_2193,In_1786,In_489);
xnor U2194 (N_2194,In_191,In_1991);
and U2195 (N_2195,In_2930,In_1472);
and U2196 (N_2196,In_2640,In_206);
nand U2197 (N_2197,In_1629,In_1893);
nor U2198 (N_2198,In_2249,In_2715);
or U2199 (N_2199,In_1352,In_1405);
nor U2200 (N_2200,In_2695,In_1516);
nand U2201 (N_2201,In_1013,In_990);
xor U2202 (N_2202,In_698,In_1086);
nor U2203 (N_2203,In_2271,In_449);
xor U2204 (N_2204,In_344,In_196);
and U2205 (N_2205,In_2242,In_416);
nor U2206 (N_2206,In_1475,In_763);
or U2207 (N_2207,In_1609,In_2477);
nand U2208 (N_2208,In_2673,In_25);
nand U2209 (N_2209,In_1970,In_491);
or U2210 (N_2210,In_2855,In_1349);
nand U2211 (N_2211,In_1058,In_468);
nor U2212 (N_2212,In_714,In_1482);
or U2213 (N_2213,In_1074,In_1371);
nor U2214 (N_2214,In_350,In_2861);
and U2215 (N_2215,In_1358,In_72);
and U2216 (N_2216,In_679,In_2236);
or U2217 (N_2217,In_2288,In_2622);
nor U2218 (N_2218,In_1699,In_554);
nor U2219 (N_2219,In_4,In_206);
nand U2220 (N_2220,In_1761,In_677);
nand U2221 (N_2221,In_464,In_623);
or U2222 (N_2222,In_995,In_2445);
nand U2223 (N_2223,In_1028,In_1237);
and U2224 (N_2224,In_731,In_2858);
nand U2225 (N_2225,In_1556,In_1047);
xnor U2226 (N_2226,In_1563,In_38);
xnor U2227 (N_2227,In_108,In_602);
nand U2228 (N_2228,In_2209,In_958);
nor U2229 (N_2229,In_646,In_1115);
nor U2230 (N_2230,In_524,In_247);
or U2231 (N_2231,In_368,In_1749);
and U2232 (N_2232,In_1472,In_1853);
nand U2233 (N_2233,In_305,In_905);
xnor U2234 (N_2234,In_612,In_228);
nand U2235 (N_2235,In_2748,In_1037);
nor U2236 (N_2236,In_2079,In_222);
nor U2237 (N_2237,In_1228,In_1362);
nand U2238 (N_2238,In_2327,In_2044);
and U2239 (N_2239,In_2962,In_502);
nand U2240 (N_2240,In_1825,In_1044);
nand U2241 (N_2241,In_371,In_1468);
or U2242 (N_2242,In_129,In_2826);
nand U2243 (N_2243,In_1226,In_2917);
nor U2244 (N_2244,In_181,In_471);
or U2245 (N_2245,In_2635,In_1780);
and U2246 (N_2246,In_2379,In_1560);
nand U2247 (N_2247,In_2920,In_2331);
nor U2248 (N_2248,In_1869,In_2300);
or U2249 (N_2249,In_2530,In_2839);
xnor U2250 (N_2250,In_1416,In_1227);
and U2251 (N_2251,In_2051,In_1923);
nand U2252 (N_2252,In_248,In_2706);
and U2253 (N_2253,In_1403,In_1048);
nand U2254 (N_2254,In_2130,In_2008);
xor U2255 (N_2255,In_2689,In_1468);
nor U2256 (N_2256,In_2866,In_1507);
and U2257 (N_2257,In_1597,In_2173);
xor U2258 (N_2258,In_331,In_589);
nand U2259 (N_2259,In_1955,In_2548);
or U2260 (N_2260,In_795,In_313);
nand U2261 (N_2261,In_436,In_2073);
nor U2262 (N_2262,In_365,In_902);
nor U2263 (N_2263,In_229,In_2842);
nand U2264 (N_2264,In_245,In_1840);
nor U2265 (N_2265,In_492,In_2290);
nand U2266 (N_2266,In_317,In_1326);
xor U2267 (N_2267,In_1215,In_1563);
or U2268 (N_2268,In_2185,In_452);
nand U2269 (N_2269,In_1300,In_1971);
or U2270 (N_2270,In_2344,In_2899);
or U2271 (N_2271,In_1238,In_1031);
nand U2272 (N_2272,In_2713,In_1935);
nor U2273 (N_2273,In_2020,In_2976);
xnor U2274 (N_2274,In_796,In_1978);
or U2275 (N_2275,In_2643,In_1569);
or U2276 (N_2276,In_541,In_1635);
nor U2277 (N_2277,In_1177,In_2997);
xor U2278 (N_2278,In_763,In_1016);
or U2279 (N_2279,In_382,In_2057);
or U2280 (N_2280,In_2662,In_74);
xor U2281 (N_2281,In_2696,In_1043);
nand U2282 (N_2282,In_2431,In_2799);
nand U2283 (N_2283,In_1036,In_171);
nand U2284 (N_2284,In_2184,In_1112);
nand U2285 (N_2285,In_2765,In_80);
xnor U2286 (N_2286,In_2764,In_114);
and U2287 (N_2287,In_2036,In_2374);
xnor U2288 (N_2288,In_680,In_2893);
nor U2289 (N_2289,In_2755,In_1012);
and U2290 (N_2290,In_1795,In_2027);
and U2291 (N_2291,In_2112,In_1201);
or U2292 (N_2292,In_747,In_488);
xor U2293 (N_2293,In_82,In_881);
xnor U2294 (N_2294,In_1477,In_1762);
or U2295 (N_2295,In_2555,In_1192);
and U2296 (N_2296,In_348,In_1661);
and U2297 (N_2297,In_1315,In_2812);
nand U2298 (N_2298,In_51,In_1418);
nor U2299 (N_2299,In_2901,In_963);
nand U2300 (N_2300,In_1027,In_2599);
nor U2301 (N_2301,In_2998,In_1703);
or U2302 (N_2302,In_2193,In_2720);
nor U2303 (N_2303,In_582,In_2805);
and U2304 (N_2304,In_471,In_1496);
nor U2305 (N_2305,In_204,In_837);
and U2306 (N_2306,In_1657,In_842);
nor U2307 (N_2307,In_1857,In_1035);
and U2308 (N_2308,In_1729,In_521);
nand U2309 (N_2309,In_2187,In_2306);
xor U2310 (N_2310,In_2617,In_2223);
nand U2311 (N_2311,In_595,In_1452);
nand U2312 (N_2312,In_963,In_178);
nor U2313 (N_2313,In_1520,In_1475);
or U2314 (N_2314,In_943,In_1136);
nand U2315 (N_2315,In_596,In_458);
and U2316 (N_2316,In_365,In_455);
and U2317 (N_2317,In_2590,In_2145);
nor U2318 (N_2318,In_341,In_1187);
nand U2319 (N_2319,In_663,In_1968);
and U2320 (N_2320,In_1670,In_2078);
and U2321 (N_2321,In_227,In_1364);
nor U2322 (N_2322,In_2111,In_488);
and U2323 (N_2323,In_627,In_722);
nor U2324 (N_2324,In_2995,In_2741);
nor U2325 (N_2325,In_1000,In_934);
xor U2326 (N_2326,In_2760,In_881);
or U2327 (N_2327,In_1596,In_491);
or U2328 (N_2328,In_2963,In_903);
and U2329 (N_2329,In_963,In_875);
nand U2330 (N_2330,In_1314,In_300);
nand U2331 (N_2331,In_1925,In_564);
or U2332 (N_2332,In_2423,In_1022);
nor U2333 (N_2333,In_2531,In_2283);
nor U2334 (N_2334,In_1548,In_1033);
xnor U2335 (N_2335,In_710,In_1615);
and U2336 (N_2336,In_2502,In_1498);
nor U2337 (N_2337,In_1965,In_791);
or U2338 (N_2338,In_188,In_1019);
or U2339 (N_2339,In_2670,In_1607);
or U2340 (N_2340,In_1880,In_1893);
or U2341 (N_2341,In_1295,In_137);
nor U2342 (N_2342,In_846,In_2062);
xor U2343 (N_2343,In_2703,In_2666);
nand U2344 (N_2344,In_2995,In_440);
nor U2345 (N_2345,In_2187,In_2703);
and U2346 (N_2346,In_2004,In_2727);
nand U2347 (N_2347,In_624,In_45);
and U2348 (N_2348,In_2607,In_923);
and U2349 (N_2349,In_1712,In_377);
xor U2350 (N_2350,In_2630,In_2077);
xnor U2351 (N_2351,In_1144,In_904);
nor U2352 (N_2352,In_750,In_2645);
or U2353 (N_2353,In_1300,In_846);
xnor U2354 (N_2354,In_389,In_86);
and U2355 (N_2355,In_2063,In_1051);
nand U2356 (N_2356,In_2848,In_1730);
nor U2357 (N_2357,In_1519,In_2434);
nand U2358 (N_2358,In_2334,In_2779);
nor U2359 (N_2359,In_1724,In_461);
xor U2360 (N_2360,In_2240,In_1381);
and U2361 (N_2361,In_119,In_2041);
nor U2362 (N_2362,In_2522,In_2400);
xor U2363 (N_2363,In_1142,In_2484);
or U2364 (N_2364,In_2483,In_1882);
nand U2365 (N_2365,In_1812,In_1272);
and U2366 (N_2366,In_286,In_182);
nor U2367 (N_2367,In_1758,In_2949);
or U2368 (N_2368,In_158,In_37);
nor U2369 (N_2369,In_1425,In_1009);
and U2370 (N_2370,In_1546,In_2343);
nor U2371 (N_2371,In_1182,In_1318);
nand U2372 (N_2372,In_1959,In_6);
nand U2373 (N_2373,In_1353,In_359);
or U2374 (N_2374,In_1810,In_65);
or U2375 (N_2375,In_883,In_2641);
or U2376 (N_2376,In_1300,In_326);
or U2377 (N_2377,In_2887,In_1778);
and U2378 (N_2378,In_2970,In_1783);
or U2379 (N_2379,In_1944,In_2628);
nor U2380 (N_2380,In_396,In_2845);
xor U2381 (N_2381,In_2974,In_2021);
nand U2382 (N_2382,In_1251,In_2893);
or U2383 (N_2383,In_1605,In_280);
xnor U2384 (N_2384,In_1364,In_2370);
xnor U2385 (N_2385,In_2723,In_1852);
and U2386 (N_2386,In_2158,In_1736);
and U2387 (N_2387,In_328,In_2994);
xor U2388 (N_2388,In_127,In_2634);
and U2389 (N_2389,In_2812,In_1746);
nor U2390 (N_2390,In_1004,In_2733);
or U2391 (N_2391,In_1716,In_1850);
nand U2392 (N_2392,In_1909,In_1850);
nand U2393 (N_2393,In_2900,In_1876);
nor U2394 (N_2394,In_2631,In_2966);
nand U2395 (N_2395,In_2855,In_1899);
nand U2396 (N_2396,In_1500,In_1129);
xor U2397 (N_2397,In_2670,In_89);
and U2398 (N_2398,In_1525,In_585);
or U2399 (N_2399,In_1738,In_1929);
nor U2400 (N_2400,In_2352,In_124);
and U2401 (N_2401,In_1238,In_976);
xnor U2402 (N_2402,In_2876,In_299);
nand U2403 (N_2403,In_1995,In_1120);
or U2404 (N_2404,In_446,In_858);
xor U2405 (N_2405,In_491,In_443);
and U2406 (N_2406,In_105,In_2008);
and U2407 (N_2407,In_1819,In_2477);
nor U2408 (N_2408,In_1883,In_1629);
and U2409 (N_2409,In_2816,In_325);
and U2410 (N_2410,In_1375,In_1996);
nand U2411 (N_2411,In_1312,In_1801);
or U2412 (N_2412,In_2418,In_2058);
and U2413 (N_2413,In_1286,In_2840);
nand U2414 (N_2414,In_1336,In_2671);
and U2415 (N_2415,In_1514,In_1796);
xnor U2416 (N_2416,In_1139,In_654);
nand U2417 (N_2417,In_2360,In_2660);
nor U2418 (N_2418,In_1825,In_816);
xnor U2419 (N_2419,In_1707,In_461);
and U2420 (N_2420,In_1935,In_2894);
or U2421 (N_2421,In_2036,In_2853);
nor U2422 (N_2422,In_2385,In_1404);
and U2423 (N_2423,In_1736,In_1511);
xor U2424 (N_2424,In_2496,In_632);
and U2425 (N_2425,In_635,In_141);
nand U2426 (N_2426,In_1631,In_1176);
nand U2427 (N_2427,In_158,In_2113);
and U2428 (N_2428,In_2266,In_1984);
xnor U2429 (N_2429,In_2288,In_1795);
nor U2430 (N_2430,In_2216,In_1609);
nor U2431 (N_2431,In_571,In_2766);
nor U2432 (N_2432,In_1814,In_1878);
xnor U2433 (N_2433,In_1957,In_666);
nand U2434 (N_2434,In_993,In_2677);
or U2435 (N_2435,In_516,In_409);
nand U2436 (N_2436,In_2699,In_2264);
or U2437 (N_2437,In_2281,In_412);
and U2438 (N_2438,In_1433,In_1369);
nand U2439 (N_2439,In_1243,In_1012);
or U2440 (N_2440,In_592,In_190);
or U2441 (N_2441,In_2235,In_1868);
xor U2442 (N_2442,In_1614,In_2131);
or U2443 (N_2443,In_2600,In_501);
or U2444 (N_2444,In_2294,In_2636);
and U2445 (N_2445,In_1217,In_994);
nor U2446 (N_2446,In_323,In_1587);
and U2447 (N_2447,In_1452,In_2431);
or U2448 (N_2448,In_1611,In_2292);
nor U2449 (N_2449,In_1049,In_1849);
or U2450 (N_2450,In_316,In_1633);
nor U2451 (N_2451,In_422,In_2375);
and U2452 (N_2452,In_2165,In_589);
nand U2453 (N_2453,In_911,In_2527);
and U2454 (N_2454,In_2560,In_486);
xor U2455 (N_2455,In_2655,In_1215);
and U2456 (N_2456,In_2184,In_2072);
nor U2457 (N_2457,In_481,In_461);
nor U2458 (N_2458,In_208,In_497);
or U2459 (N_2459,In_1523,In_1011);
or U2460 (N_2460,In_998,In_526);
or U2461 (N_2461,In_1160,In_4);
nor U2462 (N_2462,In_2476,In_1051);
xnor U2463 (N_2463,In_2518,In_2798);
nand U2464 (N_2464,In_1227,In_1788);
nor U2465 (N_2465,In_2510,In_2894);
nand U2466 (N_2466,In_2161,In_1851);
xor U2467 (N_2467,In_942,In_2397);
xor U2468 (N_2468,In_730,In_228);
nand U2469 (N_2469,In_2660,In_2762);
or U2470 (N_2470,In_2628,In_1138);
and U2471 (N_2471,In_1225,In_2);
xor U2472 (N_2472,In_695,In_2862);
and U2473 (N_2473,In_2117,In_2779);
nand U2474 (N_2474,In_1121,In_1997);
and U2475 (N_2475,In_2971,In_153);
or U2476 (N_2476,In_1072,In_2930);
xor U2477 (N_2477,In_25,In_2106);
xnor U2478 (N_2478,In_442,In_19);
xnor U2479 (N_2479,In_918,In_2835);
and U2480 (N_2480,In_1233,In_1474);
xor U2481 (N_2481,In_678,In_2011);
nor U2482 (N_2482,In_2927,In_1913);
nor U2483 (N_2483,In_557,In_1493);
and U2484 (N_2484,In_591,In_1897);
nand U2485 (N_2485,In_1417,In_2156);
or U2486 (N_2486,In_2462,In_1708);
or U2487 (N_2487,In_1225,In_952);
nand U2488 (N_2488,In_787,In_341);
nor U2489 (N_2489,In_147,In_252);
or U2490 (N_2490,In_447,In_2916);
or U2491 (N_2491,In_2875,In_1264);
xnor U2492 (N_2492,In_1702,In_1719);
or U2493 (N_2493,In_911,In_2787);
or U2494 (N_2494,In_2946,In_1987);
xnor U2495 (N_2495,In_1934,In_1623);
xnor U2496 (N_2496,In_2160,In_845);
or U2497 (N_2497,In_2384,In_1163);
and U2498 (N_2498,In_1403,In_1527);
nand U2499 (N_2499,In_1196,In_1519);
and U2500 (N_2500,In_2404,In_719);
or U2501 (N_2501,In_680,In_264);
or U2502 (N_2502,In_240,In_1157);
or U2503 (N_2503,In_909,In_1949);
and U2504 (N_2504,In_2896,In_659);
nand U2505 (N_2505,In_765,In_546);
nand U2506 (N_2506,In_413,In_2733);
and U2507 (N_2507,In_108,In_2811);
or U2508 (N_2508,In_1001,In_1102);
xnor U2509 (N_2509,In_2270,In_2261);
or U2510 (N_2510,In_2120,In_963);
and U2511 (N_2511,In_210,In_980);
nor U2512 (N_2512,In_2120,In_1030);
or U2513 (N_2513,In_638,In_2361);
nor U2514 (N_2514,In_2610,In_2392);
nor U2515 (N_2515,In_2203,In_1480);
or U2516 (N_2516,In_2511,In_2770);
nand U2517 (N_2517,In_2718,In_328);
nor U2518 (N_2518,In_2437,In_2483);
or U2519 (N_2519,In_1313,In_304);
or U2520 (N_2520,In_2072,In_612);
nor U2521 (N_2521,In_2226,In_2244);
nor U2522 (N_2522,In_1840,In_1342);
nand U2523 (N_2523,In_1411,In_2910);
and U2524 (N_2524,In_1868,In_660);
and U2525 (N_2525,In_2157,In_1385);
nand U2526 (N_2526,In_1470,In_368);
xnor U2527 (N_2527,In_559,In_1184);
and U2528 (N_2528,In_1261,In_2991);
nor U2529 (N_2529,In_1463,In_2118);
and U2530 (N_2530,In_1678,In_1581);
or U2531 (N_2531,In_2796,In_948);
or U2532 (N_2532,In_1067,In_2606);
and U2533 (N_2533,In_616,In_1402);
nor U2534 (N_2534,In_2136,In_1258);
or U2535 (N_2535,In_1899,In_1103);
nand U2536 (N_2536,In_1043,In_1736);
xor U2537 (N_2537,In_2483,In_2324);
and U2538 (N_2538,In_2312,In_101);
or U2539 (N_2539,In_2546,In_1013);
and U2540 (N_2540,In_1975,In_2899);
xnor U2541 (N_2541,In_1803,In_1566);
nor U2542 (N_2542,In_2838,In_2525);
nor U2543 (N_2543,In_1827,In_1741);
nor U2544 (N_2544,In_1101,In_1327);
nor U2545 (N_2545,In_1921,In_1957);
or U2546 (N_2546,In_1249,In_1264);
and U2547 (N_2547,In_2488,In_2905);
and U2548 (N_2548,In_1428,In_459);
or U2549 (N_2549,In_1732,In_1512);
xnor U2550 (N_2550,In_2158,In_2876);
xnor U2551 (N_2551,In_1676,In_2089);
and U2552 (N_2552,In_1596,In_1593);
nor U2553 (N_2553,In_2340,In_2658);
or U2554 (N_2554,In_2590,In_1143);
and U2555 (N_2555,In_2848,In_944);
nor U2556 (N_2556,In_804,In_937);
nor U2557 (N_2557,In_1800,In_2980);
or U2558 (N_2558,In_342,In_301);
xnor U2559 (N_2559,In_1819,In_1148);
or U2560 (N_2560,In_917,In_2081);
or U2561 (N_2561,In_340,In_2383);
nand U2562 (N_2562,In_1131,In_1545);
xnor U2563 (N_2563,In_1301,In_758);
and U2564 (N_2564,In_2764,In_532);
or U2565 (N_2565,In_181,In_2419);
xor U2566 (N_2566,In_2475,In_628);
nand U2567 (N_2567,In_236,In_2048);
nand U2568 (N_2568,In_2371,In_1194);
nor U2569 (N_2569,In_715,In_893);
xor U2570 (N_2570,In_2437,In_1085);
or U2571 (N_2571,In_291,In_2025);
nor U2572 (N_2572,In_1631,In_104);
and U2573 (N_2573,In_1435,In_2716);
and U2574 (N_2574,In_555,In_2824);
nand U2575 (N_2575,In_2261,In_1126);
and U2576 (N_2576,In_606,In_1036);
nand U2577 (N_2577,In_1137,In_777);
xor U2578 (N_2578,In_162,In_361);
nand U2579 (N_2579,In_2341,In_1310);
nand U2580 (N_2580,In_2545,In_2392);
xor U2581 (N_2581,In_974,In_193);
xor U2582 (N_2582,In_1253,In_372);
and U2583 (N_2583,In_1649,In_2049);
xor U2584 (N_2584,In_1391,In_882);
nor U2585 (N_2585,In_1519,In_2941);
or U2586 (N_2586,In_354,In_1077);
nor U2587 (N_2587,In_405,In_243);
nor U2588 (N_2588,In_1561,In_2683);
xnor U2589 (N_2589,In_433,In_191);
nor U2590 (N_2590,In_1975,In_90);
xnor U2591 (N_2591,In_210,In_1950);
nor U2592 (N_2592,In_2976,In_1920);
nor U2593 (N_2593,In_2212,In_1041);
and U2594 (N_2594,In_1290,In_204);
nand U2595 (N_2595,In_782,In_1530);
xnor U2596 (N_2596,In_1512,In_2906);
or U2597 (N_2597,In_768,In_2713);
nand U2598 (N_2598,In_1089,In_2052);
or U2599 (N_2599,In_1261,In_1377);
xor U2600 (N_2600,In_2299,In_436);
and U2601 (N_2601,In_949,In_2415);
and U2602 (N_2602,In_1858,In_310);
nor U2603 (N_2603,In_1017,In_1686);
or U2604 (N_2604,In_321,In_2281);
or U2605 (N_2605,In_462,In_2294);
xnor U2606 (N_2606,In_2224,In_2079);
and U2607 (N_2607,In_2883,In_1268);
and U2608 (N_2608,In_2512,In_2243);
xnor U2609 (N_2609,In_2811,In_1894);
nand U2610 (N_2610,In_1561,In_2937);
nor U2611 (N_2611,In_1924,In_1646);
nand U2612 (N_2612,In_1946,In_2124);
and U2613 (N_2613,In_2273,In_2082);
xnor U2614 (N_2614,In_265,In_2789);
or U2615 (N_2615,In_527,In_1066);
and U2616 (N_2616,In_1997,In_1865);
nor U2617 (N_2617,In_52,In_1381);
and U2618 (N_2618,In_774,In_2948);
and U2619 (N_2619,In_789,In_794);
or U2620 (N_2620,In_1267,In_1294);
and U2621 (N_2621,In_2870,In_1410);
or U2622 (N_2622,In_2534,In_542);
nor U2623 (N_2623,In_1577,In_566);
or U2624 (N_2624,In_1065,In_2427);
nand U2625 (N_2625,In_2290,In_1462);
xnor U2626 (N_2626,In_1867,In_521);
and U2627 (N_2627,In_2282,In_675);
nand U2628 (N_2628,In_1773,In_2957);
nor U2629 (N_2629,In_311,In_960);
xor U2630 (N_2630,In_465,In_634);
nand U2631 (N_2631,In_817,In_522);
xor U2632 (N_2632,In_2574,In_1069);
and U2633 (N_2633,In_1559,In_46);
or U2634 (N_2634,In_291,In_2268);
xor U2635 (N_2635,In_1194,In_1890);
and U2636 (N_2636,In_1845,In_2741);
nand U2637 (N_2637,In_1588,In_2198);
nor U2638 (N_2638,In_2944,In_2843);
nor U2639 (N_2639,In_2232,In_1012);
or U2640 (N_2640,In_2435,In_653);
nand U2641 (N_2641,In_2753,In_1375);
nand U2642 (N_2642,In_1863,In_1182);
xnor U2643 (N_2643,In_2612,In_242);
or U2644 (N_2644,In_2792,In_684);
nor U2645 (N_2645,In_453,In_1718);
nand U2646 (N_2646,In_69,In_2807);
xnor U2647 (N_2647,In_1966,In_488);
xor U2648 (N_2648,In_1744,In_41);
xor U2649 (N_2649,In_1942,In_792);
nor U2650 (N_2650,In_2679,In_2522);
nor U2651 (N_2651,In_1108,In_1063);
nor U2652 (N_2652,In_1314,In_2126);
or U2653 (N_2653,In_2785,In_457);
and U2654 (N_2654,In_2618,In_736);
or U2655 (N_2655,In_2453,In_1554);
or U2656 (N_2656,In_613,In_2703);
and U2657 (N_2657,In_1049,In_1853);
xor U2658 (N_2658,In_1614,In_905);
xnor U2659 (N_2659,In_2546,In_1427);
or U2660 (N_2660,In_2008,In_721);
xnor U2661 (N_2661,In_448,In_1498);
or U2662 (N_2662,In_1617,In_227);
nor U2663 (N_2663,In_1949,In_1436);
and U2664 (N_2664,In_2932,In_872);
or U2665 (N_2665,In_2405,In_2870);
nand U2666 (N_2666,In_1640,In_290);
and U2667 (N_2667,In_2992,In_345);
nand U2668 (N_2668,In_1042,In_853);
and U2669 (N_2669,In_867,In_160);
and U2670 (N_2670,In_831,In_2751);
and U2671 (N_2671,In_1235,In_1146);
or U2672 (N_2672,In_1479,In_1702);
nor U2673 (N_2673,In_1603,In_452);
or U2674 (N_2674,In_1306,In_51);
and U2675 (N_2675,In_608,In_2934);
nor U2676 (N_2676,In_412,In_1975);
xor U2677 (N_2677,In_2784,In_2885);
and U2678 (N_2678,In_1239,In_1027);
or U2679 (N_2679,In_2963,In_2813);
xor U2680 (N_2680,In_1486,In_2659);
nand U2681 (N_2681,In_2836,In_917);
xor U2682 (N_2682,In_1257,In_1271);
nand U2683 (N_2683,In_832,In_307);
or U2684 (N_2684,In_768,In_24);
nor U2685 (N_2685,In_615,In_603);
or U2686 (N_2686,In_1434,In_2371);
nand U2687 (N_2687,In_744,In_1086);
and U2688 (N_2688,In_1259,In_324);
or U2689 (N_2689,In_737,In_1062);
nor U2690 (N_2690,In_1153,In_664);
xnor U2691 (N_2691,In_1713,In_2322);
xor U2692 (N_2692,In_1213,In_2654);
nor U2693 (N_2693,In_2703,In_1479);
xor U2694 (N_2694,In_2767,In_457);
and U2695 (N_2695,In_1496,In_2991);
and U2696 (N_2696,In_1143,In_2033);
or U2697 (N_2697,In_2213,In_1861);
or U2698 (N_2698,In_1860,In_977);
nor U2699 (N_2699,In_2447,In_312);
and U2700 (N_2700,In_728,In_1606);
and U2701 (N_2701,In_1435,In_1542);
nand U2702 (N_2702,In_584,In_1491);
xnor U2703 (N_2703,In_2219,In_164);
or U2704 (N_2704,In_302,In_1573);
or U2705 (N_2705,In_2634,In_2929);
nand U2706 (N_2706,In_2833,In_903);
nand U2707 (N_2707,In_1732,In_1605);
nor U2708 (N_2708,In_2593,In_959);
or U2709 (N_2709,In_2876,In_1155);
and U2710 (N_2710,In_1390,In_2089);
xor U2711 (N_2711,In_560,In_348);
nor U2712 (N_2712,In_447,In_2209);
and U2713 (N_2713,In_2938,In_2257);
nor U2714 (N_2714,In_2442,In_350);
nor U2715 (N_2715,In_1312,In_2847);
xnor U2716 (N_2716,In_1726,In_236);
nor U2717 (N_2717,In_2478,In_1276);
and U2718 (N_2718,In_564,In_1013);
xor U2719 (N_2719,In_701,In_386);
and U2720 (N_2720,In_214,In_133);
or U2721 (N_2721,In_2937,In_2748);
or U2722 (N_2722,In_1078,In_319);
and U2723 (N_2723,In_2663,In_2922);
nor U2724 (N_2724,In_2012,In_1661);
nor U2725 (N_2725,In_1560,In_1235);
nor U2726 (N_2726,In_2917,In_1611);
nand U2727 (N_2727,In_665,In_1422);
and U2728 (N_2728,In_781,In_1469);
nor U2729 (N_2729,In_2169,In_2923);
or U2730 (N_2730,In_1275,In_795);
nand U2731 (N_2731,In_1044,In_1141);
or U2732 (N_2732,In_2482,In_1018);
and U2733 (N_2733,In_1404,In_1148);
or U2734 (N_2734,In_630,In_1550);
nor U2735 (N_2735,In_2272,In_824);
xnor U2736 (N_2736,In_2498,In_1951);
xor U2737 (N_2737,In_874,In_2837);
nor U2738 (N_2738,In_515,In_1029);
xnor U2739 (N_2739,In_1387,In_1568);
nor U2740 (N_2740,In_1502,In_1943);
or U2741 (N_2741,In_2273,In_1328);
xor U2742 (N_2742,In_788,In_1799);
or U2743 (N_2743,In_2701,In_1035);
nor U2744 (N_2744,In_1390,In_1309);
or U2745 (N_2745,In_379,In_1680);
nand U2746 (N_2746,In_86,In_2539);
xnor U2747 (N_2747,In_2735,In_150);
nand U2748 (N_2748,In_2739,In_1232);
and U2749 (N_2749,In_2994,In_1422);
and U2750 (N_2750,In_1862,In_376);
nor U2751 (N_2751,In_924,In_1895);
xor U2752 (N_2752,In_396,In_167);
nor U2753 (N_2753,In_2520,In_2028);
nor U2754 (N_2754,In_2145,In_1817);
nor U2755 (N_2755,In_2587,In_460);
nor U2756 (N_2756,In_2520,In_359);
and U2757 (N_2757,In_1467,In_1655);
nand U2758 (N_2758,In_1219,In_2314);
or U2759 (N_2759,In_148,In_1995);
nand U2760 (N_2760,In_604,In_979);
or U2761 (N_2761,In_454,In_1162);
and U2762 (N_2762,In_2721,In_2134);
and U2763 (N_2763,In_1720,In_981);
xnor U2764 (N_2764,In_2054,In_1302);
nor U2765 (N_2765,In_1042,In_767);
nand U2766 (N_2766,In_2439,In_706);
nand U2767 (N_2767,In_83,In_2698);
nor U2768 (N_2768,In_476,In_1856);
xnor U2769 (N_2769,In_2317,In_1632);
xnor U2770 (N_2770,In_2185,In_2974);
and U2771 (N_2771,In_2371,In_2552);
or U2772 (N_2772,In_364,In_2275);
or U2773 (N_2773,In_743,In_1816);
and U2774 (N_2774,In_507,In_410);
and U2775 (N_2775,In_1407,In_1610);
nand U2776 (N_2776,In_958,In_449);
nor U2777 (N_2777,In_2681,In_876);
nor U2778 (N_2778,In_1503,In_1405);
xor U2779 (N_2779,In_719,In_416);
or U2780 (N_2780,In_1377,In_2723);
or U2781 (N_2781,In_1230,In_1761);
nand U2782 (N_2782,In_7,In_852);
and U2783 (N_2783,In_584,In_370);
or U2784 (N_2784,In_550,In_2873);
nand U2785 (N_2785,In_1297,In_1514);
nor U2786 (N_2786,In_1105,In_438);
nor U2787 (N_2787,In_2010,In_871);
xor U2788 (N_2788,In_1524,In_2725);
nor U2789 (N_2789,In_480,In_1387);
and U2790 (N_2790,In_848,In_2707);
and U2791 (N_2791,In_1980,In_1185);
xor U2792 (N_2792,In_1652,In_943);
xnor U2793 (N_2793,In_2914,In_2117);
xnor U2794 (N_2794,In_2654,In_1551);
nor U2795 (N_2795,In_1753,In_602);
and U2796 (N_2796,In_2272,In_1745);
and U2797 (N_2797,In_736,In_1254);
or U2798 (N_2798,In_2296,In_381);
or U2799 (N_2799,In_1256,In_2520);
and U2800 (N_2800,In_1261,In_1103);
or U2801 (N_2801,In_1994,In_1701);
and U2802 (N_2802,In_2044,In_555);
or U2803 (N_2803,In_2572,In_2920);
nand U2804 (N_2804,In_2024,In_1676);
xor U2805 (N_2805,In_2884,In_1447);
or U2806 (N_2806,In_2387,In_2143);
nor U2807 (N_2807,In_1700,In_2106);
nand U2808 (N_2808,In_1904,In_2275);
xnor U2809 (N_2809,In_1838,In_2514);
nor U2810 (N_2810,In_2236,In_2799);
nand U2811 (N_2811,In_2390,In_198);
or U2812 (N_2812,In_1850,In_2096);
xnor U2813 (N_2813,In_155,In_700);
nor U2814 (N_2814,In_399,In_255);
xor U2815 (N_2815,In_1903,In_1328);
nand U2816 (N_2816,In_2249,In_2409);
or U2817 (N_2817,In_1132,In_1677);
xnor U2818 (N_2818,In_1784,In_116);
nand U2819 (N_2819,In_1090,In_658);
or U2820 (N_2820,In_2583,In_746);
and U2821 (N_2821,In_1024,In_786);
nand U2822 (N_2822,In_2376,In_1483);
nor U2823 (N_2823,In_2887,In_252);
and U2824 (N_2824,In_1556,In_2797);
xnor U2825 (N_2825,In_1541,In_1315);
nand U2826 (N_2826,In_1605,In_194);
or U2827 (N_2827,In_1023,In_1400);
nor U2828 (N_2828,In_9,In_230);
nor U2829 (N_2829,In_2021,In_1260);
and U2830 (N_2830,In_872,In_948);
nor U2831 (N_2831,In_2080,In_2533);
nor U2832 (N_2832,In_1510,In_2847);
nor U2833 (N_2833,In_2466,In_399);
xor U2834 (N_2834,In_1989,In_1446);
or U2835 (N_2835,In_2186,In_1691);
xnor U2836 (N_2836,In_104,In_591);
xnor U2837 (N_2837,In_749,In_1288);
nor U2838 (N_2838,In_2526,In_1379);
nand U2839 (N_2839,In_2931,In_2901);
xnor U2840 (N_2840,In_688,In_2622);
nor U2841 (N_2841,In_783,In_1593);
nand U2842 (N_2842,In_1666,In_1985);
or U2843 (N_2843,In_1973,In_309);
or U2844 (N_2844,In_545,In_201);
nand U2845 (N_2845,In_2517,In_327);
and U2846 (N_2846,In_1943,In_1333);
nor U2847 (N_2847,In_874,In_2247);
nor U2848 (N_2848,In_816,In_834);
or U2849 (N_2849,In_2417,In_1007);
nand U2850 (N_2850,In_955,In_1925);
and U2851 (N_2851,In_307,In_347);
and U2852 (N_2852,In_2134,In_2217);
xor U2853 (N_2853,In_652,In_658);
and U2854 (N_2854,In_2656,In_577);
and U2855 (N_2855,In_738,In_172);
and U2856 (N_2856,In_2880,In_2650);
nor U2857 (N_2857,In_548,In_2413);
or U2858 (N_2858,In_617,In_645);
nor U2859 (N_2859,In_1313,In_1613);
and U2860 (N_2860,In_2229,In_2761);
nor U2861 (N_2861,In_567,In_156);
nand U2862 (N_2862,In_2934,In_847);
nand U2863 (N_2863,In_1580,In_1859);
nor U2864 (N_2864,In_2751,In_749);
xor U2865 (N_2865,In_1505,In_1022);
or U2866 (N_2866,In_1078,In_2279);
nor U2867 (N_2867,In_2512,In_763);
or U2868 (N_2868,In_560,In_2708);
nand U2869 (N_2869,In_618,In_2180);
xor U2870 (N_2870,In_351,In_190);
nor U2871 (N_2871,In_786,In_2438);
xnor U2872 (N_2872,In_924,In_1161);
xnor U2873 (N_2873,In_235,In_1261);
nor U2874 (N_2874,In_717,In_918);
or U2875 (N_2875,In_155,In_706);
nand U2876 (N_2876,In_2422,In_2406);
and U2877 (N_2877,In_1492,In_127);
xor U2878 (N_2878,In_1952,In_2906);
or U2879 (N_2879,In_824,In_2387);
or U2880 (N_2880,In_1553,In_2320);
nand U2881 (N_2881,In_387,In_641);
and U2882 (N_2882,In_138,In_1052);
or U2883 (N_2883,In_712,In_733);
and U2884 (N_2884,In_587,In_2292);
and U2885 (N_2885,In_175,In_1655);
xnor U2886 (N_2886,In_2473,In_603);
nand U2887 (N_2887,In_2034,In_2333);
or U2888 (N_2888,In_2804,In_1854);
xnor U2889 (N_2889,In_2360,In_2435);
or U2890 (N_2890,In_1757,In_1446);
or U2891 (N_2891,In_1870,In_2109);
nand U2892 (N_2892,In_307,In_2483);
nor U2893 (N_2893,In_124,In_58);
xnor U2894 (N_2894,In_1744,In_771);
and U2895 (N_2895,In_1439,In_161);
xnor U2896 (N_2896,In_1362,In_2980);
xnor U2897 (N_2897,In_2783,In_108);
nand U2898 (N_2898,In_855,In_1469);
nor U2899 (N_2899,In_2869,In_849);
and U2900 (N_2900,In_1053,In_417);
and U2901 (N_2901,In_2454,In_2867);
nand U2902 (N_2902,In_101,In_2719);
xor U2903 (N_2903,In_2953,In_2158);
and U2904 (N_2904,In_2210,In_1395);
xnor U2905 (N_2905,In_1336,In_2933);
nor U2906 (N_2906,In_1865,In_1347);
and U2907 (N_2907,In_1093,In_1850);
or U2908 (N_2908,In_2969,In_179);
or U2909 (N_2909,In_1377,In_1060);
or U2910 (N_2910,In_1522,In_686);
nand U2911 (N_2911,In_330,In_2436);
xor U2912 (N_2912,In_1730,In_2417);
and U2913 (N_2913,In_2796,In_2521);
nor U2914 (N_2914,In_681,In_2550);
or U2915 (N_2915,In_623,In_61);
nor U2916 (N_2916,In_1541,In_1654);
xor U2917 (N_2917,In_2610,In_1549);
nor U2918 (N_2918,In_596,In_601);
and U2919 (N_2919,In_1838,In_74);
xor U2920 (N_2920,In_526,In_881);
xor U2921 (N_2921,In_1514,In_2445);
xnor U2922 (N_2922,In_2783,In_808);
xnor U2923 (N_2923,In_306,In_961);
and U2924 (N_2924,In_280,In_1747);
and U2925 (N_2925,In_911,In_2859);
nand U2926 (N_2926,In_851,In_1992);
and U2927 (N_2927,In_1216,In_2814);
or U2928 (N_2928,In_97,In_1888);
xnor U2929 (N_2929,In_706,In_1187);
and U2930 (N_2930,In_1103,In_2115);
nor U2931 (N_2931,In_1161,In_1182);
and U2932 (N_2932,In_1335,In_2718);
nand U2933 (N_2933,In_575,In_690);
xor U2934 (N_2934,In_784,In_1727);
or U2935 (N_2935,In_1603,In_1984);
nand U2936 (N_2936,In_182,In_841);
or U2937 (N_2937,In_269,In_2572);
and U2938 (N_2938,In_2673,In_578);
nand U2939 (N_2939,In_236,In_660);
nor U2940 (N_2940,In_783,In_1097);
nand U2941 (N_2941,In_250,In_1642);
nand U2942 (N_2942,In_2178,In_2227);
or U2943 (N_2943,In_2889,In_2044);
or U2944 (N_2944,In_1283,In_411);
nor U2945 (N_2945,In_1101,In_981);
xor U2946 (N_2946,In_516,In_219);
nor U2947 (N_2947,In_660,In_1677);
nor U2948 (N_2948,In_246,In_1314);
nor U2949 (N_2949,In_0,In_2770);
or U2950 (N_2950,In_1650,In_36);
and U2951 (N_2951,In_2056,In_1372);
and U2952 (N_2952,In_2598,In_1186);
or U2953 (N_2953,In_1884,In_868);
xor U2954 (N_2954,In_54,In_1125);
nand U2955 (N_2955,In_2492,In_381);
and U2956 (N_2956,In_1977,In_1886);
or U2957 (N_2957,In_1841,In_928);
nor U2958 (N_2958,In_228,In_2603);
or U2959 (N_2959,In_1790,In_399);
and U2960 (N_2960,In_246,In_513);
nand U2961 (N_2961,In_821,In_1178);
nand U2962 (N_2962,In_2066,In_27);
xor U2963 (N_2963,In_1201,In_2111);
xor U2964 (N_2964,In_1320,In_1375);
xor U2965 (N_2965,In_2227,In_670);
nor U2966 (N_2966,In_2167,In_2054);
or U2967 (N_2967,In_2040,In_1678);
and U2968 (N_2968,In_2837,In_2404);
nor U2969 (N_2969,In_2481,In_2431);
nor U2970 (N_2970,In_77,In_253);
xnor U2971 (N_2971,In_543,In_1134);
and U2972 (N_2972,In_2469,In_1120);
or U2973 (N_2973,In_974,In_192);
nand U2974 (N_2974,In_1959,In_1516);
xor U2975 (N_2975,In_211,In_2293);
or U2976 (N_2976,In_2461,In_2583);
nand U2977 (N_2977,In_1602,In_1847);
and U2978 (N_2978,In_2552,In_1925);
nor U2979 (N_2979,In_1734,In_1986);
nor U2980 (N_2980,In_2657,In_129);
nor U2981 (N_2981,In_2711,In_2722);
nand U2982 (N_2982,In_2987,In_2645);
nand U2983 (N_2983,In_2769,In_496);
or U2984 (N_2984,In_649,In_1477);
and U2985 (N_2985,In_2188,In_1133);
and U2986 (N_2986,In_928,In_2875);
nor U2987 (N_2987,In_2995,In_2730);
xor U2988 (N_2988,In_2976,In_386);
and U2989 (N_2989,In_1779,In_765);
and U2990 (N_2990,In_1708,In_1138);
nor U2991 (N_2991,In_2224,In_2070);
or U2992 (N_2992,In_818,In_61);
and U2993 (N_2993,In_2574,In_1735);
nor U2994 (N_2994,In_1752,In_879);
and U2995 (N_2995,In_2294,In_662);
nand U2996 (N_2996,In_697,In_741);
nand U2997 (N_2997,In_1732,In_1490);
xor U2998 (N_2998,In_2975,In_1893);
and U2999 (N_2999,In_1593,In_2931);
nor U3000 (N_3000,In_2804,In_486);
or U3001 (N_3001,In_1352,In_1897);
or U3002 (N_3002,In_1668,In_722);
or U3003 (N_3003,In_773,In_268);
nand U3004 (N_3004,In_512,In_193);
or U3005 (N_3005,In_746,In_469);
nor U3006 (N_3006,In_194,In_2423);
nand U3007 (N_3007,In_590,In_2883);
nand U3008 (N_3008,In_1270,In_1777);
nand U3009 (N_3009,In_619,In_2778);
nand U3010 (N_3010,In_1993,In_1540);
nor U3011 (N_3011,In_2004,In_1049);
or U3012 (N_3012,In_2686,In_57);
and U3013 (N_3013,In_2126,In_808);
nand U3014 (N_3014,In_2800,In_865);
and U3015 (N_3015,In_2446,In_1897);
xor U3016 (N_3016,In_181,In_2445);
or U3017 (N_3017,In_1150,In_2363);
xor U3018 (N_3018,In_487,In_2967);
xor U3019 (N_3019,In_2500,In_2901);
or U3020 (N_3020,In_2090,In_2589);
nor U3021 (N_3021,In_2768,In_1317);
nand U3022 (N_3022,In_2850,In_1090);
nand U3023 (N_3023,In_1480,In_2575);
nor U3024 (N_3024,In_1330,In_2825);
or U3025 (N_3025,In_1316,In_1765);
xor U3026 (N_3026,In_2832,In_1009);
or U3027 (N_3027,In_1714,In_2578);
nor U3028 (N_3028,In_919,In_1491);
nand U3029 (N_3029,In_1860,In_587);
and U3030 (N_3030,In_2392,In_2872);
xor U3031 (N_3031,In_1135,In_672);
or U3032 (N_3032,In_2017,In_589);
or U3033 (N_3033,In_140,In_2260);
or U3034 (N_3034,In_2158,In_1677);
or U3035 (N_3035,In_1773,In_2586);
nand U3036 (N_3036,In_2160,In_2007);
nor U3037 (N_3037,In_2033,In_2456);
nand U3038 (N_3038,In_2862,In_1010);
xnor U3039 (N_3039,In_1796,In_805);
nor U3040 (N_3040,In_1454,In_2021);
xnor U3041 (N_3041,In_2552,In_1529);
and U3042 (N_3042,In_2336,In_1743);
nor U3043 (N_3043,In_2434,In_2719);
and U3044 (N_3044,In_1703,In_2512);
or U3045 (N_3045,In_2212,In_2713);
nor U3046 (N_3046,In_2990,In_1533);
nand U3047 (N_3047,In_2910,In_1033);
and U3048 (N_3048,In_1740,In_2553);
nor U3049 (N_3049,In_797,In_1809);
nor U3050 (N_3050,In_754,In_1341);
xnor U3051 (N_3051,In_2799,In_1175);
xnor U3052 (N_3052,In_1561,In_1438);
nand U3053 (N_3053,In_2526,In_1074);
and U3054 (N_3054,In_2142,In_1686);
and U3055 (N_3055,In_2404,In_128);
xor U3056 (N_3056,In_2626,In_2495);
nand U3057 (N_3057,In_2662,In_1026);
nand U3058 (N_3058,In_1634,In_2596);
or U3059 (N_3059,In_1977,In_1056);
nand U3060 (N_3060,In_1289,In_1964);
or U3061 (N_3061,In_2887,In_2595);
and U3062 (N_3062,In_542,In_511);
nor U3063 (N_3063,In_668,In_1886);
or U3064 (N_3064,In_2460,In_1536);
and U3065 (N_3065,In_2081,In_530);
or U3066 (N_3066,In_136,In_682);
nand U3067 (N_3067,In_287,In_1808);
or U3068 (N_3068,In_493,In_1721);
or U3069 (N_3069,In_1297,In_701);
or U3070 (N_3070,In_1106,In_2136);
nand U3071 (N_3071,In_2813,In_374);
and U3072 (N_3072,In_352,In_2138);
xor U3073 (N_3073,In_788,In_151);
xnor U3074 (N_3074,In_1746,In_1863);
and U3075 (N_3075,In_861,In_1765);
nand U3076 (N_3076,In_2015,In_1608);
nor U3077 (N_3077,In_2050,In_2374);
nor U3078 (N_3078,In_1774,In_1816);
and U3079 (N_3079,In_2466,In_1681);
and U3080 (N_3080,In_1387,In_4);
and U3081 (N_3081,In_985,In_60);
xnor U3082 (N_3082,In_2091,In_891);
nor U3083 (N_3083,In_1958,In_2610);
and U3084 (N_3084,In_2636,In_2789);
nor U3085 (N_3085,In_2705,In_2581);
xnor U3086 (N_3086,In_742,In_443);
xor U3087 (N_3087,In_552,In_2718);
xnor U3088 (N_3088,In_2031,In_1829);
or U3089 (N_3089,In_1244,In_2054);
nand U3090 (N_3090,In_851,In_2126);
nand U3091 (N_3091,In_1695,In_1703);
nand U3092 (N_3092,In_446,In_2228);
or U3093 (N_3093,In_2353,In_1579);
xnor U3094 (N_3094,In_156,In_2297);
or U3095 (N_3095,In_2518,In_2806);
or U3096 (N_3096,In_2883,In_982);
xnor U3097 (N_3097,In_680,In_455);
nand U3098 (N_3098,In_2661,In_2702);
or U3099 (N_3099,In_2694,In_1259);
nor U3100 (N_3100,In_1872,In_2799);
xor U3101 (N_3101,In_689,In_2963);
and U3102 (N_3102,In_2783,In_2439);
nand U3103 (N_3103,In_855,In_2326);
and U3104 (N_3104,In_514,In_1140);
xnor U3105 (N_3105,In_702,In_2214);
and U3106 (N_3106,In_615,In_2974);
or U3107 (N_3107,In_1578,In_2180);
nand U3108 (N_3108,In_626,In_2326);
nand U3109 (N_3109,In_2072,In_1729);
or U3110 (N_3110,In_2147,In_614);
nor U3111 (N_3111,In_476,In_2682);
nand U3112 (N_3112,In_474,In_2515);
nor U3113 (N_3113,In_2204,In_1047);
nor U3114 (N_3114,In_560,In_878);
and U3115 (N_3115,In_1349,In_1630);
or U3116 (N_3116,In_1909,In_1496);
xnor U3117 (N_3117,In_2293,In_1827);
and U3118 (N_3118,In_1300,In_1105);
nand U3119 (N_3119,In_328,In_661);
xnor U3120 (N_3120,In_232,In_307);
and U3121 (N_3121,In_938,In_2079);
nor U3122 (N_3122,In_1539,In_2619);
nand U3123 (N_3123,In_1099,In_1292);
and U3124 (N_3124,In_2040,In_2297);
nand U3125 (N_3125,In_1611,In_1372);
or U3126 (N_3126,In_2775,In_2628);
or U3127 (N_3127,In_2403,In_2208);
or U3128 (N_3128,In_2536,In_205);
or U3129 (N_3129,In_2326,In_585);
and U3130 (N_3130,In_1532,In_2898);
nand U3131 (N_3131,In_256,In_597);
nand U3132 (N_3132,In_938,In_36);
xnor U3133 (N_3133,In_2996,In_28);
xnor U3134 (N_3134,In_1361,In_1926);
nor U3135 (N_3135,In_531,In_889);
and U3136 (N_3136,In_450,In_1228);
xor U3137 (N_3137,In_1971,In_1874);
nand U3138 (N_3138,In_2055,In_211);
nand U3139 (N_3139,In_255,In_256);
nand U3140 (N_3140,In_2348,In_101);
or U3141 (N_3141,In_2650,In_1808);
xor U3142 (N_3142,In_712,In_947);
nor U3143 (N_3143,In_1754,In_758);
nand U3144 (N_3144,In_2575,In_674);
and U3145 (N_3145,In_69,In_2486);
nand U3146 (N_3146,In_2472,In_1205);
or U3147 (N_3147,In_2068,In_388);
xnor U3148 (N_3148,In_2295,In_2173);
or U3149 (N_3149,In_847,In_2809);
xor U3150 (N_3150,In_2307,In_2601);
and U3151 (N_3151,In_516,In_1624);
nand U3152 (N_3152,In_27,In_1774);
xnor U3153 (N_3153,In_791,In_1779);
nand U3154 (N_3154,In_1332,In_322);
nand U3155 (N_3155,In_1845,In_1457);
xnor U3156 (N_3156,In_431,In_1680);
nand U3157 (N_3157,In_2740,In_1922);
or U3158 (N_3158,In_1277,In_164);
nand U3159 (N_3159,In_1243,In_1014);
nand U3160 (N_3160,In_291,In_2598);
or U3161 (N_3161,In_1896,In_2056);
xor U3162 (N_3162,In_1086,In_2430);
or U3163 (N_3163,In_2313,In_440);
nor U3164 (N_3164,In_565,In_592);
or U3165 (N_3165,In_1071,In_657);
or U3166 (N_3166,In_2978,In_1192);
nor U3167 (N_3167,In_123,In_2918);
nand U3168 (N_3168,In_544,In_2330);
and U3169 (N_3169,In_165,In_2361);
nor U3170 (N_3170,In_2019,In_758);
and U3171 (N_3171,In_114,In_602);
and U3172 (N_3172,In_2852,In_1417);
or U3173 (N_3173,In_2434,In_2548);
nor U3174 (N_3174,In_1720,In_2629);
nand U3175 (N_3175,In_841,In_23);
xnor U3176 (N_3176,In_2094,In_737);
nand U3177 (N_3177,In_241,In_2483);
nand U3178 (N_3178,In_1038,In_2512);
nand U3179 (N_3179,In_91,In_2883);
nand U3180 (N_3180,In_2696,In_1316);
or U3181 (N_3181,In_600,In_1117);
nand U3182 (N_3182,In_2124,In_1762);
and U3183 (N_3183,In_491,In_266);
xor U3184 (N_3184,In_256,In_2359);
xnor U3185 (N_3185,In_482,In_1137);
nand U3186 (N_3186,In_2580,In_449);
nor U3187 (N_3187,In_2124,In_1688);
or U3188 (N_3188,In_1549,In_993);
and U3189 (N_3189,In_700,In_610);
nand U3190 (N_3190,In_544,In_2639);
nor U3191 (N_3191,In_1871,In_27);
and U3192 (N_3192,In_1526,In_2611);
or U3193 (N_3193,In_2338,In_239);
xor U3194 (N_3194,In_1894,In_2960);
xnor U3195 (N_3195,In_953,In_1644);
and U3196 (N_3196,In_1253,In_2551);
and U3197 (N_3197,In_2142,In_2743);
and U3198 (N_3198,In_949,In_2248);
nor U3199 (N_3199,In_2572,In_568);
and U3200 (N_3200,In_1296,In_880);
or U3201 (N_3201,In_2334,In_699);
xnor U3202 (N_3202,In_2033,In_680);
or U3203 (N_3203,In_437,In_2386);
and U3204 (N_3204,In_2257,In_1632);
or U3205 (N_3205,In_1828,In_1607);
xor U3206 (N_3206,In_2767,In_1864);
or U3207 (N_3207,In_2143,In_2838);
nand U3208 (N_3208,In_1319,In_2684);
xor U3209 (N_3209,In_1659,In_1662);
nand U3210 (N_3210,In_800,In_2193);
or U3211 (N_3211,In_451,In_26);
or U3212 (N_3212,In_471,In_2690);
nor U3213 (N_3213,In_1553,In_660);
xnor U3214 (N_3214,In_2422,In_281);
nor U3215 (N_3215,In_2046,In_614);
and U3216 (N_3216,In_806,In_703);
or U3217 (N_3217,In_1990,In_2865);
nor U3218 (N_3218,In_79,In_737);
and U3219 (N_3219,In_1304,In_523);
nor U3220 (N_3220,In_902,In_144);
or U3221 (N_3221,In_1987,In_1081);
and U3222 (N_3222,In_2922,In_265);
xor U3223 (N_3223,In_1022,In_878);
and U3224 (N_3224,In_1666,In_2322);
nor U3225 (N_3225,In_686,In_181);
xor U3226 (N_3226,In_2893,In_979);
xnor U3227 (N_3227,In_2643,In_1202);
and U3228 (N_3228,In_2926,In_2570);
and U3229 (N_3229,In_1790,In_2772);
xnor U3230 (N_3230,In_1228,In_2581);
and U3231 (N_3231,In_254,In_1596);
and U3232 (N_3232,In_2040,In_2952);
nor U3233 (N_3233,In_2541,In_2186);
or U3234 (N_3234,In_103,In_2490);
nand U3235 (N_3235,In_561,In_383);
xnor U3236 (N_3236,In_1555,In_1849);
or U3237 (N_3237,In_385,In_2422);
nand U3238 (N_3238,In_264,In_786);
or U3239 (N_3239,In_83,In_835);
xor U3240 (N_3240,In_686,In_1016);
or U3241 (N_3241,In_1536,In_2878);
nand U3242 (N_3242,In_2710,In_1472);
nor U3243 (N_3243,In_2892,In_356);
or U3244 (N_3244,In_2252,In_2181);
or U3245 (N_3245,In_328,In_1741);
xor U3246 (N_3246,In_413,In_2354);
or U3247 (N_3247,In_2030,In_1857);
or U3248 (N_3248,In_792,In_1600);
nor U3249 (N_3249,In_1748,In_707);
and U3250 (N_3250,In_1133,In_184);
nand U3251 (N_3251,In_2230,In_1722);
nor U3252 (N_3252,In_2074,In_2078);
xor U3253 (N_3253,In_1819,In_1203);
nor U3254 (N_3254,In_458,In_2829);
and U3255 (N_3255,In_303,In_1629);
xor U3256 (N_3256,In_275,In_1757);
or U3257 (N_3257,In_1723,In_1859);
and U3258 (N_3258,In_202,In_1608);
or U3259 (N_3259,In_958,In_2994);
xor U3260 (N_3260,In_1890,In_2981);
nand U3261 (N_3261,In_262,In_2623);
nand U3262 (N_3262,In_65,In_12);
xnor U3263 (N_3263,In_842,In_1391);
xor U3264 (N_3264,In_1199,In_1932);
nand U3265 (N_3265,In_1397,In_481);
nand U3266 (N_3266,In_296,In_151);
nor U3267 (N_3267,In_2689,In_2350);
nor U3268 (N_3268,In_2109,In_1588);
or U3269 (N_3269,In_80,In_591);
nand U3270 (N_3270,In_1492,In_2516);
nand U3271 (N_3271,In_493,In_2777);
or U3272 (N_3272,In_2511,In_628);
xor U3273 (N_3273,In_293,In_2633);
nand U3274 (N_3274,In_1094,In_1280);
nand U3275 (N_3275,In_2007,In_728);
or U3276 (N_3276,In_2507,In_1326);
nand U3277 (N_3277,In_327,In_2228);
nor U3278 (N_3278,In_2904,In_790);
or U3279 (N_3279,In_1669,In_1745);
xnor U3280 (N_3280,In_272,In_1618);
and U3281 (N_3281,In_1035,In_2356);
xor U3282 (N_3282,In_1046,In_2034);
xnor U3283 (N_3283,In_1002,In_2009);
or U3284 (N_3284,In_697,In_1745);
or U3285 (N_3285,In_1,In_1174);
xnor U3286 (N_3286,In_2953,In_8);
nand U3287 (N_3287,In_645,In_23);
nand U3288 (N_3288,In_1411,In_1240);
nand U3289 (N_3289,In_1760,In_1074);
nor U3290 (N_3290,In_2118,In_2216);
xnor U3291 (N_3291,In_767,In_156);
or U3292 (N_3292,In_1607,In_1753);
or U3293 (N_3293,In_1764,In_2054);
xor U3294 (N_3294,In_934,In_1267);
xor U3295 (N_3295,In_1111,In_130);
and U3296 (N_3296,In_644,In_375);
nand U3297 (N_3297,In_351,In_2962);
nor U3298 (N_3298,In_69,In_19);
or U3299 (N_3299,In_1452,In_709);
xnor U3300 (N_3300,In_1601,In_1913);
nor U3301 (N_3301,In_131,In_1534);
and U3302 (N_3302,In_2817,In_1236);
nand U3303 (N_3303,In_1727,In_586);
nand U3304 (N_3304,In_1749,In_1294);
xor U3305 (N_3305,In_2925,In_2670);
and U3306 (N_3306,In_2771,In_2686);
and U3307 (N_3307,In_2296,In_1075);
nand U3308 (N_3308,In_1185,In_1420);
and U3309 (N_3309,In_1756,In_2492);
xnor U3310 (N_3310,In_2547,In_2228);
nor U3311 (N_3311,In_392,In_2227);
nor U3312 (N_3312,In_431,In_1670);
nor U3313 (N_3313,In_2045,In_1542);
and U3314 (N_3314,In_1756,In_10);
xor U3315 (N_3315,In_1576,In_342);
nand U3316 (N_3316,In_2335,In_853);
or U3317 (N_3317,In_2345,In_411);
and U3318 (N_3318,In_2309,In_2130);
nand U3319 (N_3319,In_1815,In_1517);
or U3320 (N_3320,In_2028,In_1091);
xor U3321 (N_3321,In_1163,In_175);
nand U3322 (N_3322,In_1355,In_1490);
nand U3323 (N_3323,In_2461,In_1282);
and U3324 (N_3324,In_2643,In_614);
nor U3325 (N_3325,In_1549,In_492);
xor U3326 (N_3326,In_2697,In_1971);
or U3327 (N_3327,In_2558,In_782);
or U3328 (N_3328,In_1311,In_2469);
or U3329 (N_3329,In_2423,In_738);
nand U3330 (N_3330,In_1176,In_799);
nand U3331 (N_3331,In_201,In_1140);
nor U3332 (N_3332,In_1694,In_1229);
and U3333 (N_3333,In_1179,In_777);
or U3334 (N_3334,In_2212,In_2169);
xor U3335 (N_3335,In_1074,In_1629);
xor U3336 (N_3336,In_883,In_2484);
nand U3337 (N_3337,In_2522,In_2052);
xnor U3338 (N_3338,In_2649,In_2609);
or U3339 (N_3339,In_2214,In_832);
or U3340 (N_3340,In_1794,In_2884);
or U3341 (N_3341,In_2258,In_1988);
and U3342 (N_3342,In_1053,In_832);
or U3343 (N_3343,In_2020,In_295);
xor U3344 (N_3344,In_2977,In_2287);
xnor U3345 (N_3345,In_1345,In_1956);
xnor U3346 (N_3346,In_1075,In_2589);
xnor U3347 (N_3347,In_622,In_273);
xnor U3348 (N_3348,In_1127,In_2172);
xor U3349 (N_3349,In_189,In_590);
xnor U3350 (N_3350,In_351,In_2048);
or U3351 (N_3351,In_2974,In_2564);
or U3352 (N_3352,In_816,In_1129);
nand U3353 (N_3353,In_2762,In_2411);
and U3354 (N_3354,In_1667,In_299);
and U3355 (N_3355,In_1012,In_2879);
nand U3356 (N_3356,In_2438,In_1211);
nor U3357 (N_3357,In_98,In_55);
xnor U3358 (N_3358,In_1205,In_1324);
nand U3359 (N_3359,In_1797,In_2740);
and U3360 (N_3360,In_707,In_586);
xnor U3361 (N_3361,In_2184,In_1698);
or U3362 (N_3362,In_259,In_2163);
or U3363 (N_3363,In_2061,In_2564);
and U3364 (N_3364,In_2507,In_1047);
nand U3365 (N_3365,In_678,In_2775);
and U3366 (N_3366,In_1727,In_964);
xor U3367 (N_3367,In_2967,In_548);
nand U3368 (N_3368,In_1216,In_1996);
nor U3369 (N_3369,In_1356,In_1343);
nor U3370 (N_3370,In_814,In_2900);
xnor U3371 (N_3371,In_1165,In_429);
or U3372 (N_3372,In_712,In_1295);
nand U3373 (N_3373,In_586,In_1395);
xor U3374 (N_3374,In_2445,In_1342);
nor U3375 (N_3375,In_1414,In_1172);
nand U3376 (N_3376,In_2125,In_2181);
or U3377 (N_3377,In_2669,In_784);
nand U3378 (N_3378,In_1745,In_1002);
nor U3379 (N_3379,In_2524,In_2336);
nand U3380 (N_3380,In_2813,In_1497);
nor U3381 (N_3381,In_2165,In_15);
or U3382 (N_3382,In_2737,In_454);
and U3383 (N_3383,In_2128,In_2473);
nand U3384 (N_3384,In_656,In_35);
and U3385 (N_3385,In_1628,In_2170);
xnor U3386 (N_3386,In_1765,In_1374);
and U3387 (N_3387,In_106,In_1041);
xor U3388 (N_3388,In_1399,In_2426);
nand U3389 (N_3389,In_1439,In_913);
and U3390 (N_3390,In_738,In_1552);
and U3391 (N_3391,In_2193,In_1735);
nand U3392 (N_3392,In_2299,In_2315);
or U3393 (N_3393,In_1647,In_2336);
nor U3394 (N_3394,In_1054,In_2793);
nor U3395 (N_3395,In_1534,In_1770);
nand U3396 (N_3396,In_990,In_1165);
and U3397 (N_3397,In_1651,In_862);
nor U3398 (N_3398,In_1247,In_2572);
xor U3399 (N_3399,In_410,In_643);
nand U3400 (N_3400,In_651,In_1103);
xor U3401 (N_3401,In_1141,In_1431);
and U3402 (N_3402,In_1134,In_2846);
xor U3403 (N_3403,In_276,In_1659);
nand U3404 (N_3404,In_2176,In_2771);
and U3405 (N_3405,In_2676,In_311);
nor U3406 (N_3406,In_798,In_2090);
xor U3407 (N_3407,In_2526,In_1278);
or U3408 (N_3408,In_2481,In_1262);
nand U3409 (N_3409,In_2213,In_40);
xor U3410 (N_3410,In_2767,In_430);
xor U3411 (N_3411,In_495,In_2782);
and U3412 (N_3412,In_2810,In_2058);
nor U3413 (N_3413,In_2305,In_2418);
nand U3414 (N_3414,In_534,In_2208);
nor U3415 (N_3415,In_485,In_2282);
and U3416 (N_3416,In_1039,In_946);
xnor U3417 (N_3417,In_2870,In_1477);
xor U3418 (N_3418,In_2590,In_1841);
nor U3419 (N_3419,In_371,In_2147);
nor U3420 (N_3420,In_1818,In_121);
nor U3421 (N_3421,In_2975,In_1070);
and U3422 (N_3422,In_2913,In_2518);
xnor U3423 (N_3423,In_2571,In_217);
nor U3424 (N_3424,In_263,In_2295);
nor U3425 (N_3425,In_2783,In_2366);
nor U3426 (N_3426,In_116,In_1291);
nand U3427 (N_3427,In_928,In_1598);
and U3428 (N_3428,In_2689,In_2427);
and U3429 (N_3429,In_1734,In_1847);
nor U3430 (N_3430,In_1778,In_1690);
or U3431 (N_3431,In_2372,In_2236);
or U3432 (N_3432,In_2875,In_1652);
or U3433 (N_3433,In_936,In_286);
nor U3434 (N_3434,In_998,In_1298);
and U3435 (N_3435,In_2499,In_1057);
or U3436 (N_3436,In_2753,In_1408);
or U3437 (N_3437,In_576,In_381);
xnor U3438 (N_3438,In_1714,In_526);
or U3439 (N_3439,In_547,In_1185);
xor U3440 (N_3440,In_2624,In_1970);
and U3441 (N_3441,In_1004,In_1094);
nand U3442 (N_3442,In_255,In_889);
xnor U3443 (N_3443,In_458,In_634);
nand U3444 (N_3444,In_236,In_2045);
xnor U3445 (N_3445,In_2946,In_959);
nand U3446 (N_3446,In_1312,In_1821);
xnor U3447 (N_3447,In_1973,In_1791);
nand U3448 (N_3448,In_1877,In_86);
and U3449 (N_3449,In_2936,In_1434);
or U3450 (N_3450,In_1346,In_262);
nand U3451 (N_3451,In_1695,In_2198);
nor U3452 (N_3452,In_2061,In_133);
xor U3453 (N_3453,In_646,In_2241);
nor U3454 (N_3454,In_2993,In_2238);
or U3455 (N_3455,In_1429,In_244);
nor U3456 (N_3456,In_756,In_1710);
and U3457 (N_3457,In_2694,In_621);
and U3458 (N_3458,In_1098,In_2388);
or U3459 (N_3459,In_1130,In_515);
xnor U3460 (N_3460,In_1385,In_903);
or U3461 (N_3461,In_1972,In_2966);
or U3462 (N_3462,In_1265,In_1253);
and U3463 (N_3463,In_2762,In_1569);
and U3464 (N_3464,In_323,In_1061);
nand U3465 (N_3465,In_2045,In_613);
nor U3466 (N_3466,In_2481,In_2459);
xnor U3467 (N_3467,In_1797,In_726);
xnor U3468 (N_3468,In_2959,In_2364);
or U3469 (N_3469,In_1694,In_2086);
and U3470 (N_3470,In_242,In_654);
xnor U3471 (N_3471,In_1383,In_180);
xnor U3472 (N_3472,In_1521,In_989);
and U3473 (N_3473,In_1165,In_2414);
nor U3474 (N_3474,In_1790,In_1472);
and U3475 (N_3475,In_2236,In_92);
nor U3476 (N_3476,In_858,In_1850);
or U3477 (N_3477,In_2166,In_2253);
nand U3478 (N_3478,In_1114,In_1537);
xor U3479 (N_3479,In_52,In_2096);
or U3480 (N_3480,In_425,In_2772);
or U3481 (N_3481,In_1502,In_2955);
or U3482 (N_3482,In_236,In_1554);
nor U3483 (N_3483,In_1137,In_789);
nand U3484 (N_3484,In_2147,In_2139);
nand U3485 (N_3485,In_2724,In_1408);
and U3486 (N_3486,In_2750,In_68);
and U3487 (N_3487,In_369,In_2994);
xor U3488 (N_3488,In_943,In_992);
xor U3489 (N_3489,In_2989,In_1585);
nand U3490 (N_3490,In_900,In_2240);
or U3491 (N_3491,In_2090,In_1312);
xnor U3492 (N_3492,In_2077,In_1890);
nor U3493 (N_3493,In_221,In_2562);
xnor U3494 (N_3494,In_2609,In_2986);
nand U3495 (N_3495,In_2151,In_880);
nand U3496 (N_3496,In_1114,In_2610);
or U3497 (N_3497,In_2224,In_220);
nand U3498 (N_3498,In_2123,In_2154);
nor U3499 (N_3499,In_1833,In_1675);
nand U3500 (N_3500,In_1689,In_649);
nor U3501 (N_3501,In_26,In_141);
xor U3502 (N_3502,In_689,In_2829);
or U3503 (N_3503,In_1446,In_1689);
xnor U3504 (N_3504,In_1939,In_1682);
and U3505 (N_3505,In_2507,In_2003);
nor U3506 (N_3506,In_2612,In_1080);
nand U3507 (N_3507,In_471,In_86);
and U3508 (N_3508,In_2919,In_1431);
xor U3509 (N_3509,In_857,In_754);
and U3510 (N_3510,In_2957,In_2032);
nor U3511 (N_3511,In_2607,In_2981);
and U3512 (N_3512,In_2010,In_1976);
nand U3513 (N_3513,In_1660,In_1074);
or U3514 (N_3514,In_2781,In_2613);
nor U3515 (N_3515,In_1149,In_2292);
nor U3516 (N_3516,In_219,In_2770);
nor U3517 (N_3517,In_1081,In_143);
nand U3518 (N_3518,In_2850,In_2626);
nor U3519 (N_3519,In_1899,In_2667);
nand U3520 (N_3520,In_767,In_160);
nor U3521 (N_3521,In_2979,In_1553);
xor U3522 (N_3522,In_2258,In_673);
nand U3523 (N_3523,In_2710,In_1930);
nor U3524 (N_3524,In_48,In_2558);
nor U3525 (N_3525,In_721,In_669);
nor U3526 (N_3526,In_266,In_1310);
or U3527 (N_3527,In_1131,In_838);
and U3528 (N_3528,In_655,In_255);
nor U3529 (N_3529,In_1307,In_2129);
and U3530 (N_3530,In_2031,In_67);
nor U3531 (N_3531,In_204,In_1936);
xor U3532 (N_3532,In_2027,In_742);
nor U3533 (N_3533,In_1631,In_1551);
xnor U3534 (N_3534,In_514,In_2901);
nor U3535 (N_3535,In_2753,In_1625);
nand U3536 (N_3536,In_421,In_2882);
nor U3537 (N_3537,In_2348,In_2619);
xor U3538 (N_3538,In_722,In_110);
or U3539 (N_3539,In_1268,In_1231);
xnor U3540 (N_3540,In_1203,In_1004);
nand U3541 (N_3541,In_2930,In_2308);
nor U3542 (N_3542,In_1662,In_1950);
or U3543 (N_3543,In_65,In_1932);
xor U3544 (N_3544,In_606,In_655);
nand U3545 (N_3545,In_1257,In_2013);
or U3546 (N_3546,In_1106,In_2236);
nand U3547 (N_3547,In_1150,In_585);
or U3548 (N_3548,In_1435,In_1714);
and U3549 (N_3549,In_1835,In_2970);
nor U3550 (N_3550,In_1022,In_2761);
and U3551 (N_3551,In_1427,In_2382);
or U3552 (N_3552,In_1381,In_34);
nor U3553 (N_3553,In_2116,In_761);
nor U3554 (N_3554,In_1066,In_2796);
nor U3555 (N_3555,In_735,In_36);
xor U3556 (N_3556,In_2827,In_1743);
and U3557 (N_3557,In_660,In_426);
and U3558 (N_3558,In_1330,In_1485);
xnor U3559 (N_3559,In_2840,In_2387);
nand U3560 (N_3560,In_1979,In_1534);
xnor U3561 (N_3561,In_673,In_2330);
or U3562 (N_3562,In_1936,In_1013);
or U3563 (N_3563,In_2361,In_316);
xnor U3564 (N_3564,In_2576,In_912);
or U3565 (N_3565,In_759,In_2675);
nor U3566 (N_3566,In_808,In_983);
nor U3567 (N_3567,In_1382,In_2255);
nand U3568 (N_3568,In_2706,In_504);
or U3569 (N_3569,In_965,In_2455);
or U3570 (N_3570,In_1644,In_343);
nor U3571 (N_3571,In_1943,In_1560);
and U3572 (N_3572,In_395,In_522);
or U3573 (N_3573,In_2913,In_946);
nor U3574 (N_3574,In_152,In_631);
nor U3575 (N_3575,In_2087,In_2054);
nor U3576 (N_3576,In_2294,In_2101);
or U3577 (N_3577,In_180,In_851);
and U3578 (N_3578,In_2669,In_93);
nand U3579 (N_3579,In_1888,In_2239);
xor U3580 (N_3580,In_1606,In_1207);
and U3581 (N_3581,In_1093,In_2201);
and U3582 (N_3582,In_248,In_2765);
and U3583 (N_3583,In_698,In_1331);
nor U3584 (N_3584,In_562,In_2691);
xnor U3585 (N_3585,In_614,In_2155);
and U3586 (N_3586,In_1568,In_2788);
and U3587 (N_3587,In_1433,In_1685);
nor U3588 (N_3588,In_936,In_429);
xor U3589 (N_3589,In_840,In_117);
and U3590 (N_3590,In_567,In_2594);
nor U3591 (N_3591,In_1102,In_1508);
nand U3592 (N_3592,In_947,In_1001);
or U3593 (N_3593,In_1112,In_2648);
nor U3594 (N_3594,In_502,In_1999);
xor U3595 (N_3595,In_2790,In_1138);
and U3596 (N_3596,In_2436,In_1270);
or U3597 (N_3597,In_1136,In_967);
xnor U3598 (N_3598,In_302,In_2846);
xor U3599 (N_3599,In_1630,In_2491);
and U3600 (N_3600,In_836,In_953);
nand U3601 (N_3601,In_2708,In_1873);
nor U3602 (N_3602,In_2616,In_2657);
nand U3603 (N_3603,In_2840,In_2874);
nand U3604 (N_3604,In_1984,In_1285);
xor U3605 (N_3605,In_47,In_2204);
nor U3606 (N_3606,In_1375,In_2953);
xor U3607 (N_3607,In_2724,In_954);
xor U3608 (N_3608,In_296,In_2433);
nand U3609 (N_3609,In_2153,In_1656);
nand U3610 (N_3610,In_2038,In_1671);
or U3611 (N_3611,In_195,In_1833);
xnor U3612 (N_3612,In_54,In_1477);
and U3613 (N_3613,In_1674,In_661);
or U3614 (N_3614,In_2527,In_1108);
xor U3615 (N_3615,In_755,In_2029);
nand U3616 (N_3616,In_1140,In_2294);
and U3617 (N_3617,In_210,In_412);
nand U3618 (N_3618,In_312,In_225);
xnor U3619 (N_3619,In_1765,In_692);
xor U3620 (N_3620,In_1223,In_639);
nor U3621 (N_3621,In_1769,In_2341);
xnor U3622 (N_3622,In_2432,In_1238);
and U3623 (N_3623,In_2210,In_1113);
nor U3624 (N_3624,In_1970,In_157);
and U3625 (N_3625,In_1871,In_1446);
nor U3626 (N_3626,In_2406,In_2411);
nand U3627 (N_3627,In_2815,In_2378);
xor U3628 (N_3628,In_2294,In_1638);
nor U3629 (N_3629,In_2179,In_1885);
and U3630 (N_3630,In_2975,In_1080);
nor U3631 (N_3631,In_1150,In_2554);
and U3632 (N_3632,In_1109,In_289);
nand U3633 (N_3633,In_2783,In_2900);
and U3634 (N_3634,In_1446,In_2225);
or U3635 (N_3635,In_173,In_2147);
and U3636 (N_3636,In_2322,In_2105);
nor U3637 (N_3637,In_1154,In_242);
and U3638 (N_3638,In_1870,In_335);
or U3639 (N_3639,In_2850,In_1317);
nor U3640 (N_3640,In_825,In_2807);
or U3641 (N_3641,In_51,In_1823);
xor U3642 (N_3642,In_1399,In_917);
nor U3643 (N_3643,In_197,In_1446);
nor U3644 (N_3644,In_1550,In_2383);
and U3645 (N_3645,In_3,In_2434);
and U3646 (N_3646,In_177,In_857);
xor U3647 (N_3647,In_1717,In_162);
xor U3648 (N_3648,In_1228,In_753);
xnor U3649 (N_3649,In_1500,In_433);
or U3650 (N_3650,In_1184,In_2934);
nand U3651 (N_3651,In_2175,In_2846);
nor U3652 (N_3652,In_2022,In_1295);
or U3653 (N_3653,In_2307,In_2353);
xor U3654 (N_3654,In_2417,In_2580);
nand U3655 (N_3655,In_2456,In_795);
and U3656 (N_3656,In_381,In_292);
nor U3657 (N_3657,In_1602,In_266);
nand U3658 (N_3658,In_701,In_1364);
nand U3659 (N_3659,In_2837,In_2953);
nand U3660 (N_3660,In_1714,In_647);
nor U3661 (N_3661,In_376,In_2666);
and U3662 (N_3662,In_2935,In_1552);
and U3663 (N_3663,In_2573,In_537);
xnor U3664 (N_3664,In_1306,In_659);
and U3665 (N_3665,In_1022,In_1236);
or U3666 (N_3666,In_4,In_991);
nor U3667 (N_3667,In_2392,In_1891);
and U3668 (N_3668,In_1382,In_1085);
xnor U3669 (N_3669,In_708,In_580);
and U3670 (N_3670,In_2744,In_1667);
nor U3671 (N_3671,In_2073,In_758);
nor U3672 (N_3672,In_1287,In_916);
and U3673 (N_3673,In_2207,In_1714);
and U3674 (N_3674,In_2552,In_936);
xor U3675 (N_3675,In_80,In_1236);
and U3676 (N_3676,In_2207,In_994);
nor U3677 (N_3677,In_299,In_1209);
or U3678 (N_3678,In_1686,In_873);
or U3679 (N_3679,In_1615,In_1527);
nor U3680 (N_3680,In_609,In_2955);
xnor U3681 (N_3681,In_2246,In_1879);
xnor U3682 (N_3682,In_1979,In_795);
xor U3683 (N_3683,In_827,In_2026);
xnor U3684 (N_3684,In_501,In_2329);
xor U3685 (N_3685,In_2055,In_628);
or U3686 (N_3686,In_857,In_513);
or U3687 (N_3687,In_2906,In_315);
and U3688 (N_3688,In_797,In_1995);
and U3689 (N_3689,In_1717,In_268);
nor U3690 (N_3690,In_821,In_1999);
xor U3691 (N_3691,In_2829,In_1043);
or U3692 (N_3692,In_1687,In_2250);
nor U3693 (N_3693,In_1746,In_1412);
or U3694 (N_3694,In_1905,In_1076);
and U3695 (N_3695,In_2357,In_2383);
nor U3696 (N_3696,In_784,In_383);
or U3697 (N_3697,In_1508,In_2602);
xnor U3698 (N_3698,In_2515,In_2838);
and U3699 (N_3699,In_1550,In_555);
or U3700 (N_3700,In_2109,In_2300);
and U3701 (N_3701,In_111,In_1555);
nor U3702 (N_3702,In_2165,In_2596);
and U3703 (N_3703,In_2259,In_723);
xor U3704 (N_3704,In_593,In_1816);
nand U3705 (N_3705,In_1323,In_2767);
nand U3706 (N_3706,In_2914,In_2662);
xor U3707 (N_3707,In_2380,In_1607);
nand U3708 (N_3708,In_775,In_2751);
nor U3709 (N_3709,In_2827,In_2981);
or U3710 (N_3710,In_551,In_593);
nand U3711 (N_3711,In_437,In_689);
or U3712 (N_3712,In_1321,In_60);
xnor U3713 (N_3713,In_2106,In_551);
or U3714 (N_3714,In_9,In_1255);
and U3715 (N_3715,In_2021,In_2397);
or U3716 (N_3716,In_576,In_969);
and U3717 (N_3717,In_859,In_454);
nor U3718 (N_3718,In_2529,In_2153);
xnor U3719 (N_3719,In_276,In_74);
nand U3720 (N_3720,In_288,In_2136);
xor U3721 (N_3721,In_2312,In_2859);
and U3722 (N_3722,In_1740,In_1695);
xnor U3723 (N_3723,In_1430,In_1721);
nor U3724 (N_3724,In_2062,In_1830);
xnor U3725 (N_3725,In_288,In_1891);
or U3726 (N_3726,In_1475,In_1858);
nand U3727 (N_3727,In_1379,In_1310);
and U3728 (N_3728,In_910,In_2451);
nor U3729 (N_3729,In_1480,In_739);
or U3730 (N_3730,In_234,In_2556);
or U3731 (N_3731,In_198,In_401);
nand U3732 (N_3732,In_2667,In_1729);
nor U3733 (N_3733,In_1879,In_1471);
or U3734 (N_3734,In_1324,In_1657);
nor U3735 (N_3735,In_1952,In_1237);
nand U3736 (N_3736,In_2799,In_872);
and U3737 (N_3737,In_2875,In_2521);
xor U3738 (N_3738,In_2128,In_474);
nand U3739 (N_3739,In_1611,In_873);
or U3740 (N_3740,In_911,In_2474);
or U3741 (N_3741,In_1597,In_1873);
xnor U3742 (N_3742,In_731,In_2762);
or U3743 (N_3743,In_2858,In_2816);
nand U3744 (N_3744,In_1714,In_436);
or U3745 (N_3745,In_1636,In_1867);
or U3746 (N_3746,In_1985,In_786);
nand U3747 (N_3747,In_199,In_1043);
and U3748 (N_3748,In_1260,In_482);
or U3749 (N_3749,In_1806,In_64);
or U3750 (N_3750,In_436,In_2312);
nor U3751 (N_3751,In_1503,In_1582);
xor U3752 (N_3752,In_2515,In_864);
nand U3753 (N_3753,In_1594,In_1540);
nand U3754 (N_3754,In_1111,In_913);
xor U3755 (N_3755,In_506,In_122);
and U3756 (N_3756,In_1474,In_1436);
and U3757 (N_3757,In_2301,In_1822);
nand U3758 (N_3758,In_939,In_2942);
nand U3759 (N_3759,In_2949,In_1337);
and U3760 (N_3760,In_2614,In_1325);
xor U3761 (N_3761,In_507,In_1755);
nand U3762 (N_3762,In_1252,In_1386);
nor U3763 (N_3763,In_1571,In_521);
nor U3764 (N_3764,In_2489,In_2829);
xor U3765 (N_3765,In_695,In_2655);
and U3766 (N_3766,In_473,In_994);
nand U3767 (N_3767,In_1921,In_1698);
nand U3768 (N_3768,In_617,In_1012);
nor U3769 (N_3769,In_1527,In_2256);
or U3770 (N_3770,In_2385,In_377);
nor U3771 (N_3771,In_888,In_820);
nor U3772 (N_3772,In_1253,In_790);
and U3773 (N_3773,In_959,In_1435);
xor U3774 (N_3774,In_1336,In_1847);
and U3775 (N_3775,In_2130,In_1667);
nand U3776 (N_3776,In_1994,In_971);
and U3777 (N_3777,In_2940,In_1664);
nand U3778 (N_3778,In_1473,In_1285);
or U3779 (N_3779,In_382,In_2674);
and U3780 (N_3780,In_1992,In_749);
or U3781 (N_3781,In_657,In_2002);
xor U3782 (N_3782,In_2477,In_564);
xnor U3783 (N_3783,In_782,In_1613);
xnor U3784 (N_3784,In_2738,In_2972);
xor U3785 (N_3785,In_184,In_2426);
nor U3786 (N_3786,In_2086,In_2949);
and U3787 (N_3787,In_2613,In_2341);
or U3788 (N_3788,In_1965,In_2641);
nand U3789 (N_3789,In_770,In_2904);
nand U3790 (N_3790,In_651,In_1375);
nand U3791 (N_3791,In_1680,In_2189);
nand U3792 (N_3792,In_1148,In_1180);
nand U3793 (N_3793,In_2022,In_2674);
nor U3794 (N_3794,In_487,In_2694);
xnor U3795 (N_3795,In_542,In_1950);
nand U3796 (N_3796,In_168,In_2869);
nor U3797 (N_3797,In_2585,In_1548);
xor U3798 (N_3798,In_143,In_659);
and U3799 (N_3799,In_1835,In_171);
or U3800 (N_3800,In_742,In_1217);
nand U3801 (N_3801,In_196,In_1335);
xor U3802 (N_3802,In_1499,In_2663);
xor U3803 (N_3803,In_2881,In_2567);
nor U3804 (N_3804,In_2889,In_2916);
or U3805 (N_3805,In_2515,In_1142);
nor U3806 (N_3806,In_2193,In_2804);
or U3807 (N_3807,In_294,In_994);
nand U3808 (N_3808,In_2913,In_2328);
nand U3809 (N_3809,In_2074,In_2274);
nor U3810 (N_3810,In_379,In_799);
xor U3811 (N_3811,In_1603,In_1681);
nand U3812 (N_3812,In_1731,In_189);
xor U3813 (N_3813,In_1194,In_2648);
nor U3814 (N_3814,In_2619,In_1266);
or U3815 (N_3815,In_1890,In_500);
nand U3816 (N_3816,In_898,In_2652);
or U3817 (N_3817,In_1730,In_1558);
and U3818 (N_3818,In_1613,In_978);
xor U3819 (N_3819,In_943,In_1251);
or U3820 (N_3820,In_934,In_977);
nand U3821 (N_3821,In_616,In_820);
and U3822 (N_3822,In_2583,In_1920);
or U3823 (N_3823,In_574,In_810);
and U3824 (N_3824,In_658,In_1184);
or U3825 (N_3825,In_65,In_617);
nand U3826 (N_3826,In_2260,In_76);
and U3827 (N_3827,In_2058,In_903);
and U3828 (N_3828,In_2706,In_1423);
and U3829 (N_3829,In_2005,In_1051);
and U3830 (N_3830,In_75,In_2780);
nor U3831 (N_3831,In_2446,In_1686);
xnor U3832 (N_3832,In_1167,In_397);
nor U3833 (N_3833,In_1742,In_1660);
nor U3834 (N_3834,In_2829,In_846);
nor U3835 (N_3835,In_2425,In_406);
xor U3836 (N_3836,In_279,In_1965);
and U3837 (N_3837,In_2526,In_1176);
and U3838 (N_3838,In_1956,In_2923);
xor U3839 (N_3839,In_2421,In_336);
nor U3840 (N_3840,In_1637,In_1443);
or U3841 (N_3841,In_2004,In_2247);
and U3842 (N_3842,In_337,In_2761);
nand U3843 (N_3843,In_2710,In_2364);
and U3844 (N_3844,In_1575,In_2400);
or U3845 (N_3845,In_2232,In_436);
and U3846 (N_3846,In_1826,In_360);
nor U3847 (N_3847,In_2844,In_2377);
and U3848 (N_3848,In_2517,In_532);
nand U3849 (N_3849,In_1653,In_409);
or U3850 (N_3850,In_105,In_442);
or U3851 (N_3851,In_1370,In_168);
and U3852 (N_3852,In_169,In_1533);
or U3853 (N_3853,In_1027,In_2319);
and U3854 (N_3854,In_591,In_2714);
or U3855 (N_3855,In_2509,In_2061);
and U3856 (N_3856,In_1003,In_817);
or U3857 (N_3857,In_511,In_2005);
and U3858 (N_3858,In_275,In_265);
and U3859 (N_3859,In_352,In_383);
and U3860 (N_3860,In_2206,In_1954);
nor U3861 (N_3861,In_1943,In_1999);
nor U3862 (N_3862,In_1695,In_670);
and U3863 (N_3863,In_2960,In_2837);
or U3864 (N_3864,In_2277,In_1236);
and U3865 (N_3865,In_301,In_2416);
nand U3866 (N_3866,In_1994,In_1539);
nand U3867 (N_3867,In_260,In_2244);
xor U3868 (N_3868,In_772,In_596);
xnor U3869 (N_3869,In_1684,In_290);
xnor U3870 (N_3870,In_2549,In_2232);
xnor U3871 (N_3871,In_2467,In_2043);
nand U3872 (N_3872,In_638,In_2300);
nand U3873 (N_3873,In_554,In_1898);
and U3874 (N_3874,In_1200,In_2273);
nand U3875 (N_3875,In_2311,In_1150);
and U3876 (N_3876,In_760,In_1999);
or U3877 (N_3877,In_184,In_1764);
nand U3878 (N_3878,In_2090,In_2521);
nor U3879 (N_3879,In_2376,In_1462);
and U3880 (N_3880,In_1312,In_1866);
and U3881 (N_3881,In_2415,In_2701);
xnor U3882 (N_3882,In_1536,In_1219);
and U3883 (N_3883,In_832,In_642);
or U3884 (N_3884,In_383,In_2130);
or U3885 (N_3885,In_518,In_230);
and U3886 (N_3886,In_2064,In_1599);
or U3887 (N_3887,In_860,In_1607);
nor U3888 (N_3888,In_1977,In_2259);
and U3889 (N_3889,In_1087,In_2473);
or U3890 (N_3890,In_2795,In_313);
xor U3891 (N_3891,In_639,In_582);
nand U3892 (N_3892,In_2589,In_2708);
xnor U3893 (N_3893,In_2560,In_1574);
xor U3894 (N_3894,In_994,In_1987);
nand U3895 (N_3895,In_1060,In_1248);
nor U3896 (N_3896,In_1820,In_851);
nor U3897 (N_3897,In_2606,In_2375);
nand U3898 (N_3898,In_1287,In_893);
nor U3899 (N_3899,In_321,In_1896);
or U3900 (N_3900,In_635,In_2925);
nand U3901 (N_3901,In_1102,In_302);
xnor U3902 (N_3902,In_1289,In_2113);
and U3903 (N_3903,In_89,In_1868);
or U3904 (N_3904,In_563,In_934);
xnor U3905 (N_3905,In_489,In_1357);
xor U3906 (N_3906,In_1631,In_2965);
and U3907 (N_3907,In_1387,In_1142);
nand U3908 (N_3908,In_724,In_286);
xor U3909 (N_3909,In_314,In_117);
nand U3910 (N_3910,In_1936,In_2216);
and U3911 (N_3911,In_591,In_1786);
or U3912 (N_3912,In_907,In_1953);
nand U3913 (N_3913,In_1110,In_906);
nand U3914 (N_3914,In_1215,In_829);
xnor U3915 (N_3915,In_724,In_294);
or U3916 (N_3916,In_1485,In_428);
nand U3917 (N_3917,In_2007,In_2793);
xor U3918 (N_3918,In_616,In_602);
and U3919 (N_3919,In_2407,In_2812);
nand U3920 (N_3920,In_215,In_2465);
xnor U3921 (N_3921,In_1419,In_30);
or U3922 (N_3922,In_631,In_1858);
and U3923 (N_3923,In_1912,In_2230);
or U3924 (N_3924,In_1313,In_1057);
xnor U3925 (N_3925,In_1301,In_2403);
or U3926 (N_3926,In_2809,In_1460);
or U3927 (N_3927,In_1396,In_2387);
and U3928 (N_3928,In_2471,In_1854);
and U3929 (N_3929,In_502,In_50);
xor U3930 (N_3930,In_1988,In_2002);
and U3931 (N_3931,In_1766,In_2940);
nor U3932 (N_3932,In_2440,In_1893);
nand U3933 (N_3933,In_2136,In_1652);
xor U3934 (N_3934,In_2178,In_875);
nor U3935 (N_3935,In_2791,In_111);
nand U3936 (N_3936,In_1843,In_1701);
xnor U3937 (N_3937,In_1645,In_1913);
or U3938 (N_3938,In_750,In_1286);
xor U3939 (N_3939,In_1434,In_1712);
nand U3940 (N_3940,In_1066,In_1445);
or U3941 (N_3941,In_1505,In_1791);
nand U3942 (N_3942,In_1807,In_716);
or U3943 (N_3943,In_2899,In_733);
and U3944 (N_3944,In_1284,In_767);
xnor U3945 (N_3945,In_27,In_539);
and U3946 (N_3946,In_951,In_518);
nor U3947 (N_3947,In_88,In_1192);
xor U3948 (N_3948,In_916,In_1019);
nand U3949 (N_3949,In_2053,In_532);
xor U3950 (N_3950,In_574,In_680);
nand U3951 (N_3951,In_2751,In_561);
nand U3952 (N_3952,In_2930,In_1305);
xor U3953 (N_3953,In_673,In_904);
or U3954 (N_3954,In_381,In_356);
nor U3955 (N_3955,In_1922,In_2389);
nor U3956 (N_3956,In_2444,In_940);
nor U3957 (N_3957,In_1054,In_2073);
xor U3958 (N_3958,In_515,In_1187);
xnor U3959 (N_3959,In_694,In_436);
nand U3960 (N_3960,In_326,In_345);
nand U3961 (N_3961,In_2901,In_189);
xnor U3962 (N_3962,In_438,In_2042);
nand U3963 (N_3963,In_1927,In_540);
nand U3964 (N_3964,In_2896,In_1054);
nor U3965 (N_3965,In_2827,In_2510);
xnor U3966 (N_3966,In_803,In_1219);
or U3967 (N_3967,In_844,In_1012);
xnor U3968 (N_3968,In_1234,In_348);
and U3969 (N_3969,In_2144,In_2493);
nand U3970 (N_3970,In_2605,In_1376);
nand U3971 (N_3971,In_517,In_2768);
xnor U3972 (N_3972,In_1852,In_572);
nor U3973 (N_3973,In_2897,In_2026);
nand U3974 (N_3974,In_424,In_1516);
xor U3975 (N_3975,In_1014,In_209);
xor U3976 (N_3976,In_524,In_1697);
and U3977 (N_3977,In_691,In_2786);
xnor U3978 (N_3978,In_621,In_947);
nor U3979 (N_3979,In_412,In_2247);
or U3980 (N_3980,In_1501,In_694);
nor U3981 (N_3981,In_1787,In_393);
xnor U3982 (N_3982,In_172,In_631);
and U3983 (N_3983,In_590,In_2470);
nor U3984 (N_3984,In_399,In_998);
or U3985 (N_3985,In_2796,In_940);
nand U3986 (N_3986,In_827,In_1772);
or U3987 (N_3987,In_76,In_3);
and U3988 (N_3988,In_1236,In_2121);
or U3989 (N_3989,In_2534,In_946);
nor U3990 (N_3990,In_2460,In_1758);
nor U3991 (N_3991,In_2554,In_1533);
nor U3992 (N_3992,In_1639,In_1767);
nand U3993 (N_3993,In_933,In_1747);
and U3994 (N_3994,In_2096,In_2207);
and U3995 (N_3995,In_220,In_1216);
xnor U3996 (N_3996,In_1616,In_307);
xnor U3997 (N_3997,In_544,In_1944);
xnor U3998 (N_3998,In_907,In_2907);
nand U3999 (N_3999,In_2214,In_2521);
or U4000 (N_4000,In_2613,In_238);
nor U4001 (N_4001,In_2078,In_1233);
nand U4002 (N_4002,In_1227,In_825);
nor U4003 (N_4003,In_2545,In_1711);
nor U4004 (N_4004,In_2533,In_556);
nand U4005 (N_4005,In_1282,In_440);
xnor U4006 (N_4006,In_1785,In_2689);
nand U4007 (N_4007,In_1767,In_2998);
and U4008 (N_4008,In_961,In_1574);
nor U4009 (N_4009,In_1039,In_1862);
xor U4010 (N_4010,In_2209,In_1466);
or U4011 (N_4011,In_2327,In_2443);
or U4012 (N_4012,In_2329,In_1789);
and U4013 (N_4013,In_875,In_737);
nand U4014 (N_4014,In_1838,In_1910);
and U4015 (N_4015,In_1050,In_1564);
or U4016 (N_4016,In_1799,In_2605);
nand U4017 (N_4017,In_2134,In_1303);
and U4018 (N_4018,In_2755,In_1730);
xor U4019 (N_4019,In_1484,In_1281);
xor U4020 (N_4020,In_1101,In_61);
xor U4021 (N_4021,In_1106,In_2473);
or U4022 (N_4022,In_762,In_1325);
nor U4023 (N_4023,In_2810,In_2552);
or U4024 (N_4024,In_2498,In_2198);
nor U4025 (N_4025,In_2351,In_2297);
and U4026 (N_4026,In_2671,In_1932);
xor U4027 (N_4027,In_1942,In_2282);
and U4028 (N_4028,In_2564,In_1487);
xnor U4029 (N_4029,In_2852,In_2196);
and U4030 (N_4030,In_2043,In_1830);
and U4031 (N_4031,In_2960,In_1235);
or U4032 (N_4032,In_761,In_1041);
nor U4033 (N_4033,In_471,In_443);
nor U4034 (N_4034,In_1335,In_717);
or U4035 (N_4035,In_1763,In_2957);
or U4036 (N_4036,In_906,In_1548);
nor U4037 (N_4037,In_2983,In_2938);
nor U4038 (N_4038,In_1945,In_2179);
or U4039 (N_4039,In_2302,In_1865);
nand U4040 (N_4040,In_1747,In_2769);
or U4041 (N_4041,In_594,In_1052);
nor U4042 (N_4042,In_2952,In_800);
and U4043 (N_4043,In_724,In_1331);
xor U4044 (N_4044,In_1720,In_1768);
and U4045 (N_4045,In_2372,In_1465);
nor U4046 (N_4046,In_2015,In_510);
nor U4047 (N_4047,In_1461,In_2360);
xnor U4048 (N_4048,In_445,In_284);
or U4049 (N_4049,In_2679,In_936);
and U4050 (N_4050,In_2501,In_2745);
xor U4051 (N_4051,In_1163,In_2985);
nor U4052 (N_4052,In_2579,In_2321);
xor U4053 (N_4053,In_1876,In_2124);
and U4054 (N_4054,In_2613,In_1044);
xor U4055 (N_4055,In_1993,In_1550);
xor U4056 (N_4056,In_1586,In_385);
nor U4057 (N_4057,In_510,In_1310);
or U4058 (N_4058,In_2754,In_2999);
or U4059 (N_4059,In_2600,In_2258);
nand U4060 (N_4060,In_1411,In_1830);
nand U4061 (N_4061,In_955,In_2262);
and U4062 (N_4062,In_2079,In_1365);
nand U4063 (N_4063,In_1450,In_1991);
and U4064 (N_4064,In_2195,In_2549);
and U4065 (N_4065,In_1093,In_1674);
xnor U4066 (N_4066,In_2114,In_1029);
and U4067 (N_4067,In_2477,In_1659);
or U4068 (N_4068,In_2412,In_2006);
nor U4069 (N_4069,In_2566,In_2456);
nor U4070 (N_4070,In_457,In_2878);
and U4071 (N_4071,In_220,In_2041);
and U4072 (N_4072,In_2481,In_1150);
or U4073 (N_4073,In_1830,In_2496);
xnor U4074 (N_4074,In_1979,In_1508);
or U4075 (N_4075,In_2203,In_2234);
or U4076 (N_4076,In_1461,In_2261);
or U4077 (N_4077,In_1420,In_2585);
xnor U4078 (N_4078,In_2959,In_2039);
and U4079 (N_4079,In_623,In_2836);
xor U4080 (N_4080,In_2273,In_468);
or U4081 (N_4081,In_1644,In_2192);
and U4082 (N_4082,In_637,In_1356);
or U4083 (N_4083,In_1070,In_2571);
nand U4084 (N_4084,In_1735,In_2801);
or U4085 (N_4085,In_2282,In_2192);
nand U4086 (N_4086,In_2715,In_1806);
nor U4087 (N_4087,In_2477,In_2439);
and U4088 (N_4088,In_971,In_452);
xor U4089 (N_4089,In_938,In_1217);
xnor U4090 (N_4090,In_1509,In_1154);
nand U4091 (N_4091,In_2859,In_1716);
and U4092 (N_4092,In_2612,In_1229);
and U4093 (N_4093,In_2804,In_2299);
xor U4094 (N_4094,In_1119,In_1438);
nor U4095 (N_4095,In_1188,In_2892);
and U4096 (N_4096,In_1576,In_799);
or U4097 (N_4097,In_2210,In_91);
nand U4098 (N_4098,In_1451,In_399);
nor U4099 (N_4099,In_632,In_1320);
xnor U4100 (N_4100,In_78,In_30);
or U4101 (N_4101,In_1270,In_111);
and U4102 (N_4102,In_130,In_941);
nand U4103 (N_4103,In_2934,In_1867);
nor U4104 (N_4104,In_474,In_69);
nor U4105 (N_4105,In_1511,In_32);
or U4106 (N_4106,In_954,In_2174);
or U4107 (N_4107,In_2911,In_173);
or U4108 (N_4108,In_1470,In_2871);
nand U4109 (N_4109,In_2652,In_502);
nor U4110 (N_4110,In_87,In_1419);
nand U4111 (N_4111,In_2692,In_1386);
xnor U4112 (N_4112,In_2344,In_515);
nor U4113 (N_4113,In_633,In_1935);
nor U4114 (N_4114,In_2413,In_2314);
nand U4115 (N_4115,In_2004,In_1033);
nand U4116 (N_4116,In_2910,In_2879);
nor U4117 (N_4117,In_1476,In_717);
xor U4118 (N_4118,In_1943,In_761);
nand U4119 (N_4119,In_2390,In_1004);
and U4120 (N_4120,In_1857,In_1943);
and U4121 (N_4121,In_1729,In_2370);
and U4122 (N_4122,In_1365,In_1700);
and U4123 (N_4123,In_325,In_619);
or U4124 (N_4124,In_74,In_2954);
nor U4125 (N_4125,In_1399,In_2842);
nand U4126 (N_4126,In_2547,In_1397);
nor U4127 (N_4127,In_2623,In_2392);
nand U4128 (N_4128,In_2450,In_1588);
nand U4129 (N_4129,In_2415,In_504);
xor U4130 (N_4130,In_111,In_2863);
xor U4131 (N_4131,In_1302,In_930);
and U4132 (N_4132,In_451,In_82);
nor U4133 (N_4133,In_660,In_2041);
nor U4134 (N_4134,In_795,In_1098);
nand U4135 (N_4135,In_441,In_86);
xor U4136 (N_4136,In_669,In_2768);
xnor U4137 (N_4137,In_650,In_697);
or U4138 (N_4138,In_2920,In_2996);
nor U4139 (N_4139,In_2636,In_2828);
nor U4140 (N_4140,In_456,In_778);
xor U4141 (N_4141,In_805,In_516);
xor U4142 (N_4142,In_1261,In_1231);
nor U4143 (N_4143,In_2413,In_503);
and U4144 (N_4144,In_2514,In_2767);
nor U4145 (N_4145,In_582,In_732);
nand U4146 (N_4146,In_1769,In_597);
nor U4147 (N_4147,In_1361,In_1904);
xor U4148 (N_4148,In_1206,In_1459);
nand U4149 (N_4149,In_2829,In_848);
and U4150 (N_4150,In_2392,In_1614);
nand U4151 (N_4151,In_1286,In_2552);
xor U4152 (N_4152,In_2979,In_2025);
xor U4153 (N_4153,In_1502,In_2153);
or U4154 (N_4154,In_866,In_464);
nor U4155 (N_4155,In_1060,In_706);
nor U4156 (N_4156,In_2340,In_1812);
xnor U4157 (N_4157,In_1333,In_981);
or U4158 (N_4158,In_2606,In_2520);
and U4159 (N_4159,In_2235,In_1914);
xnor U4160 (N_4160,In_603,In_1197);
xnor U4161 (N_4161,In_2795,In_2640);
and U4162 (N_4162,In_142,In_865);
xnor U4163 (N_4163,In_1687,In_2376);
and U4164 (N_4164,In_1235,In_2110);
nand U4165 (N_4165,In_1414,In_1136);
nand U4166 (N_4166,In_2534,In_1028);
and U4167 (N_4167,In_1568,In_2197);
or U4168 (N_4168,In_2528,In_2977);
nor U4169 (N_4169,In_2328,In_517);
xnor U4170 (N_4170,In_2262,In_1957);
xor U4171 (N_4171,In_1009,In_1963);
xnor U4172 (N_4172,In_191,In_1459);
and U4173 (N_4173,In_140,In_1816);
or U4174 (N_4174,In_1559,In_1339);
and U4175 (N_4175,In_2013,In_2212);
nand U4176 (N_4176,In_2937,In_99);
and U4177 (N_4177,In_2592,In_1006);
nand U4178 (N_4178,In_2421,In_64);
and U4179 (N_4179,In_2077,In_690);
xor U4180 (N_4180,In_1369,In_496);
and U4181 (N_4181,In_1381,In_2687);
and U4182 (N_4182,In_1525,In_811);
nor U4183 (N_4183,In_919,In_39);
nor U4184 (N_4184,In_1705,In_912);
nor U4185 (N_4185,In_2848,In_2412);
xor U4186 (N_4186,In_48,In_684);
nand U4187 (N_4187,In_2051,In_746);
nand U4188 (N_4188,In_885,In_492);
xor U4189 (N_4189,In_1118,In_351);
nand U4190 (N_4190,In_1865,In_1200);
nand U4191 (N_4191,In_2783,In_2644);
nor U4192 (N_4192,In_2617,In_2410);
nand U4193 (N_4193,In_2193,In_2501);
and U4194 (N_4194,In_2459,In_134);
nand U4195 (N_4195,In_1333,In_1778);
xor U4196 (N_4196,In_2321,In_1515);
nand U4197 (N_4197,In_1582,In_2382);
or U4198 (N_4198,In_210,In_2868);
xor U4199 (N_4199,In_2693,In_1810);
and U4200 (N_4200,In_127,In_2035);
and U4201 (N_4201,In_1349,In_567);
nor U4202 (N_4202,In_1048,In_2946);
nor U4203 (N_4203,In_2348,In_2663);
or U4204 (N_4204,In_1585,In_2767);
xnor U4205 (N_4205,In_1163,In_1757);
nand U4206 (N_4206,In_2890,In_2087);
nand U4207 (N_4207,In_1795,In_614);
or U4208 (N_4208,In_440,In_2873);
and U4209 (N_4209,In_1328,In_162);
and U4210 (N_4210,In_257,In_2724);
or U4211 (N_4211,In_1830,In_2081);
and U4212 (N_4212,In_1907,In_2370);
or U4213 (N_4213,In_2267,In_326);
xor U4214 (N_4214,In_2132,In_1707);
or U4215 (N_4215,In_128,In_2245);
xnor U4216 (N_4216,In_1767,In_1261);
nor U4217 (N_4217,In_885,In_2679);
and U4218 (N_4218,In_460,In_714);
or U4219 (N_4219,In_2204,In_1061);
xor U4220 (N_4220,In_417,In_833);
and U4221 (N_4221,In_1732,In_152);
and U4222 (N_4222,In_787,In_396);
or U4223 (N_4223,In_1713,In_2299);
or U4224 (N_4224,In_1527,In_2610);
xnor U4225 (N_4225,In_2255,In_2406);
or U4226 (N_4226,In_2881,In_220);
or U4227 (N_4227,In_1947,In_722);
nor U4228 (N_4228,In_1594,In_1816);
nor U4229 (N_4229,In_1056,In_2484);
or U4230 (N_4230,In_2671,In_2378);
xor U4231 (N_4231,In_2514,In_84);
and U4232 (N_4232,In_1834,In_657);
nor U4233 (N_4233,In_1110,In_1258);
nand U4234 (N_4234,In_2281,In_2798);
or U4235 (N_4235,In_2792,In_803);
nand U4236 (N_4236,In_953,In_11);
or U4237 (N_4237,In_672,In_2827);
or U4238 (N_4238,In_1812,In_481);
nand U4239 (N_4239,In_1411,In_2893);
xor U4240 (N_4240,In_1864,In_1104);
nand U4241 (N_4241,In_2507,In_1374);
and U4242 (N_4242,In_2230,In_1843);
or U4243 (N_4243,In_2224,In_2276);
nor U4244 (N_4244,In_902,In_1120);
nor U4245 (N_4245,In_2111,In_121);
nor U4246 (N_4246,In_197,In_1459);
nor U4247 (N_4247,In_1975,In_1471);
or U4248 (N_4248,In_51,In_1642);
nand U4249 (N_4249,In_43,In_3);
nor U4250 (N_4250,In_1595,In_309);
nor U4251 (N_4251,In_1635,In_2970);
nand U4252 (N_4252,In_1254,In_2400);
xnor U4253 (N_4253,In_1943,In_219);
xnor U4254 (N_4254,In_828,In_2384);
nand U4255 (N_4255,In_2405,In_2633);
nor U4256 (N_4256,In_2184,In_2012);
nand U4257 (N_4257,In_2038,In_2512);
nor U4258 (N_4258,In_1364,In_2256);
or U4259 (N_4259,In_601,In_263);
or U4260 (N_4260,In_2087,In_1031);
and U4261 (N_4261,In_1608,In_1567);
and U4262 (N_4262,In_1482,In_1165);
and U4263 (N_4263,In_590,In_2135);
nor U4264 (N_4264,In_240,In_2285);
xnor U4265 (N_4265,In_1543,In_1398);
and U4266 (N_4266,In_2524,In_243);
or U4267 (N_4267,In_1216,In_2502);
and U4268 (N_4268,In_1263,In_1583);
nand U4269 (N_4269,In_1898,In_2134);
or U4270 (N_4270,In_649,In_1983);
xnor U4271 (N_4271,In_457,In_2360);
and U4272 (N_4272,In_1633,In_1453);
or U4273 (N_4273,In_2049,In_1576);
and U4274 (N_4274,In_2572,In_2483);
nor U4275 (N_4275,In_161,In_1205);
and U4276 (N_4276,In_1830,In_2499);
and U4277 (N_4277,In_40,In_2033);
or U4278 (N_4278,In_723,In_2343);
or U4279 (N_4279,In_1550,In_376);
and U4280 (N_4280,In_1404,In_868);
nor U4281 (N_4281,In_699,In_1321);
nand U4282 (N_4282,In_2023,In_113);
xnor U4283 (N_4283,In_2094,In_817);
xnor U4284 (N_4284,In_828,In_1361);
and U4285 (N_4285,In_494,In_2408);
nor U4286 (N_4286,In_2292,In_2543);
or U4287 (N_4287,In_1957,In_2787);
nor U4288 (N_4288,In_1589,In_446);
nand U4289 (N_4289,In_1877,In_909);
xor U4290 (N_4290,In_598,In_2690);
or U4291 (N_4291,In_990,In_2473);
xor U4292 (N_4292,In_2804,In_2446);
or U4293 (N_4293,In_2411,In_524);
or U4294 (N_4294,In_199,In_626);
or U4295 (N_4295,In_2970,In_2079);
nand U4296 (N_4296,In_2582,In_2243);
nand U4297 (N_4297,In_507,In_1838);
xnor U4298 (N_4298,In_2569,In_2058);
nor U4299 (N_4299,In_531,In_590);
and U4300 (N_4300,In_1957,In_2696);
nand U4301 (N_4301,In_1736,In_1359);
nand U4302 (N_4302,In_1089,In_494);
xnor U4303 (N_4303,In_479,In_2743);
and U4304 (N_4304,In_2661,In_113);
and U4305 (N_4305,In_1756,In_976);
xor U4306 (N_4306,In_1426,In_1195);
nor U4307 (N_4307,In_519,In_2846);
or U4308 (N_4308,In_1294,In_664);
or U4309 (N_4309,In_151,In_2994);
or U4310 (N_4310,In_1661,In_2300);
or U4311 (N_4311,In_1555,In_2715);
or U4312 (N_4312,In_155,In_1389);
or U4313 (N_4313,In_87,In_1553);
nor U4314 (N_4314,In_2394,In_2129);
nand U4315 (N_4315,In_470,In_41);
nor U4316 (N_4316,In_2403,In_1561);
and U4317 (N_4317,In_2255,In_1593);
and U4318 (N_4318,In_1003,In_2452);
or U4319 (N_4319,In_853,In_2689);
nand U4320 (N_4320,In_2124,In_1908);
xor U4321 (N_4321,In_1396,In_383);
nand U4322 (N_4322,In_35,In_108);
and U4323 (N_4323,In_2296,In_2156);
and U4324 (N_4324,In_2848,In_2061);
nor U4325 (N_4325,In_521,In_2903);
and U4326 (N_4326,In_1462,In_2432);
nand U4327 (N_4327,In_165,In_2249);
nand U4328 (N_4328,In_1298,In_1213);
and U4329 (N_4329,In_2736,In_2968);
xor U4330 (N_4330,In_2186,In_2191);
nand U4331 (N_4331,In_2469,In_112);
nand U4332 (N_4332,In_2140,In_2848);
nand U4333 (N_4333,In_224,In_568);
nand U4334 (N_4334,In_1654,In_1849);
xnor U4335 (N_4335,In_2600,In_1796);
xor U4336 (N_4336,In_229,In_564);
nor U4337 (N_4337,In_913,In_1745);
or U4338 (N_4338,In_408,In_2198);
nand U4339 (N_4339,In_2403,In_2425);
nor U4340 (N_4340,In_2766,In_79);
nand U4341 (N_4341,In_1923,In_1802);
and U4342 (N_4342,In_2700,In_2707);
xnor U4343 (N_4343,In_1140,In_1143);
nand U4344 (N_4344,In_2797,In_1461);
xnor U4345 (N_4345,In_2607,In_2679);
and U4346 (N_4346,In_1767,In_2438);
nor U4347 (N_4347,In_1440,In_2525);
and U4348 (N_4348,In_2468,In_934);
and U4349 (N_4349,In_240,In_2678);
xor U4350 (N_4350,In_741,In_2616);
or U4351 (N_4351,In_1727,In_752);
nor U4352 (N_4352,In_2399,In_257);
and U4353 (N_4353,In_661,In_2700);
xor U4354 (N_4354,In_1324,In_2193);
and U4355 (N_4355,In_590,In_577);
xor U4356 (N_4356,In_984,In_105);
and U4357 (N_4357,In_2980,In_1577);
xnor U4358 (N_4358,In_2175,In_634);
xnor U4359 (N_4359,In_2254,In_1537);
and U4360 (N_4360,In_741,In_82);
and U4361 (N_4361,In_2942,In_921);
nor U4362 (N_4362,In_2084,In_2610);
nand U4363 (N_4363,In_180,In_1479);
or U4364 (N_4364,In_2828,In_2930);
nor U4365 (N_4365,In_2771,In_694);
nor U4366 (N_4366,In_612,In_2711);
xor U4367 (N_4367,In_2466,In_1442);
xnor U4368 (N_4368,In_2176,In_903);
and U4369 (N_4369,In_2424,In_131);
or U4370 (N_4370,In_1093,In_2512);
nor U4371 (N_4371,In_2195,In_2261);
nor U4372 (N_4372,In_1656,In_1334);
nand U4373 (N_4373,In_2263,In_2215);
nor U4374 (N_4374,In_724,In_1291);
xor U4375 (N_4375,In_2320,In_2710);
xor U4376 (N_4376,In_1662,In_1713);
nor U4377 (N_4377,In_1261,In_1338);
nand U4378 (N_4378,In_1875,In_97);
xor U4379 (N_4379,In_2183,In_442);
nand U4380 (N_4380,In_2353,In_2147);
and U4381 (N_4381,In_1981,In_2474);
nand U4382 (N_4382,In_365,In_1302);
nand U4383 (N_4383,In_2418,In_1969);
or U4384 (N_4384,In_2135,In_1745);
and U4385 (N_4385,In_1320,In_2179);
xor U4386 (N_4386,In_2292,In_2194);
or U4387 (N_4387,In_77,In_309);
xor U4388 (N_4388,In_234,In_2958);
nand U4389 (N_4389,In_274,In_1824);
and U4390 (N_4390,In_833,In_211);
and U4391 (N_4391,In_884,In_2768);
and U4392 (N_4392,In_2966,In_2247);
nor U4393 (N_4393,In_2968,In_1372);
xor U4394 (N_4394,In_1451,In_1627);
or U4395 (N_4395,In_1543,In_1669);
nand U4396 (N_4396,In_1547,In_992);
nor U4397 (N_4397,In_241,In_432);
nor U4398 (N_4398,In_579,In_1097);
xnor U4399 (N_4399,In_624,In_1879);
or U4400 (N_4400,In_2897,In_687);
nand U4401 (N_4401,In_2329,In_457);
nor U4402 (N_4402,In_1713,In_1121);
or U4403 (N_4403,In_832,In_30);
xor U4404 (N_4404,In_1263,In_2180);
xnor U4405 (N_4405,In_335,In_1269);
and U4406 (N_4406,In_2646,In_1054);
nand U4407 (N_4407,In_911,In_1155);
nand U4408 (N_4408,In_1291,In_2222);
or U4409 (N_4409,In_1627,In_586);
or U4410 (N_4410,In_2923,In_2313);
xor U4411 (N_4411,In_1129,In_1566);
xnor U4412 (N_4412,In_527,In_1273);
or U4413 (N_4413,In_1863,In_2456);
nor U4414 (N_4414,In_1337,In_2659);
nand U4415 (N_4415,In_1991,In_1533);
or U4416 (N_4416,In_1309,In_2096);
or U4417 (N_4417,In_327,In_173);
or U4418 (N_4418,In_2235,In_1010);
nand U4419 (N_4419,In_1721,In_307);
nor U4420 (N_4420,In_2110,In_1911);
nor U4421 (N_4421,In_342,In_2787);
nor U4422 (N_4422,In_1223,In_1923);
or U4423 (N_4423,In_2726,In_2794);
nor U4424 (N_4424,In_1114,In_2299);
nand U4425 (N_4425,In_955,In_2045);
xor U4426 (N_4426,In_2776,In_1984);
or U4427 (N_4427,In_323,In_1340);
xnor U4428 (N_4428,In_620,In_1048);
nor U4429 (N_4429,In_1830,In_2312);
or U4430 (N_4430,In_2320,In_111);
nor U4431 (N_4431,In_955,In_194);
nand U4432 (N_4432,In_304,In_588);
and U4433 (N_4433,In_1939,In_2196);
nor U4434 (N_4434,In_825,In_307);
or U4435 (N_4435,In_261,In_2998);
nand U4436 (N_4436,In_1488,In_1345);
and U4437 (N_4437,In_893,In_2242);
and U4438 (N_4438,In_1522,In_2614);
nand U4439 (N_4439,In_1172,In_731);
xnor U4440 (N_4440,In_811,In_28);
nand U4441 (N_4441,In_1024,In_2890);
or U4442 (N_4442,In_1461,In_2983);
and U4443 (N_4443,In_1288,In_510);
nor U4444 (N_4444,In_2990,In_2861);
xnor U4445 (N_4445,In_1904,In_2220);
nand U4446 (N_4446,In_2519,In_800);
nor U4447 (N_4447,In_1763,In_1324);
or U4448 (N_4448,In_1705,In_2850);
nor U4449 (N_4449,In_2583,In_348);
and U4450 (N_4450,In_217,In_2150);
nor U4451 (N_4451,In_299,In_2273);
xor U4452 (N_4452,In_2673,In_958);
nor U4453 (N_4453,In_1796,In_1088);
and U4454 (N_4454,In_1579,In_1759);
or U4455 (N_4455,In_1560,In_2965);
and U4456 (N_4456,In_1635,In_2226);
and U4457 (N_4457,In_1418,In_1349);
xor U4458 (N_4458,In_1531,In_192);
nand U4459 (N_4459,In_1855,In_16);
or U4460 (N_4460,In_36,In_649);
or U4461 (N_4461,In_1114,In_458);
xor U4462 (N_4462,In_812,In_99);
and U4463 (N_4463,In_2320,In_2958);
and U4464 (N_4464,In_2769,In_856);
and U4465 (N_4465,In_1065,In_1992);
nor U4466 (N_4466,In_2221,In_390);
nand U4467 (N_4467,In_1277,In_2068);
nand U4468 (N_4468,In_2388,In_663);
and U4469 (N_4469,In_1419,In_2211);
nor U4470 (N_4470,In_2286,In_2151);
or U4471 (N_4471,In_1418,In_1370);
xor U4472 (N_4472,In_639,In_1137);
or U4473 (N_4473,In_1186,In_1012);
nor U4474 (N_4474,In_2577,In_2891);
nor U4475 (N_4475,In_605,In_2520);
nand U4476 (N_4476,In_2519,In_1954);
and U4477 (N_4477,In_1165,In_1794);
nand U4478 (N_4478,In_1585,In_2581);
nor U4479 (N_4479,In_1529,In_193);
and U4480 (N_4480,In_2950,In_2913);
and U4481 (N_4481,In_2491,In_2939);
nor U4482 (N_4482,In_138,In_2947);
nor U4483 (N_4483,In_2692,In_1723);
nand U4484 (N_4484,In_2994,In_751);
nand U4485 (N_4485,In_907,In_314);
or U4486 (N_4486,In_2127,In_266);
or U4487 (N_4487,In_1883,In_867);
and U4488 (N_4488,In_794,In_1694);
nor U4489 (N_4489,In_59,In_1330);
xor U4490 (N_4490,In_544,In_1784);
and U4491 (N_4491,In_810,In_709);
or U4492 (N_4492,In_860,In_1472);
and U4493 (N_4493,In_927,In_2822);
and U4494 (N_4494,In_1952,In_2414);
xor U4495 (N_4495,In_410,In_2043);
nand U4496 (N_4496,In_2073,In_1610);
xor U4497 (N_4497,In_1124,In_2987);
xnor U4498 (N_4498,In_801,In_2360);
xor U4499 (N_4499,In_2274,In_2960);
nor U4500 (N_4500,In_1375,In_148);
xnor U4501 (N_4501,In_950,In_1743);
xor U4502 (N_4502,In_2594,In_267);
nor U4503 (N_4503,In_2787,In_2752);
xor U4504 (N_4504,In_2233,In_168);
and U4505 (N_4505,In_2710,In_2960);
nor U4506 (N_4506,In_1957,In_1271);
or U4507 (N_4507,In_1350,In_460);
nand U4508 (N_4508,In_1224,In_2028);
and U4509 (N_4509,In_2682,In_1590);
nor U4510 (N_4510,In_1901,In_190);
nor U4511 (N_4511,In_2494,In_2700);
nor U4512 (N_4512,In_257,In_2184);
xnor U4513 (N_4513,In_422,In_1455);
xor U4514 (N_4514,In_1429,In_1089);
or U4515 (N_4515,In_1164,In_1834);
nor U4516 (N_4516,In_2404,In_3);
nand U4517 (N_4517,In_2525,In_318);
or U4518 (N_4518,In_379,In_1295);
nand U4519 (N_4519,In_2362,In_2628);
or U4520 (N_4520,In_2382,In_2679);
and U4521 (N_4521,In_571,In_61);
or U4522 (N_4522,In_2892,In_1635);
or U4523 (N_4523,In_2014,In_1096);
nand U4524 (N_4524,In_1076,In_1661);
nor U4525 (N_4525,In_592,In_751);
nor U4526 (N_4526,In_2364,In_1718);
xor U4527 (N_4527,In_2075,In_541);
and U4528 (N_4528,In_446,In_2786);
or U4529 (N_4529,In_2002,In_887);
or U4530 (N_4530,In_2416,In_2025);
nor U4531 (N_4531,In_1313,In_290);
nor U4532 (N_4532,In_1041,In_1789);
nand U4533 (N_4533,In_1729,In_345);
nand U4534 (N_4534,In_1768,In_1844);
and U4535 (N_4535,In_29,In_1069);
nor U4536 (N_4536,In_1162,In_1022);
nand U4537 (N_4537,In_1400,In_2167);
nand U4538 (N_4538,In_1994,In_1254);
and U4539 (N_4539,In_165,In_2796);
or U4540 (N_4540,In_1308,In_2778);
xor U4541 (N_4541,In_2333,In_2273);
or U4542 (N_4542,In_2586,In_644);
nand U4543 (N_4543,In_1375,In_2109);
and U4544 (N_4544,In_440,In_1222);
nand U4545 (N_4545,In_2007,In_2673);
xnor U4546 (N_4546,In_2630,In_1636);
and U4547 (N_4547,In_885,In_1416);
nor U4548 (N_4548,In_2186,In_2025);
nor U4549 (N_4549,In_1397,In_255);
or U4550 (N_4550,In_1226,In_356);
nand U4551 (N_4551,In_188,In_1980);
nor U4552 (N_4552,In_2557,In_357);
nand U4553 (N_4553,In_1486,In_1933);
and U4554 (N_4554,In_1768,In_2775);
or U4555 (N_4555,In_663,In_1349);
nor U4556 (N_4556,In_2239,In_1503);
and U4557 (N_4557,In_1518,In_2704);
xor U4558 (N_4558,In_2456,In_285);
and U4559 (N_4559,In_2212,In_1655);
or U4560 (N_4560,In_1138,In_2329);
nand U4561 (N_4561,In_928,In_2618);
nor U4562 (N_4562,In_2305,In_1936);
or U4563 (N_4563,In_2842,In_1061);
xnor U4564 (N_4564,In_1878,In_1226);
nor U4565 (N_4565,In_2268,In_66);
xor U4566 (N_4566,In_2017,In_385);
xor U4567 (N_4567,In_2507,In_2780);
or U4568 (N_4568,In_1753,In_250);
or U4569 (N_4569,In_2551,In_2350);
xnor U4570 (N_4570,In_763,In_2049);
or U4571 (N_4571,In_470,In_430);
nor U4572 (N_4572,In_1441,In_2483);
nand U4573 (N_4573,In_2255,In_1780);
and U4574 (N_4574,In_2869,In_1690);
nor U4575 (N_4575,In_1472,In_1535);
and U4576 (N_4576,In_1677,In_2748);
xor U4577 (N_4577,In_1504,In_2250);
and U4578 (N_4578,In_2597,In_1471);
nand U4579 (N_4579,In_1282,In_1539);
and U4580 (N_4580,In_10,In_1895);
xnor U4581 (N_4581,In_2142,In_632);
xor U4582 (N_4582,In_206,In_1790);
and U4583 (N_4583,In_1964,In_324);
xor U4584 (N_4584,In_787,In_504);
xnor U4585 (N_4585,In_1532,In_114);
or U4586 (N_4586,In_2211,In_2947);
or U4587 (N_4587,In_487,In_1085);
or U4588 (N_4588,In_2693,In_478);
nor U4589 (N_4589,In_356,In_1281);
or U4590 (N_4590,In_1759,In_932);
nor U4591 (N_4591,In_1481,In_1277);
nor U4592 (N_4592,In_2488,In_1440);
nor U4593 (N_4593,In_407,In_2419);
nand U4594 (N_4594,In_976,In_2522);
nand U4595 (N_4595,In_7,In_1904);
xnor U4596 (N_4596,In_1188,In_1254);
xor U4597 (N_4597,In_1941,In_2524);
nor U4598 (N_4598,In_1518,In_1227);
and U4599 (N_4599,In_1114,In_587);
nand U4600 (N_4600,In_1656,In_118);
nor U4601 (N_4601,In_1224,In_461);
xnor U4602 (N_4602,In_2233,In_1608);
nor U4603 (N_4603,In_1070,In_254);
xor U4604 (N_4604,In_1566,In_2623);
or U4605 (N_4605,In_1067,In_308);
nand U4606 (N_4606,In_2612,In_1228);
nand U4607 (N_4607,In_2224,In_2026);
nand U4608 (N_4608,In_2124,In_1569);
or U4609 (N_4609,In_303,In_2174);
and U4610 (N_4610,In_2822,In_1422);
xor U4611 (N_4611,In_1869,In_2914);
nand U4612 (N_4612,In_799,In_1453);
and U4613 (N_4613,In_1394,In_2524);
nor U4614 (N_4614,In_1211,In_626);
or U4615 (N_4615,In_880,In_224);
or U4616 (N_4616,In_349,In_2740);
nand U4617 (N_4617,In_2939,In_1128);
xor U4618 (N_4618,In_1662,In_1373);
or U4619 (N_4619,In_1512,In_362);
and U4620 (N_4620,In_5,In_2258);
nand U4621 (N_4621,In_406,In_2669);
nand U4622 (N_4622,In_141,In_1237);
and U4623 (N_4623,In_1030,In_616);
and U4624 (N_4624,In_1527,In_1235);
or U4625 (N_4625,In_2684,In_1584);
xor U4626 (N_4626,In_244,In_30);
nor U4627 (N_4627,In_2018,In_2745);
and U4628 (N_4628,In_2962,In_1967);
xor U4629 (N_4629,In_1553,In_725);
nor U4630 (N_4630,In_1499,In_1099);
xnor U4631 (N_4631,In_1548,In_1915);
nand U4632 (N_4632,In_2555,In_823);
xor U4633 (N_4633,In_1482,In_2792);
nor U4634 (N_4634,In_684,In_891);
nand U4635 (N_4635,In_575,In_245);
and U4636 (N_4636,In_2639,In_1758);
xnor U4637 (N_4637,In_324,In_1157);
nand U4638 (N_4638,In_459,In_1486);
or U4639 (N_4639,In_2902,In_2045);
and U4640 (N_4640,In_833,In_517);
or U4641 (N_4641,In_544,In_503);
and U4642 (N_4642,In_2402,In_2422);
nand U4643 (N_4643,In_2575,In_359);
xnor U4644 (N_4644,In_553,In_564);
and U4645 (N_4645,In_2752,In_2702);
nand U4646 (N_4646,In_1739,In_588);
nor U4647 (N_4647,In_1200,In_1439);
nor U4648 (N_4648,In_2454,In_1063);
and U4649 (N_4649,In_713,In_2236);
nor U4650 (N_4650,In_1840,In_928);
and U4651 (N_4651,In_1629,In_420);
or U4652 (N_4652,In_385,In_2029);
nand U4653 (N_4653,In_679,In_2940);
nor U4654 (N_4654,In_394,In_2262);
xor U4655 (N_4655,In_2103,In_347);
or U4656 (N_4656,In_906,In_1143);
nand U4657 (N_4657,In_2217,In_2427);
and U4658 (N_4658,In_1044,In_845);
and U4659 (N_4659,In_2351,In_777);
nand U4660 (N_4660,In_876,In_257);
nor U4661 (N_4661,In_1981,In_1654);
nand U4662 (N_4662,In_2068,In_725);
xor U4663 (N_4663,In_1405,In_2785);
nand U4664 (N_4664,In_1147,In_1030);
xor U4665 (N_4665,In_277,In_137);
and U4666 (N_4666,In_46,In_2005);
nand U4667 (N_4667,In_2371,In_686);
nand U4668 (N_4668,In_1477,In_71);
or U4669 (N_4669,In_406,In_2210);
xnor U4670 (N_4670,In_586,In_2963);
xor U4671 (N_4671,In_34,In_1359);
or U4672 (N_4672,In_2008,In_2201);
and U4673 (N_4673,In_425,In_1429);
nand U4674 (N_4674,In_1827,In_2109);
nor U4675 (N_4675,In_619,In_1461);
nand U4676 (N_4676,In_2105,In_41);
and U4677 (N_4677,In_899,In_169);
nand U4678 (N_4678,In_1921,In_406);
nor U4679 (N_4679,In_2337,In_2212);
xnor U4680 (N_4680,In_2877,In_2861);
nor U4681 (N_4681,In_1946,In_880);
nand U4682 (N_4682,In_810,In_659);
nor U4683 (N_4683,In_2113,In_707);
nand U4684 (N_4684,In_484,In_571);
or U4685 (N_4685,In_135,In_1889);
nand U4686 (N_4686,In_870,In_633);
nand U4687 (N_4687,In_643,In_2459);
or U4688 (N_4688,In_155,In_775);
nor U4689 (N_4689,In_1698,In_380);
xnor U4690 (N_4690,In_1430,In_1184);
or U4691 (N_4691,In_146,In_2034);
nand U4692 (N_4692,In_1194,In_481);
nand U4693 (N_4693,In_1562,In_2131);
xor U4694 (N_4694,In_2981,In_1814);
nor U4695 (N_4695,In_1107,In_2368);
nand U4696 (N_4696,In_1533,In_324);
or U4697 (N_4697,In_1524,In_1847);
and U4698 (N_4698,In_1830,In_1746);
and U4699 (N_4699,In_343,In_1456);
or U4700 (N_4700,In_2653,In_1424);
nor U4701 (N_4701,In_1673,In_1310);
nor U4702 (N_4702,In_1021,In_907);
nand U4703 (N_4703,In_470,In_453);
nand U4704 (N_4704,In_1081,In_259);
and U4705 (N_4705,In_855,In_2824);
and U4706 (N_4706,In_2260,In_2433);
xnor U4707 (N_4707,In_2125,In_2652);
and U4708 (N_4708,In_925,In_1596);
nand U4709 (N_4709,In_2250,In_2497);
nand U4710 (N_4710,In_805,In_2980);
or U4711 (N_4711,In_2275,In_2286);
nor U4712 (N_4712,In_1586,In_258);
and U4713 (N_4713,In_2110,In_185);
and U4714 (N_4714,In_859,In_2828);
and U4715 (N_4715,In_1107,In_242);
or U4716 (N_4716,In_2968,In_2217);
and U4717 (N_4717,In_586,In_239);
nor U4718 (N_4718,In_1804,In_2629);
or U4719 (N_4719,In_637,In_2733);
nor U4720 (N_4720,In_1050,In_2868);
nor U4721 (N_4721,In_1776,In_317);
xor U4722 (N_4722,In_1104,In_2047);
nor U4723 (N_4723,In_475,In_2455);
nand U4724 (N_4724,In_2669,In_508);
xnor U4725 (N_4725,In_1323,In_1627);
nand U4726 (N_4726,In_2814,In_1792);
or U4727 (N_4727,In_1598,In_251);
or U4728 (N_4728,In_942,In_2947);
or U4729 (N_4729,In_2077,In_506);
xor U4730 (N_4730,In_1789,In_2515);
nor U4731 (N_4731,In_518,In_2934);
and U4732 (N_4732,In_441,In_2457);
and U4733 (N_4733,In_2070,In_2529);
or U4734 (N_4734,In_2325,In_1611);
xnor U4735 (N_4735,In_2585,In_724);
nand U4736 (N_4736,In_2688,In_1775);
nor U4737 (N_4737,In_1700,In_599);
or U4738 (N_4738,In_863,In_1424);
or U4739 (N_4739,In_1540,In_2761);
nand U4740 (N_4740,In_1667,In_1528);
and U4741 (N_4741,In_208,In_474);
or U4742 (N_4742,In_2447,In_2699);
nand U4743 (N_4743,In_2982,In_2746);
and U4744 (N_4744,In_900,In_1165);
xor U4745 (N_4745,In_2620,In_288);
nor U4746 (N_4746,In_1654,In_2552);
or U4747 (N_4747,In_1006,In_1692);
xor U4748 (N_4748,In_2559,In_2305);
and U4749 (N_4749,In_1219,In_1695);
and U4750 (N_4750,In_163,In_1320);
or U4751 (N_4751,In_1228,In_595);
or U4752 (N_4752,In_249,In_1930);
or U4753 (N_4753,In_1082,In_1112);
xor U4754 (N_4754,In_2927,In_1050);
xor U4755 (N_4755,In_2998,In_185);
nor U4756 (N_4756,In_1897,In_241);
nand U4757 (N_4757,In_691,In_1414);
xor U4758 (N_4758,In_2340,In_433);
or U4759 (N_4759,In_2358,In_1382);
nor U4760 (N_4760,In_1643,In_2526);
nand U4761 (N_4761,In_609,In_1099);
and U4762 (N_4762,In_2392,In_929);
nand U4763 (N_4763,In_495,In_2741);
or U4764 (N_4764,In_262,In_142);
nand U4765 (N_4765,In_1135,In_2630);
nand U4766 (N_4766,In_850,In_171);
and U4767 (N_4767,In_76,In_2184);
nand U4768 (N_4768,In_296,In_2854);
or U4769 (N_4769,In_794,In_2333);
nor U4770 (N_4770,In_915,In_22);
or U4771 (N_4771,In_529,In_231);
nand U4772 (N_4772,In_435,In_638);
nor U4773 (N_4773,In_2263,In_2926);
and U4774 (N_4774,In_843,In_1986);
and U4775 (N_4775,In_2424,In_1634);
nand U4776 (N_4776,In_65,In_220);
and U4777 (N_4777,In_553,In_1868);
xnor U4778 (N_4778,In_362,In_2437);
nand U4779 (N_4779,In_2933,In_1873);
nor U4780 (N_4780,In_1534,In_1254);
or U4781 (N_4781,In_2342,In_2653);
and U4782 (N_4782,In_639,In_1850);
and U4783 (N_4783,In_2043,In_1014);
and U4784 (N_4784,In_682,In_81);
xnor U4785 (N_4785,In_2809,In_1684);
nor U4786 (N_4786,In_38,In_2899);
or U4787 (N_4787,In_1552,In_374);
and U4788 (N_4788,In_982,In_591);
nand U4789 (N_4789,In_1199,In_2985);
nand U4790 (N_4790,In_2003,In_1332);
xnor U4791 (N_4791,In_2267,In_11);
or U4792 (N_4792,In_191,In_1707);
xnor U4793 (N_4793,In_1596,In_926);
nor U4794 (N_4794,In_510,In_2494);
nor U4795 (N_4795,In_1363,In_85);
nor U4796 (N_4796,In_2878,In_2573);
nand U4797 (N_4797,In_769,In_1794);
nor U4798 (N_4798,In_168,In_1964);
xor U4799 (N_4799,In_1266,In_1902);
or U4800 (N_4800,In_1142,In_2986);
nor U4801 (N_4801,In_2127,In_488);
nand U4802 (N_4802,In_2989,In_254);
nor U4803 (N_4803,In_927,In_2220);
or U4804 (N_4804,In_1263,In_269);
nand U4805 (N_4805,In_248,In_2892);
nor U4806 (N_4806,In_367,In_2276);
nor U4807 (N_4807,In_63,In_2015);
xor U4808 (N_4808,In_125,In_2584);
xor U4809 (N_4809,In_2922,In_776);
nor U4810 (N_4810,In_402,In_2872);
nand U4811 (N_4811,In_1633,In_800);
or U4812 (N_4812,In_390,In_1918);
or U4813 (N_4813,In_2400,In_1502);
nor U4814 (N_4814,In_1326,In_1540);
nor U4815 (N_4815,In_620,In_449);
nor U4816 (N_4816,In_457,In_977);
xnor U4817 (N_4817,In_1111,In_1669);
and U4818 (N_4818,In_2214,In_2433);
nand U4819 (N_4819,In_2237,In_223);
nor U4820 (N_4820,In_2036,In_96);
xor U4821 (N_4821,In_641,In_879);
nand U4822 (N_4822,In_1186,In_2369);
nor U4823 (N_4823,In_568,In_1458);
xnor U4824 (N_4824,In_1224,In_1166);
and U4825 (N_4825,In_1447,In_1901);
xnor U4826 (N_4826,In_1135,In_2263);
and U4827 (N_4827,In_2936,In_37);
nand U4828 (N_4828,In_1785,In_2523);
or U4829 (N_4829,In_2455,In_2807);
and U4830 (N_4830,In_1977,In_1291);
or U4831 (N_4831,In_90,In_2079);
and U4832 (N_4832,In_2369,In_34);
or U4833 (N_4833,In_2073,In_2961);
or U4834 (N_4834,In_1559,In_961);
or U4835 (N_4835,In_2733,In_389);
and U4836 (N_4836,In_562,In_959);
and U4837 (N_4837,In_2932,In_2326);
and U4838 (N_4838,In_1041,In_1383);
nor U4839 (N_4839,In_2293,In_2629);
xor U4840 (N_4840,In_1391,In_2439);
nor U4841 (N_4841,In_447,In_1652);
or U4842 (N_4842,In_1000,In_1228);
xor U4843 (N_4843,In_934,In_1193);
xnor U4844 (N_4844,In_291,In_523);
or U4845 (N_4845,In_2612,In_1596);
and U4846 (N_4846,In_1616,In_2705);
or U4847 (N_4847,In_18,In_533);
nand U4848 (N_4848,In_2746,In_1766);
nand U4849 (N_4849,In_1595,In_1282);
xnor U4850 (N_4850,In_413,In_603);
and U4851 (N_4851,In_1487,In_730);
or U4852 (N_4852,In_509,In_1086);
nand U4853 (N_4853,In_2616,In_1693);
nand U4854 (N_4854,In_1969,In_1546);
or U4855 (N_4855,In_1511,In_2637);
nand U4856 (N_4856,In_1687,In_63);
nor U4857 (N_4857,In_1728,In_1376);
nand U4858 (N_4858,In_193,In_2124);
or U4859 (N_4859,In_974,In_2027);
nor U4860 (N_4860,In_2609,In_463);
nand U4861 (N_4861,In_2154,In_2701);
and U4862 (N_4862,In_290,In_1367);
and U4863 (N_4863,In_2079,In_1664);
nor U4864 (N_4864,In_2859,In_611);
nor U4865 (N_4865,In_1769,In_795);
and U4866 (N_4866,In_1852,In_617);
and U4867 (N_4867,In_124,In_2390);
nor U4868 (N_4868,In_130,In_2028);
and U4869 (N_4869,In_977,In_2789);
nand U4870 (N_4870,In_1815,In_807);
or U4871 (N_4871,In_754,In_2826);
nand U4872 (N_4872,In_942,In_153);
nor U4873 (N_4873,In_1100,In_228);
xor U4874 (N_4874,In_2278,In_2675);
and U4875 (N_4875,In_2837,In_1329);
and U4876 (N_4876,In_2582,In_2915);
or U4877 (N_4877,In_159,In_121);
xnor U4878 (N_4878,In_2910,In_1780);
or U4879 (N_4879,In_1260,In_519);
nand U4880 (N_4880,In_1860,In_2668);
and U4881 (N_4881,In_99,In_2874);
nor U4882 (N_4882,In_1623,In_245);
or U4883 (N_4883,In_2751,In_1903);
xor U4884 (N_4884,In_1949,In_1387);
nor U4885 (N_4885,In_1534,In_2840);
nand U4886 (N_4886,In_2518,In_2531);
nor U4887 (N_4887,In_1899,In_816);
and U4888 (N_4888,In_1717,In_1680);
nor U4889 (N_4889,In_1262,In_753);
xnor U4890 (N_4890,In_2787,In_902);
nand U4891 (N_4891,In_748,In_2567);
xor U4892 (N_4892,In_221,In_2450);
nor U4893 (N_4893,In_1664,In_1447);
nor U4894 (N_4894,In_1166,In_287);
xnor U4895 (N_4895,In_2018,In_2827);
nand U4896 (N_4896,In_1009,In_100);
or U4897 (N_4897,In_660,In_2309);
or U4898 (N_4898,In_1667,In_2062);
xor U4899 (N_4899,In_1180,In_189);
xnor U4900 (N_4900,In_193,In_2048);
nand U4901 (N_4901,In_2251,In_33);
and U4902 (N_4902,In_223,In_1563);
and U4903 (N_4903,In_982,In_2805);
and U4904 (N_4904,In_2541,In_2423);
and U4905 (N_4905,In_2226,In_2980);
and U4906 (N_4906,In_995,In_644);
or U4907 (N_4907,In_2209,In_249);
and U4908 (N_4908,In_1039,In_637);
xor U4909 (N_4909,In_180,In_2455);
and U4910 (N_4910,In_170,In_1060);
nor U4911 (N_4911,In_2604,In_2189);
and U4912 (N_4912,In_495,In_2416);
nor U4913 (N_4913,In_1949,In_2847);
nor U4914 (N_4914,In_77,In_2390);
xor U4915 (N_4915,In_937,In_2795);
or U4916 (N_4916,In_1874,In_2772);
and U4917 (N_4917,In_1199,In_695);
nand U4918 (N_4918,In_2022,In_254);
nor U4919 (N_4919,In_1879,In_1896);
nor U4920 (N_4920,In_2632,In_617);
and U4921 (N_4921,In_1112,In_2715);
and U4922 (N_4922,In_1458,In_63);
nand U4923 (N_4923,In_268,In_1581);
nor U4924 (N_4924,In_600,In_1514);
and U4925 (N_4925,In_2050,In_759);
and U4926 (N_4926,In_2559,In_2310);
and U4927 (N_4927,In_1671,In_2300);
or U4928 (N_4928,In_518,In_2939);
nor U4929 (N_4929,In_1728,In_2497);
or U4930 (N_4930,In_1498,In_2056);
or U4931 (N_4931,In_2181,In_367);
nand U4932 (N_4932,In_2879,In_1227);
and U4933 (N_4933,In_22,In_1869);
xor U4934 (N_4934,In_2932,In_1597);
xnor U4935 (N_4935,In_990,In_793);
or U4936 (N_4936,In_1774,In_2666);
nand U4937 (N_4937,In_2341,In_2054);
or U4938 (N_4938,In_1627,In_167);
or U4939 (N_4939,In_764,In_2435);
nand U4940 (N_4940,In_1812,In_277);
or U4941 (N_4941,In_2309,In_140);
nand U4942 (N_4942,In_1476,In_222);
nor U4943 (N_4943,In_741,In_2942);
nand U4944 (N_4944,In_34,In_715);
nand U4945 (N_4945,In_392,In_1539);
xnor U4946 (N_4946,In_2198,In_2066);
xnor U4947 (N_4947,In_1921,In_311);
or U4948 (N_4948,In_1399,In_2612);
or U4949 (N_4949,In_1833,In_1928);
nor U4950 (N_4950,In_2175,In_1508);
nor U4951 (N_4951,In_1400,In_1746);
nor U4952 (N_4952,In_608,In_578);
nand U4953 (N_4953,In_997,In_2799);
xnor U4954 (N_4954,In_1866,In_2409);
xor U4955 (N_4955,In_2518,In_1859);
nand U4956 (N_4956,In_1472,In_69);
nor U4957 (N_4957,In_1446,In_698);
nand U4958 (N_4958,In_2774,In_231);
nand U4959 (N_4959,In_371,In_1353);
nor U4960 (N_4960,In_1503,In_472);
and U4961 (N_4961,In_2606,In_327);
nand U4962 (N_4962,In_1706,In_1474);
nand U4963 (N_4963,In_807,In_2490);
nand U4964 (N_4964,In_33,In_223);
xor U4965 (N_4965,In_1768,In_45);
xor U4966 (N_4966,In_2467,In_1039);
nand U4967 (N_4967,In_1992,In_2273);
nand U4968 (N_4968,In_1806,In_1421);
xor U4969 (N_4969,In_2801,In_547);
nor U4970 (N_4970,In_2368,In_872);
and U4971 (N_4971,In_2040,In_1400);
nand U4972 (N_4972,In_1474,In_1825);
nor U4973 (N_4973,In_919,In_1221);
nand U4974 (N_4974,In_2594,In_1570);
nand U4975 (N_4975,In_445,In_2060);
and U4976 (N_4976,In_2258,In_2252);
nand U4977 (N_4977,In_1870,In_444);
xor U4978 (N_4978,In_1970,In_1392);
and U4979 (N_4979,In_2650,In_1825);
or U4980 (N_4980,In_206,In_74);
nor U4981 (N_4981,In_1833,In_206);
and U4982 (N_4982,In_239,In_2901);
or U4983 (N_4983,In_1223,In_68);
nand U4984 (N_4984,In_2468,In_1799);
xnor U4985 (N_4985,In_1547,In_426);
nor U4986 (N_4986,In_1676,In_1314);
nor U4987 (N_4987,In_77,In_2908);
or U4988 (N_4988,In_1886,In_418);
xnor U4989 (N_4989,In_212,In_985);
or U4990 (N_4990,In_1906,In_2674);
or U4991 (N_4991,In_2420,In_124);
nor U4992 (N_4992,In_1215,In_1624);
or U4993 (N_4993,In_680,In_427);
or U4994 (N_4994,In_2982,In_1131);
and U4995 (N_4995,In_1490,In_1245);
xor U4996 (N_4996,In_123,In_1484);
nor U4997 (N_4997,In_1330,In_273);
nor U4998 (N_4998,In_1385,In_1908);
nand U4999 (N_4999,In_665,In_37);
nor U5000 (N_5000,In_1654,In_447);
nand U5001 (N_5001,In_1833,In_1008);
or U5002 (N_5002,In_981,In_637);
or U5003 (N_5003,In_2605,In_789);
nor U5004 (N_5004,In_1355,In_225);
nor U5005 (N_5005,In_2493,In_2320);
nor U5006 (N_5006,In_1378,In_856);
and U5007 (N_5007,In_2911,In_1739);
xnor U5008 (N_5008,In_1411,In_687);
nor U5009 (N_5009,In_2961,In_2060);
nand U5010 (N_5010,In_243,In_2499);
and U5011 (N_5011,In_1758,In_2744);
and U5012 (N_5012,In_2487,In_362);
or U5013 (N_5013,In_1187,In_2139);
xnor U5014 (N_5014,In_72,In_2814);
and U5015 (N_5015,In_954,In_2419);
xnor U5016 (N_5016,In_2250,In_2736);
and U5017 (N_5017,In_279,In_1713);
nor U5018 (N_5018,In_2159,In_734);
nand U5019 (N_5019,In_2566,In_848);
xor U5020 (N_5020,In_712,In_492);
nand U5021 (N_5021,In_2175,In_328);
xnor U5022 (N_5022,In_2109,In_539);
xor U5023 (N_5023,In_1048,In_2219);
nor U5024 (N_5024,In_1020,In_1178);
nor U5025 (N_5025,In_919,In_1000);
and U5026 (N_5026,In_2550,In_1296);
nor U5027 (N_5027,In_1802,In_1492);
nand U5028 (N_5028,In_619,In_2253);
xnor U5029 (N_5029,In_164,In_2705);
and U5030 (N_5030,In_997,In_2955);
and U5031 (N_5031,In_1529,In_2238);
nor U5032 (N_5032,In_1220,In_505);
xor U5033 (N_5033,In_1514,In_909);
nor U5034 (N_5034,In_2668,In_159);
and U5035 (N_5035,In_2637,In_2216);
and U5036 (N_5036,In_403,In_1323);
and U5037 (N_5037,In_24,In_977);
or U5038 (N_5038,In_1892,In_182);
xnor U5039 (N_5039,In_1525,In_28);
nor U5040 (N_5040,In_636,In_1662);
nand U5041 (N_5041,In_2143,In_2639);
or U5042 (N_5042,In_502,In_1718);
xor U5043 (N_5043,In_375,In_964);
nand U5044 (N_5044,In_679,In_87);
nor U5045 (N_5045,In_1512,In_468);
nand U5046 (N_5046,In_2192,In_430);
nor U5047 (N_5047,In_53,In_388);
nand U5048 (N_5048,In_1319,In_1633);
or U5049 (N_5049,In_1600,In_2558);
and U5050 (N_5050,In_2745,In_326);
and U5051 (N_5051,In_1876,In_812);
nor U5052 (N_5052,In_2321,In_450);
nand U5053 (N_5053,In_1811,In_775);
nand U5054 (N_5054,In_2655,In_1732);
or U5055 (N_5055,In_583,In_1961);
and U5056 (N_5056,In_2289,In_1984);
xnor U5057 (N_5057,In_103,In_963);
and U5058 (N_5058,In_803,In_129);
xor U5059 (N_5059,In_2505,In_2355);
xnor U5060 (N_5060,In_80,In_1244);
nand U5061 (N_5061,In_1072,In_2030);
and U5062 (N_5062,In_2244,In_73);
nor U5063 (N_5063,In_301,In_730);
nand U5064 (N_5064,In_2485,In_2180);
xor U5065 (N_5065,In_2445,In_1110);
nor U5066 (N_5066,In_1533,In_1104);
nand U5067 (N_5067,In_553,In_2841);
or U5068 (N_5068,In_949,In_673);
or U5069 (N_5069,In_1359,In_442);
xor U5070 (N_5070,In_2438,In_509);
and U5071 (N_5071,In_775,In_2948);
nand U5072 (N_5072,In_1339,In_1647);
nor U5073 (N_5073,In_752,In_2126);
and U5074 (N_5074,In_2558,In_1221);
or U5075 (N_5075,In_2325,In_2039);
nand U5076 (N_5076,In_1627,In_2868);
and U5077 (N_5077,In_75,In_1404);
xnor U5078 (N_5078,In_109,In_2855);
or U5079 (N_5079,In_38,In_1968);
nor U5080 (N_5080,In_1211,In_656);
xor U5081 (N_5081,In_2559,In_727);
or U5082 (N_5082,In_2642,In_2912);
and U5083 (N_5083,In_1447,In_209);
nor U5084 (N_5084,In_1313,In_1653);
xnor U5085 (N_5085,In_191,In_1630);
xor U5086 (N_5086,In_1034,In_2088);
nand U5087 (N_5087,In_2294,In_2827);
xor U5088 (N_5088,In_535,In_174);
or U5089 (N_5089,In_1836,In_2180);
or U5090 (N_5090,In_214,In_2697);
or U5091 (N_5091,In_2601,In_709);
xor U5092 (N_5092,In_1509,In_1695);
xor U5093 (N_5093,In_2327,In_1881);
nand U5094 (N_5094,In_1446,In_2033);
and U5095 (N_5095,In_2368,In_1415);
nand U5096 (N_5096,In_1000,In_397);
or U5097 (N_5097,In_438,In_2803);
nor U5098 (N_5098,In_1488,In_1995);
and U5099 (N_5099,In_351,In_2459);
nand U5100 (N_5100,In_1662,In_1399);
and U5101 (N_5101,In_2346,In_393);
nand U5102 (N_5102,In_456,In_2422);
nor U5103 (N_5103,In_2906,In_2108);
xor U5104 (N_5104,In_1593,In_1811);
or U5105 (N_5105,In_1754,In_309);
or U5106 (N_5106,In_945,In_1427);
nor U5107 (N_5107,In_2929,In_179);
nor U5108 (N_5108,In_2904,In_2161);
and U5109 (N_5109,In_1016,In_2569);
nand U5110 (N_5110,In_2065,In_2684);
and U5111 (N_5111,In_1904,In_913);
nor U5112 (N_5112,In_362,In_1163);
and U5113 (N_5113,In_1634,In_2089);
xor U5114 (N_5114,In_2752,In_1071);
nor U5115 (N_5115,In_2619,In_73);
nand U5116 (N_5116,In_639,In_2695);
and U5117 (N_5117,In_224,In_520);
nand U5118 (N_5118,In_633,In_1002);
and U5119 (N_5119,In_717,In_405);
or U5120 (N_5120,In_2581,In_868);
nand U5121 (N_5121,In_2412,In_2743);
nand U5122 (N_5122,In_2434,In_2204);
xor U5123 (N_5123,In_1144,In_1922);
nor U5124 (N_5124,In_1658,In_1461);
or U5125 (N_5125,In_834,In_2725);
xnor U5126 (N_5126,In_2041,In_1952);
and U5127 (N_5127,In_987,In_2723);
and U5128 (N_5128,In_941,In_818);
or U5129 (N_5129,In_2828,In_2741);
xnor U5130 (N_5130,In_574,In_1429);
and U5131 (N_5131,In_2396,In_855);
and U5132 (N_5132,In_965,In_1542);
and U5133 (N_5133,In_2733,In_1201);
nand U5134 (N_5134,In_1567,In_515);
or U5135 (N_5135,In_1176,In_68);
or U5136 (N_5136,In_2758,In_1537);
nand U5137 (N_5137,In_1099,In_2688);
and U5138 (N_5138,In_1427,In_1956);
nand U5139 (N_5139,In_510,In_507);
xor U5140 (N_5140,In_2036,In_1340);
and U5141 (N_5141,In_2267,In_2190);
nor U5142 (N_5142,In_78,In_2089);
nor U5143 (N_5143,In_2599,In_2850);
nor U5144 (N_5144,In_457,In_2075);
nand U5145 (N_5145,In_2733,In_1452);
or U5146 (N_5146,In_2146,In_1636);
xnor U5147 (N_5147,In_1652,In_754);
nor U5148 (N_5148,In_1984,In_1169);
nand U5149 (N_5149,In_248,In_1367);
and U5150 (N_5150,In_1794,In_2555);
nor U5151 (N_5151,In_1518,In_716);
nor U5152 (N_5152,In_1239,In_2496);
xor U5153 (N_5153,In_562,In_37);
and U5154 (N_5154,In_2388,In_271);
nand U5155 (N_5155,In_2503,In_323);
xnor U5156 (N_5156,In_1946,In_10);
nor U5157 (N_5157,In_2370,In_1855);
nor U5158 (N_5158,In_2601,In_745);
nand U5159 (N_5159,In_1026,In_9);
or U5160 (N_5160,In_1712,In_2609);
xor U5161 (N_5161,In_1075,In_2866);
nand U5162 (N_5162,In_81,In_1106);
and U5163 (N_5163,In_1115,In_304);
nand U5164 (N_5164,In_629,In_2215);
and U5165 (N_5165,In_578,In_1032);
or U5166 (N_5166,In_140,In_1983);
xor U5167 (N_5167,In_2196,In_1819);
or U5168 (N_5168,In_940,In_1195);
or U5169 (N_5169,In_222,In_2832);
and U5170 (N_5170,In_287,In_2214);
and U5171 (N_5171,In_2607,In_926);
nor U5172 (N_5172,In_2074,In_2052);
xnor U5173 (N_5173,In_1660,In_2154);
nor U5174 (N_5174,In_2936,In_2391);
nor U5175 (N_5175,In_2805,In_197);
nor U5176 (N_5176,In_1835,In_2818);
xor U5177 (N_5177,In_2923,In_423);
xor U5178 (N_5178,In_1660,In_784);
nor U5179 (N_5179,In_183,In_2094);
xor U5180 (N_5180,In_1510,In_1255);
or U5181 (N_5181,In_1356,In_734);
or U5182 (N_5182,In_2218,In_906);
nor U5183 (N_5183,In_574,In_712);
nor U5184 (N_5184,In_2026,In_50);
xor U5185 (N_5185,In_641,In_2246);
nand U5186 (N_5186,In_98,In_1261);
or U5187 (N_5187,In_1062,In_1164);
and U5188 (N_5188,In_667,In_2764);
nor U5189 (N_5189,In_1157,In_1021);
nand U5190 (N_5190,In_785,In_1548);
nor U5191 (N_5191,In_2147,In_1348);
nand U5192 (N_5192,In_2536,In_2789);
nor U5193 (N_5193,In_268,In_778);
xnor U5194 (N_5194,In_693,In_2852);
nand U5195 (N_5195,In_2581,In_1308);
nor U5196 (N_5196,In_1206,In_78);
and U5197 (N_5197,In_253,In_41);
nor U5198 (N_5198,In_2767,In_2829);
and U5199 (N_5199,In_1450,In_1440);
xnor U5200 (N_5200,In_2289,In_1546);
or U5201 (N_5201,In_2515,In_269);
and U5202 (N_5202,In_2340,In_2517);
xnor U5203 (N_5203,In_41,In_2891);
or U5204 (N_5204,In_2589,In_2282);
or U5205 (N_5205,In_2830,In_1286);
and U5206 (N_5206,In_1939,In_1819);
and U5207 (N_5207,In_776,In_1788);
nor U5208 (N_5208,In_2563,In_689);
xnor U5209 (N_5209,In_1572,In_2879);
nand U5210 (N_5210,In_2066,In_198);
or U5211 (N_5211,In_2244,In_1711);
nor U5212 (N_5212,In_1431,In_300);
and U5213 (N_5213,In_212,In_1599);
xnor U5214 (N_5214,In_1764,In_663);
nand U5215 (N_5215,In_2643,In_1637);
and U5216 (N_5216,In_1847,In_2358);
nand U5217 (N_5217,In_2048,In_1904);
nor U5218 (N_5218,In_1934,In_2954);
nor U5219 (N_5219,In_1433,In_818);
nor U5220 (N_5220,In_1084,In_2256);
and U5221 (N_5221,In_473,In_791);
nor U5222 (N_5222,In_308,In_1250);
xnor U5223 (N_5223,In_1935,In_1671);
or U5224 (N_5224,In_1717,In_2127);
or U5225 (N_5225,In_2085,In_1805);
and U5226 (N_5226,In_2075,In_421);
nor U5227 (N_5227,In_719,In_295);
nand U5228 (N_5228,In_647,In_691);
or U5229 (N_5229,In_2125,In_459);
xnor U5230 (N_5230,In_1286,In_1359);
and U5231 (N_5231,In_1864,In_2400);
nor U5232 (N_5232,In_2153,In_1600);
nand U5233 (N_5233,In_1570,In_466);
nand U5234 (N_5234,In_1007,In_2612);
and U5235 (N_5235,In_1996,In_2153);
or U5236 (N_5236,In_984,In_2177);
or U5237 (N_5237,In_730,In_460);
nand U5238 (N_5238,In_2344,In_747);
or U5239 (N_5239,In_2666,In_86);
xnor U5240 (N_5240,In_2818,In_1481);
and U5241 (N_5241,In_1757,In_2193);
or U5242 (N_5242,In_2124,In_2063);
and U5243 (N_5243,In_1073,In_235);
or U5244 (N_5244,In_346,In_2873);
xor U5245 (N_5245,In_194,In_1237);
and U5246 (N_5246,In_935,In_2674);
xnor U5247 (N_5247,In_2583,In_2912);
xnor U5248 (N_5248,In_117,In_1611);
xor U5249 (N_5249,In_2490,In_225);
xnor U5250 (N_5250,In_714,In_2199);
nand U5251 (N_5251,In_1808,In_866);
or U5252 (N_5252,In_2157,In_2166);
nand U5253 (N_5253,In_1400,In_1936);
nand U5254 (N_5254,In_568,In_2018);
nand U5255 (N_5255,In_2890,In_1181);
nor U5256 (N_5256,In_135,In_2327);
nand U5257 (N_5257,In_359,In_1818);
or U5258 (N_5258,In_2341,In_2778);
xnor U5259 (N_5259,In_2825,In_2168);
nand U5260 (N_5260,In_1899,In_2055);
nor U5261 (N_5261,In_1663,In_1280);
xnor U5262 (N_5262,In_1508,In_1981);
xnor U5263 (N_5263,In_2223,In_368);
nor U5264 (N_5264,In_2047,In_2014);
nor U5265 (N_5265,In_2698,In_2457);
and U5266 (N_5266,In_867,In_413);
and U5267 (N_5267,In_1602,In_2163);
xnor U5268 (N_5268,In_952,In_2959);
nor U5269 (N_5269,In_2740,In_716);
xor U5270 (N_5270,In_1726,In_514);
or U5271 (N_5271,In_2883,In_2932);
nand U5272 (N_5272,In_1008,In_528);
nor U5273 (N_5273,In_2101,In_701);
nand U5274 (N_5274,In_1870,In_2305);
nor U5275 (N_5275,In_2505,In_529);
nor U5276 (N_5276,In_1309,In_2195);
and U5277 (N_5277,In_2288,In_1674);
and U5278 (N_5278,In_1592,In_821);
or U5279 (N_5279,In_796,In_2601);
or U5280 (N_5280,In_2602,In_1333);
nor U5281 (N_5281,In_1862,In_634);
and U5282 (N_5282,In_2546,In_201);
or U5283 (N_5283,In_2840,In_340);
nand U5284 (N_5284,In_836,In_783);
xor U5285 (N_5285,In_783,In_534);
xor U5286 (N_5286,In_1556,In_2609);
nand U5287 (N_5287,In_2047,In_2764);
nand U5288 (N_5288,In_48,In_2766);
nor U5289 (N_5289,In_1528,In_827);
nand U5290 (N_5290,In_226,In_1305);
nor U5291 (N_5291,In_1850,In_776);
and U5292 (N_5292,In_402,In_2581);
nand U5293 (N_5293,In_1884,In_748);
and U5294 (N_5294,In_506,In_803);
xor U5295 (N_5295,In_1477,In_1851);
nand U5296 (N_5296,In_1709,In_1231);
nor U5297 (N_5297,In_1705,In_1711);
or U5298 (N_5298,In_794,In_2990);
xnor U5299 (N_5299,In_2169,In_1441);
and U5300 (N_5300,In_1579,In_767);
or U5301 (N_5301,In_1868,In_1841);
nor U5302 (N_5302,In_782,In_2790);
nor U5303 (N_5303,In_2124,In_1490);
and U5304 (N_5304,In_1428,In_738);
xnor U5305 (N_5305,In_677,In_872);
nand U5306 (N_5306,In_492,In_2298);
nand U5307 (N_5307,In_858,In_2357);
nand U5308 (N_5308,In_2845,In_307);
nand U5309 (N_5309,In_2753,In_757);
xor U5310 (N_5310,In_1871,In_803);
and U5311 (N_5311,In_2349,In_2558);
nand U5312 (N_5312,In_50,In_1808);
xor U5313 (N_5313,In_2132,In_461);
xnor U5314 (N_5314,In_2463,In_1553);
and U5315 (N_5315,In_609,In_2293);
and U5316 (N_5316,In_635,In_2171);
xnor U5317 (N_5317,In_1701,In_567);
or U5318 (N_5318,In_2550,In_1969);
nand U5319 (N_5319,In_2500,In_44);
nand U5320 (N_5320,In_2845,In_2167);
xnor U5321 (N_5321,In_268,In_2756);
xor U5322 (N_5322,In_992,In_2026);
xnor U5323 (N_5323,In_2237,In_2767);
and U5324 (N_5324,In_1594,In_2365);
nand U5325 (N_5325,In_551,In_1027);
xor U5326 (N_5326,In_1567,In_2368);
xnor U5327 (N_5327,In_1415,In_2141);
or U5328 (N_5328,In_1361,In_1234);
nor U5329 (N_5329,In_1613,In_2727);
nand U5330 (N_5330,In_2388,In_2798);
nand U5331 (N_5331,In_2316,In_2992);
and U5332 (N_5332,In_2767,In_84);
nor U5333 (N_5333,In_2214,In_2981);
nand U5334 (N_5334,In_2834,In_1172);
nor U5335 (N_5335,In_2765,In_2301);
nor U5336 (N_5336,In_839,In_2387);
xnor U5337 (N_5337,In_2733,In_2071);
or U5338 (N_5338,In_2271,In_1386);
or U5339 (N_5339,In_819,In_2320);
or U5340 (N_5340,In_2813,In_1298);
nor U5341 (N_5341,In_1639,In_1755);
and U5342 (N_5342,In_466,In_316);
nor U5343 (N_5343,In_2486,In_1982);
or U5344 (N_5344,In_2688,In_2424);
xnor U5345 (N_5345,In_426,In_2412);
nor U5346 (N_5346,In_2721,In_2753);
and U5347 (N_5347,In_194,In_2900);
nand U5348 (N_5348,In_2725,In_1784);
and U5349 (N_5349,In_521,In_1306);
and U5350 (N_5350,In_421,In_605);
nor U5351 (N_5351,In_1728,In_2820);
or U5352 (N_5352,In_1056,In_529);
or U5353 (N_5353,In_420,In_2569);
nor U5354 (N_5354,In_1706,In_1100);
nand U5355 (N_5355,In_2022,In_836);
nand U5356 (N_5356,In_705,In_1950);
nor U5357 (N_5357,In_1804,In_1799);
and U5358 (N_5358,In_742,In_1533);
nor U5359 (N_5359,In_2151,In_677);
nor U5360 (N_5360,In_2195,In_844);
nor U5361 (N_5361,In_1448,In_774);
nor U5362 (N_5362,In_2683,In_2123);
xnor U5363 (N_5363,In_232,In_1097);
nand U5364 (N_5364,In_2357,In_2147);
nand U5365 (N_5365,In_306,In_415);
nand U5366 (N_5366,In_1033,In_1012);
nor U5367 (N_5367,In_1949,In_956);
and U5368 (N_5368,In_2444,In_2669);
nor U5369 (N_5369,In_951,In_754);
nor U5370 (N_5370,In_642,In_860);
nand U5371 (N_5371,In_743,In_1773);
or U5372 (N_5372,In_1795,In_117);
and U5373 (N_5373,In_1984,In_1523);
xor U5374 (N_5374,In_2980,In_1517);
or U5375 (N_5375,In_1249,In_2540);
and U5376 (N_5376,In_2686,In_2559);
xnor U5377 (N_5377,In_1482,In_1417);
nor U5378 (N_5378,In_173,In_1366);
nor U5379 (N_5379,In_867,In_969);
and U5380 (N_5380,In_666,In_1213);
nor U5381 (N_5381,In_2893,In_2357);
or U5382 (N_5382,In_1504,In_2146);
nand U5383 (N_5383,In_1965,In_2417);
or U5384 (N_5384,In_168,In_2145);
nand U5385 (N_5385,In_93,In_1071);
or U5386 (N_5386,In_2834,In_266);
nand U5387 (N_5387,In_79,In_2004);
nand U5388 (N_5388,In_1950,In_2548);
and U5389 (N_5389,In_1726,In_2959);
and U5390 (N_5390,In_1568,In_1070);
xnor U5391 (N_5391,In_1137,In_2339);
nand U5392 (N_5392,In_2861,In_2326);
or U5393 (N_5393,In_413,In_2389);
nand U5394 (N_5394,In_2442,In_2522);
and U5395 (N_5395,In_973,In_1082);
xnor U5396 (N_5396,In_2535,In_1380);
and U5397 (N_5397,In_543,In_455);
xor U5398 (N_5398,In_1076,In_1119);
xnor U5399 (N_5399,In_2567,In_2864);
nand U5400 (N_5400,In_2689,In_1309);
or U5401 (N_5401,In_606,In_194);
and U5402 (N_5402,In_766,In_1836);
nand U5403 (N_5403,In_1762,In_2218);
nor U5404 (N_5404,In_2994,In_1949);
nor U5405 (N_5405,In_2499,In_1638);
nor U5406 (N_5406,In_2883,In_2648);
nand U5407 (N_5407,In_2466,In_1884);
and U5408 (N_5408,In_1345,In_2824);
xnor U5409 (N_5409,In_2134,In_1937);
nand U5410 (N_5410,In_344,In_1817);
or U5411 (N_5411,In_2205,In_2285);
and U5412 (N_5412,In_938,In_2148);
nor U5413 (N_5413,In_1427,In_264);
or U5414 (N_5414,In_1715,In_2363);
nor U5415 (N_5415,In_1390,In_2101);
nor U5416 (N_5416,In_1484,In_1419);
nor U5417 (N_5417,In_947,In_271);
xnor U5418 (N_5418,In_544,In_1142);
and U5419 (N_5419,In_1612,In_1530);
or U5420 (N_5420,In_2300,In_777);
xnor U5421 (N_5421,In_1911,In_1280);
nor U5422 (N_5422,In_1242,In_2290);
nor U5423 (N_5423,In_2001,In_1846);
nand U5424 (N_5424,In_249,In_117);
nor U5425 (N_5425,In_290,In_1142);
or U5426 (N_5426,In_2114,In_2250);
nor U5427 (N_5427,In_1588,In_1113);
or U5428 (N_5428,In_2497,In_2033);
nand U5429 (N_5429,In_531,In_1695);
xor U5430 (N_5430,In_319,In_1422);
nor U5431 (N_5431,In_2208,In_1323);
xnor U5432 (N_5432,In_90,In_2258);
xor U5433 (N_5433,In_157,In_2853);
and U5434 (N_5434,In_574,In_1124);
nand U5435 (N_5435,In_1904,In_2492);
nor U5436 (N_5436,In_1644,In_2638);
nor U5437 (N_5437,In_477,In_2890);
nand U5438 (N_5438,In_1251,In_183);
or U5439 (N_5439,In_1336,In_1768);
nor U5440 (N_5440,In_1708,In_477);
nor U5441 (N_5441,In_444,In_1946);
nand U5442 (N_5442,In_817,In_1781);
or U5443 (N_5443,In_2128,In_2997);
nand U5444 (N_5444,In_2550,In_1674);
or U5445 (N_5445,In_1274,In_2156);
nand U5446 (N_5446,In_1336,In_1058);
nand U5447 (N_5447,In_1207,In_192);
nand U5448 (N_5448,In_2705,In_896);
or U5449 (N_5449,In_1600,In_749);
nor U5450 (N_5450,In_2590,In_1710);
nor U5451 (N_5451,In_1950,In_764);
or U5452 (N_5452,In_603,In_1507);
or U5453 (N_5453,In_986,In_2587);
or U5454 (N_5454,In_271,In_2199);
nor U5455 (N_5455,In_2519,In_1344);
xor U5456 (N_5456,In_2127,In_1183);
nand U5457 (N_5457,In_88,In_1127);
xor U5458 (N_5458,In_1785,In_1615);
nand U5459 (N_5459,In_2578,In_308);
nor U5460 (N_5460,In_2200,In_1967);
nor U5461 (N_5461,In_107,In_1730);
or U5462 (N_5462,In_2101,In_528);
or U5463 (N_5463,In_386,In_523);
or U5464 (N_5464,In_357,In_2604);
or U5465 (N_5465,In_2905,In_69);
and U5466 (N_5466,In_678,In_1685);
and U5467 (N_5467,In_2403,In_759);
nor U5468 (N_5468,In_1781,In_524);
xnor U5469 (N_5469,In_1060,In_2017);
nand U5470 (N_5470,In_473,In_2494);
nand U5471 (N_5471,In_38,In_2957);
or U5472 (N_5472,In_2674,In_2629);
xor U5473 (N_5473,In_328,In_2664);
xnor U5474 (N_5474,In_2655,In_2702);
nand U5475 (N_5475,In_825,In_1051);
or U5476 (N_5476,In_2561,In_1151);
nor U5477 (N_5477,In_261,In_2163);
and U5478 (N_5478,In_627,In_1547);
nand U5479 (N_5479,In_1563,In_2561);
and U5480 (N_5480,In_913,In_170);
and U5481 (N_5481,In_2244,In_2637);
nand U5482 (N_5482,In_1119,In_930);
xor U5483 (N_5483,In_2768,In_2215);
and U5484 (N_5484,In_45,In_1115);
xor U5485 (N_5485,In_390,In_1201);
and U5486 (N_5486,In_2017,In_2026);
nand U5487 (N_5487,In_1609,In_1274);
and U5488 (N_5488,In_1615,In_1754);
xor U5489 (N_5489,In_243,In_1518);
nor U5490 (N_5490,In_2786,In_2090);
nor U5491 (N_5491,In_1624,In_2164);
nor U5492 (N_5492,In_1431,In_1101);
nand U5493 (N_5493,In_493,In_209);
and U5494 (N_5494,In_585,In_119);
or U5495 (N_5495,In_1773,In_2537);
or U5496 (N_5496,In_1705,In_1493);
or U5497 (N_5497,In_934,In_1363);
xnor U5498 (N_5498,In_1215,In_2424);
or U5499 (N_5499,In_2756,In_2961);
and U5500 (N_5500,In_304,In_1817);
xnor U5501 (N_5501,In_2891,In_2800);
xor U5502 (N_5502,In_1778,In_2392);
xnor U5503 (N_5503,In_2527,In_1783);
xor U5504 (N_5504,In_862,In_403);
nor U5505 (N_5505,In_611,In_2970);
nor U5506 (N_5506,In_2348,In_1674);
and U5507 (N_5507,In_2879,In_2635);
or U5508 (N_5508,In_2092,In_830);
xnor U5509 (N_5509,In_287,In_38);
and U5510 (N_5510,In_1953,In_3);
nor U5511 (N_5511,In_2746,In_2843);
or U5512 (N_5512,In_1447,In_81);
nand U5513 (N_5513,In_368,In_1475);
xor U5514 (N_5514,In_1141,In_586);
nand U5515 (N_5515,In_2540,In_1932);
xnor U5516 (N_5516,In_1852,In_2242);
nand U5517 (N_5517,In_983,In_644);
nor U5518 (N_5518,In_146,In_2314);
xor U5519 (N_5519,In_2200,In_2448);
xor U5520 (N_5520,In_2421,In_136);
xnor U5521 (N_5521,In_535,In_2582);
and U5522 (N_5522,In_2002,In_1873);
and U5523 (N_5523,In_1281,In_954);
nor U5524 (N_5524,In_2749,In_1584);
and U5525 (N_5525,In_306,In_2219);
or U5526 (N_5526,In_470,In_2205);
nand U5527 (N_5527,In_2792,In_1965);
and U5528 (N_5528,In_1958,In_1453);
nor U5529 (N_5529,In_263,In_237);
nor U5530 (N_5530,In_1846,In_1531);
nor U5531 (N_5531,In_1747,In_1428);
nor U5532 (N_5532,In_27,In_830);
xnor U5533 (N_5533,In_1528,In_1419);
nand U5534 (N_5534,In_368,In_2090);
or U5535 (N_5535,In_2456,In_1347);
xor U5536 (N_5536,In_363,In_2467);
xor U5537 (N_5537,In_385,In_2144);
nand U5538 (N_5538,In_743,In_2016);
and U5539 (N_5539,In_2899,In_549);
nand U5540 (N_5540,In_1375,In_1488);
nor U5541 (N_5541,In_2342,In_496);
and U5542 (N_5542,In_2193,In_1591);
nand U5543 (N_5543,In_1503,In_435);
nand U5544 (N_5544,In_1281,In_27);
and U5545 (N_5545,In_1049,In_111);
or U5546 (N_5546,In_2565,In_204);
nor U5547 (N_5547,In_2645,In_2416);
and U5548 (N_5548,In_2363,In_873);
nand U5549 (N_5549,In_1835,In_2888);
and U5550 (N_5550,In_11,In_515);
nor U5551 (N_5551,In_1129,In_1387);
nor U5552 (N_5552,In_261,In_1106);
and U5553 (N_5553,In_515,In_2742);
nand U5554 (N_5554,In_1750,In_46);
or U5555 (N_5555,In_1655,In_2609);
xnor U5556 (N_5556,In_198,In_1280);
or U5557 (N_5557,In_2608,In_2850);
and U5558 (N_5558,In_2636,In_1082);
and U5559 (N_5559,In_2809,In_2422);
nand U5560 (N_5560,In_2908,In_1498);
xor U5561 (N_5561,In_562,In_377);
nor U5562 (N_5562,In_2337,In_200);
nor U5563 (N_5563,In_894,In_889);
nand U5564 (N_5564,In_145,In_291);
xor U5565 (N_5565,In_1155,In_2820);
or U5566 (N_5566,In_2692,In_1886);
xor U5567 (N_5567,In_924,In_2839);
nand U5568 (N_5568,In_2379,In_1940);
and U5569 (N_5569,In_1333,In_1345);
nand U5570 (N_5570,In_1418,In_647);
or U5571 (N_5571,In_2051,In_75);
and U5572 (N_5572,In_2843,In_1388);
or U5573 (N_5573,In_2875,In_1313);
nor U5574 (N_5574,In_1285,In_2439);
xnor U5575 (N_5575,In_1794,In_2899);
nor U5576 (N_5576,In_524,In_2786);
and U5577 (N_5577,In_564,In_1378);
xnor U5578 (N_5578,In_722,In_150);
xor U5579 (N_5579,In_71,In_2315);
nor U5580 (N_5580,In_2379,In_2711);
xor U5581 (N_5581,In_172,In_1661);
xnor U5582 (N_5582,In_380,In_2935);
nand U5583 (N_5583,In_605,In_2590);
xnor U5584 (N_5584,In_1653,In_2984);
xor U5585 (N_5585,In_489,In_558);
xor U5586 (N_5586,In_1006,In_1200);
xnor U5587 (N_5587,In_604,In_2220);
or U5588 (N_5588,In_2823,In_2814);
xor U5589 (N_5589,In_1785,In_1165);
and U5590 (N_5590,In_2756,In_15);
nand U5591 (N_5591,In_2356,In_1498);
and U5592 (N_5592,In_1807,In_2068);
and U5593 (N_5593,In_936,In_731);
or U5594 (N_5594,In_941,In_2484);
or U5595 (N_5595,In_2454,In_1366);
nand U5596 (N_5596,In_2741,In_820);
and U5597 (N_5597,In_2911,In_919);
nor U5598 (N_5598,In_1126,In_1598);
or U5599 (N_5599,In_1415,In_1533);
or U5600 (N_5600,In_462,In_2338);
nor U5601 (N_5601,In_2477,In_1959);
nor U5602 (N_5602,In_1159,In_2147);
nor U5603 (N_5603,In_954,In_667);
nand U5604 (N_5604,In_2008,In_1452);
or U5605 (N_5605,In_1050,In_1202);
nor U5606 (N_5606,In_1113,In_146);
and U5607 (N_5607,In_1064,In_1247);
nor U5608 (N_5608,In_2885,In_1667);
or U5609 (N_5609,In_2492,In_2806);
nand U5610 (N_5610,In_2825,In_2332);
xnor U5611 (N_5611,In_2871,In_1027);
and U5612 (N_5612,In_2117,In_2627);
nand U5613 (N_5613,In_861,In_176);
or U5614 (N_5614,In_894,In_2134);
nand U5615 (N_5615,In_2238,In_1748);
or U5616 (N_5616,In_1302,In_1655);
xnor U5617 (N_5617,In_1190,In_894);
or U5618 (N_5618,In_298,In_2369);
nor U5619 (N_5619,In_278,In_1657);
nand U5620 (N_5620,In_122,In_350);
or U5621 (N_5621,In_540,In_854);
and U5622 (N_5622,In_2092,In_424);
nor U5623 (N_5623,In_1127,In_868);
nor U5624 (N_5624,In_2980,In_2985);
xor U5625 (N_5625,In_1542,In_2271);
xnor U5626 (N_5626,In_225,In_952);
and U5627 (N_5627,In_2782,In_1912);
nor U5628 (N_5628,In_921,In_1770);
nand U5629 (N_5629,In_629,In_1396);
xor U5630 (N_5630,In_2921,In_2641);
xor U5631 (N_5631,In_662,In_2398);
nor U5632 (N_5632,In_1380,In_148);
or U5633 (N_5633,In_2568,In_1474);
nand U5634 (N_5634,In_258,In_1792);
or U5635 (N_5635,In_1570,In_647);
xor U5636 (N_5636,In_2045,In_1791);
xnor U5637 (N_5637,In_869,In_1320);
nand U5638 (N_5638,In_2507,In_2638);
xor U5639 (N_5639,In_1019,In_2431);
nor U5640 (N_5640,In_2723,In_1440);
xor U5641 (N_5641,In_1286,In_1600);
and U5642 (N_5642,In_2700,In_712);
nand U5643 (N_5643,In_1850,In_2790);
nor U5644 (N_5644,In_2353,In_571);
nor U5645 (N_5645,In_854,In_1380);
nor U5646 (N_5646,In_1090,In_1467);
nand U5647 (N_5647,In_1785,In_2665);
or U5648 (N_5648,In_1572,In_682);
and U5649 (N_5649,In_58,In_2344);
and U5650 (N_5650,In_1640,In_1681);
nor U5651 (N_5651,In_1899,In_2342);
or U5652 (N_5652,In_2001,In_2692);
nor U5653 (N_5653,In_1921,In_65);
and U5654 (N_5654,In_2337,In_683);
nor U5655 (N_5655,In_1928,In_2571);
nor U5656 (N_5656,In_8,In_2400);
nand U5657 (N_5657,In_871,In_694);
and U5658 (N_5658,In_768,In_816);
or U5659 (N_5659,In_852,In_1179);
nand U5660 (N_5660,In_1898,In_1970);
or U5661 (N_5661,In_807,In_2731);
or U5662 (N_5662,In_855,In_1236);
xor U5663 (N_5663,In_1979,In_582);
or U5664 (N_5664,In_22,In_1323);
nand U5665 (N_5665,In_984,In_2924);
nor U5666 (N_5666,In_1142,In_2411);
xor U5667 (N_5667,In_333,In_2252);
or U5668 (N_5668,In_161,In_335);
nand U5669 (N_5669,In_1585,In_1979);
nor U5670 (N_5670,In_2000,In_1457);
and U5671 (N_5671,In_2475,In_574);
nor U5672 (N_5672,In_928,In_2364);
or U5673 (N_5673,In_2453,In_386);
nand U5674 (N_5674,In_639,In_2394);
and U5675 (N_5675,In_118,In_1509);
xor U5676 (N_5676,In_2987,In_585);
xnor U5677 (N_5677,In_1773,In_1614);
or U5678 (N_5678,In_1932,In_113);
xor U5679 (N_5679,In_346,In_1870);
and U5680 (N_5680,In_2398,In_2518);
or U5681 (N_5681,In_1372,In_2354);
and U5682 (N_5682,In_286,In_444);
xnor U5683 (N_5683,In_2561,In_2432);
xnor U5684 (N_5684,In_2213,In_2257);
nand U5685 (N_5685,In_2395,In_527);
and U5686 (N_5686,In_2778,In_2651);
nand U5687 (N_5687,In_216,In_2690);
nand U5688 (N_5688,In_2620,In_354);
nand U5689 (N_5689,In_334,In_2432);
xor U5690 (N_5690,In_2399,In_119);
nand U5691 (N_5691,In_1476,In_2786);
and U5692 (N_5692,In_674,In_319);
xor U5693 (N_5693,In_2212,In_2686);
xnor U5694 (N_5694,In_988,In_754);
nand U5695 (N_5695,In_781,In_1504);
nor U5696 (N_5696,In_1267,In_135);
nor U5697 (N_5697,In_2955,In_2917);
nand U5698 (N_5698,In_1030,In_288);
and U5699 (N_5699,In_1316,In_1526);
and U5700 (N_5700,In_652,In_139);
nor U5701 (N_5701,In_2283,In_513);
nor U5702 (N_5702,In_1138,In_281);
and U5703 (N_5703,In_1157,In_2505);
or U5704 (N_5704,In_1648,In_2385);
and U5705 (N_5705,In_1928,In_1829);
or U5706 (N_5706,In_2259,In_22);
or U5707 (N_5707,In_1658,In_1902);
and U5708 (N_5708,In_174,In_2950);
and U5709 (N_5709,In_1291,In_2210);
or U5710 (N_5710,In_501,In_2096);
and U5711 (N_5711,In_1362,In_2710);
or U5712 (N_5712,In_1991,In_2976);
and U5713 (N_5713,In_2643,In_429);
xor U5714 (N_5714,In_913,In_2391);
nor U5715 (N_5715,In_2101,In_1395);
nor U5716 (N_5716,In_786,In_1952);
or U5717 (N_5717,In_2214,In_2331);
or U5718 (N_5718,In_1542,In_2682);
xnor U5719 (N_5719,In_1450,In_119);
nand U5720 (N_5720,In_2445,In_2061);
or U5721 (N_5721,In_1418,In_2935);
and U5722 (N_5722,In_558,In_2535);
xnor U5723 (N_5723,In_2113,In_2903);
nand U5724 (N_5724,In_1833,In_2206);
or U5725 (N_5725,In_2659,In_1123);
xnor U5726 (N_5726,In_593,In_1572);
or U5727 (N_5727,In_1064,In_228);
nand U5728 (N_5728,In_429,In_821);
nor U5729 (N_5729,In_1582,In_1756);
and U5730 (N_5730,In_2812,In_1168);
nor U5731 (N_5731,In_13,In_674);
and U5732 (N_5732,In_2004,In_2187);
or U5733 (N_5733,In_2680,In_1444);
xnor U5734 (N_5734,In_27,In_2090);
nand U5735 (N_5735,In_1013,In_1020);
nand U5736 (N_5736,In_527,In_907);
xnor U5737 (N_5737,In_1851,In_1927);
or U5738 (N_5738,In_938,In_1719);
nand U5739 (N_5739,In_698,In_401);
xor U5740 (N_5740,In_610,In_2329);
or U5741 (N_5741,In_759,In_1764);
and U5742 (N_5742,In_47,In_345);
nor U5743 (N_5743,In_2543,In_1034);
or U5744 (N_5744,In_53,In_147);
or U5745 (N_5745,In_2894,In_272);
nand U5746 (N_5746,In_669,In_2746);
or U5747 (N_5747,In_327,In_1017);
or U5748 (N_5748,In_73,In_2672);
xnor U5749 (N_5749,In_2092,In_2854);
and U5750 (N_5750,In_331,In_2240);
and U5751 (N_5751,In_51,In_2429);
nor U5752 (N_5752,In_2860,In_629);
nand U5753 (N_5753,In_2175,In_2249);
nand U5754 (N_5754,In_2014,In_2738);
and U5755 (N_5755,In_500,In_2963);
nor U5756 (N_5756,In_456,In_1254);
and U5757 (N_5757,In_2661,In_2591);
and U5758 (N_5758,In_212,In_928);
nor U5759 (N_5759,In_2741,In_2700);
and U5760 (N_5760,In_2224,In_1550);
xor U5761 (N_5761,In_1491,In_448);
and U5762 (N_5762,In_1718,In_2132);
xor U5763 (N_5763,In_539,In_1519);
nor U5764 (N_5764,In_185,In_1146);
xnor U5765 (N_5765,In_339,In_2658);
and U5766 (N_5766,In_2733,In_2629);
xor U5767 (N_5767,In_637,In_1315);
nand U5768 (N_5768,In_651,In_139);
nor U5769 (N_5769,In_1434,In_685);
nand U5770 (N_5770,In_703,In_2409);
and U5771 (N_5771,In_2114,In_2521);
and U5772 (N_5772,In_1796,In_2530);
xnor U5773 (N_5773,In_1047,In_2748);
nor U5774 (N_5774,In_413,In_499);
nor U5775 (N_5775,In_1986,In_1760);
or U5776 (N_5776,In_876,In_677);
nand U5777 (N_5777,In_1128,In_2656);
nand U5778 (N_5778,In_2765,In_2749);
nand U5779 (N_5779,In_1797,In_1263);
and U5780 (N_5780,In_985,In_281);
xor U5781 (N_5781,In_673,In_2607);
nand U5782 (N_5782,In_2314,In_813);
or U5783 (N_5783,In_296,In_983);
or U5784 (N_5784,In_1885,In_2951);
xnor U5785 (N_5785,In_2766,In_154);
and U5786 (N_5786,In_1335,In_1329);
or U5787 (N_5787,In_2528,In_1833);
nand U5788 (N_5788,In_1601,In_2308);
and U5789 (N_5789,In_2990,In_2444);
and U5790 (N_5790,In_844,In_439);
nor U5791 (N_5791,In_93,In_692);
xor U5792 (N_5792,In_1952,In_1663);
xor U5793 (N_5793,In_2237,In_2864);
nor U5794 (N_5794,In_2581,In_1359);
or U5795 (N_5795,In_1177,In_1664);
nor U5796 (N_5796,In_2952,In_577);
nor U5797 (N_5797,In_1214,In_58);
or U5798 (N_5798,In_2229,In_2573);
xor U5799 (N_5799,In_2401,In_1174);
nand U5800 (N_5800,In_1488,In_2535);
and U5801 (N_5801,In_1255,In_556);
nor U5802 (N_5802,In_1156,In_81);
xor U5803 (N_5803,In_459,In_2897);
and U5804 (N_5804,In_481,In_274);
or U5805 (N_5805,In_1107,In_2363);
xnor U5806 (N_5806,In_1695,In_1954);
or U5807 (N_5807,In_290,In_1334);
nand U5808 (N_5808,In_2823,In_2736);
xnor U5809 (N_5809,In_675,In_2118);
or U5810 (N_5810,In_2237,In_554);
nor U5811 (N_5811,In_2600,In_1408);
or U5812 (N_5812,In_908,In_2251);
and U5813 (N_5813,In_1838,In_786);
nand U5814 (N_5814,In_2004,In_2159);
or U5815 (N_5815,In_1906,In_2616);
nor U5816 (N_5816,In_1157,In_188);
xor U5817 (N_5817,In_935,In_418);
nor U5818 (N_5818,In_670,In_1019);
nand U5819 (N_5819,In_2147,In_199);
or U5820 (N_5820,In_167,In_1825);
or U5821 (N_5821,In_1502,In_2114);
xnor U5822 (N_5822,In_948,In_2385);
or U5823 (N_5823,In_1715,In_1420);
xnor U5824 (N_5824,In_2730,In_515);
xor U5825 (N_5825,In_1281,In_914);
nor U5826 (N_5826,In_2798,In_2606);
or U5827 (N_5827,In_2835,In_1774);
or U5828 (N_5828,In_2833,In_439);
nor U5829 (N_5829,In_1278,In_2755);
or U5830 (N_5830,In_2928,In_479);
nand U5831 (N_5831,In_1644,In_2894);
nand U5832 (N_5832,In_220,In_2381);
xnor U5833 (N_5833,In_2406,In_2857);
nand U5834 (N_5834,In_525,In_1717);
and U5835 (N_5835,In_2416,In_2573);
xor U5836 (N_5836,In_2083,In_2526);
and U5837 (N_5837,In_531,In_79);
or U5838 (N_5838,In_800,In_1125);
nand U5839 (N_5839,In_1510,In_1594);
and U5840 (N_5840,In_1412,In_46);
nor U5841 (N_5841,In_1315,In_2032);
and U5842 (N_5842,In_2203,In_1947);
xnor U5843 (N_5843,In_2201,In_992);
or U5844 (N_5844,In_1871,In_107);
nor U5845 (N_5845,In_2495,In_1374);
nand U5846 (N_5846,In_1528,In_728);
nand U5847 (N_5847,In_1391,In_1642);
nor U5848 (N_5848,In_2585,In_416);
and U5849 (N_5849,In_2323,In_2062);
nand U5850 (N_5850,In_1987,In_1326);
xnor U5851 (N_5851,In_91,In_1476);
xor U5852 (N_5852,In_319,In_639);
or U5853 (N_5853,In_2422,In_1885);
nor U5854 (N_5854,In_1538,In_2392);
and U5855 (N_5855,In_1715,In_1531);
and U5856 (N_5856,In_1471,In_2122);
nor U5857 (N_5857,In_424,In_408);
xor U5858 (N_5858,In_1500,In_435);
and U5859 (N_5859,In_1315,In_2938);
nand U5860 (N_5860,In_617,In_2489);
nor U5861 (N_5861,In_460,In_1096);
or U5862 (N_5862,In_2626,In_1764);
and U5863 (N_5863,In_2938,In_2043);
xnor U5864 (N_5864,In_920,In_622);
nor U5865 (N_5865,In_2987,In_858);
or U5866 (N_5866,In_1130,In_1940);
nor U5867 (N_5867,In_2768,In_1741);
or U5868 (N_5868,In_2231,In_557);
xnor U5869 (N_5869,In_1546,In_900);
nor U5870 (N_5870,In_1002,In_548);
xnor U5871 (N_5871,In_2450,In_693);
xor U5872 (N_5872,In_2197,In_2129);
nand U5873 (N_5873,In_358,In_567);
nor U5874 (N_5874,In_2198,In_1529);
xnor U5875 (N_5875,In_2533,In_341);
and U5876 (N_5876,In_1656,In_1864);
or U5877 (N_5877,In_690,In_2863);
xnor U5878 (N_5878,In_828,In_1798);
nor U5879 (N_5879,In_2215,In_2891);
or U5880 (N_5880,In_2400,In_1961);
nand U5881 (N_5881,In_1642,In_1720);
or U5882 (N_5882,In_1926,In_2389);
nand U5883 (N_5883,In_1965,In_998);
or U5884 (N_5884,In_749,In_389);
xor U5885 (N_5885,In_889,In_2801);
or U5886 (N_5886,In_2936,In_1198);
and U5887 (N_5887,In_1464,In_978);
nor U5888 (N_5888,In_1643,In_1758);
and U5889 (N_5889,In_2372,In_866);
nand U5890 (N_5890,In_1707,In_1679);
xor U5891 (N_5891,In_2290,In_1151);
nand U5892 (N_5892,In_1450,In_261);
or U5893 (N_5893,In_2876,In_359);
or U5894 (N_5894,In_196,In_776);
or U5895 (N_5895,In_1937,In_863);
and U5896 (N_5896,In_2344,In_372);
and U5897 (N_5897,In_2970,In_1079);
nand U5898 (N_5898,In_1962,In_2893);
and U5899 (N_5899,In_1075,In_68);
nor U5900 (N_5900,In_836,In_1982);
or U5901 (N_5901,In_460,In_508);
nand U5902 (N_5902,In_2448,In_1080);
and U5903 (N_5903,In_2547,In_2362);
or U5904 (N_5904,In_2543,In_2343);
nand U5905 (N_5905,In_2735,In_2418);
nand U5906 (N_5906,In_898,In_2116);
nor U5907 (N_5907,In_1487,In_2420);
nor U5908 (N_5908,In_2191,In_990);
or U5909 (N_5909,In_2402,In_1464);
xnor U5910 (N_5910,In_2993,In_1457);
and U5911 (N_5911,In_2445,In_1451);
nand U5912 (N_5912,In_2643,In_688);
nand U5913 (N_5913,In_1169,In_601);
or U5914 (N_5914,In_1410,In_1387);
xnor U5915 (N_5915,In_983,In_1139);
nor U5916 (N_5916,In_2162,In_540);
nor U5917 (N_5917,In_1156,In_2029);
nor U5918 (N_5918,In_571,In_2378);
or U5919 (N_5919,In_1715,In_2394);
nand U5920 (N_5920,In_2314,In_59);
nand U5921 (N_5921,In_842,In_2839);
nand U5922 (N_5922,In_2,In_525);
and U5923 (N_5923,In_1200,In_1989);
nand U5924 (N_5924,In_841,In_1635);
or U5925 (N_5925,In_1168,In_2502);
nand U5926 (N_5926,In_1889,In_194);
xor U5927 (N_5927,In_975,In_2960);
or U5928 (N_5928,In_717,In_61);
or U5929 (N_5929,In_2771,In_1840);
and U5930 (N_5930,In_2673,In_754);
nor U5931 (N_5931,In_2348,In_1453);
nand U5932 (N_5932,In_707,In_2777);
nor U5933 (N_5933,In_656,In_2537);
and U5934 (N_5934,In_751,In_2787);
xnor U5935 (N_5935,In_879,In_2165);
and U5936 (N_5936,In_2734,In_92);
nand U5937 (N_5937,In_2157,In_822);
and U5938 (N_5938,In_1353,In_2926);
or U5939 (N_5939,In_982,In_496);
nand U5940 (N_5940,In_276,In_2837);
and U5941 (N_5941,In_2689,In_1250);
nand U5942 (N_5942,In_1808,In_2068);
nor U5943 (N_5943,In_29,In_1348);
and U5944 (N_5944,In_1825,In_1579);
and U5945 (N_5945,In_1950,In_1099);
nand U5946 (N_5946,In_1204,In_408);
or U5947 (N_5947,In_2660,In_1065);
nor U5948 (N_5948,In_2185,In_1261);
and U5949 (N_5949,In_52,In_1485);
xor U5950 (N_5950,In_1961,In_1491);
nand U5951 (N_5951,In_947,In_2613);
and U5952 (N_5952,In_591,In_2164);
or U5953 (N_5953,In_210,In_1482);
nand U5954 (N_5954,In_1641,In_2805);
nor U5955 (N_5955,In_2463,In_2150);
nor U5956 (N_5956,In_2164,In_2894);
nor U5957 (N_5957,In_543,In_2918);
nand U5958 (N_5958,In_1816,In_709);
or U5959 (N_5959,In_1372,In_1157);
nor U5960 (N_5960,In_1092,In_1529);
nand U5961 (N_5961,In_1037,In_914);
xor U5962 (N_5962,In_2734,In_1180);
nor U5963 (N_5963,In_1938,In_219);
and U5964 (N_5964,In_881,In_946);
nor U5965 (N_5965,In_1008,In_2394);
xnor U5966 (N_5966,In_1852,In_2037);
nand U5967 (N_5967,In_1745,In_2959);
or U5968 (N_5968,In_542,In_1671);
xor U5969 (N_5969,In_2721,In_141);
and U5970 (N_5970,In_1901,In_1050);
xor U5971 (N_5971,In_1236,In_628);
or U5972 (N_5972,In_2795,In_1272);
nand U5973 (N_5973,In_2002,In_1798);
and U5974 (N_5974,In_65,In_172);
and U5975 (N_5975,In_2038,In_612);
nor U5976 (N_5976,In_2360,In_632);
and U5977 (N_5977,In_2566,In_311);
or U5978 (N_5978,In_1905,In_232);
and U5979 (N_5979,In_2489,In_1989);
xnor U5980 (N_5980,In_1896,In_838);
xnor U5981 (N_5981,In_868,In_1578);
nand U5982 (N_5982,In_2988,In_1254);
nand U5983 (N_5983,In_632,In_2364);
and U5984 (N_5984,In_2712,In_574);
xor U5985 (N_5985,In_297,In_2725);
and U5986 (N_5986,In_1927,In_77);
nand U5987 (N_5987,In_1641,In_36);
nor U5988 (N_5988,In_2075,In_236);
or U5989 (N_5989,In_2841,In_444);
nand U5990 (N_5990,In_948,In_2619);
and U5991 (N_5991,In_1797,In_2367);
nand U5992 (N_5992,In_1135,In_833);
nor U5993 (N_5993,In_1587,In_591);
nand U5994 (N_5994,In_205,In_1843);
nor U5995 (N_5995,In_951,In_721);
nor U5996 (N_5996,In_1736,In_2273);
and U5997 (N_5997,In_346,In_1437);
nor U5998 (N_5998,In_1311,In_1477);
nor U5999 (N_5999,In_1921,In_1421);
nand U6000 (N_6000,In_2159,In_2048);
and U6001 (N_6001,In_338,In_1510);
xnor U6002 (N_6002,In_339,In_200);
or U6003 (N_6003,In_315,In_2608);
nor U6004 (N_6004,In_222,In_979);
xor U6005 (N_6005,In_541,In_1050);
nor U6006 (N_6006,In_2304,In_65);
or U6007 (N_6007,In_798,In_231);
and U6008 (N_6008,In_1199,In_2314);
or U6009 (N_6009,In_615,In_1218);
xnor U6010 (N_6010,In_1365,In_2601);
and U6011 (N_6011,In_2193,In_2313);
or U6012 (N_6012,In_1486,In_2528);
and U6013 (N_6013,In_1288,In_527);
and U6014 (N_6014,In_2603,In_2768);
xor U6015 (N_6015,In_1120,In_2482);
or U6016 (N_6016,In_1054,In_1785);
nand U6017 (N_6017,In_1281,In_493);
xor U6018 (N_6018,In_156,In_1128);
nand U6019 (N_6019,In_156,In_806);
and U6020 (N_6020,In_2211,In_2750);
or U6021 (N_6021,In_776,In_772);
xor U6022 (N_6022,In_1283,In_326);
and U6023 (N_6023,In_767,In_2440);
or U6024 (N_6024,In_2021,In_632);
nand U6025 (N_6025,In_326,In_187);
and U6026 (N_6026,In_586,In_2277);
or U6027 (N_6027,In_437,In_835);
nand U6028 (N_6028,In_310,In_1409);
or U6029 (N_6029,In_2312,In_2857);
nor U6030 (N_6030,In_537,In_720);
nor U6031 (N_6031,In_899,In_502);
nand U6032 (N_6032,In_440,In_1859);
nand U6033 (N_6033,In_138,In_849);
xor U6034 (N_6034,In_619,In_1173);
or U6035 (N_6035,In_2560,In_715);
and U6036 (N_6036,In_1909,In_1258);
nand U6037 (N_6037,In_2587,In_914);
nand U6038 (N_6038,In_2916,In_1697);
or U6039 (N_6039,In_2484,In_1171);
and U6040 (N_6040,In_1167,In_2318);
nand U6041 (N_6041,In_2920,In_1891);
or U6042 (N_6042,In_2763,In_1163);
nand U6043 (N_6043,In_107,In_782);
or U6044 (N_6044,In_957,In_292);
and U6045 (N_6045,In_1062,In_2870);
nor U6046 (N_6046,In_553,In_460);
and U6047 (N_6047,In_1132,In_1853);
or U6048 (N_6048,In_1270,In_832);
xnor U6049 (N_6049,In_486,In_1162);
nor U6050 (N_6050,In_1432,In_838);
nand U6051 (N_6051,In_897,In_1293);
xor U6052 (N_6052,In_756,In_1772);
nand U6053 (N_6053,In_342,In_742);
nor U6054 (N_6054,In_2878,In_1776);
xnor U6055 (N_6055,In_1306,In_1785);
nor U6056 (N_6056,In_1073,In_2918);
and U6057 (N_6057,In_593,In_486);
nor U6058 (N_6058,In_2032,In_589);
xor U6059 (N_6059,In_2784,In_2675);
nor U6060 (N_6060,In_149,In_1496);
nand U6061 (N_6061,In_2885,In_1783);
or U6062 (N_6062,In_191,In_2481);
nand U6063 (N_6063,In_2319,In_2528);
or U6064 (N_6064,In_838,In_2283);
and U6065 (N_6065,In_389,In_1538);
xnor U6066 (N_6066,In_1442,In_208);
xor U6067 (N_6067,In_750,In_1488);
xnor U6068 (N_6068,In_2130,In_317);
nor U6069 (N_6069,In_68,In_186);
nor U6070 (N_6070,In_2607,In_1378);
xnor U6071 (N_6071,In_182,In_613);
nor U6072 (N_6072,In_2423,In_2137);
nand U6073 (N_6073,In_1841,In_110);
xor U6074 (N_6074,In_2443,In_2611);
or U6075 (N_6075,In_2745,In_2200);
nand U6076 (N_6076,In_1336,In_2497);
nand U6077 (N_6077,In_228,In_2787);
or U6078 (N_6078,In_2659,In_2795);
nand U6079 (N_6079,In_2471,In_651);
and U6080 (N_6080,In_982,In_1498);
or U6081 (N_6081,In_379,In_1442);
and U6082 (N_6082,In_926,In_1627);
and U6083 (N_6083,In_1920,In_2354);
nor U6084 (N_6084,In_873,In_2311);
xnor U6085 (N_6085,In_2114,In_57);
nand U6086 (N_6086,In_261,In_2528);
nor U6087 (N_6087,In_1128,In_166);
or U6088 (N_6088,In_2755,In_257);
and U6089 (N_6089,In_408,In_1129);
or U6090 (N_6090,In_1341,In_410);
or U6091 (N_6091,In_2818,In_890);
nand U6092 (N_6092,In_2197,In_2834);
nor U6093 (N_6093,In_2486,In_457);
and U6094 (N_6094,In_1950,In_1535);
nor U6095 (N_6095,In_2596,In_959);
nor U6096 (N_6096,In_1779,In_2631);
xnor U6097 (N_6097,In_2498,In_892);
or U6098 (N_6098,In_2360,In_955);
and U6099 (N_6099,In_2499,In_312);
and U6100 (N_6100,In_1827,In_1794);
and U6101 (N_6101,In_1520,In_1436);
nor U6102 (N_6102,In_1610,In_2674);
or U6103 (N_6103,In_1799,In_2211);
or U6104 (N_6104,In_2063,In_1769);
and U6105 (N_6105,In_992,In_1849);
xor U6106 (N_6106,In_1175,In_2856);
and U6107 (N_6107,In_1574,In_350);
or U6108 (N_6108,In_695,In_113);
nor U6109 (N_6109,In_2007,In_2849);
xnor U6110 (N_6110,In_471,In_1828);
xor U6111 (N_6111,In_2965,In_2584);
nand U6112 (N_6112,In_1971,In_1345);
xor U6113 (N_6113,In_2822,In_2802);
nand U6114 (N_6114,In_1407,In_1272);
xor U6115 (N_6115,In_794,In_174);
nor U6116 (N_6116,In_1594,In_1127);
nor U6117 (N_6117,In_1616,In_2823);
nor U6118 (N_6118,In_1272,In_276);
and U6119 (N_6119,In_2332,In_728);
nand U6120 (N_6120,In_1870,In_1714);
or U6121 (N_6121,In_2174,In_1513);
and U6122 (N_6122,In_77,In_336);
and U6123 (N_6123,In_1282,In_1874);
xor U6124 (N_6124,In_2791,In_2240);
xnor U6125 (N_6125,In_1203,In_1095);
nand U6126 (N_6126,In_2787,In_1513);
and U6127 (N_6127,In_115,In_38);
xor U6128 (N_6128,In_2324,In_2548);
nand U6129 (N_6129,In_593,In_1969);
xnor U6130 (N_6130,In_1276,In_1146);
xor U6131 (N_6131,In_1458,In_570);
and U6132 (N_6132,In_99,In_1203);
or U6133 (N_6133,In_1136,In_1400);
nor U6134 (N_6134,In_1911,In_1221);
nand U6135 (N_6135,In_1845,In_859);
nand U6136 (N_6136,In_2047,In_484);
xnor U6137 (N_6137,In_2973,In_1151);
nor U6138 (N_6138,In_429,In_1292);
or U6139 (N_6139,In_32,In_1397);
and U6140 (N_6140,In_2593,In_2558);
or U6141 (N_6141,In_2687,In_2761);
or U6142 (N_6142,In_230,In_1796);
or U6143 (N_6143,In_838,In_458);
xnor U6144 (N_6144,In_2118,In_691);
nand U6145 (N_6145,In_2680,In_1681);
and U6146 (N_6146,In_1195,In_2361);
and U6147 (N_6147,In_205,In_223);
or U6148 (N_6148,In_1100,In_318);
nand U6149 (N_6149,In_125,In_2243);
nor U6150 (N_6150,In_736,In_141);
or U6151 (N_6151,In_1765,In_2419);
or U6152 (N_6152,In_570,In_2047);
or U6153 (N_6153,In_794,In_1377);
nand U6154 (N_6154,In_1881,In_238);
nand U6155 (N_6155,In_1255,In_2501);
xor U6156 (N_6156,In_1504,In_2264);
nand U6157 (N_6157,In_2487,In_925);
nand U6158 (N_6158,In_1502,In_2322);
xor U6159 (N_6159,In_2979,In_1430);
xor U6160 (N_6160,In_2419,In_934);
xor U6161 (N_6161,In_2456,In_542);
xnor U6162 (N_6162,In_190,In_2638);
nand U6163 (N_6163,In_2619,In_304);
xor U6164 (N_6164,In_1748,In_1457);
and U6165 (N_6165,In_1275,In_1296);
or U6166 (N_6166,In_1054,In_1862);
or U6167 (N_6167,In_2106,In_2634);
or U6168 (N_6168,In_878,In_2237);
xor U6169 (N_6169,In_1804,In_2860);
and U6170 (N_6170,In_1734,In_1065);
nand U6171 (N_6171,In_405,In_271);
nand U6172 (N_6172,In_147,In_2345);
nor U6173 (N_6173,In_1891,In_1109);
or U6174 (N_6174,In_2180,In_2381);
and U6175 (N_6175,In_939,In_459);
xor U6176 (N_6176,In_581,In_1082);
or U6177 (N_6177,In_562,In_2062);
nand U6178 (N_6178,In_1050,In_563);
nand U6179 (N_6179,In_489,In_2658);
and U6180 (N_6180,In_379,In_2385);
nor U6181 (N_6181,In_890,In_859);
and U6182 (N_6182,In_1629,In_2154);
xor U6183 (N_6183,In_62,In_2754);
or U6184 (N_6184,In_1539,In_1738);
nor U6185 (N_6185,In_1972,In_2532);
nand U6186 (N_6186,In_2330,In_2317);
xor U6187 (N_6187,In_142,In_2148);
or U6188 (N_6188,In_527,In_1092);
xor U6189 (N_6189,In_1009,In_2211);
nor U6190 (N_6190,In_2419,In_508);
or U6191 (N_6191,In_946,In_2210);
xor U6192 (N_6192,In_230,In_685);
nor U6193 (N_6193,In_887,In_2993);
nor U6194 (N_6194,In_412,In_522);
nor U6195 (N_6195,In_1548,In_1203);
nor U6196 (N_6196,In_96,In_1022);
nand U6197 (N_6197,In_2927,In_68);
nor U6198 (N_6198,In_447,In_2360);
and U6199 (N_6199,In_919,In_184);
and U6200 (N_6200,In_1108,In_987);
nand U6201 (N_6201,In_1995,In_2018);
xor U6202 (N_6202,In_173,In_1178);
xor U6203 (N_6203,In_1291,In_2526);
or U6204 (N_6204,In_964,In_2292);
nor U6205 (N_6205,In_2174,In_2954);
xnor U6206 (N_6206,In_2566,In_2532);
or U6207 (N_6207,In_2618,In_2357);
nand U6208 (N_6208,In_187,In_485);
nand U6209 (N_6209,In_2663,In_2377);
nor U6210 (N_6210,In_1244,In_2562);
xor U6211 (N_6211,In_2303,In_2432);
xnor U6212 (N_6212,In_1703,In_175);
nor U6213 (N_6213,In_2567,In_1021);
xor U6214 (N_6214,In_1508,In_979);
nand U6215 (N_6215,In_2210,In_2259);
xnor U6216 (N_6216,In_951,In_2161);
nor U6217 (N_6217,In_662,In_2953);
nor U6218 (N_6218,In_52,In_1720);
nor U6219 (N_6219,In_1217,In_1621);
xor U6220 (N_6220,In_346,In_1024);
nor U6221 (N_6221,In_821,In_1311);
nand U6222 (N_6222,In_2807,In_1417);
and U6223 (N_6223,In_2117,In_2550);
nor U6224 (N_6224,In_1501,In_1641);
or U6225 (N_6225,In_2283,In_1108);
nor U6226 (N_6226,In_1116,In_2552);
and U6227 (N_6227,In_2403,In_1403);
and U6228 (N_6228,In_2397,In_1374);
nor U6229 (N_6229,In_19,In_1969);
nand U6230 (N_6230,In_2184,In_1506);
xnor U6231 (N_6231,In_2643,In_350);
nand U6232 (N_6232,In_1621,In_2152);
nor U6233 (N_6233,In_472,In_2978);
or U6234 (N_6234,In_1722,In_1036);
nor U6235 (N_6235,In_1481,In_142);
xor U6236 (N_6236,In_2062,In_649);
nor U6237 (N_6237,In_1642,In_929);
or U6238 (N_6238,In_115,In_2375);
nor U6239 (N_6239,In_1156,In_1129);
nand U6240 (N_6240,In_845,In_2232);
and U6241 (N_6241,In_1782,In_2546);
and U6242 (N_6242,In_870,In_2755);
nand U6243 (N_6243,In_1429,In_818);
nor U6244 (N_6244,In_72,In_1141);
and U6245 (N_6245,In_2676,In_543);
and U6246 (N_6246,In_487,In_1742);
nor U6247 (N_6247,In_2456,In_1039);
nor U6248 (N_6248,In_295,In_2303);
nand U6249 (N_6249,In_736,In_1135);
xnor U6250 (N_6250,In_1681,In_2108);
xnor U6251 (N_6251,In_382,In_2164);
nand U6252 (N_6252,In_633,In_1004);
nand U6253 (N_6253,In_2000,In_1733);
nor U6254 (N_6254,In_2849,In_1893);
nor U6255 (N_6255,In_2080,In_981);
or U6256 (N_6256,In_421,In_1551);
and U6257 (N_6257,In_484,In_2032);
nand U6258 (N_6258,In_46,In_2069);
nor U6259 (N_6259,In_1544,In_365);
xor U6260 (N_6260,In_2082,In_2287);
and U6261 (N_6261,In_2574,In_2800);
nand U6262 (N_6262,In_55,In_237);
or U6263 (N_6263,In_611,In_2454);
or U6264 (N_6264,In_2386,In_713);
nor U6265 (N_6265,In_1348,In_613);
nor U6266 (N_6266,In_758,In_1938);
or U6267 (N_6267,In_773,In_1276);
nor U6268 (N_6268,In_2025,In_1682);
or U6269 (N_6269,In_2833,In_2985);
nor U6270 (N_6270,In_810,In_2379);
and U6271 (N_6271,In_23,In_408);
nand U6272 (N_6272,In_2314,In_2066);
and U6273 (N_6273,In_793,In_1992);
xor U6274 (N_6274,In_2671,In_322);
nand U6275 (N_6275,In_1890,In_2963);
nand U6276 (N_6276,In_196,In_1685);
xnor U6277 (N_6277,In_2508,In_923);
xor U6278 (N_6278,In_1892,In_1478);
nor U6279 (N_6279,In_2227,In_2018);
nand U6280 (N_6280,In_1016,In_2496);
nor U6281 (N_6281,In_1105,In_684);
and U6282 (N_6282,In_1475,In_359);
xnor U6283 (N_6283,In_15,In_2817);
xnor U6284 (N_6284,In_688,In_69);
xnor U6285 (N_6285,In_2119,In_684);
and U6286 (N_6286,In_1985,In_2484);
xor U6287 (N_6287,In_454,In_2578);
and U6288 (N_6288,In_846,In_136);
and U6289 (N_6289,In_1282,In_1076);
or U6290 (N_6290,In_1964,In_103);
xnor U6291 (N_6291,In_383,In_2353);
xnor U6292 (N_6292,In_1203,In_953);
or U6293 (N_6293,In_1239,In_2974);
nor U6294 (N_6294,In_2816,In_1150);
nand U6295 (N_6295,In_193,In_630);
nor U6296 (N_6296,In_1028,In_1589);
nor U6297 (N_6297,In_1981,In_746);
xor U6298 (N_6298,In_360,In_942);
or U6299 (N_6299,In_1477,In_449);
or U6300 (N_6300,In_98,In_50);
xor U6301 (N_6301,In_46,In_2426);
xor U6302 (N_6302,In_872,In_2525);
and U6303 (N_6303,In_937,In_828);
and U6304 (N_6304,In_1840,In_2574);
or U6305 (N_6305,In_2152,In_479);
and U6306 (N_6306,In_2652,In_1859);
or U6307 (N_6307,In_1057,In_1609);
xnor U6308 (N_6308,In_926,In_1423);
or U6309 (N_6309,In_1889,In_1673);
nand U6310 (N_6310,In_1067,In_2384);
nand U6311 (N_6311,In_575,In_983);
nand U6312 (N_6312,In_502,In_1621);
nor U6313 (N_6313,In_2832,In_865);
or U6314 (N_6314,In_423,In_1624);
or U6315 (N_6315,In_2743,In_1004);
xor U6316 (N_6316,In_2800,In_1941);
and U6317 (N_6317,In_246,In_1091);
nand U6318 (N_6318,In_1040,In_2790);
xnor U6319 (N_6319,In_1909,In_1151);
or U6320 (N_6320,In_1291,In_2828);
nor U6321 (N_6321,In_801,In_2798);
nor U6322 (N_6322,In_2456,In_521);
nand U6323 (N_6323,In_1730,In_2651);
nand U6324 (N_6324,In_1644,In_2905);
or U6325 (N_6325,In_1347,In_1556);
or U6326 (N_6326,In_1269,In_313);
or U6327 (N_6327,In_1964,In_952);
xnor U6328 (N_6328,In_1112,In_568);
or U6329 (N_6329,In_2645,In_1844);
xor U6330 (N_6330,In_2847,In_115);
xor U6331 (N_6331,In_86,In_2903);
nor U6332 (N_6332,In_2935,In_428);
xnor U6333 (N_6333,In_2179,In_17);
nor U6334 (N_6334,In_1806,In_2938);
or U6335 (N_6335,In_1278,In_1665);
and U6336 (N_6336,In_2595,In_581);
xnor U6337 (N_6337,In_276,In_69);
and U6338 (N_6338,In_1403,In_1180);
nand U6339 (N_6339,In_2814,In_752);
nand U6340 (N_6340,In_978,In_2993);
and U6341 (N_6341,In_2397,In_1278);
or U6342 (N_6342,In_2123,In_837);
xor U6343 (N_6343,In_1697,In_1235);
nor U6344 (N_6344,In_1168,In_1688);
or U6345 (N_6345,In_2513,In_2082);
or U6346 (N_6346,In_231,In_244);
and U6347 (N_6347,In_2332,In_856);
xor U6348 (N_6348,In_1473,In_691);
nor U6349 (N_6349,In_2679,In_1534);
nand U6350 (N_6350,In_1271,In_2730);
or U6351 (N_6351,In_429,In_1187);
or U6352 (N_6352,In_1210,In_2956);
xnor U6353 (N_6353,In_2790,In_2110);
xor U6354 (N_6354,In_2814,In_1028);
xor U6355 (N_6355,In_2478,In_487);
or U6356 (N_6356,In_97,In_112);
and U6357 (N_6357,In_2092,In_1326);
xor U6358 (N_6358,In_380,In_2213);
xnor U6359 (N_6359,In_4,In_887);
or U6360 (N_6360,In_398,In_445);
or U6361 (N_6361,In_2692,In_297);
nand U6362 (N_6362,In_1351,In_1758);
and U6363 (N_6363,In_758,In_110);
or U6364 (N_6364,In_2874,In_330);
and U6365 (N_6365,In_1845,In_131);
xnor U6366 (N_6366,In_429,In_720);
or U6367 (N_6367,In_282,In_2209);
nor U6368 (N_6368,In_371,In_265);
or U6369 (N_6369,In_2420,In_82);
or U6370 (N_6370,In_2736,In_2281);
xnor U6371 (N_6371,In_764,In_1745);
nor U6372 (N_6372,In_469,In_1366);
xor U6373 (N_6373,In_2712,In_2856);
nor U6374 (N_6374,In_1494,In_1900);
nor U6375 (N_6375,In_2544,In_931);
nand U6376 (N_6376,In_2675,In_2627);
nand U6377 (N_6377,In_380,In_2522);
nand U6378 (N_6378,In_531,In_1251);
nand U6379 (N_6379,In_1138,In_1751);
or U6380 (N_6380,In_2502,In_1437);
nor U6381 (N_6381,In_1614,In_2986);
nand U6382 (N_6382,In_1651,In_1575);
xnor U6383 (N_6383,In_2365,In_1815);
nand U6384 (N_6384,In_2571,In_2410);
or U6385 (N_6385,In_1725,In_714);
nor U6386 (N_6386,In_111,In_1941);
or U6387 (N_6387,In_2787,In_1989);
or U6388 (N_6388,In_913,In_1811);
or U6389 (N_6389,In_2774,In_2175);
xnor U6390 (N_6390,In_202,In_2980);
nand U6391 (N_6391,In_869,In_2156);
or U6392 (N_6392,In_1953,In_1627);
or U6393 (N_6393,In_2835,In_1847);
or U6394 (N_6394,In_2232,In_951);
or U6395 (N_6395,In_1151,In_2173);
and U6396 (N_6396,In_2881,In_453);
xor U6397 (N_6397,In_457,In_1836);
nand U6398 (N_6398,In_1749,In_2530);
and U6399 (N_6399,In_2663,In_2396);
nor U6400 (N_6400,In_2469,In_1043);
nand U6401 (N_6401,In_1217,In_2158);
or U6402 (N_6402,In_2662,In_916);
xnor U6403 (N_6403,In_902,In_795);
nand U6404 (N_6404,In_979,In_2163);
xor U6405 (N_6405,In_1562,In_2369);
or U6406 (N_6406,In_1956,In_1743);
or U6407 (N_6407,In_1616,In_1888);
or U6408 (N_6408,In_847,In_877);
and U6409 (N_6409,In_2783,In_431);
nand U6410 (N_6410,In_475,In_1743);
xor U6411 (N_6411,In_67,In_2021);
and U6412 (N_6412,In_2820,In_2038);
and U6413 (N_6413,In_128,In_177);
nand U6414 (N_6414,In_2794,In_965);
and U6415 (N_6415,In_1587,In_1639);
or U6416 (N_6416,In_2403,In_2887);
and U6417 (N_6417,In_1059,In_1198);
nor U6418 (N_6418,In_439,In_1006);
and U6419 (N_6419,In_2362,In_1664);
and U6420 (N_6420,In_2763,In_1909);
nor U6421 (N_6421,In_203,In_2150);
or U6422 (N_6422,In_282,In_663);
and U6423 (N_6423,In_142,In_1256);
nor U6424 (N_6424,In_854,In_2413);
or U6425 (N_6425,In_1730,In_2392);
nor U6426 (N_6426,In_47,In_809);
nor U6427 (N_6427,In_1782,In_817);
or U6428 (N_6428,In_813,In_154);
or U6429 (N_6429,In_360,In_1195);
or U6430 (N_6430,In_2550,In_829);
or U6431 (N_6431,In_2845,In_1192);
and U6432 (N_6432,In_299,In_2923);
or U6433 (N_6433,In_2921,In_1282);
nand U6434 (N_6434,In_2816,In_2191);
nor U6435 (N_6435,In_84,In_2854);
xnor U6436 (N_6436,In_1603,In_2326);
nor U6437 (N_6437,In_73,In_2214);
xor U6438 (N_6438,In_2115,In_1573);
nor U6439 (N_6439,In_2170,In_2283);
and U6440 (N_6440,In_505,In_921);
xor U6441 (N_6441,In_110,In_602);
and U6442 (N_6442,In_1152,In_641);
nand U6443 (N_6443,In_2974,In_1294);
nor U6444 (N_6444,In_1445,In_1500);
nor U6445 (N_6445,In_2056,In_2153);
nor U6446 (N_6446,In_868,In_2767);
and U6447 (N_6447,In_2401,In_1915);
xor U6448 (N_6448,In_2098,In_415);
or U6449 (N_6449,In_1797,In_322);
nand U6450 (N_6450,In_2411,In_2845);
xor U6451 (N_6451,In_2080,In_1922);
and U6452 (N_6452,In_2780,In_1220);
xor U6453 (N_6453,In_2329,In_771);
nand U6454 (N_6454,In_1364,In_1258);
and U6455 (N_6455,In_144,In_1086);
and U6456 (N_6456,In_647,In_138);
nor U6457 (N_6457,In_1958,In_2244);
nand U6458 (N_6458,In_737,In_723);
and U6459 (N_6459,In_827,In_2531);
and U6460 (N_6460,In_1012,In_1205);
nor U6461 (N_6461,In_938,In_1927);
nor U6462 (N_6462,In_2243,In_988);
or U6463 (N_6463,In_2175,In_570);
nand U6464 (N_6464,In_2835,In_621);
nand U6465 (N_6465,In_2435,In_368);
xor U6466 (N_6466,In_81,In_1820);
xor U6467 (N_6467,In_1307,In_1027);
xor U6468 (N_6468,In_209,In_627);
and U6469 (N_6469,In_2538,In_2025);
nand U6470 (N_6470,In_2366,In_2884);
nor U6471 (N_6471,In_2120,In_2520);
nand U6472 (N_6472,In_1769,In_1596);
nand U6473 (N_6473,In_416,In_2665);
nand U6474 (N_6474,In_470,In_1312);
or U6475 (N_6475,In_1398,In_2096);
nand U6476 (N_6476,In_1266,In_1820);
xor U6477 (N_6477,In_941,In_439);
and U6478 (N_6478,In_995,In_2055);
and U6479 (N_6479,In_1467,In_1179);
and U6480 (N_6480,In_1193,In_2201);
nand U6481 (N_6481,In_2949,In_1547);
and U6482 (N_6482,In_2643,In_160);
or U6483 (N_6483,In_1346,In_1979);
nand U6484 (N_6484,In_1431,In_242);
nand U6485 (N_6485,In_2069,In_2495);
and U6486 (N_6486,In_2280,In_1780);
nor U6487 (N_6487,In_1421,In_2360);
xnor U6488 (N_6488,In_2267,In_2550);
nand U6489 (N_6489,In_2256,In_1777);
xnor U6490 (N_6490,In_1512,In_2631);
nor U6491 (N_6491,In_1951,In_2173);
xnor U6492 (N_6492,In_2969,In_702);
xor U6493 (N_6493,In_1110,In_461);
nand U6494 (N_6494,In_736,In_1595);
nand U6495 (N_6495,In_2042,In_1100);
and U6496 (N_6496,In_1794,In_60);
nand U6497 (N_6497,In_2785,In_496);
and U6498 (N_6498,In_1705,In_1598);
xnor U6499 (N_6499,In_617,In_1129);
xnor U6500 (N_6500,In_1831,In_193);
and U6501 (N_6501,In_2466,In_472);
or U6502 (N_6502,In_127,In_2090);
and U6503 (N_6503,In_2661,In_1947);
xor U6504 (N_6504,In_2739,In_1153);
nand U6505 (N_6505,In_2379,In_1133);
xor U6506 (N_6506,In_1472,In_2460);
and U6507 (N_6507,In_1755,In_2643);
nand U6508 (N_6508,In_1855,In_2245);
nor U6509 (N_6509,In_1619,In_2574);
xor U6510 (N_6510,In_2764,In_398);
xor U6511 (N_6511,In_295,In_1224);
or U6512 (N_6512,In_2897,In_1450);
nand U6513 (N_6513,In_2120,In_37);
and U6514 (N_6514,In_535,In_2351);
and U6515 (N_6515,In_411,In_1388);
and U6516 (N_6516,In_1603,In_2428);
or U6517 (N_6517,In_2006,In_2718);
nor U6518 (N_6518,In_1141,In_1521);
nand U6519 (N_6519,In_1063,In_1952);
xnor U6520 (N_6520,In_167,In_2637);
nor U6521 (N_6521,In_1546,In_1431);
nand U6522 (N_6522,In_1290,In_272);
xnor U6523 (N_6523,In_108,In_1390);
nand U6524 (N_6524,In_1820,In_1476);
nand U6525 (N_6525,In_1287,In_153);
xor U6526 (N_6526,In_2541,In_267);
and U6527 (N_6527,In_514,In_2256);
xnor U6528 (N_6528,In_1525,In_1608);
nor U6529 (N_6529,In_2223,In_418);
nand U6530 (N_6530,In_459,In_748);
nor U6531 (N_6531,In_1647,In_1334);
nand U6532 (N_6532,In_2330,In_1687);
nor U6533 (N_6533,In_63,In_1835);
or U6534 (N_6534,In_1748,In_228);
and U6535 (N_6535,In_266,In_658);
and U6536 (N_6536,In_2369,In_2894);
nand U6537 (N_6537,In_1994,In_634);
nand U6538 (N_6538,In_1208,In_1851);
xnor U6539 (N_6539,In_2704,In_2232);
nand U6540 (N_6540,In_2303,In_1461);
nand U6541 (N_6541,In_1322,In_978);
or U6542 (N_6542,In_1414,In_1207);
and U6543 (N_6543,In_733,In_1844);
or U6544 (N_6544,In_2565,In_2831);
and U6545 (N_6545,In_1171,In_607);
or U6546 (N_6546,In_2677,In_169);
xnor U6547 (N_6547,In_1492,In_2994);
nor U6548 (N_6548,In_2161,In_652);
and U6549 (N_6549,In_1513,In_1956);
nor U6550 (N_6550,In_1810,In_1282);
and U6551 (N_6551,In_1954,In_160);
xor U6552 (N_6552,In_51,In_668);
or U6553 (N_6553,In_550,In_1464);
and U6554 (N_6554,In_2595,In_1190);
and U6555 (N_6555,In_2586,In_2608);
xnor U6556 (N_6556,In_62,In_1336);
nor U6557 (N_6557,In_1124,In_1363);
xnor U6558 (N_6558,In_662,In_2994);
xnor U6559 (N_6559,In_381,In_186);
nand U6560 (N_6560,In_2540,In_653);
or U6561 (N_6561,In_1041,In_1601);
and U6562 (N_6562,In_304,In_1177);
nand U6563 (N_6563,In_1737,In_1100);
or U6564 (N_6564,In_1509,In_2052);
nand U6565 (N_6565,In_1820,In_1100);
and U6566 (N_6566,In_2146,In_1574);
or U6567 (N_6567,In_2595,In_4);
nand U6568 (N_6568,In_1118,In_1368);
or U6569 (N_6569,In_2922,In_1400);
nand U6570 (N_6570,In_2464,In_1094);
nand U6571 (N_6571,In_989,In_984);
nand U6572 (N_6572,In_1421,In_2955);
or U6573 (N_6573,In_568,In_657);
xor U6574 (N_6574,In_2441,In_1237);
xor U6575 (N_6575,In_514,In_143);
or U6576 (N_6576,In_956,In_2558);
nor U6577 (N_6577,In_999,In_2192);
or U6578 (N_6578,In_369,In_460);
nor U6579 (N_6579,In_278,In_2721);
nand U6580 (N_6580,In_2897,In_2855);
nand U6581 (N_6581,In_1141,In_1621);
nor U6582 (N_6582,In_849,In_2637);
xnor U6583 (N_6583,In_1325,In_2448);
nor U6584 (N_6584,In_1319,In_1190);
nand U6585 (N_6585,In_2898,In_1877);
and U6586 (N_6586,In_636,In_1528);
or U6587 (N_6587,In_2865,In_1137);
nor U6588 (N_6588,In_2106,In_956);
nand U6589 (N_6589,In_2579,In_2868);
nor U6590 (N_6590,In_2066,In_2085);
nand U6591 (N_6591,In_2198,In_564);
nor U6592 (N_6592,In_1912,In_1541);
or U6593 (N_6593,In_2888,In_1851);
nand U6594 (N_6594,In_663,In_2916);
and U6595 (N_6595,In_1248,In_423);
or U6596 (N_6596,In_901,In_1963);
nand U6597 (N_6597,In_126,In_97);
nor U6598 (N_6598,In_2271,In_2413);
nand U6599 (N_6599,In_90,In_1144);
or U6600 (N_6600,In_2629,In_2415);
nor U6601 (N_6601,In_133,In_2950);
xnor U6602 (N_6602,In_1872,In_1185);
or U6603 (N_6603,In_2444,In_2579);
and U6604 (N_6604,In_879,In_2538);
or U6605 (N_6605,In_195,In_1117);
or U6606 (N_6606,In_1908,In_483);
nand U6607 (N_6607,In_1500,In_1654);
xnor U6608 (N_6608,In_1435,In_1770);
or U6609 (N_6609,In_836,In_1150);
nand U6610 (N_6610,In_705,In_699);
or U6611 (N_6611,In_2287,In_2400);
nor U6612 (N_6612,In_495,In_2475);
and U6613 (N_6613,In_591,In_711);
or U6614 (N_6614,In_2947,In_1712);
nand U6615 (N_6615,In_1684,In_1465);
or U6616 (N_6616,In_131,In_830);
xor U6617 (N_6617,In_2042,In_1150);
and U6618 (N_6618,In_2417,In_2206);
nor U6619 (N_6619,In_2959,In_2467);
nor U6620 (N_6620,In_313,In_735);
or U6621 (N_6621,In_1752,In_1903);
nand U6622 (N_6622,In_259,In_2736);
nand U6623 (N_6623,In_899,In_178);
nand U6624 (N_6624,In_2379,In_2162);
xnor U6625 (N_6625,In_535,In_2840);
nor U6626 (N_6626,In_2355,In_1904);
xor U6627 (N_6627,In_396,In_729);
nor U6628 (N_6628,In_870,In_2253);
nand U6629 (N_6629,In_2112,In_361);
nor U6630 (N_6630,In_135,In_200);
nand U6631 (N_6631,In_818,In_2342);
and U6632 (N_6632,In_2194,In_200);
nor U6633 (N_6633,In_2432,In_2453);
or U6634 (N_6634,In_444,In_708);
and U6635 (N_6635,In_1873,In_781);
xnor U6636 (N_6636,In_62,In_546);
nor U6637 (N_6637,In_2875,In_246);
or U6638 (N_6638,In_2587,In_1243);
or U6639 (N_6639,In_318,In_1712);
nor U6640 (N_6640,In_2109,In_2048);
or U6641 (N_6641,In_596,In_1433);
or U6642 (N_6642,In_1618,In_947);
nor U6643 (N_6643,In_70,In_590);
nor U6644 (N_6644,In_2322,In_2045);
nor U6645 (N_6645,In_1886,In_2738);
and U6646 (N_6646,In_680,In_1065);
nand U6647 (N_6647,In_151,In_2181);
or U6648 (N_6648,In_1434,In_2921);
and U6649 (N_6649,In_2282,In_2012);
or U6650 (N_6650,In_475,In_2130);
nor U6651 (N_6651,In_1938,In_2968);
or U6652 (N_6652,In_1208,In_2627);
xor U6653 (N_6653,In_537,In_376);
nand U6654 (N_6654,In_1706,In_2363);
or U6655 (N_6655,In_188,In_1701);
and U6656 (N_6656,In_1850,In_1659);
or U6657 (N_6657,In_813,In_1132);
nand U6658 (N_6658,In_1007,In_1165);
or U6659 (N_6659,In_1286,In_2700);
nor U6660 (N_6660,In_1537,In_2135);
and U6661 (N_6661,In_864,In_1084);
and U6662 (N_6662,In_1706,In_447);
nor U6663 (N_6663,In_1615,In_2910);
nand U6664 (N_6664,In_2140,In_1137);
xnor U6665 (N_6665,In_876,In_164);
nor U6666 (N_6666,In_809,In_1222);
and U6667 (N_6667,In_1335,In_1421);
and U6668 (N_6668,In_298,In_1422);
nor U6669 (N_6669,In_309,In_1219);
nor U6670 (N_6670,In_2643,In_16);
xnor U6671 (N_6671,In_1210,In_2702);
nor U6672 (N_6672,In_685,In_2076);
nand U6673 (N_6673,In_1989,In_987);
and U6674 (N_6674,In_861,In_2107);
and U6675 (N_6675,In_380,In_1601);
and U6676 (N_6676,In_2603,In_1518);
nor U6677 (N_6677,In_2524,In_619);
or U6678 (N_6678,In_319,In_2144);
or U6679 (N_6679,In_1525,In_757);
nor U6680 (N_6680,In_2209,In_1893);
or U6681 (N_6681,In_2262,In_864);
or U6682 (N_6682,In_1391,In_134);
or U6683 (N_6683,In_365,In_1247);
xnor U6684 (N_6684,In_1589,In_2374);
or U6685 (N_6685,In_1112,In_640);
and U6686 (N_6686,In_354,In_376);
or U6687 (N_6687,In_2266,In_2509);
nand U6688 (N_6688,In_2981,In_2924);
nor U6689 (N_6689,In_2223,In_2690);
or U6690 (N_6690,In_331,In_862);
xnor U6691 (N_6691,In_34,In_706);
or U6692 (N_6692,In_2740,In_965);
and U6693 (N_6693,In_245,In_1369);
nor U6694 (N_6694,In_571,In_2904);
nor U6695 (N_6695,In_2116,In_2526);
or U6696 (N_6696,In_346,In_2398);
nand U6697 (N_6697,In_2605,In_438);
or U6698 (N_6698,In_2770,In_2333);
or U6699 (N_6699,In_2416,In_2880);
nor U6700 (N_6700,In_2798,In_1893);
xor U6701 (N_6701,In_2678,In_2089);
nor U6702 (N_6702,In_1117,In_1248);
or U6703 (N_6703,In_2368,In_2503);
xnor U6704 (N_6704,In_2981,In_504);
and U6705 (N_6705,In_398,In_181);
nor U6706 (N_6706,In_2380,In_893);
or U6707 (N_6707,In_486,In_49);
nand U6708 (N_6708,In_1790,In_2418);
and U6709 (N_6709,In_2994,In_244);
and U6710 (N_6710,In_2733,In_74);
or U6711 (N_6711,In_243,In_525);
xnor U6712 (N_6712,In_1317,In_994);
and U6713 (N_6713,In_1310,In_473);
nor U6714 (N_6714,In_2582,In_1787);
xor U6715 (N_6715,In_1897,In_1918);
or U6716 (N_6716,In_898,In_2402);
nor U6717 (N_6717,In_2790,In_2581);
xor U6718 (N_6718,In_1825,In_2521);
nand U6719 (N_6719,In_219,In_1522);
xor U6720 (N_6720,In_2422,In_2489);
nand U6721 (N_6721,In_429,In_2860);
or U6722 (N_6722,In_883,In_347);
nor U6723 (N_6723,In_1241,In_425);
xor U6724 (N_6724,In_441,In_2957);
nor U6725 (N_6725,In_197,In_1737);
and U6726 (N_6726,In_2729,In_947);
nand U6727 (N_6727,In_1704,In_212);
or U6728 (N_6728,In_22,In_2330);
and U6729 (N_6729,In_257,In_1091);
nand U6730 (N_6730,In_636,In_925);
nor U6731 (N_6731,In_682,In_2016);
and U6732 (N_6732,In_865,In_822);
nand U6733 (N_6733,In_163,In_2408);
nor U6734 (N_6734,In_1700,In_556);
or U6735 (N_6735,In_1617,In_2624);
nand U6736 (N_6736,In_2431,In_2493);
nor U6737 (N_6737,In_1267,In_2324);
nand U6738 (N_6738,In_60,In_2267);
or U6739 (N_6739,In_824,In_536);
nor U6740 (N_6740,In_1243,In_539);
nor U6741 (N_6741,In_317,In_2817);
nor U6742 (N_6742,In_2794,In_530);
and U6743 (N_6743,In_488,In_845);
or U6744 (N_6744,In_657,In_725);
nor U6745 (N_6745,In_2252,In_2487);
nand U6746 (N_6746,In_2973,In_1295);
nand U6747 (N_6747,In_2651,In_2541);
nand U6748 (N_6748,In_402,In_634);
nand U6749 (N_6749,In_482,In_750);
nor U6750 (N_6750,In_1737,In_847);
and U6751 (N_6751,In_1040,In_2557);
nand U6752 (N_6752,In_545,In_441);
xnor U6753 (N_6753,In_2308,In_2114);
nand U6754 (N_6754,In_2829,In_242);
and U6755 (N_6755,In_2205,In_155);
nand U6756 (N_6756,In_2139,In_1655);
or U6757 (N_6757,In_2379,In_2429);
and U6758 (N_6758,In_2250,In_719);
xnor U6759 (N_6759,In_2196,In_1498);
nor U6760 (N_6760,In_805,In_15);
nor U6761 (N_6761,In_1200,In_2718);
and U6762 (N_6762,In_1732,In_1780);
nor U6763 (N_6763,In_714,In_1487);
nand U6764 (N_6764,In_923,In_218);
nor U6765 (N_6765,In_2230,In_1749);
or U6766 (N_6766,In_1277,In_2370);
xor U6767 (N_6767,In_1482,In_1087);
nor U6768 (N_6768,In_338,In_388);
and U6769 (N_6769,In_69,In_2319);
nand U6770 (N_6770,In_1119,In_1458);
nand U6771 (N_6771,In_1144,In_2941);
xnor U6772 (N_6772,In_2074,In_681);
xor U6773 (N_6773,In_1589,In_2458);
and U6774 (N_6774,In_2488,In_1222);
or U6775 (N_6775,In_2920,In_444);
or U6776 (N_6776,In_1614,In_2967);
xnor U6777 (N_6777,In_975,In_671);
or U6778 (N_6778,In_1452,In_1606);
nor U6779 (N_6779,In_2941,In_37);
xor U6780 (N_6780,In_1126,In_2477);
nor U6781 (N_6781,In_1925,In_1361);
nand U6782 (N_6782,In_178,In_415);
and U6783 (N_6783,In_1956,In_2469);
and U6784 (N_6784,In_1213,In_1291);
and U6785 (N_6785,In_2246,In_1180);
nand U6786 (N_6786,In_2096,In_294);
xor U6787 (N_6787,In_1488,In_682);
or U6788 (N_6788,In_630,In_254);
and U6789 (N_6789,In_1518,In_2081);
nor U6790 (N_6790,In_2448,In_2959);
nor U6791 (N_6791,In_1673,In_14);
and U6792 (N_6792,In_2537,In_2816);
or U6793 (N_6793,In_2579,In_310);
nor U6794 (N_6794,In_590,In_388);
nand U6795 (N_6795,In_1106,In_1445);
nand U6796 (N_6796,In_772,In_854);
or U6797 (N_6797,In_1655,In_2807);
or U6798 (N_6798,In_713,In_2101);
nand U6799 (N_6799,In_659,In_974);
or U6800 (N_6800,In_670,In_2543);
nor U6801 (N_6801,In_511,In_365);
or U6802 (N_6802,In_1185,In_1858);
nand U6803 (N_6803,In_1779,In_2028);
nor U6804 (N_6804,In_2961,In_1045);
nor U6805 (N_6805,In_2201,In_2024);
and U6806 (N_6806,In_1382,In_233);
nor U6807 (N_6807,In_1167,In_2487);
nand U6808 (N_6808,In_2113,In_1324);
nand U6809 (N_6809,In_324,In_742);
nand U6810 (N_6810,In_1809,In_1661);
xnor U6811 (N_6811,In_633,In_189);
or U6812 (N_6812,In_14,In_183);
or U6813 (N_6813,In_2209,In_2372);
nor U6814 (N_6814,In_2971,In_1078);
nor U6815 (N_6815,In_715,In_1686);
and U6816 (N_6816,In_548,In_673);
or U6817 (N_6817,In_1812,In_1987);
xnor U6818 (N_6818,In_1448,In_2698);
xor U6819 (N_6819,In_2269,In_836);
or U6820 (N_6820,In_747,In_708);
nor U6821 (N_6821,In_715,In_453);
xor U6822 (N_6822,In_2248,In_2412);
xnor U6823 (N_6823,In_2128,In_517);
or U6824 (N_6824,In_627,In_933);
nand U6825 (N_6825,In_2942,In_2675);
or U6826 (N_6826,In_2286,In_337);
and U6827 (N_6827,In_1376,In_904);
or U6828 (N_6828,In_830,In_2564);
xor U6829 (N_6829,In_425,In_294);
xor U6830 (N_6830,In_1606,In_1534);
or U6831 (N_6831,In_1474,In_953);
or U6832 (N_6832,In_191,In_255);
or U6833 (N_6833,In_105,In_2127);
nand U6834 (N_6834,In_1933,In_172);
nor U6835 (N_6835,In_914,In_2568);
nand U6836 (N_6836,In_467,In_887);
xnor U6837 (N_6837,In_1451,In_2429);
xor U6838 (N_6838,In_1008,In_2284);
or U6839 (N_6839,In_255,In_533);
xor U6840 (N_6840,In_1723,In_959);
nand U6841 (N_6841,In_1977,In_697);
xnor U6842 (N_6842,In_2018,In_299);
or U6843 (N_6843,In_1372,In_766);
nor U6844 (N_6844,In_1228,In_619);
xnor U6845 (N_6845,In_315,In_1015);
and U6846 (N_6846,In_2355,In_1208);
xnor U6847 (N_6847,In_654,In_478);
and U6848 (N_6848,In_985,In_1671);
nor U6849 (N_6849,In_222,In_2823);
nand U6850 (N_6850,In_1239,In_2281);
xor U6851 (N_6851,In_2813,In_924);
xnor U6852 (N_6852,In_1456,In_1910);
nor U6853 (N_6853,In_2399,In_623);
or U6854 (N_6854,In_984,In_529);
nand U6855 (N_6855,In_2166,In_1573);
nand U6856 (N_6856,In_2339,In_685);
nand U6857 (N_6857,In_748,In_1294);
or U6858 (N_6858,In_1160,In_2349);
xor U6859 (N_6859,In_616,In_1421);
xnor U6860 (N_6860,In_2211,In_527);
and U6861 (N_6861,In_1948,In_1705);
nand U6862 (N_6862,In_1055,In_2493);
and U6863 (N_6863,In_207,In_1674);
or U6864 (N_6864,In_1903,In_2941);
and U6865 (N_6865,In_554,In_2934);
and U6866 (N_6866,In_1330,In_342);
xor U6867 (N_6867,In_39,In_2205);
nand U6868 (N_6868,In_2088,In_1872);
and U6869 (N_6869,In_820,In_1441);
nand U6870 (N_6870,In_1710,In_2368);
xnor U6871 (N_6871,In_2508,In_36);
nand U6872 (N_6872,In_2968,In_1191);
and U6873 (N_6873,In_1444,In_1365);
xor U6874 (N_6874,In_93,In_1630);
nor U6875 (N_6875,In_2647,In_1245);
nor U6876 (N_6876,In_2763,In_2441);
and U6877 (N_6877,In_1199,In_68);
or U6878 (N_6878,In_2205,In_1304);
xor U6879 (N_6879,In_316,In_613);
nand U6880 (N_6880,In_478,In_2518);
nor U6881 (N_6881,In_635,In_472);
and U6882 (N_6882,In_1994,In_2694);
xor U6883 (N_6883,In_732,In_2384);
nand U6884 (N_6884,In_426,In_1367);
or U6885 (N_6885,In_898,In_1619);
and U6886 (N_6886,In_1983,In_176);
xor U6887 (N_6887,In_1901,In_583);
xnor U6888 (N_6888,In_1470,In_1063);
and U6889 (N_6889,In_1151,In_305);
or U6890 (N_6890,In_1954,In_562);
nor U6891 (N_6891,In_2839,In_1485);
nand U6892 (N_6892,In_944,In_1134);
nor U6893 (N_6893,In_2834,In_29);
and U6894 (N_6894,In_2625,In_453);
nand U6895 (N_6895,In_2922,In_2600);
nand U6896 (N_6896,In_2424,In_851);
and U6897 (N_6897,In_527,In_980);
xor U6898 (N_6898,In_1085,In_2286);
and U6899 (N_6899,In_2062,In_1277);
and U6900 (N_6900,In_885,In_1945);
or U6901 (N_6901,In_1107,In_2215);
nand U6902 (N_6902,In_1473,In_2774);
nor U6903 (N_6903,In_2256,In_2812);
and U6904 (N_6904,In_1895,In_930);
or U6905 (N_6905,In_2852,In_2969);
nor U6906 (N_6906,In_2361,In_1460);
xnor U6907 (N_6907,In_972,In_1897);
and U6908 (N_6908,In_2886,In_1164);
nand U6909 (N_6909,In_2350,In_2805);
nand U6910 (N_6910,In_1340,In_562);
nor U6911 (N_6911,In_2229,In_378);
nand U6912 (N_6912,In_1302,In_1526);
xnor U6913 (N_6913,In_2770,In_1285);
nor U6914 (N_6914,In_1842,In_1414);
nand U6915 (N_6915,In_2681,In_1758);
nor U6916 (N_6916,In_972,In_2119);
nor U6917 (N_6917,In_483,In_2074);
nand U6918 (N_6918,In_2397,In_1295);
nand U6919 (N_6919,In_86,In_2123);
or U6920 (N_6920,In_2664,In_2188);
and U6921 (N_6921,In_1019,In_2694);
and U6922 (N_6922,In_1919,In_1018);
or U6923 (N_6923,In_2582,In_2998);
nor U6924 (N_6924,In_2674,In_2006);
nor U6925 (N_6925,In_2803,In_693);
and U6926 (N_6926,In_983,In_2620);
xor U6927 (N_6927,In_271,In_1864);
and U6928 (N_6928,In_1012,In_1415);
xnor U6929 (N_6929,In_1417,In_1281);
or U6930 (N_6930,In_303,In_1025);
nand U6931 (N_6931,In_2656,In_2115);
xnor U6932 (N_6932,In_1307,In_1188);
or U6933 (N_6933,In_73,In_2901);
xnor U6934 (N_6934,In_2617,In_80);
or U6935 (N_6935,In_876,In_926);
and U6936 (N_6936,In_1299,In_85);
and U6937 (N_6937,In_2016,In_2170);
nand U6938 (N_6938,In_1597,In_2291);
xnor U6939 (N_6939,In_140,In_692);
and U6940 (N_6940,In_75,In_2790);
nand U6941 (N_6941,In_615,In_1229);
nand U6942 (N_6942,In_1511,In_1765);
xor U6943 (N_6943,In_2039,In_2230);
nand U6944 (N_6944,In_2255,In_977);
xor U6945 (N_6945,In_429,In_580);
and U6946 (N_6946,In_1562,In_1499);
and U6947 (N_6947,In_1115,In_1613);
nand U6948 (N_6948,In_2322,In_1614);
and U6949 (N_6949,In_2709,In_1553);
nand U6950 (N_6950,In_494,In_560);
or U6951 (N_6951,In_2285,In_1238);
nand U6952 (N_6952,In_1618,In_1602);
nor U6953 (N_6953,In_681,In_2795);
and U6954 (N_6954,In_1795,In_417);
nor U6955 (N_6955,In_2365,In_447);
xor U6956 (N_6956,In_821,In_871);
nor U6957 (N_6957,In_224,In_420);
nor U6958 (N_6958,In_2545,In_2937);
or U6959 (N_6959,In_346,In_1116);
nor U6960 (N_6960,In_2825,In_1384);
xnor U6961 (N_6961,In_1437,In_2189);
xnor U6962 (N_6962,In_1981,In_850);
nand U6963 (N_6963,In_1051,In_1454);
xnor U6964 (N_6964,In_1544,In_1309);
xnor U6965 (N_6965,In_799,In_147);
nand U6966 (N_6966,In_1286,In_517);
xor U6967 (N_6967,In_843,In_1220);
and U6968 (N_6968,In_2667,In_1811);
nor U6969 (N_6969,In_1868,In_256);
and U6970 (N_6970,In_2816,In_1925);
xnor U6971 (N_6971,In_313,In_1054);
xnor U6972 (N_6972,In_1464,In_707);
nor U6973 (N_6973,In_763,In_329);
and U6974 (N_6974,In_2103,In_1293);
or U6975 (N_6975,In_1438,In_1101);
or U6976 (N_6976,In_2627,In_594);
or U6977 (N_6977,In_2223,In_710);
or U6978 (N_6978,In_116,In_1507);
nor U6979 (N_6979,In_1228,In_1997);
xor U6980 (N_6980,In_1330,In_1655);
nor U6981 (N_6981,In_2787,In_2898);
and U6982 (N_6982,In_2830,In_2154);
xnor U6983 (N_6983,In_793,In_2707);
or U6984 (N_6984,In_79,In_980);
and U6985 (N_6985,In_1976,In_418);
nand U6986 (N_6986,In_1717,In_1564);
nand U6987 (N_6987,In_1871,In_1491);
or U6988 (N_6988,In_396,In_613);
nor U6989 (N_6989,In_1102,In_629);
nand U6990 (N_6990,In_1013,In_850);
or U6991 (N_6991,In_611,In_1015);
xor U6992 (N_6992,In_2069,In_2446);
nor U6993 (N_6993,In_2945,In_2650);
xnor U6994 (N_6994,In_873,In_2265);
and U6995 (N_6995,In_1471,In_724);
nor U6996 (N_6996,In_2081,In_2616);
and U6997 (N_6997,In_2733,In_1634);
or U6998 (N_6998,In_1352,In_2055);
xor U6999 (N_6999,In_2890,In_1074);
nor U7000 (N_7000,In_2730,In_601);
and U7001 (N_7001,In_644,In_403);
or U7002 (N_7002,In_421,In_1633);
xnor U7003 (N_7003,In_1007,In_1171);
and U7004 (N_7004,In_734,In_1417);
and U7005 (N_7005,In_2296,In_2375);
and U7006 (N_7006,In_2163,In_2220);
xor U7007 (N_7007,In_1153,In_787);
nand U7008 (N_7008,In_2228,In_2788);
nand U7009 (N_7009,In_1843,In_767);
nand U7010 (N_7010,In_277,In_2272);
or U7011 (N_7011,In_109,In_1916);
and U7012 (N_7012,In_2310,In_299);
and U7013 (N_7013,In_2842,In_1973);
nor U7014 (N_7014,In_1521,In_303);
nand U7015 (N_7015,In_2950,In_2693);
and U7016 (N_7016,In_813,In_2689);
xor U7017 (N_7017,In_2692,In_1640);
xnor U7018 (N_7018,In_1210,In_817);
nand U7019 (N_7019,In_1652,In_82);
or U7020 (N_7020,In_2717,In_1413);
and U7021 (N_7021,In_2273,In_2669);
nand U7022 (N_7022,In_2384,In_2438);
xor U7023 (N_7023,In_1113,In_322);
xor U7024 (N_7024,In_2420,In_2852);
xnor U7025 (N_7025,In_711,In_2034);
xnor U7026 (N_7026,In_952,In_1914);
nor U7027 (N_7027,In_1990,In_2595);
nand U7028 (N_7028,In_873,In_2055);
and U7029 (N_7029,In_80,In_1211);
or U7030 (N_7030,In_1501,In_11);
or U7031 (N_7031,In_406,In_1617);
and U7032 (N_7032,In_355,In_197);
or U7033 (N_7033,In_1284,In_59);
or U7034 (N_7034,In_1148,In_495);
nand U7035 (N_7035,In_1254,In_2087);
xnor U7036 (N_7036,In_151,In_2566);
and U7037 (N_7037,In_68,In_2615);
nor U7038 (N_7038,In_2509,In_227);
and U7039 (N_7039,In_352,In_1141);
nor U7040 (N_7040,In_1450,In_1525);
or U7041 (N_7041,In_487,In_1466);
or U7042 (N_7042,In_178,In_2762);
nand U7043 (N_7043,In_2254,In_573);
nand U7044 (N_7044,In_2005,In_2476);
or U7045 (N_7045,In_922,In_2859);
nand U7046 (N_7046,In_1516,In_971);
xnor U7047 (N_7047,In_378,In_1666);
or U7048 (N_7048,In_1883,In_613);
or U7049 (N_7049,In_10,In_67);
xor U7050 (N_7050,In_666,In_1712);
and U7051 (N_7051,In_2366,In_971);
nor U7052 (N_7052,In_2706,In_2423);
nor U7053 (N_7053,In_1469,In_1475);
nand U7054 (N_7054,In_1343,In_733);
nor U7055 (N_7055,In_1148,In_2297);
nor U7056 (N_7056,In_807,In_2656);
nand U7057 (N_7057,In_2321,In_819);
or U7058 (N_7058,In_907,In_1152);
nand U7059 (N_7059,In_1856,In_1504);
xor U7060 (N_7060,In_1603,In_2839);
or U7061 (N_7061,In_2593,In_2169);
nor U7062 (N_7062,In_1694,In_7);
nor U7063 (N_7063,In_77,In_810);
xor U7064 (N_7064,In_2431,In_1973);
nand U7065 (N_7065,In_1633,In_1249);
and U7066 (N_7066,In_173,In_248);
nor U7067 (N_7067,In_2466,In_553);
or U7068 (N_7068,In_524,In_321);
nor U7069 (N_7069,In_2400,In_6);
or U7070 (N_7070,In_2915,In_2653);
and U7071 (N_7071,In_2344,In_1546);
and U7072 (N_7072,In_483,In_33);
and U7073 (N_7073,In_1533,In_1996);
nand U7074 (N_7074,In_1189,In_1831);
or U7075 (N_7075,In_915,In_2753);
nor U7076 (N_7076,In_2762,In_273);
nand U7077 (N_7077,In_1500,In_1690);
and U7078 (N_7078,In_2892,In_1610);
and U7079 (N_7079,In_714,In_5);
xnor U7080 (N_7080,In_188,In_2561);
and U7081 (N_7081,In_1140,In_1687);
nand U7082 (N_7082,In_123,In_1521);
nand U7083 (N_7083,In_2077,In_2374);
nor U7084 (N_7084,In_125,In_624);
xnor U7085 (N_7085,In_2161,In_1768);
and U7086 (N_7086,In_1709,In_516);
nor U7087 (N_7087,In_2022,In_2667);
nand U7088 (N_7088,In_2396,In_1826);
nor U7089 (N_7089,In_2671,In_965);
nor U7090 (N_7090,In_1,In_780);
or U7091 (N_7091,In_865,In_2808);
nand U7092 (N_7092,In_19,In_2153);
or U7093 (N_7093,In_1237,In_373);
and U7094 (N_7094,In_2622,In_599);
xor U7095 (N_7095,In_355,In_1276);
nand U7096 (N_7096,In_1001,In_2495);
or U7097 (N_7097,In_2090,In_1047);
xnor U7098 (N_7098,In_2660,In_1019);
or U7099 (N_7099,In_586,In_1275);
and U7100 (N_7100,In_925,In_1565);
nand U7101 (N_7101,In_2704,In_2558);
or U7102 (N_7102,In_1153,In_1507);
xnor U7103 (N_7103,In_2694,In_1646);
nand U7104 (N_7104,In_652,In_2448);
nand U7105 (N_7105,In_1531,In_2133);
xor U7106 (N_7106,In_160,In_1828);
xor U7107 (N_7107,In_1481,In_1966);
and U7108 (N_7108,In_1030,In_57);
nand U7109 (N_7109,In_2299,In_2764);
nor U7110 (N_7110,In_590,In_1186);
xor U7111 (N_7111,In_1620,In_2854);
nor U7112 (N_7112,In_36,In_1843);
nand U7113 (N_7113,In_784,In_2665);
nand U7114 (N_7114,In_2955,In_1662);
nor U7115 (N_7115,In_2093,In_1006);
nand U7116 (N_7116,In_873,In_813);
or U7117 (N_7117,In_1337,In_2002);
nand U7118 (N_7118,In_1439,In_2102);
xor U7119 (N_7119,In_1951,In_2580);
xnor U7120 (N_7120,In_2473,In_538);
and U7121 (N_7121,In_2977,In_399);
xor U7122 (N_7122,In_1047,In_56);
xor U7123 (N_7123,In_2540,In_333);
nor U7124 (N_7124,In_1056,In_774);
nor U7125 (N_7125,In_1880,In_53);
nand U7126 (N_7126,In_599,In_612);
xor U7127 (N_7127,In_1714,In_2651);
nor U7128 (N_7128,In_2874,In_2397);
nor U7129 (N_7129,In_496,In_1415);
nand U7130 (N_7130,In_2882,In_2781);
nand U7131 (N_7131,In_2725,In_344);
and U7132 (N_7132,In_1980,In_198);
nor U7133 (N_7133,In_1251,In_2638);
xor U7134 (N_7134,In_1610,In_1901);
xnor U7135 (N_7135,In_2989,In_1671);
and U7136 (N_7136,In_756,In_2025);
nand U7137 (N_7137,In_1443,In_2421);
nor U7138 (N_7138,In_1719,In_2552);
and U7139 (N_7139,In_1342,In_222);
or U7140 (N_7140,In_1235,In_1694);
nor U7141 (N_7141,In_542,In_2511);
xnor U7142 (N_7142,In_2419,In_2835);
nor U7143 (N_7143,In_185,In_888);
and U7144 (N_7144,In_1741,In_862);
or U7145 (N_7145,In_324,In_2215);
nor U7146 (N_7146,In_2062,In_1306);
nor U7147 (N_7147,In_1220,In_2370);
xor U7148 (N_7148,In_592,In_1883);
and U7149 (N_7149,In_2544,In_1542);
nor U7150 (N_7150,In_45,In_2057);
or U7151 (N_7151,In_840,In_1186);
nand U7152 (N_7152,In_2791,In_1039);
and U7153 (N_7153,In_2520,In_2684);
nor U7154 (N_7154,In_1805,In_2736);
or U7155 (N_7155,In_921,In_2210);
xor U7156 (N_7156,In_1949,In_2260);
and U7157 (N_7157,In_712,In_434);
or U7158 (N_7158,In_351,In_1568);
nor U7159 (N_7159,In_2269,In_1354);
nor U7160 (N_7160,In_2878,In_2308);
or U7161 (N_7161,In_1466,In_1860);
xor U7162 (N_7162,In_233,In_632);
and U7163 (N_7163,In_1033,In_2220);
xor U7164 (N_7164,In_1467,In_504);
xnor U7165 (N_7165,In_1867,In_1168);
and U7166 (N_7166,In_253,In_162);
nand U7167 (N_7167,In_1106,In_2633);
and U7168 (N_7168,In_954,In_1999);
nand U7169 (N_7169,In_447,In_1332);
nand U7170 (N_7170,In_2579,In_621);
and U7171 (N_7171,In_2468,In_877);
nor U7172 (N_7172,In_1258,In_2591);
nor U7173 (N_7173,In_1688,In_2684);
and U7174 (N_7174,In_2555,In_1763);
nor U7175 (N_7175,In_2236,In_2554);
nand U7176 (N_7176,In_1893,In_1577);
nand U7177 (N_7177,In_289,In_209);
or U7178 (N_7178,In_773,In_1522);
xor U7179 (N_7179,In_2424,In_1381);
nand U7180 (N_7180,In_1469,In_439);
xnor U7181 (N_7181,In_2550,In_968);
and U7182 (N_7182,In_2701,In_2335);
nand U7183 (N_7183,In_2183,In_512);
and U7184 (N_7184,In_1793,In_777);
nor U7185 (N_7185,In_1135,In_2605);
xor U7186 (N_7186,In_2867,In_81);
nand U7187 (N_7187,In_571,In_2885);
and U7188 (N_7188,In_1069,In_1809);
nand U7189 (N_7189,In_2660,In_716);
and U7190 (N_7190,In_2734,In_375);
and U7191 (N_7191,In_849,In_1053);
and U7192 (N_7192,In_2173,In_2616);
nor U7193 (N_7193,In_1073,In_877);
and U7194 (N_7194,In_2353,In_1278);
nand U7195 (N_7195,In_930,In_327);
xnor U7196 (N_7196,In_589,In_2672);
nor U7197 (N_7197,In_837,In_1685);
xor U7198 (N_7198,In_366,In_1516);
xnor U7199 (N_7199,In_562,In_484);
nand U7200 (N_7200,In_2518,In_1787);
or U7201 (N_7201,In_1211,In_2581);
and U7202 (N_7202,In_259,In_2114);
nor U7203 (N_7203,In_508,In_642);
and U7204 (N_7204,In_2422,In_2592);
nor U7205 (N_7205,In_1351,In_422);
nor U7206 (N_7206,In_1065,In_524);
xor U7207 (N_7207,In_1540,In_350);
or U7208 (N_7208,In_497,In_1264);
xor U7209 (N_7209,In_1166,In_2928);
xnor U7210 (N_7210,In_468,In_2703);
xor U7211 (N_7211,In_1957,In_2072);
nand U7212 (N_7212,In_817,In_2342);
nor U7213 (N_7213,In_1276,In_2069);
and U7214 (N_7214,In_1104,In_1359);
nor U7215 (N_7215,In_540,In_1107);
nand U7216 (N_7216,In_2413,In_1287);
nor U7217 (N_7217,In_2325,In_2830);
nor U7218 (N_7218,In_2530,In_1345);
xnor U7219 (N_7219,In_2344,In_1176);
nand U7220 (N_7220,In_1893,In_470);
nor U7221 (N_7221,In_316,In_388);
xor U7222 (N_7222,In_2367,In_1976);
nor U7223 (N_7223,In_1236,In_2130);
or U7224 (N_7224,In_2369,In_2315);
nor U7225 (N_7225,In_1536,In_1837);
xor U7226 (N_7226,In_455,In_2983);
xnor U7227 (N_7227,In_641,In_1055);
xnor U7228 (N_7228,In_1245,In_2120);
and U7229 (N_7229,In_352,In_2070);
xnor U7230 (N_7230,In_2522,In_1848);
or U7231 (N_7231,In_2384,In_1243);
or U7232 (N_7232,In_2268,In_1249);
or U7233 (N_7233,In_895,In_2651);
nor U7234 (N_7234,In_881,In_2692);
xnor U7235 (N_7235,In_2944,In_1246);
nand U7236 (N_7236,In_1493,In_2083);
and U7237 (N_7237,In_1089,In_1739);
or U7238 (N_7238,In_790,In_2336);
and U7239 (N_7239,In_932,In_1393);
nor U7240 (N_7240,In_625,In_1405);
and U7241 (N_7241,In_2023,In_100);
nand U7242 (N_7242,In_376,In_1069);
or U7243 (N_7243,In_2592,In_1183);
nor U7244 (N_7244,In_2398,In_2714);
nand U7245 (N_7245,In_2174,In_2318);
nand U7246 (N_7246,In_1980,In_2927);
or U7247 (N_7247,In_486,In_1970);
nand U7248 (N_7248,In_255,In_1055);
nand U7249 (N_7249,In_650,In_110);
xnor U7250 (N_7250,In_2933,In_1112);
nor U7251 (N_7251,In_2320,In_1080);
or U7252 (N_7252,In_1960,In_2348);
or U7253 (N_7253,In_1276,In_2795);
nor U7254 (N_7254,In_2563,In_793);
nand U7255 (N_7255,In_1760,In_258);
xor U7256 (N_7256,In_1664,In_2834);
nand U7257 (N_7257,In_1751,In_799);
xnor U7258 (N_7258,In_889,In_2303);
xor U7259 (N_7259,In_1459,In_2153);
nand U7260 (N_7260,In_2702,In_2891);
xnor U7261 (N_7261,In_2040,In_1494);
nand U7262 (N_7262,In_1203,In_602);
or U7263 (N_7263,In_2345,In_76);
or U7264 (N_7264,In_232,In_147);
and U7265 (N_7265,In_351,In_1005);
xnor U7266 (N_7266,In_2284,In_2949);
and U7267 (N_7267,In_1318,In_1486);
nand U7268 (N_7268,In_1943,In_1529);
nand U7269 (N_7269,In_1045,In_805);
or U7270 (N_7270,In_15,In_880);
xnor U7271 (N_7271,In_2165,In_294);
nand U7272 (N_7272,In_2458,In_561);
nor U7273 (N_7273,In_1487,In_171);
nor U7274 (N_7274,In_161,In_491);
nor U7275 (N_7275,In_421,In_1555);
nand U7276 (N_7276,In_2896,In_2674);
and U7277 (N_7277,In_1458,In_433);
nand U7278 (N_7278,In_1286,In_1459);
and U7279 (N_7279,In_1518,In_808);
nand U7280 (N_7280,In_1253,In_2268);
nand U7281 (N_7281,In_1273,In_1247);
nor U7282 (N_7282,In_2882,In_1686);
and U7283 (N_7283,In_1298,In_546);
xnor U7284 (N_7284,In_1118,In_2453);
and U7285 (N_7285,In_970,In_1425);
or U7286 (N_7286,In_2094,In_808);
nor U7287 (N_7287,In_1932,In_19);
nor U7288 (N_7288,In_1360,In_402);
and U7289 (N_7289,In_2802,In_629);
nor U7290 (N_7290,In_1965,In_2458);
and U7291 (N_7291,In_2641,In_339);
nand U7292 (N_7292,In_1605,In_1125);
xnor U7293 (N_7293,In_1804,In_2327);
xnor U7294 (N_7294,In_1302,In_27);
xnor U7295 (N_7295,In_2084,In_1965);
xor U7296 (N_7296,In_839,In_15);
or U7297 (N_7297,In_2421,In_1807);
and U7298 (N_7298,In_2640,In_2518);
xnor U7299 (N_7299,In_160,In_2314);
xnor U7300 (N_7300,In_259,In_2700);
xnor U7301 (N_7301,In_2063,In_1391);
and U7302 (N_7302,In_2390,In_1486);
nor U7303 (N_7303,In_2777,In_524);
nor U7304 (N_7304,In_1287,In_1719);
xor U7305 (N_7305,In_757,In_2754);
or U7306 (N_7306,In_2457,In_847);
or U7307 (N_7307,In_16,In_814);
nand U7308 (N_7308,In_1201,In_2531);
nor U7309 (N_7309,In_274,In_2986);
or U7310 (N_7310,In_954,In_1448);
and U7311 (N_7311,In_1345,In_2934);
or U7312 (N_7312,In_1690,In_2787);
xnor U7313 (N_7313,In_310,In_1289);
nand U7314 (N_7314,In_117,In_1618);
and U7315 (N_7315,In_2279,In_2118);
or U7316 (N_7316,In_624,In_737);
xnor U7317 (N_7317,In_2202,In_1567);
or U7318 (N_7318,In_2835,In_231);
nor U7319 (N_7319,In_1378,In_1677);
and U7320 (N_7320,In_1603,In_1327);
and U7321 (N_7321,In_1845,In_2483);
xor U7322 (N_7322,In_72,In_1119);
nor U7323 (N_7323,In_507,In_2122);
xor U7324 (N_7324,In_1236,In_953);
xor U7325 (N_7325,In_2551,In_1910);
xor U7326 (N_7326,In_827,In_2525);
and U7327 (N_7327,In_2562,In_2896);
or U7328 (N_7328,In_214,In_2698);
nand U7329 (N_7329,In_2225,In_229);
nand U7330 (N_7330,In_2180,In_2153);
xor U7331 (N_7331,In_511,In_578);
and U7332 (N_7332,In_2916,In_439);
and U7333 (N_7333,In_1927,In_1283);
or U7334 (N_7334,In_1155,In_1447);
or U7335 (N_7335,In_1951,In_2743);
nor U7336 (N_7336,In_2109,In_1468);
or U7337 (N_7337,In_2083,In_2483);
or U7338 (N_7338,In_374,In_2478);
xor U7339 (N_7339,In_2450,In_125);
nor U7340 (N_7340,In_386,In_231);
xor U7341 (N_7341,In_371,In_529);
and U7342 (N_7342,In_2346,In_2310);
and U7343 (N_7343,In_1882,In_2724);
xnor U7344 (N_7344,In_2958,In_2575);
and U7345 (N_7345,In_1767,In_1831);
nor U7346 (N_7346,In_1135,In_48);
and U7347 (N_7347,In_555,In_2983);
xnor U7348 (N_7348,In_2509,In_1801);
or U7349 (N_7349,In_756,In_1070);
xnor U7350 (N_7350,In_1686,In_1729);
and U7351 (N_7351,In_118,In_86);
nor U7352 (N_7352,In_116,In_790);
xor U7353 (N_7353,In_134,In_2632);
nand U7354 (N_7354,In_1660,In_948);
and U7355 (N_7355,In_585,In_461);
and U7356 (N_7356,In_1052,In_1873);
nand U7357 (N_7357,In_857,In_2091);
or U7358 (N_7358,In_657,In_495);
and U7359 (N_7359,In_497,In_579);
and U7360 (N_7360,In_1823,In_2498);
and U7361 (N_7361,In_1802,In_2125);
xor U7362 (N_7362,In_1264,In_1880);
and U7363 (N_7363,In_2266,In_1482);
nor U7364 (N_7364,In_841,In_191);
xnor U7365 (N_7365,In_78,In_108);
nand U7366 (N_7366,In_2666,In_296);
nor U7367 (N_7367,In_1350,In_669);
nand U7368 (N_7368,In_1953,In_2681);
or U7369 (N_7369,In_1943,In_1266);
xnor U7370 (N_7370,In_1496,In_917);
xor U7371 (N_7371,In_104,In_2713);
xnor U7372 (N_7372,In_2643,In_792);
nor U7373 (N_7373,In_2229,In_1031);
and U7374 (N_7374,In_1824,In_2266);
nand U7375 (N_7375,In_246,In_1500);
and U7376 (N_7376,In_2147,In_57);
nand U7377 (N_7377,In_2565,In_1877);
nand U7378 (N_7378,In_244,In_2343);
nor U7379 (N_7379,In_1137,In_467);
or U7380 (N_7380,In_1559,In_336);
or U7381 (N_7381,In_2764,In_148);
nor U7382 (N_7382,In_604,In_2012);
xor U7383 (N_7383,In_213,In_1705);
nor U7384 (N_7384,In_225,In_749);
nand U7385 (N_7385,In_1082,In_993);
or U7386 (N_7386,In_2851,In_908);
nor U7387 (N_7387,In_2710,In_1090);
nor U7388 (N_7388,In_72,In_1584);
nand U7389 (N_7389,In_809,In_799);
or U7390 (N_7390,In_225,In_1431);
nand U7391 (N_7391,In_2848,In_535);
nand U7392 (N_7392,In_731,In_2226);
and U7393 (N_7393,In_1708,In_576);
and U7394 (N_7394,In_446,In_25);
and U7395 (N_7395,In_163,In_2832);
xor U7396 (N_7396,In_916,In_2201);
nand U7397 (N_7397,In_447,In_2203);
nand U7398 (N_7398,In_1479,In_2322);
or U7399 (N_7399,In_2601,In_2513);
nor U7400 (N_7400,In_2187,In_2305);
xnor U7401 (N_7401,In_2628,In_1854);
nor U7402 (N_7402,In_1698,In_982);
xnor U7403 (N_7403,In_2226,In_318);
nor U7404 (N_7404,In_1964,In_473);
and U7405 (N_7405,In_2743,In_805);
or U7406 (N_7406,In_2416,In_2965);
and U7407 (N_7407,In_2383,In_2874);
nand U7408 (N_7408,In_721,In_204);
nor U7409 (N_7409,In_1958,In_344);
nor U7410 (N_7410,In_2150,In_1121);
nand U7411 (N_7411,In_2413,In_444);
and U7412 (N_7412,In_1619,In_241);
or U7413 (N_7413,In_1051,In_1202);
and U7414 (N_7414,In_2872,In_535);
nand U7415 (N_7415,In_2819,In_429);
nand U7416 (N_7416,In_922,In_2210);
nor U7417 (N_7417,In_1352,In_414);
nand U7418 (N_7418,In_1219,In_938);
nand U7419 (N_7419,In_1162,In_2409);
and U7420 (N_7420,In_2396,In_1291);
nor U7421 (N_7421,In_782,In_764);
xnor U7422 (N_7422,In_2018,In_2359);
or U7423 (N_7423,In_1469,In_290);
nor U7424 (N_7424,In_1402,In_2127);
and U7425 (N_7425,In_880,In_2203);
nand U7426 (N_7426,In_2936,In_1837);
xor U7427 (N_7427,In_1187,In_716);
and U7428 (N_7428,In_352,In_544);
nor U7429 (N_7429,In_2147,In_2451);
nand U7430 (N_7430,In_2971,In_2424);
nor U7431 (N_7431,In_2709,In_4);
nand U7432 (N_7432,In_1674,In_2302);
nor U7433 (N_7433,In_2064,In_1095);
and U7434 (N_7434,In_291,In_1137);
or U7435 (N_7435,In_778,In_124);
nor U7436 (N_7436,In_2779,In_2071);
xor U7437 (N_7437,In_2430,In_1398);
xnor U7438 (N_7438,In_54,In_1337);
nand U7439 (N_7439,In_1055,In_769);
nor U7440 (N_7440,In_2702,In_2156);
xnor U7441 (N_7441,In_203,In_931);
nand U7442 (N_7442,In_571,In_704);
xor U7443 (N_7443,In_1694,In_1101);
and U7444 (N_7444,In_104,In_520);
and U7445 (N_7445,In_1482,In_987);
nor U7446 (N_7446,In_328,In_609);
nand U7447 (N_7447,In_557,In_1299);
and U7448 (N_7448,In_2363,In_1011);
xnor U7449 (N_7449,In_557,In_603);
or U7450 (N_7450,In_1875,In_956);
or U7451 (N_7451,In_709,In_150);
or U7452 (N_7452,In_2231,In_2062);
nand U7453 (N_7453,In_2249,In_2651);
nand U7454 (N_7454,In_1977,In_2083);
xor U7455 (N_7455,In_1429,In_1216);
and U7456 (N_7456,In_74,In_2371);
or U7457 (N_7457,In_960,In_1173);
and U7458 (N_7458,In_723,In_2178);
nand U7459 (N_7459,In_657,In_1291);
nor U7460 (N_7460,In_485,In_1878);
nor U7461 (N_7461,In_2948,In_862);
nand U7462 (N_7462,In_310,In_10);
xnor U7463 (N_7463,In_260,In_2435);
and U7464 (N_7464,In_1172,In_2190);
and U7465 (N_7465,In_1158,In_2575);
or U7466 (N_7466,In_480,In_624);
and U7467 (N_7467,In_727,In_2684);
nor U7468 (N_7468,In_645,In_2503);
or U7469 (N_7469,In_2260,In_2919);
or U7470 (N_7470,In_2431,In_668);
xor U7471 (N_7471,In_769,In_1251);
nand U7472 (N_7472,In_2328,In_1913);
or U7473 (N_7473,In_1357,In_2915);
nor U7474 (N_7474,In_1624,In_1701);
and U7475 (N_7475,In_2188,In_156);
xor U7476 (N_7476,In_2405,In_2107);
xor U7477 (N_7477,In_1095,In_1395);
nor U7478 (N_7478,In_2006,In_2171);
nand U7479 (N_7479,In_1048,In_2812);
or U7480 (N_7480,In_1389,In_2942);
nor U7481 (N_7481,In_1932,In_1276);
nand U7482 (N_7482,In_381,In_920);
and U7483 (N_7483,In_2472,In_2029);
nor U7484 (N_7484,In_1712,In_626);
or U7485 (N_7485,In_2916,In_154);
nand U7486 (N_7486,In_963,In_189);
nor U7487 (N_7487,In_840,In_1815);
nand U7488 (N_7488,In_2167,In_2432);
nand U7489 (N_7489,In_1721,In_582);
xor U7490 (N_7490,In_2389,In_1132);
nand U7491 (N_7491,In_1500,In_768);
nand U7492 (N_7492,In_1013,In_1164);
nand U7493 (N_7493,In_1309,In_747);
xor U7494 (N_7494,In_2485,In_1635);
nand U7495 (N_7495,In_204,In_660);
nor U7496 (N_7496,In_54,In_2898);
xnor U7497 (N_7497,In_9,In_2543);
nor U7498 (N_7498,In_1766,In_2808);
nor U7499 (N_7499,In_2809,In_2603);
xor U7500 (N_7500,In_1717,In_2516);
or U7501 (N_7501,In_2446,In_2697);
nor U7502 (N_7502,In_2028,In_1610);
nand U7503 (N_7503,In_1199,In_1108);
xor U7504 (N_7504,In_1750,In_713);
nor U7505 (N_7505,In_859,In_1326);
or U7506 (N_7506,In_2465,In_1685);
or U7507 (N_7507,In_1227,In_2094);
nand U7508 (N_7508,In_1217,In_2105);
nor U7509 (N_7509,In_2622,In_1474);
and U7510 (N_7510,In_2661,In_923);
xnor U7511 (N_7511,In_1070,In_475);
nor U7512 (N_7512,In_2607,In_2741);
or U7513 (N_7513,In_2471,In_2519);
nor U7514 (N_7514,In_2395,In_2169);
or U7515 (N_7515,In_1524,In_962);
nand U7516 (N_7516,In_844,In_2018);
nor U7517 (N_7517,In_2846,In_880);
xor U7518 (N_7518,In_531,In_1195);
nor U7519 (N_7519,In_1991,In_1960);
or U7520 (N_7520,In_645,In_1351);
nand U7521 (N_7521,In_1314,In_631);
xnor U7522 (N_7522,In_1415,In_2949);
and U7523 (N_7523,In_2699,In_1619);
xor U7524 (N_7524,In_324,In_1398);
xor U7525 (N_7525,In_1900,In_1882);
nor U7526 (N_7526,In_925,In_621);
nor U7527 (N_7527,In_1679,In_1350);
nor U7528 (N_7528,In_2678,In_2003);
nor U7529 (N_7529,In_1663,In_37);
and U7530 (N_7530,In_2452,In_2845);
xor U7531 (N_7531,In_2066,In_2264);
nand U7532 (N_7532,In_1784,In_2049);
or U7533 (N_7533,In_503,In_1583);
and U7534 (N_7534,In_2232,In_1810);
and U7535 (N_7535,In_298,In_2022);
nor U7536 (N_7536,In_2119,In_1161);
and U7537 (N_7537,In_406,In_392);
or U7538 (N_7538,In_776,In_740);
xnor U7539 (N_7539,In_1679,In_1751);
xor U7540 (N_7540,In_1314,In_1958);
xnor U7541 (N_7541,In_1275,In_1157);
xor U7542 (N_7542,In_2218,In_456);
or U7543 (N_7543,In_260,In_1368);
nand U7544 (N_7544,In_768,In_802);
xor U7545 (N_7545,In_1609,In_2366);
or U7546 (N_7546,In_572,In_2242);
nor U7547 (N_7547,In_2144,In_1318);
nor U7548 (N_7548,In_661,In_150);
xor U7549 (N_7549,In_182,In_2622);
xor U7550 (N_7550,In_4,In_173);
nand U7551 (N_7551,In_1902,In_1835);
nand U7552 (N_7552,In_267,In_1571);
or U7553 (N_7553,In_1599,In_2459);
or U7554 (N_7554,In_2069,In_57);
nor U7555 (N_7555,In_422,In_1027);
nor U7556 (N_7556,In_232,In_2751);
or U7557 (N_7557,In_2979,In_344);
nor U7558 (N_7558,In_305,In_2904);
nor U7559 (N_7559,In_2226,In_2615);
nand U7560 (N_7560,In_187,In_1975);
nor U7561 (N_7561,In_1697,In_2848);
and U7562 (N_7562,In_1059,In_2429);
and U7563 (N_7563,In_643,In_955);
xnor U7564 (N_7564,In_89,In_1757);
or U7565 (N_7565,In_916,In_1226);
xor U7566 (N_7566,In_2284,In_2602);
nand U7567 (N_7567,In_2739,In_1349);
and U7568 (N_7568,In_1591,In_1043);
nor U7569 (N_7569,In_754,In_2495);
and U7570 (N_7570,In_730,In_231);
xnor U7571 (N_7571,In_2006,In_1643);
and U7572 (N_7572,In_1311,In_1860);
xor U7573 (N_7573,In_1127,In_1541);
nand U7574 (N_7574,In_1381,In_1293);
nor U7575 (N_7575,In_2937,In_2464);
xnor U7576 (N_7576,In_1886,In_1291);
and U7577 (N_7577,In_854,In_396);
xnor U7578 (N_7578,In_1300,In_2107);
xor U7579 (N_7579,In_2330,In_2462);
nor U7580 (N_7580,In_1534,In_1805);
nand U7581 (N_7581,In_2494,In_1343);
nand U7582 (N_7582,In_394,In_230);
and U7583 (N_7583,In_2618,In_1265);
and U7584 (N_7584,In_2103,In_1879);
or U7585 (N_7585,In_1554,In_1078);
and U7586 (N_7586,In_2012,In_26);
or U7587 (N_7587,In_2896,In_2947);
xnor U7588 (N_7588,In_311,In_1058);
nand U7589 (N_7589,In_2495,In_2257);
and U7590 (N_7590,In_873,In_2644);
xnor U7591 (N_7591,In_1641,In_463);
nor U7592 (N_7592,In_1973,In_412);
nor U7593 (N_7593,In_1979,In_606);
and U7594 (N_7594,In_1737,In_1154);
and U7595 (N_7595,In_367,In_2537);
nand U7596 (N_7596,In_2149,In_2924);
nand U7597 (N_7597,In_1420,In_1566);
xor U7598 (N_7598,In_861,In_1964);
nor U7599 (N_7599,In_282,In_1967);
xor U7600 (N_7600,In_1047,In_1622);
nand U7601 (N_7601,In_327,In_1734);
and U7602 (N_7602,In_1888,In_711);
xor U7603 (N_7603,In_2524,In_967);
nand U7604 (N_7604,In_433,In_949);
and U7605 (N_7605,In_1830,In_1405);
nor U7606 (N_7606,In_962,In_2031);
xor U7607 (N_7607,In_138,In_1693);
and U7608 (N_7608,In_1479,In_2938);
and U7609 (N_7609,In_383,In_2694);
and U7610 (N_7610,In_1135,In_1780);
and U7611 (N_7611,In_2595,In_1015);
or U7612 (N_7612,In_297,In_2477);
or U7613 (N_7613,In_1858,In_1258);
xor U7614 (N_7614,In_1661,In_2917);
xnor U7615 (N_7615,In_1517,In_1229);
nand U7616 (N_7616,In_2855,In_217);
and U7617 (N_7617,In_2978,In_2252);
xnor U7618 (N_7618,In_1392,In_775);
nor U7619 (N_7619,In_400,In_2786);
and U7620 (N_7620,In_2791,In_2523);
xnor U7621 (N_7621,In_989,In_2734);
and U7622 (N_7622,In_2781,In_1407);
and U7623 (N_7623,In_1367,In_1223);
and U7624 (N_7624,In_759,In_1346);
nor U7625 (N_7625,In_1843,In_2743);
and U7626 (N_7626,In_1670,In_973);
and U7627 (N_7627,In_1672,In_2120);
or U7628 (N_7628,In_768,In_1376);
or U7629 (N_7629,In_1599,In_209);
nand U7630 (N_7630,In_674,In_2284);
or U7631 (N_7631,In_979,In_1255);
and U7632 (N_7632,In_2705,In_2841);
and U7633 (N_7633,In_392,In_2161);
and U7634 (N_7634,In_1673,In_2883);
nor U7635 (N_7635,In_86,In_1399);
nand U7636 (N_7636,In_353,In_1205);
or U7637 (N_7637,In_794,In_1840);
nand U7638 (N_7638,In_668,In_1675);
nand U7639 (N_7639,In_1923,In_1498);
nand U7640 (N_7640,In_1948,In_235);
or U7641 (N_7641,In_235,In_1061);
or U7642 (N_7642,In_2900,In_1773);
xor U7643 (N_7643,In_2692,In_2458);
nor U7644 (N_7644,In_2856,In_2509);
nor U7645 (N_7645,In_117,In_30);
nand U7646 (N_7646,In_2305,In_2185);
or U7647 (N_7647,In_2440,In_234);
or U7648 (N_7648,In_2005,In_1857);
nand U7649 (N_7649,In_429,In_2454);
nand U7650 (N_7650,In_1490,In_383);
and U7651 (N_7651,In_2130,In_2233);
nor U7652 (N_7652,In_2134,In_1020);
and U7653 (N_7653,In_369,In_2279);
xor U7654 (N_7654,In_24,In_2906);
xnor U7655 (N_7655,In_616,In_1312);
nor U7656 (N_7656,In_1966,In_601);
xnor U7657 (N_7657,In_10,In_917);
or U7658 (N_7658,In_325,In_941);
nor U7659 (N_7659,In_1898,In_1499);
and U7660 (N_7660,In_1969,In_1817);
or U7661 (N_7661,In_2752,In_902);
xor U7662 (N_7662,In_1285,In_1850);
nor U7663 (N_7663,In_662,In_1322);
nor U7664 (N_7664,In_1751,In_1165);
nor U7665 (N_7665,In_2737,In_536);
and U7666 (N_7666,In_1606,In_843);
or U7667 (N_7667,In_2993,In_1517);
and U7668 (N_7668,In_340,In_1564);
nand U7669 (N_7669,In_2853,In_2868);
nand U7670 (N_7670,In_2091,In_2997);
nor U7671 (N_7671,In_1977,In_858);
xor U7672 (N_7672,In_160,In_2820);
nand U7673 (N_7673,In_462,In_72);
and U7674 (N_7674,In_857,In_2388);
xor U7675 (N_7675,In_862,In_1282);
and U7676 (N_7676,In_1454,In_2586);
nor U7677 (N_7677,In_951,In_1236);
nor U7678 (N_7678,In_2223,In_1810);
nor U7679 (N_7679,In_1342,In_1807);
nand U7680 (N_7680,In_2578,In_156);
nor U7681 (N_7681,In_948,In_2303);
nand U7682 (N_7682,In_843,In_485);
nand U7683 (N_7683,In_1271,In_1481);
nand U7684 (N_7684,In_1292,In_75);
nor U7685 (N_7685,In_1645,In_2370);
and U7686 (N_7686,In_2464,In_725);
and U7687 (N_7687,In_1559,In_2670);
and U7688 (N_7688,In_283,In_2704);
or U7689 (N_7689,In_142,In_1420);
nor U7690 (N_7690,In_917,In_1146);
nor U7691 (N_7691,In_2422,In_1954);
or U7692 (N_7692,In_2245,In_1183);
or U7693 (N_7693,In_802,In_1024);
nor U7694 (N_7694,In_1504,In_431);
nand U7695 (N_7695,In_2421,In_2500);
nor U7696 (N_7696,In_1939,In_2154);
nor U7697 (N_7697,In_871,In_179);
nor U7698 (N_7698,In_371,In_2591);
nand U7699 (N_7699,In_1798,In_2124);
nor U7700 (N_7700,In_2685,In_1210);
xnor U7701 (N_7701,In_983,In_2664);
nand U7702 (N_7702,In_97,In_2675);
and U7703 (N_7703,In_1172,In_548);
xnor U7704 (N_7704,In_9,In_1696);
nand U7705 (N_7705,In_1464,In_1637);
and U7706 (N_7706,In_2861,In_2268);
nor U7707 (N_7707,In_1423,In_2487);
xor U7708 (N_7708,In_1208,In_2942);
xor U7709 (N_7709,In_1449,In_11);
nor U7710 (N_7710,In_1919,In_10);
nand U7711 (N_7711,In_1419,In_2580);
xnor U7712 (N_7712,In_2259,In_1907);
or U7713 (N_7713,In_1131,In_1513);
xnor U7714 (N_7714,In_1269,In_1208);
nand U7715 (N_7715,In_396,In_1830);
nor U7716 (N_7716,In_675,In_1938);
nor U7717 (N_7717,In_2838,In_2225);
nor U7718 (N_7718,In_2018,In_1691);
xnor U7719 (N_7719,In_155,In_926);
nand U7720 (N_7720,In_1972,In_440);
xnor U7721 (N_7721,In_2775,In_5);
or U7722 (N_7722,In_2993,In_1134);
xnor U7723 (N_7723,In_1389,In_2912);
or U7724 (N_7724,In_97,In_786);
and U7725 (N_7725,In_545,In_166);
and U7726 (N_7726,In_1316,In_2855);
nor U7727 (N_7727,In_2025,In_1718);
nor U7728 (N_7728,In_2703,In_2963);
nand U7729 (N_7729,In_898,In_352);
xor U7730 (N_7730,In_1103,In_1333);
and U7731 (N_7731,In_2385,In_1681);
or U7732 (N_7732,In_2829,In_2792);
nand U7733 (N_7733,In_1370,In_2895);
or U7734 (N_7734,In_2272,In_2901);
and U7735 (N_7735,In_857,In_1054);
or U7736 (N_7736,In_1129,In_372);
nand U7737 (N_7737,In_822,In_256);
and U7738 (N_7738,In_1476,In_2897);
xor U7739 (N_7739,In_1726,In_415);
nor U7740 (N_7740,In_1728,In_2829);
and U7741 (N_7741,In_521,In_1592);
and U7742 (N_7742,In_2001,In_866);
and U7743 (N_7743,In_2733,In_2033);
nand U7744 (N_7744,In_1704,In_1752);
nor U7745 (N_7745,In_2334,In_1727);
nand U7746 (N_7746,In_1975,In_1841);
nand U7747 (N_7747,In_734,In_337);
nor U7748 (N_7748,In_1552,In_257);
and U7749 (N_7749,In_383,In_1131);
xnor U7750 (N_7750,In_78,In_1288);
or U7751 (N_7751,In_2249,In_499);
nor U7752 (N_7752,In_1519,In_1828);
xor U7753 (N_7753,In_2103,In_2870);
nor U7754 (N_7754,In_1722,In_2732);
and U7755 (N_7755,In_2939,In_958);
nand U7756 (N_7756,In_382,In_1039);
or U7757 (N_7757,In_502,In_1732);
nor U7758 (N_7758,In_2233,In_1076);
nand U7759 (N_7759,In_2563,In_676);
nor U7760 (N_7760,In_1927,In_2392);
and U7761 (N_7761,In_1988,In_1207);
xor U7762 (N_7762,In_1927,In_1835);
nor U7763 (N_7763,In_2131,In_212);
xnor U7764 (N_7764,In_1887,In_2140);
nor U7765 (N_7765,In_1000,In_647);
nor U7766 (N_7766,In_14,In_1374);
and U7767 (N_7767,In_1288,In_2739);
and U7768 (N_7768,In_1025,In_961);
and U7769 (N_7769,In_1894,In_2952);
or U7770 (N_7770,In_780,In_2850);
or U7771 (N_7771,In_314,In_552);
or U7772 (N_7772,In_1386,In_2461);
xor U7773 (N_7773,In_845,In_1823);
and U7774 (N_7774,In_1518,In_1093);
nand U7775 (N_7775,In_2624,In_774);
xor U7776 (N_7776,In_1023,In_2666);
and U7777 (N_7777,In_2734,In_2357);
or U7778 (N_7778,In_900,In_1691);
and U7779 (N_7779,In_2519,In_1590);
or U7780 (N_7780,In_1413,In_2482);
or U7781 (N_7781,In_1639,In_372);
or U7782 (N_7782,In_2407,In_1286);
nand U7783 (N_7783,In_2857,In_273);
xor U7784 (N_7784,In_2758,In_356);
nor U7785 (N_7785,In_2138,In_612);
or U7786 (N_7786,In_580,In_172);
nand U7787 (N_7787,In_2810,In_2435);
or U7788 (N_7788,In_1615,In_452);
nand U7789 (N_7789,In_1266,In_2079);
xor U7790 (N_7790,In_1658,In_1129);
and U7791 (N_7791,In_2027,In_1981);
xnor U7792 (N_7792,In_583,In_1497);
nand U7793 (N_7793,In_191,In_2291);
nand U7794 (N_7794,In_699,In_1316);
nor U7795 (N_7795,In_1240,In_1273);
nor U7796 (N_7796,In_2795,In_1173);
or U7797 (N_7797,In_718,In_591);
nand U7798 (N_7798,In_511,In_2847);
xor U7799 (N_7799,In_889,In_2701);
xor U7800 (N_7800,In_1254,In_2231);
xnor U7801 (N_7801,In_1650,In_103);
xnor U7802 (N_7802,In_2287,In_513);
or U7803 (N_7803,In_2747,In_722);
and U7804 (N_7804,In_2936,In_83);
and U7805 (N_7805,In_2127,In_3);
and U7806 (N_7806,In_1136,In_464);
nand U7807 (N_7807,In_178,In_1839);
xor U7808 (N_7808,In_2749,In_2865);
or U7809 (N_7809,In_39,In_453);
nor U7810 (N_7810,In_499,In_727);
and U7811 (N_7811,In_1346,In_976);
nand U7812 (N_7812,In_847,In_1152);
xor U7813 (N_7813,In_178,In_2017);
and U7814 (N_7814,In_1108,In_1479);
or U7815 (N_7815,In_2691,In_2406);
nor U7816 (N_7816,In_1266,In_1649);
or U7817 (N_7817,In_1681,In_193);
or U7818 (N_7818,In_196,In_518);
and U7819 (N_7819,In_321,In_2062);
xnor U7820 (N_7820,In_2489,In_1455);
nor U7821 (N_7821,In_2331,In_2799);
xor U7822 (N_7822,In_2160,In_1032);
nor U7823 (N_7823,In_2144,In_86);
nand U7824 (N_7824,In_1198,In_236);
nor U7825 (N_7825,In_1969,In_938);
nand U7826 (N_7826,In_226,In_2978);
and U7827 (N_7827,In_2619,In_571);
xor U7828 (N_7828,In_2407,In_2890);
nand U7829 (N_7829,In_66,In_2298);
xnor U7830 (N_7830,In_2003,In_1861);
nand U7831 (N_7831,In_1657,In_215);
nor U7832 (N_7832,In_242,In_411);
xor U7833 (N_7833,In_2259,In_581);
xor U7834 (N_7834,In_896,In_546);
nor U7835 (N_7835,In_2196,In_2039);
and U7836 (N_7836,In_436,In_1277);
xor U7837 (N_7837,In_1543,In_780);
or U7838 (N_7838,In_2362,In_942);
or U7839 (N_7839,In_2452,In_1922);
or U7840 (N_7840,In_2158,In_1756);
and U7841 (N_7841,In_1214,In_1157);
or U7842 (N_7842,In_2852,In_2941);
xor U7843 (N_7843,In_1057,In_2348);
and U7844 (N_7844,In_306,In_1378);
nor U7845 (N_7845,In_2593,In_2279);
nor U7846 (N_7846,In_1998,In_1554);
nand U7847 (N_7847,In_1005,In_1998);
xor U7848 (N_7848,In_722,In_970);
nand U7849 (N_7849,In_373,In_1868);
nor U7850 (N_7850,In_1343,In_210);
nor U7851 (N_7851,In_2215,In_2220);
xor U7852 (N_7852,In_1447,In_2432);
nor U7853 (N_7853,In_651,In_385);
or U7854 (N_7854,In_1021,In_2554);
nor U7855 (N_7855,In_2662,In_2879);
nand U7856 (N_7856,In_77,In_1140);
nor U7857 (N_7857,In_2516,In_1950);
xnor U7858 (N_7858,In_1819,In_2215);
and U7859 (N_7859,In_785,In_1299);
and U7860 (N_7860,In_2523,In_1261);
and U7861 (N_7861,In_1428,In_641);
nand U7862 (N_7862,In_2879,In_2870);
xor U7863 (N_7863,In_1690,In_2853);
xnor U7864 (N_7864,In_2284,In_1659);
or U7865 (N_7865,In_1141,In_1057);
nand U7866 (N_7866,In_1959,In_1351);
and U7867 (N_7867,In_421,In_1098);
and U7868 (N_7868,In_350,In_2221);
xor U7869 (N_7869,In_2999,In_1078);
nand U7870 (N_7870,In_735,In_2621);
nand U7871 (N_7871,In_456,In_1250);
nor U7872 (N_7872,In_2392,In_1683);
nor U7873 (N_7873,In_836,In_1128);
nand U7874 (N_7874,In_2688,In_2882);
nor U7875 (N_7875,In_725,In_213);
nand U7876 (N_7876,In_399,In_2623);
nand U7877 (N_7877,In_2969,In_1541);
or U7878 (N_7878,In_1408,In_765);
or U7879 (N_7879,In_187,In_2094);
nor U7880 (N_7880,In_785,In_2887);
xnor U7881 (N_7881,In_2311,In_1785);
and U7882 (N_7882,In_665,In_2089);
nand U7883 (N_7883,In_1339,In_2954);
nand U7884 (N_7884,In_1333,In_1517);
and U7885 (N_7885,In_1404,In_2236);
nand U7886 (N_7886,In_608,In_777);
nand U7887 (N_7887,In_23,In_519);
or U7888 (N_7888,In_2645,In_1256);
and U7889 (N_7889,In_291,In_1218);
nor U7890 (N_7890,In_2441,In_2321);
and U7891 (N_7891,In_724,In_1678);
or U7892 (N_7892,In_1463,In_2435);
and U7893 (N_7893,In_788,In_481);
xor U7894 (N_7894,In_2555,In_666);
and U7895 (N_7895,In_2404,In_486);
nor U7896 (N_7896,In_2974,In_542);
nand U7897 (N_7897,In_1077,In_2088);
or U7898 (N_7898,In_2949,In_2099);
and U7899 (N_7899,In_2824,In_1342);
and U7900 (N_7900,In_2106,In_621);
and U7901 (N_7901,In_2403,In_88);
nor U7902 (N_7902,In_244,In_1531);
or U7903 (N_7903,In_214,In_345);
and U7904 (N_7904,In_2424,In_1122);
nor U7905 (N_7905,In_191,In_2114);
xnor U7906 (N_7906,In_2952,In_2246);
xor U7907 (N_7907,In_2425,In_2944);
nand U7908 (N_7908,In_2621,In_861);
xor U7909 (N_7909,In_2203,In_1678);
or U7910 (N_7910,In_1255,In_1482);
xnor U7911 (N_7911,In_2353,In_2235);
nor U7912 (N_7912,In_1557,In_1366);
xor U7913 (N_7913,In_634,In_2027);
nand U7914 (N_7914,In_2898,In_289);
nor U7915 (N_7915,In_655,In_2722);
or U7916 (N_7916,In_766,In_952);
or U7917 (N_7917,In_79,In_1558);
nand U7918 (N_7918,In_2209,In_2991);
nor U7919 (N_7919,In_1958,In_126);
nand U7920 (N_7920,In_2320,In_2713);
xnor U7921 (N_7921,In_1295,In_1119);
xor U7922 (N_7922,In_2654,In_2399);
or U7923 (N_7923,In_1242,In_1224);
or U7924 (N_7924,In_2910,In_1314);
or U7925 (N_7925,In_2161,In_1430);
xor U7926 (N_7926,In_2916,In_2814);
and U7927 (N_7927,In_1159,In_2108);
or U7928 (N_7928,In_2800,In_2073);
and U7929 (N_7929,In_2184,In_1343);
nor U7930 (N_7930,In_2036,In_1283);
nand U7931 (N_7931,In_29,In_886);
nand U7932 (N_7932,In_195,In_229);
and U7933 (N_7933,In_1428,In_1558);
xnor U7934 (N_7934,In_1853,In_2029);
xor U7935 (N_7935,In_1901,In_1479);
or U7936 (N_7936,In_1235,In_1222);
xor U7937 (N_7937,In_1810,In_21);
nor U7938 (N_7938,In_31,In_2317);
nand U7939 (N_7939,In_1610,In_844);
or U7940 (N_7940,In_1850,In_523);
nor U7941 (N_7941,In_1748,In_14);
xor U7942 (N_7942,In_1495,In_910);
xnor U7943 (N_7943,In_766,In_181);
and U7944 (N_7944,In_362,In_1751);
nand U7945 (N_7945,In_1082,In_1403);
nand U7946 (N_7946,In_1321,In_2012);
and U7947 (N_7947,In_2101,In_2577);
and U7948 (N_7948,In_2568,In_2896);
xor U7949 (N_7949,In_1168,In_1279);
nand U7950 (N_7950,In_2501,In_1366);
nor U7951 (N_7951,In_431,In_1116);
nor U7952 (N_7952,In_1037,In_2393);
nor U7953 (N_7953,In_898,In_55);
or U7954 (N_7954,In_2774,In_532);
and U7955 (N_7955,In_854,In_1988);
and U7956 (N_7956,In_296,In_1366);
or U7957 (N_7957,In_863,In_2122);
nand U7958 (N_7958,In_2776,In_1924);
and U7959 (N_7959,In_1999,In_202);
xor U7960 (N_7960,In_1595,In_565);
and U7961 (N_7961,In_697,In_626);
and U7962 (N_7962,In_809,In_1610);
xnor U7963 (N_7963,In_1933,In_924);
nor U7964 (N_7964,In_2469,In_1930);
nand U7965 (N_7965,In_347,In_466);
nor U7966 (N_7966,In_2713,In_136);
nand U7967 (N_7967,In_197,In_667);
nand U7968 (N_7968,In_874,In_2527);
xnor U7969 (N_7969,In_666,In_1192);
or U7970 (N_7970,In_9,In_1578);
and U7971 (N_7971,In_1031,In_1097);
or U7972 (N_7972,In_1080,In_960);
and U7973 (N_7973,In_2433,In_1642);
xnor U7974 (N_7974,In_934,In_2457);
nand U7975 (N_7975,In_1243,In_2313);
and U7976 (N_7976,In_2313,In_520);
nor U7977 (N_7977,In_816,In_363);
xnor U7978 (N_7978,In_2241,In_772);
nand U7979 (N_7979,In_2974,In_1868);
or U7980 (N_7980,In_487,In_241);
and U7981 (N_7981,In_2282,In_2540);
nor U7982 (N_7982,In_2376,In_1338);
and U7983 (N_7983,In_318,In_259);
xnor U7984 (N_7984,In_2463,In_991);
or U7985 (N_7985,In_1264,In_1185);
and U7986 (N_7986,In_1048,In_1312);
nor U7987 (N_7987,In_1950,In_1461);
nor U7988 (N_7988,In_1695,In_572);
or U7989 (N_7989,In_598,In_1769);
or U7990 (N_7990,In_1201,In_2692);
nor U7991 (N_7991,In_1189,In_2419);
xor U7992 (N_7992,In_1017,In_2040);
or U7993 (N_7993,In_375,In_1343);
xor U7994 (N_7994,In_53,In_1368);
nand U7995 (N_7995,In_1660,In_305);
or U7996 (N_7996,In_2886,In_414);
nor U7997 (N_7997,In_2133,In_2234);
or U7998 (N_7998,In_1689,In_1744);
and U7999 (N_7999,In_1826,In_346);
or U8000 (N_8000,In_545,In_484);
nand U8001 (N_8001,In_1549,In_982);
nor U8002 (N_8002,In_2908,In_1181);
xnor U8003 (N_8003,In_14,In_860);
and U8004 (N_8004,In_2601,In_2027);
nor U8005 (N_8005,In_1928,In_1184);
and U8006 (N_8006,In_1177,In_1534);
nand U8007 (N_8007,In_14,In_2728);
xor U8008 (N_8008,In_259,In_2619);
nand U8009 (N_8009,In_991,In_2854);
or U8010 (N_8010,In_538,In_1414);
and U8011 (N_8011,In_1856,In_800);
and U8012 (N_8012,In_2685,In_805);
or U8013 (N_8013,In_1443,In_2768);
nor U8014 (N_8014,In_2704,In_793);
nand U8015 (N_8015,In_2289,In_2811);
and U8016 (N_8016,In_2182,In_441);
nor U8017 (N_8017,In_1794,In_778);
and U8018 (N_8018,In_2079,In_2447);
and U8019 (N_8019,In_1494,In_2513);
nand U8020 (N_8020,In_2845,In_385);
nor U8021 (N_8021,In_2278,In_2354);
and U8022 (N_8022,In_2269,In_2010);
and U8023 (N_8023,In_1021,In_2121);
nor U8024 (N_8024,In_1949,In_1534);
and U8025 (N_8025,In_2518,In_2530);
nand U8026 (N_8026,In_604,In_2153);
and U8027 (N_8027,In_1654,In_2474);
or U8028 (N_8028,In_2670,In_1088);
nor U8029 (N_8029,In_2721,In_611);
and U8030 (N_8030,In_2970,In_869);
xnor U8031 (N_8031,In_2389,In_1047);
nor U8032 (N_8032,In_2151,In_2930);
or U8033 (N_8033,In_700,In_942);
nand U8034 (N_8034,In_60,In_1486);
or U8035 (N_8035,In_2865,In_2280);
nand U8036 (N_8036,In_600,In_975);
or U8037 (N_8037,In_643,In_1466);
nor U8038 (N_8038,In_1027,In_1686);
nand U8039 (N_8039,In_2293,In_385);
or U8040 (N_8040,In_1603,In_1491);
and U8041 (N_8041,In_1775,In_669);
or U8042 (N_8042,In_748,In_466);
nor U8043 (N_8043,In_641,In_392);
and U8044 (N_8044,In_1588,In_1833);
nand U8045 (N_8045,In_1262,In_1729);
xnor U8046 (N_8046,In_2727,In_959);
nand U8047 (N_8047,In_1402,In_938);
and U8048 (N_8048,In_1623,In_344);
and U8049 (N_8049,In_441,In_446);
and U8050 (N_8050,In_1621,In_2722);
or U8051 (N_8051,In_1042,In_1691);
xor U8052 (N_8052,In_11,In_1684);
and U8053 (N_8053,In_306,In_2126);
xnor U8054 (N_8054,In_76,In_2480);
nor U8055 (N_8055,In_604,In_984);
and U8056 (N_8056,In_2829,In_1448);
or U8057 (N_8057,In_2270,In_1225);
and U8058 (N_8058,In_670,In_554);
or U8059 (N_8059,In_932,In_1048);
nor U8060 (N_8060,In_507,In_313);
nor U8061 (N_8061,In_319,In_208);
or U8062 (N_8062,In_1795,In_1133);
nor U8063 (N_8063,In_66,In_1172);
or U8064 (N_8064,In_1296,In_1244);
nand U8065 (N_8065,In_1559,In_118);
and U8066 (N_8066,In_1070,In_1016);
xor U8067 (N_8067,In_1056,In_2989);
nand U8068 (N_8068,In_2602,In_1680);
xor U8069 (N_8069,In_2810,In_1298);
nor U8070 (N_8070,In_1693,In_1551);
and U8071 (N_8071,In_397,In_709);
nand U8072 (N_8072,In_237,In_2782);
nor U8073 (N_8073,In_1087,In_2535);
or U8074 (N_8074,In_1861,In_1675);
and U8075 (N_8075,In_836,In_1733);
or U8076 (N_8076,In_1362,In_1559);
or U8077 (N_8077,In_1559,In_2560);
or U8078 (N_8078,In_1901,In_2810);
and U8079 (N_8079,In_2527,In_1819);
nor U8080 (N_8080,In_1064,In_1228);
nand U8081 (N_8081,In_1016,In_2507);
nand U8082 (N_8082,In_85,In_112);
and U8083 (N_8083,In_1326,In_1542);
xor U8084 (N_8084,In_1687,In_837);
nand U8085 (N_8085,In_1642,In_1833);
and U8086 (N_8086,In_1436,In_411);
or U8087 (N_8087,In_2927,In_2424);
nor U8088 (N_8088,In_1020,In_972);
nor U8089 (N_8089,In_1378,In_268);
nor U8090 (N_8090,In_1064,In_2900);
nand U8091 (N_8091,In_2625,In_2721);
xor U8092 (N_8092,In_1566,In_1442);
and U8093 (N_8093,In_2207,In_266);
or U8094 (N_8094,In_549,In_6);
nor U8095 (N_8095,In_2523,In_2402);
nor U8096 (N_8096,In_507,In_752);
xor U8097 (N_8097,In_1371,In_785);
or U8098 (N_8098,In_1952,In_2509);
and U8099 (N_8099,In_530,In_2168);
nand U8100 (N_8100,In_730,In_1646);
nand U8101 (N_8101,In_1082,In_2518);
and U8102 (N_8102,In_2159,In_1601);
or U8103 (N_8103,In_2097,In_2013);
xor U8104 (N_8104,In_128,In_1321);
and U8105 (N_8105,In_1263,In_2133);
or U8106 (N_8106,In_2500,In_2542);
xnor U8107 (N_8107,In_1853,In_967);
nand U8108 (N_8108,In_2934,In_2614);
xnor U8109 (N_8109,In_998,In_1740);
nor U8110 (N_8110,In_1854,In_1964);
xor U8111 (N_8111,In_792,In_1303);
and U8112 (N_8112,In_40,In_2714);
nor U8113 (N_8113,In_2964,In_935);
nor U8114 (N_8114,In_2043,In_405);
and U8115 (N_8115,In_1168,In_443);
nand U8116 (N_8116,In_1714,In_2362);
and U8117 (N_8117,In_1348,In_2946);
or U8118 (N_8118,In_2997,In_382);
or U8119 (N_8119,In_379,In_1898);
nor U8120 (N_8120,In_1238,In_800);
nand U8121 (N_8121,In_2886,In_2685);
and U8122 (N_8122,In_2094,In_2851);
nand U8123 (N_8123,In_933,In_1841);
and U8124 (N_8124,In_2222,In_2076);
and U8125 (N_8125,In_2320,In_2189);
or U8126 (N_8126,In_1589,In_2985);
nand U8127 (N_8127,In_184,In_1490);
or U8128 (N_8128,In_1601,In_2688);
or U8129 (N_8129,In_2787,In_88);
and U8130 (N_8130,In_1719,In_1024);
nand U8131 (N_8131,In_1139,In_1337);
and U8132 (N_8132,In_2250,In_97);
and U8133 (N_8133,In_967,In_2506);
or U8134 (N_8134,In_2853,In_1529);
or U8135 (N_8135,In_1445,In_933);
nor U8136 (N_8136,In_2238,In_1206);
xnor U8137 (N_8137,In_1532,In_1378);
nand U8138 (N_8138,In_804,In_162);
nand U8139 (N_8139,In_2042,In_1525);
or U8140 (N_8140,In_2412,In_2600);
xor U8141 (N_8141,In_1664,In_2574);
or U8142 (N_8142,In_1887,In_2306);
xor U8143 (N_8143,In_739,In_1912);
xnor U8144 (N_8144,In_2907,In_2168);
nor U8145 (N_8145,In_2129,In_1991);
xnor U8146 (N_8146,In_1339,In_476);
nor U8147 (N_8147,In_1017,In_367);
nand U8148 (N_8148,In_941,In_1746);
xnor U8149 (N_8149,In_2643,In_2880);
nand U8150 (N_8150,In_1242,In_2635);
and U8151 (N_8151,In_312,In_629);
nand U8152 (N_8152,In_1046,In_1270);
nand U8153 (N_8153,In_722,In_1020);
or U8154 (N_8154,In_1260,In_459);
nor U8155 (N_8155,In_1826,In_530);
xor U8156 (N_8156,In_1133,In_242);
nor U8157 (N_8157,In_2553,In_2356);
or U8158 (N_8158,In_2096,In_1951);
xnor U8159 (N_8159,In_1431,In_2390);
and U8160 (N_8160,In_2533,In_1310);
or U8161 (N_8161,In_2257,In_1742);
and U8162 (N_8162,In_541,In_1200);
xnor U8163 (N_8163,In_1186,In_1741);
xnor U8164 (N_8164,In_2139,In_1417);
xor U8165 (N_8165,In_1079,In_519);
nand U8166 (N_8166,In_1194,In_87);
and U8167 (N_8167,In_1871,In_2733);
nor U8168 (N_8168,In_20,In_160);
and U8169 (N_8169,In_809,In_1782);
or U8170 (N_8170,In_62,In_1344);
xor U8171 (N_8171,In_1081,In_638);
or U8172 (N_8172,In_262,In_1637);
xnor U8173 (N_8173,In_1046,In_2143);
xor U8174 (N_8174,In_171,In_895);
or U8175 (N_8175,In_2992,In_1283);
or U8176 (N_8176,In_990,In_825);
nand U8177 (N_8177,In_426,In_2636);
and U8178 (N_8178,In_854,In_1029);
and U8179 (N_8179,In_1279,In_2869);
nand U8180 (N_8180,In_459,In_744);
and U8181 (N_8181,In_1673,In_851);
nand U8182 (N_8182,In_1925,In_971);
nor U8183 (N_8183,In_2553,In_2028);
and U8184 (N_8184,In_773,In_2314);
nor U8185 (N_8185,In_2024,In_184);
or U8186 (N_8186,In_1141,In_1117);
and U8187 (N_8187,In_894,In_594);
and U8188 (N_8188,In_2474,In_2576);
or U8189 (N_8189,In_730,In_2346);
nor U8190 (N_8190,In_277,In_468);
or U8191 (N_8191,In_23,In_123);
nor U8192 (N_8192,In_1456,In_74);
and U8193 (N_8193,In_657,In_2392);
and U8194 (N_8194,In_2187,In_278);
nand U8195 (N_8195,In_2189,In_978);
nand U8196 (N_8196,In_1400,In_2099);
nor U8197 (N_8197,In_907,In_1473);
xor U8198 (N_8198,In_1394,In_1365);
nand U8199 (N_8199,In_1636,In_2496);
nor U8200 (N_8200,In_922,In_1573);
nand U8201 (N_8201,In_1236,In_367);
and U8202 (N_8202,In_2796,In_2665);
nand U8203 (N_8203,In_1364,In_686);
xor U8204 (N_8204,In_344,In_1205);
nor U8205 (N_8205,In_488,In_2668);
or U8206 (N_8206,In_2886,In_801);
nor U8207 (N_8207,In_1619,In_2755);
or U8208 (N_8208,In_1846,In_1109);
and U8209 (N_8209,In_2020,In_1180);
nor U8210 (N_8210,In_1928,In_1308);
and U8211 (N_8211,In_1390,In_2436);
nor U8212 (N_8212,In_1376,In_1012);
xor U8213 (N_8213,In_434,In_1022);
xor U8214 (N_8214,In_1838,In_2497);
nor U8215 (N_8215,In_1879,In_2306);
xnor U8216 (N_8216,In_1387,In_2796);
xor U8217 (N_8217,In_1450,In_256);
or U8218 (N_8218,In_2744,In_140);
nor U8219 (N_8219,In_2195,In_2667);
and U8220 (N_8220,In_2991,In_2750);
and U8221 (N_8221,In_2193,In_155);
nor U8222 (N_8222,In_2035,In_2973);
and U8223 (N_8223,In_1338,In_742);
or U8224 (N_8224,In_64,In_2016);
and U8225 (N_8225,In_2697,In_656);
nor U8226 (N_8226,In_2589,In_293);
nor U8227 (N_8227,In_859,In_581);
nand U8228 (N_8228,In_1509,In_2856);
nand U8229 (N_8229,In_1523,In_1688);
or U8230 (N_8230,In_1059,In_986);
nand U8231 (N_8231,In_1225,In_1151);
nand U8232 (N_8232,In_1552,In_791);
xnor U8233 (N_8233,In_435,In_1646);
or U8234 (N_8234,In_2050,In_2786);
nor U8235 (N_8235,In_2414,In_771);
nor U8236 (N_8236,In_171,In_1548);
nor U8237 (N_8237,In_129,In_1876);
nor U8238 (N_8238,In_94,In_1403);
and U8239 (N_8239,In_2834,In_752);
nand U8240 (N_8240,In_1390,In_2548);
xor U8241 (N_8241,In_1371,In_747);
and U8242 (N_8242,In_1144,In_30);
xor U8243 (N_8243,In_171,In_495);
or U8244 (N_8244,In_1315,In_1104);
and U8245 (N_8245,In_2188,In_313);
nand U8246 (N_8246,In_294,In_2895);
xnor U8247 (N_8247,In_1404,In_2562);
xnor U8248 (N_8248,In_93,In_120);
or U8249 (N_8249,In_560,In_887);
nor U8250 (N_8250,In_1851,In_1746);
nand U8251 (N_8251,In_2309,In_2481);
xor U8252 (N_8252,In_2449,In_2791);
and U8253 (N_8253,In_234,In_779);
and U8254 (N_8254,In_2263,In_2718);
or U8255 (N_8255,In_2776,In_2943);
nand U8256 (N_8256,In_2898,In_2245);
nor U8257 (N_8257,In_2794,In_2020);
nand U8258 (N_8258,In_776,In_1188);
xor U8259 (N_8259,In_852,In_2395);
and U8260 (N_8260,In_1485,In_2216);
nand U8261 (N_8261,In_840,In_1431);
xor U8262 (N_8262,In_562,In_189);
xnor U8263 (N_8263,In_277,In_2692);
or U8264 (N_8264,In_2816,In_1858);
nor U8265 (N_8265,In_2911,In_171);
or U8266 (N_8266,In_604,In_1407);
nor U8267 (N_8267,In_730,In_2807);
xnor U8268 (N_8268,In_1853,In_2392);
or U8269 (N_8269,In_507,In_2998);
nand U8270 (N_8270,In_1763,In_1790);
or U8271 (N_8271,In_1534,In_650);
or U8272 (N_8272,In_1397,In_2569);
nand U8273 (N_8273,In_1189,In_504);
and U8274 (N_8274,In_1982,In_2893);
xnor U8275 (N_8275,In_1932,In_1280);
and U8276 (N_8276,In_1034,In_1814);
or U8277 (N_8277,In_2460,In_1719);
xnor U8278 (N_8278,In_1187,In_2235);
nor U8279 (N_8279,In_238,In_1369);
and U8280 (N_8280,In_2882,In_1233);
xnor U8281 (N_8281,In_1931,In_499);
or U8282 (N_8282,In_2919,In_1956);
xnor U8283 (N_8283,In_887,In_67);
nor U8284 (N_8284,In_242,In_383);
nand U8285 (N_8285,In_2436,In_845);
or U8286 (N_8286,In_1162,In_122);
nand U8287 (N_8287,In_714,In_1419);
or U8288 (N_8288,In_1396,In_2167);
or U8289 (N_8289,In_1442,In_2368);
and U8290 (N_8290,In_2391,In_1393);
xor U8291 (N_8291,In_2219,In_138);
or U8292 (N_8292,In_568,In_2078);
or U8293 (N_8293,In_151,In_780);
xnor U8294 (N_8294,In_985,In_801);
or U8295 (N_8295,In_493,In_1002);
or U8296 (N_8296,In_1410,In_209);
or U8297 (N_8297,In_2117,In_1110);
nor U8298 (N_8298,In_600,In_2928);
nand U8299 (N_8299,In_2763,In_558);
or U8300 (N_8300,In_1961,In_550);
xnor U8301 (N_8301,In_626,In_729);
xnor U8302 (N_8302,In_2574,In_69);
or U8303 (N_8303,In_1613,In_2996);
nand U8304 (N_8304,In_300,In_2447);
nor U8305 (N_8305,In_136,In_9);
nand U8306 (N_8306,In_182,In_9);
and U8307 (N_8307,In_1414,In_302);
and U8308 (N_8308,In_2991,In_780);
xor U8309 (N_8309,In_2370,In_562);
nor U8310 (N_8310,In_2188,In_1292);
nand U8311 (N_8311,In_1969,In_408);
and U8312 (N_8312,In_1042,In_984);
xor U8313 (N_8313,In_1265,In_2523);
nand U8314 (N_8314,In_2141,In_332);
or U8315 (N_8315,In_2310,In_731);
nor U8316 (N_8316,In_216,In_1703);
xnor U8317 (N_8317,In_2501,In_2154);
nand U8318 (N_8318,In_2315,In_2184);
or U8319 (N_8319,In_892,In_79);
or U8320 (N_8320,In_692,In_930);
xnor U8321 (N_8321,In_2224,In_923);
nor U8322 (N_8322,In_825,In_2255);
or U8323 (N_8323,In_2383,In_1115);
nand U8324 (N_8324,In_751,In_1424);
nand U8325 (N_8325,In_1669,In_2206);
or U8326 (N_8326,In_196,In_1688);
nand U8327 (N_8327,In_1526,In_138);
or U8328 (N_8328,In_1161,In_447);
xnor U8329 (N_8329,In_889,In_1244);
nor U8330 (N_8330,In_2335,In_2153);
nand U8331 (N_8331,In_693,In_1525);
xnor U8332 (N_8332,In_710,In_2665);
and U8333 (N_8333,In_1942,In_154);
and U8334 (N_8334,In_2123,In_1838);
nor U8335 (N_8335,In_1644,In_1017);
and U8336 (N_8336,In_1837,In_253);
or U8337 (N_8337,In_813,In_1543);
or U8338 (N_8338,In_2916,In_884);
xor U8339 (N_8339,In_2763,In_2705);
xor U8340 (N_8340,In_849,In_1511);
and U8341 (N_8341,In_2702,In_937);
and U8342 (N_8342,In_1841,In_1177);
and U8343 (N_8343,In_996,In_196);
nor U8344 (N_8344,In_996,In_448);
nor U8345 (N_8345,In_2690,In_1826);
xnor U8346 (N_8346,In_1657,In_2502);
xnor U8347 (N_8347,In_1305,In_1236);
nand U8348 (N_8348,In_2085,In_2505);
xor U8349 (N_8349,In_1568,In_1449);
or U8350 (N_8350,In_462,In_2577);
nand U8351 (N_8351,In_16,In_765);
nand U8352 (N_8352,In_1304,In_2670);
xnor U8353 (N_8353,In_1294,In_2282);
xnor U8354 (N_8354,In_2474,In_112);
xor U8355 (N_8355,In_1283,In_1437);
or U8356 (N_8356,In_409,In_440);
or U8357 (N_8357,In_1735,In_995);
xnor U8358 (N_8358,In_1672,In_921);
nand U8359 (N_8359,In_2877,In_1958);
nand U8360 (N_8360,In_251,In_2971);
xnor U8361 (N_8361,In_1867,In_1371);
nand U8362 (N_8362,In_1413,In_1147);
or U8363 (N_8363,In_1899,In_393);
nand U8364 (N_8364,In_2358,In_2520);
or U8365 (N_8365,In_1838,In_621);
xor U8366 (N_8366,In_771,In_895);
nand U8367 (N_8367,In_1141,In_315);
nand U8368 (N_8368,In_2399,In_2505);
xnor U8369 (N_8369,In_334,In_2829);
and U8370 (N_8370,In_1631,In_955);
and U8371 (N_8371,In_1565,In_188);
xnor U8372 (N_8372,In_1169,In_1122);
nand U8373 (N_8373,In_156,In_1398);
or U8374 (N_8374,In_1001,In_1572);
and U8375 (N_8375,In_961,In_523);
nand U8376 (N_8376,In_1763,In_266);
xor U8377 (N_8377,In_2799,In_735);
xor U8378 (N_8378,In_305,In_1844);
nand U8379 (N_8379,In_1882,In_2395);
nand U8380 (N_8380,In_1976,In_1933);
and U8381 (N_8381,In_267,In_954);
xor U8382 (N_8382,In_902,In_1295);
nand U8383 (N_8383,In_2113,In_2421);
xor U8384 (N_8384,In_815,In_1187);
xor U8385 (N_8385,In_2697,In_1820);
xnor U8386 (N_8386,In_1176,In_2075);
xnor U8387 (N_8387,In_2279,In_878);
nor U8388 (N_8388,In_1324,In_983);
xnor U8389 (N_8389,In_39,In_1788);
nor U8390 (N_8390,In_35,In_963);
or U8391 (N_8391,In_114,In_659);
nor U8392 (N_8392,In_1647,In_2459);
or U8393 (N_8393,In_2645,In_2526);
nor U8394 (N_8394,In_796,In_174);
xnor U8395 (N_8395,In_1466,In_537);
or U8396 (N_8396,In_1531,In_1111);
xnor U8397 (N_8397,In_2846,In_569);
nor U8398 (N_8398,In_2124,In_449);
or U8399 (N_8399,In_2438,In_1558);
and U8400 (N_8400,In_585,In_1805);
xnor U8401 (N_8401,In_1708,In_2216);
xor U8402 (N_8402,In_1627,In_376);
nand U8403 (N_8403,In_234,In_2989);
nand U8404 (N_8404,In_2378,In_565);
and U8405 (N_8405,In_420,In_2614);
or U8406 (N_8406,In_2583,In_1314);
or U8407 (N_8407,In_2633,In_352);
xnor U8408 (N_8408,In_4,In_526);
xnor U8409 (N_8409,In_1424,In_1483);
nand U8410 (N_8410,In_1912,In_1621);
nand U8411 (N_8411,In_2334,In_588);
or U8412 (N_8412,In_2345,In_255);
xnor U8413 (N_8413,In_393,In_351);
xnor U8414 (N_8414,In_1281,In_82);
and U8415 (N_8415,In_2445,In_65);
nor U8416 (N_8416,In_1570,In_1639);
xnor U8417 (N_8417,In_52,In_519);
nand U8418 (N_8418,In_749,In_1502);
and U8419 (N_8419,In_2182,In_1303);
nand U8420 (N_8420,In_669,In_674);
nor U8421 (N_8421,In_2530,In_1245);
and U8422 (N_8422,In_1675,In_2748);
nor U8423 (N_8423,In_2012,In_643);
xnor U8424 (N_8424,In_2170,In_815);
and U8425 (N_8425,In_764,In_1180);
nand U8426 (N_8426,In_2699,In_473);
xor U8427 (N_8427,In_1144,In_1842);
xor U8428 (N_8428,In_2860,In_1068);
nand U8429 (N_8429,In_2880,In_2218);
nand U8430 (N_8430,In_2433,In_2324);
or U8431 (N_8431,In_2463,In_1263);
nand U8432 (N_8432,In_2734,In_1263);
xor U8433 (N_8433,In_885,In_1797);
or U8434 (N_8434,In_1750,In_1211);
or U8435 (N_8435,In_1059,In_2540);
nor U8436 (N_8436,In_2975,In_2025);
nor U8437 (N_8437,In_669,In_1459);
and U8438 (N_8438,In_559,In_959);
or U8439 (N_8439,In_1260,In_1122);
nor U8440 (N_8440,In_2320,In_2138);
and U8441 (N_8441,In_1224,In_100);
and U8442 (N_8442,In_660,In_1454);
xor U8443 (N_8443,In_1872,In_2577);
xor U8444 (N_8444,In_2925,In_300);
nand U8445 (N_8445,In_1608,In_2144);
or U8446 (N_8446,In_2502,In_1125);
nor U8447 (N_8447,In_320,In_1623);
and U8448 (N_8448,In_1064,In_1112);
or U8449 (N_8449,In_1569,In_2117);
or U8450 (N_8450,In_1179,In_2284);
and U8451 (N_8451,In_925,In_2266);
and U8452 (N_8452,In_2020,In_1532);
xor U8453 (N_8453,In_747,In_2149);
and U8454 (N_8454,In_2147,In_2239);
and U8455 (N_8455,In_519,In_2755);
and U8456 (N_8456,In_2752,In_429);
xor U8457 (N_8457,In_1573,In_1698);
nor U8458 (N_8458,In_586,In_565);
or U8459 (N_8459,In_289,In_925);
and U8460 (N_8460,In_1552,In_1104);
nand U8461 (N_8461,In_873,In_717);
or U8462 (N_8462,In_893,In_240);
nor U8463 (N_8463,In_1149,In_1259);
xor U8464 (N_8464,In_1316,In_553);
nand U8465 (N_8465,In_2761,In_880);
xnor U8466 (N_8466,In_2254,In_1006);
and U8467 (N_8467,In_2098,In_520);
or U8468 (N_8468,In_295,In_1008);
and U8469 (N_8469,In_1304,In_647);
and U8470 (N_8470,In_517,In_1472);
nand U8471 (N_8471,In_1190,In_931);
xnor U8472 (N_8472,In_2399,In_2447);
nand U8473 (N_8473,In_173,In_254);
or U8474 (N_8474,In_2543,In_2945);
nor U8475 (N_8475,In_562,In_2299);
and U8476 (N_8476,In_2570,In_942);
xnor U8477 (N_8477,In_1611,In_1866);
nor U8478 (N_8478,In_1781,In_550);
and U8479 (N_8479,In_1481,In_1608);
nor U8480 (N_8480,In_2742,In_1620);
nor U8481 (N_8481,In_184,In_716);
and U8482 (N_8482,In_1241,In_1975);
nor U8483 (N_8483,In_1575,In_2496);
or U8484 (N_8484,In_1453,In_2300);
or U8485 (N_8485,In_728,In_2279);
nor U8486 (N_8486,In_1595,In_1886);
or U8487 (N_8487,In_1805,In_2230);
xor U8488 (N_8488,In_455,In_1300);
nand U8489 (N_8489,In_82,In_127);
xor U8490 (N_8490,In_314,In_1992);
or U8491 (N_8491,In_1869,In_1170);
nor U8492 (N_8492,In_2284,In_1793);
xor U8493 (N_8493,In_2479,In_2286);
xor U8494 (N_8494,In_693,In_1770);
nand U8495 (N_8495,In_2795,In_1261);
and U8496 (N_8496,In_719,In_2986);
nor U8497 (N_8497,In_640,In_2681);
or U8498 (N_8498,In_200,In_2413);
or U8499 (N_8499,In_1445,In_2929);
nand U8500 (N_8500,In_803,In_2998);
xor U8501 (N_8501,In_1897,In_247);
nor U8502 (N_8502,In_339,In_2953);
or U8503 (N_8503,In_1925,In_403);
nor U8504 (N_8504,In_30,In_2948);
and U8505 (N_8505,In_2104,In_2803);
xor U8506 (N_8506,In_793,In_1016);
nand U8507 (N_8507,In_2126,In_877);
xor U8508 (N_8508,In_518,In_1633);
nand U8509 (N_8509,In_588,In_2535);
and U8510 (N_8510,In_1919,In_2656);
and U8511 (N_8511,In_112,In_2762);
nand U8512 (N_8512,In_1698,In_1627);
nand U8513 (N_8513,In_632,In_1205);
nand U8514 (N_8514,In_1862,In_32);
or U8515 (N_8515,In_1449,In_247);
or U8516 (N_8516,In_1380,In_2442);
nand U8517 (N_8517,In_1920,In_2391);
and U8518 (N_8518,In_2605,In_2912);
nor U8519 (N_8519,In_2388,In_2474);
nor U8520 (N_8520,In_2285,In_1706);
nand U8521 (N_8521,In_1559,In_1652);
and U8522 (N_8522,In_2942,In_1367);
nand U8523 (N_8523,In_2999,In_802);
nor U8524 (N_8524,In_1998,In_1691);
or U8525 (N_8525,In_2357,In_1191);
xnor U8526 (N_8526,In_2052,In_2820);
or U8527 (N_8527,In_2599,In_2740);
and U8528 (N_8528,In_106,In_1748);
or U8529 (N_8529,In_2912,In_357);
xor U8530 (N_8530,In_1336,In_1563);
nand U8531 (N_8531,In_2787,In_2674);
and U8532 (N_8532,In_2536,In_978);
nor U8533 (N_8533,In_2090,In_2876);
nor U8534 (N_8534,In_2173,In_2881);
and U8535 (N_8535,In_530,In_2372);
and U8536 (N_8536,In_2606,In_1522);
xnor U8537 (N_8537,In_2657,In_2315);
nor U8538 (N_8538,In_2197,In_849);
or U8539 (N_8539,In_846,In_2296);
or U8540 (N_8540,In_887,In_136);
or U8541 (N_8541,In_1524,In_2340);
xor U8542 (N_8542,In_820,In_1630);
nor U8543 (N_8543,In_786,In_431);
or U8544 (N_8544,In_194,In_309);
or U8545 (N_8545,In_2906,In_408);
and U8546 (N_8546,In_822,In_831);
or U8547 (N_8547,In_1084,In_2405);
xnor U8548 (N_8548,In_1866,In_2629);
or U8549 (N_8549,In_1463,In_2600);
xnor U8550 (N_8550,In_912,In_1843);
and U8551 (N_8551,In_568,In_1933);
or U8552 (N_8552,In_2245,In_835);
nor U8553 (N_8553,In_2791,In_2917);
or U8554 (N_8554,In_2521,In_2895);
nand U8555 (N_8555,In_683,In_2816);
and U8556 (N_8556,In_281,In_157);
nor U8557 (N_8557,In_2850,In_1473);
or U8558 (N_8558,In_1444,In_1888);
nor U8559 (N_8559,In_1414,In_2576);
or U8560 (N_8560,In_2772,In_1705);
nor U8561 (N_8561,In_98,In_2951);
nor U8562 (N_8562,In_2245,In_2827);
nor U8563 (N_8563,In_2655,In_2775);
nor U8564 (N_8564,In_2833,In_2251);
or U8565 (N_8565,In_1554,In_2240);
and U8566 (N_8566,In_1540,In_2854);
and U8567 (N_8567,In_1377,In_2764);
xor U8568 (N_8568,In_45,In_1318);
or U8569 (N_8569,In_1548,In_2373);
nand U8570 (N_8570,In_738,In_2059);
or U8571 (N_8571,In_1131,In_2865);
xnor U8572 (N_8572,In_1587,In_2107);
xnor U8573 (N_8573,In_829,In_623);
nand U8574 (N_8574,In_676,In_421);
and U8575 (N_8575,In_29,In_2408);
and U8576 (N_8576,In_2154,In_840);
nand U8577 (N_8577,In_1947,In_2086);
xnor U8578 (N_8578,In_1928,In_446);
and U8579 (N_8579,In_1898,In_1143);
nand U8580 (N_8580,In_2396,In_197);
or U8581 (N_8581,In_2505,In_1141);
nand U8582 (N_8582,In_2578,In_982);
xnor U8583 (N_8583,In_708,In_1061);
xor U8584 (N_8584,In_153,In_1768);
xnor U8585 (N_8585,In_2900,In_950);
nor U8586 (N_8586,In_585,In_2749);
nand U8587 (N_8587,In_518,In_1324);
nand U8588 (N_8588,In_1740,In_651);
or U8589 (N_8589,In_9,In_2393);
and U8590 (N_8590,In_2264,In_1499);
or U8591 (N_8591,In_760,In_2025);
nor U8592 (N_8592,In_1027,In_675);
xnor U8593 (N_8593,In_2477,In_2064);
nor U8594 (N_8594,In_195,In_552);
and U8595 (N_8595,In_920,In_1954);
nand U8596 (N_8596,In_2108,In_972);
xor U8597 (N_8597,In_597,In_2415);
xnor U8598 (N_8598,In_2239,In_813);
or U8599 (N_8599,In_1534,In_972);
and U8600 (N_8600,In_605,In_1212);
nand U8601 (N_8601,In_738,In_2527);
and U8602 (N_8602,In_991,In_2195);
nor U8603 (N_8603,In_1269,In_1268);
and U8604 (N_8604,In_858,In_2644);
xnor U8605 (N_8605,In_26,In_239);
or U8606 (N_8606,In_793,In_853);
nor U8607 (N_8607,In_1916,In_1114);
and U8608 (N_8608,In_2285,In_2739);
and U8609 (N_8609,In_1069,In_2014);
xor U8610 (N_8610,In_373,In_2931);
and U8611 (N_8611,In_1270,In_1099);
and U8612 (N_8612,In_760,In_860);
nor U8613 (N_8613,In_2046,In_392);
xnor U8614 (N_8614,In_2450,In_2629);
xor U8615 (N_8615,In_0,In_574);
and U8616 (N_8616,In_1984,In_2858);
and U8617 (N_8617,In_1969,In_2362);
nand U8618 (N_8618,In_719,In_2280);
and U8619 (N_8619,In_1270,In_2152);
nor U8620 (N_8620,In_2326,In_2485);
or U8621 (N_8621,In_2526,In_1377);
nor U8622 (N_8622,In_184,In_706);
nor U8623 (N_8623,In_638,In_645);
xor U8624 (N_8624,In_4,In_2967);
or U8625 (N_8625,In_1003,In_879);
nand U8626 (N_8626,In_1853,In_354);
nor U8627 (N_8627,In_2596,In_1853);
nor U8628 (N_8628,In_2815,In_1169);
nand U8629 (N_8629,In_2766,In_2854);
xor U8630 (N_8630,In_1854,In_639);
and U8631 (N_8631,In_320,In_1535);
nor U8632 (N_8632,In_122,In_703);
and U8633 (N_8633,In_472,In_179);
xnor U8634 (N_8634,In_1319,In_133);
and U8635 (N_8635,In_1842,In_1482);
or U8636 (N_8636,In_455,In_408);
xnor U8637 (N_8637,In_1737,In_694);
and U8638 (N_8638,In_1188,In_966);
and U8639 (N_8639,In_389,In_1858);
xnor U8640 (N_8640,In_704,In_2080);
or U8641 (N_8641,In_2264,In_364);
nor U8642 (N_8642,In_2371,In_1736);
xor U8643 (N_8643,In_95,In_2972);
nand U8644 (N_8644,In_2784,In_1503);
or U8645 (N_8645,In_2441,In_2413);
xor U8646 (N_8646,In_426,In_1852);
or U8647 (N_8647,In_2508,In_1876);
xor U8648 (N_8648,In_2150,In_1174);
and U8649 (N_8649,In_1334,In_297);
nor U8650 (N_8650,In_1191,In_2348);
xnor U8651 (N_8651,In_9,In_2076);
xnor U8652 (N_8652,In_1286,In_651);
nand U8653 (N_8653,In_2035,In_49);
and U8654 (N_8654,In_651,In_2573);
and U8655 (N_8655,In_1190,In_94);
nor U8656 (N_8656,In_452,In_2773);
xnor U8657 (N_8657,In_1984,In_2184);
and U8658 (N_8658,In_2503,In_1627);
and U8659 (N_8659,In_68,In_2772);
and U8660 (N_8660,In_38,In_1365);
nand U8661 (N_8661,In_1715,In_1127);
and U8662 (N_8662,In_855,In_636);
and U8663 (N_8663,In_1439,In_966);
nor U8664 (N_8664,In_331,In_254);
or U8665 (N_8665,In_2365,In_2830);
or U8666 (N_8666,In_2840,In_697);
xor U8667 (N_8667,In_43,In_1658);
xor U8668 (N_8668,In_1041,In_1490);
nor U8669 (N_8669,In_1790,In_860);
nor U8670 (N_8670,In_2577,In_8);
and U8671 (N_8671,In_1776,In_1199);
or U8672 (N_8672,In_483,In_749);
nor U8673 (N_8673,In_372,In_446);
or U8674 (N_8674,In_544,In_133);
nor U8675 (N_8675,In_2099,In_185);
or U8676 (N_8676,In_358,In_1111);
nor U8677 (N_8677,In_1954,In_2355);
nor U8678 (N_8678,In_369,In_1734);
or U8679 (N_8679,In_2772,In_1100);
and U8680 (N_8680,In_2011,In_1096);
and U8681 (N_8681,In_99,In_1797);
xor U8682 (N_8682,In_2406,In_2227);
nand U8683 (N_8683,In_1615,In_925);
or U8684 (N_8684,In_437,In_1556);
xnor U8685 (N_8685,In_1044,In_1851);
nand U8686 (N_8686,In_1790,In_1445);
nand U8687 (N_8687,In_2783,In_2769);
xnor U8688 (N_8688,In_2240,In_2577);
nor U8689 (N_8689,In_70,In_1488);
or U8690 (N_8690,In_1411,In_1449);
and U8691 (N_8691,In_2674,In_257);
xnor U8692 (N_8692,In_1297,In_2653);
nor U8693 (N_8693,In_2957,In_1124);
nand U8694 (N_8694,In_2596,In_837);
or U8695 (N_8695,In_2722,In_2319);
or U8696 (N_8696,In_1696,In_1017);
nand U8697 (N_8697,In_1622,In_266);
nor U8698 (N_8698,In_1768,In_1288);
xor U8699 (N_8699,In_2095,In_2369);
nor U8700 (N_8700,In_978,In_846);
xnor U8701 (N_8701,In_1072,In_998);
nor U8702 (N_8702,In_2085,In_1676);
nand U8703 (N_8703,In_962,In_2781);
nor U8704 (N_8704,In_832,In_2283);
or U8705 (N_8705,In_1306,In_509);
or U8706 (N_8706,In_485,In_5);
nand U8707 (N_8707,In_1581,In_1397);
xnor U8708 (N_8708,In_2271,In_1479);
or U8709 (N_8709,In_271,In_785);
or U8710 (N_8710,In_1355,In_2966);
and U8711 (N_8711,In_2924,In_2069);
nand U8712 (N_8712,In_2061,In_2651);
or U8713 (N_8713,In_1207,In_2112);
nor U8714 (N_8714,In_851,In_699);
nor U8715 (N_8715,In_640,In_1613);
nand U8716 (N_8716,In_1990,In_545);
or U8717 (N_8717,In_304,In_2004);
nor U8718 (N_8718,In_2877,In_774);
nand U8719 (N_8719,In_2924,In_2109);
nand U8720 (N_8720,In_2645,In_836);
xor U8721 (N_8721,In_2903,In_10);
nand U8722 (N_8722,In_425,In_2108);
nor U8723 (N_8723,In_234,In_489);
xnor U8724 (N_8724,In_2910,In_797);
or U8725 (N_8725,In_2227,In_779);
and U8726 (N_8726,In_2375,In_357);
and U8727 (N_8727,In_927,In_2023);
xnor U8728 (N_8728,In_217,In_2000);
and U8729 (N_8729,In_637,In_970);
xor U8730 (N_8730,In_41,In_2704);
nand U8731 (N_8731,In_2377,In_2750);
nor U8732 (N_8732,In_199,In_2341);
nor U8733 (N_8733,In_521,In_1039);
nor U8734 (N_8734,In_993,In_1894);
xnor U8735 (N_8735,In_1271,In_260);
nand U8736 (N_8736,In_1718,In_2245);
nor U8737 (N_8737,In_1252,In_18);
nand U8738 (N_8738,In_1972,In_910);
nor U8739 (N_8739,In_2783,In_1741);
and U8740 (N_8740,In_2572,In_1982);
nor U8741 (N_8741,In_2094,In_1084);
and U8742 (N_8742,In_595,In_1153);
and U8743 (N_8743,In_2346,In_1549);
nand U8744 (N_8744,In_934,In_2609);
nand U8745 (N_8745,In_550,In_2561);
xnor U8746 (N_8746,In_834,In_1280);
or U8747 (N_8747,In_1423,In_1238);
xor U8748 (N_8748,In_760,In_665);
or U8749 (N_8749,In_2486,In_67);
nor U8750 (N_8750,In_1375,In_1126);
and U8751 (N_8751,In_475,In_2595);
xnor U8752 (N_8752,In_415,In_2974);
xor U8753 (N_8753,In_2272,In_2768);
nor U8754 (N_8754,In_2482,In_1059);
xnor U8755 (N_8755,In_2907,In_574);
xnor U8756 (N_8756,In_2660,In_2471);
nor U8757 (N_8757,In_956,In_781);
nor U8758 (N_8758,In_2584,In_2947);
and U8759 (N_8759,In_1554,In_1097);
xor U8760 (N_8760,In_1960,In_688);
and U8761 (N_8761,In_274,In_2627);
nand U8762 (N_8762,In_1783,In_2499);
nand U8763 (N_8763,In_622,In_1867);
nand U8764 (N_8764,In_785,In_1066);
and U8765 (N_8765,In_873,In_689);
and U8766 (N_8766,In_1702,In_1962);
nand U8767 (N_8767,In_2169,In_1580);
nand U8768 (N_8768,In_1973,In_821);
nand U8769 (N_8769,In_382,In_967);
and U8770 (N_8770,In_2950,In_284);
and U8771 (N_8771,In_1978,In_2518);
or U8772 (N_8772,In_1893,In_137);
nand U8773 (N_8773,In_2516,In_446);
and U8774 (N_8774,In_1244,In_216);
or U8775 (N_8775,In_1021,In_105);
and U8776 (N_8776,In_867,In_978);
and U8777 (N_8777,In_165,In_578);
xor U8778 (N_8778,In_817,In_357);
nand U8779 (N_8779,In_1321,In_1741);
and U8780 (N_8780,In_230,In_2955);
and U8781 (N_8781,In_262,In_289);
nor U8782 (N_8782,In_455,In_2844);
or U8783 (N_8783,In_2792,In_2856);
nor U8784 (N_8784,In_192,In_1085);
nand U8785 (N_8785,In_2771,In_2619);
nand U8786 (N_8786,In_1517,In_1814);
or U8787 (N_8787,In_2563,In_2442);
or U8788 (N_8788,In_1026,In_2717);
or U8789 (N_8789,In_2992,In_1714);
and U8790 (N_8790,In_837,In_1971);
xnor U8791 (N_8791,In_231,In_918);
xnor U8792 (N_8792,In_1249,In_2302);
and U8793 (N_8793,In_826,In_1673);
or U8794 (N_8794,In_1054,In_1913);
nand U8795 (N_8795,In_821,In_2538);
and U8796 (N_8796,In_1614,In_256);
xnor U8797 (N_8797,In_527,In_1367);
nor U8798 (N_8798,In_1625,In_341);
and U8799 (N_8799,In_1458,In_1879);
and U8800 (N_8800,In_397,In_2507);
nor U8801 (N_8801,In_1720,In_1368);
and U8802 (N_8802,In_2429,In_1897);
xor U8803 (N_8803,In_1604,In_2667);
nor U8804 (N_8804,In_2377,In_2602);
or U8805 (N_8805,In_1165,In_1866);
and U8806 (N_8806,In_1778,In_2038);
xnor U8807 (N_8807,In_162,In_2810);
xnor U8808 (N_8808,In_1052,In_1116);
and U8809 (N_8809,In_2406,In_2885);
nand U8810 (N_8810,In_1527,In_331);
or U8811 (N_8811,In_2,In_633);
nand U8812 (N_8812,In_1301,In_866);
xor U8813 (N_8813,In_2575,In_2036);
xnor U8814 (N_8814,In_55,In_1407);
nor U8815 (N_8815,In_2253,In_2954);
or U8816 (N_8816,In_579,In_524);
nor U8817 (N_8817,In_2538,In_1092);
nand U8818 (N_8818,In_2037,In_369);
nor U8819 (N_8819,In_1567,In_1117);
or U8820 (N_8820,In_1300,In_286);
and U8821 (N_8821,In_2257,In_1955);
xor U8822 (N_8822,In_2200,In_2165);
nand U8823 (N_8823,In_1242,In_1637);
and U8824 (N_8824,In_1393,In_1045);
nand U8825 (N_8825,In_2002,In_334);
or U8826 (N_8826,In_0,In_2952);
nand U8827 (N_8827,In_1775,In_2084);
and U8828 (N_8828,In_972,In_2791);
or U8829 (N_8829,In_1970,In_1093);
nor U8830 (N_8830,In_938,In_2578);
or U8831 (N_8831,In_1745,In_552);
and U8832 (N_8832,In_1385,In_2259);
or U8833 (N_8833,In_1010,In_2398);
and U8834 (N_8834,In_1410,In_2132);
xnor U8835 (N_8835,In_2337,In_2919);
or U8836 (N_8836,In_1217,In_1639);
nand U8837 (N_8837,In_2011,In_1813);
nand U8838 (N_8838,In_1522,In_868);
xor U8839 (N_8839,In_1817,In_1339);
nand U8840 (N_8840,In_265,In_413);
xor U8841 (N_8841,In_1209,In_1232);
and U8842 (N_8842,In_1845,In_1935);
xor U8843 (N_8843,In_775,In_2501);
xor U8844 (N_8844,In_593,In_2414);
and U8845 (N_8845,In_1467,In_444);
xnor U8846 (N_8846,In_421,In_1145);
nor U8847 (N_8847,In_1204,In_2794);
or U8848 (N_8848,In_2682,In_443);
nor U8849 (N_8849,In_1214,In_1337);
xnor U8850 (N_8850,In_1693,In_282);
and U8851 (N_8851,In_1755,In_2860);
xnor U8852 (N_8852,In_1807,In_1220);
and U8853 (N_8853,In_2628,In_508);
and U8854 (N_8854,In_386,In_2835);
nor U8855 (N_8855,In_1498,In_2556);
nand U8856 (N_8856,In_2629,In_415);
and U8857 (N_8857,In_2911,In_2764);
xor U8858 (N_8858,In_686,In_1625);
nor U8859 (N_8859,In_1340,In_1450);
and U8860 (N_8860,In_2195,In_412);
xor U8861 (N_8861,In_314,In_280);
or U8862 (N_8862,In_2178,In_2365);
xnor U8863 (N_8863,In_779,In_2361);
and U8864 (N_8864,In_149,In_1458);
nand U8865 (N_8865,In_2169,In_2034);
xnor U8866 (N_8866,In_710,In_1295);
xnor U8867 (N_8867,In_391,In_2348);
and U8868 (N_8868,In_2302,In_866);
nand U8869 (N_8869,In_1633,In_247);
or U8870 (N_8870,In_429,In_1447);
or U8871 (N_8871,In_173,In_2535);
nand U8872 (N_8872,In_1023,In_2490);
and U8873 (N_8873,In_1545,In_2861);
xor U8874 (N_8874,In_2893,In_8);
nor U8875 (N_8875,In_1563,In_2278);
or U8876 (N_8876,In_1857,In_1346);
and U8877 (N_8877,In_1262,In_2261);
and U8878 (N_8878,In_796,In_2015);
or U8879 (N_8879,In_2958,In_1305);
or U8880 (N_8880,In_2960,In_169);
or U8881 (N_8881,In_446,In_1015);
and U8882 (N_8882,In_870,In_2865);
or U8883 (N_8883,In_1620,In_932);
nand U8884 (N_8884,In_2522,In_280);
xnor U8885 (N_8885,In_1477,In_1725);
nor U8886 (N_8886,In_1858,In_381);
and U8887 (N_8887,In_237,In_318);
xor U8888 (N_8888,In_111,In_721);
nor U8889 (N_8889,In_1878,In_1428);
or U8890 (N_8890,In_2071,In_693);
xnor U8891 (N_8891,In_2158,In_2321);
xnor U8892 (N_8892,In_1823,In_2317);
or U8893 (N_8893,In_1238,In_2962);
or U8894 (N_8894,In_1061,In_799);
nor U8895 (N_8895,In_2837,In_1905);
nand U8896 (N_8896,In_1494,In_2596);
nor U8897 (N_8897,In_2006,In_461);
or U8898 (N_8898,In_2065,In_2583);
xor U8899 (N_8899,In_1632,In_1972);
or U8900 (N_8900,In_1649,In_1772);
nand U8901 (N_8901,In_2011,In_78);
xor U8902 (N_8902,In_1970,In_2393);
or U8903 (N_8903,In_1488,In_669);
nor U8904 (N_8904,In_43,In_692);
nor U8905 (N_8905,In_7,In_2062);
xor U8906 (N_8906,In_1835,In_831);
nand U8907 (N_8907,In_1055,In_307);
nand U8908 (N_8908,In_1131,In_2459);
nand U8909 (N_8909,In_1924,In_107);
xor U8910 (N_8910,In_492,In_1900);
nor U8911 (N_8911,In_663,In_2970);
or U8912 (N_8912,In_2237,In_1570);
xnor U8913 (N_8913,In_2907,In_940);
nor U8914 (N_8914,In_1661,In_1738);
xnor U8915 (N_8915,In_1206,In_1843);
xnor U8916 (N_8916,In_363,In_400);
nand U8917 (N_8917,In_2988,In_1765);
nand U8918 (N_8918,In_1509,In_2182);
or U8919 (N_8919,In_2278,In_1430);
nand U8920 (N_8920,In_1491,In_536);
or U8921 (N_8921,In_1321,In_1595);
and U8922 (N_8922,In_787,In_2054);
nand U8923 (N_8923,In_1995,In_2296);
or U8924 (N_8924,In_1099,In_1783);
or U8925 (N_8925,In_959,In_2738);
or U8926 (N_8926,In_382,In_543);
xnor U8927 (N_8927,In_393,In_2313);
and U8928 (N_8928,In_457,In_2740);
nor U8929 (N_8929,In_293,In_1851);
nor U8930 (N_8930,In_1455,In_115);
nand U8931 (N_8931,In_80,In_774);
and U8932 (N_8932,In_2095,In_1917);
or U8933 (N_8933,In_1272,In_2327);
and U8934 (N_8934,In_2581,In_2813);
nor U8935 (N_8935,In_186,In_550);
xor U8936 (N_8936,In_602,In_2444);
xor U8937 (N_8937,In_1945,In_727);
or U8938 (N_8938,In_2793,In_2808);
xnor U8939 (N_8939,In_2542,In_1962);
or U8940 (N_8940,In_2645,In_345);
xnor U8941 (N_8941,In_1762,In_2438);
xnor U8942 (N_8942,In_1562,In_89);
and U8943 (N_8943,In_2234,In_636);
nor U8944 (N_8944,In_1425,In_1870);
xor U8945 (N_8945,In_752,In_2107);
and U8946 (N_8946,In_105,In_2871);
or U8947 (N_8947,In_2569,In_193);
xnor U8948 (N_8948,In_1037,In_1530);
nor U8949 (N_8949,In_778,In_1159);
xnor U8950 (N_8950,In_2804,In_1688);
nand U8951 (N_8951,In_2944,In_1691);
and U8952 (N_8952,In_1298,In_1226);
or U8953 (N_8953,In_118,In_2630);
or U8954 (N_8954,In_1414,In_214);
and U8955 (N_8955,In_970,In_1296);
nor U8956 (N_8956,In_956,In_2941);
nand U8957 (N_8957,In_909,In_669);
xnor U8958 (N_8958,In_2545,In_572);
xnor U8959 (N_8959,In_1598,In_2882);
and U8960 (N_8960,In_2465,In_2272);
and U8961 (N_8961,In_1907,In_1805);
xor U8962 (N_8962,In_617,In_2075);
nor U8963 (N_8963,In_83,In_2497);
nand U8964 (N_8964,In_379,In_2943);
xnor U8965 (N_8965,In_1362,In_1160);
nor U8966 (N_8966,In_2204,In_191);
xnor U8967 (N_8967,In_249,In_663);
nand U8968 (N_8968,In_659,In_2001);
and U8969 (N_8969,In_1502,In_2335);
xnor U8970 (N_8970,In_1494,In_2864);
or U8971 (N_8971,In_252,In_1340);
or U8972 (N_8972,In_835,In_2542);
and U8973 (N_8973,In_2950,In_1327);
and U8974 (N_8974,In_2762,In_350);
and U8975 (N_8975,In_2207,In_177);
xnor U8976 (N_8976,In_2205,In_1394);
xor U8977 (N_8977,In_215,In_2987);
nand U8978 (N_8978,In_2734,In_767);
nand U8979 (N_8979,In_191,In_2471);
nor U8980 (N_8980,In_2058,In_2216);
nor U8981 (N_8981,In_1732,In_543);
nand U8982 (N_8982,In_480,In_1651);
and U8983 (N_8983,In_2356,In_2933);
nand U8984 (N_8984,In_1107,In_2164);
or U8985 (N_8985,In_1932,In_593);
xnor U8986 (N_8986,In_1601,In_1649);
and U8987 (N_8987,In_1132,In_972);
xnor U8988 (N_8988,In_301,In_1560);
nand U8989 (N_8989,In_318,In_1506);
nor U8990 (N_8990,In_1298,In_2618);
nor U8991 (N_8991,In_2088,In_991);
xor U8992 (N_8992,In_2763,In_1490);
or U8993 (N_8993,In_973,In_1628);
or U8994 (N_8994,In_320,In_1991);
nand U8995 (N_8995,In_1233,In_1221);
xor U8996 (N_8996,In_2587,In_1229);
or U8997 (N_8997,In_221,In_2964);
nor U8998 (N_8998,In_2362,In_2546);
and U8999 (N_8999,In_2796,In_2459);
nand U9000 (N_9000,In_1427,In_1039);
and U9001 (N_9001,In_1065,In_1256);
xor U9002 (N_9002,In_698,In_1689);
nand U9003 (N_9003,In_319,In_2377);
xor U9004 (N_9004,In_2206,In_1910);
xnor U9005 (N_9005,In_2898,In_2440);
nand U9006 (N_9006,In_2066,In_980);
xnor U9007 (N_9007,In_722,In_2666);
or U9008 (N_9008,In_2265,In_619);
or U9009 (N_9009,In_642,In_1906);
nor U9010 (N_9010,In_2334,In_259);
and U9011 (N_9011,In_2365,In_2716);
or U9012 (N_9012,In_1736,In_1864);
xor U9013 (N_9013,In_1627,In_43);
xnor U9014 (N_9014,In_659,In_432);
and U9015 (N_9015,In_471,In_2124);
or U9016 (N_9016,In_2930,In_2611);
nor U9017 (N_9017,In_2725,In_736);
and U9018 (N_9018,In_644,In_1765);
or U9019 (N_9019,In_2241,In_710);
nor U9020 (N_9020,In_347,In_1557);
or U9021 (N_9021,In_1298,In_245);
xnor U9022 (N_9022,In_1157,In_1125);
nor U9023 (N_9023,In_1873,In_2745);
nor U9024 (N_9024,In_1134,In_2318);
or U9025 (N_9025,In_1734,In_2482);
or U9026 (N_9026,In_779,In_1184);
and U9027 (N_9027,In_2498,In_2436);
nand U9028 (N_9028,In_652,In_2728);
xnor U9029 (N_9029,In_1473,In_2681);
and U9030 (N_9030,In_2157,In_1840);
nand U9031 (N_9031,In_811,In_1950);
xnor U9032 (N_9032,In_1990,In_2260);
xnor U9033 (N_9033,In_1143,In_1151);
xor U9034 (N_9034,In_1118,In_694);
or U9035 (N_9035,In_1316,In_868);
xnor U9036 (N_9036,In_1806,In_1994);
nand U9037 (N_9037,In_259,In_1116);
nor U9038 (N_9038,In_1610,In_1393);
nand U9039 (N_9039,In_1779,In_1248);
nand U9040 (N_9040,In_524,In_1210);
or U9041 (N_9041,In_1051,In_1156);
nor U9042 (N_9042,In_2393,In_80);
and U9043 (N_9043,In_244,In_1062);
or U9044 (N_9044,In_2699,In_940);
or U9045 (N_9045,In_2144,In_2443);
and U9046 (N_9046,In_2260,In_2999);
or U9047 (N_9047,In_629,In_2641);
nor U9048 (N_9048,In_2328,In_1162);
xnor U9049 (N_9049,In_2851,In_1170);
and U9050 (N_9050,In_2670,In_1107);
nand U9051 (N_9051,In_2650,In_513);
or U9052 (N_9052,In_1382,In_458);
and U9053 (N_9053,In_317,In_2858);
and U9054 (N_9054,In_2660,In_2202);
nand U9055 (N_9055,In_2664,In_2402);
xor U9056 (N_9056,In_2171,In_868);
and U9057 (N_9057,In_1958,In_1683);
or U9058 (N_9058,In_762,In_1141);
and U9059 (N_9059,In_2283,In_2538);
or U9060 (N_9060,In_543,In_192);
nor U9061 (N_9061,In_926,In_1084);
nand U9062 (N_9062,In_1206,In_1314);
nor U9063 (N_9063,In_109,In_225);
or U9064 (N_9064,In_835,In_1995);
nand U9065 (N_9065,In_2017,In_1926);
or U9066 (N_9066,In_1543,In_2570);
nand U9067 (N_9067,In_472,In_202);
nor U9068 (N_9068,In_72,In_1150);
xor U9069 (N_9069,In_1469,In_1336);
or U9070 (N_9070,In_1242,In_2038);
and U9071 (N_9071,In_1997,In_1249);
xnor U9072 (N_9072,In_5,In_1621);
and U9073 (N_9073,In_773,In_2008);
or U9074 (N_9074,In_873,In_1648);
or U9075 (N_9075,In_1434,In_945);
xor U9076 (N_9076,In_249,In_2934);
nand U9077 (N_9077,In_323,In_1345);
or U9078 (N_9078,In_2995,In_1222);
nor U9079 (N_9079,In_1100,In_686);
or U9080 (N_9080,In_765,In_703);
or U9081 (N_9081,In_683,In_2286);
and U9082 (N_9082,In_2601,In_2218);
nand U9083 (N_9083,In_1562,In_488);
and U9084 (N_9084,In_2369,In_2539);
nor U9085 (N_9085,In_2389,In_677);
or U9086 (N_9086,In_375,In_2255);
nor U9087 (N_9087,In_2372,In_2232);
nand U9088 (N_9088,In_2567,In_916);
xor U9089 (N_9089,In_2099,In_411);
xor U9090 (N_9090,In_879,In_2703);
nor U9091 (N_9091,In_2901,In_1953);
nor U9092 (N_9092,In_2053,In_1909);
xor U9093 (N_9093,In_1128,In_1533);
xnor U9094 (N_9094,In_2726,In_432);
or U9095 (N_9095,In_2618,In_371);
or U9096 (N_9096,In_2701,In_2965);
xor U9097 (N_9097,In_39,In_2152);
nand U9098 (N_9098,In_1957,In_1917);
nand U9099 (N_9099,In_749,In_1510);
and U9100 (N_9100,In_1522,In_2183);
and U9101 (N_9101,In_2162,In_1285);
and U9102 (N_9102,In_2570,In_195);
nand U9103 (N_9103,In_1909,In_1174);
or U9104 (N_9104,In_1398,In_68);
nand U9105 (N_9105,In_2536,In_1520);
xnor U9106 (N_9106,In_284,In_2176);
nor U9107 (N_9107,In_835,In_1871);
nor U9108 (N_9108,In_1788,In_1408);
xnor U9109 (N_9109,In_1437,In_308);
nor U9110 (N_9110,In_410,In_530);
nand U9111 (N_9111,In_654,In_2787);
nand U9112 (N_9112,In_2101,In_2611);
and U9113 (N_9113,In_2414,In_1785);
and U9114 (N_9114,In_2513,In_430);
xnor U9115 (N_9115,In_1002,In_2565);
and U9116 (N_9116,In_1608,In_667);
or U9117 (N_9117,In_328,In_638);
xor U9118 (N_9118,In_744,In_37);
and U9119 (N_9119,In_1389,In_2654);
nor U9120 (N_9120,In_1666,In_971);
nor U9121 (N_9121,In_8,In_585);
or U9122 (N_9122,In_1661,In_2788);
xnor U9123 (N_9123,In_2007,In_2516);
or U9124 (N_9124,In_1844,In_182);
or U9125 (N_9125,In_2904,In_1121);
nand U9126 (N_9126,In_459,In_918);
xor U9127 (N_9127,In_2310,In_600);
and U9128 (N_9128,In_2010,In_2791);
or U9129 (N_9129,In_2983,In_819);
xor U9130 (N_9130,In_2753,In_261);
nand U9131 (N_9131,In_1042,In_2931);
nor U9132 (N_9132,In_1021,In_1143);
and U9133 (N_9133,In_77,In_1195);
and U9134 (N_9134,In_317,In_2290);
xnor U9135 (N_9135,In_2534,In_96);
nand U9136 (N_9136,In_788,In_2763);
xor U9137 (N_9137,In_1874,In_385);
xor U9138 (N_9138,In_1610,In_1202);
xnor U9139 (N_9139,In_1756,In_1484);
xor U9140 (N_9140,In_2063,In_2916);
and U9141 (N_9141,In_1198,In_2489);
nor U9142 (N_9142,In_851,In_1190);
and U9143 (N_9143,In_2476,In_1762);
nor U9144 (N_9144,In_2859,In_825);
and U9145 (N_9145,In_2607,In_1685);
nor U9146 (N_9146,In_2140,In_2881);
and U9147 (N_9147,In_1557,In_2914);
xnor U9148 (N_9148,In_1679,In_539);
nand U9149 (N_9149,In_212,In_2008);
xnor U9150 (N_9150,In_1073,In_1760);
xor U9151 (N_9151,In_1977,In_356);
and U9152 (N_9152,In_193,In_2848);
nand U9153 (N_9153,In_2974,In_891);
nand U9154 (N_9154,In_894,In_2951);
nor U9155 (N_9155,In_295,In_658);
nor U9156 (N_9156,In_173,In_2520);
and U9157 (N_9157,In_850,In_134);
xor U9158 (N_9158,In_1324,In_414);
and U9159 (N_9159,In_2256,In_956);
xnor U9160 (N_9160,In_2459,In_154);
or U9161 (N_9161,In_2422,In_1359);
nor U9162 (N_9162,In_1127,In_1364);
xor U9163 (N_9163,In_174,In_2438);
xor U9164 (N_9164,In_1819,In_1838);
xor U9165 (N_9165,In_2562,In_2480);
nand U9166 (N_9166,In_40,In_2250);
nand U9167 (N_9167,In_103,In_2041);
or U9168 (N_9168,In_1593,In_817);
xor U9169 (N_9169,In_401,In_1251);
xor U9170 (N_9170,In_1255,In_2578);
nand U9171 (N_9171,In_1179,In_865);
nor U9172 (N_9172,In_1115,In_2721);
xor U9173 (N_9173,In_1722,In_75);
or U9174 (N_9174,In_1979,In_2033);
nand U9175 (N_9175,In_2092,In_1347);
and U9176 (N_9176,In_576,In_2237);
nor U9177 (N_9177,In_186,In_407);
nand U9178 (N_9178,In_1983,In_1532);
nor U9179 (N_9179,In_11,In_175);
xnor U9180 (N_9180,In_2449,In_2214);
xnor U9181 (N_9181,In_500,In_575);
or U9182 (N_9182,In_2707,In_1216);
nor U9183 (N_9183,In_1510,In_1229);
and U9184 (N_9184,In_1768,In_2813);
or U9185 (N_9185,In_2981,In_1629);
and U9186 (N_9186,In_1788,In_2165);
nand U9187 (N_9187,In_2054,In_1343);
xnor U9188 (N_9188,In_2999,In_1407);
nor U9189 (N_9189,In_1276,In_1075);
xor U9190 (N_9190,In_1494,In_2975);
nor U9191 (N_9191,In_303,In_2949);
or U9192 (N_9192,In_194,In_1115);
and U9193 (N_9193,In_568,In_2261);
nor U9194 (N_9194,In_1979,In_2116);
nor U9195 (N_9195,In_1860,In_110);
and U9196 (N_9196,In_2706,In_2513);
or U9197 (N_9197,In_870,In_2438);
or U9198 (N_9198,In_2687,In_1938);
or U9199 (N_9199,In_2644,In_246);
xor U9200 (N_9200,In_2558,In_1953);
or U9201 (N_9201,In_2417,In_146);
nand U9202 (N_9202,In_656,In_348);
or U9203 (N_9203,In_604,In_198);
or U9204 (N_9204,In_2618,In_1471);
or U9205 (N_9205,In_1544,In_788);
xor U9206 (N_9206,In_2543,In_2621);
or U9207 (N_9207,In_1035,In_1494);
nand U9208 (N_9208,In_1559,In_880);
and U9209 (N_9209,In_1990,In_1435);
nor U9210 (N_9210,In_2824,In_2832);
and U9211 (N_9211,In_1446,In_2300);
and U9212 (N_9212,In_104,In_1981);
nand U9213 (N_9213,In_2637,In_765);
and U9214 (N_9214,In_642,In_1319);
nand U9215 (N_9215,In_2386,In_2106);
and U9216 (N_9216,In_251,In_754);
or U9217 (N_9217,In_596,In_2315);
nand U9218 (N_9218,In_1990,In_1057);
xor U9219 (N_9219,In_795,In_840);
and U9220 (N_9220,In_812,In_1334);
nand U9221 (N_9221,In_2703,In_2011);
xor U9222 (N_9222,In_2817,In_938);
or U9223 (N_9223,In_677,In_979);
nor U9224 (N_9224,In_2162,In_40);
nor U9225 (N_9225,In_1348,In_2056);
and U9226 (N_9226,In_928,In_839);
nand U9227 (N_9227,In_164,In_2563);
and U9228 (N_9228,In_767,In_1347);
xor U9229 (N_9229,In_1321,In_2121);
nor U9230 (N_9230,In_1729,In_1850);
and U9231 (N_9231,In_1432,In_835);
and U9232 (N_9232,In_1658,In_707);
and U9233 (N_9233,In_973,In_1115);
xnor U9234 (N_9234,In_1831,In_1746);
nand U9235 (N_9235,In_2859,In_2514);
nand U9236 (N_9236,In_1265,In_2751);
nor U9237 (N_9237,In_1783,In_511);
and U9238 (N_9238,In_1596,In_342);
and U9239 (N_9239,In_514,In_2385);
xor U9240 (N_9240,In_2651,In_2229);
xnor U9241 (N_9241,In_1281,In_514);
nand U9242 (N_9242,In_2795,In_683);
or U9243 (N_9243,In_1247,In_2921);
nor U9244 (N_9244,In_1354,In_1737);
and U9245 (N_9245,In_670,In_397);
nor U9246 (N_9246,In_2129,In_954);
nand U9247 (N_9247,In_2342,In_1376);
and U9248 (N_9248,In_726,In_2059);
nand U9249 (N_9249,In_1020,In_1999);
and U9250 (N_9250,In_2707,In_1008);
xnor U9251 (N_9251,In_1582,In_2199);
or U9252 (N_9252,In_284,In_2922);
or U9253 (N_9253,In_1502,In_2449);
nor U9254 (N_9254,In_1848,In_2697);
nand U9255 (N_9255,In_1421,In_325);
and U9256 (N_9256,In_799,In_2753);
nand U9257 (N_9257,In_2469,In_2048);
xor U9258 (N_9258,In_120,In_996);
nand U9259 (N_9259,In_1530,In_80);
nand U9260 (N_9260,In_860,In_2085);
nor U9261 (N_9261,In_1532,In_789);
and U9262 (N_9262,In_707,In_1572);
xnor U9263 (N_9263,In_330,In_1245);
nor U9264 (N_9264,In_2771,In_1179);
or U9265 (N_9265,In_368,In_848);
or U9266 (N_9266,In_1614,In_1533);
xnor U9267 (N_9267,In_2062,In_2979);
or U9268 (N_9268,In_2773,In_1977);
or U9269 (N_9269,In_973,In_2133);
nand U9270 (N_9270,In_830,In_163);
xor U9271 (N_9271,In_290,In_661);
nand U9272 (N_9272,In_453,In_2970);
nand U9273 (N_9273,In_2721,In_2935);
nor U9274 (N_9274,In_119,In_1685);
xor U9275 (N_9275,In_1839,In_2882);
and U9276 (N_9276,In_725,In_2372);
or U9277 (N_9277,In_2328,In_1181);
nor U9278 (N_9278,In_1290,In_772);
and U9279 (N_9279,In_179,In_2686);
nor U9280 (N_9280,In_1694,In_1536);
or U9281 (N_9281,In_2271,In_1378);
or U9282 (N_9282,In_1535,In_1562);
and U9283 (N_9283,In_1394,In_2911);
or U9284 (N_9284,In_1566,In_926);
or U9285 (N_9285,In_366,In_558);
and U9286 (N_9286,In_217,In_2734);
nor U9287 (N_9287,In_2513,In_2067);
xnor U9288 (N_9288,In_1361,In_1756);
and U9289 (N_9289,In_626,In_1448);
and U9290 (N_9290,In_1604,In_83);
nor U9291 (N_9291,In_1632,In_1826);
nor U9292 (N_9292,In_112,In_31);
or U9293 (N_9293,In_1744,In_1421);
nor U9294 (N_9294,In_1198,In_779);
nor U9295 (N_9295,In_2624,In_1686);
nand U9296 (N_9296,In_928,In_2337);
nand U9297 (N_9297,In_2764,In_157);
and U9298 (N_9298,In_1290,In_1349);
and U9299 (N_9299,In_952,In_2978);
xnor U9300 (N_9300,In_2038,In_1378);
xor U9301 (N_9301,In_2503,In_370);
xor U9302 (N_9302,In_1883,In_1734);
nor U9303 (N_9303,In_2479,In_49);
nor U9304 (N_9304,In_566,In_553);
nor U9305 (N_9305,In_1262,In_1491);
xor U9306 (N_9306,In_318,In_660);
and U9307 (N_9307,In_1393,In_2688);
nand U9308 (N_9308,In_1158,In_1968);
nor U9309 (N_9309,In_1662,In_1458);
or U9310 (N_9310,In_1452,In_2178);
nand U9311 (N_9311,In_1325,In_2339);
nand U9312 (N_9312,In_1767,In_1552);
nor U9313 (N_9313,In_1673,In_1276);
or U9314 (N_9314,In_954,In_2694);
and U9315 (N_9315,In_1558,In_1665);
and U9316 (N_9316,In_626,In_674);
xor U9317 (N_9317,In_886,In_2101);
or U9318 (N_9318,In_612,In_2081);
nand U9319 (N_9319,In_2368,In_1159);
nand U9320 (N_9320,In_929,In_1584);
and U9321 (N_9321,In_1371,In_408);
nand U9322 (N_9322,In_2584,In_1256);
nor U9323 (N_9323,In_862,In_2259);
and U9324 (N_9324,In_1854,In_250);
xnor U9325 (N_9325,In_2212,In_2666);
and U9326 (N_9326,In_815,In_581);
and U9327 (N_9327,In_1496,In_946);
or U9328 (N_9328,In_2006,In_145);
or U9329 (N_9329,In_1985,In_2148);
and U9330 (N_9330,In_954,In_1356);
nand U9331 (N_9331,In_2872,In_1007);
nand U9332 (N_9332,In_2472,In_2637);
nor U9333 (N_9333,In_1388,In_2499);
nand U9334 (N_9334,In_2197,In_1498);
and U9335 (N_9335,In_928,In_1805);
nand U9336 (N_9336,In_526,In_2342);
nand U9337 (N_9337,In_2377,In_1434);
xnor U9338 (N_9338,In_792,In_2489);
or U9339 (N_9339,In_1504,In_1845);
nor U9340 (N_9340,In_2877,In_1768);
and U9341 (N_9341,In_2529,In_1052);
xor U9342 (N_9342,In_166,In_2666);
nor U9343 (N_9343,In_2775,In_1175);
nor U9344 (N_9344,In_1620,In_277);
xor U9345 (N_9345,In_783,In_242);
nand U9346 (N_9346,In_2135,In_2255);
and U9347 (N_9347,In_1751,In_2608);
nor U9348 (N_9348,In_434,In_1011);
and U9349 (N_9349,In_2905,In_285);
or U9350 (N_9350,In_422,In_1114);
or U9351 (N_9351,In_1241,In_1645);
and U9352 (N_9352,In_2691,In_2762);
and U9353 (N_9353,In_1003,In_2466);
or U9354 (N_9354,In_1426,In_2809);
or U9355 (N_9355,In_2204,In_170);
nand U9356 (N_9356,In_1544,In_859);
xor U9357 (N_9357,In_2775,In_1249);
or U9358 (N_9358,In_1298,In_2789);
nor U9359 (N_9359,In_421,In_2496);
nor U9360 (N_9360,In_864,In_545);
or U9361 (N_9361,In_474,In_2303);
xor U9362 (N_9362,In_503,In_708);
nand U9363 (N_9363,In_2577,In_2293);
xnor U9364 (N_9364,In_1747,In_1213);
and U9365 (N_9365,In_1155,In_538);
or U9366 (N_9366,In_1247,In_569);
xnor U9367 (N_9367,In_919,In_2883);
or U9368 (N_9368,In_892,In_1994);
xor U9369 (N_9369,In_1512,In_2703);
nor U9370 (N_9370,In_1035,In_2295);
or U9371 (N_9371,In_2742,In_703);
nor U9372 (N_9372,In_1687,In_129);
nand U9373 (N_9373,In_2095,In_444);
nor U9374 (N_9374,In_2652,In_1215);
and U9375 (N_9375,In_826,In_2666);
and U9376 (N_9376,In_2337,In_1960);
xor U9377 (N_9377,In_1080,In_2512);
or U9378 (N_9378,In_1742,In_189);
nor U9379 (N_9379,In_985,In_2875);
or U9380 (N_9380,In_2686,In_2785);
or U9381 (N_9381,In_859,In_125);
nor U9382 (N_9382,In_1535,In_1418);
nand U9383 (N_9383,In_871,In_1250);
nor U9384 (N_9384,In_906,In_441);
and U9385 (N_9385,In_537,In_2714);
and U9386 (N_9386,In_2267,In_2435);
nand U9387 (N_9387,In_1118,In_2555);
and U9388 (N_9388,In_460,In_2773);
nor U9389 (N_9389,In_1057,In_2098);
nor U9390 (N_9390,In_799,In_2624);
nand U9391 (N_9391,In_1914,In_2806);
and U9392 (N_9392,In_1559,In_63);
nand U9393 (N_9393,In_1858,In_143);
nand U9394 (N_9394,In_2009,In_1297);
nor U9395 (N_9395,In_955,In_1222);
nand U9396 (N_9396,In_2804,In_1420);
or U9397 (N_9397,In_645,In_1728);
nand U9398 (N_9398,In_741,In_1325);
or U9399 (N_9399,In_329,In_1464);
or U9400 (N_9400,In_915,In_1595);
nand U9401 (N_9401,In_349,In_1168);
or U9402 (N_9402,In_217,In_359);
xnor U9403 (N_9403,In_2400,In_2717);
xor U9404 (N_9404,In_1171,In_2275);
nand U9405 (N_9405,In_1820,In_367);
xor U9406 (N_9406,In_624,In_317);
nand U9407 (N_9407,In_1307,In_507);
and U9408 (N_9408,In_495,In_1688);
nand U9409 (N_9409,In_800,In_598);
nor U9410 (N_9410,In_1468,In_2472);
and U9411 (N_9411,In_1854,In_1891);
nor U9412 (N_9412,In_1260,In_258);
xor U9413 (N_9413,In_30,In_1840);
nor U9414 (N_9414,In_506,In_940);
or U9415 (N_9415,In_1432,In_2774);
xnor U9416 (N_9416,In_2396,In_1803);
xor U9417 (N_9417,In_360,In_265);
xnor U9418 (N_9418,In_2484,In_1951);
and U9419 (N_9419,In_1226,In_168);
nor U9420 (N_9420,In_564,In_2383);
or U9421 (N_9421,In_2866,In_614);
or U9422 (N_9422,In_723,In_2757);
or U9423 (N_9423,In_2419,In_2940);
and U9424 (N_9424,In_2229,In_1951);
nand U9425 (N_9425,In_2026,In_277);
nor U9426 (N_9426,In_1722,In_1228);
xnor U9427 (N_9427,In_1938,In_2106);
xor U9428 (N_9428,In_1661,In_2465);
or U9429 (N_9429,In_2725,In_1893);
and U9430 (N_9430,In_1789,In_756);
and U9431 (N_9431,In_93,In_2397);
xnor U9432 (N_9432,In_2754,In_2833);
nand U9433 (N_9433,In_2778,In_1088);
xnor U9434 (N_9434,In_1786,In_1241);
xor U9435 (N_9435,In_807,In_2316);
and U9436 (N_9436,In_960,In_2997);
or U9437 (N_9437,In_2257,In_471);
or U9438 (N_9438,In_2806,In_1998);
xor U9439 (N_9439,In_1204,In_109);
and U9440 (N_9440,In_2374,In_2778);
and U9441 (N_9441,In_1175,In_855);
xor U9442 (N_9442,In_1323,In_2098);
and U9443 (N_9443,In_2446,In_2993);
xor U9444 (N_9444,In_1903,In_1651);
nor U9445 (N_9445,In_2745,In_1006);
or U9446 (N_9446,In_1632,In_2801);
and U9447 (N_9447,In_1694,In_1485);
or U9448 (N_9448,In_1752,In_1071);
xnor U9449 (N_9449,In_909,In_1289);
or U9450 (N_9450,In_2658,In_2578);
nor U9451 (N_9451,In_2173,In_1665);
nand U9452 (N_9452,In_300,In_285);
xnor U9453 (N_9453,In_620,In_2494);
and U9454 (N_9454,In_199,In_527);
and U9455 (N_9455,In_2715,In_2657);
or U9456 (N_9456,In_2371,In_2401);
or U9457 (N_9457,In_2886,In_2963);
nand U9458 (N_9458,In_1017,In_239);
xor U9459 (N_9459,In_73,In_660);
nor U9460 (N_9460,In_618,In_426);
xor U9461 (N_9461,In_1306,In_2374);
nand U9462 (N_9462,In_2409,In_2932);
and U9463 (N_9463,In_1804,In_2157);
xor U9464 (N_9464,In_1817,In_1453);
and U9465 (N_9465,In_2139,In_69);
nor U9466 (N_9466,In_1104,In_2795);
nand U9467 (N_9467,In_739,In_2637);
and U9468 (N_9468,In_530,In_415);
nand U9469 (N_9469,In_2845,In_2280);
nand U9470 (N_9470,In_562,In_2034);
and U9471 (N_9471,In_191,In_219);
xor U9472 (N_9472,In_2051,In_2048);
and U9473 (N_9473,In_1397,In_1656);
xnor U9474 (N_9474,In_174,In_1256);
nor U9475 (N_9475,In_1638,In_2370);
or U9476 (N_9476,In_1681,In_970);
and U9477 (N_9477,In_2669,In_2362);
nand U9478 (N_9478,In_2736,In_1530);
or U9479 (N_9479,In_100,In_491);
nand U9480 (N_9480,In_999,In_1636);
and U9481 (N_9481,In_2613,In_1346);
and U9482 (N_9482,In_2133,In_2253);
and U9483 (N_9483,In_1404,In_262);
or U9484 (N_9484,In_515,In_2584);
nor U9485 (N_9485,In_2645,In_1023);
xor U9486 (N_9486,In_594,In_861);
and U9487 (N_9487,In_2234,In_84);
nand U9488 (N_9488,In_449,In_269);
nand U9489 (N_9489,In_722,In_1609);
or U9490 (N_9490,In_1128,In_321);
xnor U9491 (N_9491,In_2126,In_2354);
xnor U9492 (N_9492,In_2059,In_606);
nand U9493 (N_9493,In_1723,In_1816);
nand U9494 (N_9494,In_802,In_773);
or U9495 (N_9495,In_1521,In_1153);
nor U9496 (N_9496,In_1514,In_2410);
or U9497 (N_9497,In_2876,In_2021);
xor U9498 (N_9498,In_2543,In_653);
nand U9499 (N_9499,In_734,In_2145);
or U9500 (N_9500,In_1163,In_1936);
and U9501 (N_9501,In_2403,In_2917);
xor U9502 (N_9502,In_911,In_485);
nor U9503 (N_9503,In_815,In_282);
or U9504 (N_9504,In_236,In_2748);
xnor U9505 (N_9505,In_2259,In_2530);
xnor U9506 (N_9506,In_1243,In_354);
xnor U9507 (N_9507,In_1475,In_1926);
xor U9508 (N_9508,In_201,In_697);
and U9509 (N_9509,In_635,In_670);
or U9510 (N_9510,In_2661,In_2867);
nand U9511 (N_9511,In_1343,In_2408);
xnor U9512 (N_9512,In_2852,In_703);
nor U9513 (N_9513,In_106,In_564);
or U9514 (N_9514,In_1546,In_2619);
nand U9515 (N_9515,In_1889,In_2472);
or U9516 (N_9516,In_1033,In_583);
or U9517 (N_9517,In_212,In_1466);
nor U9518 (N_9518,In_1225,In_1934);
or U9519 (N_9519,In_1127,In_1071);
or U9520 (N_9520,In_430,In_291);
nor U9521 (N_9521,In_1749,In_547);
nor U9522 (N_9522,In_2894,In_2198);
xnor U9523 (N_9523,In_2944,In_873);
or U9524 (N_9524,In_2998,In_1113);
or U9525 (N_9525,In_888,In_1675);
or U9526 (N_9526,In_1265,In_2546);
nor U9527 (N_9527,In_2657,In_1048);
nand U9528 (N_9528,In_2876,In_190);
or U9529 (N_9529,In_2364,In_1097);
or U9530 (N_9530,In_1926,In_2073);
xor U9531 (N_9531,In_1583,In_214);
xnor U9532 (N_9532,In_519,In_2621);
xor U9533 (N_9533,In_250,In_1995);
or U9534 (N_9534,In_1838,In_1249);
xor U9535 (N_9535,In_578,In_312);
nand U9536 (N_9536,In_2491,In_2813);
nand U9537 (N_9537,In_1911,In_366);
xnor U9538 (N_9538,In_1832,In_79);
xor U9539 (N_9539,In_2880,In_2844);
or U9540 (N_9540,In_2374,In_1941);
or U9541 (N_9541,In_2429,In_1452);
nand U9542 (N_9542,In_2877,In_704);
and U9543 (N_9543,In_2678,In_1178);
nand U9544 (N_9544,In_994,In_1972);
and U9545 (N_9545,In_1770,In_1624);
nor U9546 (N_9546,In_207,In_2379);
nor U9547 (N_9547,In_1458,In_1739);
and U9548 (N_9548,In_1012,In_2745);
nor U9549 (N_9549,In_100,In_2955);
nor U9550 (N_9550,In_1989,In_667);
nor U9551 (N_9551,In_2054,In_1176);
xor U9552 (N_9552,In_2502,In_686);
xor U9553 (N_9553,In_1090,In_215);
xnor U9554 (N_9554,In_1994,In_1821);
nor U9555 (N_9555,In_186,In_1765);
and U9556 (N_9556,In_353,In_1815);
nand U9557 (N_9557,In_119,In_1989);
xor U9558 (N_9558,In_2998,In_2138);
nor U9559 (N_9559,In_1542,In_2641);
xor U9560 (N_9560,In_1253,In_1786);
nor U9561 (N_9561,In_1192,In_561);
xnor U9562 (N_9562,In_1747,In_1487);
nand U9563 (N_9563,In_530,In_1745);
or U9564 (N_9564,In_1052,In_2988);
nand U9565 (N_9565,In_1714,In_2821);
and U9566 (N_9566,In_843,In_649);
xor U9567 (N_9567,In_2581,In_1060);
nor U9568 (N_9568,In_1363,In_620);
or U9569 (N_9569,In_2729,In_1516);
nand U9570 (N_9570,In_483,In_2940);
or U9571 (N_9571,In_1301,In_2046);
xor U9572 (N_9572,In_1895,In_2675);
or U9573 (N_9573,In_870,In_2899);
nor U9574 (N_9574,In_1337,In_817);
xnor U9575 (N_9575,In_665,In_1266);
nor U9576 (N_9576,In_2065,In_2329);
xnor U9577 (N_9577,In_1640,In_2894);
xor U9578 (N_9578,In_138,In_2517);
nor U9579 (N_9579,In_1802,In_1763);
or U9580 (N_9580,In_2643,In_786);
or U9581 (N_9581,In_2918,In_2941);
nand U9582 (N_9582,In_2866,In_2756);
and U9583 (N_9583,In_1359,In_2197);
or U9584 (N_9584,In_2770,In_1224);
nor U9585 (N_9585,In_2223,In_1043);
xnor U9586 (N_9586,In_1274,In_2883);
xnor U9587 (N_9587,In_2267,In_2822);
nand U9588 (N_9588,In_314,In_309);
or U9589 (N_9589,In_1036,In_2072);
nor U9590 (N_9590,In_1216,In_478);
or U9591 (N_9591,In_624,In_1548);
and U9592 (N_9592,In_1521,In_362);
xor U9593 (N_9593,In_657,In_2397);
or U9594 (N_9594,In_2699,In_42);
nand U9595 (N_9595,In_1383,In_2845);
or U9596 (N_9596,In_2319,In_631);
or U9597 (N_9597,In_346,In_190);
nand U9598 (N_9598,In_1508,In_2217);
and U9599 (N_9599,In_1586,In_114);
xor U9600 (N_9600,In_2190,In_887);
xor U9601 (N_9601,In_513,In_2262);
or U9602 (N_9602,In_2109,In_1854);
nand U9603 (N_9603,In_1727,In_83);
nand U9604 (N_9604,In_2972,In_1898);
nand U9605 (N_9605,In_1107,In_23);
and U9606 (N_9606,In_348,In_1209);
or U9607 (N_9607,In_1540,In_2228);
nand U9608 (N_9608,In_676,In_1723);
xnor U9609 (N_9609,In_864,In_610);
nor U9610 (N_9610,In_456,In_2123);
nor U9611 (N_9611,In_1294,In_2645);
nand U9612 (N_9612,In_992,In_1156);
xnor U9613 (N_9613,In_853,In_889);
xnor U9614 (N_9614,In_47,In_1672);
xor U9615 (N_9615,In_1259,In_2209);
and U9616 (N_9616,In_1249,In_855);
and U9617 (N_9617,In_1849,In_2438);
nor U9618 (N_9618,In_814,In_241);
nand U9619 (N_9619,In_2142,In_1315);
xnor U9620 (N_9620,In_638,In_569);
or U9621 (N_9621,In_2777,In_2918);
xnor U9622 (N_9622,In_643,In_702);
or U9623 (N_9623,In_138,In_327);
nand U9624 (N_9624,In_299,In_151);
nand U9625 (N_9625,In_2535,In_1038);
and U9626 (N_9626,In_939,In_3);
nor U9627 (N_9627,In_983,In_2145);
nor U9628 (N_9628,In_1685,In_1212);
nand U9629 (N_9629,In_1793,In_1183);
xnor U9630 (N_9630,In_1810,In_701);
or U9631 (N_9631,In_204,In_2495);
and U9632 (N_9632,In_1185,In_1690);
or U9633 (N_9633,In_106,In_1950);
nand U9634 (N_9634,In_516,In_1594);
nand U9635 (N_9635,In_2249,In_739);
and U9636 (N_9636,In_1277,In_1256);
and U9637 (N_9637,In_186,In_1229);
and U9638 (N_9638,In_131,In_1014);
or U9639 (N_9639,In_226,In_1655);
nor U9640 (N_9640,In_1308,In_272);
and U9641 (N_9641,In_2014,In_1906);
nand U9642 (N_9642,In_1048,In_1867);
and U9643 (N_9643,In_588,In_560);
nor U9644 (N_9644,In_798,In_201);
nand U9645 (N_9645,In_2868,In_2253);
or U9646 (N_9646,In_396,In_1663);
nand U9647 (N_9647,In_1251,In_2682);
and U9648 (N_9648,In_1622,In_2585);
and U9649 (N_9649,In_168,In_1309);
nor U9650 (N_9650,In_1287,In_1919);
and U9651 (N_9651,In_1117,In_1982);
or U9652 (N_9652,In_2265,In_243);
nand U9653 (N_9653,In_2626,In_49);
and U9654 (N_9654,In_822,In_1330);
and U9655 (N_9655,In_1963,In_667);
or U9656 (N_9656,In_1435,In_1037);
nand U9657 (N_9657,In_596,In_2773);
nor U9658 (N_9658,In_415,In_596);
nor U9659 (N_9659,In_1464,In_1265);
nand U9660 (N_9660,In_2909,In_2165);
or U9661 (N_9661,In_2197,In_1631);
or U9662 (N_9662,In_598,In_2750);
nor U9663 (N_9663,In_932,In_185);
xor U9664 (N_9664,In_2618,In_675);
and U9665 (N_9665,In_2330,In_642);
nand U9666 (N_9666,In_883,In_2493);
and U9667 (N_9667,In_519,In_2180);
and U9668 (N_9668,In_406,In_166);
or U9669 (N_9669,In_224,In_890);
and U9670 (N_9670,In_2003,In_141);
nor U9671 (N_9671,In_1679,In_1965);
or U9672 (N_9672,In_1694,In_1840);
xnor U9673 (N_9673,In_1254,In_964);
xnor U9674 (N_9674,In_263,In_1349);
nor U9675 (N_9675,In_2579,In_579);
xor U9676 (N_9676,In_1987,In_323);
or U9677 (N_9677,In_1364,In_2472);
nor U9678 (N_9678,In_2643,In_2757);
or U9679 (N_9679,In_1150,In_2378);
xnor U9680 (N_9680,In_1769,In_85);
nand U9681 (N_9681,In_350,In_2947);
or U9682 (N_9682,In_2700,In_1884);
xor U9683 (N_9683,In_2043,In_1376);
xor U9684 (N_9684,In_1694,In_2602);
or U9685 (N_9685,In_1523,In_15);
nor U9686 (N_9686,In_2460,In_1803);
xor U9687 (N_9687,In_1796,In_2833);
xnor U9688 (N_9688,In_981,In_2345);
nand U9689 (N_9689,In_122,In_2171);
and U9690 (N_9690,In_1811,In_39);
nor U9691 (N_9691,In_344,In_409);
nand U9692 (N_9692,In_87,In_172);
nor U9693 (N_9693,In_339,In_1399);
xnor U9694 (N_9694,In_2408,In_1371);
nand U9695 (N_9695,In_660,In_1194);
xnor U9696 (N_9696,In_770,In_1558);
and U9697 (N_9697,In_176,In_984);
or U9698 (N_9698,In_375,In_1563);
nand U9699 (N_9699,In_2748,In_1080);
xor U9700 (N_9700,In_690,In_99);
nor U9701 (N_9701,In_2519,In_865);
nor U9702 (N_9702,In_461,In_2618);
xor U9703 (N_9703,In_897,In_468);
nor U9704 (N_9704,In_1420,In_1026);
or U9705 (N_9705,In_2848,In_729);
xnor U9706 (N_9706,In_1000,In_1296);
nand U9707 (N_9707,In_557,In_2437);
nand U9708 (N_9708,In_788,In_2369);
or U9709 (N_9709,In_2949,In_1912);
and U9710 (N_9710,In_2379,In_1846);
xor U9711 (N_9711,In_1071,In_2257);
and U9712 (N_9712,In_1718,In_2742);
nor U9713 (N_9713,In_62,In_463);
or U9714 (N_9714,In_363,In_2045);
or U9715 (N_9715,In_2273,In_1305);
and U9716 (N_9716,In_2705,In_2266);
nor U9717 (N_9717,In_2741,In_1077);
nor U9718 (N_9718,In_969,In_55);
or U9719 (N_9719,In_2279,In_1763);
nor U9720 (N_9720,In_547,In_1469);
xor U9721 (N_9721,In_1050,In_1353);
or U9722 (N_9722,In_2294,In_665);
nor U9723 (N_9723,In_2289,In_1585);
and U9724 (N_9724,In_1864,In_2410);
and U9725 (N_9725,In_34,In_1443);
and U9726 (N_9726,In_2389,In_447);
nand U9727 (N_9727,In_1060,In_453);
nand U9728 (N_9728,In_503,In_1224);
or U9729 (N_9729,In_2772,In_1350);
nand U9730 (N_9730,In_242,In_109);
and U9731 (N_9731,In_1935,In_2419);
and U9732 (N_9732,In_2488,In_2238);
xor U9733 (N_9733,In_651,In_145);
and U9734 (N_9734,In_480,In_477);
nand U9735 (N_9735,In_631,In_1406);
xnor U9736 (N_9736,In_1896,In_2086);
xnor U9737 (N_9737,In_1942,In_2348);
nand U9738 (N_9738,In_2153,In_528);
nor U9739 (N_9739,In_73,In_277);
nor U9740 (N_9740,In_1707,In_2952);
and U9741 (N_9741,In_142,In_555);
or U9742 (N_9742,In_266,In_787);
and U9743 (N_9743,In_1004,In_1966);
and U9744 (N_9744,In_1443,In_175);
and U9745 (N_9745,In_1166,In_1289);
nor U9746 (N_9746,In_1125,In_1273);
and U9747 (N_9747,In_2438,In_2522);
and U9748 (N_9748,In_2338,In_2202);
nand U9749 (N_9749,In_1464,In_666);
or U9750 (N_9750,In_2375,In_1129);
xor U9751 (N_9751,In_2692,In_350);
nor U9752 (N_9752,In_1528,In_2548);
nand U9753 (N_9753,In_2153,In_1379);
or U9754 (N_9754,In_1806,In_1687);
and U9755 (N_9755,In_1151,In_2196);
or U9756 (N_9756,In_1475,In_1839);
xnor U9757 (N_9757,In_432,In_2161);
or U9758 (N_9758,In_1201,In_1903);
nand U9759 (N_9759,In_1236,In_2238);
nor U9760 (N_9760,In_394,In_2594);
nand U9761 (N_9761,In_2935,In_2513);
or U9762 (N_9762,In_1818,In_1773);
nor U9763 (N_9763,In_1041,In_1554);
nor U9764 (N_9764,In_2506,In_993);
xor U9765 (N_9765,In_2090,In_1910);
nor U9766 (N_9766,In_1882,In_2131);
or U9767 (N_9767,In_2470,In_1530);
nand U9768 (N_9768,In_679,In_939);
nor U9769 (N_9769,In_2027,In_469);
and U9770 (N_9770,In_2558,In_1749);
and U9771 (N_9771,In_382,In_873);
nor U9772 (N_9772,In_2865,In_2949);
nand U9773 (N_9773,In_641,In_1267);
nand U9774 (N_9774,In_367,In_943);
nor U9775 (N_9775,In_2293,In_2357);
nor U9776 (N_9776,In_1471,In_651);
nand U9777 (N_9777,In_2053,In_503);
xor U9778 (N_9778,In_629,In_1357);
and U9779 (N_9779,In_364,In_339);
or U9780 (N_9780,In_799,In_80);
xnor U9781 (N_9781,In_2122,In_122);
xnor U9782 (N_9782,In_1936,In_1635);
nor U9783 (N_9783,In_451,In_1148);
nand U9784 (N_9784,In_314,In_2056);
and U9785 (N_9785,In_1721,In_2659);
or U9786 (N_9786,In_52,In_2926);
nand U9787 (N_9787,In_1562,In_244);
nor U9788 (N_9788,In_2084,In_2702);
xnor U9789 (N_9789,In_99,In_429);
nand U9790 (N_9790,In_1217,In_648);
or U9791 (N_9791,In_2077,In_752);
or U9792 (N_9792,In_1410,In_263);
and U9793 (N_9793,In_762,In_2717);
nor U9794 (N_9794,In_2115,In_2113);
xnor U9795 (N_9795,In_1802,In_231);
xor U9796 (N_9796,In_860,In_1459);
and U9797 (N_9797,In_1587,In_89);
nor U9798 (N_9798,In_1362,In_2619);
nor U9799 (N_9799,In_2277,In_2686);
nand U9800 (N_9800,In_226,In_1896);
and U9801 (N_9801,In_24,In_2410);
nor U9802 (N_9802,In_2962,In_590);
or U9803 (N_9803,In_2709,In_930);
nand U9804 (N_9804,In_1324,In_1057);
xor U9805 (N_9805,In_1893,In_228);
nor U9806 (N_9806,In_2477,In_1974);
or U9807 (N_9807,In_1448,In_61);
nand U9808 (N_9808,In_565,In_2647);
or U9809 (N_9809,In_1987,In_1466);
or U9810 (N_9810,In_853,In_1943);
nor U9811 (N_9811,In_2058,In_552);
nand U9812 (N_9812,In_1227,In_997);
and U9813 (N_9813,In_840,In_2890);
xnor U9814 (N_9814,In_1445,In_2715);
nor U9815 (N_9815,In_181,In_505);
or U9816 (N_9816,In_822,In_1853);
xnor U9817 (N_9817,In_1873,In_2204);
nand U9818 (N_9818,In_213,In_1088);
and U9819 (N_9819,In_93,In_651);
nor U9820 (N_9820,In_2077,In_2375);
xor U9821 (N_9821,In_1431,In_1657);
xnor U9822 (N_9822,In_294,In_1428);
nor U9823 (N_9823,In_1638,In_979);
nand U9824 (N_9824,In_877,In_775);
or U9825 (N_9825,In_1712,In_1518);
or U9826 (N_9826,In_132,In_1236);
nand U9827 (N_9827,In_183,In_2394);
and U9828 (N_9828,In_2925,In_2335);
nor U9829 (N_9829,In_1800,In_931);
and U9830 (N_9830,In_1870,In_2243);
xnor U9831 (N_9831,In_72,In_528);
nor U9832 (N_9832,In_1187,In_168);
or U9833 (N_9833,In_630,In_2958);
nor U9834 (N_9834,In_489,In_945);
xnor U9835 (N_9835,In_520,In_1527);
and U9836 (N_9836,In_2521,In_2233);
nand U9837 (N_9837,In_2220,In_2042);
xor U9838 (N_9838,In_2336,In_2642);
and U9839 (N_9839,In_2428,In_1814);
or U9840 (N_9840,In_1373,In_1444);
xnor U9841 (N_9841,In_2444,In_2475);
xor U9842 (N_9842,In_359,In_2533);
and U9843 (N_9843,In_682,In_2493);
and U9844 (N_9844,In_2682,In_2524);
nor U9845 (N_9845,In_1816,In_2881);
nand U9846 (N_9846,In_1565,In_392);
nand U9847 (N_9847,In_1577,In_1525);
or U9848 (N_9848,In_1216,In_95);
nand U9849 (N_9849,In_495,In_2726);
nand U9850 (N_9850,In_2735,In_309);
or U9851 (N_9851,In_2502,In_149);
nor U9852 (N_9852,In_2469,In_2620);
nor U9853 (N_9853,In_130,In_2464);
nand U9854 (N_9854,In_2515,In_457);
and U9855 (N_9855,In_657,In_969);
nand U9856 (N_9856,In_540,In_1713);
or U9857 (N_9857,In_1938,In_2909);
xor U9858 (N_9858,In_6,In_519);
xnor U9859 (N_9859,In_723,In_1977);
xnor U9860 (N_9860,In_2321,In_601);
nand U9861 (N_9861,In_2445,In_2975);
nor U9862 (N_9862,In_1484,In_109);
and U9863 (N_9863,In_1231,In_512);
and U9864 (N_9864,In_1729,In_1995);
nor U9865 (N_9865,In_1745,In_2304);
nand U9866 (N_9866,In_188,In_907);
and U9867 (N_9867,In_1668,In_2817);
xor U9868 (N_9868,In_2002,In_854);
nand U9869 (N_9869,In_695,In_2853);
nor U9870 (N_9870,In_2052,In_881);
nor U9871 (N_9871,In_2944,In_1582);
nor U9872 (N_9872,In_310,In_2015);
or U9873 (N_9873,In_810,In_2991);
or U9874 (N_9874,In_2383,In_2605);
nand U9875 (N_9875,In_2161,In_2389);
and U9876 (N_9876,In_1068,In_2441);
nor U9877 (N_9877,In_1003,In_2006);
nor U9878 (N_9878,In_1913,In_352);
nand U9879 (N_9879,In_1566,In_266);
nor U9880 (N_9880,In_2486,In_2059);
and U9881 (N_9881,In_2639,In_1843);
nor U9882 (N_9882,In_2614,In_476);
nor U9883 (N_9883,In_411,In_638);
xor U9884 (N_9884,In_119,In_2693);
xor U9885 (N_9885,In_1870,In_482);
or U9886 (N_9886,In_2934,In_527);
xor U9887 (N_9887,In_1951,In_1490);
and U9888 (N_9888,In_2030,In_2101);
xnor U9889 (N_9889,In_20,In_419);
or U9890 (N_9890,In_886,In_1693);
or U9891 (N_9891,In_782,In_192);
nor U9892 (N_9892,In_1931,In_1315);
nor U9893 (N_9893,In_1545,In_2675);
xnor U9894 (N_9894,In_2077,In_2121);
nor U9895 (N_9895,In_1005,In_54);
or U9896 (N_9896,In_2155,In_2873);
and U9897 (N_9897,In_2541,In_249);
nand U9898 (N_9898,In_788,In_453);
nand U9899 (N_9899,In_645,In_936);
xor U9900 (N_9900,In_66,In_1957);
nand U9901 (N_9901,In_2120,In_1389);
or U9902 (N_9902,In_2045,In_596);
and U9903 (N_9903,In_864,In_846);
nand U9904 (N_9904,In_2843,In_2827);
nor U9905 (N_9905,In_2047,In_2132);
nor U9906 (N_9906,In_1539,In_1258);
nand U9907 (N_9907,In_1000,In_2252);
xnor U9908 (N_9908,In_659,In_1539);
nor U9909 (N_9909,In_2186,In_2516);
and U9910 (N_9910,In_455,In_1637);
nor U9911 (N_9911,In_1397,In_445);
or U9912 (N_9912,In_2595,In_719);
or U9913 (N_9913,In_2314,In_1988);
and U9914 (N_9914,In_2254,In_2653);
xor U9915 (N_9915,In_395,In_2299);
xnor U9916 (N_9916,In_376,In_932);
or U9917 (N_9917,In_2051,In_2245);
nor U9918 (N_9918,In_1398,In_1067);
nor U9919 (N_9919,In_2433,In_1472);
nor U9920 (N_9920,In_38,In_1284);
or U9921 (N_9921,In_1815,In_87);
or U9922 (N_9922,In_937,In_1046);
and U9923 (N_9923,In_2326,In_2105);
xnor U9924 (N_9924,In_2913,In_2007);
or U9925 (N_9925,In_126,In_2438);
and U9926 (N_9926,In_2666,In_2942);
and U9927 (N_9927,In_1280,In_1954);
and U9928 (N_9928,In_1034,In_2932);
nand U9929 (N_9929,In_2940,In_624);
nor U9930 (N_9930,In_2951,In_2107);
or U9931 (N_9931,In_1310,In_1957);
and U9932 (N_9932,In_1490,In_795);
xor U9933 (N_9933,In_2664,In_1908);
nand U9934 (N_9934,In_1451,In_2048);
nor U9935 (N_9935,In_310,In_2108);
xnor U9936 (N_9936,In_501,In_2568);
or U9937 (N_9937,In_2483,In_1170);
xor U9938 (N_9938,In_195,In_10);
xor U9939 (N_9939,In_1475,In_409);
or U9940 (N_9940,In_2021,In_1270);
or U9941 (N_9941,In_16,In_1069);
xor U9942 (N_9942,In_1719,In_2523);
and U9943 (N_9943,In_1939,In_316);
nor U9944 (N_9944,In_525,In_2382);
nor U9945 (N_9945,In_1818,In_230);
xor U9946 (N_9946,In_1562,In_546);
and U9947 (N_9947,In_2736,In_1219);
or U9948 (N_9948,In_818,In_374);
nor U9949 (N_9949,In_1591,In_2942);
or U9950 (N_9950,In_2959,In_1894);
xor U9951 (N_9951,In_175,In_1736);
nand U9952 (N_9952,In_1147,In_797);
xor U9953 (N_9953,In_238,In_2054);
and U9954 (N_9954,In_2992,In_179);
nor U9955 (N_9955,In_2190,In_1022);
nand U9956 (N_9956,In_898,In_610);
nor U9957 (N_9957,In_1938,In_2271);
nand U9958 (N_9958,In_2318,In_1798);
or U9959 (N_9959,In_731,In_2991);
or U9960 (N_9960,In_1371,In_2462);
nor U9961 (N_9961,In_1767,In_2851);
and U9962 (N_9962,In_1861,In_77);
nor U9963 (N_9963,In_2357,In_502);
and U9964 (N_9964,In_248,In_852);
xnor U9965 (N_9965,In_2862,In_1025);
xnor U9966 (N_9966,In_354,In_1746);
nand U9967 (N_9967,In_726,In_1381);
and U9968 (N_9968,In_458,In_2646);
nand U9969 (N_9969,In_142,In_765);
nor U9970 (N_9970,In_2589,In_813);
nand U9971 (N_9971,In_2676,In_1937);
nor U9972 (N_9972,In_1473,In_2358);
xor U9973 (N_9973,In_1852,In_2720);
nand U9974 (N_9974,In_2629,In_2264);
nand U9975 (N_9975,In_516,In_595);
or U9976 (N_9976,In_1125,In_1746);
and U9977 (N_9977,In_1939,In_2454);
xnor U9978 (N_9978,In_2210,In_1859);
and U9979 (N_9979,In_1631,In_1686);
xor U9980 (N_9980,In_2301,In_127);
or U9981 (N_9981,In_2975,In_2896);
nor U9982 (N_9982,In_2349,In_1728);
xnor U9983 (N_9983,In_589,In_221);
nor U9984 (N_9984,In_1162,In_662);
or U9985 (N_9985,In_653,In_2843);
nor U9986 (N_9986,In_2941,In_502);
and U9987 (N_9987,In_2754,In_1486);
or U9988 (N_9988,In_2571,In_1139);
and U9989 (N_9989,In_1198,In_2426);
or U9990 (N_9990,In_2554,In_493);
xnor U9991 (N_9991,In_1244,In_1747);
xor U9992 (N_9992,In_2358,In_1960);
xor U9993 (N_9993,In_944,In_2620);
nand U9994 (N_9994,In_101,In_1995);
nand U9995 (N_9995,In_449,In_754);
and U9996 (N_9996,In_2582,In_189);
nand U9997 (N_9997,In_2522,In_805);
nor U9998 (N_9998,In_1508,In_2937);
or U9999 (N_9999,In_357,In_1204);
nor U10000 (N_10000,N_7674,N_7459);
xnor U10001 (N_10001,N_8042,N_2460);
nand U10002 (N_10002,N_3026,N_240);
and U10003 (N_10003,N_5238,N_395);
and U10004 (N_10004,N_1650,N_5897);
or U10005 (N_10005,N_4316,N_575);
and U10006 (N_10006,N_5075,N_6214);
xnor U10007 (N_10007,N_585,N_4737);
or U10008 (N_10008,N_9007,N_9060);
xor U10009 (N_10009,N_622,N_1453);
nand U10010 (N_10010,N_2060,N_1557);
nand U10011 (N_10011,N_1571,N_9679);
nand U10012 (N_10012,N_5470,N_4160);
xnor U10013 (N_10013,N_2188,N_6479);
xnor U10014 (N_10014,N_8364,N_9429);
or U10015 (N_10015,N_4104,N_9635);
xor U10016 (N_10016,N_6512,N_4391);
nor U10017 (N_10017,N_7873,N_3571);
xnor U10018 (N_10018,N_8781,N_3438);
nor U10019 (N_10019,N_3662,N_5375);
and U10020 (N_10020,N_3503,N_3291);
nand U10021 (N_10021,N_1320,N_2362);
nand U10022 (N_10022,N_8197,N_5262);
nor U10023 (N_10023,N_2861,N_6752);
nor U10024 (N_10024,N_4839,N_8107);
and U10025 (N_10025,N_5636,N_6806);
xnor U10026 (N_10026,N_4051,N_3371);
or U10027 (N_10027,N_9063,N_4220);
xor U10028 (N_10028,N_2465,N_426);
or U10029 (N_10029,N_6314,N_7988);
and U10030 (N_10030,N_1683,N_5842);
or U10031 (N_10031,N_9884,N_8847);
nand U10032 (N_10032,N_4854,N_2527);
or U10033 (N_10033,N_4058,N_6726);
nor U10034 (N_10034,N_9453,N_7448);
nor U10035 (N_10035,N_4233,N_4169);
nand U10036 (N_10036,N_9537,N_5824);
nand U10037 (N_10037,N_2835,N_7414);
nand U10038 (N_10038,N_7354,N_3017);
nand U10039 (N_10039,N_2241,N_4539);
xnor U10040 (N_10040,N_9921,N_3105);
or U10041 (N_10041,N_9685,N_651);
or U10042 (N_10042,N_4450,N_1166);
and U10043 (N_10043,N_4066,N_3648);
xnor U10044 (N_10044,N_785,N_6896);
xnor U10045 (N_10045,N_4670,N_8064);
or U10046 (N_10046,N_5409,N_1064);
nand U10047 (N_10047,N_4862,N_7052);
xnor U10048 (N_10048,N_1761,N_688);
and U10049 (N_10049,N_1212,N_889);
and U10050 (N_10050,N_7201,N_8973);
nand U10051 (N_10051,N_6995,N_9895);
nor U10052 (N_10052,N_9508,N_5372);
xnor U10053 (N_10053,N_9959,N_4208);
xor U10054 (N_10054,N_9006,N_4817);
or U10055 (N_10055,N_5102,N_77);
nand U10056 (N_10056,N_4632,N_758);
or U10057 (N_10057,N_8499,N_4088);
nand U10058 (N_10058,N_9170,N_9931);
nand U10059 (N_10059,N_7516,N_7018);
nor U10060 (N_10060,N_2350,N_7099);
xnor U10061 (N_10061,N_139,N_2099);
xnor U10062 (N_10062,N_9337,N_327);
or U10063 (N_10063,N_5421,N_1440);
xnor U10064 (N_10064,N_8520,N_7905);
and U10065 (N_10065,N_6059,N_9251);
nand U10066 (N_10066,N_4822,N_8626);
and U10067 (N_10067,N_2258,N_5632);
xor U10068 (N_10068,N_5302,N_248);
nor U10069 (N_10069,N_6268,N_6513);
or U10070 (N_10070,N_7687,N_8825);
or U10071 (N_10071,N_5362,N_254);
nor U10072 (N_10072,N_6568,N_8126);
nor U10073 (N_10073,N_5807,N_8482);
and U10074 (N_10074,N_5290,N_5250);
and U10075 (N_10075,N_6309,N_769);
nor U10076 (N_10076,N_9820,N_7998);
nor U10077 (N_10077,N_6390,N_5206);
and U10078 (N_10078,N_4376,N_9521);
nand U10079 (N_10079,N_4942,N_8136);
xor U10080 (N_10080,N_543,N_3252);
and U10081 (N_10081,N_6516,N_9497);
and U10082 (N_10082,N_1014,N_3716);
or U10083 (N_10083,N_1110,N_4431);
nor U10084 (N_10084,N_2256,N_9943);
xnor U10085 (N_10085,N_5571,N_8600);
and U10086 (N_10086,N_906,N_8308);
nand U10087 (N_10087,N_1396,N_7999);
xnor U10088 (N_10088,N_3844,N_9257);
xor U10089 (N_10089,N_8264,N_7779);
nor U10090 (N_10090,N_2776,N_6315);
or U10091 (N_10091,N_2616,N_2247);
nor U10092 (N_10092,N_279,N_6637);
nor U10093 (N_10093,N_7635,N_918);
or U10094 (N_10094,N_8791,N_8217);
nand U10095 (N_10095,N_5770,N_9038);
nor U10096 (N_10096,N_7663,N_3737);
or U10097 (N_10097,N_4366,N_6760);
or U10098 (N_10098,N_8530,N_4706);
and U10099 (N_10099,N_4045,N_6118);
nand U10100 (N_10100,N_6798,N_4341);
xor U10101 (N_10101,N_868,N_604);
nor U10102 (N_10102,N_9054,N_8869);
or U10103 (N_10103,N_9712,N_8398);
xor U10104 (N_10104,N_8278,N_6438);
xor U10105 (N_10105,N_6997,N_5847);
xnor U10106 (N_10106,N_9799,N_7402);
and U10107 (N_10107,N_3050,N_8204);
and U10108 (N_10108,N_8045,N_6410);
xnor U10109 (N_10109,N_5467,N_7318);
nand U10110 (N_10110,N_2212,N_1191);
xnor U10111 (N_10111,N_2988,N_3866);
nor U10112 (N_10112,N_4318,N_7132);
or U10113 (N_10113,N_4148,N_7050);
xor U10114 (N_10114,N_530,N_1519);
nand U10115 (N_10115,N_8811,N_1403);
nand U10116 (N_10116,N_4353,N_9215);
xnor U10117 (N_10117,N_4768,N_1776);
nor U10118 (N_10118,N_9912,N_4917);
nor U10119 (N_10119,N_8258,N_8368);
or U10120 (N_10120,N_1102,N_1463);
and U10121 (N_10121,N_2232,N_5772);
or U10122 (N_10122,N_5753,N_250);
or U10123 (N_10123,N_3037,N_4820);
nand U10124 (N_10124,N_9440,N_4396);
and U10125 (N_10125,N_7956,N_8070);
or U10126 (N_10126,N_3847,N_5221);
xor U10127 (N_10127,N_5501,N_2504);
and U10128 (N_10128,N_82,N_3413);
and U10129 (N_10129,N_3606,N_6199);
nand U10130 (N_10130,N_8420,N_4360);
and U10131 (N_10131,N_7966,N_3135);
and U10132 (N_10132,N_8319,N_1871);
and U10133 (N_10133,N_3172,N_2984);
and U10134 (N_10134,N_826,N_1408);
xnor U10135 (N_10135,N_2733,N_338);
nor U10136 (N_10136,N_7176,N_9082);
nand U10137 (N_10137,N_4134,N_2868);
nor U10138 (N_10138,N_315,N_5420);
or U10139 (N_10139,N_9330,N_1714);
nand U10140 (N_10140,N_2595,N_4935);
xnor U10141 (N_10141,N_2481,N_1298);
nand U10142 (N_10142,N_217,N_1036);
or U10143 (N_10143,N_4807,N_2449);
xnor U10144 (N_10144,N_2712,N_5435);
nor U10145 (N_10145,N_8215,N_5241);
or U10146 (N_10146,N_4921,N_2630);
nand U10147 (N_10147,N_546,N_7748);
xor U10148 (N_10148,N_8524,N_1919);
and U10149 (N_10149,N_2205,N_2730);
xor U10150 (N_10150,N_5949,N_3048);
or U10151 (N_10151,N_5245,N_7825);
nor U10152 (N_10152,N_3241,N_3043);
xnor U10153 (N_10153,N_1973,N_3346);
nand U10154 (N_10154,N_2574,N_8535);
xor U10155 (N_10155,N_2822,N_8369);
xnor U10156 (N_10156,N_5861,N_1658);
xor U10157 (N_10157,N_6478,N_596);
nand U10158 (N_10158,N_3286,N_1295);
and U10159 (N_10159,N_505,N_4122);
and U10160 (N_10160,N_155,N_7338);
or U10161 (N_10161,N_8519,N_7688);
xor U10162 (N_10162,N_8479,N_5103);
nor U10163 (N_10163,N_5017,N_1262);
xor U10164 (N_10164,N_5355,N_6946);
nor U10165 (N_10165,N_7276,N_6952);
nor U10166 (N_10166,N_3708,N_2934);
and U10167 (N_10167,N_8248,N_2214);
and U10168 (N_10168,N_6832,N_6860);
and U10169 (N_10169,N_2736,N_9377);
nor U10170 (N_10170,N_4269,N_9648);
and U10171 (N_10171,N_9896,N_9136);
or U10172 (N_10172,N_888,N_537);
and U10173 (N_10173,N_2443,N_4200);
nand U10174 (N_10174,N_3790,N_9660);
nand U10175 (N_10175,N_5611,N_3741);
nand U10176 (N_10176,N_911,N_2825);
nor U10177 (N_10177,N_6652,N_7352);
and U10178 (N_10178,N_3168,N_2727);
or U10179 (N_10179,N_9653,N_3430);
nand U10180 (N_10180,N_6456,N_6912);
or U10181 (N_10181,N_2851,N_1428);
nand U10182 (N_10182,N_3106,N_4146);
or U10183 (N_10183,N_1775,N_8669);
nand U10184 (N_10184,N_799,N_9318);
or U10185 (N_10185,N_5783,N_3303);
or U10186 (N_10186,N_2220,N_1265);
or U10187 (N_10187,N_2440,N_5809);
and U10188 (N_10188,N_9162,N_7003);
nor U10189 (N_10189,N_7574,N_8906);
and U10190 (N_10190,N_8988,N_1653);
xnor U10191 (N_10191,N_9425,N_3659);
nand U10192 (N_10192,N_5363,N_9245);
and U10193 (N_10193,N_5061,N_4830);
xnor U10194 (N_10194,N_7932,N_3549);
or U10195 (N_10195,N_4941,N_3758);
xnor U10196 (N_10196,N_3851,N_1046);
xnor U10197 (N_10197,N_638,N_6228);
nor U10198 (N_10198,N_1599,N_325);
or U10199 (N_10199,N_3014,N_8174);
nand U10200 (N_10200,N_3693,N_539);
or U10201 (N_10201,N_5558,N_2287);
or U10202 (N_10202,N_7800,N_7009);
and U10203 (N_10203,N_8773,N_2137);
or U10204 (N_10204,N_1097,N_4455);
nor U10205 (N_10205,N_7157,N_6854);
and U10206 (N_10206,N_2140,N_4863);
nor U10207 (N_10207,N_7639,N_6712);
xor U10208 (N_10208,N_9841,N_3518);
xor U10209 (N_10209,N_9225,N_2933);
or U10210 (N_10210,N_4782,N_145);
and U10211 (N_10211,N_8780,N_5835);
nand U10212 (N_10212,N_8028,N_1192);
nand U10213 (N_10213,N_4462,N_2124);
or U10214 (N_10214,N_3517,N_3931);
or U10215 (N_10215,N_183,N_6258);
or U10216 (N_10216,N_7922,N_9247);
xor U10217 (N_10217,N_1502,N_4998);
nor U10218 (N_10218,N_6471,N_5802);
nor U10219 (N_10219,N_8106,N_329);
xnor U10220 (N_10220,N_9471,N_6098);
nand U10221 (N_10221,N_9879,N_3062);
and U10222 (N_10222,N_5354,N_6669);
nor U10223 (N_10223,N_965,N_8382);
or U10224 (N_10224,N_5993,N_9831);
xor U10225 (N_10225,N_6373,N_9058);
or U10226 (N_10226,N_5500,N_6274);
or U10227 (N_10227,N_9370,N_4522);
xor U10228 (N_10228,N_6633,N_3437);
nor U10229 (N_10229,N_8843,N_2773);
nand U10230 (N_10230,N_7357,N_1790);
xnor U10231 (N_10231,N_4657,N_745);
or U10232 (N_10232,N_5198,N_2697);
nand U10233 (N_10233,N_6034,N_7707);
and U10234 (N_10234,N_3032,N_2589);
or U10235 (N_10235,N_3242,N_5249);
nand U10236 (N_10236,N_7026,N_1524);
nor U10237 (N_10237,N_1032,N_5064);
and U10238 (N_10238,N_1665,N_1030);
or U10239 (N_10239,N_5097,N_2715);
nor U10240 (N_10240,N_5635,N_4627);
nand U10241 (N_10241,N_9511,N_3663);
nor U10242 (N_10242,N_1578,N_2237);
nand U10243 (N_10243,N_9115,N_569);
xnor U10244 (N_10244,N_3140,N_9017);
xor U10245 (N_10245,N_4166,N_620);
nand U10246 (N_10246,N_5644,N_616);
xor U10247 (N_10247,N_1731,N_729);
or U10248 (N_10248,N_9837,N_9238);
and U10249 (N_10249,N_4060,N_87);
nor U10250 (N_10250,N_3743,N_2159);
and U10251 (N_10251,N_1646,N_6823);
nand U10252 (N_10252,N_1783,N_3886);
nand U10253 (N_10253,N_1503,N_7085);
nand U10254 (N_10254,N_427,N_1535);
xor U10255 (N_10255,N_7416,N_2548);
nor U10256 (N_10256,N_8889,N_4403);
nand U10257 (N_10257,N_9674,N_9042);
xnor U10258 (N_10258,N_4140,N_7185);
nor U10259 (N_10259,N_2898,N_6142);
nand U10260 (N_10260,N_9433,N_3519);
nor U10261 (N_10261,N_460,N_6886);
nor U10262 (N_10262,N_8567,N_5675);
or U10263 (N_10263,N_4000,N_4413);
nand U10264 (N_10264,N_8576,N_6922);
nand U10265 (N_10265,N_7440,N_1623);
and U10266 (N_10266,N_439,N_764);
nand U10267 (N_10267,N_5920,N_9600);
and U10268 (N_10268,N_360,N_1918);
nor U10269 (N_10269,N_878,N_9675);
and U10270 (N_10270,N_6959,N_603);
or U10271 (N_10271,N_9980,N_926);
nand U10272 (N_10272,N_4779,N_8166);
nand U10273 (N_10273,N_2959,N_8181);
xor U10274 (N_10274,N_3419,N_3640);
nand U10275 (N_10275,N_9978,N_8465);
xnor U10276 (N_10276,N_1442,N_4372);
nand U10277 (N_10277,N_7846,N_4042);
nand U10278 (N_10278,N_1936,N_268);
or U10279 (N_10279,N_4488,N_4944);
nand U10280 (N_10280,N_4037,N_3853);
or U10281 (N_10281,N_4349,N_4020);
nand U10282 (N_10282,N_4723,N_1544);
nand U10283 (N_10283,N_2410,N_2052);
and U10284 (N_10284,N_3927,N_6105);
xnor U10285 (N_10285,N_8110,N_9767);
nand U10286 (N_10286,N_6193,N_3442);
and U10287 (N_10287,N_3725,N_2117);
nand U10288 (N_10288,N_2412,N_847);
xnor U10289 (N_10289,N_5337,N_9088);
nor U10290 (N_10290,N_8097,N_2142);
and U10291 (N_10291,N_2725,N_9725);
xnor U10292 (N_10292,N_9644,N_5525);
nor U10293 (N_10293,N_9560,N_4019);
xnor U10294 (N_10294,N_5565,N_9081);
and U10295 (N_10295,N_5074,N_1476);
xor U10296 (N_10296,N_7705,N_347);
or U10297 (N_10297,N_1318,N_7807);
and U10298 (N_10298,N_3781,N_1848);
and U10299 (N_10299,N_3586,N_7521);
xor U10300 (N_10300,N_2732,N_1205);
or U10301 (N_10301,N_8975,N_6723);
nor U10302 (N_10302,N_3918,N_2197);
xor U10303 (N_10303,N_2301,N_3592);
xnor U10304 (N_10304,N_2886,N_9923);
nand U10305 (N_10305,N_2797,N_6562);
xor U10306 (N_10306,N_1134,N_6665);
xnor U10307 (N_10307,N_9311,N_5101);
and U10308 (N_10308,N_3331,N_2321);
nand U10309 (N_10309,N_1685,N_4999);
and U10310 (N_10310,N_8014,N_2871);
and U10311 (N_10311,N_2585,N_7245);
and U10312 (N_10312,N_3087,N_3138);
nand U10313 (N_10313,N_6650,N_5788);
or U10314 (N_10314,N_6819,N_2633);
xor U10315 (N_10315,N_1841,N_5596);
and U10316 (N_10316,N_8970,N_1123);
xor U10317 (N_10317,N_6060,N_6302);
or U10318 (N_10318,N_4302,N_9072);
and U10319 (N_10319,N_2050,N_1662);
xnor U10320 (N_10320,N_7005,N_4725);
nand U10321 (N_10321,N_5356,N_6006);
nand U10322 (N_10322,N_1632,N_6631);
or U10323 (N_10323,N_4911,N_349);
nand U10324 (N_10324,N_6826,N_2593);
and U10325 (N_10325,N_1169,N_401);
and U10326 (N_10326,N_8820,N_1126);
nor U10327 (N_10327,N_6674,N_6024);
nor U10328 (N_10328,N_3469,N_2759);
and U10329 (N_10329,N_1415,N_528);
xor U10330 (N_10330,N_7817,N_3131);
nor U10331 (N_10331,N_8818,N_8299);
nor U10332 (N_10332,N_5059,N_235);
xnor U10333 (N_10333,N_5643,N_2354);
or U10334 (N_10334,N_7739,N_6559);
or U10335 (N_10335,N_495,N_7889);
nand U10336 (N_10336,N_5982,N_3669);
nand U10337 (N_10337,N_4738,N_3505);
nor U10338 (N_10338,N_7415,N_3121);
xor U10339 (N_10339,N_6550,N_4966);
and U10340 (N_10340,N_7827,N_9048);
nand U10341 (N_10341,N_1344,N_5175);
and U10342 (N_10342,N_400,N_425);
nor U10343 (N_10343,N_3879,N_5285);
xnor U10344 (N_10344,N_4116,N_4115);
and U10345 (N_10345,N_7378,N_6040);
nand U10346 (N_10346,N_8372,N_6709);
nand U10347 (N_10347,N_3902,N_303);
xnor U10348 (N_10348,N_9845,N_357);
and U10349 (N_10349,N_5167,N_177);
nor U10350 (N_10350,N_7881,N_1617);
nand U10351 (N_10351,N_9632,N_378);
xnor U10352 (N_10352,N_3095,N_1361);
or U10353 (N_10353,N_2459,N_655);
and U10354 (N_10354,N_3223,N_4456);
xor U10355 (N_10355,N_405,N_6621);
nor U10356 (N_10356,N_756,N_4305);
nand U10357 (N_10357,N_7594,N_9129);
nor U10358 (N_10358,N_3694,N_7493);
or U10359 (N_10359,N_6519,N_940);
or U10360 (N_10360,N_60,N_9045);
xnor U10361 (N_10361,N_4608,N_992);
nand U10362 (N_10362,N_2468,N_6226);
nor U10363 (N_10363,N_5845,N_5545);
or U10364 (N_10364,N_7148,N_7504);
nor U10365 (N_10365,N_9652,N_7184);
and U10366 (N_10366,N_9785,N_853);
nor U10367 (N_10367,N_3072,N_7653);
nor U10368 (N_10368,N_3178,N_5553);
xor U10369 (N_10369,N_4300,N_8610);
or U10370 (N_10370,N_5322,N_831);
nor U10371 (N_10371,N_6965,N_3219);
xnor U10372 (N_10372,N_4016,N_2857);
nor U10373 (N_10373,N_6173,N_6615);
xnor U10374 (N_10374,N_1937,N_3246);
and U10375 (N_10375,N_7231,N_387);
nand U10376 (N_10376,N_4384,N_4358);
xnor U10377 (N_10377,N_3093,N_7279);
nor U10378 (N_10378,N_2512,N_8884);
nor U10379 (N_10379,N_1928,N_753);
xor U10380 (N_10380,N_7063,N_5287);
nor U10381 (N_10381,N_6042,N_8060);
nor U10382 (N_10382,N_1855,N_557);
nor U10383 (N_10383,N_635,N_952);
and U10384 (N_10384,N_4479,N_2338);
xor U10385 (N_10385,N_2671,N_8370);
xnor U10386 (N_10386,N_2767,N_7427);
or U10387 (N_10387,N_1000,N_6945);
nand U10388 (N_10388,N_2516,N_5577);
nand U10389 (N_10389,N_4809,N_6257);
or U10390 (N_10390,N_3320,N_9645);
xor U10391 (N_10391,N_9727,N_365);
nor U10392 (N_10392,N_8742,N_9207);
and U10393 (N_10393,N_4713,N_3221);
and U10394 (N_10394,N_4348,N_7893);
or U10395 (N_10395,N_9463,N_2058);
or U10396 (N_10396,N_6841,N_8763);
xnor U10397 (N_10397,N_4252,N_5471);
xor U10398 (N_10398,N_7668,N_4765);
xor U10399 (N_10399,N_7866,N_5006);
nand U10400 (N_10400,N_8565,N_6102);
nor U10401 (N_10401,N_8671,N_8296);
nor U10402 (N_10402,N_9360,N_8102);
nand U10403 (N_10403,N_7820,N_801);
nor U10404 (N_10404,N_5342,N_9084);
xor U10405 (N_10405,N_2742,N_1300);
and U10406 (N_10406,N_7951,N_278);
nand U10407 (N_10407,N_3577,N_2351);
nor U10408 (N_10408,N_6644,N_9441);
or U10409 (N_10409,N_4852,N_9589);
xnor U10410 (N_10410,N_4621,N_9539);
or U10411 (N_10411,N_5416,N_4028);
and U10412 (N_10412,N_4730,N_512);
nor U10413 (N_10413,N_3158,N_2919);
and U10414 (N_10414,N_7780,N_8597);
xnor U10415 (N_10415,N_1523,N_9176);
xor U10416 (N_10416,N_2384,N_6140);
nand U10417 (N_10417,N_1121,N_9774);
nor U10418 (N_10418,N_483,N_4549);
nand U10419 (N_10419,N_2326,N_5508);
xor U10420 (N_10420,N_75,N_3588);
xor U10421 (N_10421,N_9741,N_5091);
nor U10422 (N_10422,N_9812,N_6321);
nand U10423 (N_10423,N_4218,N_4010);
nor U10424 (N_10424,N_8427,N_7614);
and U10425 (N_10425,N_3159,N_9814);
or U10426 (N_10426,N_1712,N_5374);
nand U10427 (N_10427,N_2790,N_8901);
nand U10428 (N_10428,N_4271,N_4119);
or U10429 (N_10429,N_9480,N_4990);
nor U10430 (N_10430,N_9705,N_3333);
nor U10431 (N_10431,N_3933,N_2833);
and U10432 (N_10432,N_3324,N_7204);
nand U10433 (N_10433,N_469,N_9783);
nor U10434 (N_10434,N_9313,N_4424);
or U10435 (N_10435,N_1616,N_8409);
nand U10436 (N_10436,N_3650,N_1324);
or U10437 (N_10437,N_7172,N_5656);
nand U10438 (N_10438,N_659,N_2128);
xnor U10439 (N_10439,N_6463,N_98);
nor U10440 (N_10440,N_5233,N_8173);
and U10441 (N_10441,N_7559,N_1387);
or U10442 (N_10442,N_2122,N_5036);
and U10443 (N_10443,N_8358,N_8155);
nor U10444 (N_10444,N_6523,N_5978);
or U10445 (N_10445,N_6235,N_3373);
and U10446 (N_10446,N_6980,N_4049);
and U10447 (N_10447,N_2969,N_1496);
or U10448 (N_10448,N_7535,N_8048);
xnor U10449 (N_10449,N_9570,N_833);
xor U10450 (N_10450,N_4150,N_4663);
nor U10451 (N_10451,N_9466,N_5505);
nor U10452 (N_10452,N_802,N_507);
nor U10453 (N_10453,N_5434,N_4865);
and U10454 (N_10454,N_6211,N_1574);
and U10455 (N_10455,N_4943,N_4147);
or U10456 (N_10456,N_8084,N_2612);
nand U10457 (N_10457,N_2908,N_4856);
nand U10458 (N_10458,N_658,N_6973);
or U10459 (N_10459,N_9158,N_3778);
xnor U10460 (N_10460,N_8668,N_6785);
and U10461 (N_10461,N_4317,N_3185);
and U10462 (N_10462,N_6987,N_5210);
nor U10463 (N_10463,N_1129,N_9066);
nand U10464 (N_10464,N_6927,N_4013);
nor U10465 (N_10465,N_3712,N_2261);
and U10466 (N_10466,N_2300,N_2881);
nand U10467 (N_10467,N_3965,N_6490);
xnor U10468 (N_10468,N_9264,N_1067);
xnor U10469 (N_10469,N_6192,N_725);
or U10470 (N_10470,N_3770,N_4986);
nor U10471 (N_10471,N_5584,N_9011);
xor U10472 (N_10472,N_8253,N_982);
xnor U10473 (N_10473,N_4778,N_1314);
and U10474 (N_10474,N_5874,N_5089);
or U10475 (N_10475,N_1782,N_4715);
or U10476 (N_10476,N_2274,N_9346);
and U10477 (N_10477,N_6573,N_5479);
nand U10478 (N_10478,N_1537,N_2450);
nor U10479 (N_10479,N_8690,N_2796);
and U10480 (N_10480,N_2346,N_2550);
nor U10481 (N_10481,N_9714,N_2694);
nand U10482 (N_10482,N_6285,N_2946);
and U10483 (N_10483,N_9324,N_1719);
nand U10484 (N_10484,N_7896,N_6700);
nand U10485 (N_10485,N_3354,N_4410);
and U10486 (N_10486,N_6080,N_3937);
nand U10487 (N_10487,N_8683,N_5157);
and U10488 (N_10488,N_549,N_938);
xor U10489 (N_10489,N_404,N_1017);
xor U10490 (N_10490,N_8114,N_7280);
and U10491 (N_10491,N_8870,N_6452);
and U10492 (N_10492,N_6857,N_1518);
or U10493 (N_10493,N_9854,N_8919);
and U10494 (N_10494,N_3019,N_2523);
nor U10495 (N_10495,N_7702,N_3739);
nand U10496 (N_10496,N_7164,N_3114);
xor U10497 (N_10497,N_8283,N_164);
nand U10498 (N_10498,N_991,N_630);
and U10499 (N_10499,N_7979,N_7666);
nand U10500 (N_10500,N_8207,N_3245);
or U10501 (N_10501,N_1267,N_8609);
xor U10502 (N_10502,N_4240,N_2187);
xor U10503 (N_10503,N_3506,N_4833);
nand U10504 (N_10504,N_1155,N_815);
nand U10505 (N_10505,N_2850,N_6205);
nor U10506 (N_10506,N_9743,N_6430);
nor U10507 (N_10507,N_8738,N_470);
or U10508 (N_10508,N_7523,N_7657);
xnor U10509 (N_10509,N_3885,N_3192);
xnor U10510 (N_10510,N_4421,N_7370);
nor U10511 (N_10511,N_6457,N_1236);
xor U10512 (N_10512,N_9413,N_6141);
or U10513 (N_10513,N_66,N_8801);
and U10514 (N_10514,N_7710,N_7806);
nand U10515 (N_10515,N_5070,N_5647);
nand U10516 (N_10516,N_7275,N_8834);
nand U10517 (N_10517,N_1629,N_4155);
nor U10518 (N_10518,N_3594,N_397);
or U10519 (N_10519,N_9780,N_8375);
nor U10520 (N_10520,N_5131,N_6347);
nand U10521 (N_10521,N_2763,N_9860);
nand U10522 (N_10522,N_9593,N_5489);
xor U10523 (N_10523,N_1716,N_5696);
xor U10524 (N_10524,N_7061,N_8685);
nor U10525 (N_10525,N_8894,N_4864);
nor U10526 (N_10526,N_7233,N_2386);
nor U10527 (N_10527,N_957,N_4620);
nand U10528 (N_10528,N_8552,N_8031);
and U10529 (N_10529,N_5922,N_997);
nor U10530 (N_10530,N_2655,N_124);
xnor U10531 (N_10531,N_5276,N_6326);
xnor U10532 (N_10532,N_9828,N_9694);
xnor U10533 (N_10533,N_9667,N_5455);
xnor U10534 (N_10534,N_5575,N_5130);
nand U10535 (N_10535,N_1509,N_7088);
and U10536 (N_10536,N_1770,N_6587);
and U10537 (N_10537,N_1058,N_9962);
xnor U10538 (N_10538,N_6009,N_1119);
nand U10539 (N_10539,N_1373,N_1901);
or U10540 (N_10540,N_4468,N_9216);
and U10541 (N_10541,N_8282,N_6354);
or U10542 (N_10542,N_4340,N_6203);
and U10543 (N_10543,N_1799,N_6108);
xor U10544 (N_10544,N_6379,N_1418);
nor U10545 (N_10545,N_7685,N_1293);
nor U10546 (N_10546,N_9187,N_3022);
or U10547 (N_10547,N_4562,N_9716);
nand U10548 (N_10548,N_9367,N_2364);
nand U10549 (N_10549,N_9052,N_9760);
xnor U10550 (N_10550,N_4368,N_2458);
xor U10551 (N_10551,N_6520,N_5943);
and U10552 (N_10552,N_8508,N_1642);
nor U10553 (N_10553,N_9108,N_8703);
nand U10554 (N_10554,N_590,N_7718);
and U10555 (N_10555,N_4326,N_9513);
nor U10556 (N_10556,N_1831,N_5811);
and U10557 (N_10557,N_7126,N_817);
and U10558 (N_10558,N_9899,N_2359);
xor U10559 (N_10559,N_383,N_810);
or U10560 (N_10560,N_6915,N_2577);
or U10561 (N_10561,N_3280,N_8717);
or U10562 (N_10562,N_8624,N_3007);
nor U10563 (N_10563,N_3583,N_457);
and U10564 (N_10564,N_5723,N_7105);
nand U10565 (N_10565,N_3476,N_8035);
xnor U10566 (N_10566,N_6646,N_7189);
nand U10567 (N_10567,N_6605,N_2030);
nor U10568 (N_10568,N_5825,N_6779);
and U10569 (N_10569,N_8677,N_4185);
or U10570 (N_10570,N_7805,N_3490);
nand U10571 (N_10571,N_3426,N_3336);
or U10572 (N_10572,N_1638,N_3630);
nor U10573 (N_10573,N_930,N_3624);
nor U10574 (N_10574,N_227,N_9973);
nand U10575 (N_10575,N_5660,N_1281);
xor U10576 (N_10576,N_9979,N_3416);
nor U10577 (N_10577,N_2924,N_8183);
nand U10578 (N_10578,N_6135,N_4286);
or U10579 (N_10579,N_8252,N_5775);
nand U10580 (N_10580,N_5078,N_9435);
xor U10581 (N_10581,N_4527,N_6744);
or U10582 (N_10582,N_1215,N_525);
xor U10583 (N_10583,N_5963,N_277);
xnor U10584 (N_10584,N_6904,N_1147);
and U10585 (N_10585,N_5286,N_3963);
nand U10586 (N_10586,N_2786,N_8905);
xor U10587 (N_10587,N_8182,N_5555);
and U10588 (N_10588,N_3309,N_2744);
nor U10589 (N_10589,N_2087,N_4596);
or U10590 (N_10590,N_5578,N_5358);
and U10591 (N_10591,N_9246,N_3243);
xnor U10592 (N_10592,N_1633,N_2662);
and U10593 (N_10593,N_3104,N_6642);
or U10594 (N_10594,N_2620,N_1494);
nand U10595 (N_10595,N_5303,N_2615);
and U10596 (N_10596,N_2150,N_3433);
and U10597 (N_10597,N_566,N_8396);
and U10598 (N_10598,N_195,N_6783);
xor U10599 (N_10599,N_3389,N_2526);
nand U10600 (N_10600,N_2395,N_923);
and U10601 (N_10601,N_513,N_4573);
and U10602 (N_10602,N_5365,N_9911);
nor U10603 (N_10603,N_4581,N_9878);
xor U10604 (N_10604,N_5832,N_9152);
nor U10605 (N_10605,N_8450,N_707);
xnor U10606 (N_10606,N_5773,N_2324);
and U10607 (N_10607,N_7057,N_9900);
or U10608 (N_10608,N_1596,N_324);
xor U10609 (N_10609,N_9277,N_4594);
nor U10610 (N_10610,N_9558,N_6038);
and U10611 (N_10611,N_4988,N_12);
or U10612 (N_10612,N_6816,N_1459);
xnor U10613 (N_10613,N_450,N_1047);
or U10614 (N_10614,N_7781,N_9597);
nor U10615 (N_10615,N_6998,N_7065);
nand U10616 (N_10616,N_4477,N_4975);
or U10617 (N_10617,N_4261,N_4676);
or U10618 (N_10618,N_9771,N_6620);
xor U10619 (N_10619,N_1213,N_3360);
nand U10620 (N_10620,N_3302,N_7092);
and U10621 (N_10621,N_5349,N_5009);
and U10622 (N_10622,N_9203,N_7048);
nand U10623 (N_10623,N_8900,N_2545);
and U10624 (N_10624,N_2101,N_2841);
nor U10625 (N_10625,N_4823,N_5899);
and U10626 (N_10626,N_8627,N_5726);
and U10627 (N_10627,N_193,N_1306);
xor U10628 (N_10628,N_9886,N_5714);
xnor U10629 (N_10629,N_1343,N_3784);
nor U10630 (N_10630,N_8904,N_9398);
xor U10631 (N_10631,N_9278,N_9350);
xnor U10632 (N_10632,N_1707,N_9954);
and U10633 (N_10633,N_5697,N_1028);
nor U10634 (N_10634,N_2992,N_5684);
nand U10635 (N_10635,N_4236,N_4542);
nor U10636 (N_10636,N_5418,N_6951);
or U10637 (N_10637,N_581,N_6544);
nor U10638 (N_10638,N_9120,N_9706);
nand U10639 (N_10639,N_6840,N_7071);
xor U10640 (N_10640,N_1885,N_2906);
nand U10641 (N_10641,N_1887,N_4469);
nor U10642 (N_10642,N_4536,N_3388);
and U10643 (N_10643,N_9499,N_1217);
xor U10644 (N_10644,N_6966,N_5984);
nand U10645 (N_10645,N_8598,N_8436);
nand U10646 (N_10646,N_5977,N_6176);
nand U10647 (N_10647,N_5626,N_5995);
nand U10648 (N_10648,N_9454,N_9975);
or U10649 (N_10649,N_8122,N_8859);
nor U10650 (N_10650,N_8865,N_2675);
and U10651 (N_10651,N_1128,N_2086);
and U10652 (N_10652,N_748,N_678);
nand U10653 (N_10653,N_4215,N_7539);
or U10654 (N_10654,N_7973,N_8458);
nor U10655 (N_10655,N_550,N_2867);
xnor U10656 (N_10656,N_8327,N_3316);
and U10657 (N_10657,N_8490,N_318);
nand U10658 (N_10658,N_111,N_5678);
nand U10659 (N_10659,N_1150,N_1567);
or U10660 (N_10660,N_7310,N_3710);
and U10661 (N_10661,N_796,N_7424);
and U10662 (N_10662,N_4685,N_2441);
xor U10663 (N_10663,N_5251,N_7302);
nand U10664 (N_10664,N_1462,N_3152);
or U10665 (N_10665,N_3189,N_3423);
nor U10666 (N_10666,N_446,N_7226);
and U10667 (N_10667,N_3378,N_1194);
and U10668 (N_10668,N_4766,N_376);
and U10669 (N_10669,N_5925,N_7242);
nor U10670 (N_10670,N_3231,N_628);
nand U10671 (N_10671,N_203,N_2471);
or U10672 (N_10672,N_3567,N_5954);
nand U10673 (N_10673,N_2446,N_2889);
nand U10674 (N_10674,N_7968,N_5084);
or U10675 (N_10675,N_4915,N_3209);
xnor U10676 (N_10676,N_5542,N_6749);
or U10677 (N_10677,N_136,N_4309);
nand U10678 (N_10678,N_3734,N_5702);
nor U10679 (N_10679,N_4953,N_7485);
xnor U10680 (N_10680,N_8157,N_104);
and U10681 (N_10681,N_1362,N_8062);
xnor U10682 (N_10682,N_8313,N_4081);
and U10683 (N_10683,N_7696,N_8251);
or U10684 (N_10684,N_4069,N_9617);
or U10685 (N_10685,N_5243,N_3085);
or U10686 (N_10686,N_5520,N_1363);
nand U10687 (N_10687,N_4630,N_9684);
nor U10688 (N_10688,N_9477,N_9897);
xnor U10689 (N_10689,N_5368,N_6893);
xnor U10690 (N_10690,N_2454,N_1700);
or U10691 (N_10691,N_6133,N_4755);
or U10692 (N_10692,N_1814,N_461);
nor U10693 (N_10693,N_3480,N_2784);
nor U10694 (N_10694,N_3895,N_8057);
or U10695 (N_10695,N_4913,N_9117);
and U10696 (N_10696,N_9728,N_366);
nor U10697 (N_10697,N_4775,N_3552);
xnor U10698 (N_10698,N_5460,N_908);
nor U10699 (N_10699,N_5361,N_9003);
xor U10700 (N_10700,N_2007,N_9121);
or U10701 (N_10701,N_776,N_5895);
nor U10702 (N_10702,N_9012,N_2093);
xor U10703 (N_10703,N_1709,N_8815);
xnor U10704 (N_10704,N_2913,N_3560);
xnor U10705 (N_10705,N_3939,N_7845);
nand U10706 (N_10706,N_969,N_7002);
nor U10707 (N_10707,N_8116,N_2996);
nand U10708 (N_10708,N_2439,N_8964);
and U10709 (N_10709,N_1961,N_3464);
nor U10710 (N_10710,N_6685,N_1520);
nand U10711 (N_10711,N_4687,N_168);
nor U10712 (N_10712,N_6150,N_4306);
or U10713 (N_10713,N_6172,N_3250);
nand U10714 (N_10714,N_9101,N_7910);
nand U10715 (N_10715,N_7054,N_9388);
nand U10716 (N_10716,N_3041,N_7384);
and U10717 (N_10717,N_4009,N_7471);
nand U10718 (N_10718,N_9307,N_9185);
nor U10719 (N_10719,N_6282,N_6994);
or U10720 (N_10720,N_7359,N_9059);
and U10721 (N_10721,N_7439,N_3133);
xor U10722 (N_10722,N_8534,N_7100);
nand U10723 (N_10723,N_531,N_3634);
and U10724 (N_10724,N_7170,N_4736);
xnor U10725 (N_10725,N_3768,N_5708);
and U10726 (N_10726,N_4282,N_876);
or U10727 (N_10727,N_5352,N_2332);
xnor U10728 (N_10728,N_7266,N_7209);
nand U10729 (N_10729,N_6195,N_8410);
xnor U10730 (N_10730,N_4142,N_3239);
xor U10731 (N_10731,N_5923,N_4297);
nor U10732 (N_10732,N_7714,N_2021);
nor U10733 (N_10733,N_2936,N_2228);
xnor U10734 (N_10734,N_180,N_6788);
xnor U10735 (N_10735,N_8945,N_8958);
xor U10736 (N_10736,N_6267,N_131);
or U10737 (N_10737,N_9719,N_2613);
nor U10738 (N_10738,N_4031,N_7970);
or U10739 (N_10739,N_3115,N_820);
xnor U10740 (N_10740,N_451,N_6567);
nand U10741 (N_10741,N_5369,N_7325);
and U10742 (N_10742,N_3574,N_8751);
nand U10743 (N_10743,N_3791,N_6164);
nand U10744 (N_10744,N_1890,N_6773);
nand U10745 (N_10745,N_2765,N_6557);
xnor U10746 (N_10746,N_5573,N_4654);
xnor U10747 (N_10747,N_7802,N_9288);
xor U10748 (N_10748,N_8216,N_4065);
xor U10749 (N_10749,N_2792,N_594);
and U10750 (N_10750,N_3646,N_4507);
xor U10751 (N_10751,N_8577,N_3459);
xor U10752 (N_10752,N_6413,N_2668);
nand U10753 (N_10753,N_542,N_4125);
or U10754 (N_10754,N_1974,N_218);
xor U10755 (N_10755,N_20,N_2966);
nor U10756 (N_10756,N_1860,N_4827);
nor U10757 (N_10757,N_1971,N_36);
nor U10758 (N_10758,N_2186,N_5905);
nand U10759 (N_10759,N_1422,N_59);
nand U10760 (N_10760,N_5217,N_1449);
nor U10761 (N_10761,N_3997,N_7584);
nor U10762 (N_10762,N_924,N_8074);
nor U10763 (N_10763,N_4258,N_8651);
xnor U10764 (N_10764,N_8198,N_1332);
xnor U10765 (N_10765,N_6691,N_7248);
and U10766 (N_10766,N_2431,N_7525);
nand U10767 (N_10767,N_4756,N_3482);
nor U10768 (N_10768,N_3652,N_9478);
nand U10769 (N_10769,N_1592,N_3500);
xor U10770 (N_10770,N_7617,N_9380);
nor U10771 (N_10771,N_3538,N_7683);
nor U10772 (N_10772,N_6504,N_7239);
and U10773 (N_10773,N_7649,N_6988);
xnor U10774 (N_10774,N_4230,N_8632);
or U10775 (N_10775,N_2141,N_6962);
nor U10776 (N_10776,N_8804,N_256);
and U10777 (N_10777,N_4232,N_3311);
nor U10778 (N_10778,N_4859,N_8999);
or U10779 (N_10779,N_1029,N_6932);
nor U10780 (N_10780,N_4484,N_685);
or U10781 (N_10781,N_744,N_4401);
nand U10782 (N_10782,N_7497,N_2132);
nand U10783 (N_10783,N_1336,N_996);
or U10784 (N_10784,N_1357,N_319);
or U10785 (N_10785,N_6511,N_3752);
xor U10786 (N_10786,N_5653,N_1536);
or U10787 (N_10787,N_271,N_6907);
nor U10788 (N_10788,N_4094,N_961);
and U10789 (N_10789,N_1856,N_521);
or U10790 (N_10790,N_4383,N_4678);
nand U10791 (N_10791,N_7701,N_6436);
nand U10792 (N_10792,N_4443,N_6259);
nand U10793 (N_10793,N_9825,N_8356);
nor U10794 (N_10794,N_135,N_1691);
and U10795 (N_10795,N_7576,N_1892);
xor U10796 (N_10796,N_5607,N_1285);
nor U10797 (N_10797,N_5387,N_2100);
nand U10798 (N_10798,N_4530,N_2304);
nand U10799 (N_10799,N_8923,N_4958);
nand U10800 (N_10800,N_6677,N_7721);
nor U10801 (N_10801,N_8463,N_6085);
nand U10802 (N_10802,N_2964,N_2909);
nand U10803 (N_10803,N_7274,N_5889);
and U10804 (N_10804,N_2054,N_6177);
xor U10805 (N_10805,N_8666,N_559);
or U10806 (N_10806,N_9568,N_9300);
and U10807 (N_10807,N_9709,N_7282);
and U10808 (N_10808,N_2762,N_8043);
or U10809 (N_10809,N_3899,N_4875);
xnor U10810 (N_10810,N_2066,N_3656);
nor U10811 (N_10811,N_8940,N_3386);
xor U10812 (N_10812,N_2607,N_2540);
or U10813 (N_10813,N_6179,N_6584);
and U10814 (N_10814,N_5110,N_1744);
or U10815 (N_10815,N_207,N_2757);
and U10816 (N_10816,N_146,N_8426);
or U10817 (N_10817,N_3653,N_7958);
or U10818 (N_10818,N_5439,N_442);
nor U10819 (N_10819,N_4747,N_3481);
nand U10820 (N_10820,N_2252,N_618);
nand U10821 (N_10821,N_9159,N_4221);
nand U10822 (N_10822,N_6262,N_8557);
xnor U10823 (N_10823,N_3760,N_2089);
or U10824 (N_10824,N_5743,N_8593);
and U10825 (N_10825,N_3259,N_8606);
xor U10826 (N_10826,N_6364,N_9525);
nor U10827 (N_10827,N_5712,N_6658);
or U10828 (N_10828,N_4453,N_3638);
or U10829 (N_10829,N_5271,N_1545);
and U10830 (N_10830,N_897,N_6409);
nor U10831 (N_10831,N_8782,N_8280);
nand U10832 (N_10832,N_5871,N_9545);
nand U10833 (N_10833,N_5332,N_7957);
and U10834 (N_10834,N_5204,N_8206);
and U10835 (N_10835,N_3400,N_305);
and U10836 (N_10836,N_7670,N_999);
nand U10837 (N_10837,N_5863,N_9409);
nand U10838 (N_10838,N_5158,N_1849);
or U10839 (N_10839,N_68,N_8360);
and U10840 (N_10840,N_2090,N_1602);
nand U10841 (N_10841,N_6756,N_9966);
or U10842 (N_10842,N_4588,N_3564);
nand U10843 (N_10843,N_8186,N_6154);
nand U10844 (N_10844,N_4127,N_6450);
and U10845 (N_10845,N_4050,N_4514);
nand U10846 (N_10846,N_2049,N_1334);
nor U10847 (N_10847,N_8281,N_7241);
or U10848 (N_10848,N_4246,N_806);
and U10849 (N_10849,N_3310,N_1404);
or U10850 (N_10850,N_213,N_6362);
or U10851 (N_10851,N_8871,N_6906);
and U10852 (N_10852,N_2896,N_3625);
or U10853 (N_10853,N_795,N_7680);
or U10854 (N_10854,N_4387,N_6256);
xor U10855 (N_10855,N_144,N_5057);
nand U10856 (N_10856,N_4254,N_6608);
nor U10857 (N_10857,N_4078,N_1794);
xnor U10858 (N_10858,N_3934,N_9702);
nor U10859 (N_10859,N_6780,N_8235);
and U10860 (N_10860,N_5463,N_8411);
nand U10861 (N_10861,N_264,N_9544);
nand U10862 (N_10862,N_9583,N_2900);
or U10863 (N_10863,N_7826,N_9414);
nand U10864 (N_10864,N_4937,N_7225);
and U10865 (N_10865,N_4936,N_2284);
and U10866 (N_10866,N_9984,N_9877);
xor U10867 (N_10867,N_7089,N_4523);
and U10868 (N_10868,N_1643,N_9062);
and U10869 (N_10869,N_6299,N_7182);
nor U10870 (N_10870,N_1264,N_7761);
nor U10871 (N_10871,N_5213,N_3949);
nand U10872 (N_10872,N_4321,N_4397);
and U10873 (N_10873,N_5561,N_5419);
nor U10874 (N_10874,N_5588,N_7068);
xor U10875 (N_10875,N_4983,N_7984);
nor U10876 (N_10876,N_6887,N_977);
xor U10877 (N_10877,N_7363,N_6345);
and U10878 (N_10878,N_572,N_7021);
xnor U10879 (N_10879,N_4813,N_1533);
nand U10880 (N_10880,N_1399,N_9439);
xor U10881 (N_10881,N_5793,N_9802);
and U10882 (N_10882,N_1922,N_371);
or U10883 (N_10883,N_8119,N_9177);
or U10884 (N_10884,N_118,N_2103);
nor U10885 (N_10885,N_834,N_9218);
or U10886 (N_10886,N_2555,N_7212);
or U10887 (N_10887,N_2660,N_4598);
or U10888 (N_10888,N_4452,N_5642);
nand U10889 (N_10889,N_710,N_6106);
or U10890 (N_10890,N_7937,N_7919);
and U10891 (N_10891,N_6352,N_960);
or U10892 (N_10892,N_3146,N_295);
and U10893 (N_10893,N_2251,N_3440);
nand U10894 (N_10894,N_9365,N_5828);
or U10895 (N_10895,N_6549,N_9806);
and U10896 (N_10896,N_7436,N_8478);
or U10897 (N_10897,N_4219,N_8888);
nor U10898 (N_10898,N_3974,N_746);
nor U10899 (N_10899,N_627,N_7195);
xor U10900 (N_10900,N_8393,N_2365);
or U10901 (N_10901,N_127,N_7713);
xnor U10902 (N_10902,N_9189,N_4695);
or U10903 (N_10903,N_5859,N_1631);
or U10904 (N_10904,N_7735,N_642);
nand U10905 (N_10905,N_9394,N_5855);
xor U10906 (N_10906,N_9903,N_8345);
and U10907 (N_10907,N_1681,N_4167);
nor U10908 (N_10908,N_8244,N_308);
and U10909 (N_10909,N_2941,N_4681);
and U10910 (N_10910,N_6891,N_2230);
and U10911 (N_10911,N_2019,N_5265);
xnor U10912 (N_10912,N_3972,N_8546);
nor U10913 (N_10913,N_1797,N_4591);
or U10914 (N_10914,N_5933,N_9594);
xnor U10915 (N_10915,N_8223,N_7457);
nand U10916 (N_10916,N_2444,N_6543);
nand U10917 (N_10917,N_1439,N_1550);
and U10918 (N_10918,N_718,N_9862);
xor U10919 (N_10919,N_5124,N_1385);
nand U10920 (N_10920,N_6977,N_3387);
and U10921 (N_10921,N_4241,N_6517);
or U10922 (N_10922,N_9763,N_6003);
nand U10923 (N_10923,N_1202,N_6958);
and U10924 (N_10924,N_2724,N_9103);
and U10925 (N_10925,N_7655,N_7502);
nand U10926 (N_10926,N_5957,N_2659);
and U10927 (N_10927,N_803,N_8298);
or U10928 (N_10928,N_7982,N_1190);
xnor U10929 (N_10929,N_8893,N_647);
nor U10930 (N_10930,N_565,N_5983);
nand U10931 (N_10931,N_5996,N_7885);
nor U10932 (N_10932,N_5396,N_9666);
nand U10933 (N_10933,N_6942,N_2121);
xnor U10934 (N_10934,N_4073,N_4639);
and U10935 (N_10935,N_5394,N_4906);
xnor U10936 (N_10936,N_9296,N_8719);
nand U10937 (N_10937,N_2204,N_1843);
xor U10938 (N_10938,N_7654,N_2123);
xnor U10939 (N_10939,N_6890,N_8682);
xnor U10940 (N_10940,N_7297,N_2062);
nand U10941 (N_10941,N_5627,N_8001);
nor U10942 (N_10942,N_693,N_3044);
and U10943 (N_10943,N_5550,N_1867);
nor U10944 (N_10944,N_7740,N_6878);
nor U10945 (N_10945,N_4448,N_4490);
and U10946 (N_10946,N_3608,N_6066);
nand U10947 (N_10947,N_3558,N_9408);
nand U10948 (N_10948,N_7789,N_3039);
or U10949 (N_10949,N_5366,N_9578);
nor U10950 (N_10950,N_3053,N_8089);
nand U10951 (N_10951,N_5300,N_5808);
xor U10952 (N_10952,N_5546,N_8256);
and U10953 (N_10953,N_8694,N_6378);
nor U10954 (N_10954,N_2367,N_1635);
or U10955 (N_10955,N_8574,N_9153);
nand U10956 (N_10956,N_4799,N_3979);
or U10957 (N_10957,N_7388,N_9948);
or U10958 (N_10958,N_3762,N_4841);
nor U10959 (N_10959,N_3005,N_3077);
nand U10960 (N_10960,N_4493,N_2091);
nand U10961 (N_10961,N_3203,N_6184);
and U10962 (N_10962,N_8321,N_7112);
or U10963 (N_10963,N_215,N_681);
xor U10964 (N_10964,N_9581,N_2508);
nor U10965 (N_10965,N_2466,N_5344);
nor U10966 (N_10966,N_7328,N_5739);
nand U10967 (N_10967,N_4194,N_4460);
or U10968 (N_10968,N_6221,N_534);
nor U10969 (N_10969,N_5261,N_8800);
nor U10970 (N_10970,N_2846,N_63);
xor U10971 (N_10971,N_4041,N_5671);
xor U10972 (N_10972,N_1068,N_7821);
and U10973 (N_10973,N_3826,N_5095);
xor U10974 (N_10974,N_65,N_156);
or U10975 (N_10975,N_1413,N_3173);
nand U10976 (N_10976,N_314,N_7948);
nand U10977 (N_10977,N_5662,N_9404);
xnor U10978 (N_10978,N_9838,N_5657);
nand U10979 (N_10979,N_6764,N_9470);
nor U10980 (N_10980,N_7996,N_7785);
nor U10981 (N_10981,N_2079,N_9205);
and U10982 (N_10982,N_126,N_2146);
or U10983 (N_10983,N_4910,N_626);
or U10984 (N_10984,N_5780,N_1105);
or U10985 (N_10985,N_913,N_2134);
and U10986 (N_10986,N_6776,N_2782);
nor U10987 (N_10987,N_1820,N_3267);
nand U10988 (N_10988,N_2820,N_1221);
or U10989 (N_10989,N_7861,N_9967);
or U10990 (N_10990,N_6470,N_3996);
xor U10991 (N_10991,N_6671,N_752);
or U10992 (N_10992,N_3099,N_3822);
xor U10993 (N_10993,N_8931,N_6162);
xor U10994 (N_10994,N_5913,N_6761);
xor U10995 (N_10995,N_6152,N_6459);
nand U10996 (N_10996,N_9526,N_8689);
xor U10997 (N_10997,N_7983,N_2192);
or U10998 (N_10998,N_6071,N_1995);
xnor U10999 (N_10999,N_1606,N_4646);
nand U11000 (N_11000,N_9805,N_8168);
nor U11001 (N_11001,N_3468,N_5170);
xnor U11002 (N_11002,N_1007,N_9639);
or U11003 (N_11003,N_3905,N_6574);
and U11004 (N_11004,N_971,N_3499);
and U11005 (N_11005,N_4414,N_8255);
and U11006 (N_11006,N_6229,N_3925);
or U11007 (N_11007,N_5538,N_1647);
nand U11008 (N_11008,N_1828,N_4614);
xor U11009 (N_11009,N_2336,N_239);
and U11010 (N_11010,N_9971,N_6837);
xnor U11011 (N_11011,N_1504,N_5860);
xnor U11012 (N_11012,N_703,N_1610);
or U11013 (N_11013,N_7079,N_8103);
nor U11014 (N_11014,N_83,N_2862);
or U11015 (N_11015,N_7165,N_4566);
or U11016 (N_11016,N_2832,N_3195);
or U11017 (N_11017,N_1380,N_4821);
xor U11018 (N_11018,N_1837,N_6772);
and U11019 (N_11019,N_1585,N_1703);
nor U11020 (N_11020,N_4881,N_9629);
nor U11021 (N_11021,N_270,N_8007);
xnor U11022 (N_11022,N_5769,N_5032);
nand U11023 (N_11023,N_6708,N_5298);
or U11024 (N_11024,N_9253,N_7304);
and U11025 (N_11025,N_3010,N_9020);
nor U11026 (N_11026,N_6297,N_4303);
and U11027 (N_11027,N_8394,N_2845);
xor U11028 (N_11028,N_8004,N_762);
nor U11029 (N_11029,N_1327,N_1376);
xnor U11030 (N_11030,N_5034,N_9457);
or U11031 (N_11031,N_5386,N_577);
or U11032 (N_11032,N_5581,N_8016);
or U11033 (N_11033,N_170,N_4087);
and U11034 (N_11034,N_6809,N_7742);
nor U11035 (N_11035,N_9144,N_5836);
nand U11036 (N_11036,N_788,N_5968);
and U11037 (N_11037,N_8986,N_8538);
and U11038 (N_11038,N_2472,N_9579);
and U11039 (N_11039,N_9509,N_2026);
or U11040 (N_11040,N_1401,N_4933);
or U11041 (N_11041,N_7776,N_8856);
or U11042 (N_11042,N_1446,N_9664);
nand U11043 (N_11043,N_4029,N_5119);
or U11044 (N_11044,N_4965,N_1070);
nor U11045 (N_11045,N_1483,N_3090);
or U11046 (N_11046,N_1167,N_6208);
nor U11047 (N_11047,N_6882,N_7757);
and U11048 (N_11048,N_4128,N_6127);
and U11049 (N_11049,N_3983,N_1248);
or U11050 (N_11050,N_6547,N_6866);
nand U11051 (N_11051,N_7804,N_7814);
or U11052 (N_11052,N_7652,N_6989);
nor U11053 (N_11053,N_2938,N_1317);
xor U11054 (N_11054,N_9506,N_9173);
and U11055 (N_11055,N_5559,N_3489);
xor U11056 (N_11056,N_2129,N_358);
or U11057 (N_11057,N_7618,N_1627);
or U11058 (N_11058,N_8240,N_9672);
and U11059 (N_11059,N_373,N_9992);
xor U11060 (N_11060,N_8329,N_2807);
or U11061 (N_11061,N_134,N_8851);
xor U11062 (N_11062,N_292,N_3296);
and U11063 (N_11063,N_5864,N_9874);
nand U11064 (N_11064,N_5881,N_6775);
and U11065 (N_11065,N_9476,N_697);
and U11066 (N_11066,N_1789,N_152);
or U11067 (N_11067,N_5522,N_3278);
or U11068 (N_11068,N_8429,N_7636);
nand U11069 (N_11069,N_1570,N_3738);
nand U11070 (N_11070,N_1738,N_6935);
xor U11071 (N_11071,N_6482,N_9229);
or U11072 (N_11072,N_1779,N_3610);
xor U11073 (N_11073,N_5282,N_8944);
and U11074 (N_11074,N_7947,N_1981);
and U11075 (N_11075,N_3929,N_8000);
nor U11076 (N_11076,N_9057,N_6894);
and U11077 (N_11077,N_7879,N_5377);
xnor U11078 (N_11078,N_7732,N_6802);
xnor U11079 (N_11079,N_2164,N_9485);
xnor U11080 (N_11080,N_9662,N_7428);
and U11081 (N_11081,N_1251,N_3914);
nor U11082 (N_11082,N_3269,N_8101);
or U11083 (N_11083,N_8821,N_1913);
or U11084 (N_11084,N_7629,N_981);
nor U11085 (N_11085,N_9935,N_726);
nor U11086 (N_11086,N_2223,N_5576);
and U11087 (N_11087,N_8288,N_4606);
nor U11088 (N_11088,N_8640,N_8117);
nor U11089 (N_11089,N_8475,N_7117);
nand U11090 (N_11090,N_7492,N_2196);
nor U11091 (N_11091,N_8832,N_1906);
xnor U11092 (N_11092,N_2138,N_2578);
and U11093 (N_11093,N_8966,N_6423);
nor U11094 (N_11094,N_3801,N_452);
xor U11095 (N_11095,N_6429,N_7078);
nand U11096 (N_11096,N_8860,N_5380);
xnor U11097 (N_11097,N_4098,N_4741);
and U11098 (N_11098,N_3599,N_8128);
or U11099 (N_11099,N_669,N_3935);
xnor U11100 (N_11100,N_6595,N_5159);
nand U11101 (N_11101,N_1634,N_4440);
or U11102 (N_11102,N_9591,N_2915);
nand U11103 (N_11103,N_9695,N_1870);
or U11104 (N_11104,N_2823,N_9009);
xnor U11105 (N_11105,N_2379,N_6166);
nor U11106 (N_11106,N_7746,N_854);
and U11107 (N_11107,N_2193,N_4818);
nand U11108 (N_11108,N_6319,N_563);
nor U11109 (N_11109,N_3704,N_242);
and U11110 (N_11110,N_4592,N_5502);
or U11111 (N_11111,N_1579,N_4518);
nand U11112 (N_11112,N_1873,N_5495);
nand U11113 (N_11113,N_6933,N_2397);
nor U11114 (N_11114,N_4919,N_4901);
nand U11115 (N_11115,N_2666,N_672);
nand U11116 (N_11116,N_7320,N_6333);
nand U11117 (N_11117,N_7532,N_6575);
and U11118 (N_11118,N_3136,N_7890);
nand U11119 (N_11119,N_8224,N_3756);
or U11120 (N_11120,N_3753,N_8221);
or U11121 (N_11121,N_3234,N_9611);
nand U11122 (N_11122,N_2962,N_9075);
or U11123 (N_11123,N_8591,N_8935);
and U11124 (N_11124,N_6805,N_5735);
nand U11125 (N_11125,N_1352,N_1724);
nand U11126 (N_11126,N_1083,N_9349);
nand U11127 (N_11127,N_328,N_4511);
nand U11128 (N_11128,N_5613,N_1268);
and U11129 (N_11129,N_662,N_9592);
or U11130 (N_11130,N_8575,N_1072);
or U11131 (N_11131,N_1037,N_716);
nor U11132 (N_11132,N_2391,N_3314);
nor U11133 (N_11133,N_3970,N_2259);
nand U11134 (N_11134,N_8829,N_5073);
nand U11135 (N_11135,N_6443,N_2292);
and U11136 (N_11136,N_8687,N_1511);
and U11137 (N_11137,N_5296,N_9751);
nor U11138 (N_11138,N_2737,N_5289);
xnor U11139 (N_11139,N_9363,N_3842);
or U11140 (N_11140,N_5579,N_4163);
nor U11141 (N_11141,N_5081,N_1622);
nor U11142 (N_11142,N_2700,N_6206);
or U11143 (N_11143,N_9647,N_7235);
nor U11144 (N_11144,N_6369,N_4675);
xor U11145 (N_11145,N_480,N_3922);
and U11146 (N_11146,N_3264,N_777);
nand U11147 (N_11147,N_3647,N_6609);
and U11148 (N_11148,N_3553,N_7484);
nor U11149 (N_11149,N_1607,N_5464);
nor U11150 (N_11150,N_7765,N_8659);
nand U11151 (N_11151,N_9166,N_5706);
nor U11152 (N_11152,N_9148,N_591);
nand U11153 (N_11153,N_4570,N_4711);
nand U11154 (N_11154,N_2571,N_7145);
nand U11155 (N_11155,N_713,N_7356);
nand U11156 (N_11156,N_6983,N_4091);
or U11157 (N_11157,N_8745,N_3471);
or U11158 (N_11158,N_6666,N_9556);
nor U11159 (N_11159,N_3352,N_2085);
xor U11160 (N_11160,N_5945,N_1766);
or U11161 (N_11161,N_323,N_9740);
and U11162 (N_11162,N_7135,N_5002);
and U11163 (N_11163,N_392,N_3782);
nand U11164 (N_11164,N_2238,N_862);
xnor U11165 (N_11165,N_4485,N_9641);
or U11166 (N_11166,N_336,N_1240);
or U11167 (N_11167,N_3211,N_5193);
nor U11168 (N_11168,N_265,N_4075);
and U11169 (N_11169,N_5533,N_9430);
nand U11170 (N_11170,N_4432,N_1491);
or U11171 (N_11171,N_8294,N_9029);
nor U11172 (N_11172,N_6334,N_6069);
xnor U11173 (N_11173,N_8276,N_551);
nand U11174 (N_11174,N_8228,N_8290);
and U11175 (N_11175,N_7083,N_8836);
nand U11176 (N_11176,N_3861,N_9034);
or U11177 (N_11177,N_2215,N_4024);
nor U11178 (N_11178,N_9090,N_3123);
and U11179 (N_11179,N_4212,N_316);
nor U11180 (N_11180,N_1546,N_2816);
and U11181 (N_11181,N_4930,N_3686);
and U11182 (N_11182,N_1612,N_8978);
or U11183 (N_11183,N_3723,N_5350);
and U11184 (N_11184,N_9939,N_2874);
and U11185 (N_11185,N_4408,N_7470);
or U11186 (N_11186,N_6697,N_1758);
xor U11187 (N_11187,N_1807,N_1367);
xnor U11188 (N_11188,N_9242,N_2353);
nand U11189 (N_11189,N_3823,N_122);
xnor U11190 (N_11190,N_6397,N_8359);
nor U11191 (N_11191,N_8377,N_4702);
xnor U11192 (N_11192,N_7876,N_8892);
nand U11193 (N_11193,N_3002,N_7531);
nand U11194 (N_11194,N_6741,N_839);
nor U11195 (N_11195,N_9569,N_7220);
nor U11196 (N_11196,N_6062,N_8726);
nand U11197 (N_11197,N_3709,N_6400);
or U11198 (N_11198,N_3290,N_3376);
and U11199 (N_11199,N_1803,N_282);
or U11200 (N_11200,N_5658,N_532);
nor U11201 (N_11201,N_7013,N_5901);
nand U11202 (N_11202,N_4920,N_6799);
nor U11203 (N_11203,N_9765,N_6279);
nor U11204 (N_11204,N_5921,N_7626);
nand U11205 (N_11205,N_9309,N_8551);
nand U11206 (N_11206,N_8401,N_9951);
and U11207 (N_11207,N_1868,N_237);
or U11208 (N_11208,N_8922,N_503);
or U11209 (N_11209,N_4395,N_9);
or U11210 (N_11210,N_4355,N_9686);
nor U11211 (N_11211,N_8445,N_9582);
nand U11212 (N_11212,N_2877,N_8346);
or U11213 (N_11213,N_1846,N_8455);
nand U11214 (N_11214,N_3212,N_8528);
and U11215 (N_11215,N_1861,N_9585);
nand U11216 (N_11216,N_5086,N_9876);
and U11217 (N_11217,N_57,N_6505);
nor U11218 (N_11218,N_9001,N_6847);
nor U11219 (N_11219,N_2383,N_9849);
xnor U11220 (N_11220,N_830,N_9037);
or U11221 (N_11221,N_6976,N_3870);
xor U11222 (N_11222,N_2539,N_3001);
or U11223 (N_11223,N_7795,N_3384);
xor U11224 (N_11224,N_4739,N_6810);
nor U11225 (N_11225,N_8297,N_6553);
nor U11226 (N_11226,N_6215,N_8071);
xnor U11227 (N_11227,N_8980,N_210);
and U11228 (N_11228,N_9451,N_5202);
nor U11229 (N_11229,N_4312,N_948);
and U11230 (N_11230,N_2680,N_4929);
nand U11231 (N_11231,N_5511,N_1710);
and U11232 (N_11232,N_644,N_2236);
and U11233 (N_11233,N_7345,N_9536);
nand U11234 (N_11234,N_8452,N_1172);
or U11235 (N_11235,N_3809,N_1252);
and U11236 (N_11236,N_1312,N_4712);
nor U11237 (N_11237,N_5222,N_942);
and U11238 (N_11238,N_6884,N_980);
nor U11239 (N_11239,N_4607,N_7803);
nor U11240 (N_11240,N_4158,N_2012);
and U11241 (N_11241,N_3850,N_6125);
nor U11242 (N_11242,N_3713,N_7299);
xor U11243 (N_11243,N_3559,N_9138);
nand U11244 (N_11244,N_2372,N_7406);
and U11245 (N_11245,N_9232,N_6663);
xnor U11246 (N_11246,N_5330,N_18);
and U11247 (N_11247,N_7976,N_4754);
nor U11248 (N_11248,N_6232,N_2818);
nor U11249 (N_11249,N_760,N_2264);
and U11250 (N_11250,N_9969,N_7946);
nor U11251 (N_11251,N_9891,N_6940);
nor U11252 (N_11252,N_4532,N_5844);
nand U11253 (N_11253,N_1498,N_3255);
and U11254 (N_11254,N_1548,N_4916);
nor U11255 (N_11255,N_9759,N_2566);
or U11256 (N_11256,N_5385,N_8875);
or U11257 (N_11257,N_9092,N_2068);
nand U11258 (N_11258,N_9226,N_6588);
nand U11259 (N_11259,N_1934,N_1830);
and U11260 (N_11260,N_6725,N_8716);
nor U11261 (N_11261,N_3055,N_6625);
and U11262 (N_11262,N_1600,N_4417);
or U11263 (N_11263,N_2393,N_6359);
or U11264 (N_11264,N_6240,N_3948);
nor U11265 (N_11265,N_3372,N_3461);
and U11266 (N_11266,N_2240,N_1586);
and U11267 (N_11267,N_4057,N_3257);
nor U11268 (N_11268,N_3298,N_5754);
or U11269 (N_11269,N_2345,N_3665);
nand U11270 (N_11270,N_5516,N_4243);
and U11271 (N_11271,N_9945,N_2965);
nand U11272 (N_11272,N_8506,N_2638);
nor U11273 (N_11273,N_7110,N_6272);
nor U11274 (N_11274,N_5024,N_851);
xor U11275 (N_11275,N_759,N_9008);
nor U11276 (N_11276,N_5120,N_2983);
and U11277 (N_11277,N_4068,N_5848);
and U11278 (N_11278,N_9527,N_509);
or U11279 (N_11279,N_8059,N_6630);
and U11280 (N_11280,N_6053,N_2401);
or U11281 (N_11281,N_2380,N_1816);
nand U11282 (N_11282,N_7333,N_3460);
xor U11283 (N_11283,N_4262,N_8485);
or U11284 (N_11284,N_3323,N_7486);
xnor U11285 (N_11285,N_4618,N_4470);
nand U11286 (N_11286,N_1143,N_2027);
xnor U11287 (N_11287,N_6996,N_1874);
nor U11288 (N_11288,N_9085,N_4672);
or U11289 (N_11289,N_4335,N_7903);
xnor U11290 (N_11290,N_2456,N_1112);
nand U11291 (N_11291,N_3023,N_822);
or U11292 (N_11292,N_5334,N_4550);
and U11293 (N_11293,N_738,N_9972);
or U11294 (N_11294,N_9047,N_5096);
and U11295 (N_11295,N_8969,N_8879);
nand U11296 (N_11296,N_8765,N_9787);
xnor U11297 (N_11297,N_4989,N_7483);
and U11298 (N_11298,N_2761,N_9764);
nor U11299 (N_11299,N_6635,N_6207);
or U11300 (N_11300,N_6699,N_8082);
nand U11301 (N_11301,N_7134,N_9422);
nor U11302 (N_11302,N_8234,N_7114);
nor U11303 (N_11303,N_6564,N_3513);
nand U11304 (N_11304,N_5936,N_9366);
and U11305 (N_11305,N_964,N_7010);
and U11306 (N_11306,N_2657,N_9934);
nor U11307 (N_11307,N_5634,N_6236);
xnor U11308 (N_11308,N_8525,N_7137);
nor U11309 (N_11309,N_2683,N_571);
nor U11310 (N_11310,N_9141,N_2623);
nor U11311 (N_11311,N_8178,N_4797);
xnor U11312 (N_11312,N_4428,N_4268);
nand U11313 (N_11313,N_6566,N_4957);
or U11314 (N_11314,N_988,N_7348);
nor U11315 (N_11315,N_5215,N_5224);
and U11316 (N_11316,N_9255,N_5453);
xnor U11317 (N_11317,N_6288,N_7277);
and U11318 (N_11318,N_5554,N_7868);
nand U11319 (N_11319,N_3955,N_8285);
or U11320 (N_11320,N_529,N_1305);
nor U11321 (N_11321,N_3329,N_4743);
and U11322 (N_11322,N_4814,N_666);
xor U11323 (N_11323,N_7985,N_6978);
nand U11324 (N_11324,N_398,N_791);
and U11325 (N_11325,N_7887,N_6190);
or U11326 (N_11326,N_5417,N_3409);
xnor U11327 (N_11327,N_7413,N_9964);
or U11328 (N_11328,N_1226,N_123);
nor U11329 (N_11329,N_7341,N_41);
or U11330 (N_11330,N_8607,N_9067);
nor U11331 (N_11331,N_6921,N_3622);
nand U11332 (N_11332,N_8542,N_5220);
nand U11333 (N_11333,N_7032,N_335);
and U11334 (N_11334,N_2040,N_9336);
or U11335 (N_11335,N_2470,N_1573);
xor U11336 (N_11336,N_1541,N_2044);
nand U11337 (N_11337,N_5557,N_4251);
or U11338 (N_11338,N_3837,N_4939);
nor U11339 (N_11339,N_8295,N_6383);
xor U11340 (N_11340,N_7597,N_1443);
nand U11341 (N_11341,N_8371,N_3921);
and U11342 (N_11342,N_4378,N_2360);
or U11343 (N_11343,N_7633,N_1748);
nor U11344 (N_11344,N_6499,N_7638);
xnor U11345 (N_11345,N_2549,N_6185);
and U11346 (N_11346,N_8537,N_990);
nand U11347 (N_11347,N_9095,N_6337);
or U11348 (N_11348,N_1696,N_223);
nand U11349 (N_11349,N_448,N_3);
or U11350 (N_11350,N_261,N_9853);
or U11351 (N_11351,N_3497,N_9193);
nor U11352 (N_11352,N_9222,N_623);
nand U11353 (N_11353,N_5929,N_9797);
xor U11354 (N_11354,N_4893,N_8230);
and U11355 (N_11355,N_7040,N_5907);
nand U11356 (N_11356,N_2432,N_186);
and U11357 (N_11357,N_9810,N_8808);
nor U11358 (N_11358,N_333,N_5535);
nand U11359 (N_11359,N_4497,N_3967);
or U11360 (N_11360,N_4285,N_4560);
or U11361 (N_11361,N_1996,N_9322);
xnor U11362 (N_11362,N_2083,N_1717);
or U11363 (N_11363,N_6812,N_8798);
xnor U11364 (N_11364,N_7257,N_4784);
nand U11365 (N_11365,N_9790,N_2849);
nor U11366 (N_11366,N_5713,N_8937);
nor U11367 (N_11367,N_4557,N_8728);
or U11368 (N_11368,N_3443,N_3351);
nand U11369 (N_11369,N_9941,N_6654);
xor U11370 (N_11370,N_2573,N_2249);
nor U11371 (N_11371,N_970,N_2254);
nor U11372 (N_11372,N_3880,N_3418);
nor U11373 (N_11373,N_3951,N_7712);
and U11374 (N_11374,N_6678,N_5058);
or U11375 (N_11375,N_71,N_7039);
nand U11376 (N_11376,N_76,N_5944);
or U11377 (N_11377,N_9803,N_9383);
xnor U11378 (N_11378,N_3343,N_6768);
xnor U11379 (N_11379,N_8284,N_6737);
xnor U11380 (N_11380,N_8012,N_7692);
nor U11381 (N_11381,N_6010,N_7551);
xor U11382 (N_11382,N_8003,N_5345);
nor U11383 (N_11383,N_6861,N_7337);
xnor U11384 (N_11384,N_3247,N_8599);
nor U11385 (N_11385,N_4501,N_1844);
and U11386 (N_11386,N_7031,N_8673);
and U11387 (N_11387,N_6690,N_6748);
xor U11388 (N_11388,N_9204,N_4018);
nor U11389 (N_11389,N_2417,N_8928);
nor U11390 (N_11390,N_1313,N_3153);
nor U11391 (N_11391,N_114,N_1910);
nor U11392 (N_11392,N_4535,N_915);
nor U11393 (N_11393,N_3603,N_3284);
nand U11394 (N_11394,N_32,N_8496);
xnor U11395 (N_11395,N_5701,N_7289);
and U11396 (N_11396,N_2977,N_1127);
nor U11397 (N_11397,N_4361,N_5728);
nand U11398 (N_11398,N_5834,N_4613);
nor U11399 (N_11399,N_6981,N_167);
or U11400 (N_11400,N_8638,N_1991);
or U11401 (N_11401,N_3926,N_7358);
nand U11402 (N_11402,N_6619,N_1395);
xor U11403 (N_11403,N_197,N_7526);
or U11404 (N_11404,N_9210,N_5540);
nand U11405 (N_11405,N_699,N_8140);
xnor U11406 (N_11406,N_928,N_7590);
or U11407 (N_11407,N_9977,N_2643);
and U11408 (N_11408,N_7323,N_9274);
nor U11409 (N_11409,N_8476,N_4472);
or U11410 (N_11410,N_3362,N_3793);
nand U11411 (N_11411,N_8941,N_5336);
nor U11412 (N_11412,N_6556,N_5734);
and U11413 (N_11413,N_5512,N_3154);
or U11414 (N_11414,N_7724,N_5226);
or U11415 (N_11415,N_7447,N_2888);
nand U11416 (N_11416,N_5469,N_430);
or U11417 (N_11417,N_1705,N_19);
xor U11418 (N_11418,N_4239,N_6787);
nand U11419 (N_11419,N_5312,N_9817);
and U11420 (N_11420,N_3986,N_2497);
nor U11421 (N_11421,N_6045,N_2794);
nand U11422 (N_11422,N_7730,N_2702);
nor U11423 (N_11423,N_3126,N_4445);
nand U11424 (N_11424,N_1052,N_9392);
nand U11425 (N_11425,N_440,N_9563);
and U11426 (N_11426,N_1495,N_7344);
nand U11427 (N_11427,N_6762,N_3350);
nand U11428 (N_11428,N_8670,N_3194);
or U11429 (N_11429,N_1931,N_2722);
xor U11430 (N_11430,N_6763,N_2008);
nand U11431 (N_11431,N_3486,N_3660);
and U11432 (N_11432,N_320,N_5719);
and U11433 (N_11433,N_4757,N_7046);
nor U11434 (N_11434,N_5766,N_6350);
nand U11435 (N_11435,N_224,N_6733);
and U11436 (N_11436,N_9190,N_8699);
nand U11437 (N_11437,N_4411,N_5031);
and U11438 (N_11438,N_5989,N_7856);
nand U11439 (N_11439,N_9894,N_4399);
nor U11440 (N_11440,N_8350,N_1986);
nand U11441 (N_11441,N_3128,N_2598);
nand U11442 (N_11442,N_30,N_1138);
nand U11443 (N_11443,N_2746,N_6858);
nand U11444 (N_11444,N_3395,N_9777);
nor U11445 (N_11445,N_6614,N_8292);
and U11446 (N_11446,N_2057,N_3892);
nand U11447 (N_11447,N_4021,N_3304);
or U11448 (N_11448,N_2149,N_8805);
nand U11449 (N_11449,N_9586,N_4339);
nor U11450 (N_11450,N_216,N_4336);
nor U11451 (N_11451,N_6916,N_7849);
or U11452 (N_11452,N_2798,N_1562);
nor U11453 (N_11453,N_8816,N_7387);
or U11454 (N_11454,N_2843,N_2780);
or U11455 (N_11455,N_6842,N_5357);
nand U11456 (N_11456,N_1686,N_2147);
or U11457 (N_11457,N_1760,N_7243);
or U11458 (N_11458,N_5146,N_1589);
or U11459 (N_11459,N_1020,N_2831);
xnor U11460 (N_11460,N_5582,N_7555);
and U11461 (N_11461,N_4992,N_423);
and U11462 (N_11462,N_932,N_7190);
xnor U11463 (N_11463,N_9194,N_8693);
and U11464 (N_11464,N_6355,N_69);
or U11465 (N_11465,N_695,N_9924);
xor U11466 (N_11466,N_6874,N_2622);
xnor U11467 (N_11467,N_7774,N_813);
or U11468 (N_11468,N_9724,N_3375);
nand U11469 (N_11469,N_4734,N_3202);
nand U11470 (N_11470,N_7528,N_8613);
nand U11471 (N_11471,N_5507,N_399);
nor U11472 (N_11472,N_5543,N_8950);
nor U11473 (N_11473,N_561,N_5727);
and U11474 (N_11474,N_7127,N_4576);
or U11475 (N_11475,N_6765,N_7544);
xor U11476 (N_11476,N_1474,N_7900);
nand U11477 (N_11477,N_3111,N_1572);
nand U11478 (N_11478,N_6616,N_8710);
xor U11479 (N_11479,N_9111,N_2023);
and U11480 (N_11480,N_6330,N_3472);
nand U11481 (N_11481,N_9882,N_7522);
or U11482 (N_11482,N_6969,N_116);
and U11483 (N_11483,N_4751,N_5560);
xor U11484 (N_11484,N_5171,N_579);
or U11485 (N_11485,N_8180,N_9223);
and U11486 (N_11486,N_5038,N_2298);
nor U11487 (N_11487,N_8141,N_7627);
and U11488 (N_11488,N_7463,N_5778);
nor U11489 (N_11489,N_1566,N_3514);
xnor U11490 (N_11490,N_6729,N_5827);
or U11491 (N_11491,N_3008,N_3909);
xnor U11492 (N_11492,N_9533,N_1587);
and U11493 (N_11493,N_3984,N_6270);
and U11494 (N_11494,N_2,N_958);
nor U11495 (N_11495,N_6371,N_129);
xor U11496 (N_11496,N_7545,N_863);
xor U11497 (N_11497,N_9942,N_4324);
or U11498 (N_11498,N_6790,N_6130);
or U11499 (N_11499,N_9041,N_5838);
nand U11500 (N_11500,N_5749,N_5951);
or U11501 (N_11501,N_4373,N_523);
or U11502 (N_11502,N_7930,N_8625);
nor U11503 (N_11503,N_966,N_4553);
nand U11504 (N_11504,N_3783,N_6963);
and U11505 (N_11505,N_6375,N_4649);
nand U11506 (N_11506,N_6473,N_2787);
nand U11507 (N_11507,N_8771,N_6865);
and U11508 (N_11508,N_7960,N_9165);
or U11509 (N_11509,N_46,N_7660);
nand U11510 (N_11510,N_141,N_6707);
nand U11511 (N_11511,N_2170,N_9436);
nor U11512 (N_11512,N_5196,N_8704);
nand U11513 (N_11513,N_3821,N_9256);
nand U11514 (N_11514,N_1073,N_348);
nor U11515 (N_11515,N_4011,N_6862);
nor U11516 (N_11516,N_9214,N_5730);
xnor U11517 (N_11517,N_3863,N_6311);
or U11518 (N_11518,N_7173,N_6672);
xnor U11519 (N_11519,N_150,N_8934);
or U11520 (N_11520,N_9922,N_6049);
nor U11521 (N_11521,N_2501,N_6853);
xnor U11522 (N_11522,N_1479,N_2564);
and U11523 (N_11523,N_7931,N_5379);
or U11524 (N_11524,N_7339,N_6181);
and U11525 (N_11525,N_5275,N_8979);
xnor U11526 (N_11526,N_6001,N_417);
or U11527 (N_11527,N_4508,N_8796);
xnor U11528 (N_11528,N_2392,N_3496);
or U11529 (N_11529,N_891,N_7331);
nand U11530 (N_11530,N_4682,N_6743);
nor U11531 (N_11531,N_7425,N_1353);
and U11532 (N_11532,N_6848,N_4347);
nand U11533 (N_11533,N_2743,N_7223);
or U11534 (N_11534,N_8320,N_3913);
nand U11535 (N_11535,N_5720,N_1140);
or U11536 (N_11536,N_3271,N_3377);
and U11537 (N_11537,N_4837,N_306);
xnor U11538 (N_11538,N_4956,N_1968);
and U11539 (N_11539,N_7191,N_5694);
xor U11540 (N_11540,N_747,N_1652);
nor U11541 (N_11541,N_8018,N_7723);
or U11542 (N_11542,N_2696,N_7273);
nand U11543 (N_11543,N_9030,N_3991);
nor U11544 (N_11544,N_6115,N_8545);
nor U11545 (N_11545,N_1481,N_7143);
nor U11546 (N_11546,N_9791,N_4487);
nor U11547 (N_11547,N_8921,N_2704);
xor U11548 (N_11548,N_9901,N_9387);
nand U11549 (N_11549,N_220,N_2930);
and U11550 (N_11550,N_3530,N_5214);
xnor U11551 (N_11551,N_5595,N_21);
and U11552 (N_11552,N_5796,N_4840);
xor U11553 (N_11553,N_4526,N_608);
xnor U11554 (N_11554,N_8354,N_6676);
nand U11555 (N_11555,N_7605,N_5532);
and U11556 (N_11556,N_67,N_3118);
xor U11557 (N_11557,N_2201,N_2294);
xnor U11558 (N_11558,N_4847,N_1679);
nor U11559 (N_11559,N_6331,N_6960);
xor U11560 (N_11560,N_6416,N_9080);
xor U11561 (N_11561,N_2234,N_7131);
nor U11562 (N_11562,N_7969,N_2503);
xnor U11563 (N_11563,N_9174,N_870);
nor U11564 (N_11564,N_6687,N_3764);
xor U11565 (N_11565,N_4645,N_8330);
or U11566 (N_11566,N_2663,N_6178);
nand U11567 (N_11567,N_9997,N_3649);
xor U11568 (N_11568,N_3591,N_4330);
nor U11569 (N_11569,N_1777,N_9472);
and U11570 (N_11570,N_3341,N_4892);
or U11571 (N_11571,N_5033,N_5465);
nand U11572 (N_11572,N_1659,N_4273);
nor U11573 (N_11573,N_3867,N_6277);
and U11574 (N_11574,N_3575,N_5504);
nand U11575 (N_11575,N_3568,N_4278);
nor U11576 (N_11576,N_8326,N_8637);
nand U11577 (N_11577,N_4973,N_3992);
or U11578 (N_11578,N_8067,N_6521);
or U11579 (N_11579,N_6668,N_7972);
and U11580 (N_11580,N_564,N_8193);
or U11581 (N_11581,N_2041,N_9866);
xor U11582 (N_11582,N_8322,N_2546);
xnor U11583 (N_11583,N_3078,N_1307);
xor U11584 (N_11584,N_9316,N_8680);
nor U11585 (N_11585,N_9983,N_3907);
nand U11586 (N_11586,N_7438,N_5970);
and U11587 (N_11587,N_2319,N_4669);
nor U11588 (N_11588,N_7482,N_9109);
or U11589 (N_11589,N_5155,N_1);
and U11590 (N_11590,N_2637,N_9145);
and U11591 (N_11591,N_2131,N_8383);
nand U11592 (N_11592,N_7149,N_8286);
nand U11593 (N_11593,N_6592,N_5331);
nor U11594 (N_11594,N_6791,N_6394);
xnor U11595 (N_11595,N_1042,N_5691);
xnor U11596 (N_11596,N_4442,N_2325);
and U11597 (N_11597,N_201,N_7162);
nor U11598 (N_11598,N_9114,N_7709);
or U11599 (N_11599,N_7412,N_8176);
and U11600 (N_11600,N_661,N_6830);
and U11601 (N_11601,N_99,N_4585);
and U11602 (N_11602,N_1882,N_7598);
or U11603 (N_11603,N_3428,N_800);
and U11604 (N_11604,N_2852,N_8453);
and U11605 (N_11605,N_8054,N_7656);
or U11606 (N_11606,N_8165,N_9739);
or U11607 (N_11607,N_3888,N_3800);
xor U11608 (N_11608,N_7433,N_3340);
and U11609 (N_11609,N_735,N_5373);
and U11610 (N_11610,N_4441,N_441);
nor U11611 (N_11611,N_6480,N_7686);
or U11612 (N_11612,N_8435,N_7155);
nor U11613 (N_11613,N_1249,N_7107);
nor U11614 (N_11614,N_4584,N_9314);
nand U11615 (N_11615,N_7012,N_4857);
xnor U11616 (N_11616,N_7501,N_9637);
xnor U11617 (N_11617,N_2484,N_3287);
nor U11618 (N_11618,N_4382,N_1976);
xor U11619 (N_11619,N_2269,N_6151);
and U11620 (N_11620,N_782,N_3220);
or U11621 (N_11621,N_5786,N_1788);
nand U11622 (N_11622,N_3092,N_4422);
and U11623 (N_11623,N_3862,N_3076);
or U11624 (N_11624,N_1603,N_2708);
nor U11625 (N_11625,N_1412,N_860);
xnor U11626 (N_11626,N_6624,N_2388);
and U11627 (N_11627,N_4699,N_8850);
nor U11628 (N_11628,N_4777,N_3803);
nand U11629 (N_11629,N_4168,N_2748);
or U11630 (N_11630,N_4386,N_4248);
xnor U11631 (N_11631,N_1740,N_975);
nand U11632 (N_11632,N_7490,N_842);
and U11633 (N_11633,N_8561,N_3031);
nand U11634 (N_11634,N_6385,N_4089);
nor U11635 (N_11635,N_9023,N_4263);
and U11636 (N_11636,N_7578,N_8088);
or U11637 (N_11637,N_1651,N_6241);
or U11638 (N_11638,N_4922,N_2160);
and U11639 (N_11639,N_3609,N_7285);
and U11640 (N_11640,N_3187,N_7064);
and U11641 (N_11641,N_9618,N_3293);
and U11642 (N_11642,N_9268,N_8835);
nand U11643 (N_11643,N_408,N_7024);
nand U11644 (N_11644,N_9512,N_5762);
or U11645 (N_11645,N_1018,N_9024);
or U11646 (N_11646,N_8984,N_8963);
nor U11647 (N_11647,N_2389,N_2541);
and U11648 (N_11648,N_6316,N_2070);
nor U11649 (N_11649,N_7534,N_3664);
or U11650 (N_11650,N_6943,N_1781);
or U11651 (N_11651,N_2658,N_8723);
xnor U11652 (N_11652,N_5950,N_6425);
nand U11653 (N_11653,N_6072,N_3679);
nor U11654 (N_11654,N_8013,N_7444);
nor U11655 (N_11655,N_1929,N_7381);
nor U11656 (N_11656,N_2222,N_8029);
xnor U11657 (N_11657,N_8926,N_1750);
nor U11658 (N_11658,N_1720,N_1620);
nand U11659 (N_11659,N_7451,N_9294);
xor U11660 (N_11660,N_5190,N_502);
nor U11661 (N_11661,N_7615,N_8709);
xor U11662 (N_11662,N_6357,N_605);
or U11663 (N_11663,N_4763,N_3830);
xor U11664 (N_11664,N_6030,N_154);
nand U11665 (N_11665,N_172,N_2701);
nand U11666 (N_11666,N_5293,N_7734);
nand U11667 (N_11667,N_4971,N_4036);
xnor U11668 (N_11668,N_1156,N_9104);
nor U11669 (N_11669,N_4788,N_2878);
and U11670 (N_11670,N_8732,N_7442);
or U11671 (N_11671,N_6554,N_9775);
or U11672 (N_11672,N_6200,N_2955);
and U11673 (N_11673,N_1615,N_4667);
xor U11674 (N_11674,N_8400,N_1209);
nand U11675 (N_11675,N_7481,N_3915);
xor U11676 (N_11676,N_8200,N_1805);
or U11677 (N_11677,N_612,N_7941);
xnor U11678 (N_11678,N_6041,N_1729);
and U11679 (N_11679,N_5452,N_5049);
nand U11680 (N_11680,N_4,N_2172);
nand U11681 (N_11681,N_9234,N_9968);
or U11682 (N_11682,N_3509,N_6696);
nor U11683 (N_11683,N_5683,N_8578);
xnor U11684 (N_11684,N_1053,N_1301);
nor U11685 (N_11685,N_7033,N_1304);
nor U11686 (N_11686,N_4295,N_5179);
or U11687 (N_11687,N_7454,N_9169);
nor U11688 (N_11688,N_7383,N_1593);
and U11689 (N_11689,N_7520,N_2098);
or U11690 (N_11690,N_8480,N_8645);
nor U11691 (N_11691,N_7142,N_9927);
nand U11692 (N_11692,N_1802,N_4829);
xnor U11693 (N_11693,N_4032,N_4184);
or U11694 (N_11694,N_6021,N_266);
and U11695 (N_11695,N_3515,N_8873);
nand U11696 (N_11696,N_2437,N_5397);
and U11697 (N_11697,N_1626,N_3745);
nand U11698 (N_11698,N_5148,N_7272);
nand U11699 (N_11699,N_2998,N_687);
and U11700 (N_11700,N_6593,N_6143);
xnor U11701 (N_11701,N_8586,N_2632);
nor U11702 (N_11702,N_9707,N_602);
xor U11703 (N_11703,N_7449,N_7524);
nor U11704 (N_11704,N_2136,N_3089);
nand U11705 (N_11705,N_6800,N_296);
xor U11706 (N_11706,N_7240,N_9335);
nor U11707 (N_11707,N_3495,N_3325);
and U11708 (N_11708,N_9887,N_1732);
or U11709 (N_11709,N_8536,N_7234);
or U11710 (N_11710,N_944,N_4225);
nand U11711 (N_11711,N_5869,N_309);
nand U11712 (N_11712,N_4139,N_1094);
xor U11713 (N_11713,N_4828,N_1389);
xnor U11714 (N_11714,N_5450,N_6686);
nor U11715 (N_11715,N_3675,N_1384);
nor U11716 (N_11716,N_6956,N_7924);
nor U11717 (N_11717,N_7955,N_1234);
or U11718 (N_11718,N_1914,N_6064);
xnor U11719 (N_11719,N_7183,N_1753);
and U11720 (N_11720,N_8509,N_8130);
and U11721 (N_11721,N_2673,N_5426);
or U11722 (N_11722,N_9285,N_8553);
nand U11723 (N_11723,N_985,N_6431);
xnor U11724 (N_11724,N_5569,N_3475);
and U11725 (N_11725,N_4903,N_8195);
and U11726 (N_11726,N_2355,N_9326);
and U11727 (N_11727,N_5474,N_9000);
and U11728 (N_11728,N_9628,N_6974);
nor U11729 (N_11729,N_3348,N_148);
or U11730 (N_11730,N_1745,N_498);
xor U11731 (N_11731,N_8518,N_9280);
and U11732 (N_11732,N_7178,N_7865);
and U11733 (N_11733,N_5428,N_169);
nor U11734 (N_11734,N_8909,N_7199);
and U11735 (N_11735,N_6101,N_7719);
or U11736 (N_11736,N_8085,N_717);
xnor U11737 (N_11737,N_691,N_7147);
xnor U11738 (N_11738,N_1104,N_3370);
or U11739 (N_11739,N_4149,N_1424);
xor U11740 (N_11740,N_4994,N_5654);
nand U11741 (N_11741,N_5631,N_8079);
xor U11742 (N_11742,N_2095,N_100);
xor U11743 (N_11743,N_4601,N_7620);
and U11744 (N_11744,N_9554,N_4666);
nor U11745 (N_11745,N_1246,N_6492);
xnor U11746 (N_11746,N_7496,N_1131);
or U11747 (N_11747,N_9918,N_7840);
or U11748 (N_11748,N_1232,N_6528);
or U11749 (N_11749,N_2561,N_5444);
or U11750 (N_11750,N_5711,N_1872);
nor U11751 (N_11751,N_4638,N_5100);
nor U11752 (N_11752,N_3893,N_3281);
or U11753 (N_11753,N_3401,N_3786);
xnor U11754 (N_11754,N_5497,N_8779);
nor U11755 (N_11755,N_3744,N_3458);
or U11756 (N_11756,N_2935,N_9553);
nand U11757 (N_11757,N_9873,N_232);
or U11758 (N_11758,N_8150,N_1322);
nor U11759 (N_11759,N_3952,N_1272);
and U11760 (N_11760,N_8708,N_274);
xor U11761 (N_11761,N_3073,N_2297);
nor U11762 (N_11762,N_653,N_6924);
nand U11763 (N_11763,N_995,N_2958);
xnor U11764 (N_11764,N_6065,N_4290);
nand U11765 (N_11765,N_2610,N_3183);
xor U11766 (N_11766,N_6526,N_6596);
and U11767 (N_11767,N_637,N_4308);
nand U11768 (N_11768,N_2519,N_7122);
nor U11769 (N_11769,N_3449,N_1282);
and U11770 (N_11770,N_3279,N_922);
and U11771 (N_11771,N_5232,N_3968);
nor U11772 (N_11772,N_606,N_4046);
nand U11773 (N_11773,N_5051,N_5795);
and U11774 (N_11774,N_4402,N_1829);
and U11775 (N_11775,N_4529,N_8570);
nor U11776 (N_11776,N_7197,N_1569);
xnor U11777 (N_11777,N_1135,N_9325);
nand U11778 (N_11778,N_7554,N_1414);
nand U11779 (N_11779,N_7364,N_5291);
and U11780 (N_11780,N_5878,N_3898);
nor U11781 (N_11781,N_8335,N_9772);
and U11782 (N_11782,N_730,N_317);
xnor U11783 (N_11783,N_4696,N_4972);
nand U11784 (N_11784,N_8976,N_3523);
nand U11785 (N_11785,N_1875,N_8643);
nand U11786 (N_11786,N_6434,N_9137);
nor U11787 (N_11787,N_4506,N_6583);
nor U11788 (N_11788,N_4352,N_5);
nand U11789 (N_11789,N_7466,N_2303);
nor U11790 (N_11790,N_9354,N_1351);
and U11791 (N_11791,N_3012,N_5572);
and U11792 (N_11792,N_835,N_4867);
or U11793 (N_11793,N_8532,N_8724);
nor U11794 (N_11794,N_2672,N_5689);
xnor U11795 (N_11795,N_8,N_9320);
and U11796 (N_11796,N_9523,N_9859);
xor U11797 (N_11797,N_9113,N_3427);
xnor U11798 (N_11798,N_3492,N_9450);
xnor U11799 (N_11799,N_1364,N_2313);
and U11800 (N_11800,N_6412,N_6827);
and U11801 (N_11801,N_4227,N_7025);
or U11802 (N_11802,N_3321,N_1581);
nand U11803 (N_11803,N_1451,N_3817);
or U11804 (N_11804,N_5022,N_6451);
nor U11805 (N_11805,N_838,N_3299);
nor U11806 (N_11806,N_2713,N_3262);
and U11807 (N_11807,N_2310,N_3787);
or U11808 (N_11808,N_4284,N_3165);
and U11809 (N_11809,N_4234,N_1969);
and U11810 (N_11810,N_9748,N_3117);
nor U11811 (N_11811,N_3978,N_5986);
xnor U11812 (N_11812,N_6833,N_3944);
xor U11813 (N_11813,N_5254,N_7319);
nor U11814 (N_11814,N_3143,N_7907);
or U11815 (N_11815,N_2917,N_7700);
or U11816 (N_11816,N_5077,N_8657);
or U11817 (N_11817,N_6577,N_5875);
nor U11818 (N_11818,N_4811,N_463);
or U11819 (N_11819,N_1547,N_832);
nor U11820 (N_11820,N_4700,N_3671);
and U11821 (N_11821,N_7027,N_526);
nor U11822 (N_11822,N_5062,N_8911);
and U11823 (N_11823,N_1368,N_5563);
or U11824 (N_11824,N_7104,N_939);
nor U11825 (N_11825,N_5448,N_9467);
nor U11826 (N_11826,N_5292,N_5423);
and U11827 (N_11827,N_3711,N_818);
and U11828 (N_11828,N_5615,N_9016);
nand U11829 (N_11829,N_660,N_4951);
and U11830 (N_11830,N_9722,N_3054);
xor U11831 (N_11831,N_1680,N_4948);
nand U11832 (N_11832,N_4005,N_3434);
and U11833 (N_11833,N_4815,N_8220);
or U11834 (N_11834,N_3585,N_6338);
nand U11835 (N_11835,N_3431,N_9824);
and U11836 (N_11836,N_496,N_5195);
xnor U11837 (N_11837,N_6230,N_1015);
and U11838 (N_11838,N_5267,N_5140);
nand U11839 (N_11839,N_6128,N_1958);
nand U11840 (N_11840,N_6219,N_5967);
or U11841 (N_11841,N_339,N_8380);
nand U11842 (N_11842,N_9396,N_6124);
nor U11843 (N_11843,N_1695,N_9402);
nand U11844 (N_11844,N_5194,N_3122);
xnor U11845 (N_11845,N_6718,N_5594);
or U11846 (N_11846,N_3644,N_1938);
nand U11847 (N_11847,N_700,N_4362);
nand U11848 (N_11848,N_9861,N_6433);
or U11849 (N_11849,N_2885,N_1835);
xnor U11850 (N_11850,N_386,N_983);
or U11851 (N_11851,N_720,N_2800);
and U11852 (N_11852,N_595,N_912);
and U11853 (N_11853,N_5258,N_7056);
or U11854 (N_11854,N_3550,N_8146);
and U11855 (N_11855,N_2883,N_8065);
nand U11856 (N_11856,N_9846,N_6876);
and U11857 (N_11857,N_8837,N_4206);
or U11858 (N_11858,N_7371,N_2529);
or U11859 (N_11859,N_2923,N_3180);
or U11860 (N_11860,N_5182,N_9228);
and U11861 (N_11861,N_5327,N_4961);
nor U11862 (N_11862,N_1669,N_8623);
nand U11863 (N_11863,N_2339,N_6419);
xor U11864 (N_11864,N_2178,N_4398);
and U11865 (N_11865,N_5799,N_6509);
xnor U11866 (N_11866,N_117,N_4182);
and U11867 (N_11867,N_4405,N_6418);
or U11868 (N_11868,N_1076,N_1383);
xor U11869 (N_11869,N_4543,N_6286);
nor U11870 (N_11870,N_2876,N_9546);
xnor U11871 (N_11871,N_6872,N_6014);
nand U11872 (N_11872,N_5328,N_4603);
and U11873 (N_11873,N_6898,N_7997);
or U11874 (N_11874,N_176,N_9507);
nand U11875 (N_11875,N_4914,N_5624);
nor U11876 (N_11876,N_462,N_7368);
xnor U11877 (N_11877,N_5674,N_486);
or U11878 (N_11878,N_2785,N_2038);
nor U11879 (N_11879,N_1117,N_9631);
nand U11880 (N_11880,N_476,N_8785);
and U11881 (N_11881,N_8758,N_6401);
nor U11882 (N_11882,N_9784,N_968);
nor U11883 (N_11883,N_391,N_8080);
nor U11884 (N_11884,N_3184,N_6031);
or U11885 (N_11885,N_7986,N_601);
nand U11886 (N_11886,N_1930,N_3597);
nor U11887 (N_11887,N_3702,N_9779);
and U11888 (N_11888,N_6731,N_9498);
and U11889 (N_11889,N_8246,N_388);
nand U11890 (N_11890,N_4459,N_8897);
xor U11891 (N_11891,N_5053,N_7529);
nand U11892 (N_11892,N_4197,N_3639);
and U11893 (N_11893,N_7029,N_1768);
nor U11894 (N_11894,N_70,N_4112);
xor U11895 (N_11895,N_9149,N_2830);
and U11896 (N_11896,N_1158,N_2518);
or U11897 (N_11897,N_3779,N_8903);
xor U11898 (N_11898,N_9405,N_6018);
nor U11899 (N_11899,N_2772,N_3887);
or U11900 (N_11900,N_3312,N_1598);
or U11901 (N_11901,N_3846,N_7588);
and U11902 (N_11902,N_4656,N_456);
or U11903 (N_11903,N_9906,N_3900);
and U11904 (N_11904,N_3632,N_967);
xnor U11905 (N_11905,N_1796,N_1006);
or U11906 (N_11906,N_5482,N_4231);
or U11907 (N_11907,N_6020,N_5272);
and U11908 (N_11908,N_2268,N_2283);
and U11909 (N_11909,N_593,N_3912);
xor U11910 (N_11910,N_3288,N_9351);
nor U11911 (N_11911,N_9344,N_9333);
xnor U11912 (N_11912,N_2824,N_1534);
nand U11913 (N_11913,N_9851,N_9587);
or U11914 (N_11914,N_7144,N_9516);
nand U11915 (N_11915,N_3957,N_4770);
xor U11916 (N_11916,N_4776,N_8373);
xor U11917 (N_11917,N_9455,N_5338);
and U11918 (N_11918,N_188,N_789);
or U11919 (N_11919,N_6759,N_6645);
xnor U11920 (N_11920,N_6688,N_7859);
xor U11921 (N_11921,N_8094,N_9304);
nor U11922 (N_11922,N_9676,N_4789);
nand U11923 (N_11923,N_1278,N_1613);
and U11924 (N_11924,N_2653,N_3164);
and U11925 (N_11925,N_5539,N_5528);
nand U11926 (N_11926,N_7434,N_8965);
and U11927 (N_11927,N_9816,N_8112);
and U11928 (N_11928,N_5736,N_4307);
or U11929 (N_11929,N_6343,N_3673);
xnor U11930 (N_11930,N_5364,N_8469);
nand U11931 (N_11931,N_1347,N_7446);
xor U11932 (N_11932,N_8352,N_7349);
nor U11933 (N_11933,N_4753,N_872);
and U11934 (N_11934,N_7695,N_6325);
or U11935 (N_11935,N_3544,N_4272);
xnor U11936 (N_11936,N_4909,N_8639);
nand U11937 (N_11937,N_9792,N_7453);
or U11938 (N_11938,N_9704,N_770);
nor U11939 (N_11939,N_668,N_6073);
and U11940 (N_11940,N_9893,N_9208);
or U11941 (N_11941,N_6304,N_5160);
nor U11942 (N_11942,N_1818,N_3852);
or U11943 (N_11943,N_4968,N_696);
and U11944 (N_11944,N_3820,N_4393);
nand U11945 (N_11945,N_5216,N_5928);
xnor U11946 (N_11946,N_8225,N_2690);
and U11947 (N_11947,N_6182,N_5121);
or U11948 (N_11948,N_9535,N_3956);
nor U11949 (N_11949,N_3792,N_5456);
xor U11950 (N_11950,N_6758,N_7437);
xor U11951 (N_11951,N_8361,N_2636);
and U11952 (N_11952,N_902,N_8210);
xnor U11953 (N_11953,N_7703,N_8133);
nor U11954 (N_11954,N_4429,N_8218);
nor U11955 (N_11955,N_2190,N_9352);
nor U11956 (N_11956,N_9916,N_384);
and U11957 (N_11957,N_4655,N_3543);
nor U11958 (N_11958,N_8743,N_9839);
nor U11959 (N_11959,N_6445,N_5587);
nor U11960 (N_11960,N_7731,N_14);
or U11961 (N_11961,N_2064,N_8261);
and U11962 (N_11962,N_4600,N_3488);
xor U11963 (N_11963,N_7458,N_3722);
and U11964 (N_11964,N_445,N_6442);
xnor U11965 (N_11965,N_6724,N_9091);
and U11966 (N_11966,N_6586,N_4304);
nand U11967 (N_11967,N_2768,N_1965);
xor U11968 (N_11968,N_5586,N_614);
xor U11969 (N_11969,N_8916,N_2002);
or U11970 (N_11970,N_9243,N_2961);
and U11971 (N_11971,N_3875,N_4121);
xnor U11972 (N_11972,N_4908,N_8494);
and U11973 (N_11973,N_9061,N_3357);
and U11974 (N_11974,N_6875,N_811);
xnor U11975 (N_11975,N_4792,N_2570);
nand U11976 (N_11976,N_7775,N_5425);
xnor U11977 (N_11977,N_3825,N_2591);
or U11978 (N_11978,N_9415,N_3751);
and U11979 (N_11979,N_8024,N_2200);
xor U11980 (N_11980,N_8473,N_9420);
or U11981 (N_11981,N_1708,N_5348);
xnor U11982 (N_11982,N_4520,N_6139);
xor U11983 (N_11983,N_6930,N_9673);
or U11984 (N_11984,N_9917,N_4026);
nand U11985 (N_11985,N_3035,N_9298);
xnor U11986 (N_11986,N_6911,N_9303);
nand U11987 (N_11987,N_6713,N_9819);
nor U11988 (N_11988,N_5393,N_225);
and U11989 (N_11989,N_1397,N_377);
or U11990 (N_11990,N_5313,N_5648);
xnor U11991 (N_11991,N_9919,N_7603);
nand U11992 (N_11992,N_7906,N_147);
nand U11993 (N_11993,N_4152,N_2581);
or U11994 (N_11994,N_4077,N_8664);
xnor U11995 (N_11995,N_1711,N_3064);
or U11996 (N_11996,N_3683,N_778);
nand U11997 (N_11997,N_8456,N_9955);
and U11998 (N_11998,N_4733,N_8866);
nor U11999 (N_11999,N_611,N_1903);
nand U12000 (N_12000,N_8055,N_2242);
or U12001 (N_12001,N_772,N_6836);
and U12002 (N_12002,N_3894,N_3063);
nor U12003 (N_12003,N_8910,N_8874);
nor U12004 (N_12004,N_6047,N_9290);
xor U12005 (N_12005,N_5699,N_8681);
or U12006 (N_12006,N_6667,N_5732);
and U12007 (N_12007,N_909,N_3447);
and U12008 (N_12008,N_2014,N_4924);
nor U12009 (N_12009,N_5370,N_1970);
nand U12010 (N_12010,N_2112,N_2635);
nor U12011 (N_12011,N_2563,N_2048);
or U12012 (N_12012,N_3616,N_3182);
or U12013 (N_12013,N_6022,N_8595);
or U12014 (N_12014,N_1657,N_6889);
xor U12015 (N_12015,N_6502,N_4954);
or U12016 (N_12016,N_3392,N_5136);
nor U12017 (N_12017,N_6340,N_9357);
or U12018 (N_12018,N_2754,N_3903);
or U12019 (N_12019,N_9395,N_7877);
and U12020 (N_12020,N_8271,N_4333);
nand U12021 (N_12021,N_9798,N_3642);
nand U12022 (N_12022,N_485,N_7832);
xor U12023 (N_12023,N_6792,N_6489);
nor U12024 (N_12024,N_2069,N_4683);
xor U12025 (N_12025,N_2963,N_8953);
and U12026 (N_12026,N_4283,N_896);
nor U12027 (N_12027,N_2125,N_1576);
xor U12028 (N_12028,N_5045,N_8817);
nor U12029 (N_12029,N_2221,N_5223);
nor U12030 (N_12030,N_6900,N_4541);
or U12031 (N_12031,N_7367,N_2879);
nand U12032 (N_12032,N_3020,N_44);
nor U12033 (N_12033,N_9692,N_1107);
and U12034 (N_12034,N_1666,N_2596);
or U12035 (N_12035,N_7599,N_9961);
or U12036 (N_12036,N_2985,N_3773);
nor U12037 (N_12037,N_5527,N_8073);
xnor U12038 (N_12038,N_7715,N_420);
nand U12039 (N_12039,N_1277,N_5118);
nand U12040 (N_12040,N_7569,N_3380);
xor U12041 (N_12041,N_72,N_2176);
nand U12042 (N_12042,N_5079,N_1161);
nand U12043 (N_12043,N_6113,N_2954);
nor U12044 (N_12044,N_8431,N_5633);
nor U12045 (N_12045,N_6099,N_4054);
and U12046 (N_12046,N_260,N_2151);
and U12047 (N_12047,N_6271,N_632);
or U12048 (N_12048,N_6361,N_1270);
or U12049 (N_12049,N_1668,N_9557);
or U12050 (N_12050,N_8914,N_1199);
and U12051 (N_12051,N_7213,N_4871);
nand U12052 (N_12052,N_3637,N_416);
nor U12053 (N_12053,N_2649,N_2428);
nor U12054 (N_12054,N_7548,N_7084);
and U12055 (N_12055,N_6036,N_5235);
and U12056 (N_12056,N_560,N_9857);
nand U12057 (N_12057,N_3009,N_7167);
or U12058 (N_12058,N_5790,N_9488);
or U12059 (N_12059,N_7394,N_6782);
and U12060 (N_12060,N_8408,N_675);
and U12061 (N_12061,N_2273,N_158);
nand U12062 (N_12062,N_2565,N_8748);
or U12063 (N_12063,N_3542,N_5782);
nand U12064 (N_12064,N_7782,N_5990);
and U12065 (N_12065,N_6881,N_5599);
nand U12066 (N_12066,N_6255,N_8404);
or U12067 (N_12067,N_3405,N_7682);
and U12068 (N_12068,N_5952,N_8214);
nor U12069 (N_12069,N_4524,N_828);
xnor U12070 (N_12070,N_4960,N_6576);
and U12071 (N_12071,N_7410,N_7317);
nand U12072 (N_12072,N_3224,N_8898);
nand U12073 (N_12073,N_5305,N_353);
or U12074 (N_12074,N_6300,N_9530);
or U12075 (N_12075,N_3399,N_9400);
and U12076 (N_12076,N_4226,N_1111);
nor U12077 (N_12077,N_4641,N_8090);
nand U12078 (N_12078,N_4899,N_7001);
nor U12079 (N_12079,N_1309,N_3810);
xor U12080 (N_12080,N_5742,N_3315);
or U12081 (N_12081,N_9699,N_1507);
nand U12082 (N_12082,N_2006,N_6197);
nor U12083 (N_12083,N_4154,N_5477);
or U12084 (N_12084,N_5383,N_9949);
nand U12085 (N_12085,N_6611,N_3858);
nand U12086 (N_12086,N_1604,N_3033);
xnor U12087 (N_12087,N_9431,N_4192);
and U12088 (N_12088,N_1370,N_6092);
nor U12089 (N_12089,N_1722,N_1425);
nor U12090 (N_12090,N_8191,N_5402);
nor U12091 (N_12091,N_1787,N_1372);
nand U12092 (N_12092,N_7405,N_8789);
nand U12093 (N_12093,N_8312,N_2280);
and U12094 (N_12094,N_4885,N_1687);
xnor U12095 (N_12095,N_7726,N_2583);
or U12096 (N_12096,N_6821,N_9356);
xor U12097 (N_12097,N_5239,N_2530);
xor U12098 (N_12098,N_1055,N_2521);
nand U12099 (N_12099,N_7990,N_8338);
and U12100 (N_12100,N_6406,N_3049);
and U12101 (N_12101,N_9013,N_545);
nor U12102 (N_12102,N_2980,N_8918);
or U12103 (N_12103,N_2111,N_6263);
or U12104 (N_12104,N_4014,N_9093);
or U12105 (N_12105,N_763,N_4476);
nand U12106 (N_12106,N_7777,N_2469);
or U12107 (N_12107,N_9260,N_973);
xnor U12108 (N_12108,N_3532,N_6493);
nor U12109 (N_12109,N_2174,N_3456);
and U12110 (N_12110,N_2753,N_1290);
xor U12111 (N_12111,N_9680,N_1016);
nand U12112 (N_12112,N_8548,N_9708);
or U12113 (N_12113,N_6310,N_3680);
xor U12114 (N_12114,N_9607,N_7389);
or U12115 (N_12115,N_518,N_5524);
nor U12116 (N_12116,N_2088,N_2422);
xnor U12117 (N_12117,N_1989,N_3728);
xnor U12118 (N_12118,N_4044,N_1959);
xnor U12119 (N_12119,N_8399,N_6322);
nand U12120 (N_12120,N_7076,N_4732);
nand U12121 (N_12121,N_2488,N_7238);
nor U12122 (N_12122,N_8746,N_9742);
and U12123 (N_12123,N_6803,N_743);
and U12124 (N_12124,N_422,N_2562);
or U12125 (N_12125,N_6585,N_9937);
nand U12126 (N_12126,N_4494,N_2840);
nor U12127 (N_12127,N_8812,N_3724);
or U12128 (N_12128,N_4781,N_8474);
or U12129 (N_12129,N_2559,N_5065);
nand U12130 (N_12130,N_7991,N_9027);
nand U12131 (N_12131,N_9870,N_6868);
xnor U12132 (N_12132,N_5395,N_859);
nor U12133 (N_12133,N_4605,N_1214);
xor U12134 (N_12134,N_4740,N_7573);
and U12135 (N_12135,N_6491,N_5868);
nand U12136 (N_12136,N_414,N_4027);
or U12137 (N_12137,N_7086,N_7953);
nand U12138 (N_12138,N_8560,N_8078);
nor U12139 (N_12139,N_1817,N_7066);
or U12140 (N_12140,N_8522,N_1152);
nand U12141 (N_12141,N_7562,N_9726);
nor U12142 (N_12142,N_3897,N_9559);
nand U12143 (N_12143,N_3804,N_8505);
nand U12144 (N_12144,N_5760,N_6386);
and U12145 (N_12145,N_2209,N_6000);
and U12146 (N_12146,N_6838,N_1988);
xnor U12147 (N_12147,N_6308,N_3107);
nor U12148 (N_12148,N_7752,N_7743);
or U12149 (N_12149,N_9339,N_9963);
or U12150 (N_12150,N_8762,N_1819);
xnor U12151 (N_12151,N_587,N_332);
or U12152 (N_12152,N_5315,N_4624);
nand U12153 (N_12153,N_3789,N_8208);
xor U12154 (N_12154,N_6474,N_2495);
and U12155 (N_12155,N_6111,N_3545);
or U12156 (N_12156,N_9469,N_9749);
xnor U12157 (N_12157,N_3872,N_7851);
and U12158 (N_12158,N_5605,N_3878);
nor U12159 (N_12159,N_9793,N_251);
and U12160 (N_12160,N_3263,N_211);
or U12161 (N_12161,N_6284,N_6356);
nand U12162 (N_12162,N_8802,N_3069);
nor U12163 (N_12163,N_3831,N_8051);
nor U12164 (N_12164,N_8757,N_6908);
nor U12165 (N_12165,N_2493,N_6518);
nand U12166 (N_12166,N_1201,N_4708);
nor U12167 (N_12167,N_1764,N_2180);
and U12168 (N_12168,N_8924,N_1909);
nand U12169 (N_12169,N_6970,N_489);
nor U12170 (N_12170,N_5405,N_3890);
nand U12171 (N_12171,N_3966,N_1120);
and U12172 (N_12172,N_9452,N_8938);
or U12173 (N_12173,N_9998,N_5515);
or U12174 (N_12174,N_6289,N_4099);
xor U12175 (N_12175,N_3160,N_9273);
nor U12176 (N_12176,N_3742,N_1093);
and U12177 (N_12177,N_7607,N_9127);
xnor U12178 (N_12178,N_1993,N_5763);
and U12179 (N_12179,N_2500,N_8540);
or U12180 (N_12180,N_7153,N_8701);
or U12181 (N_12181,N_3236,N_704);
xor U12182 (N_12182,N_1624,N_5099);
or U12183 (N_12183,N_1486,N_2760);
nand U12184 (N_12184,N_7375,N_2682);
nor U12185 (N_12185,N_6591,N_5940);
xor U12186 (N_12186,N_6736,N_9098);
nor U12187 (N_12187,N_5597,N_6399);
xor U12188 (N_12188,N_1243,N_9809);
or U12189 (N_12189,N_3151,N_7557);
or U12190 (N_12190,N_1013,N_8053);
and U12191 (N_12191,N_5510,N_946);
nor U12192 (N_12192,N_9496,N_8783);
nand U12193 (N_12193,N_454,N_2413);
or U12194 (N_12194,N_6075,N_3204);
nor U12195 (N_12195,N_4509,N_8618);
nand U12196 (N_12196,N_7037,N_501);
and U12197 (N_12197,N_4313,N_3474);
or U12198 (N_12198,N_9730,N_5585);
nor U12199 (N_12199,N_1977,N_9348);
nor U12200 (N_12200,N_2532,N_5431);
nand U12201 (N_12201,N_4640,N_6721);
and U12202 (N_12202,N_4247,N_6402);
or U12203 (N_12203,N_5187,N_4680);
xor U12204 (N_12204,N_7430,N_1437);
or U12205 (N_12205,N_6793,N_898);
nor U12206 (N_12206,N_3785,N_3161);
or U12207 (N_12207,N_9986,N_6789);
nor U12208 (N_12208,N_8555,N_1900);
xnor U12209 (N_12209,N_9573,N_2161);
nand U12210 (N_12210,N_6196,N_7511);
nand U12211 (N_12211,N_2306,N_520);
and U12212 (N_12212,N_7429,N_4838);
xor U12213 (N_12213,N_1692,N_825);
xnor U12214 (N_12214,N_3910,N_2967);
or U12215 (N_12215,N_2755,N_9745);
and U12216 (N_12216,N_9244,N_2059);
or U12217 (N_12217,N_5562,N_8365);
or U12218 (N_12218,N_4658,N_7140);
nor U12219 (N_12219,N_8588,N_6496);
nor U12220 (N_12220,N_719,N_6755);
and U12221 (N_12221,N_5985,N_5821);
xor U12222 (N_12222,N_7869,N_5975);
nand U12223 (N_12223,N_943,N_5218);
nor U12224 (N_12224,N_3884,N_4574);
or U12225 (N_12225,N_6058,N_6126);
nor U12226 (N_12226,N_2953,N_2166);
xnor U12227 (N_12227,N_4173,N_1431);
and U12228 (N_12228,N_257,N_4653);
nor U12229 (N_12229,N_8539,N_3612);
and U12230 (N_12230,N_444,N_4203);
xor U12231 (N_12231,N_4652,N_4047);
xor U12232 (N_12232,N_4327,N_1024);
or U12233 (N_12233,N_1554,N_1706);
nand U12234 (N_12234,N_5176,N_9074);
and U12235 (N_12235,N_3435,N_3088);
xor U12236 (N_12236,N_8159,N_9211);
or U12237 (N_12237,N_4895,N_6992);
or U12238 (N_12238,N_8955,N_6680);
xor U12239 (N_12239,N_2390,N_3451);
nand U12240 (N_12240,N_7305,N_1778);
nand U12241 (N_12241,N_7152,N_4940);
nor U12242 (N_12242,N_4970,N_9562);
xnor U12243 (N_12243,N_3052,N_8794);
nor U12244 (N_12244,N_5496,N_7222);
and U12245 (N_12245,N_8202,N_7582);
or U12246 (N_12246,N_5817,N_5185);
and U12247 (N_12247,N_3636,N_790);
nor U12248 (N_12248,N_7469,N_1655);
or U12249 (N_12249,N_3374,N_5189);
or U12250 (N_12250,N_5672,N_7613);
xnor U12251 (N_12251,N_8184,N_1891);
nand U12252 (N_12252,N_6158,N_2813);
nand U12253 (N_12253,N_8862,N_9078);
nor U12254 (N_12254,N_1640,N_5621);
xnor U12255 (N_12255,N_7075,N_5765);
nand U12256 (N_12256,N_4299,N_2067);
xnor U12257 (N_12257,N_1133,N_7763);
xnor U12258 (N_12258,N_8513,N_7230);
or U12259 (N_12259,N_8437,N_6507);
or U12260 (N_12260,N_3108,N_5404);
or U12261 (N_12261,N_4883,N_9747);
nand U12262 (N_12262,N_5590,N_9157);
xor U12263 (N_12263,N_7221,N_9690);
or U12264 (N_12264,N_3082,N_3422);
xnor U12265 (N_12265,N_3808,N_7287);
nor U12266 (N_12266,N_6016,N_2016);
nor U12267 (N_12267,N_5209,N_8507);
nor U12268 (N_12268,N_3943,N_6834);
nor U12269 (N_12269,N_4030,N_6622);
or U12270 (N_12270,N_1832,N_9358);
nand U12271 (N_12271,N_5955,N_5473);
xnor U12272 (N_12272,N_5676,N_1455);
or U12273 (N_12273,N_7706,N_2865);
xnor U12274 (N_12274,N_4525,N_3166);
or U12275 (N_12275,N_2246,N_9283);
nand U12276 (N_12276,N_9319,N_8318);
or U12277 (N_12277,N_7477,N_2880);
xnor U12278 (N_12278,N_1365,N_1978);
xnor U12279 (N_12279,N_2342,N_9201);
nor U12280 (N_12280,N_837,N_7708);
nand U12281 (N_12281,N_6318,N_2802);
nor U12282 (N_12282,N_9483,N_4379);
xor U12283 (N_12283,N_8302,N_8990);
or U12284 (N_12284,N_1878,N_1310);
nor U12285 (N_12285,N_4595,N_1109);
or U12286 (N_12286,N_2039,N_9241);
nand U12287 (N_12287,N_7377,N_2741);
nand U12288 (N_12288,N_4277,N_914);
nand U12289 (N_12289,N_7593,N_5937);
or U12290 (N_12290,N_7993,N_73);
and U12291 (N_12291,N_8713,N_6903);
xnor U12292 (N_12292,N_8303,N_8564);
or U12293 (N_12293,N_861,N_8896);
and U12294 (N_12294,N_10,N_8311);
xnor U12295 (N_12295,N_9124,N_5427);
or U12296 (N_12296,N_7894,N_2430);
or U12297 (N_12297,N_9826,N_2047);
nand U12298 (N_12298,N_1517,N_2239);
nor U12299 (N_12299,N_7498,N_6129);
or U12300 (N_12300,N_7281,N_8209);
xnor U12301 (N_12301,N_9813,N_9548);
nand U12302 (N_12302,N_2855,N_7309);
or U12303 (N_12303,N_4438,N_1458);
nand U12304 (N_12304,N_3394,N_1229);
or U12305 (N_12305,N_8731,N_1148);
nand U12306 (N_12306,N_3018,N_1676);
nand U12307 (N_12307,N_1532,N_8650);
nor U12308 (N_12308,N_3385,N_8768);
nand U12309 (N_12309,N_9872,N_4473);
or U12310 (N_12310,N_850,N_2265);
nor U12311 (N_12311,N_5837,N_2394);
nand U12312 (N_12312,N_9755,N_9735);
xor U12313 (N_12313,N_7830,N_3718);
and U12314 (N_12314,N_4575,N_3113);
nor U12315 (N_12315,N_7284,N_6524);
nand U12316 (N_12316,N_8277,N_5947);
xor U12317 (N_12317,N_8838,N_7174);
nand U12318 (N_12318,N_2063,N_3733);
xor U12319 (N_12319,N_3455,N_3232);
and U12320 (N_12320,N_2036,N_5461);
or U12321 (N_12321,N_8635,N_2947);
or U12322 (N_12322,N_5247,N_8658);
nand U12323 (N_12323,N_8267,N_5122);
xor U12324 (N_12324,N_8041,N_1333);
or U12325 (N_12325,N_1492,N_3381);
nor U12326 (N_12326,N_6990,N_1990);
or U12327 (N_12327,N_5503,N_5277);
nor U12328 (N_12328,N_6639,N_4216);
nand U12329 (N_12329,N_4334,N_5200);
or U12330 (N_12330,N_1984,N_3003);
nor U12331 (N_12331,N_3682,N_588);
and U12332 (N_12332,N_1559,N_6651);
or U12333 (N_12333,N_7138,N_8674);
nand U12334 (N_12334,N_6427,N_8447);
xnor U12335 (N_12335,N_6027,N_272);
xor U12336 (N_12336,N_1146,N_4279);
or U12337 (N_12337,N_3692,N_3643);
nand U12338 (N_12338,N_686,N_7764);
nor U12339 (N_12339,N_1950,N_6161);
nor U12340 (N_12340,N_7995,N_7612);
or U12341 (N_12341,N_9438,N_4294);
nand U12342 (N_12342,N_3605,N_2734);
and U12343 (N_12343,N_7568,N_7136);
or U12344 (N_12344,N_9481,N_9621);
nand U12345 (N_12345,N_6561,N_9595);
and U12346 (N_12346,N_2918,N_4181);
nor U12347 (N_12347,N_4093,N_5015);
or U12348 (N_12348,N_3735,N_5098);
and U12349 (N_12349,N_3958,N_7671);
or U12350 (N_12350,N_1784,N_9447);
or U12351 (N_12351,N_3127,N_5776);
nor U12352 (N_12352,N_1288,N_6469);
or U12353 (N_12353,N_7518,N_519);
nor U12354 (N_12354,N_6695,N_5813);
and U12355 (N_12355,N_7809,N_5476);
xnor U12356 (N_12356,N_9744,N_6804);
and U12357 (N_12357,N_7841,N_4423);
nor U12358 (N_12358,N_3541,N_4363);
xor U12359 (N_12359,N_9434,N_4111);
nor U12360 (N_12360,N_259,N_8803);
or U12361 (N_12361,N_9151,N_4938);
and U12362 (N_12362,N_4554,N_396);
nand U12363 (N_12363,N_6074,N_4665);
xnor U12364 (N_12364,N_2158,N_9026);
and U12365 (N_12365,N_9182,N_3147);
xor U12366 (N_12366,N_1386,N_7938);
nand U12367 (N_12367,N_5308,N_6029);
nand U12368 (N_12368,N_121,N_1661);
xnor U12369 (N_12369,N_950,N_85);
or U12370 (N_12370,N_8047,N_1238);
xnor U12371 (N_12371,N_9183,N_2810);
nand U12372 (N_12372,N_4467,N_6769);
nor U12373 (N_12373,N_3305,N_7441);
xor U12374 (N_12374,N_8098,N_244);
xor U12375 (N_12375,N_9397,N_3328);
and U12376 (N_12376,N_5862,N_6168);
xor U12377 (N_12377,N_7697,N_4375);
and U12378 (N_12378,N_8946,N_8487);
and U12379 (N_12379,N_2361,N_1144);
or U12380 (N_12380,N_58,N_5637);
and U12381 (N_12381,N_7699,N_7077);
nor U12382 (N_12382,N_5926,N_3156);
xor U12383 (N_12383,N_5199,N_8880);
nor U12384 (N_12384,N_8951,N_2077);
nand U12385 (N_12385,N_6467,N_6249);
nand U12386 (N_12386,N_5623,N_7154);
and U12387 (N_12387,N_8442,N_690);
xor U12388 (N_12388,N_1864,N_5622);
or U12389 (N_12389,N_6244,N_7210);
xnor U12390 (N_12390,N_3995,N_554);
nand U12391 (N_12391,N_4926,N_7766);
nand U12392 (N_12392,N_1916,N_8314);
or U12393 (N_12393,N_9188,N_8895);
xnor U12394 (N_12394,N_7884,N_1049);
or U12395 (N_12395,N_8920,N_7994);
nor U12396 (N_12396,N_921,N_4265);
xor U12397 (N_12397,N_4552,N_8162);
nor U12398 (N_12398,N_3462,N_7637);
and U12399 (N_12399,N_1222,N_2945);
or U12400 (N_12400,N_3672,N_9733);
nand U12401 (N_12401,N_1513,N_9161);
nand U12402 (N_12402,N_1915,N_6348);
and U12403 (N_12403,N_9046,N_4735);
and U12404 (N_12404,N_2406,N_3214);
nor U12405 (N_12405,N_8138,N_110);
and U12406 (N_12406,N_5408,N_5797);
nor U12407 (N_12407,N_827,N_2322);
and U12408 (N_12408,N_9355,N_3366);
nand U12409 (N_12409,N_4762,N_3141);
and U12410 (N_12410,N_5761,N_9202);
nor U12411 (N_12411,N_5339,N_4325);
nand U12412 (N_12412,N_1292,N_1795);
nor U12413 (N_12413,N_8247,N_7098);
nand U12414 (N_12414,N_6510,N_1780);
nor U12415 (N_12415,N_994,N_1099);
and U12416 (N_12416,N_8619,N_4947);
xnor U12417 (N_12417,N_1912,N_9649);
and U12418 (N_12418,N_6506,N_5886);
or U12419 (N_12419,N_8491,N_6720);
or U12420 (N_12420,N_7676,N_4291);
and U12421 (N_12421,N_6455,N_8192);
nor U12422 (N_12422,N_779,N_5526);
nor U12423 (N_12423,N_3338,N_6138);
and U12424 (N_12424,N_96,N_7640);
nor U12425 (N_12425,N_7464,N_9258);
nor U12426 (N_12426,N_2102,N_9443);
and U12427 (N_12427,N_4465,N_5974);
or U12428 (N_12428,N_1583,N_1741);
nor U12429 (N_12429,N_1505,N_3799);
nor U12430 (N_12430,N_4877,N_8917);
xnor U12431 (N_12431,N_5771,N_8439);
and U12432 (N_12432,N_2120,N_4810);
nand U12433 (N_12433,N_3463,N_2374);
xnor U12434 (N_12434,N_1060,N_6855);
or U12435 (N_12435,N_524,N_8864);
or U12436 (N_12436,N_6283,N_7691);
xor U12437 (N_12437,N_1009,N_8612);
nor U12438 (N_12438,N_3551,N_3946);
nand U12439 (N_12439,N_8446,N_7460);
nand U12440 (N_12440,N_1791,N_3854);
xnor U12441 (N_12441,N_6360,N_5485);
or U12442 (N_12442,N_2716,N_1568);
and U12443 (N_12443,N_7069,N_3763);
and U12444 (N_12444,N_1388,N_4178);
or U12445 (N_12445,N_1342,N_429);
nand U12446 (N_12446,N_8498,N_9890);
xnor U12447 (N_12447,N_9988,N_4748);
nand U12448 (N_12448,N_6777,N_6088);
or U12449 (N_12449,N_6037,N_9909);
nand U12450 (N_12450,N_1879,N_6747);
or U12451 (N_12451,N_2162,N_7206);
nand U12452 (N_12452,N_6234,N_8622);
and U12453 (N_12453,N_5659,N_3470);
nor U12454 (N_12454,N_3404,N_7891);
nand U12455 (N_12455,N_723,N_7041);
nand U12456 (N_12456,N_6376,N_3871);
nor U12457 (N_12457,N_9510,N_7962);
nand U12458 (N_12458,N_200,N_7646);
or U12459 (N_12459,N_1736,N_5710);
nand U12460 (N_12460,N_1785,N_7566);
xor U12461 (N_12461,N_269,N_344);
nand U12462 (N_12462,N_8722,N_1409);
nor U12463 (N_12463,N_3096,N_7159);
nand U12464 (N_12464,N_9213,N_8617);
xor U12465 (N_12465,N_1527,N_4193);
nor U12466 (N_12466,N_1597,N_4774);
or U12467 (N_12467,N_5781,N_3557);
nand U12468 (N_12468,N_6869,N_610);
and U12469 (N_12469,N_1923,N_6839);
or U12470 (N_12470,N_4345,N_8581);
and U12471 (N_12471,N_241,N_8957);
or U12472 (N_12472,N_7515,N_431);
or U12473 (N_12473,N_2815,N_8187);
nand U12474 (N_12474,N_6706,N_8005);
or U12475 (N_12475,N_5703,N_2642);
nor U12476 (N_12476,N_3429,N_2309);
nand U12477 (N_12477,N_2619,N_9384);
or U12478 (N_12478,N_649,N_1894);
nand U12479 (N_12479,N_4565,N_4869);
and U12480 (N_12480,N_1137,N_3059);
nand U12481 (N_12481,N_7878,N_1756);
nand U12482 (N_12482,N_449,N_9261);
nand U12483 (N_12483,N_2604,N_3369);
or U12484 (N_12484,N_3698,N_6148);
nor U12485 (N_12485,N_7014,N_9341);
or U12486 (N_12486,N_2999,N_7059);
xnor U12487 (N_12487,N_9926,N_8543);
nor U12488 (N_12488,N_9788,N_1378);
and U12489 (N_12489,N_4281,N_381);
or U12490 (N_12490,N_6701,N_6704);
nand U12491 (N_12491,N_7207,N_1315);
nand U12492 (N_12492,N_3769,N_6488);
xor U12493 (N_12493,N_7396,N_5857);
and U12494 (N_12494,N_4110,N_2216);
and U12495 (N_12495,N_3112,N_3466);
or U12496 (N_12496,N_8239,N_3798);
nor U12497 (N_12497,N_9033,N_2994);
nor U12498 (N_12498,N_3116,N_2618);
xor U12499 (N_12499,N_6156,N_5764);
nand U12500 (N_12500,N_2783,N_4136);
or U12501 (N_12501,N_3344,N_1590);
nand U12502 (N_12502,N_5803,N_3124);
and U12503 (N_12503,N_9212,N_4615);
nor U12504 (N_12504,N_3705,N_4135);
nor U12505 (N_12505,N_5248,N_673);
nor U12506 (N_12506,N_3042,N_3215);
nor U12507 (N_12507,N_8433,N_4555);
nor U12508 (N_12508,N_8987,N_159);
nand U12509 (N_12509,N_128,N_6751);
or U12510 (N_12510,N_5264,N_5454);
or U12511 (N_12511,N_8799,N_5536);
nand U12512 (N_12512,N_6254,N_9199);
nand U12513 (N_12513,N_9406,N_8849);
nor U12514 (N_12514,N_368,N_4038);
nor U12515 (N_12515,N_2032,N_1667);
or U12516 (N_12516,N_7082,N_7119);
or U12517 (N_12517,N_3237,N_7744);
xor U12518 (N_12518,N_5228,N_4890);
nor U12519 (N_12519,N_8254,N_2206);
nor U12520 (N_12520,N_6067,N_7156);
nand U12521 (N_12521,N_1031,N_1325);
xnor U12522 (N_12522,N_9070,N_3144);
and U12523 (N_12523,N_6953,N_4878);
nor U12524 (N_12524,N_4351,N_9602);
or U12525 (N_12525,N_229,N_3363);
nand U12526 (N_12526,N_3200,N_9815);
nor U12527 (N_12527,N_4255,N_7641);
xor U12528 (N_12528,N_6871,N_1975);
xor U12529 (N_12529,N_8956,N_4430);
nand U12530 (N_12530,N_9460,N_8500);
xor U12531 (N_12531,N_5896,N_7081);
or U12532 (N_12532,N_1165,N_9844);
xor U12533 (N_12533,N_4800,N_9756);
nor U12534 (N_12534,N_1698,N_1284);
and U12535 (N_12535,N_5946,N_5916);
and U12536 (N_12536,N_8787,N_8362);
or U12537 (N_12537,N_267,N_8902);
and U12538 (N_12538,N_464,N_7036);
xor U12539 (N_12539,N_9822,N_4250);
or U12540 (N_12540,N_5259,N_4661);
nand U12541 (N_12541,N_9952,N_3750);
or U12542 (N_12542,N_3038,N_2348);
or U12543 (N_12543,N_2416,N_1326);
xor U12544 (N_12544,N_4688,N_1048);
or U12545 (N_12545,N_8397,N_4404);
nor U12546 (N_12546,N_5335,N_1225);
nor U12547 (N_12547,N_2914,N_3748);
or U12548 (N_12548,N_2707,N_1184);
nor U12549 (N_12549,N_6548,N_8720);
xor U12550 (N_12550,N_2198,N_5343);
nand U12551 (N_12551,N_3359,N_3334);
nand U12552 (N_12552,N_1393,N_8649);
nand U12553 (N_12553,N_447,N_1421);
and U12554 (N_12554,N_7316,N_2534);
or U12555 (N_12555,N_8792,N_2884);
and U12556 (N_12556,N_724,N_1895);
nor U12557 (N_12557,N_6312,N_5991);
nand U12558 (N_12558,N_955,N_7915);
or U12559 (N_12559,N_6365,N_552);
nor U12560 (N_12560,N_6186,N_4912);
and U12561 (N_12561,N_1230,N_6486);
nor U12562 (N_12562,N_8497,N_4583);
nor U12563 (N_12563,N_4690,N_3251);
or U12564 (N_12564,N_2506,N_4486);
and U12565 (N_12565,N_1311,N_2075);
or U12566 (N_12566,N_2956,N_7095);
or U12567 (N_12567,N_9928,N_4131);
nor U12568 (N_12568,N_4377,N_2267);
xnor U12569 (N_12569,N_6498,N_1471);
nand U12570 (N_12570,N_1994,N_6171);
and U12571 (N_12571,N_7622,N_3841);
and U12572 (N_12572,N_187,N_5014);
nand U12573 (N_12573,N_8877,N_6100);
and U12574 (N_12574,N_2706,N_2480);
nor U12575 (N_12575,N_5651,N_1992);
or U12576 (N_12576,N_951,N_7857);
nor U12577 (N_12577,N_2318,N_8169);
nand U12578 (N_12578,N_2349,N_6238);
nand U12579 (N_12579,N_8807,N_731);
xor U12580 (N_12580,N_2266,N_8824);
nor U12581 (N_12581,N_8032,N_7020);
nor U12582 (N_12582,N_7784,N_1168);
nand U12583 (N_12583,N_5142,N_1063);
or U12584 (N_12584,N_3274,N_5048);
or U12585 (N_12585,N_6508,N_6484);
xnor U12586 (N_12586,N_7992,N_7301);
or U12587 (N_12587,N_6328,N_9868);
and U12588 (N_12588,N_2226,N_3687);
and U12589 (N_12589,N_9681,N_8460);
and U12590 (N_12590,N_3546,N_4500);
and U12591 (N_12591,N_7602,N_6250);
or U12592 (N_12592,N_8786,N_5005);
or U12593 (N_12593,N_6627,N_3706);
or U12594 (N_12594,N_9946,N_6638);
xnor U12595 (N_12595,N_4995,N_5618);
and U12596 (N_12596,N_5650,N_3391);
or U12597 (N_12597,N_7391,N_4210);
xnor U12598 (N_12598,N_8672,N_873);
or U12599 (N_12599,N_6081,N_619);
nor U12600 (N_12600,N_2863,N_8568);
xor U12601 (N_12601,N_9154,N_1809);
or U12602 (N_12602,N_2558,N_1897);
xnor U12603 (N_12603,N_9836,N_5649);
or U12604 (N_12604,N_7510,N_2640);
xor U12605 (N_12605,N_1276,N_5737);
and U12606 (N_12606,N_6581,N_6503);
nand U12607 (N_12607,N_2805,N_7336);
xor U12608 (N_12608,N_6925,N_7000);
xor U12609 (N_12609,N_9131,N_9577);
or U12610 (N_12610,N_6565,N_2177);
xnor U12611 (N_12611,N_7512,N_4085);
nor U12612 (N_12612,N_1866,N_3397);
or U12613 (N_12613,N_4189,N_8153);
or U12614 (N_12614,N_7141,N_1946);
nand U12615 (N_12615,N_8759,N_9623);
and U12616 (N_12616,N_7870,N_313);
or U12617 (N_12617,N_9863,N_1022);
and U12618 (N_12618,N_4664,N_3547);
nor U12619 (N_12619,N_8954,N_3525);
or U12620 (N_12620,N_4267,N_805);
nand U12621 (N_12621,N_9588,N_1088);
xnor U12622 (N_12622,N_5178,N_8493);
xnor U12623 (N_12623,N_4123,N_5389);
xnor U12624 (N_12624,N_2385,N_9386);
nor U12625 (N_12625,N_2560,N_1354);
and U12626 (N_12626,N_7929,N_5441);
xor U12627 (N_12627,N_9295,N_1308);
or U12628 (N_12628,N_4633,N_8511);
nor U12629 (N_12629,N_2279,N_823);
and U12630 (N_12630,N_8219,N_9930);
xor U12631 (N_12631,N_636,N_7108);
nand U12632 (N_12632,N_5257,N_2442);
xor U12633 (N_12633,N_8315,N_7750);
xor U12634 (N_12634,N_5429,N_3864);
nand U12635 (N_12635,N_848,N_7047);
and U12636 (N_12636,N_6083,N_1880);
or U12637 (N_12637,N_1174,N_54);
and U12638 (N_12638,N_9317,N_26);
xnor U12639 (N_12639,N_2414,N_1164);
or U12640 (N_12640,N_3527,N_6795);
nor U12641 (N_12641,N_701,N_4904);
nor U12642 (N_12642,N_2487,N_5457);
xor U12643 (N_12643,N_9171,N_8466);
or U12644 (N_12644,N_1500,N_5440);
nor U12645 (N_12645,N_6873,N_8403);
xnor U12646 (N_12646,N_1082,N_4798);
nor U12647 (N_12647,N_7246,N_4137);
nand U12648 (N_12648,N_9657,N_4407);
xor U12649 (N_12649,N_5041,N_4338);
xor U12650 (N_12650,N_5854,N_1043);
xnor U12651 (N_12651,N_3208,N_6629);
or U12652 (N_12652,N_9987,N_5682);
and U12653 (N_12653,N_8992,N_7312);
xor U12654 (N_12654,N_3244,N_1296);
nor U12655 (N_12655,N_4105,N_689);
nand U12656 (N_12656,N_8406,N_8105);
nor U12657 (N_12657,N_5979,N_3487);
nand U12658 (N_12658,N_1684,N_1983);
nand U12659 (N_12659,N_9004,N_7175);
or U12660 (N_12660,N_7229,N_3097);
and U12661 (N_12661,N_5149,N_8336);
or U12662 (N_12662,N_7509,N_4332);
nor U12663 (N_12663,N_2990,N_9659);
nor U12664 (N_12664,N_7456,N_2387);
nand U12665 (N_12665,N_8793,N_5717);
or U12666 (N_12666,N_8556,N_8145);
and U12667 (N_12667,N_6303,N_2135);
xor U12668 (N_12668,N_419,N_3869);
xor U12669 (N_12669,N_2290,N_466);
and U12670 (N_12670,N_5602,N_935);
xnor U12671 (N_12671,N_209,N_4437);
nand U12672 (N_12672,N_9486,N_1948);
and U12673 (N_12673,N_7667,N_6253);
nor U12674 (N_12674,N_9670,N_5867);
nand U12675 (N_12675,N_2552,N_8989);
nand U12676 (N_12676,N_402,N_8876);
and U12677 (N_12677,N_2873,N_4174);
nand U12678 (N_12678,N_2171,N_3617);
nand U12679 (N_12679,N_434,N_2756);
or U12680 (N_12680,N_5152,N_2971);
nor U12681 (N_12681,N_488,N_7669);
and U12682 (N_12682,N_5367,N_1274);
or U12683 (N_12683,N_852,N_4744);
xor U12684 (N_12684,N_1862,N_6539);
nor U12685 (N_12685,N_8752,N_4369);
and U12686 (N_12686,N_9807,N_3889);
and U12687 (N_12687,N_4997,N_6460);
and U12688 (N_12688,N_9323,N_7923);
or U12689 (N_12689,N_8594,N_321);
and U12690 (N_12690,N_238,N_1480);
xnor U12691 (N_12691,N_2903,N_5147);
nor U12692 (N_12692,N_4489,N_5004);
nand U12693 (N_12693,N_6655,N_8777);
and U12694 (N_12694,N_2426,N_6273);
and U12695 (N_12695,N_8392,N_5941);
nor U12696 (N_12696,N_7801,N_9133);
and U12697 (N_12697,N_6820,N_8468);
and U12698 (N_12698,N_1081,N_5446);
nor U12699 (N_12699,N_95,N_9858);
xnor U12700 (N_12700,N_9646,N_3856);
nor U12701 (N_12701,N_4040,N_8310);
nor U12702 (N_12702,N_9287,N_8199);
nand U12703 (N_12703,N_2408,N_9456);
or U12704 (N_12704,N_5768,N_2199);
and U12705 (N_12705,N_4928,N_2312);
nor U12706 (N_12706,N_9542,N_2243);
or U12707 (N_12707,N_7129,N_7062);
or U12708 (N_12708,N_5888,N_3614);
xnor U12709 (N_12709,N_3766,N_8331);
nor U12710 (N_12710,N_2311,N_5037);
xor U12711 (N_12711,N_6260,N_5580);
nand U12712 (N_12712,N_4650,N_2286);
and U12713 (N_12713,N_6454,N_2165);
or U12714 (N_12714,N_3051,N_3859);
and U12715 (N_12715,N_3528,N_8633);
xnor U12716 (N_12716,N_8831,N_4558);
or U12717 (N_12717,N_7853,N_5574);
and U12718 (N_12718,N_4952,N_2710);
or U12719 (N_12719,N_5319,N_5568);
xor U12720 (N_12720,N_4979,N_2995);
and U12721 (N_12721,N_198,N_9179);
or U12722 (N_12722,N_2182,N_4415);
nor U12723 (N_12723,N_9614,N_5246);
nand U12724 (N_12724,N_3623,N_7372);
or U12725 (N_12725,N_231,N_8655);
nor U12726 (N_12726,N_6174,N_5133);
nor U12727 (N_12727,N_2860,N_3717);
nand U12728 (N_12728,N_1106,N_8887);
or U12729 (N_12729,N_3685,N_4171);
nand U12730 (N_12730,N_7904,N_179);
nand U12731 (N_12731,N_7373,N_583);
and U12732 (N_12732,N_7422,N_1269);
nand U12733 (N_12733,N_5007,N_8243);
nand U12734 (N_12734,N_3188,N_8233);
xnor U12735 (N_12735,N_4117,N_3465);
nor U12736 (N_12736,N_7237,N_9734);
xor U12737 (N_12737,N_9599,N_7909);
or U12738 (N_12738,N_7914,N_2520);
or U12739 (N_12739,N_5025,N_6934);
nor U12740 (N_12740,N_8353,N_3601);
or U12741 (N_12741,N_1390,N_2371);
nor U12742 (N_12742,N_94,N_2148);
xor U12743 (N_12743,N_954,N_6336);
nor U12744 (N_12744,N_2105,N_6579);
nor U12745 (N_12745,N_1206,N_8764);
and U12746 (N_12746,N_905,N_1261);
xor U12747 (N_12747,N_8211,N_245);
nand U12748 (N_12748,N_3726,N_52);
and U12749 (N_12749,N_6391,N_5628);
nand U12750 (N_12750,N_4955,N_1611);
xor U12751 (N_12751,N_5488,N_6052);
nor U12752 (N_12752,N_9789,N_3425);
nand U12753 (N_12753,N_6972,N_5746);
xor U12754 (N_12754,N_9833,N_7480);
and U12755 (N_12755,N_6910,N_2502);
and U12756 (N_12756,N_3301,N_1721);
xor U12757 (N_12757,N_9312,N_9697);
xor U12758 (N_12758,N_1538,N_1465);
nor U12759 (N_12759,N_6163,N_1280);
xnor U12760 (N_12760,N_5667,N_6008);
nand U12761 (N_12761,N_8111,N_8982);
xnor U12762 (N_12762,N_4475,N_3047);
and U12763 (N_12763,N_5751,N_3729);
nand U12764 (N_12764,N_5411,N_843);
or U12765 (N_12765,N_1565,N_2463);
xnor U12766 (N_12766,N_9417,N_6307);
nand U12767 (N_12767,N_9888,N_1654);
or U12768 (N_12768,N_7262,N_7139);
xnor U12769 (N_12769,N_4717,N_5128);
and U12770 (N_12770,N_7772,N_679);
or U12771 (N_12771,N_2018,N_2127);
xor U12772 (N_12772,N_2606,N_2848);
nand U12773 (N_12773,N_2597,N_7860);
nor U12774 (N_12774,N_9610,N_8149);
nor U12775 (N_12775,N_3828,N_4310);
nor U12776 (N_12776,N_6169,N_9071);
nor U12777 (N_12777,N_7747,N_4932);
xnor U12778 (N_12778,N_856,N_3412);
xor U12779 (N_12779,N_9410,N_5741);
and U12780 (N_12780,N_8179,N_341);
xor U12781 (N_12781,N_9970,N_5197);
xnor U12782 (N_12782,N_1725,N_9529);
nor U12783 (N_12783,N_8809,N_7769);
nand U12784 (N_12784,N_6883,N_4426);
or U12785 (N_12785,N_2275,N_9925);
nor U12786 (N_12786,N_1426,N_7102);
or U12787 (N_12787,N_962,N_4235);
nor U12788 (N_12788,N_4889,N_3157);
xnor U12789 (N_12789,N_9938,N_288);
xnor U12790 (N_12790,N_8402,N_705);
nor U12791 (N_12791,N_7296,N_4616);
and U12792 (N_12792,N_7811,N_9269);
xor U12793 (N_12793,N_6711,N_663);
nor U12794 (N_12794,N_7346,N_78);
or U12795 (N_12795,N_4064,N_2514);
nand U12796 (N_12796,N_7060,N_1677);
and U12797 (N_12797,N_6560,N_6339);
xor U12798 (N_12798,N_7409,N_1771);
and U12799 (N_12799,N_1023,N_5478);
xnor U12800 (N_12800,N_5988,N_1208);
and U12801 (N_12801,N_1898,N_5812);
and U12802 (N_12802,N_6086,N_9119);
nor U12803 (N_12803,N_4898,N_6012);
and U12804 (N_12804,N_39,N_3865);
or U12805 (N_12805,N_1375,N_7933);
xor U12806 (N_12806,N_8083,N_4199);
and U12807 (N_12807,N_8050,N_3598);
nand U12808 (N_12808,N_6242,N_9110);
nand U12809 (N_12809,N_3883,N_3840);
nor U12810 (N_12810,N_3403,N_1171);
nor U12811 (N_12811,N_3177,N_5483);
nor U12812 (N_12812,N_7263,N_7311);
xnor U12813 (N_12813,N_3641,N_4096);
and U12814 (N_12814,N_8020,N_3198);
nand U12815 (N_12815,N_406,N_6494);
or U12816 (N_12816,N_3668,N_1087);
and U12817 (N_12817,N_2108,N_5619);
and U12818 (N_12818,N_7500,N_9601);
or U12819 (N_12819,N_6941,N_1348);
nor U12820 (N_12820,N_4315,N_7270);
nor U12821 (N_12821,N_4761,N_6435);
and U12822 (N_12822,N_844,N_3013);
xnor U12823 (N_12823,N_5316,N_4048);
nand U12824 (N_12824,N_4454,N_1154);
or U12825 (N_12825,N_7759,N_1649);
nor U12826 (N_12826,N_2175,N_8761);
nor U12827 (N_12827,N_2285,N_3589);
nor U12828 (N_12828,N_5851,N_5443);
or U12829 (N_12829,N_5882,N_3604);
nand U12830 (N_12830,N_6218,N_3415);
nor U12831 (N_12831,N_2949,N_5853);
xor U12832 (N_12832,N_4548,N_4759);
and U12833 (N_12833,N_2752,N_9035);
nor U12834 (N_12834,N_5677,N_7007);
and U12835 (N_12835,N_1886,N_2781);
and U12836 (N_12836,N_5548,N_2155);
nand U12837 (N_12837,N_6155,N_1163);
xor U12838 (N_12838,N_3318,N_1374);
xnor U12839 (N_12839,N_1854,N_9731);
xnor U12840 (N_12840,N_6774,N_5961);
or U12841 (N_12841,N_3973,N_192);
xor U12842 (N_12842,N_2537,N_9032);
xor U12843 (N_12843,N_8711,N_6093);
and U12844 (N_12844,N_9019,N_204);
or U12845 (N_12845,N_775,N_6794);
and U12846 (N_12846,N_5600,N_8629);
xor U12847 (N_12847,N_4388,N_2293);
and U12848 (N_12848,N_3368,N_2809);
nand U12849 (N_12849,N_6522,N_5959);
nand U12850 (N_12850,N_7543,N_4346);
xor U12851 (N_12851,N_1177,N_6213);
and U12852 (N_12852,N_9538,N_652);
nand U12853 (N_12853,N_1987,N_3479);
xor U12854 (N_12854,N_1926,N_5932);
xnor U12855 (N_12855,N_9374,N_6856);
nor U12856 (N_12856,N_7514,N_5449);
nand U12857 (N_12857,N_343,N_9021);
or U12858 (N_12858,N_2952,N_140);
nor U12859 (N_12859,N_2055,N_1718);
nor U12860 (N_12860,N_4783,N_8270);
nor U12861 (N_12861,N_5255,N_7008);
nor U12862 (N_12862,N_3446,N_890);
or U12863 (N_12863,N_297,N_3467);
and U12864 (N_12864,N_7465,N_8515);
nor U12865 (N_12865,N_5914,N_643);
or U12866 (N_12866,N_1674,N_3812);
and U12867 (N_12867,N_1466,N_5168);
xnor U12868 (N_12868,N_6767,N_9869);
xor U12869 (N_12869,N_8885,N_4843);
nand U12870 (N_12870,N_1749,N_4151);
nor U12871 (N_12871,N_9150,N_8030);
nor U12872 (N_12872,N_6487,N_3954);
xnor U12873 (N_12873,N_6497,N_4694);
or U12874 (N_12874,N_7527,N_6363);
or U12875 (N_12875,N_7109,N_276);
nor U12876 (N_12876,N_646,N_1614);
nand U12877 (N_12877,N_2013,N_8422);
xor U12878 (N_12878,N_5163,N_6610);
nand U12879 (N_12879,N_3715,N_2184);
nand U12880 (N_12880,N_9175,N_3225);
nand U12881 (N_12881,N_4223,N_7);
xnor U12882 (N_12882,N_120,N_7188);
xnor U12883 (N_12883,N_4544,N_9840);
and U12884 (N_12884,N_6784,N_9331);
xnor U12885 (N_12885,N_6829,N_4772);
or U12886 (N_12886,N_433,N_5134);
nor U12887 (N_12887,N_1091,N_7202);
nand U12888 (N_12888,N_2647,N_1175);
and U12889 (N_12889,N_1636,N_9347);
nor U12890 (N_12890,N_4785,N_840);
nand U12891 (N_12891,N_7844,N_7693);
nand U12892 (N_12892,N_8425,N_2771);
nand U12893 (N_12893,N_9881,N_1435);
and U12894 (N_12894,N_8344,N_5353);
nor U12895 (N_12895,N_7379,N_8249);
or U12896 (N_12896,N_2477,N_5801);
nor U12897 (N_12897,N_394,N_1297);
xnor U12898 (N_12898,N_1955,N_3289);
and U12899 (N_12899,N_5141,N_4582);
nand U12900 (N_12900,N_5865,N_5341);
and U12901 (N_12901,N_511,N_1869);
and U12902 (N_12902,N_6578,N_692);
and U12903 (N_12903,N_5917,N_6039);
nor U12904 (N_12904,N_3936,N_1080);
xor U12905 (N_12905,N_1980,N_1066);
or U12906 (N_12906,N_6266,N_1730);
and U12907 (N_12907,N_7322,N_8702);
and U12908 (N_12908,N_3142,N_7631);
xnor U12909 (N_12909,N_7886,N_9818);
nand U12910 (N_12910,N_6153,N_9459);
and U12911 (N_12911,N_8033,N_2893);
xnor U12912 (N_12912,N_3994,N_2411);
nor U12913 (N_12913,N_9310,N_8262);
xnor U12914 (N_12914,N_9584,N_8949);
nand U12915 (N_12915,N_7495,N_8968);
xor U12916 (N_12916,N_1876,N_1952);
nor U12917 (N_12917,N_2235,N_5910);
nor U12918 (N_12918,N_6728,N_6107);
and U12919 (N_12919,N_8550,N_7560);
nor U12920 (N_12920,N_6675,N_1263);
nor U12921 (N_12921,N_3962,N_4876);
nand U12922 (N_12922,N_9180,N_9710);
nor U12923 (N_12923,N_1044,N_6209);
and U12924 (N_12924,N_7630,N_2718);
nand U12925 (N_12925,N_5401,N_2316);
nand U12926 (N_12926,N_2592,N_5849);
and U12927 (N_12927,N_4461,N_1441);
nor U12928 (N_12928,N_236,N_5870);
nand U12929 (N_12929,N_7055,N_1092);
xor U12930 (N_12930,N_4071,N_3727);
xnor U12931 (N_12931,N_3175,N_1021);
or U12932 (N_12932,N_1531,N_8289);
nor U12933 (N_12933,N_4359,N_5153);
or U12934 (N_12934,N_2434,N_8580);
nor U12935 (N_12935,N_9551,N_4425);
nand U12936 (N_12936,N_5436,N_3587);
or U12937 (N_12937,N_6781,N_9691);
or U12938 (N_12938,N_283,N_8492);
or U12939 (N_12939,N_7797,N_7793);
nand U12940 (N_12940,N_2473,N_3260);
nand U12941 (N_12941,N_9068,N_4579);
xor U12942 (N_12942,N_7420,N_1951);
nand U12943 (N_12943,N_3300,N_253);
nand U12944 (N_12944,N_4773,N_3938);
and U12945 (N_12945,N_2498,N_4842);
nor U12946 (N_12946,N_3103,N_2451);
xor U12947 (N_12947,N_1575,N_6395);
and U12948 (N_12948,N_4012,N_8644);
xnor U12949 (N_12949,N_1954,N_5521);
and U12950 (N_12950,N_5301,N_6656);
xnor U12951 (N_12951,N_3254,N_178);
nand U12952 (N_12952,N_7549,N_6472);
xnor U12953 (N_12953,N_3109,N_4229);
and U12954 (N_12954,N_5608,N_1130);
nand U12955 (N_12955,N_7916,N_6096);
xor U12956 (N_12956,N_9651,N_1742);
or U12957 (N_12957,N_6477,N_6428);
nand U12958 (N_12958,N_5604,N_5268);
and U12959 (N_12959,N_1027,N_9106);
xor U12960 (N_12960,N_84,N_4519);
nor U12961 (N_12961,N_6905,N_2189);
or U12962 (N_12962,N_8164,N_9723);
and U12963 (N_12963,N_7927,N_7530);
nand U12964 (N_12964,N_5614,N_5144);
xnor U12965 (N_12965,N_7847,N_6982);
nand U12966 (N_12966,N_6351,N_5616);
and U12967 (N_12967,N_5116,N_3573);
xor U12968 (N_12968,N_9407,N_4746);
or U12969 (N_12969,N_7080,N_7215);
or U12970 (N_12970,N_9371,N_3218);
or U12971 (N_12971,N_6971,N_5039);
and U12972 (N_12972,N_5866,N_4623);
xor U12973 (N_12973,N_7690,N_4224);
xor U12974 (N_12974,N_8819,N_866);
or U12975 (N_12975,N_9834,N_4280);
xor U12976 (N_12976,N_8813,N_3674);
and U12977 (N_12977,N_8775,N_4551);
nor U12978 (N_12978,N_7443,N_2738);
nor U12979 (N_12979,N_5451,N_4354);
xnor U12980 (N_12980,N_284,N_1911);
and U12981 (N_12981,N_2072,N_5641);
xor U12982 (N_12982,N_1406,N_5777);
or U12983 (N_12983,N_362,N_1008);
and U12984 (N_12984,N_4950,N_8942);
or U12985 (N_12985,N_8648,N_22);
or U12986 (N_12986,N_7662,N_165);
nor U12987 (N_12987,N_8913,N_5493);
and U12988 (N_12988,N_9721,N_3417);
nand U12989 (N_12989,N_9249,N_4374);
nor U12990 (N_12990,N_6050,N_4053);
xor U12991 (N_12991,N_807,N_9634);
nor U12992 (N_12992,N_2745,N_50);
xnor U12993 (N_12993,N_9143,N_3011);
nand U12994 (N_12994,N_4634,N_814);
and U12995 (N_12995,N_9369,N_5207);
nand U12996 (N_12996,N_2586,N_6404);
nand U12997 (N_12997,N_9248,N_3600);
nand U12998 (N_12998,N_5903,N_7507);
nand U12999 (N_12999,N_142,N_1735);
xor U13000 (N_13000,N_2693,N_6745);
xor U13001 (N_13001,N_8691,N_599);
nor U13002 (N_13002,N_797,N_9389);
xnor U13003 (N_13003,N_5462,N_4834);
nand U13004 (N_13004,N_3721,N_6157);
nor U13005 (N_13005,N_8388,N_7395);
or U13006 (N_13006,N_2000,N_8044);
xor U13007 (N_13007,N_5592,N_4866);
and U13008 (N_13008,N_514,N_3855);
nand U13009 (N_13009,N_2110,N_9996);
xnor U13010 (N_13010,N_3819,N_294);
or U13011 (N_13011,N_4855,N_711);
nand U13012 (N_13012,N_1005,N_4298);
nand U13013 (N_13013,N_8158,N_9191);
xor U13014 (N_13014,N_2644,N_8389);
or U13015 (N_13015,N_9965,N_8739);
and U13016 (N_13016,N_322,N_6598);
or U13017 (N_13017,N_1360,N_4517);
xor U13018 (N_13018,N_1187,N_2892);
xnor U13019 (N_13019,N_1757,N_9112);
nor U13020 (N_13020,N_2866,N_9250);
nand U13021 (N_13021,N_2579,N_7399);
nand U13022 (N_13022,N_7533,N_5704);
nand U13023 (N_13023,N_2538,N_6275);
nand U13024 (N_13024,N_7049,N_5517);
nor U13025 (N_13025,N_7058,N_6217);
nor U13026 (N_13026,N_9552,N_4101);
or U13027 (N_13027,N_7538,N_4365);
xor U13028 (N_13028,N_49,N_3942);
or U13029 (N_13029,N_2842,N_5242);
xor U13030 (N_13030,N_9039,N_291);
xor U13031 (N_13031,N_1136,N_4505);
or U13032 (N_13032,N_28,N_767);
nand U13033 (N_13033,N_6448,N_8688);
and U13034 (N_13034,N_2363,N_2376);
and U13035 (N_13035,N_3904,N_5722);
nand U13036 (N_13036,N_1704,N_728);
or U13037 (N_13037,N_9263,N_867);
nor U13038 (N_13038,N_1838,N_3473);
nor U13039 (N_13039,N_5447,N_7925);
and U13040 (N_13040,N_7783,N_2037);
nand U13041 (N_13041,N_7115,N_1478);
and U13042 (N_13042,N_3205,N_8063);
or U13043 (N_13043,N_768,N_2631);
or U13044 (N_13044,N_3080,N_2152);
nand U13045 (N_13045,N_4350,N_7595);
and U13046 (N_13046,N_2543,N_7038);
and U13047 (N_13047,N_3537,N_2043);
xnor U13048 (N_13048,N_1237,N_4153);
nand U13049 (N_13049,N_3681,N_1183);
nor U13050 (N_13050,N_2328,N_7292);
nor U13051 (N_13051,N_3578,N_4934);
and U13052 (N_13052,N_2507,N_5318);
and U13053 (N_13053,N_4540,N_3740);
and U13054 (N_13054,N_3066,N_2208);
xor U13055 (N_13055,N_8608,N_5082);
or U13056 (N_13056,N_548,N_9015);
nand U13057 (N_13057,N_4276,N_2891);
or U13058 (N_13058,N_4891,N_676);
xnor U13059 (N_13059,N_246,N_8081);
nand U13060 (N_13060,N_7004,N_1840);
xor U13061 (N_13061,N_5063,N_3919);
nand U13062 (N_13062,N_3829,N_5406);
or U13063 (N_13063,N_5969,N_3068);
and U13064 (N_13064,N_6366,N_6026);
xnor U13065 (N_13065,N_9981,N_2728);
and U13066 (N_13066,N_6716,N_8061);
or U13067 (N_13067,N_9139,N_7632);
and U13068 (N_13068,N_2944,N_7935);
nand U13069 (N_13069,N_9689,N_2457);
nor U13070 (N_13070,N_5212,N_3034);
nor U13071 (N_13071,N_7186,N_9910);
or U13072 (N_13072,N_9502,N_6822);
or U13073 (N_13073,N_4850,N_1529);
or U13074 (N_13074,N_1618,N_7921);
xor U13075 (N_13075,N_901,N_2921);
nor U13076 (N_13076,N_5893,N_8592);
nand U13077 (N_13077,N_8962,N_8072);
or U13078 (N_13078,N_5709,N_7945);
and U13079 (N_13079,N_453,N_412);
and U13080 (N_13080,N_4545,N_2667);
nor U13081 (N_13081,N_3602,N_6880);
nand U13082 (N_13082,N_8132,N_9811);
nor U13083 (N_13083,N_5685,N_62);
nand U13084 (N_13084,N_438,N_102);
xnor U13085 (N_13085,N_677,N_1358);
xnor U13086 (N_13086,N_1956,N_5652);
nand U13087 (N_13087,N_8740,N_88);
nor U13088 (N_13088,N_2296,N_4001);
xor U13089 (N_13089,N_2225,N_8152);
nor U13090 (N_13090,N_6778,N_7028);
or U13091 (N_13091,N_9622,N_7290);
nor U13092 (N_13092,N_337,N_5930);
xnor U13093 (N_13093,N_8260,N_1460);
xnor U13094 (N_13094,N_5266,N_9566);
nand U13095 (N_13095,N_6693,N_3277);
or U13096 (N_13096,N_6796,N_3611);
nor U13097 (N_13097,N_2717,N_2687);
xor U13098 (N_13098,N_6466,N_4722);
nand U13099 (N_13099,N_153,N_3270);
or U13100 (N_13100,N_4629,N_9683);
or U13101 (N_13101,N_8663,N_1427);
or U13102 (N_13102,N_8470,N_9994);
or U13103 (N_13103,N_4844,N_6694);
and U13104 (N_13104,N_3171,N_5472);
and U13105 (N_13105,N_7011,N_4709);
nand U13106 (N_13106,N_2522,N_6531);
or U13107 (N_13107,N_9289,N_7643);
or U13108 (N_13108,N_656,N_7474);
and U13109 (N_13109,N_9865,N_3071);
or U13110 (N_13110,N_3285,N_3802);
or U13111 (N_13111,N_361,N_8788);
nand U13112 (N_13112,N_1319,N_9340);
or U13113 (N_13113,N_5432,N_9418);
or U13114 (N_13114,N_6089,N_5407);
nor U13115 (N_13115,N_389,N_5252);
and U13116 (N_13116,N_9227,N_937);
xnor U13117 (N_13117,N_2533,N_8991);
or U13118 (N_13118,N_4977,N_504);
or U13119 (N_13119,N_1933,N_5738);
or U13120 (N_13120,N_9976,N_1516);
xor U13121 (N_13121,N_4804,N_1510);
and U13122 (N_13122,N_3670,N_4172);
nand U13123 (N_13123,N_8641,N_4084);
and U13124 (N_13124,N_6225,N_3129);
or U13125 (N_13125,N_9864,N_7882);
or U13126 (N_13126,N_5934,N_8066);
nand U13127 (N_13127,N_9461,N_2340);
or U13128 (N_13128,N_4061,N_2233);
and U13129 (N_13129,N_5830,N_4674);
or U13130 (N_13130,N_2479,N_2289);
and U13131 (N_13131,N_5056,N_8512);
nand U13132 (N_13132,N_8087,N_2817);
or U13133 (N_13133,N_6084,N_2689);
and U13134 (N_13134,N_9500,N_9746);
nand U13135 (N_13135,N_8741,N_7264);
or U13136 (N_13136,N_3720,N_1257);
and U13137 (N_13137,N_1291,N_5475);
nor U13138 (N_13138,N_6850,N_5088);
and U13139 (N_13139,N_1726,N_3067);
or U13140 (N_13140,N_8985,N_7863);
xnor U13141 (N_13141,N_3795,N_35);
xor U13142 (N_13142,N_1932,N_8993);
and U13143 (N_13143,N_7120,N_3701);
or U13144 (N_13144,N_7771,N_9561);
nor U13145 (N_13145,N_6110,N_4556);
nor U13146 (N_13146,N_9056,N_5137);
nor U13147 (N_13147,N_4668,N_3408);
nand U13148 (N_13148,N_6222,N_8839);
and U13149 (N_13149,N_5422,N_6681);
nand U13150 (N_13150,N_7704,N_7161);
and U13151 (N_13151,N_6742,N_7303);
xnor U13152 (N_13152,N_5609,N_6224);
nor U13153 (N_13153,N_2114,N_4201);
or U13154 (N_13154,N_4480,N_6813);
nand U13155 (N_13155,N_2231,N_904);
and U13156 (N_13156,N_8760,N_2144);
nor U13157 (N_13157,N_5029,N_2897);
nand U13158 (N_13158,N_1256,N_5506);
or U13159 (N_13159,N_8407,N_1115);
xor U13160 (N_13160,N_8160,N_536);
nor U13161 (N_13161,N_7537,N_4745);
or U13162 (N_13162,N_1410,N_7556);
and U13163 (N_13163,N_6068,N_6589);
or U13164 (N_13164,N_1162,N_9574);
nand U13165 (N_13165,N_5459,N_1953);
nor U13166 (N_13166,N_6673,N_1902);
or U13167 (N_13167,N_1630,N_4586);
xnor U13168 (N_13168,N_7874,N_108);
nand U13169 (N_13169,N_8840,N_5552);
or U13170 (N_13170,N_6097,N_2739);
xor U13171 (N_13171,N_7193,N_7181);
or U13172 (N_13172,N_7291,N_9642);
or U13173 (N_13173,N_1004,N_1675);
nand U13174 (N_13174,N_5606,N_1694);
nand U13175 (N_13175,N_2278,N_7295);
and U13176 (N_13176,N_9762,N_6019);
or U13177 (N_13177,N_4689,N_4872);
nand U13178 (N_13178,N_9638,N_3780);
xnor U13179 (N_13179,N_1069,N_7017);
and U13180 (N_13180,N_6750,N_5646);
nor U13181 (N_13181,N_2679,N_2749);
nor U13182 (N_13182,N_9616,N_8156);
xor U13183 (N_13183,N_3448,N_3081);
xnor U13184 (N_13184,N_7505,N_671);
or U13185 (N_13185,N_9221,N_5972);
nor U13186 (N_13186,N_5000,N_6032);
and U13187 (N_13187,N_1279,N_61);
or U13188 (N_13188,N_3945,N_8734);
nor U13189 (N_13189,N_784,N_331);
nor U13190 (N_13190,N_4086,N_641);
or U13191 (N_13191,N_4264,N_4389);
xnor U13192 (N_13192,N_1339,N_7978);
and U13193 (N_13193,N_5317,N_2928);
nor U13194 (N_13194,N_5663,N_418);
nand U13195 (N_13195,N_7335,N_355);
and U13196 (N_13196,N_1619,N_6327);
nand U13197 (N_13197,N_7314,N_1739);
and U13198 (N_13198,N_2139,N_2482);
or U13199 (N_13199,N_7397,N_5299);
xnor U13200 (N_13200,N_6046,N_2907);
or U13201 (N_13201,N_4976,N_1964);
nand U13202 (N_13202,N_5898,N_5169);
and U13203 (N_13203,N_9076,N_7954);
nand U13204 (N_13204,N_2750,N_1077);
and U13205 (N_13205,N_7698,N_736);
xor U13206 (N_13206,N_8092,N_6527);
xnor U13207 (N_13207,N_9543,N_293);
xor U13208 (N_13208,N_1962,N_7883);
or U13209 (N_13209,N_2116,N_2425);
nor U13210 (N_13210,N_6682,N_2207);
xnor U13211 (N_13211,N_7392,N_2250);
xor U13212 (N_13212,N_9880,N_6892);
xnor U13213 (N_13213,N_2948,N_1377);
nor U13214 (N_13214,N_2314,N_2467);
xnor U13215 (N_13215,N_38,N_2614);
or U13216 (N_13216,N_2793,N_132);
xnor U13217 (N_13217,N_7822,N_5829);
and U13218 (N_13218,N_3860,N_4416);
nand U13219 (N_13219,N_8883,N_436);
xnor U13220 (N_13220,N_2588,N_4905);
xnor U13221 (N_13221,N_4198,N_5673);
or U13222 (N_13222,N_9612,N_3332);
and U13223 (N_13223,N_1664,N_8384);
and U13224 (N_13224,N_1273,N_4034);
nor U13225 (N_13225,N_5371,N_6);
xor U13226 (N_13226,N_8139,N_6926);
nand U13227 (N_13227,N_7503,N_9936);
nor U13228 (N_13228,N_1690,N_6944);
or U13229 (N_13229,N_5700,N_7799);
xnor U13230 (N_13230,N_2042,N_8093);
or U13231 (N_13231,N_219,N_6077);
nor U13232 (N_13232,N_1200,N_7265);
xor U13233 (N_13233,N_2911,N_2937);
nor U13234 (N_13234,N_7479,N_7839);
or U13235 (N_13235,N_4228,N_2769);
or U13236 (N_13236,N_3848,N_4635);
and U13237 (N_13237,N_2872,N_6754);
xor U13238 (N_13238,N_8863,N_3873);
nor U13239 (N_13239,N_9301,N_4580);
nand U13240 (N_13240,N_2369,N_7472);
nor U13241 (N_13241,N_5666,N_2795);
xnor U13242 (N_13242,N_8744,N_8601);
xnor U13243 (N_13243,N_3874,N_4003);
nand U13244 (N_13244,N_8927,N_8236);
or U13245 (N_13245,N_5231,N_9445);
or U13246 (N_13246,N_8172,N_786);
xnor U13247 (N_13247,N_8806,N_3699);
and U13248 (N_13248,N_8339,N_7445);
and U13249 (N_13249,N_3065,N_6600);
or U13250 (N_13250,N_2033,N_4824);
xor U13251 (N_13251,N_4510,N_4482);
and U13252 (N_13252,N_2723,N_3436);
nor U13253 (N_13253,N_3896,N_5234);
nor U13254 (N_13254,N_4059,N_8753);
nor U13255 (N_13255,N_2894,N_7166);
xnor U13256 (N_13256,N_8347,N_1908);
nor U13257 (N_13257,N_6961,N_2356);
nand U13258 (N_13258,N_6570,N_742);
and U13259 (N_13259,N_4923,N_9915);
nand U13260 (N_13260,N_3258,N_9465);
nand U13261 (N_13261,N_1621,N_299);
and U13262 (N_13262,N_773,N_3119);
nor U13263 (N_13263,N_5191,N_6188);
xnor U13264 (N_13264,N_3424,N_1553);
nor U13265 (N_13265,N_5537,N_9361);
nand U13266 (N_13266,N_2626,N_2557);
and U13267 (N_13267,N_1896,N_7070);
or U13268 (N_13268,N_5203,N_7917);
nand U13269 (N_13269,N_4175,N_9608);
nand U13270 (N_13270,N_2119,N_8040);
and U13271 (N_13271,N_2916,N_7834);
and U13272 (N_13272,N_8514,N_2004);
xnor U13273 (N_13273,N_2071,N_3120);
and U13274 (N_13274,N_3025,N_4720);
nor U13275 (N_13275,N_2005,N_7741);
nand U13276 (N_13276,N_7651,N_9715);
xnor U13277 (N_13277,N_8614,N_2133);
nor U13278 (N_13278,N_9087,N_8692);
nand U13279 (N_13279,N_933,N_9907);
and U13280 (N_13280,N_5960,N_2904);
xnor U13281 (N_13281,N_8454,N_3626);
xor U13282 (N_13282,N_1521,N_3193);
or U13283 (N_13283,N_4390,N_3345);
nor U13284 (N_13284,N_4211,N_6703);
nor U13285 (N_13285,N_9421,N_3091);
and U13286 (N_13286,N_4572,N_1289);
or U13287 (N_13287,N_1825,N_2244);
nor U13288 (N_13288,N_9487,N_4381);
or U13289 (N_13289,N_2801,N_4707);
xnor U13290 (N_13290,N_6212,N_9230);
xnor U13291 (N_13291,N_1560,N_8037);
nor U13292 (N_13292,N_7902,N_5042);
and U13293 (N_13293,N_6895,N_475);
or U13294 (N_13294,N_2168,N_4819);
or U13295 (N_13295,N_4319,N_4067);
and U13296 (N_13296,N_8390,N_9252);
xor U13297 (N_13297,N_5725,N_1405);
nor U13298 (N_13298,N_7855,N_4138);
and U13299 (N_13299,N_1957,N_8516);
or U13300 (N_13300,N_1552,N_625);
nand U13301 (N_13301,N_650,N_9800);
and U13302 (N_13302,N_8822,N_5415);
and U13303 (N_13303,N_6342,N_8293);
or U13304 (N_13304,N_880,N_6109);
and U13305 (N_13305,N_1883,N_5603);
or U13306 (N_13306,N_5347,N_1526);
xnor U13307 (N_13307,N_7227,N_2427);
nand U13308 (N_13308,N_6004,N_1207);
nand U13309 (N_13309,N_907,N_6387);
xor U13310 (N_13310,N_56,N_6136);
nor U13311 (N_13311,N_576,N_3485);
nand U13312 (N_13312,N_8367,N_3982);
nor U13313 (N_13313,N_9172,N_9932);
nand U13314 (N_13314,N_2407,N_5965);
and U13315 (N_13315,N_1050,N_8306);
nand U13316 (N_13316,N_3510,N_9195);
or U13317 (N_13317,N_929,N_5466);
nor U13318 (N_13318,N_3057,N_9532);
or U13319 (N_13319,N_4329,N_3349);
and U13320 (N_13320,N_9375,N_8317);
nand U13321 (N_13321,N_1071,N_2812);
or U13322 (N_13322,N_6002,N_6358);
nand U13323 (N_13323,N_3772,N_8438);
or U13324 (N_13324,N_6292,N_6647);
xnor U13325 (N_13325,N_4043,N_4357);
xnor U13326 (N_13326,N_7431,N_936);
nand U13327 (N_13327,N_8642,N_3308);
and U13328 (N_13328,N_8376,N_573);
and U13329 (N_13329,N_8077,N_2045);
nand U13330 (N_13330,N_8307,N_2381);
xor U13331 (N_13331,N_3767,N_3520);
xnor U13332 (N_13332,N_877,N_3661);
and U13333 (N_13333,N_9362,N_7564);
nand U13334 (N_13334,N_4256,N_1259);
nor U13335 (N_13335,N_3631,N_6398);
nand U13336 (N_13336,N_171,N_2029);
or U13337 (N_13337,N_8579,N_8002);
xnor U13338 (N_13338,N_721,N_6968);
and U13339 (N_13339,N_4143,N_7552);
nand U13340 (N_13340,N_106,N_5805);
or U13341 (N_13341,N_5547,N_5810);
or U13342 (N_13342,N_2081,N_6571);
nor U13343 (N_13343,N_1366,N_3570);
and U13344 (N_13344,N_5784,N_5601);
nor U13345 (N_13345,N_2082,N_4253);
or U13346 (N_13346,N_4861,N_2017);
xor U13347 (N_13347,N_2344,N_6899);
or U13348 (N_13348,N_7369,N_9490);
or U13349 (N_13349,N_9135,N_1294);
nand U13350 (N_13350,N_3569,N_1467);
nor U13351 (N_13351,N_2315,N_3029);
nand U13352 (N_13352,N_5891,N_4647);
or U13353 (N_13353,N_2343,N_3134);
nor U13354 (N_13354,N_5698,N_6626);
nand U13355 (N_13355,N_3590,N_1888);
or U13356 (N_13356,N_7288,N_7151);
nor U13357 (N_13357,N_8634,N_6269);
nor U13358 (N_13358,N_3566,N_4023);
nand U13359 (N_13359,N_2611,N_1605);
and U13360 (N_13360,N_262,N_2829);
and U13361 (N_13361,N_6815,N_3491);
nor U13362 (N_13362,N_1271,N_9168);
or U13363 (N_13363,N_4848,N_7200);
nand U13364 (N_13364,N_2337,N_9328);
or U13365 (N_13365,N_1178,N_3881);
nand U13366 (N_13366,N_3155,N_3529);
nand U13367 (N_13367,N_4626,N_2277);
xnor U13368 (N_13368,N_437,N_7672);
and U13369 (N_13369,N_5161,N_6936);
nand U13370 (N_13370,N_191,N_6617);
nand U13371 (N_13371,N_1752,N_7044);
xnor U13372 (N_13372,N_9892,N_1160);
or U13373 (N_13373,N_1490,N_6828);
and U13374 (N_13374,N_2646,N_9576);
xor U13375 (N_13375,N_458,N_6475);
xor U13376 (N_13376,N_4259,N_1450);
nor U13377 (N_13377,N_5841,N_9237);
or U13378 (N_13378,N_7169,N_2951);
and U13379 (N_13379,N_4328,N_3971);
xor U13380 (N_13380,N_2827,N_3814);
and U13381 (N_13381,N_535,N_9079);
and U13382 (N_13382,N_3916,N_8379);
and U13383 (N_13383,N_8343,N_9381);
or U13384 (N_13384,N_7661,N_5804);
nand U13385 (N_13385,N_4102,N_664);
or U13386 (N_13386,N_9781,N_8337);
xor U13387 (N_13387,N_1762,N_2115);
nand U13388 (N_13388,N_9519,N_8527);
nand U13389 (N_13389,N_8590,N_390);
nor U13390 (N_13390,N_9458,N_8960);
nand U13391 (N_13391,N_3393,N_5815);
nand U13392 (N_13392,N_7324,N_2181);
and U13393 (N_13393,N_2699,N_4113);
nand U13394 (N_13394,N_657,N_1241);
xnor U13395 (N_13395,N_7918,N_8981);
xor U13396 (N_13396,N_1402,N_3774);
and U13397 (N_13397,N_364,N_9956);
and U13398 (N_13398,N_4662,N_1551);
or U13399 (N_13399,N_3330,N_1142);
and U13400 (N_13400,N_2080,N_7401);
nor U13401 (N_13401,N_9867,N_5733);
nand U13402 (N_13402,N_482,N_6458);
nand U13403 (N_13403,N_5030,N_9373);
nor U13404 (N_13404,N_5748,N_8995);
nor U13405 (N_13405,N_5003,N_5403);
xor U13406 (N_13406,N_8886,N_9796);
and U13407 (N_13407,N_6923,N_7928);
and U13408 (N_13408,N_47,N_2513);
nand U13409 (N_13409,N_7268,N_516);
nand U13410 (N_13410,N_4693,N_5392);
nand U13411 (N_13411,N_9505,N_7871);
xnor U13412 (N_13412,N_5534,N_9515);
and U13413 (N_13413,N_4323,N_5320);
nor U13414 (N_13414,N_2609,N_8899);
or U13415 (N_13415,N_7944,N_8022);
or U13416 (N_13416,N_5071,N_1260);
nand U13417 (N_13417,N_3365,N_1204);
xor U13418 (N_13418,N_2678,N_5752);
nor U13419 (N_13419,N_17,N_1591);
nor U13420 (N_13420,N_8587,N_5360);
and U13421 (N_13421,N_9549,N_1688);
and U13422 (N_13422,N_3757,N_9732);
nor U13423 (N_13423,N_7920,N_4463);
nand U13424 (N_13424,N_290,N_4791);
nand U13425 (N_13425,N_6714,N_1508);
xnor U13426 (N_13426,N_1253,N_2594);
xor U13427 (N_13427,N_212,N_2491);
and U13428 (N_13428,N_1609,N_4760);
or U13429 (N_13429,N_3806,N_6007);
nor U13430 (N_13430,N_1323,N_6640);
xor U13431 (N_13431,N_6623,N_6210);
and U13432 (N_13432,N_9495,N_8274);
nand U13433 (N_13433,N_682,N_5530);
or U13434 (N_13434,N_359,N_2270);
or U13435 (N_13435,N_7911,N_3775);
xor U13436 (N_13436,N_8569,N_9625);
xnor U13437 (N_13437,N_5931,N_5883);
xnor U13438 (N_13438,N_9390,N_9757);
nand U13439 (N_13439,N_2705,N_6863);
and U13440 (N_13440,N_9902,N_8714);
and U13441 (N_13441,N_2436,N_2330);
and U13442 (N_13442,N_3322,N_3998);
nand U13443 (N_13443,N_2703,N_7608);
and U13444 (N_13444,N_175,N_8972);
nand U13445 (N_13445,N_9002,N_1468);
nand U13446 (N_13446,N_226,N_9146);
nand U13447 (N_13447,N_1482,N_9100);
nor U13448 (N_13448,N_2670,N_5126);
and U13449 (N_13449,N_8144,N_2073);
and U13450 (N_13450,N_286,N_9524);
nor U13451 (N_13451,N_2217,N_9665);
xor U13452 (N_13452,N_3765,N_7407);
xor U13453 (N_13453,N_5311,N_101);
and U13454 (N_13454,N_4538,N_527);
xnor U13455 (N_13455,N_4492,N_7236);
and U13456 (N_13456,N_2847,N_9766);
xor U13457 (N_13457,N_3794,N_6984);
nor U13458 (N_13458,N_6054,N_7621);
or U13459 (N_13459,N_93,N_2218);
nand U13460 (N_13460,N_9254,N_8828);
xnor U13461 (N_13461,N_8750,N_74);
or U13462 (N_13462,N_1759,N_354);
nand U13463 (N_13463,N_5072,N_7074);
and U13464 (N_13464,N_7087,N_9411);
and U13465 (N_13465,N_7778,N_6043);
nor U13466 (N_13466,N_6462,N_3677);
xnor U13467 (N_13467,N_794,N_8853);
or U13468 (N_13468,N_4534,N_510);
nand U13469 (N_13469,N_5230,N_4874);
nor U13470 (N_13470,N_541,N_9282);
and U13471 (N_13471,N_5219,N_8125);
nor U13472 (N_13472,N_138,N_8939);
or U13473 (N_13473,N_5670,N_6076);
xor U13474 (N_13474,N_3170,N_3990);
nor U13475 (N_13475,N_7374,N_9014);
nand U13476 (N_13476,N_3985,N_8848);
or U13477 (N_13477,N_7546,N_1108);
nand U13478 (N_13478,N_7208,N_2305);
xnor U13479 (N_13479,N_2229,N_3980);
and U13480 (N_13480,N_7267,N_4130);
or U13481 (N_13481,N_544,N_7623);
and U13482 (N_13482,N_6807,N_8457);
or U13483 (N_13483,N_8095,N_3882);
or U13484 (N_13484,N_2163,N_4204);
nand U13485 (N_13485,N_5564,N_6634);
and U13486 (N_13486,N_5117,N_8523);
xor U13487 (N_13487,N_5567,N_8908);
xnor U13488 (N_13488,N_7616,N_9272);
nand U13489 (N_13489,N_6929,N_2092);
or U13490 (N_13490,N_9125,N_7253);
and U13491 (N_13491,N_5892,N_9192);
or U13492 (N_13492,N_9332,N_4144);
nand U13493 (N_13493,N_9308,N_8328);
or U13494 (N_13494,N_273,N_7053);
or U13495 (N_13495,N_7452,N_804);
nor U13496 (N_13496,N_4337,N_5818);
nand U13497 (N_13497,N_80,N_6612);
nand U13498 (N_13498,N_7592,N_1464);
nor U13499 (N_13499,N_3813,N_6835);
nand U13500 (N_13500,N_3327,N_9503);
or U13501 (N_13501,N_9974,N_5942);
xnor U13502 (N_13502,N_5927,N_8994);
xnor U13503 (N_13503,N_2001,N_3565);
nand U13504 (N_13504,N_7261,N_3688);
nor U13505 (N_13505,N_2489,N_97);
nand U13506 (N_13506,N_6298,N_9089);
nor U13507 (N_13507,N_4165,N_2078);
nor U13508 (N_13508,N_5745,N_9929);
or U13509 (N_13509,N_7403,N_3238);
nand U13510 (N_13510,N_7689,N_2509);
nor U13511 (N_13511,N_6261,N_40);
nand U13512 (N_13512,N_5083,N_3444);
xnor U13513 (N_13513,N_4991,N_3684);
and U13514 (N_13514,N_196,N_8104);
nand U13515 (N_13515,N_3110,N_162);
nand U13516 (N_13516,N_6202,N_6239);
and U13517 (N_13517,N_2806,N_7558);
xor U13518 (N_13518,N_9598,N_2774);
or U13519 (N_13519,N_1436,N_5956);
xnor U13520 (N_13520,N_8034,N_3297);
nor U13521 (N_13521,N_2628,N_125);
and U13522 (N_13522,N_5911,N_6540);
or U13523 (N_13523,N_4812,N_5617);
nand U13524 (N_13524,N_3229,N_9271);
xor U13525 (N_13525,N_883,N_3098);
nand U13526 (N_13526,N_2418,N_6679);
nor U13527 (N_13527,N_403,N_7180);
nand U13528 (N_13528,N_9711,N_4157);
and U13529 (N_13529,N_1286,N_9905);
nand U13530 (N_13530,N_4062,N_9738);
nand U13531 (N_13531,N_2320,N_9801);
and U13532 (N_13532,N_4079,N_1223);
nor U13533 (N_13533,N_6476,N_8414);
nand U13534 (N_13534,N_8858,N_7073);
and U13535 (N_13535,N_6975,N_5484);
and U13536 (N_13536,N_7678,N_694);
or U13537 (N_13537,N_4868,N_3908);
and U13538 (N_13538,N_4237,N_1786);
or U13539 (N_13539,N_3719,N_2779);
or U13540 (N_13540,N_9995,N_4495);
and U13541 (N_13541,N_4380,N_648);
or U13542 (N_13542,N_9167,N_9196);
xnor U13543 (N_13543,N_5399,N_6194);
or U13544 (N_13544,N_5010,N_4449);
or U13545 (N_13545,N_8596,N_8415);
or U13546 (N_13546,N_1417,N_998);
nand U13547 (N_13547,N_7892,N_2639);
nand U13548 (N_13548,N_9077,N_7355);
or U13549 (N_13549,N_3197,N_2819);
or U13550 (N_13550,N_3102,N_3959);
or U13551 (N_13551,N_9468,N_9875);
xor U13552 (N_13552,N_6294,N_1485);
nor U13553 (N_13553,N_9270,N_7411);
xor U13554 (N_13554,N_2931,N_8996);
nand U13555 (N_13555,N_1114,N_6722);
nor U13556 (N_13556,N_255,N_4035);
nand U13557 (N_13557,N_8412,N_7269);
nand U13558 (N_13558,N_5192,N_829);
or U13559 (N_13559,N_8882,N_7224);
nand U13560 (N_13560,N_472,N_345);
or U13561 (N_13561,N_8131,N_7754);
xor U13562 (N_13562,N_1316,N_7517);
and U13563 (N_13563,N_3849,N_2455);
or U13564 (N_13564,N_9160,N_5731);
nor U13565 (N_13565,N_5718,N_2227);
or U13566 (N_13566,N_1203,N_7895);
and U13567 (N_13567,N_7810,N_5273);
xor U13568 (N_13568,N_4521,N_2572);
and U13569 (N_13569,N_2510,N_5523);
nand U13570 (N_13570,N_6440,N_6048);
xor U13571 (N_13571,N_6439,N_27);
and U13572 (N_13572,N_4191,N_1382);
nor U13573 (N_13573,N_7609,N_7581);
nand U13574 (N_13574,N_7090,N_1542);
nor U13575 (N_13575,N_5915,N_9155);
nor U13576 (N_13576,N_5127,N_5309);
nor U13577 (N_13577,N_1103,N_949);
or U13578 (N_13578,N_115,N_7606);
nor U13579 (N_13579,N_8096,N_8715);
and U13580 (N_13580,N_3746,N_5724);
or U13581 (N_13581,N_2652,N_3004);
or U13582 (N_13582,N_7733,N_3556);
xnor U13583 (N_13583,N_310,N_4993);
nor U13584 (N_13584,N_7476,N_3176);
nor U13585 (N_13585,N_7455,N_1303);
and U13586 (N_13586,N_2003,N_6055);
nand U13587 (N_13587,N_1216,N_3703);
and U13588 (N_13588,N_3046,N_5529);
or U13589 (N_13589,N_1793,N_9827);
xor U13590 (N_13590,N_5690,N_1737);
or U13591 (N_13591,N_8572,N_7382);
or U13592 (N_13592,N_5381,N_9843);
nor U13593 (N_13593,N_4006,N_7563);
and U13594 (N_13594,N_7684,N_3512);
or U13595 (N_13595,N_4222,N_474);
nand U13596 (N_13596,N_9343,N_2544);
nor U13597 (N_13597,N_6392,N_956);
nor U13598 (N_13598,N_1019,N_5111);
nand U13599 (N_13599,N_2686,N_4718);
nor U13600 (N_13600,N_5047,N_2758);
nand U13601 (N_13601,N_7553,N_8695);
and U13602 (N_13602,N_3452,N_9555);
nor U13603 (N_13603,N_4249,N_8148);
and U13604 (N_13604,N_1493,N_1180);
xor U13605 (N_13605,N_8163,N_7283);
nor U13606 (N_13606,N_5324,N_4478);
nor U13607 (N_13607,N_6144,N_8707);
nor U13608 (N_13608,N_4780,N_6159);
nor U13609 (N_13609,N_484,N_6901);
xor U13610 (N_13610,N_5113,N_5240);
and U13611 (N_13611,N_3615,N_2625);
nand U13612 (N_13612,N_4832,N_1335);
and U13613 (N_13613,N_7506,N_8867);
nor U13614 (N_13614,N_5295,N_4564);
and U13615 (N_13615,N_5589,N_9668);
nand U13616 (N_13616,N_3074,N_2853);
nand U13617 (N_13617,N_249,N_24);
nand U13618 (N_13618,N_8878,N_4790);
nor U13619 (N_13619,N_6170,N_5556);
nor U13620 (N_13620,N_4503,N_9442);
nor U13621 (N_13621,N_5758,N_4835);
or U13622 (N_13622,N_4589,N_3179);
nor U13623 (N_13623,N_2415,N_9989);
nand U13624 (N_13624,N_1865,N_6189);
or U13625 (N_13625,N_9603,N_9696);
or U13626 (N_13626,N_5885,N_2927);
and U13627 (N_13627,N_4464,N_375);
or U13628 (N_13628,N_4563,N_8386);
nand U13629 (N_13629,N_3524,N_8769);
nand U13630 (N_13630,N_9044,N_8948);
nor U13631 (N_13631,N_4752,N_9605);
nor U13632 (N_13632,N_792,N_8810);
and U13633 (N_13633,N_7770,N_9770);
xnor U13634 (N_13634,N_3024,N_6643);
or U13635 (N_13635,N_5001,N_2814);
nand U13636 (N_13636,N_3868,N_5340);
and U13637 (N_13637,N_2126,N_4769);
or U13638 (N_13638,N_5105,N_4420);
nor U13639 (N_13639,N_1101,N_8189);
nand U13640 (N_13640,N_5912,N_9565);
nand U13641 (N_13641,N_7762,N_8241);
or U13642 (N_13642,N_2811,N_2826);
xor U13643 (N_13643,N_7327,N_2253);
xor U13644 (N_13644,N_9235,N_3410);
or U13645 (N_13645,N_1645,N_8416);
xor U13646 (N_13646,N_7313,N_161);
xnor U13647 (N_13647,N_893,N_7286);
and U13648 (N_13648,N_4082,N_8113);
nor U13649 (N_13649,N_1699,N_9769);
nor U13650 (N_13650,N_8621,N_3836);
nor U13651 (N_13651,N_2698,N_4056);
nand U13652 (N_13652,N_8907,N_130);
nor U13653 (N_13653,N_6500,N_9293);
or U13654 (N_13654,N_5688,N_3696);
nor U13655 (N_13655,N_8541,N_4900);
xor U13656 (N_13656,N_8017,N_3580);
nand U13657 (N_13657,N_3358,N_3248);
nor U13658 (N_13658,N_7307,N_4392);
or U13659 (N_13659,N_163,N_1089);
xnor U13660 (N_13660,N_5909,N_6346);
and U13661 (N_13661,N_5177,N_9985);
xnor U13662 (N_13662,N_5027,N_2634);
nand U13663 (N_13663,N_4080,N_1025);
nor U13664 (N_13664,N_8737,N_3975);
or U13665 (N_13665,N_7864,N_1033);
nor U13666 (N_13666,N_2524,N_2858);
nor U13667 (N_13667,N_5879,N_2729);
nor U13668 (N_13668,N_9236,N_2009);
nor U13669 (N_13669,N_8245,N_2665);
xor U13670 (N_13670,N_5973,N_5491);
nor U13671 (N_13671,N_7096,N_5154);
nand U13672 (N_13672,N_9240,N_2424);
xor U13673 (N_13673,N_1811,N_8823);
nor U13674 (N_13674,N_1924,N_4962);
xnor U13675 (N_13675,N_3125,N_7294);
nor U13676 (N_13676,N_8025,N_7254);
and U13677 (N_13677,N_6606,N_1941);
xnor U13678 (N_13678,N_771,N_4886);
nor U13679 (N_13679,N_4092,N_6546);
nor U13680 (N_13680,N_2576,N_1196);
xor U13681 (N_13681,N_2536,N_7912);
nor U13682 (N_13682,N_1477,N_6344);
nand U13683 (N_13683,N_4644,N_2979);
nor U13684 (N_13684,N_1713,N_2262);
nand U13685 (N_13685,N_2778,N_7168);
or U13686 (N_13686,N_8983,N_3845);
and U13687 (N_13687,N_9958,N_9231);
xnor U13688 (N_13688,N_7828,N_64);
and U13689 (N_13689,N_1061,N_9885);
and U13690 (N_13690,N_1564,N_1540);
nand U13691 (N_13691,N_8971,N_6103);
and U13692 (N_13692,N_2211,N_684);
and U13693 (N_13693,N_4180,N_3695);
xor U13694 (N_13694,N_4721,N_8855);
nor U13695 (N_13695,N_6551,N_9484);
and U13696 (N_13696,N_112,N_7103);
xnor U13697 (N_13697,N_8222,N_5066);
nand U13698 (N_13698,N_1824,N_3186);
xor U13699 (N_13699,N_4409,N_9040);
and U13700 (N_13700,N_858,N_2617);
and U13701 (N_13701,N_3816,N_7380);
nand U13702 (N_13702,N_4698,N_6087);
or U13703 (N_13703,N_2651,N_5164);
nor U13704 (N_13704,N_5620,N_633);
nor U13705 (N_13705,N_5665,N_9284);
nor U13706 (N_13706,N_1379,N_875);
xor U13707 (N_13707,N_1656,N_3707);
nor U13708 (N_13708,N_8562,N_667);
nand U13709 (N_13709,N_8449,N_1195);
and U13710 (N_13710,N_8351,N_4825);
and U13711 (N_13711,N_3411,N_1543);
or U13712 (N_13712,N_4177,N_9262);
nand U13713 (N_13713,N_1577,N_7016);
and U13714 (N_13714,N_2403,N_2547);
nand U13715 (N_13715,N_6670,N_7790);
nor U13716 (N_13716,N_2600,N_2308);
nor U13717 (N_13717,N_9281,N_4750);
nand U13718 (N_13718,N_9786,N_92);
nor U13719 (N_13719,N_615,N_1054);
nand U13720 (N_13720,N_7959,N_2505);
nand U13721 (N_13721,N_7596,N_9596);
or U13722 (N_13722,N_2887,N_2692);
nand U13723 (N_13723,N_812,N_2685);
xor U13724 (N_13724,N_3226,N_4108);
nor U13725 (N_13725,N_3021,N_2535);
and U13726 (N_13726,N_9661,N_9504);
xor U13727 (N_13727,N_3555,N_9572);
or U13728 (N_13728,N_9671,N_37);
nand U13729 (N_13729,N_6057,N_479);
and U13730 (N_13730,N_5123,N_7350);
nand U13731 (N_13731,N_8582,N_5833);
nor U13732 (N_13732,N_302,N_4845);
or U13733 (N_13733,N_8451,N_4217);
xor U13734 (N_13734,N_8585,N_3754);
or U13735 (N_13735,N_8483,N_5227);
or U13736 (N_13736,N_5280,N_8120);
nand U13737 (N_13737,N_4293,N_4187);
nor U13738 (N_13738,N_5186,N_2423);
or U13739 (N_13739,N_4729,N_947);
and U13740 (N_13740,N_382,N_5826);
or U13741 (N_13741,N_4498,N_2864);
nor U13742 (N_13742,N_8891,N_7330);
xnor U13743 (N_13743,N_6648,N_6380);
nor U13744 (N_13744,N_8108,N_9640);
or U13745 (N_13745,N_7819,N_3657);
nor U13746 (N_13746,N_9224,N_8776);
nor U13747 (N_13747,N_4095,N_2799);
and U13748 (N_13748,N_4984,N_7808);
nor U13749 (N_13749,N_3150,N_7271);
xor U13750 (N_13750,N_7600,N_6137);
nand U13751 (N_13751,N_3036,N_8549);
and U13752 (N_13752,N_7196,N_6447);
nor U13753 (N_13753,N_4612,N_8631);
and U13754 (N_13754,N_8212,N_5918);
and U13755 (N_13755,N_2358,N_1125);
xor U13756 (N_13756,N_4170,N_6660);
or U13757 (N_13757,N_3317,N_9908);
nor U13758 (N_13758,N_6280,N_3356);
or U13759 (N_13759,N_45,N_4244);
or U13760 (N_13760,N_2912,N_9564);
nand U13761 (N_13761,N_3736,N_4371);
or U13762 (N_13762,N_629,N_3989);
or U13763 (N_13763,N_8533,N_1944);
nand U13764 (N_13764,N_7824,N_8616);
and U13765 (N_13765,N_1999,N_2972);
xnor U13766 (N_13766,N_1672,N_849);
xor U13767 (N_13767,N_311,N_9643);
nor U13768 (N_13768,N_1582,N_3027);
nor U13769 (N_13769,N_11,N_8544);
and U13770 (N_13770,N_7332,N_3045);
or U13771 (N_13771,N_287,N_3761);
xnor U13772 (N_13772,N_7491,N_2202);
nand U13773 (N_13773,N_7404,N_1210);
xnor U13774 (N_13774,N_5840,N_1648);
nand U13775 (N_13775,N_6684,N_8418);
xor U13776 (N_13776,N_8712,N_7308);
nor U13777 (N_13777,N_4314,N_222);
nor U13778 (N_13778,N_9855,N_7831);
and U13779 (N_13779,N_13,N_4083);
nand U13780 (N_13780,N_3941,N_1040);
or U13781 (N_13781,N_885,N_1170);
nand U13782 (N_13782,N_7842,N_8194);
nor U13783 (N_13783,N_540,N_7351);
xor U13784 (N_13784,N_2991,N_9094);
or U13785 (N_13785,N_4196,N_5499);
and U13786 (N_13786,N_1345,N_3132);
or U13787 (N_13787,N_1808,N_7836);
nor U13788 (N_13788,N_7426,N_737);
xnor U13789 (N_13789,N_9701,N_4129);
or U13790 (N_13790,N_421,N_6028);
xnor U13791 (N_13791,N_9737,N_9493);
and U13792 (N_13792,N_4758,N_3827);
and U13793 (N_13793,N_5090,N_4120);
and U13794 (N_13794,N_6329,N_2603);
and U13795 (N_13795,N_4692,N_2939);
or U13796 (N_13796,N_6485,N_8603);
xor U13797 (N_13797,N_7030,N_9399);
nand U13798 (N_13798,N_9517,N_1842);
xnor U13799 (N_13799,N_6957,N_4637);
nand U13800 (N_13800,N_9982,N_8947);
and U13801 (N_13801,N_2542,N_1833);
and U13802 (N_13802,N_4659,N_2608);
nand U13803 (N_13803,N_5112,N_781);
nand U13804 (N_13804,N_3273,N_3364);
and U13805 (N_13805,N_424,N_8784);
or U13806 (N_13806,N_6563,N_6246);
nand U13807 (N_13807,N_4176,N_9889);
nand U13808 (N_13808,N_3502,N_5980);
and U13809 (N_13809,N_2357,N_1329);
nand U13810 (N_13810,N_7738,N_9338);
xor U13811 (N_13811,N_2567,N_2654);
nand U13812 (N_13812,N_1555,N_8510);
nor U13813 (N_13813,N_9401,N_8205);
nand U13814 (N_13814,N_4418,N_6939);
nor U13815 (N_13815,N_8015,N_7901);
nor U13816 (N_13816,N_2942,N_774);
nand U13817 (N_13817,N_9489,N_9914);
nor U13818 (N_13818,N_4691,N_7963);
and U13819 (N_13819,N_2569,N_5570);
nor U13820 (N_13820,N_5779,N_2248);
and U13821 (N_13821,N_8529,N_2688);
nor U13822 (N_13822,N_4801,N_9427);
or U13823 (N_13823,N_5486,N_3805);
nand U13824 (N_13824,N_9571,N_3075);
nor U13825 (N_13825,N_1889,N_2282);
and U13826 (N_13826,N_9393,N_7589);
nor U13827 (N_13827,N_1773,N_2624);
or U13828 (N_13828,N_8652,N_9073);
and U13829 (N_13829,N_9518,N_6044);
or U13830 (N_13830,N_3924,N_2515);
xnor U13831 (N_13831,N_4435,N_3454);
nor U13832 (N_13832,N_9580,N_6902);
nand U13833 (N_13833,N_9795,N_7950);
nor U13834 (N_13834,N_5150,N_1452);
nand U13835 (N_13835,N_1255,N_6368);
or U13836 (N_13836,N_9053,N_1823);
and U13837 (N_13837,N_5412,N_727);
nand U13838 (N_13838,N_3839,N_7232);
and U13839 (N_13839,N_2645,N_1765);
or U13840 (N_13840,N_5716,N_5236);
xnor U13841 (N_13841,N_2448,N_7677);
nand U13842 (N_13842,N_5237,N_9990);
or U13843 (N_13843,N_8142,N_6991);
xnor U13844 (N_13844,N_6739,N_7315);
or U13845 (N_13845,N_8503,N_8374);
xnor U13846 (N_13846,N_4796,N_4996);
nand U13847 (N_13847,N_4873,N_8654);
nor U13848 (N_13848,N_374,N_4451);
or U13849 (N_13849,N_7386,N_7943);
xor U13850 (N_13850,N_6735,N_8461);
xnor U13851 (N_13851,N_5384,N_974);
nand U13852 (N_13852,N_7611,N_8213);
nor U13853 (N_13853,N_8502,N_8448);
or U13854 (N_13854,N_2854,N_8154);
nor U13855 (N_13855,N_6734,N_4946);
or U13856 (N_13856,N_3689,N_9126);
nand U13857 (N_13857,N_1826,N_7177);
or U13858 (N_13858,N_754,N_7965);
nand U13859 (N_13859,N_6201,N_8143);
xor U13860 (N_13860,N_8405,N_9514);
or U13861 (N_13861,N_3058,N_6601);
and U13862 (N_13862,N_7198,N_7716);
nor U13863 (N_13863,N_2556,N_7219);
or U13864 (N_13864,N_3563,N_2076);
xnor U13865 (N_13865,N_5410,N_4561);
nor U13866 (N_13866,N_8430,N_3216);
nand U13867 (N_13867,N_4406,N_9687);
or U13868 (N_13868,N_2329,N_4090);
nand U13869 (N_13869,N_5011,N_8378);
xnor U13870 (N_13870,N_715,N_9130);
nor U13871 (N_13871,N_1220,N_2157);
xnor U13872 (N_13872,N_9018,N_2764);
xnor U13873 (N_13873,N_7093,N_6123);
nand U13874 (N_13874,N_1227,N_5800);
nand U13875 (N_13875,N_6305,N_4604);
nand U13876 (N_13876,N_9086,N_3222);
or U13877 (N_13877,N_4504,N_7489);
xnor U13878 (N_13878,N_181,N_8628);
nor U13879 (N_13879,N_2584,N_4114);
xor U13880 (N_13880,N_9097,N_624);
nor U13881 (N_13881,N_894,N_2551);
xor U13882 (N_13882,N_592,N_6851);
or U13883 (N_13883,N_5981,N_8814);
xnor U13884 (N_13884,N_3326,N_9829);
nor U13885 (N_13885,N_7974,N_1728);
nor U13886 (N_13886,N_1853,N_9178);
nor U13887 (N_13887,N_4546,N_3256);
and U13888 (N_13888,N_3319,N_4145);
xnor U13889 (N_13889,N_9540,N_2789);
and U13890 (N_13890,N_2929,N_7228);
nand U13891 (N_13891,N_1473,N_5541);
or U13892 (N_13892,N_8287,N_7940);
and U13893 (N_13893,N_6928,N_7123);
and U13894 (N_13894,N_808,N_5297);
or U13895 (N_13895,N_1118,N_109);
or U13896 (N_13896,N_5757,N_3911);
and U13897 (N_13897,N_6599,N_871);
xnor U13898 (N_13898,N_5756,N_1857);
or U13899 (N_13899,N_356,N_9299);
or U13900 (N_13900,N_7218,N_5274);
or U13901 (N_13901,N_8615,N_1454);
and U13902 (N_13902,N_7794,N_6468);
nand U13903 (N_13903,N_4897,N_4288);
nand U13904 (N_13904,N_9219,N_3654);
nand U13905 (N_13905,N_8201,N_8846);
nand U13906 (N_13906,N_5831,N_3283);
nand U13907 (N_13907,N_8665,N_5679);
nand U13908 (N_13908,N_2327,N_3396);
nand U13909 (N_13909,N_6446,N_5669);
or U13910 (N_13910,N_9050,N_1972);
xnor U13911 (N_13911,N_1925,N_3201);
or U13912 (N_13912,N_993,N_640);
xor U13913 (N_13913,N_879,N_5846);
and U13914 (N_13914,N_2420,N_5021);
and U13915 (N_13915,N_304,N_8123);
or U13916 (N_13916,N_5480,N_3891);
nand U13917 (N_13917,N_8291,N_1416);
or U13918 (N_13918,N_413,N_3697);
nand U13919 (N_13919,N_9693,N_7717);
xnor U13920 (N_13920,N_1302,N_7862);
or U13921 (N_13921,N_9933,N_8930);
nor U13922 (N_13922,N_9464,N_7659);
or U13923 (N_13923,N_631,N_4439);
nor U13924 (N_13924,N_6051,N_4771);
xnor U13925 (N_13925,N_1747,N_9132);
and U13926 (N_13926,N_5430,N_6534);
nand U13927 (N_13927,N_8305,N_8484);
nor U13928 (N_13928,N_934,N_3162);
or U13929 (N_13929,N_8091,N_477);
and U13930 (N_13930,N_8052,N_4342);
nor U13931 (N_13931,N_1859,N_6757);
nor U13932 (N_13932,N_2022,N_5013);
and U13933 (N_13933,N_7858,N_555);
and U13934 (N_13934,N_4749,N_7758);
nand U13935 (N_13935,N_4004,N_9385);
and U13936 (N_13936,N_6415,N_6349);
xor U13937 (N_13937,N_570,N_1836);
or U13938 (N_13938,N_7729,N_9852);
and U13939 (N_13939,N_2943,N_1682);
and U13940 (N_13940,N_137,N_6033);
and U13941 (N_13941,N_1660,N_8027);
or U13942 (N_13942,N_1943,N_1881);
nor U13943 (N_13943,N_6216,N_4213);
nand U13944 (N_13944,N_4697,N_5873);
and U13945 (N_13945,N_5492,N_3655);
nor U13946 (N_13946,N_1804,N_5894);
and U13947 (N_13947,N_7067,N_8729);
nand U13948 (N_13948,N_1772,N_6035);
or U13949 (N_13949,N_7216,N_6845);
and U13950 (N_13950,N_3993,N_7192);
xnor U13951 (N_13951,N_6613,N_1116);
nor U13952 (N_13952,N_1157,N_1608);
nand U13953 (N_13953,N_2492,N_8265);
nand U13954 (N_13954,N_3595,N_3439);
nor U13955 (N_13955,N_1949,N_9842);
nor U13956 (N_13956,N_4419,N_4481);
and U13957 (N_13957,N_6223,N_568);
and U13958 (N_13958,N_2601,N_1641);
nand U13959 (N_13959,N_5085,N_7203);
xor U13960 (N_13960,N_5744,N_7468);
or U13961 (N_13961,N_6424,N_8357);
or U13962 (N_13962,N_9036,N_698);
xor U13963 (N_13963,N_9754,N_2553);
nor U13964 (N_13964,N_6013,N_2981);
and U13965 (N_13965,N_900,N_7816);
nand U13966 (N_13966,N_2333,N_5948);
nand U13967 (N_13967,N_2173,N_1407);
nand U13968 (N_13968,N_6252,N_346);
or U13969 (N_13969,N_6730,N_3511);
and U13970 (N_13970,N_5284,N_7926);
or U13971 (N_13971,N_607,N_4063);
nor U13972 (N_13972,N_5205,N_1141);
or U13973 (N_13973,N_1038,N_9275);
nand U13974 (N_13974,N_6746,N_598);
and U13975 (N_13975,N_6552,N_2331);
and U13976 (N_13976,N_4458,N_8250);
nand U13977 (N_13977,N_6078,N_7340);
nor U13978 (N_13978,N_8517,N_280);
nor U13979 (N_13979,N_499,N_9491);
or U13980 (N_13980,N_6204,N_5715);
xnor U13981 (N_13981,N_5938,N_6481);
nand U13982 (N_13982,N_1702,N_4660);
xnor U13983 (N_13983,N_5906,N_9531);
or U13984 (N_13984,N_6131,N_8868);
and U13985 (N_13985,N_4434,N_761);
nor U13986 (N_13986,N_432,N_3450);
xnor U13987 (N_13987,N_8434,N_8237);
or U13988 (N_13988,N_7321,N_4055);
and U13989 (N_13989,N_4894,N_6382);
xnor U13990 (N_13990,N_6317,N_1432);
and U13991 (N_13991,N_9520,N_7023);
and U13992 (N_13992,N_3521,N_6095);
and U13993 (N_13993,N_8852,N_1132);
or U13994 (N_13994,N_6937,N_2975);
xor U13995 (N_13995,N_1499,N_1096);
and U13996 (N_13996,N_8349,N_9099);
nand U13997 (N_13997,N_2976,N_7815);
xor U13998 (N_13998,N_1392,N_8137);
and U13999 (N_13999,N_4100,N_2195);
and U14000 (N_14000,N_4133,N_5433);
or U14001 (N_14001,N_8443,N_7256);
nor U14002 (N_14002,N_9835,N_7829);
xor U14003 (N_14003,N_1723,N_3163);
and U14004 (N_14004,N_113,N_8547);
xnor U14005 (N_14005,N_2368,N_7768);
xor U14006 (N_14006,N_3940,N_1845);
and U14007 (N_14007,N_3295,N_8755);
nor U14008 (N_14008,N_809,N_1475);
and U14009 (N_14009,N_5822,N_4870);
nor U14010 (N_14010,N_855,N_1010);
nand U14011 (N_14011,N_8324,N_2720);
xor U14012 (N_14012,N_712,N_8733);
or U14013 (N_14013,N_8009,N_680);
nor U14014 (N_14014,N_6628,N_1185);
nor U14015 (N_14015,N_7400,N_1349);
xnor U14016 (N_14016,N_3645,N_8526);
or U14017 (N_14017,N_7513,N_89);
nor U14018 (N_14018,N_7187,N_1940);
xnor U14019 (N_14019,N_4320,N_5043);
nand U14020 (N_14020,N_2709,N_1098);
nand U14021 (N_14021,N_2677,N_798);
nand U14022 (N_14022,N_7760,N_1628);
xnor U14023 (N_14023,N_199,N_4945);
and U14024 (N_14024,N_899,N_674);
nand U14025 (N_14025,N_8440,N_2859);
nand U14026 (N_14026,N_6437,N_3421);
nand U14027 (N_14027,N_7111,N_7601);
nand U14028 (N_14028,N_5201,N_9297);
or U14029 (N_14029,N_5109,N_4207);
nand U14030 (N_14030,N_6594,N_1062);
and U14031 (N_14031,N_2402,N_4590);
nand U14032 (N_14032,N_4569,N_986);
or U14033 (N_14033,N_3266,N_2590);
nand U14034 (N_14034,N_5962,N_8464);
or U14035 (N_14035,N_783,N_884);
xnor U14036 (N_14036,N_3040,N_582);
or U14037 (N_14037,N_1153,N_7408);
nand U14038 (N_14038,N_4617,N_1470);
or U14039 (N_14039,N_1338,N_6370);
nor U14040 (N_14040,N_5908,N_9913);
nand U14041 (N_14041,N_3999,N_3494);
xnor U14042 (N_14042,N_3961,N_7561);
nand U14043 (N_14043,N_1863,N_7571);
or U14044 (N_14044,N_8667,N_8857);
nor U14045 (N_14045,N_8933,N_3988);
nor U14046 (N_14046,N_1982,N_5012);
xor U14047 (N_14047,N_9055,N_7179);
and U14048 (N_14048,N_547,N_340);
and U14049 (N_14049,N_6885,N_3987);
xnor U14050 (N_14050,N_6529,N_4124);
or U14051 (N_14051,N_15,N_6597);
nand U14052 (N_14052,N_6198,N_6689);
and U14053 (N_14053,N_490,N_1065);
and U14054 (N_14054,N_8932,N_1588);
nor U14055 (N_14055,N_8341,N_821);
or U14056 (N_14056,N_6530,N_281);
and U14057 (N_14057,N_6541,N_465);
nand U14058 (N_14058,N_2185,N_9043);
and U14059 (N_14059,N_8127,N_7106);
xnor U14060 (N_14060,N_5035,N_5785);
nand U14061 (N_14061,N_7645,N_3199);
nor U14062 (N_14062,N_2869,N_5890);
and U14063 (N_14063,N_1420,N_1218);
and U14064 (N_14064,N_9025,N_9292);
or U14065 (N_14065,N_8010,N_1967);
nor U14066 (N_14066,N_6388,N_3207);
and U14067 (N_14067,N_9904,N_8563);
nand U14068 (N_14068,N_7423,N_6323);
and U14069 (N_14069,N_1727,N_1522);
nand U14070 (N_14070,N_1525,N_9028);
nor U14071 (N_14071,N_1979,N_920);
or U14072 (N_14072,N_9856,N_1763);
and U14073 (N_14073,N_8413,N_6165);
and U14074 (N_14074,N_3533,N_5069);
nand U14075 (N_14075,N_3759,N_6278);
and U14076 (N_14076,N_7366,N_6632);
and U14077 (N_14077,N_2053,N_5437);
xnor U14078 (N_14078,N_4805,N_3070);
xor U14079 (N_14079,N_4022,N_1715);
xor U14080 (N_14080,N_2034,N_2024);
nand U14081 (N_14081,N_5279,N_2153);
or U14082 (N_14082,N_9677,N_8019);
xor U14083 (N_14083,N_6119,N_350);
xor U14084 (N_14084,N_3815,N_258);
xor U14085 (N_14085,N_8135,N_2462);
nand U14086 (N_14086,N_927,N_3540);
nand U14087 (N_14087,N_4577,N_5400);
nand U14088 (N_14088,N_556,N_5787);
nand U14089 (N_14089,N_7473,N_3818);
xor U14090 (N_14090,N_8355,N_275);
nand U14091 (N_14091,N_7385,N_5544);
xnor U14092 (N_14092,N_8471,N_4879);
nand U14093 (N_14093,N_2803,N_9107);
xor U14094 (N_14094,N_6293,N_6237);
nor U14095 (N_14095,N_9156,N_7171);
nor U14096 (N_14096,N_34,N_330);
xnor U14097 (N_14097,N_8115,N_29);
xor U14098 (N_14098,N_6180,N_1689);
nand U14099 (N_14099,N_8721,N_3584);
nand U14100 (N_14100,N_2084,N_1457);
or U14101 (N_14101,N_9920,N_6407);
nand U14102 (N_14102,N_7755,N_4531);
nor U14103 (N_14103,N_7205,N_1231);
nor U14104 (N_14104,N_3788,N_1447);
nand U14105 (N_14105,N_5953,N_6414);
nand U14106 (N_14106,N_8395,N_9379);
nor U14107 (N_14107,N_8309,N_589);
xor U14108 (N_14108,N_2922,N_3562);
nand U14109 (N_14109,N_7342,N_5173);
nand U14110 (N_14110,N_7475,N_5856);
and U14111 (N_14111,N_8272,N_1122);
xnor U14112 (N_14112,N_3306,N_3561);
nand U14113 (N_14113,N_2641,N_4625);
or U14114 (N_14114,N_8584,N_2788);
xnor U14115 (N_14115,N_3420,N_1086);
and U14116 (N_14116,N_5310,N_1998);
xnor U14117 (N_14117,N_208,N_9773);
and U14118 (N_14118,N_6811,N_1189);
nand U14119 (N_14119,N_3554,N_5976);
or U14120 (N_14120,N_9064,N_886);
xnor U14121 (N_14121,N_7727,N_2143);
or U14122 (N_14122,N_6381,N_8259);
xor U14123 (N_14123,N_2494,N_2957);
and U14124 (N_14124,N_6295,N_2028);
xnor U14125 (N_14125,N_9720,N_1847);
nor U14126 (N_14126,N_5143,N_8175);
xor U14127 (N_14127,N_8366,N_4684);
nor U14128 (N_14128,N_3834,N_3249);
or U14129 (N_14129,N_4787,N_1188);
nor U14130 (N_14130,N_7673,N_7848);
and U14131 (N_14131,N_4981,N_881);
nand U14132 (N_14132,N_334,N_6056);
and U14133 (N_14133,N_2531,N_1858);
nor U14134 (N_14134,N_6692,N_6950);
and U14135 (N_14135,N_9302,N_1484);
and U14136 (N_14136,N_6572,N_8419);
xor U14137 (N_14137,N_945,N_23);
or U14138 (N_14138,N_1039,N_9416);
and U14139 (N_14139,N_6112,N_2011);
or U14140 (N_14140,N_3457,N_6393);
xor U14141 (N_14141,N_2219,N_2438);
or U14142 (N_14142,N_6867,N_411);
and U14143 (N_14143,N_925,N_2575);
or U14144 (N_14144,N_8486,N_8611);
nand U14145 (N_14145,N_7899,N_8861);
nand U14146 (N_14146,N_2676,N_3292);
nor U14147 (N_14147,N_5080,N_8845);
and U14148 (N_14148,N_5998,N_3261);
nand U14149 (N_14149,N_3596,N_1920);
or U14150 (N_14150,N_9823,N_300);
xnor U14151 (N_14151,N_7989,N_7247);
nand U14152 (N_14152,N_2950,N_1355);
nor U14153 (N_14153,N_7586,N_3240);
nor U14154 (N_14154,N_757,N_8038);
or U14155 (N_14155,N_1330,N_8008);
xnor U14156 (N_14156,N_3282,N_8100);
nand U14157 (N_14157,N_6441,N_5884);
nor U14158 (N_14158,N_5509,N_979);
or U14159 (N_14159,N_1235,N_53);
xor U14160 (N_14160,N_2370,N_3920);
or U14161 (N_14161,N_205,N_380);
nand U14162 (N_14162,N_1075,N_1056);
nor U14163 (N_14163,N_1356,N_9953);
and U14164 (N_14164,N_5326,N_5487);
xnor U14165 (N_14165,N_4370,N_1497);
or U14166 (N_14166,N_4412,N_9575);
and U14167 (N_14167,N_7610,N_9778);
and U14168 (N_14168,N_3621,N_9306);
or U14169 (N_14169,N_3313,N_892);
xor U14170 (N_14170,N_4266,N_6335);
xor U14171 (N_14171,N_9534,N_2399);
nand U14172 (N_14172,N_2486,N_385);
xor U14173 (N_14173,N_2691,N_5638);
nor U14174 (N_14174,N_750,N_6948);
nand U14175 (N_14175,N_2352,N_9198);
nor U14176 (N_14176,N_8842,N_8177);
and U14177 (N_14177,N_8967,N_8129);
or U14178 (N_14178,N_1340,N_3006);
and U14179 (N_14179,N_6501,N_6167);
nor U14180 (N_14180,N_751,N_2993);
or U14181 (N_14181,N_1625,N_2901);
and U14182 (N_14182,N_1337,N_2528);
nand U14183 (N_14183,N_4033,N_9898);
nor U14184 (N_14184,N_5424,N_7580);
nor U14185 (N_14185,N_4457,N_6465);
nor U14186 (N_14186,N_6604,N_7194);
xor U14187 (N_14187,N_2731,N_6537);
nand U14188 (N_14188,N_7867,N_7751);
nand U14189 (N_14189,N_6313,N_8049);
and U14190 (N_14190,N_1283,N_6444);
xnor U14191 (N_14191,N_7850,N_5351);
or U14192 (N_14192,N_8797,N_733);
nor U14193 (N_14193,N_5115,N_9606);
or U14194 (N_14194,N_1074,N_7583);
xnor U14195 (N_14195,N_2478,N_3700);
nand U14196 (N_14196,N_7647,N_2377);
and U14197 (N_14197,N_1233,N_4671);
and U14198 (N_14198,N_3342,N_2260);
nand U14199 (N_14199,N_9376,N_4719);
nor U14200 (N_14200,N_4126,N_4628);
or U14201 (N_14201,N_9947,N_6114);
nor U14202 (N_14202,N_7211,N_6146);
nand U14203 (N_14203,N_874,N_2627);
nor U14204 (N_14204,N_7818,N_5820);
nor U14205 (N_14205,N_468,N_2317);
xnor U14206 (N_14206,N_9768,N_5092);
and U14207 (N_14207,N_4008,N_6870);
nor U14208 (N_14208,N_467,N_1514);
xnor U14209 (N_14209,N_7728,N_2167);
or U14210 (N_14210,N_9752,N_4597);
xnor U14211 (N_14211,N_2770,N_1079);
or U14212 (N_14212,N_8566,N_2097);
xnor U14213 (N_14213,N_8795,N_2056);
nor U14214 (N_14214,N_4161,N_3627);
nor U14215 (N_14215,N_3964,N_9620);
xor U14216 (N_14216,N_1331,N_2447);
or U14217 (N_14217,N_3579,N_3145);
and U14218 (N_14218,N_9005,N_3526);
xnor U14219 (N_14219,N_7034,N_3508);
or U14220 (N_14220,N_3833,N_407);
or U14221 (N_14221,N_2582,N_7908);
and U14222 (N_14222,N_5551,N_3977);
nand U14223 (N_14223,N_9782,N_8263);
or U14224 (N_14224,N_7756,N_3953);
nand U14225 (N_14225,N_5307,N_7450);
nand U14226 (N_14226,N_2837,N_3137);
and U14227 (N_14227,N_9528,N_741);
nor U14228 (N_14228,N_654,N_4076);
nand U14229 (N_14229,N_538,N_342);
and U14230 (N_14230,N_2664,N_6931);
nand U14231 (N_14231,N_9118,N_2272);
nor U14232 (N_14232,N_2263,N_8841);
or U14233 (N_14233,N_8679,N_5664);
xor U14234 (N_14234,N_5094,N_1966);
xnor U14235 (N_14235,N_4052,N_3522);
xnor U14236 (N_14236,N_5612,N_2194);
xor U14237 (N_14237,N_1149,N_5629);
xor U14238 (N_14238,N_5288,N_43);
nand U14239 (N_14239,N_8647,N_9423);
nand U14240 (N_14240,N_7964,N_9624);
and U14241 (N_14241,N_1244,N_9944);
and U14242 (N_14242,N_1445,N_7259);
and U14243 (N_14243,N_1539,N_7971);
or U14244 (N_14244,N_8697,N_7837);
nor U14245 (N_14245,N_3406,N_9940);
or U14246 (N_14246,N_9321,N_221);
and U14247 (N_14247,N_2997,N_7577);
xnor U14248 (N_14248,N_8039,N_7022);
nor U14249 (N_14249,N_8778,N_8023);
nor U14250 (N_14250,N_4190,N_2382);
nand U14251 (N_14251,N_9474,N_1899);
and U14252 (N_14252,N_6306,N_4795);
or U14253 (N_14253,N_5388,N_372);
and U14254 (N_14254,N_5162,N_1228);
xnor U14255 (N_14255,N_8620,N_8767);
xnor U14256 (N_14256,N_9184,N_190);
nor U14257 (N_14257,N_2378,N_6396);
or U14258 (N_14258,N_2490,N_1800);
and U14259 (N_14259,N_2483,N_1812);
or U14260 (N_14260,N_4499,N_1398);
nor U14261 (N_14261,N_2323,N_522);
nor U14262 (N_14262,N_4270,N_6384);
nand U14263 (N_14263,N_6732,N_9804);
and U14264 (N_14264,N_2920,N_4311);
and U14265 (N_14265,N_5132,N_8602);
and U14266 (N_14266,N_8467,N_9279);
and U14267 (N_14267,N_2517,N_1792);
nand U14268 (N_14268,N_857,N_7244);
nand U14269 (N_14269,N_2836,N_2684);
and U14270 (N_14270,N_1549,N_1639);
nor U14271 (N_14271,N_3478,N_8573);
xor U14272 (N_14272,N_6353,N_4767);
or U14273 (N_14273,N_8872,N_7980);
nor U14274 (N_14274,N_7585,N_7365);
xor U14275 (N_14275,N_3079,N_6175);
or U14276 (N_14276,N_1670,N_972);
nor U14277 (N_14277,N_8334,N_7042);
and U14278 (N_14278,N_455,N_9883);
and U14279 (N_14279,N_307,N_1673);
xnor U14280 (N_14280,N_9266,N_3572);
nand U14281 (N_14281,N_8747,N_2747);
nand U14282 (N_14282,N_1051,N_4568);
or U14283 (N_14283,N_2404,N_9305);
and U14284 (N_14284,N_9342,N_166);
xnor U14285 (N_14285,N_7736,N_5270);
nand U14286 (N_14286,N_8521,N_5413);
nand U14287 (N_14287,N_6117,N_7658);
nor U14288 (N_14288,N_578,N_6825);
nor U14289 (N_14289,N_8660,N_1250);
nor U14290 (N_14290,N_3181,N_5858);
or U14291 (N_14291,N_2213,N_9541);
xnor U14292 (N_14292,N_9102,N_8678);
and U14293 (N_14293,N_2347,N_1035);
nor U14294 (N_14294,N_247,N_2726);
or U14295 (N_14295,N_25,N_9830);
or U14296 (N_14296,N_3083,N_4109);
nor U14297 (N_14297,N_2875,N_2183);
or U14298 (N_14298,N_1506,N_3353);
and U14299 (N_14299,N_2485,N_1159);
xor U14300 (N_14300,N_6290,N_3620);
xor U14301 (N_14301,N_4860,N_3367);
and U14302 (N_14302,N_6817,N_6740);
xor U14303 (N_14303,N_7798,N_8774);
and U14304 (N_14304,N_3876,N_6590);
nand U14305 (N_14305,N_5304,N_5707);
and U14306 (N_14306,N_4836,N_4516);
nand U14307 (N_14307,N_2476,N_6698);
and U14308 (N_14308,N_7118,N_5378);
and U14309 (N_14309,N_194,N_1239);
nand U14310 (N_14310,N_9065,N_7398);
xnor U14311 (N_14311,N_7665,N_9630);
and U14312 (N_14312,N_6426,N_3838);
nor U14313 (N_14313,N_2882,N_3857);
and U14314 (N_14314,N_5880,N_3811);
and U14315 (N_14315,N_8554,N_9428);
or U14316 (N_14316,N_3086,N_7975);
nor U14317 (N_14317,N_617,N_1275);
nand U14318 (N_14318,N_7888,N_3534);
and U14319 (N_14319,N_6545,N_1381);
nand U14320 (N_14320,N_1850,N_4162);
xor U14321 (N_14321,N_2429,N_5135);
or U14322 (N_14322,N_8323,N_8772);
nor U14323 (N_14323,N_4292,N_5987);
and U14324 (N_14324,N_7967,N_4602);
nor U14325 (N_14325,N_7376,N_185);
or U14326 (N_14326,N_9522,N_8459);
nor U14327 (N_14327,N_6920,N_3613);
or U14328 (N_14328,N_1755,N_6421);
or U14329 (N_14329,N_7540,N_3453);
nand U14330 (N_14330,N_984,N_8229);
nand U14331 (N_14331,N_6408,N_1423);
or U14332 (N_14332,N_8304,N_1113);
xor U14333 (N_14333,N_9181,N_9134);
nor U14334 (N_14334,N_1472,N_48);
xor U14335 (N_14335,N_7872,N_7329);
nand U14336 (N_14336,N_5020,N_3276);
nor U14337 (N_14337,N_1594,N_5028);
nor U14338 (N_14338,N_8462,N_639);
nand U14339 (N_14339,N_6664,N_987);
or U14340 (N_14340,N_2669,N_8109);
and U14341 (N_14341,N_1746,N_780);
or U14342 (N_14342,N_2035,N_2905);
and U14343 (N_14343,N_6918,N_609);
xor U14344 (N_14344,N_7494,N_7217);
xor U14345 (N_14345,N_5798,N_3628);
and U14346 (N_14346,N_5887,N_1198);
or U14347 (N_14347,N_3932,N_6301);
or U14348 (N_14348,N_500,N_6245);
and U14349 (N_14349,N_6276,N_3477);
nand U14350 (N_14350,N_8961,N_182);
xor U14351 (N_14351,N_9444,N_8363);
or U14352 (N_14352,N_7432,N_2621);
xnor U14353 (N_14353,N_4274,N_2334);
nor U14354 (N_14354,N_5087,N_4015);
nand U14355 (N_14355,N_4195,N_4209);
xnor U14356 (N_14356,N_6808,N_8504);
nor U14357 (N_14357,N_9547,N_580);
xor U14358 (N_14358,N_4918,N_824);
nand U14359 (N_14359,N_5767,N_2856);
nor U14360 (N_14360,N_5106,N_9164);
nor U14361 (N_14361,N_2025,N_4985);
and U14362 (N_14362,N_4987,N_4849);
and U14363 (N_14363,N_4343,N_3516);
or U14364 (N_14364,N_6831,N_5789);
or U14365 (N_14365,N_363,N_9713);
nand U14366 (N_14366,N_7158,N_8636);
nand U14367 (N_14367,N_6116,N_3196);
xnor U14368 (N_14368,N_3923,N_3015);
xor U14369 (N_14369,N_1827,N_9957);
nor U14370 (N_14370,N_8754,N_2838);
nand U14371 (N_14371,N_5359,N_2605);
xor U14372 (N_14372,N_5253,N_8844);
xor U14373 (N_14373,N_1182,N_9832);
and U14374 (N_14374,N_9999,N_910);
or U14375 (N_14375,N_6846,N_1438);
and U14376 (N_14376,N_3084,N_33);
or U14377 (N_14377,N_7745,N_5382);
xor U14378 (N_14378,N_8630,N_9613);
nand U14379 (N_14379,N_5747,N_3190);
nor U14380 (N_14380,N_4515,N_2191);
nor U14381 (N_14381,N_119,N_6341);
or U14382 (N_14382,N_8974,N_734);
and U14383 (N_14383,N_3981,N_4802);
or U14384 (N_14384,N_7550,N_7579);
and U14385 (N_14385,N_5229,N_9412);
and U14386 (N_14386,N_4214,N_5183);
and U14387 (N_14387,N_7675,N_1328);
nor U14388 (N_14388,N_3906,N_1997);
nor U14389 (N_14389,N_5165,N_6967);
nor U14390 (N_14390,N_4831,N_5054);
nor U14391 (N_14391,N_6849,N_6449);
and U14392 (N_14392,N_9233,N_5281);
nand U14393 (N_14393,N_6938,N_7362);
nor U14394 (N_14394,N_8749,N_2291);
nand U14395 (N_14395,N_5151,N_6683);
nand U14396 (N_14396,N_4466,N_8559);
nand U14397 (N_14397,N_7838,N_7360);
nand U14398 (N_14398,N_1942,N_7720);
xnor U14399 (N_14399,N_5816,N_4107);
and U14400 (N_14400,N_5044,N_5442);
xnor U14401 (N_14401,N_4188,N_5016);
nor U14402 (N_14402,N_214,N_4025);
and U14403 (N_14403,N_8185,N_4496);
or U14404 (N_14404,N_9590,N_5306);
and U14405 (N_14405,N_7565,N_3191);
and U14406 (N_14406,N_9950,N_3950);
and U14407 (N_14407,N_351,N_379);
nand U14408 (N_14408,N_8727,N_7334);
or U14409 (N_14409,N_1085,N_8696);
and U14410 (N_14410,N_8026,N_2932);
xor U14411 (N_14411,N_6947,N_714);
nand U14412 (N_14412,N_5792,N_5244);
nand U14413 (N_14413,N_9682,N_1839);
nand U14414 (N_14414,N_6231,N_508);
and U14415 (N_14415,N_5843,N_7664);
xnor U14416 (N_14416,N_1012,N_5876);
and U14417 (N_14417,N_2839,N_7788);
or U14418 (N_14418,N_133,N_2409);
nand U14419 (N_14419,N_369,N_9700);
and U14420 (N_14420,N_6786,N_6955);
nand U14421 (N_14421,N_9991,N_4097);
nand U14422 (N_14422,N_3441,N_8167);
nand U14423 (N_14423,N_6753,N_5794);
nor U14424 (N_14424,N_1341,N_6919);
xor U14425 (N_14425,N_2154,N_2257);
nor U14426 (N_14426,N_6536,N_6770);
nand U14427 (N_14427,N_1488,N_553);
and U14428 (N_14428,N_7813,N_8124);
nor U14429 (N_14429,N_4156,N_8227);
xnor U14430 (N_14430,N_2020,N_1530);
xor U14431 (N_14431,N_8472,N_2453);
or U14432 (N_14432,N_2599,N_1671);
xor U14433 (N_14433,N_895,N_9022);
xnor U14434 (N_14434,N_1433,N_7913);
or U14435 (N_14435,N_6017,N_7260);
nand U14436 (N_14436,N_1419,N_8890);
or U14437 (N_14437,N_533,N_6964);
or U14438 (N_14438,N_8698,N_8646);
xnor U14439 (N_14439,N_4447,N_1884);
nor U14440 (N_14440,N_3028,N_1002);
or U14441 (N_14441,N_865,N_567);
nor U14442 (N_14442,N_1193,N_4002);
or U14443 (N_14443,N_7163,N_285);
nor U14444 (N_14444,N_3398,N_443);
nor U14445 (N_14445,N_864,N_4851);
and U14446 (N_14446,N_6514,N_1801);
or U14447 (N_14447,N_1258,N_7124);
xnor U14448 (N_14448,N_9776,N_4205);
nand U14449 (N_14449,N_7749,N_3749);
or U14450 (N_14450,N_3824,N_7567);
nand U14451 (N_14451,N_2366,N_7125);
and U14452 (N_14452,N_5992,N_7542);
nor U14453 (N_14453,N_8735,N_4039);
and U14454 (N_14454,N_6233,N_7150);
or U14455 (N_14455,N_765,N_8332);
xnor U14456 (N_14456,N_2808,N_4593);
nor U14457 (N_14457,N_9753,N_7019);
nor U14458 (N_14458,N_3100,N_3347);
and U14459 (N_14459,N_1580,N_708);
nand U14460 (N_14460,N_8952,N_6641);
nor U14461 (N_14461,N_8268,N_7648);
nand U14462 (N_14462,N_481,N_7604);
xnor U14463 (N_14463,N_4963,N_5900);
nor U14464 (N_14464,N_3227,N_7461);
nand U14465 (N_14465,N_7418,N_8238);
xor U14466 (N_14466,N_1011,N_1815);
nor U14467 (N_14467,N_9703,N_252);
or U14468 (N_14468,N_7725,N_107);
nand U14469 (N_14469,N_6121,N_9382);
nand U14470 (N_14470,N_8684,N_6569);
nor U14471 (N_14471,N_5398,N_665);
or U14472 (N_14472,N_1489,N_9848);
xor U14473 (N_14473,N_9083,N_3658);
or U14474 (N_14474,N_5414,N_6422);
nand U14475 (N_14475,N_1429,N_2396);
xor U14476 (N_14476,N_841,N_7298);
xnor U14477 (N_14477,N_4446,N_1371);
nor U14478 (N_14478,N_1851,N_1430);
nor U14479 (N_14479,N_8833,N_6291);
nand U14480 (N_14480,N_473,N_1181);
or U14481 (N_14481,N_6715,N_613);
xor U14482 (N_14482,N_5125,N_9615);
xor U14483 (N_14483,N_8147,N_7045);
xnor U14484 (N_14484,N_1697,N_4356);
or U14485 (N_14485,N_7478,N_4118);
xnor U14486 (N_14486,N_9010,N_6657);
or U14487 (N_14487,N_1391,N_6411);
and U14488 (N_14488,N_8226,N_4070);
nand U14489 (N_14489,N_5023,N_5076);
or U14490 (N_14490,N_9633,N_8333);
nor U14491 (N_14491,N_3629,N_6495);
and U14492 (N_14492,N_8151,N_8488);
nand U14493 (N_14493,N_9871,N_2681);
nor U14494 (N_14494,N_7812,N_5333);
or U14495 (N_14495,N_8558,N_3379);
xor U14496 (N_14496,N_5180,N_2130);
xnor U14497 (N_14497,N_3272,N_8915);
or U14498 (N_14498,N_5019,N_8275);
or U14499 (N_14499,N_5872,N_5188);
and U14500 (N_14500,N_487,N_9761);
xor U14501 (N_14501,N_2474,N_103);
nand U14502 (N_14502,N_8242,N_515);
nand U14503 (N_14503,N_9267,N_3928);
xor U14504 (N_14504,N_9163,N_2989);
or U14505 (N_14505,N_9729,N_5026);
nand U14506 (N_14506,N_5774,N_941);
xor U14507 (N_14507,N_1733,N_3230);
or U14508 (N_14508,N_2511,N_3960);
nor U14509 (N_14509,N_5325,N_2419);
and U14510 (N_14510,N_1346,N_5376);
or U14511 (N_14511,N_8121,N_3548);
nand U14512 (N_14512,N_5283,N_4858);
or U14513 (N_14513,N_3167,N_5018);
nor U14514 (N_14514,N_5055,N_5852);
nand U14515 (N_14515,N_3976,N_4578);
nor U14516 (N_14516,N_9960,N_621);
nor U14517 (N_14517,N_1084,N_816);
nand U14518 (N_14518,N_9808,N_8021);
or U14519 (N_14519,N_6183,N_5260);
or U14520 (N_14520,N_160,N_5067);
or U14521 (N_14521,N_7015,N_9669);
or U14522 (N_14522,N_5695,N_2302);
nor U14523 (N_14523,N_7487,N_7547);
nor U14524 (N_14524,N_9206,N_7679);
and U14525 (N_14525,N_2107,N_5046);
and U14526 (N_14526,N_5321,N_8279);
and U14527 (N_14527,N_7252,N_6879);
and U14528 (N_14528,N_3235,N_5346);
or U14529 (N_14529,N_6122,N_5181);
or U14530 (N_14530,N_2255,N_7792);
xnor U14531 (N_14531,N_5630,N_4559);
nand U14532 (N_14532,N_6483,N_1595);
or U14533 (N_14533,N_8099,N_4896);
nor U14534 (N_14534,N_3691,N_206);
nor U14535 (N_14535,N_6251,N_1563);
xor U14536 (N_14536,N_2714,N_1219);
nand U14537 (N_14537,N_8943,N_7961);
xor U14538 (N_14538,N_6719,N_1100);
and U14539 (N_14539,N_7146,N_7694);
or U14540 (N_14540,N_2568,N_4742);
nand U14541 (N_14541,N_1369,N_2895);
and U14542 (N_14542,N_4980,N_81);
and U14543 (N_14543,N_4238,N_9475);
nand U14544 (N_14544,N_3796,N_497);
nand U14545 (N_14545,N_4710,N_4400);
or U14546 (N_14546,N_6525,N_5518);
xnor U14547 (N_14547,N_9736,N_8348);
nand U14548 (N_14548,N_1754,N_2435);
and U14549 (N_14549,N_9031,N_9051);
nand U14550 (N_14550,N_5755,N_2982);
xnor U14551 (N_14551,N_7634,N_4716);
nor U14552 (N_14552,N_4444,N_5850);
nor U14553 (N_14553,N_6090,N_5438);
nand U14554 (N_14554,N_2844,N_1045);
nor U14555 (N_14555,N_7949,N_8929);
or U14556 (N_14556,N_953,N_2307);
and U14557 (N_14557,N_9446,N_1556);
or U14558 (N_14558,N_517,N_4622);
nand U14559 (N_14559,N_1877,N_9364);
nor U14560 (N_14560,N_3676,N_3947);
nor U14561 (N_14561,N_5814,N_1769);
xnor U14562 (N_14562,N_6145,N_9403);
nor U14563 (N_14563,N_2721,N_5052);
nor U14564 (N_14564,N_586,N_4289);
or U14565 (N_14565,N_6160,N_2777);
nor U14566 (N_14566,N_7681,N_7852);
nor U14567 (N_14567,N_352,N_3678);
and U14568 (N_14568,N_2276,N_8423);
nor U14569 (N_14569,N_3294,N_5819);
and U14570 (N_14570,N_916,N_6005);
and U14571 (N_14571,N_4528,N_4880);
or U14572 (N_14572,N_793,N_2648);
and U14573 (N_14573,N_1810,N_9501);
and U14574 (N_14574,N_2925,N_5323);
nand U14575 (N_14575,N_2179,N_6015);
xor U14576 (N_14576,N_5966,N_978);
nand U14577 (N_14577,N_7499,N_4179);
or U14578 (N_14578,N_3210,N_9200);
and U14579 (N_14579,N_3030,N_7419);
and U14580 (N_14580,N_9128,N_4186);
xor U14581 (N_14581,N_1663,N_597);
nor U14582 (N_14582,N_5174,N_1985);
nor U14583 (N_14583,N_1637,N_8231);
xor U14584 (N_14584,N_976,N_2106);
nor U14585 (N_14585,N_6986,N_6417);
nor U14586 (N_14586,N_5490,N_8171);
or U14587 (N_14587,N_1947,N_5610);
xor U14588 (N_14588,N_3414,N_7898);
or U14589 (N_14589,N_6320,N_184);
xor U14590 (N_14590,N_5566,N_8011);
nor U14591 (N_14591,N_7570,N_149);
nor U14592 (N_14592,N_8830,N_4103);
nor U14593 (N_14593,N_6432,N_5498);
nor U14594 (N_14594,N_2986,N_7833);
nor U14595 (N_14595,N_2711,N_4888);
nor U14596 (N_14596,N_4322,N_9329);
nand U14597 (N_14597,N_9993,N_7823);
and U14598 (N_14598,N_963,N_6372);
xor U14599 (N_14599,N_9604,N_5390);
nand U14600 (N_14600,N_1501,N_722);
xnor U14601 (N_14601,N_7897,N_8428);
nor U14602 (N_14602,N_6582,N_3619);
xor U14603 (N_14603,N_6949,N_3835);
or U14604 (N_14604,N_8232,N_6374);
xor U14605 (N_14605,N_3576,N_6332);
nand U14606 (N_14606,N_1852,N_6063);
and U14607 (N_14607,N_8925,N_8161);
nand U14608 (N_14608,N_3061,N_8421);
nor U14609 (N_14609,N_6535,N_2602);
xnor U14610 (N_14610,N_5971,N_3432);
nor U14611 (N_14611,N_8604,N_8075);
xor U14612 (N_14612,N_5108,N_2445);
nor U14613 (N_14613,N_7390,N_5997);
nor U14614 (N_14614,N_4513,N_9698);
xor U14615 (N_14615,N_989,N_3268);
nand U14616 (N_14616,N_4726,N_6538);
xnor U14617 (N_14617,N_7160,N_2375);
nand U14618 (N_14618,N_1905,N_2400);
nand U14619 (N_14619,N_6852,N_7133);
xor U14620 (N_14620,N_6248,N_1266);
nand U14621 (N_14621,N_7796,N_6864);
nand U14622 (N_14622,N_7767,N_9462);
and U14623 (N_14623,N_491,N_917);
and U14624 (N_14624,N_4882,N_1960);
and U14625 (N_14625,N_2295,N_1057);
nor U14626 (N_14626,N_8881,N_5263);
or U14627 (N_14627,N_8571,N_8424);
xnor U14628 (N_14628,N_6542,N_5877);
and U14629 (N_14629,N_8827,N_2828);
or U14630 (N_14630,N_9217,N_6985);
nor U14631 (N_14631,N_4949,N_7711);
xor U14632 (N_14632,N_8134,N_3355);
xor U14633 (N_14633,N_1945,N_2899);
and U14634 (N_14634,N_4287,N_6618);
nor U14635 (N_14635,N_9494,N_1834);
xnor U14636 (N_14636,N_9717,N_3228);
and U14637 (N_14637,N_5729,N_8006);
nor U14638 (N_14638,N_787,N_7624);
and U14639 (N_14639,N_7854,N_9678);
and U14640 (N_14640,N_1394,N_289);
nand U14641 (N_14641,N_887,N_7091);
and U14642 (N_14642,N_3901,N_8441);
nand U14643 (N_14643,N_574,N_6264);
or U14644 (N_14644,N_4978,N_3582);
nor U14645 (N_14645,N_7488,N_9718);
or U14646 (N_14646,N_9140,N_6324);
and U14647 (N_14647,N_4619,N_3877);
nand U14648 (N_14648,N_6603,N_2405);
nor U14649 (N_14649,N_1224,N_1287);
and U14650 (N_14650,N_8997,N_4164);
xor U14651 (N_14651,N_9448,N_584);
nor U14652 (N_14652,N_2421,N_4931);
or U14653 (N_14653,N_1487,N_6147);
or U14654 (N_14654,N_2452,N_3382);
nor U14655 (N_14655,N_5329,N_702);
nor U14656 (N_14656,N_3206,N_1242);
and U14657 (N_14657,N_9794,N_3339);
or U14658 (N_14658,N_1456,N_1151);
nand U14659 (N_14659,N_5680,N_2791);
nand U14660 (N_14660,N_6061,N_3747);
nor U14661 (N_14661,N_2335,N_1798);
and U14662 (N_14662,N_4007,N_7942);
nor U14663 (N_14663,N_2271,N_7625);
or U14664 (N_14664,N_9654,N_3777);
and U14665 (N_14665,N_415,N_9391);
or U14666 (N_14666,N_7121,N_7101);
or U14667 (N_14667,N_91,N_5740);
or U14668 (N_14668,N_2775,N_5093);
nand U14669 (N_14669,N_6888,N_8998);
and U14670 (N_14670,N_6649,N_869);
or U14671 (N_14671,N_3149,N_6661);
or U14672 (N_14672,N_9345,N_3776);
and U14673 (N_14673,N_6367,N_3253);
nand U14674 (N_14674,N_7467,N_2987);
xor U14675 (N_14675,N_3633,N_8300);
nor U14676 (N_14676,N_7773,N_2870);
or U14677 (N_14677,N_1904,N_6913);
and U14678 (N_14678,N_3493,N_2299);
or U14679 (N_14679,N_8686,N_670);
nor U14680 (N_14680,N_1528,N_6104);
nand U14681 (N_14681,N_5129,N_6766);
or U14682 (N_14682,N_755,N_202);
or U14683 (N_14683,N_326,N_7880);
xnor U14684 (N_14684,N_9658,N_1767);
xnor U14685 (N_14685,N_8481,N_8653);
and U14686 (N_14686,N_5314,N_2118);
nor U14687 (N_14687,N_2096,N_8266);
and U14688 (N_14688,N_6082,N_1644);
nor U14689 (N_14689,N_8531,N_8725);
or U14690 (N_14690,N_6247,N_9197);
or U14691 (N_14691,N_5640,N_4436);
and U14692 (N_14692,N_4703,N_9209);
and U14693 (N_14693,N_6070,N_7541);
nand U14694 (N_14694,N_1145,N_819);
and U14695 (N_14695,N_5759,N_5839);
and U14696 (N_14696,N_2656,N_5999);
and U14697 (N_14697,N_6287,N_79);
nand U14698 (N_14698,N_6220,N_4502);
and U14699 (N_14699,N_6079,N_5184);
or U14700 (N_14700,N_1139,N_173);
or U14701 (N_14701,N_6025,N_7300);
and U14702 (N_14702,N_4367,N_4571);
xnor U14703 (N_14703,N_9847,N_5687);
and U14704 (N_14704,N_6814,N_6602);
nand U14705 (N_14705,N_3483,N_1743);
and U14706 (N_14706,N_4884,N_2341);
nand U14707 (N_14707,N_3337,N_683);
nor U14708 (N_14708,N_1176,N_7987);
nor U14709 (N_14709,N_16,N_4887);
or U14710 (N_14710,N_2650,N_5939);
xor U14711 (N_14711,N_6461,N_4611);
nor U14712 (N_14712,N_5924,N_9147);
nand U14713 (N_14713,N_2104,N_6859);
nor U14714 (N_14714,N_709,N_5531);
nand U14715 (N_14715,N_5208,N_7835);
and U14716 (N_14716,N_2587,N_7939);
xor U14717 (N_14717,N_4260,N_6824);
xnor U14718 (N_14718,N_9220,N_4394);
nor U14719 (N_14719,N_5294,N_9368);
and U14720 (N_14720,N_4846,N_6653);
xor U14721 (N_14721,N_558,N_9239);
xnor U14722 (N_14722,N_3618,N_4808);
and U14723 (N_14723,N_5060,N_3174);
and U14724 (N_14724,N_1774,N_7435);
or U14725 (N_14725,N_3666,N_5269);
and U14726 (N_14726,N_2821,N_882);
and U14727 (N_14727,N_9449,N_7072);
xnor U14728 (N_14728,N_1678,N_3593);
and U14729 (N_14729,N_6844,N_4547);
or U14730 (N_14730,N_8046,N_5114);
xor U14731 (N_14731,N_9424,N_6405);
and U14732 (N_14732,N_3635,N_766);
xnor U14733 (N_14733,N_3169,N_233);
or U14734 (N_14734,N_1806,N_428);
nand U14735 (N_14735,N_7249,N_4764);
xor U14736 (N_14736,N_5139,N_5225);
xor U14737 (N_14737,N_8495,N_7255);
or U14738 (N_14738,N_3730,N_9550);
xor U14739 (N_14739,N_7347,N_959);
nand U14740 (N_14740,N_3361,N_1124);
or U14741 (N_14741,N_5391,N_90);
nor U14742 (N_14742,N_8854,N_3539);
or U14743 (N_14743,N_2203,N_1927);
nor U14744 (N_14744,N_1350,N_2398);
and U14745 (N_14745,N_9656,N_9286);
xor U14746 (N_14746,N_6705,N_6191);
nand U14747 (N_14747,N_1963,N_6265);
xnor U14748 (N_14748,N_1197,N_739);
nand U14749 (N_14749,N_4474,N_3335);
nor U14750 (N_14750,N_7619,N_1359);
xnor U14751 (N_14751,N_5514,N_8076);
and U14752 (N_14752,N_5681,N_3016);
nand U14753 (N_14753,N_3383,N_8605);
xor U14754 (N_14754,N_2464,N_1939);
or U14755 (N_14755,N_7753,N_4642);
nor U14756 (N_14756,N_4364,N_1907);
xnor U14757 (N_14757,N_9378,N_9265);
nor U14758 (N_14758,N_9353,N_8718);
and U14759 (N_14759,N_5481,N_1893);
nor U14760 (N_14760,N_7536,N_4677);
or U14761 (N_14761,N_2740,N_8432);
nor U14762 (N_14762,N_9315,N_9688);
nor U14763 (N_14763,N_9049,N_5958);
or U14764 (N_14764,N_7326,N_1821);
nor U14765 (N_14765,N_9758,N_732);
xnor U14766 (N_14766,N_2094,N_5823);
nand U14767 (N_14767,N_2373,N_1917);
xor U14768 (N_14768,N_6281,N_8977);
or U14769 (N_14769,N_8273,N_2046);
xor U14770 (N_14770,N_3307,N_6914);
or U14771 (N_14771,N_4793,N_2074);
and U14772 (N_14772,N_3130,N_8058);
or U14773 (N_14773,N_8661,N_6843);
and U14774 (N_14774,N_1254,N_6738);
nor U14775 (N_14775,N_1411,N_3732);
and U14776 (N_14776,N_9432,N_7293);
or U14777 (N_14777,N_298,N_2902);
or U14778 (N_14778,N_8381,N_2910);
nand U14779 (N_14779,N_1400,N_6917);
nand U14780 (N_14780,N_1041,N_3690);
xor U14781 (N_14781,N_51,N_2890);
or U14782 (N_14782,N_8706,N_1444);
xor U14783 (N_14783,N_4686,N_3213);
xor U14784 (N_14784,N_7258,N_5494);
and U14785 (N_14785,N_6818,N_4132);
or U14786 (N_14786,N_8316,N_6464);
nor U14787 (N_14787,N_234,N_9419);
nor U14788 (N_14788,N_8385,N_1461);
xnor U14789 (N_14789,N_174,N_5598);
and U14790 (N_14790,N_634,N_6797);
nor U14791 (N_14791,N_6023,N_8675);
or U14792 (N_14792,N_7875,N_6149);
and U14793 (N_14793,N_7977,N_2031);
nor U14794 (N_14794,N_4826,N_2461);
and U14795 (N_14795,N_7421,N_8676);
xor U14796 (N_14796,N_3531,N_2065);
nor U14797 (N_14797,N_8340,N_6227);
or U14798 (N_14798,N_1693,N_5593);
and U14799 (N_14799,N_1003,N_2804);
and U14800 (N_14800,N_6533,N_2629);
nand U14801 (N_14801,N_5721,N_3843);
nor U14802 (N_14802,N_4727,N_7250);
nand U14803 (N_14803,N_4974,N_9105);
xor U14804 (N_14804,N_6243,N_6094);
nor U14805 (N_14805,N_492,N_1469);
and U14806 (N_14806,N_5468,N_3536);
xnor U14807 (N_14807,N_9627,N_2499);
or U14808 (N_14808,N_5935,N_5172);
xnor U14809 (N_14809,N_3731,N_6909);
nand U14810 (N_14810,N_1186,N_2145);
nor U14811 (N_14811,N_2973,N_6389);
nor U14812 (N_14812,N_2210,N_6296);
nand U14813 (N_14813,N_4636,N_5008);
or U14814 (N_14814,N_86,N_2751);
nor U14815 (N_14815,N_6187,N_5278);
or U14816 (N_14816,N_2496,N_7128);
xnor U14817 (N_14817,N_5519,N_6877);
and U14818 (N_14818,N_6727,N_6403);
nand U14819 (N_14819,N_2968,N_5625);
nor U14820 (N_14820,N_5902,N_5705);
nand U14821 (N_14821,N_4927,N_493);
nor U14822 (N_14822,N_4794,N_3217);
and U14823 (N_14823,N_6702,N_8188);
nor U14824 (N_14824,N_1299,N_8583);
nand U14825 (N_14825,N_143,N_9663);
and U14826 (N_14826,N_5645,N_1179);
or U14827 (N_14827,N_7787,N_9655);
and U14828 (N_14828,N_4106,N_370);
or U14829 (N_14829,N_494,N_7094);
and U14830 (N_14830,N_5107,N_3607);
and U14831 (N_14831,N_1561,N_6558);
and U14832 (N_14832,N_7130,N_8069);
nand U14833 (N_14833,N_7508,N_4714);
and U14834 (N_14834,N_4651,N_4806);
and U14835 (N_14835,N_189,N_4631);
xnor U14836 (N_14836,N_4902,N_3148);
nor U14837 (N_14837,N_7642,N_4245);
xnor U14838 (N_14838,N_3484,N_8301);
xnor U14839 (N_14839,N_4643,N_4159);
xnor U14840 (N_14840,N_1034,N_8391);
nor U14841 (N_14841,N_5750,N_1026);
nand U14842 (N_14842,N_9636,N_6515);
nand U14843 (N_14843,N_5919,N_4679);
xor U14844 (N_14844,N_9069,N_5145);
and U14845 (N_14845,N_7353,N_471);
nor U14846 (N_14846,N_1822,N_8056);
and U14847 (N_14847,N_4803,N_2109);
and U14848 (N_14848,N_4967,N_4074);
xor U14849 (N_14849,N_4705,N_5964);
or U14850 (N_14850,N_6771,N_5583);
nand U14851 (N_14851,N_7113,N_4959);
or U14852 (N_14852,N_8477,N_7519);
nor U14853 (N_14853,N_312,N_4331);
xor U14854 (N_14854,N_7650,N_706);
xor U14855 (N_14855,N_506,N_4471);
xnor U14856 (N_14856,N_6580,N_8257);
nor U14857 (N_14857,N_919,N_740);
nor U14858 (N_14858,N_7278,N_8736);
nand U14859 (N_14859,N_3807,N_7214);
and U14860 (N_14860,N_4853,N_4609);
nand U14861 (N_14861,N_6120,N_7572);
nand U14862 (N_14862,N_7628,N_409);
nor U14863 (N_14863,N_8656,N_6710);
xor U14864 (N_14864,N_9437,N_7116);
and U14865 (N_14865,N_5068,N_7591);
xnor U14866 (N_14866,N_9473,N_1512);
xor U14867 (N_14867,N_5686,N_7043);
and U14868 (N_14868,N_4344,N_3000);
or U14869 (N_14869,N_5639,N_4512);
nand U14870 (N_14870,N_9609,N_3139);
and U14871 (N_14871,N_8036,N_7936);
nor U14872 (N_14872,N_9116,N_3755);
nand U14873 (N_14873,N_6134,N_2674);
xnor U14874 (N_14874,N_4385,N_4296);
and U14875 (N_14875,N_459,N_2766);
nor U14876 (N_14876,N_4301,N_3501);
xor U14877 (N_14877,N_7737,N_7251);
or U14878 (N_14878,N_1584,N_7934);
nand U14879 (N_14879,N_3667,N_3771);
nand U14880 (N_14880,N_3056,N_55);
and U14881 (N_14881,N_7393,N_846);
nand U14882 (N_14882,N_4925,N_3265);
nand U14883 (N_14883,N_1001,N_2281);
xnor U14884 (N_14884,N_4907,N_4599);
or U14885 (N_14885,N_1434,N_4724);
nor U14886 (N_14886,N_3930,N_8203);
and U14887 (N_14887,N_9142,N_2169);
and U14888 (N_14888,N_3651,N_8190);
or U14889 (N_14889,N_1701,N_8790);
and U14890 (N_14890,N_8489,N_151);
nand U14891 (N_14891,N_4242,N_6532);
or U14892 (N_14892,N_7306,N_9650);
or U14893 (N_14893,N_3917,N_4731);
nor U14894 (N_14894,N_9359,N_8589);
xor U14895 (N_14895,N_7981,N_3969);
nor U14896 (N_14896,N_6897,N_4587);
or U14897 (N_14897,N_8826,N_5661);
xor U14898 (N_14898,N_5994,N_31);
xor U14899 (N_14899,N_1813,N_4202);
nand U14900 (N_14900,N_2661,N_8501);
and U14901 (N_14901,N_8068,N_8325);
or U14902 (N_14902,N_9626,N_9567);
xnor U14903 (N_14903,N_4183,N_5655);
or U14904 (N_14904,N_1245,N_8700);
nor U14905 (N_14905,N_6377,N_6607);
or U14906 (N_14906,N_2288,N_3714);
nand U14907 (N_14907,N_6801,N_2719);
nand U14908 (N_14908,N_7786,N_2834);
nor U14909 (N_14909,N_3101,N_3094);
nor U14910 (N_14910,N_8269,N_2061);
and U14911 (N_14911,N_8444,N_243);
nor U14912 (N_14912,N_7035,N_4433);
xnor U14913 (N_14913,N_9821,N_3407);
nor U14914 (N_14914,N_228,N_6011);
xnor U14915 (N_14915,N_9334,N_4969);
and U14916 (N_14916,N_0,N_7097);
nand U14917 (N_14917,N_9327,N_845);
or U14918 (N_14918,N_6659,N_4533);
nor U14919 (N_14919,N_8936,N_1935);
or U14920 (N_14920,N_5904,N_4701);
or U14921 (N_14921,N_3390,N_2015);
xnor U14922 (N_14922,N_3832,N_8417);
nand U14923 (N_14923,N_2735,N_4275);
or U14924 (N_14924,N_1173,N_4673);
nor U14925 (N_14925,N_230,N_5156);
nand U14926 (N_14926,N_5138,N_2156);
xor U14927 (N_14927,N_8118,N_2525);
nor U14928 (N_14928,N_301,N_3504);
nor U14929 (N_14929,N_2113,N_6132);
or U14930 (N_14930,N_7462,N_5458);
and U14931 (N_14931,N_1059,N_9482);
or U14932 (N_14932,N_4648,N_2974);
xnor U14933 (N_14933,N_7791,N_1751);
xnor U14934 (N_14934,N_6662,N_645);
and U14935 (N_14935,N_2695,N_3581);
nor U14936 (N_14936,N_2940,N_1734);
and U14937 (N_14937,N_1321,N_4728);
nand U14938 (N_14938,N_9122,N_7343);
xor U14939 (N_14939,N_1515,N_2554);
or U14940 (N_14940,N_6979,N_6420);
nor U14941 (N_14941,N_5211,N_7006);
xnor U14942 (N_14942,N_3498,N_157);
and U14943 (N_14943,N_6091,N_5445);
nor U14944 (N_14944,N_2926,N_2245);
nor U14945 (N_14945,N_8959,N_931);
or U14946 (N_14946,N_836,N_4816);
and U14947 (N_14947,N_4427,N_9619);
nand U14948 (N_14948,N_600,N_3275);
and U14949 (N_14949,N_7587,N_4610);
nor U14950 (N_14950,N_1211,N_105);
and U14951 (N_14951,N_562,N_8196);
nand U14952 (N_14952,N_5591,N_367);
and U14953 (N_14953,N_4964,N_4567);
xnor U14954 (N_14954,N_4483,N_1078);
xnor U14955 (N_14955,N_5040,N_3507);
and U14956 (N_14956,N_5791,N_4017);
nor U14957 (N_14957,N_9123,N_6636);
nor U14958 (N_14958,N_8342,N_42);
xor U14959 (N_14959,N_8770,N_7843);
xor U14960 (N_14960,N_5256,N_4982);
nor U14961 (N_14961,N_3402,N_5693);
and U14962 (N_14962,N_2580,N_5549);
nand U14963 (N_14963,N_7361,N_2978);
nand U14964 (N_14964,N_5166,N_903);
nor U14965 (N_14965,N_3535,N_435);
or U14966 (N_14966,N_7575,N_6555);
nand U14967 (N_14967,N_5668,N_2010);
or U14968 (N_14968,N_2970,N_393);
nand U14969 (N_14969,N_9850,N_1090);
xnor U14970 (N_14970,N_9492,N_9750);
and U14971 (N_14971,N_8086,N_2475);
xnor U14972 (N_14972,N_8756,N_6993);
nor U14973 (N_14973,N_5806,N_2224);
nor U14974 (N_14974,N_3060,N_5513);
xnor U14975 (N_14975,N_7644,N_9291);
xnor U14976 (N_14976,N_9186,N_7417);
xnor U14977 (N_14977,N_478,N_9096);
or U14978 (N_14978,N_6717,N_1448);
xor U14979 (N_14979,N_9276,N_4141);
and U14980 (N_14980,N_263,N_8766);
nand U14981 (N_14981,N_9372,N_7952);
nor U14982 (N_14982,N_8170,N_3797);
and U14983 (N_14983,N_4704,N_6453);
and U14984 (N_14984,N_3233,N_5692);
or U14985 (N_14985,N_9426,N_6954);
or U14986 (N_14986,N_4786,N_8662);
nand U14987 (N_14987,N_2433,N_9479);
nor U14988 (N_14988,N_4072,N_2051);
and U14989 (N_14989,N_8705,N_4257);
nand U14990 (N_14990,N_410,N_8387);
nor U14991 (N_14991,N_1247,N_1601);
and U14992 (N_14992,N_1921,N_2960);
and U14993 (N_14993,N_5104,N_4537);
nor U14994 (N_14994,N_3445,N_6999);
xnor U14995 (N_14995,N_7722,N_8730);
or U14996 (N_14996,N_5050,N_4491);
nand U14997 (N_14997,N_8912,N_7051);
and U14998 (N_14998,N_1095,N_1558);
nand U14999 (N_14999,N_749,N_9259);
and U15000 (N_15000,N_9511,N_932);
xnor U15001 (N_15001,N_7216,N_8336);
and U15002 (N_15002,N_3934,N_5274);
nand U15003 (N_15003,N_682,N_8431);
and U15004 (N_15004,N_1079,N_6340);
and U15005 (N_15005,N_5992,N_9843);
or U15006 (N_15006,N_8160,N_9485);
nand U15007 (N_15007,N_7984,N_9370);
nor U15008 (N_15008,N_1902,N_2139);
or U15009 (N_15009,N_4669,N_74);
xor U15010 (N_15010,N_1191,N_2409);
or U15011 (N_15011,N_8905,N_4430);
xor U15012 (N_15012,N_8903,N_3882);
or U15013 (N_15013,N_8278,N_2488);
xnor U15014 (N_15014,N_7549,N_1506);
xnor U15015 (N_15015,N_6946,N_7108);
or U15016 (N_15016,N_9627,N_2537);
nand U15017 (N_15017,N_1468,N_5505);
xor U15018 (N_15018,N_5968,N_1997);
xor U15019 (N_15019,N_8986,N_5690);
nand U15020 (N_15020,N_9929,N_3944);
nor U15021 (N_15021,N_1420,N_9281);
nor U15022 (N_15022,N_3582,N_536);
nor U15023 (N_15023,N_4441,N_384);
xor U15024 (N_15024,N_2952,N_5711);
and U15025 (N_15025,N_7432,N_2171);
nand U15026 (N_15026,N_3884,N_5595);
and U15027 (N_15027,N_5775,N_1438);
nand U15028 (N_15028,N_6679,N_7965);
nor U15029 (N_15029,N_8311,N_1409);
nor U15030 (N_15030,N_7612,N_9417);
and U15031 (N_15031,N_848,N_6626);
and U15032 (N_15032,N_6269,N_2988);
nor U15033 (N_15033,N_776,N_8107);
nor U15034 (N_15034,N_8907,N_3755);
nand U15035 (N_15035,N_349,N_5005);
nor U15036 (N_15036,N_7783,N_6378);
xor U15037 (N_15037,N_757,N_4294);
and U15038 (N_15038,N_3932,N_1775);
nand U15039 (N_15039,N_7486,N_7702);
or U15040 (N_15040,N_8449,N_8999);
nor U15041 (N_15041,N_2454,N_8869);
nor U15042 (N_15042,N_9468,N_36);
xnor U15043 (N_15043,N_2849,N_1766);
xnor U15044 (N_15044,N_4494,N_3032);
or U15045 (N_15045,N_7864,N_9009);
xnor U15046 (N_15046,N_9941,N_826);
and U15047 (N_15047,N_3624,N_3564);
xor U15048 (N_15048,N_1233,N_2189);
xor U15049 (N_15049,N_6045,N_2404);
xnor U15050 (N_15050,N_6582,N_4001);
or U15051 (N_15051,N_5422,N_7800);
nor U15052 (N_15052,N_4040,N_7945);
xnor U15053 (N_15053,N_8683,N_2461);
xor U15054 (N_15054,N_8494,N_3981);
and U15055 (N_15055,N_5719,N_1651);
xor U15056 (N_15056,N_8232,N_4173);
xor U15057 (N_15057,N_7131,N_2405);
nand U15058 (N_15058,N_7209,N_266);
xnor U15059 (N_15059,N_3109,N_6409);
nor U15060 (N_15060,N_8139,N_5061);
xor U15061 (N_15061,N_6071,N_5752);
xor U15062 (N_15062,N_5841,N_1013);
or U15063 (N_15063,N_817,N_3955);
or U15064 (N_15064,N_9063,N_3367);
nand U15065 (N_15065,N_5078,N_3949);
xnor U15066 (N_15066,N_1901,N_8844);
xor U15067 (N_15067,N_7811,N_1024);
nor U15068 (N_15068,N_5243,N_6157);
or U15069 (N_15069,N_2828,N_1223);
xor U15070 (N_15070,N_6584,N_5171);
xor U15071 (N_15071,N_5752,N_8434);
nand U15072 (N_15072,N_9238,N_2931);
and U15073 (N_15073,N_8172,N_4827);
nor U15074 (N_15074,N_604,N_7577);
and U15075 (N_15075,N_356,N_6536);
or U15076 (N_15076,N_5199,N_6537);
or U15077 (N_15077,N_6332,N_9274);
or U15078 (N_15078,N_3222,N_2051);
and U15079 (N_15079,N_9489,N_8019);
and U15080 (N_15080,N_8528,N_8335);
and U15081 (N_15081,N_9987,N_1450);
or U15082 (N_15082,N_6296,N_1582);
nand U15083 (N_15083,N_5936,N_4844);
nor U15084 (N_15084,N_468,N_572);
or U15085 (N_15085,N_3079,N_1079);
nor U15086 (N_15086,N_4757,N_4706);
nor U15087 (N_15087,N_1989,N_1276);
xnor U15088 (N_15088,N_2370,N_5234);
or U15089 (N_15089,N_6130,N_9686);
nand U15090 (N_15090,N_2256,N_4052);
and U15091 (N_15091,N_7332,N_2471);
or U15092 (N_15092,N_5666,N_2440);
and U15093 (N_15093,N_7856,N_2037);
or U15094 (N_15094,N_3106,N_1502);
nand U15095 (N_15095,N_9899,N_8395);
and U15096 (N_15096,N_3179,N_858);
xnor U15097 (N_15097,N_2311,N_1056);
and U15098 (N_15098,N_4059,N_872);
nor U15099 (N_15099,N_6212,N_7876);
nor U15100 (N_15100,N_936,N_1943);
or U15101 (N_15101,N_3622,N_1248);
nand U15102 (N_15102,N_3082,N_2687);
xor U15103 (N_15103,N_9964,N_3445);
nand U15104 (N_15104,N_6174,N_9543);
xor U15105 (N_15105,N_6963,N_6334);
or U15106 (N_15106,N_4578,N_2303);
nor U15107 (N_15107,N_8067,N_9158);
and U15108 (N_15108,N_9154,N_707);
nand U15109 (N_15109,N_1050,N_9354);
nor U15110 (N_15110,N_3698,N_2793);
nand U15111 (N_15111,N_142,N_3856);
nand U15112 (N_15112,N_9153,N_6329);
nor U15113 (N_15113,N_5072,N_2184);
nor U15114 (N_15114,N_7518,N_3775);
xnor U15115 (N_15115,N_4425,N_8524);
nand U15116 (N_15116,N_5092,N_859);
nand U15117 (N_15117,N_7564,N_3564);
xnor U15118 (N_15118,N_8644,N_7210);
nand U15119 (N_15119,N_8986,N_4934);
and U15120 (N_15120,N_9192,N_7244);
xor U15121 (N_15121,N_4299,N_1714);
and U15122 (N_15122,N_2934,N_2851);
or U15123 (N_15123,N_3143,N_6480);
xor U15124 (N_15124,N_3174,N_8750);
nand U15125 (N_15125,N_9429,N_8919);
xor U15126 (N_15126,N_5338,N_7252);
nor U15127 (N_15127,N_5563,N_1020);
or U15128 (N_15128,N_9764,N_507);
or U15129 (N_15129,N_8502,N_5073);
nand U15130 (N_15130,N_5168,N_4220);
xnor U15131 (N_15131,N_8894,N_1561);
xor U15132 (N_15132,N_9383,N_4789);
and U15133 (N_15133,N_4751,N_633);
nor U15134 (N_15134,N_4524,N_2604);
or U15135 (N_15135,N_7846,N_4945);
nor U15136 (N_15136,N_1948,N_1559);
or U15137 (N_15137,N_3771,N_9287);
or U15138 (N_15138,N_6346,N_7912);
or U15139 (N_15139,N_5020,N_8837);
nand U15140 (N_15140,N_1079,N_5208);
nand U15141 (N_15141,N_1365,N_8599);
nand U15142 (N_15142,N_5224,N_4804);
xnor U15143 (N_15143,N_5066,N_9964);
or U15144 (N_15144,N_794,N_7124);
xor U15145 (N_15145,N_709,N_2503);
or U15146 (N_15146,N_942,N_7059);
or U15147 (N_15147,N_565,N_9163);
nor U15148 (N_15148,N_3669,N_9719);
xor U15149 (N_15149,N_6412,N_6838);
nor U15150 (N_15150,N_2169,N_455);
and U15151 (N_15151,N_3325,N_8699);
and U15152 (N_15152,N_5490,N_4567);
and U15153 (N_15153,N_3768,N_8577);
or U15154 (N_15154,N_6872,N_3794);
or U15155 (N_15155,N_2998,N_9035);
and U15156 (N_15156,N_7544,N_9241);
xor U15157 (N_15157,N_3853,N_7073);
nor U15158 (N_15158,N_8195,N_804);
nor U15159 (N_15159,N_1822,N_5187);
nand U15160 (N_15160,N_6490,N_7867);
nand U15161 (N_15161,N_7475,N_2670);
and U15162 (N_15162,N_8457,N_9790);
and U15163 (N_15163,N_245,N_6317);
nor U15164 (N_15164,N_9747,N_9498);
and U15165 (N_15165,N_6099,N_3216);
or U15166 (N_15166,N_5732,N_196);
or U15167 (N_15167,N_3904,N_8458);
and U15168 (N_15168,N_9016,N_594);
or U15169 (N_15169,N_5694,N_3990);
nand U15170 (N_15170,N_9748,N_8756);
and U15171 (N_15171,N_7646,N_5970);
xor U15172 (N_15172,N_3859,N_7901);
nand U15173 (N_15173,N_2250,N_4164);
nor U15174 (N_15174,N_7017,N_3299);
nor U15175 (N_15175,N_8387,N_7465);
xnor U15176 (N_15176,N_4233,N_6493);
nand U15177 (N_15177,N_1590,N_1745);
nor U15178 (N_15178,N_2606,N_9547);
nor U15179 (N_15179,N_9263,N_8472);
or U15180 (N_15180,N_6615,N_338);
nand U15181 (N_15181,N_3512,N_1993);
nand U15182 (N_15182,N_2176,N_1109);
nor U15183 (N_15183,N_4507,N_8958);
or U15184 (N_15184,N_8975,N_3434);
xor U15185 (N_15185,N_5353,N_4);
nand U15186 (N_15186,N_7866,N_373);
xor U15187 (N_15187,N_2170,N_3694);
xnor U15188 (N_15188,N_1219,N_6513);
nor U15189 (N_15189,N_2111,N_9592);
xnor U15190 (N_15190,N_8714,N_8722);
or U15191 (N_15191,N_330,N_7801);
nand U15192 (N_15192,N_9846,N_5992);
and U15193 (N_15193,N_7668,N_6922);
nor U15194 (N_15194,N_8856,N_1029);
and U15195 (N_15195,N_512,N_17);
and U15196 (N_15196,N_1198,N_6991);
or U15197 (N_15197,N_4202,N_3374);
nand U15198 (N_15198,N_9574,N_1334);
xnor U15199 (N_15199,N_1815,N_3416);
nor U15200 (N_15200,N_9056,N_9356);
xor U15201 (N_15201,N_2040,N_4935);
xnor U15202 (N_15202,N_7674,N_9405);
and U15203 (N_15203,N_8806,N_1151);
nand U15204 (N_15204,N_6393,N_9497);
nor U15205 (N_15205,N_8669,N_2458);
and U15206 (N_15206,N_9965,N_8580);
nand U15207 (N_15207,N_5829,N_5112);
xor U15208 (N_15208,N_430,N_5403);
and U15209 (N_15209,N_971,N_8370);
xor U15210 (N_15210,N_323,N_5057);
xor U15211 (N_15211,N_361,N_7322);
or U15212 (N_15212,N_4421,N_6974);
xor U15213 (N_15213,N_2233,N_5947);
or U15214 (N_15214,N_5098,N_3856);
xor U15215 (N_15215,N_3677,N_3185);
and U15216 (N_15216,N_9642,N_4866);
or U15217 (N_15217,N_8791,N_5917);
nor U15218 (N_15218,N_3603,N_8482);
nor U15219 (N_15219,N_3075,N_1307);
nand U15220 (N_15220,N_1650,N_7013);
and U15221 (N_15221,N_3293,N_8552);
and U15222 (N_15222,N_5308,N_3161);
nor U15223 (N_15223,N_7938,N_8689);
nor U15224 (N_15224,N_2149,N_3263);
nand U15225 (N_15225,N_5993,N_7758);
and U15226 (N_15226,N_8638,N_2015);
and U15227 (N_15227,N_2712,N_2522);
nor U15228 (N_15228,N_2693,N_1380);
xor U15229 (N_15229,N_682,N_939);
xor U15230 (N_15230,N_8169,N_4210);
or U15231 (N_15231,N_4250,N_2479);
nand U15232 (N_15232,N_8983,N_2448);
nor U15233 (N_15233,N_1478,N_4060);
and U15234 (N_15234,N_8534,N_4327);
xnor U15235 (N_15235,N_3013,N_5956);
nor U15236 (N_15236,N_4622,N_1263);
and U15237 (N_15237,N_160,N_588);
nand U15238 (N_15238,N_1964,N_9300);
or U15239 (N_15239,N_2116,N_2541);
nand U15240 (N_15240,N_3350,N_9656);
or U15241 (N_15241,N_8759,N_6691);
and U15242 (N_15242,N_3388,N_1257);
or U15243 (N_15243,N_9227,N_3598);
and U15244 (N_15244,N_9988,N_7407);
and U15245 (N_15245,N_9030,N_3959);
or U15246 (N_15246,N_5567,N_3718);
or U15247 (N_15247,N_5515,N_861);
or U15248 (N_15248,N_8349,N_6592);
or U15249 (N_15249,N_7386,N_5099);
or U15250 (N_15250,N_7774,N_8536);
xor U15251 (N_15251,N_1666,N_8949);
nor U15252 (N_15252,N_1037,N_4897);
and U15253 (N_15253,N_5505,N_3357);
nor U15254 (N_15254,N_3722,N_5638);
or U15255 (N_15255,N_546,N_401);
nor U15256 (N_15256,N_2975,N_3567);
or U15257 (N_15257,N_3034,N_6157);
nor U15258 (N_15258,N_6389,N_7468);
nand U15259 (N_15259,N_5364,N_2681);
or U15260 (N_15260,N_185,N_6009);
nand U15261 (N_15261,N_8081,N_8017);
nor U15262 (N_15262,N_9623,N_8367);
nor U15263 (N_15263,N_4835,N_1105);
nor U15264 (N_15264,N_5494,N_4232);
nor U15265 (N_15265,N_3470,N_2137);
xor U15266 (N_15266,N_9341,N_4676);
or U15267 (N_15267,N_7894,N_3562);
nand U15268 (N_15268,N_7927,N_1260);
and U15269 (N_15269,N_6792,N_5694);
xnor U15270 (N_15270,N_9808,N_3788);
and U15271 (N_15271,N_9836,N_8993);
nand U15272 (N_15272,N_3907,N_3767);
nand U15273 (N_15273,N_2963,N_2119);
nand U15274 (N_15274,N_7621,N_1774);
nand U15275 (N_15275,N_2610,N_5453);
and U15276 (N_15276,N_5959,N_5566);
nand U15277 (N_15277,N_5478,N_2746);
nor U15278 (N_15278,N_9814,N_8355);
or U15279 (N_15279,N_3125,N_8769);
nand U15280 (N_15280,N_8453,N_6309);
nor U15281 (N_15281,N_8170,N_2971);
nor U15282 (N_15282,N_9662,N_7059);
and U15283 (N_15283,N_9722,N_9876);
nor U15284 (N_15284,N_2984,N_6884);
or U15285 (N_15285,N_3388,N_1896);
or U15286 (N_15286,N_4647,N_3264);
nor U15287 (N_15287,N_5528,N_290);
xor U15288 (N_15288,N_5172,N_3137);
nand U15289 (N_15289,N_5926,N_7796);
nor U15290 (N_15290,N_1161,N_4046);
nand U15291 (N_15291,N_1012,N_837);
or U15292 (N_15292,N_3074,N_6677);
and U15293 (N_15293,N_6170,N_6311);
or U15294 (N_15294,N_9581,N_236);
nand U15295 (N_15295,N_3643,N_9846);
nor U15296 (N_15296,N_9337,N_4895);
nand U15297 (N_15297,N_4458,N_2962);
xor U15298 (N_15298,N_2062,N_7332);
and U15299 (N_15299,N_1330,N_8840);
or U15300 (N_15300,N_8692,N_8700);
nor U15301 (N_15301,N_5274,N_3848);
and U15302 (N_15302,N_1293,N_3637);
xnor U15303 (N_15303,N_2621,N_8458);
and U15304 (N_15304,N_245,N_632);
and U15305 (N_15305,N_4109,N_6831);
nor U15306 (N_15306,N_7429,N_7687);
and U15307 (N_15307,N_6631,N_1843);
nor U15308 (N_15308,N_5177,N_8093);
nor U15309 (N_15309,N_1345,N_5373);
or U15310 (N_15310,N_4670,N_7479);
nand U15311 (N_15311,N_1587,N_1485);
or U15312 (N_15312,N_5541,N_3870);
nor U15313 (N_15313,N_6356,N_3583);
or U15314 (N_15314,N_5987,N_4341);
nand U15315 (N_15315,N_909,N_8856);
xor U15316 (N_15316,N_4633,N_1026);
nand U15317 (N_15317,N_4283,N_6392);
xnor U15318 (N_15318,N_8396,N_1653);
nand U15319 (N_15319,N_4511,N_2167);
or U15320 (N_15320,N_5934,N_9324);
xor U15321 (N_15321,N_1078,N_1694);
nand U15322 (N_15322,N_3658,N_9597);
xor U15323 (N_15323,N_5146,N_5816);
or U15324 (N_15324,N_2997,N_2480);
and U15325 (N_15325,N_9481,N_9329);
nor U15326 (N_15326,N_5141,N_6271);
and U15327 (N_15327,N_3847,N_2088);
xor U15328 (N_15328,N_7629,N_9744);
or U15329 (N_15329,N_5346,N_6715);
or U15330 (N_15330,N_6745,N_3256);
nand U15331 (N_15331,N_599,N_279);
or U15332 (N_15332,N_307,N_3894);
xnor U15333 (N_15333,N_8945,N_9512);
or U15334 (N_15334,N_3291,N_7164);
or U15335 (N_15335,N_6128,N_6683);
nor U15336 (N_15336,N_3616,N_6350);
nand U15337 (N_15337,N_4863,N_6995);
and U15338 (N_15338,N_4885,N_7938);
and U15339 (N_15339,N_4335,N_3916);
nor U15340 (N_15340,N_755,N_4734);
nand U15341 (N_15341,N_7734,N_7067);
xor U15342 (N_15342,N_6950,N_2824);
nor U15343 (N_15343,N_1780,N_7421);
nand U15344 (N_15344,N_8950,N_2123);
xnor U15345 (N_15345,N_8896,N_8370);
nand U15346 (N_15346,N_4180,N_6887);
nor U15347 (N_15347,N_9884,N_2179);
nand U15348 (N_15348,N_7558,N_7956);
nor U15349 (N_15349,N_7660,N_8844);
nor U15350 (N_15350,N_3813,N_4270);
and U15351 (N_15351,N_946,N_604);
and U15352 (N_15352,N_479,N_9347);
xor U15353 (N_15353,N_3165,N_5135);
and U15354 (N_15354,N_4389,N_7472);
xnor U15355 (N_15355,N_340,N_4673);
or U15356 (N_15356,N_1932,N_7002);
nor U15357 (N_15357,N_3656,N_7587);
or U15358 (N_15358,N_9829,N_7622);
nor U15359 (N_15359,N_1577,N_2718);
and U15360 (N_15360,N_3092,N_3213);
nand U15361 (N_15361,N_1094,N_3312);
nor U15362 (N_15362,N_4124,N_7706);
nor U15363 (N_15363,N_4034,N_3013);
nor U15364 (N_15364,N_1856,N_5204);
nor U15365 (N_15365,N_3296,N_8018);
xor U15366 (N_15366,N_5009,N_2270);
or U15367 (N_15367,N_2,N_8847);
xnor U15368 (N_15368,N_1703,N_2394);
and U15369 (N_15369,N_2215,N_1111);
nor U15370 (N_15370,N_9462,N_3437);
and U15371 (N_15371,N_7772,N_5429);
nand U15372 (N_15372,N_2023,N_8316);
nor U15373 (N_15373,N_7967,N_14);
nand U15374 (N_15374,N_8771,N_3682);
or U15375 (N_15375,N_5744,N_835);
and U15376 (N_15376,N_4520,N_518);
xnor U15377 (N_15377,N_6102,N_3676);
xnor U15378 (N_15378,N_3402,N_254);
xnor U15379 (N_15379,N_7271,N_6582);
xnor U15380 (N_15380,N_1246,N_2889);
xor U15381 (N_15381,N_3544,N_8709);
nor U15382 (N_15382,N_893,N_9031);
nand U15383 (N_15383,N_2318,N_9825);
xor U15384 (N_15384,N_7739,N_3760);
xnor U15385 (N_15385,N_31,N_8310);
and U15386 (N_15386,N_4868,N_1193);
or U15387 (N_15387,N_943,N_5538);
xnor U15388 (N_15388,N_7671,N_3474);
or U15389 (N_15389,N_6729,N_6361);
nor U15390 (N_15390,N_9238,N_5278);
or U15391 (N_15391,N_679,N_1824);
nor U15392 (N_15392,N_9560,N_5853);
or U15393 (N_15393,N_7455,N_5521);
or U15394 (N_15394,N_5953,N_876);
xnor U15395 (N_15395,N_4072,N_1110);
and U15396 (N_15396,N_8537,N_9141);
xnor U15397 (N_15397,N_4095,N_8495);
or U15398 (N_15398,N_1369,N_4473);
nor U15399 (N_15399,N_3726,N_9789);
and U15400 (N_15400,N_355,N_7791);
and U15401 (N_15401,N_5392,N_847);
or U15402 (N_15402,N_2531,N_6203);
xor U15403 (N_15403,N_1077,N_2721);
and U15404 (N_15404,N_5217,N_353);
nand U15405 (N_15405,N_218,N_6968);
xor U15406 (N_15406,N_8106,N_9316);
nand U15407 (N_15407,N_5831,N_3854);
nand U15408 (N_15408,N_5842,N_5884);
and U15409 (N_15409,N_309,N_3375);
and U15410 (N_15410,N_2164,N_9799);
nand U15411 (N_15411,N_9468,N_273);
or U15412 (N_15412,N_7631,N_533);
nor U15413 (N_15413,N_683,N_4017);
xnor U15414 (N_15414,N_585,N_8111);
xor U15415 (N_15415,N_7884,N_5986);
or U15416 (N_15416,N_1758,N_2191);
or U15417 (N_15417,N_9630,N_1667);
xor U15418 (N_15418,N_9380,N_2666);
and U15419 (N_15419,N_4349,N_6139);
nand U15420 (N_15420,N_5603,N_582);
nor U15421 (N_15421,N_1856,N_2435);
xor U15422 (N_15422,N_4375,N_1742);
or U15423 (N_15423,N_8269,N_9433);
and U15424 (N_15424,N_6613,N_1341);
xor U15425 (N_15425,N_7590,N_1979);
and U15426 (N_15426,N_704,N_944);
and U15427 (N_15427,N_1368,N_652);
and U15428 (N_15428,N_9743,N_6514);
nor U15429 (N_15429,N_1409,N_4608);
nor U15430 (N_15430,N_7859,N_2065);
nor U15431 (N_15431,N_5917,N_5874);
and U15432 (N_15432,N_9422,N_291);
nor U15433 (N_15433,N_4377,N_6525);
xor U15434 (N_15434,N_5709,N_1776);
xor U15435 (N_15435,N_4542,N_7212);
nand U15436 (N_15436,N_7612,N_705);
and U15437 (N_15437,N_4008,N_9349);
nor U15438 (N_15438,N_8258,N_901);
nor U15439 (N_15439,N_6170,N_2628);
or U15440 (N_15440,N_3523,N_454);
nor U15441 (N_15441,N_5867,N_7901);
or U15442 (N_15442,N_9879,N_2281);
xor U15443 (N_15443,N_3799,N_6174);
nor U15444 (N_15444,N_6945,N_3196);
and U15445 (N_15445,N_4934,N_3129);
or U15446 (N_15446,N_6127,N_3041);
nor U15447 (N_15447,N_8269,N_6075);
nor U15448 (N_15448,N_8871,N_1441);
nor U15449 (N_15449,N_7197,N_681);
or U15450 (N_15450,N_4722,N_2485);
and U15451 (N_15451,N_45,N_6569);
and U15452 (N_15452,N_7381,N_7363);
and U15453 (N_15453,N_6954,N_5214);
nor U15454 (N_15454,N_8702,N_2468);
or U15455 (N_15455,N_5800,N_2071);
nor U15456 (N_15456,N_5510,N_7455);
or U15457 (N_15457,N_4140,N_5033);
and U15458 (N_15458,N_4797,N_8414);
nand U15459 (N_15459,N_2365,N_6754);
and U15460 (N_15460,N_8252,N_4595);
and U15461 (N_15461,N_4732,N_7727);
and U15462 (N_15462,N_8773,N_6965);
xnor U15463 (N_15463,N_7953,N_5709);
xnor U15464 (N_15464,N_5431,N_5673);
xnor U15465 (N_15465,N_4394,N_3414);
nand U15466 (N_15466,N_6880,N_3995);
xor U15467 (N_15467,N_826,N_8430);
and U15468 (N_15468,N_5803,N_1778);
and U15469 (N_15469,N_5306,N_9017);
xnor U15470 (N_15470,N_7831,N_1744);
or U15471 (N_15471,N_7203,N_708);
xor U15472 (N_15472,N_8806,N_3913);
or U15473 (N_15473,N_4416,N_7344);
nor U15474 (N_15474,N_7147,N_1794);
and U15475 (N_15475,N_5008,N_8358);
nand U15476 (N_15476,N_1518,N_9695);
nor U15477 (N_15477,N_788,N_3186);
or U15478 (N_15478,N_7146,N_9772);
and U15479 (N_15479,N_2829,N_2317);
and U15480 (N_15480,N_1107,N_6727);
xor U15481 (N_15481,N_5078,N_4864);
or U15482 (N_15482,N_9197,N_2544);
and U15483 (N_15483,N_9643,N_5204);
or U15484 (N_15484,N_8914,N_4992);
xor U15485 (N_15485,N_4844,N_7350);
and U15486 (N_15486,N_8849,N_8823);
or U15487 (N_15487,N_4531,N_4961);
or U15488 (N_15488,N_1968,N_8664);
and U15489 (N_15489,N_8044,N_6749);
or U15490 (N_15490,N_7144,N_8);
nor U15491 (N_15491,N_1644,N_2173);
or U15492 (N_15492,N_4415,N_4102);
nand U15493 (N_15493,N_1668,N_4405);
and U15494 (N_15494,N_1815,N_2310);
xnor U15495 (N_15495,N_4703,N_8625);
xor U15496 (N_15496,N_6237,N_4291);
and U15497 (N_15497,N_5358,N_8486);
nand U15498 (N_15498,N_6751,N_1870);
and U15499 (N_15499,N_4261,N_1015);
or U15500 (N_15500,N_1358,N_3630);
nand U15501 (N_15501,N_1572,N_6407);
nand U15502 (N_15502,N_5423,N_1065);
xor U15503 (N_15503,N_5391,N_2285);
nand U15504 (N_15504,N_987,N_3489);
xor U15505 (N_15505,N_2852,N_2776);
and U15506 (N_15506,N_8964,N_7943);
xnor U15507 (N_15507,N_7051,N_3943);
xor U15508 (N_15508,N_5736,N_1929);
or U15509 (N_15509,N_6855,N_5273);
xnor U15510 (N_15510,N_7890,N_1516);
and U15511 (N_15511,N_6200,N_4972);
xor U15512 (N_15512,N_9160,N_9173);
xnor U15513 (N_15513,N_4830,N_9010);
nor U15514 (N_15514,N_6594,N_8785);
nor U15515 (N_15515,N_6472,N_4470);
and U15516 (N_15516,N_3813,N_9635);
nor U15517 (N_15517,N_4845,N_3134);
nor U15518 (N_15518,N_8977,N_239);
xor U15519 (N_15519,N_1279,N_66);
xnor U15520 (N_15520,N_4253,N_1887);
and U15521 (N_15521,N_3022,N_4441);
nand U15522 (N_15522,N_6393,N_6372);
nand U15523 (N_15523,N_1473,N_3048);
and U15524 (N_15524,N_9254,N_6501);
nor U15525 (N_15525,N_226,N_65);
or U15526 (N_15526,N_4354,N_3113);
and U15527 (N_15527,N_5460,N_4802);
and U15528 (N_15528,N_6746,N_968);
nand U15529 (N_15529,N_9253,N_8556);
and U15530 (N_15530,N_3660,N_7778);
or U15531 (N_15531,N_8083,N_8555);
or U15532 (N_15532,N_3430,N_8346);
nor U15533 (N_15533,N_6503,N_118);
nor U15534 (N_15534,N_1099,N_9723);
or U15535 (N_15535,N_4914,N_4037);
nor U15536 (N_15536,N_3349,N_6278);
or U15537 (N_15537,N_3352,N_8652);
xor U15538 (N_15538,N_3178,N_6434);
and U15539 (N_15539,N_9749,N_9959);
nand U15540 (N_15540,N_9108,N_259);
nor U15541 (N_15541,N_7939,N_3087);
nor U15542 (N_15542,N_5770,N_6732);
or U15543 (N_15543,N_500,N_5262);
nand U15544 (N_15544,N_6700,N_3834);
xnor U15545 (N_15545,N_5717,N_9102);
and U15546 (N_15546,N_7386,N_2780);
or U15547 (N_15547,N_1712,N_5843);
nor U15548 (N_15548,N_7252,N_1319);
xnor U15549 (N_15549,N_8322,N_4263);
or U15550 (N_15550,N_2631,N_7264);
or U15551 (N_15551,N_2090,N_3510);
xnor U15552 (N_15552,N_9187,N_3279);
or U15553 (N_15553,N_6997,N_8085);
nand U15554 (N_15554,N_605,N_331);
nand U15555 (N_15555,N_8088,N_5733);
or U15556 (N_15556,N_2404,N_5687);
and U15557 (N_15557,N_8457,N_5153);
xnor U15558 (N_15558,N_2866,N_5753);
and U15559 (N_15559,N_4406,N_3091);
and U15560 (N_15560,N_2212,N_3180);
or U15561 (N_15561,N_9026,N_6528);
nand U15562 (N_15562,N_7526,N_835);
or U15563 (N_15563,N_35,N_4388);
or U15564 (N_15564,N_8342,N_5636);
nor U15565 (N_15565,N_5865,N_835);
nor U15566 (N_15566,N_7964,N_5434);
and U15567 (N_15567,N_5563,N_9092);
xnor U15568 (N_15568,N_9173,N_3385);
nand U15569 (N_15569,N_3088,N_1564);
nor U15570 (N_15570,N_9795,N_5843);
nor U15571 (N_15571,N_7068,N_6915);
and U15572 (N_15572,N_7735,N_1961);
xnor U15573 (N_15573,N_9332,N_4583);
nand U15574 (N_15574,N_6634,N_3503);
xnor U15575 (N_15575,N_8644,N_8393);
xor U15576 (N_15576,N_2370,N_6795);
and U15577 (N_15577,N_7661,N_1548);
xor U15578 (N_15578,N_2836,N_3015);
nor U15579 (N_15579,N_6804,N_8568);
nor U15580 (N_15580,N_595,N_1851);
nor U15581 (N_15581,N_8905,N_1528);
nand U15582 (N_15582,N_5820,N_68);
nor U15583 (N_15583,N_446,N_2905);
nand U15584 (N_15584,N_9716,N_4717);
nor U15585 (N_15585,N_1011,N_2720);
nand U15586 (N_15586,N_9249,N_7033);
nor U15587 (N_15587,N_1331,N_7655);
or U15588 (N_15588,N_8240,N_4632);
or U15589 (N_15589,N_8763,N_8189);
nor U15590 (N_15590,N_6849,N_5499);
and U15591 (N_15591,N_6029,N_4854);
xor U15592 (N_15592,N_8675,N_9869);
or U15593 (N_15593,N_2431,N_1433);
xor U15594 (N_15594,N_1094,N_5717);
xor U15595 (N_15595,N_1772,N_8681);
or U15596 (N_15596,N_4854,N_9070);
or U15597 (N_15597,N_3456,N_8355);
nand U15598 (N_15598,N_3748,N_7595);
and U15599 (N_15599,N_7208,N_656);
nor U15600 (N_15600,N_6048,N_3557);
or U15601 (N_15601,N_1532,N_1722);
and U15602 (N_15602,N_126,N_3885);
and U15603 (N_15603,N_4283,N_1279);
or U15604 (N_15604,N_4719,N_5855);
and U15605 (N_15605,N_8615,N_2403);
nand U15606 (N_15606,N_1976,N_1359);
xnor U15607 (N_15607,N_6724,N_2214);
nand U15608 (N_15608,N_5675,N_9385);
nor U15609 (N_15609,N_5702,N_5339);
and U15610 (N_15610,N_6167,N_1067);
nor U15611 (N_15611,N_1208,N_5870);
nor U15612 (N_15612,N_416,N_5759);
and U15613 (N_15613,N_2347,N_8058);
xnor U15614 (N_15614,N_456,N_8200);
or U15615 (N_15615,N_4335,N_6377);
and U15616 (N_15616,N_8177,N_4867);
xor U15617 (N_15617,N_8684,N_1495);
nand U15618 (N_15618,N_8429,N_1650);
or U15619 (N_15619,N_2836,N_6912);
or U15620 (N_15620,N_6200,N_7014);
xnor U15621 (N_15621,N_7441,N_782);
or U15622 (N_15622,N_5621,N_3369);
and U15623 (N_15623,N_4283,N_7465);
nand U15624 (N_15624,N_8291,N_2800);
xor U15625 (N_15625,N_2929,N_6453);
xor U15626 (N_15626,N_8148,N_154);
nor U15627 (N_15627,N_4461,N_197);
or U15628 (N_15628,N_1135,N_6137);
and U15629 (N_15629,N_8854,N_2636);
or U15630 (N_15630,N_8202,N_5108);
nand U15631 (N_15631,N_4426,N_6598);
or U15632 (N_15632,N_9706,N_2608);
xor U15633 (N_15633,N_7799,N_3038);
nand U15634 (N_15634,N_1506,N_4561);
nor U15635 (N_15635,N_2620,N_5266);
and U15636 (N_15636,N_9509,N_2917);
xnor U15637 (N_15637,N_2815,N_430);
and U15638 (N_15638,N_9948,N_3483);
nand U15639 (N_15639,N_6683,N_975);
and U15640 (N_15640,N_3688,N_6966);
nor U15641 (N_15641,N_3499,N_4575);
nand U15642 (N_15642,N_6025,N_6071);
xor U15643 (N_15643,N_1967,N_7836);
xnor U15644 (N_15644,N_5886,N_671);
nor U15645 (N_15645,N_8356,N_6361);
or U15646 (N_15646,N_2723,N_6847);
or U15647 (N_15647,N_380,N_3357);
nand U15648 (N_15648,N_743,N_276);
nand U15649 (N_15649,N_4095,N_3289);
nor U15650 (N_15650,N_444,N_6954);
xor U15651 (N_15651,N_9019,N_7923);
xor U15652 (N_15652,N_205,N_7826);
xor U15653 (N_15653,N_4326,N_5713);
and U15654 (N_15654,N_9423,N_3108);
xor U15655 (N_15655,N_9730,N_3569);
nor U15656 (N_15656,N_8483,N_3842);
nand U15657 (N_15657,N_8463,N_1160);
and U15658 (N_15658,N_977,N_5369);
nor U15659 (N_15659,N_3307,N_9105);
or U15660 (N_15660,N_3126,N_7751);
xor U15661 (N_15661,N_8301,N_6299);
and U15662 (N_15662,N_2950,N_9026);
nor U15663 (N_15663,N_391,N_6759);
and U15664 (N_15664,N_8313,N_4391);
xor U15665 (N_15665,N_4424,N_2553);
xor U15666 (N_15666,N_6874,N_5518);
nor U15667 (N_15667,N_6143,N_2833);
nand U15668 (N_15668,N_6366,N_5543);
and U15669 (N_15669,N_7444,N_2782);
or U15670 (N_15670,N_1173,N_5133);
and U15671 (N_15671,N_6495,N_5701);
and U15672 (N_15672,N_7899,N_9914);
nor U15673 (N_15673,N_8176,N_969);
xor U15674 (N_15674,N_9429,N_6265);
and U15675 (N_15675,N_3132,N_615);
and U15676 (N_15676,N_8011,N_4724);
and U15677 (N_15677,N_1153,N_3568);
xnor U15678 (N_15678,N_2252,N_5689);
or U15679 (N_15679,N_2664,N_2540);
or U15680 (N_15680,N_3807,N_9323);
xnor U15681 (N_15681,N_6492,N_9083);
xnor U15682 (N_15682,N_9812,N_2425);
nand U15683 (N_15683,N_5524,N_5908);
xor U15684 (N_15684,N_329,N_5514);
xor U15685 (N_15685,N_4319,N_7718);
or U15686 (N_15686,N_1578,N_2487);
nor U15687 (N_15687,N_5469,N_9361);
and U15688 (N_15688,N_7854,N_376);
xor U15689 (N_15689,N_2212,N_4174);
and U15690 (N_15690,N_772,N_5422);
and U15691 (N_15691,N_3779,N_8795);
xor U15692 (N_15692,N_3567,N_6887);
xor U15693 (N_15693,N_221,N_3899);
nand U15694 (N_15694,N_5206,N_7749);
nor U15695 (N_15695,N_2066,N_5202);
nor U15696 (N_15696,N_8068,N_9473);
nand U15697 (N_15697,N_6367,N_6743);
nor U15698 (N_15698,N_3182,N_6443);
nand U15699 (N_15699,N_7608,N_9127);
nor U15700 (N_15700,N_4074,N_6309);
xnor U15701 (N_15701,N_7623,N_6766);
or U15702 (N_15702,N_48,N_3468);
nor U15703 (N_15703,N_596,N_1704);
or U15704 (N_15704,N_5213,N_8840);
or U15705 (N_15705,N_185,N_5446);
or U15706 (N_15706,N_7508,N_8525);
nand U15707 (N_15707,N_1517,N_2422);
xnor U15708 (N_15708,N_7798,N_8023);
and U15709 (N_15709,N_1029,N_8296);
and U15710 (N_15710,N_8773,N_6733);
nand U15711 (N_15711,N_7575,N_5694);
or U15712 (N_15712,N_4563,N_145);
nand U15713 (N_15713,N_678,N_9070);
nand U15714 (N_15714,N_688,N_3706);
nor U15715 (N_15715,N_9508,N_1855);
xor U15716 (N_15716,N_3987,N_7509);
or U15717 (N_15717,N_7242,N_689);
nor U15718 (N_15718,N_4741,N_7336);
nor U15719 (N_15719,N_1271,N_4352);
xor U15720 (N_15720,N_3429,N_9340);
nor U15721 (N_15721,N_5271,N_9563);
or U15722 (N_15722,N_4694,N_4945);
nand U15723 (N_15723,N_9460,N_5939);
or U15724 (N_15724,N_2740,N_9010);
nor U15725 (N_15725,N_342,N_2757);
nand U15726 (N_15726,N_331,N_8622);
nor U15727 (N_15727,N_4096,N_1522);
nor U15728 (N_15728,N_2330,N_2708);
nor U15729 (N_15729,N_5697,N_7149);
nand U15730 (N_15730,N_9880,N_1512);
xor U15731 (N_15731,N_1471,N_5575);
xnor U15732 (N_15732,N_4711,N_107);
and U15733 (N_15733,N_7768,N_1352);
nor U15734 (N_15734,N_4189,N_4347);
xnor U15735 (N_15735,N_7940,N_2072);
or U15736 (N_15736,N_2737,N_1008);
and U15737 (N_15737,N_7257,N_1269);
nor U15738 (N_15738,N_8000,N_7057);
nor U15739 (N_15739,N_9341,N_2215);
and U15740 (N_15740,N_8254,N_3190);
nand U15741 (N_15741,N_6232,N_8611);
and U15742 (N_15742,N_5337,N_3093);
xor U15743 (N_15743,N_5071,N_866);
and U15744 (N_15744,N_2253,N_5912);
nand U15745 (N_15745,N_7474,N_8135);
nor U15746 (N_15746,N_581,N_6931);
nand U15747 (N_15747,N_3099,N_5652);
nor U15748 (N_15748,N_249,N_3591);
nor U15749 (N_15749,N_5554,N_4826);
and U15750 (N_15750,N_4113,N_7761);
or U15751 (N_15751,N_6899,N_6858);
nor U15752 (N_15752,N_9642,N_6315);
xor U15753 (N_15753,N_2642,N_1220);
or U15754 (N_15754,N_3543,N_3551);
nand U15755 (N_15755,N_915,N_1295);
or U15756 (N_15756,N_2228,N_1403);
xor U15757 (N_15757,N_4586,N_6577);
nor U15758 (N_15758,N_7973,N_7609);
nand U15759 (N_15759,N_4441,N_9596);
and U15760 (N_15760,N_8795,N_7525);
and U15761 (N_15761,N_1423,N_4361);
and U15762 (N_15762,N_3975,N_3898);
and U15763 (N_15763,N_3001,N_383);
or U15764 (N_15764,N_891,N_6071);
xnor U15765 (N_15765,N_8627,N_9299);
or U15766 (N_15766,N_7213,N_6759);
xnor U15767 (N_15767,N_5169,N_5060);
and U15768 (N_15768,N_2812,N_9712);
xnor U15769 (N_15769,N_3317,N_2662);
and U15770 (N_15770,N_4636,N_4674);
and U15771 (N_15771,N_2000,N_9573);
or U15772 (N_15772,N_9465,N_3633);
nand U15773 (N_15773,N_8001,N_3116);
nor U15774 (N_15774,N_1212,N_6934);
nand U15775 (N_15775,N_2578,N_7950);
nor U15776 (N_15776,N_6975,N_7961);
nor U15777 (N_15777,N_5390,N_6668);
and U15778 (N_15778,N_9967,N_4914);
or U15779 (N_15779,N_998,N_9450);
or U15780 (N_15780,N_360,N_2237);
nand U15781 (N_15781,N_9038,N_8373);
nand U15782 (N_15782,N_1872,N_9943);
and U15783 (N_15783,N_1246,N_5515);
nor U15784 (N_15784,N_7246,N_3462);
nor U15785 (N_15785,N_1200,N_6395);
or U15786 (N_15786,N_7545,N_198);
nand U15787 (N_15787,N_314,N_6177);
and U15788 (N_15788,N_9721,N_1301);
nand U15789 (N_15789,N_6483,N_3211);
nor U15790 (N_15790,N_2961,N_5586);
or U15791 (N_15791,N_6768,N_519);
and U15792 (N_15792,N_4412,N_5605);
and U15793 (N_15793,N_2427,N_1412);
and U15794 (N_15794,N_1481,N_326);
xor U15795 (N_15795,N_7345,N_9865);
nor U15796 (N_15796,N_3508,N_8945);
or U15797 (N_15797,N_1322,N_5400);
xnor U15798 (N_15798,N_9871,N_2246);
or U15799 (N_15799,N_5565,N_405);
and U15800 (N_15800,N_3427,N_657);
and U15801 (N_15801,N_9624,N_8708);
nor U15802 (N_15802,N_4519,N_7111);
nand U15803 (N_15803,N_6050,N_244);
nor U15804 (N_15804,N_7592,N_4478);
nand U15805 (N_15805,N_5606,N_3217);
nand U15806 (N_15806,N_2882,N_1797);
or U15807 (N_15807,N_9371,N_3887);
xnor U15808 (N_15808,N_4443,N_2946);
nor U15809 (N_15809,N_2873,N_7895);
nor U15810 (N_15810,N_1797,N_4896);
nand U15811 (N_15811,N_8383,N_3724);
nand U15812 (N_15812,N_7033,N_7552);
xnor U15813 (N_15813,N_7459,N_2497);
or U15814 (N_15814,N_534,N_3847);
nor U15815 (N_15815,N_572,N_3953);
nor U15816 (N_15816,N_1908,N_7929);
xor U15817 (N_15817,N_5322,N_7303);
nor U15818 (N_15818,N_5943,N_245);
nor U15819 (N_15819,N_5163,N_730);
xnor U15820 (N_15820,N_5292,N_546);
nor U15821 (N_15821,N_9292,N_5461);
xor U15822 (N_15822,N_8109,N_3744);
and U15823 (N_15823,N_1574,N_6266);
nand U15824 (N_15824,N_1045,N_6156);
xnor U15825 (N_15825,N_3085,N_8744);
xor U15826 (N_15826,N_128,N_7121);
or U15827 (N_15827,N_1032,N_5652);
xnor U15828 (N_15828,N_5724,N_3221);
and U15829 (N_15829,N_7582,N_2036);
nor U15830 (N_15830,N_4718,N_3214);
or U15831 (N_15831,N_5229,N_9853);
nor U15832 (N_15832,N_748,N_4071);
nand U15833 (N_15833,N_5589,N_8161);
nand U15834 (N_15834,N_6166,N_3770);
or U15835 (N_15835,N_6772,N_2506);
xor U15836 (N_15836,N_3837,N_5905);
and U15837 (N_15837,N_4583,N_3851);
nand U15838 (N_15838,N_6934,N_4746);
nor U15839 (N_15839,N_6445,N_5901);
nand U15840 (N_15840,N_6736,N_2337);
or U15841 (N_15841,N_6972,N_5677);
nor U15842 (N_15842,N_5337,N_1282);
nand U15843 (N_15843,N_3800,N_3661);
nand U15844 (N_15844,N_6694,N_2461);
nand U15845 (N_15845,N_5185,N_6600);
nor U15846 (N_15846,N_346,N_6793);
xnor U15847 (N_15847,N_8215,N_2598);
or U15848 (N_15848,N_5288,N_2132);
xor U15849 (N_15849,N_5298,N_6273);
or U15850 (N_15850,N_4788,N_2534);
nand U15851 (N_15851,N_7247,N_8699);
and U15852 (N_15852,N_8887,N_4623);
nand U15853 (N_15853,N_3640,N_6590);
nand U15854 (N_15854,N_2104,N_4232);
and U15855 (N_15855,N_8693,N_5283);
xor U15856 (N_15856,N_3516,N_5480);
or U15857 (N_15857,N_2772,N_1635);
nand U15858 (N_15858,N_9397,N_6464);
xor U15859 (N_15859,N_7089,N_6948);
or U15860 (N_15860,N_3916,N_5816);
nor U15861 (N_15861,N_1328,N_9247);
xor U15862 (N_15862,N_7060,N_5788);
or U15863 (N_15863,N_1458,N_1613);
or U15864 (N_15864,N_6043,N_7676);
and U15865 (N_15865,N_1025,N_2542);
or U15866 (N_15866,N_2589,N_6310);
nand U15867 (N_15867,N_1684,N_7272);
nand U15868 (N_15868,N_5922,N_7694);
nand U15869 (N_15869,N_3591,N_5170);
nor U15870 (N_15870,N_2977,N_8406);
or U15871 (N_15871,N_9549,N_4670);
or U15872 (N_15872,N_8868,N_2224);
nor U15873 (N_15873,N_8831,N_6591);
nor U15874 (N_15874,N_626,N_843);
or U15875 (N_15875,N_5846,N_3689);
or U15876 (N_15876,N_6495,N_448);
nor U15877 (N_15877,N_767,N_9214);
nand U15878 (N_15878,N_9559,N_9353);
nand U15879 (N_15879,N_81,N_6935);
and U15880 (N_15880,N_271,N_4437);
nand U15881 (N_15881,N_3595,N_5961);
nor U15882 (N_15882,N_3542,N_1749);
nor U15883 (N_15883,N_7102,N_6948);
nand U15884 (N_15884,N_8697,N_2943);
or U15885 (N_15885,N_4950,N_7697);
or U15886 (N_15886,N_6832,N_6639);
xor U15887 (N_15887,N_3373,N_5434);
xnor U15888 (N_15888,N_9244,N_6034);
or U15889 (N_15889,N_9024,N_9731);
xnor U15890 (N_15890,N_2681,N_792);
or U15891 (N_15891,N_6809,N_8004);
or U15892 (N_15892,N_5276,N_5118);
nor U15893 (N_15893,N_3275,N_8433);
or U15894 (N_15894,N_8556,N_1859);
xnor U15895 (N_15895,N_2906,N_6922);
and U15896 (N_15896,N_4665,N_7709);
or U15897 (N_15897,N_5132,N_5026);
nand U15898 (N_15898,N_7274,N_571);
nor U15899 (N_15899,N_4417,N_5408);
or U15900 (N_15900,N_4837,N_7208);
nor U15901 (N_15901,N_2911,N_6953);
or U15902 (N_15902,N_8778,N_883);
or U15903 (N_15903,N_8835,N_1521);
nand U15904 (N_15904,N_8911,N_2948);
nand U15905 (N_15905,N_9704,N_2956);
and U15906 (N_15906,N_8727,N_578);
nor U15907 (N_15907,N_3051,N_7974);
xnor U15908 (N_15908,N_8682,N_6311);
and U15909 (N_15909,N_8237,N_6808);
nor U15910 (N_15910,N_8164,N_5444);
and U15911 (N_15911,N_4289,N_3563);
xor U15912 (N_15912,N_642,N_6913);
nand U15913 (N_15913,N_4825,N_877);
nor U15914 (N_15914,N_2825,N_9312);
or U15915 (N_15915,N_6968,N_3234);
and U15916 (N_15916,N_2879,N_7373);
xnor U15917 (N_15917,N_9920,N_3558);
and U15918 (N_15918,N_9288,N_5555);
nor U15919 (N_15919,N_4188,N_8432);
and U15920 (N_15920,N_2840,N_5591);
nand U15921 (N_15921,N_7367,N_9578);
and U15922 (N_15922,N_6964,N_9586);
nor U15923 (N_15923,N_5704,N_1036);
xnor U15924 (N_15924,N_603,N_4081);
xnor U15925 (N_15925,N_7565,N_1237);
nand U15926 (N_15926,N_9050,N_7285);
nor U15927 (N_15927,N_8134,N_2653);
nand U15928 (N_15928,N_3362,N_5586);
xnor U15929 (N_15929,N_7440,N_3207);
or U15930 (N_15930,N_1455,N_5421);
and U15931 (N_15931,N_2848,N_522);
xnor U15932 (N_15932,N_5848,N_8868);
nand U15933 (N_15933,N_4608,N_1190);
or U15934 (N_15934,N_9944,N_8931);
xor U15935 (N_15935,N_7354,N_7808);
xor U15936 (N_15936,N_6403,N_9878);
or U15937 (N_15937,N_7659,N_8496);
xor U15938 (N_15938,N_9339,N_395);
nand U15939 (N_15939,N_379,N_5583);
xnor U15940 (N_15940,N_8972,N_9660);
and U15941 (N_15941,N_8430,N_604);
xnor U15942 (N_15942,N_8087,N_6266);
or U15943 (N_15943,N_6952,N_9768);
xnor U15944 (N_15944,N_9071,N_8896);
nor U15945 (N_15945,N_365,N_7394);
or U15946 (N_15946,N_8153,N_8305);
or U15947 (N_15947,N_754,N_9971);
nand U15948 (N_15948,N_984,N_5281);
xor U15949 (N_15949,N_7968,N_8908);
nor U15950 (N_15950,N_4714,N_2700);
or U15951 (N_15951,N_2394,N_7483);
nand U15952 (N_15952,N_50,N_7555);
nand U15953 (N_15953,N_4789,N_4773);
or U15954 (N_15954,N_270,N_1155);
xor U15955 (N_15955,N_5920,N_3773);
and U15956 (N_15956,N_6927,N_9109);
xnor U15957 (N_15957,N_2654,N_7883);
xor U15958 (N_15958,N_3064,N_6869);
xor U15959 (N_15959,N_5565,N_2332);
nor U15960 (N_15960,N_6376,N_6865);
xor U15961 (N_15961,N_3738,N_7618);
xor U15962 (N_15962,N_1175,N_3987);
and U15963 (N_15963,N_9535,N_9005);
nor U15964 (N_15964,N_2464,N_4294);
or U15965 (N_15965,N_1269,N_2702);
nand U15966 (N_15966,N_8240,N_6637);
nor U15967 (N_15967,N_1422,N_2635);
and U15968 (N_15968,N_7727,N_9980);
and U15969 (N_15969,N_4043,N_4869);
nor U15970 (N_15970,N_8667,N_9175);
nand U15971 (N_15971,N_3262,N_1951);
or U15972 (N_15972,N_7738,N_8370);
or U15973 (N_15973,N_568,N_5995);
xnor U15974 (N_15974,N_7148,N_2313);
and U15975 (N_15975,N_9972,N_6110);
nor U15976 (N_15976,N_2495,N_6210);
xnor U15977 (N_15977,N_3998,N_3010);
nand U15978 (N_15978,N_3125,N_4640);
or U15979 (N_15979,N_6719,N_1022);
xnor U15980 (N_15980,N_737,N_9824);
nor U15981 (N_15981,N_2553,N_3231);
and U15982 (N_15982,N_3426,N_9365);
nor U15983 (N_15983,N_873,N_2736);
nor U15984 (N_15984,N_8574,N_4903);
or U15985 (N_15985,N_2550,N_4694);
or U15986 (N_15986,N_7886,N_82);
nand U15987 (N_15987,N_2125,N_3340);
nor U15988 (N_15988,N_5006,N_904);
and U15989 (N_15989,N_7317,N_1282);
or U15990 (N_15990,N_245,N_6069);
or U15991 (N_15991,N_5957,N_7826);
xor U15992 (N_15992,N_4741,N_8169);
nand U15993 (N_15993,N_4317,N_6790);
and U15994 (N_15994,N_9094,N_4416);
or U15995 (N_15995,N_7836,N_3599);
xnor U15996 (N_15996,N_8536,N_8114);
and U15997 (N_15997,N_9293,N_6150);
and U15998 (N_15998,N_4791,N_7163);
and U15999 (N_15999,N_8890,N_3406);
nor U16000 (N_16000,N_4120,N_9349);
nand U16001 (N_16001,N_297,N_8857);
or U16002 (N_16002,N_7967,N_8023);
or U16003 (N_16003,N_7412,N_709);
nor U16004 (N_16004,N_3850,N_359);
xnor U16005 (N_16005,N_6452,N_8162);
and U16006 (N_16006,N_4576,N_4354);
and U16007 (N_16007,N_8466,N_5896);
or U16008 (N_16008,N_7917,N_1495);
or U16009 (N_16009,N_1742,N_4513);
nor U16010 (N_16010,N_2850,N_1623);
nor U16011 (N_16011,N_5337,N_8392);
nand U16012 (N_16012,N_8873,N_2707);
xnor U16013 (N_16013,N_6065,N_9735);
nor U16014 (N_16014,N_7177,N_2714);
xor U16015 (N_16015,N_7719,N_4370);
nor U16016 (N_16016,N_8670,N_3312);
xor U16017 (N_16017,N_7945,N_7292);
or U16018 (N_16018,N_6984,N_1032);
nand U16019 (N_16019,N_1708,N_3869);
and U16020 (N_16020,N_5007,N_4978);
and U16021 (N_16021,N_8148,N_211);
nor U16022 (N_16022,N_9891,N_4914);
xor U16023 (N_16023,N_9815,N_3623);
nor U16024 (N_16024,N_8500,N_1286);
or U16025 (N_16025,N_8551,N_6768);
or U16026 (N_16026,N_4284,N_68);
or U16027 (N_16027,N_3105,N_4771);
or U16028 (N_16028,N_4805,N_547);
xor U16029 (N_16029,N_7169,N_7988);
or U16030 (N_16030,N_5065,N_1144);
nand U16031 (N_16031,N_3982,N_9713);
nor U16032 (N_16032,N_6857,N_3415);
nand U16033 (N_16033,N_6471,N_1542);
nor U16034 (N_16034,N_5915,N_6327);
xnor U16035 (N_16035,N_8826,N_569);
and U16036 (N_16036,N_3928,N_466);
or U16037 (N_16037,N_3137,N_6934);
and U16038 (N_16038,N_196,N_3918);
or U16039 (N_16039,N_6450,N_9973);
nor U16040 (N_16040,N_236,N_1859);
xnor U16041 (N_16041,N_2315,N_388);
nand U16042 (N_16042,N_7455,N_3254);
xor U16043 (N_16043,N_7001,N_7461);
and U16044 (N_16044,N_8822,N_473);
nor U16045 (N_16045,N_2875,N_8297);
and U16046 (N_16046,N_2920,N_6942);
xor U16047 (N_16047,N_9484,N_9348);
or U16048 (N_16048,N_8981,N_3209);
nand U16049 (N_16049,N_744,N_1703);
xor U16050 (N_16050,N_5083,N_945);
or U16051 (N_16051,N_7090,N_8456);
xnor U16052 (N_16052,N_758,N_3700);
xor U16053 (N_16053,N_4178,N_2162);
or U16054 (N_16054,N_5044,N_8807);
or U16055 (N_16055,N_5914,N_9595);
xnor U16056 (N_16056,N_2289,N_9487);
xor U16057 (N_16057,N_467,N_1053);
nor U16058 (N_16058,N_5548,N_8743);
or U16059 (N_16059,N_643,N_3652);
nor U16060 (N_16060,N_9973,N_9903);
and U16061 (N_16061,N_1285,N_785);
nor U16062 (N_16062,N_527,N_6341);
nand U16063 (N_16063,N_5991,N_9961);
and U16064 (N_16064,N_1542,N_1818);
nand U16065 (N_16065,N_6965,N_5398);
xor U16066 (N_16066,N_1225,N_7240);
or U16067 (N_16067,N_87,N_9834);
nand U16068 (N_16068,N_2339,N_3877);
and U16069 (N_16069,N_4270,N_3406);
nand U16070 (N_16070,N_7293,N_793);
nand U16071 (N_16071,N_941,N_1108);
nand U16072 (N_16072,N_6974,N_8187);
and U16073 (N_16073,N_3241,N_4709);
nand U16074 (N_16074,N_5069,N_119);
nand U16075 (N_16075,N_9182,N_2459);
and U16076 (N_16076,N_1325,N_6356);
and U16077 (N_16077,N_5832,N_1327);
nand U16078 (N_16078,N_2177,N_5910);
or U16079 (N_16079,N_6793,N_9499);
nor U16080 (N_16080,N_4872,N_7091);
or U16081 (N_16081,N_3763,N_6919);
nor U16082 (N_16082,N_4717,N_2044);
xnor U16083 (N_16083,N_9265,N_6630);
nor U16084 (N_16084,N_4584,N_8514);
nor U16085 (N_16085,N_9087,N_6903);
or U16086 (N_16086,N_1744,N_1296);
and U16087 (N_16087,N_979,N_9710);
xnor U16088 (N_16088,N_5424,N_4975);
xnor U16089 (N_16089,N_2395,N_5457);
xnor U16090 (N_16090,N_3357,N_592);
xnor U16091 (N_16091,N_7308,N_7947);
nand U16092 (N_16092,N_2600,N_3262);
or U16093 (N_16093,N_5218,N_5968);
nand U16094 (N_16094,N_6953,N_8392);
nand U16095 (N_16095,N_5096,N_5613);
or U16096 (N_16096,N_232,N_6996);
or U16097 (N_16097,N_8078,N_3139);
and U16098 (N_16098,N_7547,N_5895);
or U16099 (N_16099,N_1308,N_3815);
xnor U16100 (N_16100,N_2648,N_2326);
nor U16101 (N_16101,N_6548,N_2440);
nand U16102 (N_16102,N_152,N_4686);
or U16103 (N_16103,N_48,N_8232);
nor U16104 (N_16104,N_3761,N_3519);
nor U16105 (N_16105,N_7625,N_3534);
nor U16106 (N_16106,N_6005,N_9349);
and U16107 (N_16107,N_1370,N_5700);
nor U16108 (N_16108,N_2574,N_3250);
xor U16109 (N_16109,N_8269,N_2799);
nor U16110 (N_16110,N_5179,N_8133);
nor U16111 (N_16111,N_6190,N_7819);
or U16112 (N_16112,N_5167,N_3864);
and U16113 (N_16113,N_1846,N_9651);
and U16114 (N_16114,N_174,N_5735);
or U16115 (N_16115,N_2290,N_6339);
and U16116 (N_16116,N_25,N_4836);
and U16117 (N_16117,N_4760,N_2258);
or U16118 (N_16118,N_4147,N_6706);
nand U16119 (N_16119,N_9271,N_1201);
or U16120 (N_16120,N_2202,N_4513);
nand U16121 (N_16121,N_9471,N_2489);
or U16122 (N_16122,N_3638,N_5609);
nor U16123 (N_16123,N_4085,N_3604);
nand U16124 (N_16124,N_5900,N_3918);
or U16125 (N_16125,N_1166,N_446);
nand U16126 (N_16126,N_8823,N_4031);
nand U16127 (N_16127,N_5706,N_1954);
xnor U16128 (N_16128,N_8702,N_4118);
xnor U16129 (N_16129,N_9212,N_15);
xor U16130 (N_16130,N_5284,N_5238);
nor U16131 (N_16131,N_7313,N_4719);
nand U16132 (N_16132,N_852,N_2980);
and U16133 (N_16133,N_5362,N_1669);
nor U16134 (N_16134,N_200,N_7071);
xor U16135 (N_16135,N_8972,N_7494);
and U16136 (N_16136,N_2585,N_9475);
or U16137 (N_16137,N_6486,N_6574);
nand U16138 (N_16138,N_6095,N_7668);
xnor U16139 (N_16139,N_9957,N_957);
nor U16140 (N_16140,N_6747,N_6073);
and U16141 (N_16141,N_5771,N_4760);
nor U16142 (N_16142,N_882,N_4735);
xor U16143 (N_16143,N_4256,N_8596);
nand U16144 (N_16144,N_4590,N_3166);
or U16145 (N_16145,N_1144,N_4098);
xnor U16146 (N_16146,N_9579,N_3758);
nand U16147 (N_16147,N_3452,N_7939);
xnor U16148 (N_16148,N_2503,N_7405);
nand U16149 (N_16149,N_784,N_7617);
and U16150 (N_16150,N_6641,N_1199);
nor U16151 (N_16151,N_2479,N_5421);
nor U16152 (N_16152,N_6130,N_2562);
nand U16153 (N_16153,N_9169,N_92);
nand U16154 (N_16154,N_5342,N_8946);
nor U16155 (N_16155,N_4862,N_1512);
xor U16156 (N_16156,N_5157,N_3071);
nand U16157 (N_16157,N_4779,N_4726);
nand U16158 (N_16158,N_3125,N_2478);
and U16159 (N_16159,N_6835,N_6443);
and U16160 (N_16160,N_6732,N_4652);
nor U16161 (N_16161,N_8392,N_657);
xor U16162 (N_16162,N_1335,N_5560);
and U16163 (N_16163,N_3287,N_5252);
nor U16164 (N_16164,N_1556,N_3040);
and U16165 (N_16165,N_9128,N_9865);
and U16166 (N_16166,N_1715,N_5549);
xor U16167 (N_16167,N_1133,N_6082);
nand U16168 (N_16168,N_2685,N_6388);
xnor U16169 (N_16169,N_4869,N_7703);
nor U16170 (N_16170,N_815,N_8270);
nor U16171 (N_16171,N_3216,N_236);
xnor U16172 (N_16172,N_8665,N_3833);
nor U16173 (N_16173,N_9700,N_7659);
nor U16174 (N_16174,N_5232,N_4396);
or U16175 (N_16175,N_4085,N_4421);
and U16176 (N_16176,N_3363,N_4486);
and U16177 (N_16177,N_2563,N_5435);
nor U16178 (N_16178,N_5186,N_4961);
xnor U16179 (N_16179,N_8216,N_1451);
or U16180 (N_16180,N_9576,N_4864);
xnor U16181 (N_16181,N_4777,N_2151);
nand U16182 (N_16182,N_9959,N_9211);
nor U16183 (N_16183,N_9468,N_1409);
or U16184 (N_16184,N_8610,N_7482);
or U16185 (N_16185,N_5035,N_1033);
or U16186 (N_16186,N_5893,N_3309);
nand U16187 (N_16187,N_9861,N_4074);
or U16188 (N_16188,N_1270,N_9684);
xor U16189 (N_16189,N_4786,N_7715);
or U16190 (N_16190,N_9236,N_4259);
and U16191 (N_16191,N_224,N_4123);
and U16192 (N_16192,N_5571,N_6052);
nor U16193 (N_16193,N_9628,N_8306);
and U16194 (N_16194,N_4627,N_1845);
and U16195 (N_16195,N_4737,N_405);
nor U16196 (N_16196,N_8603,N_8162);
nand U16197 (N_16197,N_5241,N_6679);
nand U16198 (N_16198,N_3313,N_2001);
and U16199 (N_16199,N_3516,N_2947);
nor U16200 (N_16200,N_3652,N_306);
nand U16201 (N_16201,N_6293,N_2391);
nand U16202 (N_16202,N_454,N_4481);
and U16203 (N_16203,N_5521,N_7737);
nor U16204 (N_16204,N_1583,N_2390);
and U16205 (N_16205,N_4438,N_4407);
nor U16206 (N_16206,N_8983,N_7823);
nand U16207 (N_16207,N_25,N_3178);
and U16208 (N_16208,N_8850,N_4452);
and U16209 (N_16209,N_6024,N_7545);
or U16210 (N_16210,N_2576,N_2158);
or U16211 (N_16211,N_2331,N_6402);
and U16212 (N_16212,N_4796,N_7718);
and U16213 (N_16213,N_2680,N_4623);
nand U16214 (N_16214,N_7480,N_9985);
nand U16215 (N_16215,N_7640,N_7118);
or U16216 (N_16216,N_2624,N_4517);
nor U16217 (N_16217,N_9388,N_6091);
or U16218 (N_16218,N_680,N_2227);
and U16219 (N_16219,N_7769,N_1929);
and U16220 (N_16220,N_1596,N_2639);
xnor U16221 (N_16221,N_7763,N_4468);
xor U16222 (N_16222,N_8032,N_9034);
nor U16223 (N_16223,N_7041,N_32);
nand U16224 (N_16224,N_4400,N_4326);
and U16225 (N_16225,N_5926,N_6594);
nor U16226 (N_16226,N_6144,N_8869);
and U16227 (N_16227,N_8987,N_8417);
or U16228 (N_16228,N_5773,N_5689);
nor U16229 (N_16229,N_1643,N_4234);
nor U16230 (N_16230,N_5650,N_921);
nor U16231 (N_16231,N_3861,N_3768);
and U16232 (N_16232,N_701,N_8772);
xnor U16233 (N_16233,N_1136,N_5988);
or U16234 (N_16234,N_4021,N_5576);
nand U16235 (N_16235,N_1165,N_5252);
and U16236 (N_16236,N_4382,N_7997);
or U16237 (N_16237,N_775,N_8619);
xor U16238 (N_16238,N_4392,N_4911);
xor U16239 (N_16239,N_9954,N_7700);
and U16240 (N_16240,N_3067,N_44);
and U16241 (N_16241,N_893,N_4004);
and U16242 (N_16242,N_1842,N_7410);
nand U16243 (N_16243,N_5044,N_1950);
or U16244 (N_16244,N_316,N_9107);
or U16245 (N_16245,N_3671,N_1387);
and U16246 (N_16246,N_6476,N_3990);
nor U16247 (N_16247,N_7322,N_6723);
or U16248 (N_16248,N_8827,N_9781);
or U16249 (N_16249,N_4345,N_8571);
nand U16250 (N_16250,N_8600,N_9020);
nand U16251 (N_16251,N_5603,N_5527);
nand U16252 (N_16252,N_3114,N_3811);
nor U16253 (N_16253,N_1030,N_8834);
or U16254 (N_16254,N_4050,N_6405);
and U16255 (N_16255,N_4791,N_9110);
nand U16256 (N_16256,N_435,N_7952);
or U16257 (N_16257,N_9554,N_8906);
xnor U16258 (N_16258,N_5627,N_1928);
nor U16259 (N_16259,N_1534,N_2551);
xnor U16260 (N_16260,N_1980,N_9878);
nand U16261 (N_16261,N_5182,N_9602);
or U16262 (N_16262,N_8272,N_2682);
nand U16263 (N_16263,N_3143,N_1603);
or U16264 (N_16264,N_8620,N_6847);
or U16265 (N_16265,N_5275,N_9247);
or U16266 (N_16266,N_6511,N_3248);
nor U16267 (N_16267,N_8685,N_4089);
nor U16268 (N_16268,N_3855,N_5579);
xnor U16269 (N_16269,N_2822,N_50);
and U16270 (N_16270,N_6712,N_7387);
xnor U16271 (N_16271,N_1844,N_3255);
and U16272 (N_16272,N_1513,N_6742);
or U16273 (N_16273,N_1902,N_3209);
nand U16274 (N_16274,N_7498,N_2480);
xnor U16275 (N_16275,N_7971,N_86);
nor U16276 (N_16276,N_509,N_8492);
and U16277 (N_16277,N_9848,N_6903);
nor U16278 (N_16278,N_8319,N_3567);
or U16279 (N_16279,N_7324,N_2123);
and U16280 (N_16280,N_3396,N_3684);
xnor U16281 (N_16281,N_1927,N_5905);
nand U16282 (N_16282,N_2330,N_2336);
or U16283 (N_16283,N_3858,N_998);
nor U16284 (N_16284,N_3816,N_5212);
nand U16285 (N_16285,N_8429,N_1556);
nor U16286 (N_16286,N_8357,N_3221);
xor U16287 (N_16287,N_4577,N_4231);
or U16288 (N_16288,N_5858,N_2126);
xor U16289 (N_16289,N_5583,N_5076);
and U16290 (N_16290,N_7007,N_3464);
nand U16291 (N_16291,N_8092,N_1393);
nand U16292 (N_16292,N_8966,N_4132);
xor U16293 (N_16293,N_9380,N_8789);
or U16294 (N_16294,N_5732,N_4584);
and U16295 (N_16295,N_8251,N_1925);
or U16296 (N_16296,N_1476,N_483);
and U16297 (N_16297,N_5709,N_8579);
and U16298 (N_16298,N_4928,N_9534);
nand U16299 (N_16299,N_1024,N_4108);
and U16300 (N_16300,N_7432,N_5602);
nor U16301 (N_16301,N_2225,N_7938);
nand U16302 (N_16302,N_6554,N_5493);
xor U16303 (N_16303,N_3981,N_7503);
nor U16304 (N_16304,N_5915,N_6744);
or U16305 (N_16305,N_4950,N_8761);
or U16306 (N_16306,N_1073,N_876);
nor U16307 (N_16307,N_8398,N_4573);
or U16308 (N_16308,N_6457,N_7740);
and U16309 (N_16309,N_2839,N_1324);
and U16310 (N_16310,N_4262,N_7881);
nor U16311 (N_16311,N_80,N_4704);
and U16312 (N_16312,N_3761,N_9941);
xnor U16313 (N_16313,N_761,N_5657);
nand U16314 (N_16314,N_7118,N_4172);
nor U16315 (N_16315,N_2859,N_9629);
xor U16316 (N_16316,N_8967,N_6052);
nand U16317 (N_16317,N_7806,N_468);
xor U16318 (N_16318,N_6755,N_113);
nor U16319 (N_16319,N_8187,N_9826);
nand U16320 (N_16320,N_6333,N_8589);
nor U16321 (N_16321,N_5195,N_3536);
and U16322 (N_16322,N_1368,N_2274);
and U16323 (N_16323,N_4935,N_7773);
xnor U16324 (N_16324,N_3119,N_4038);
xnor U16325 (N_16325,N_9633,N_3311);
nor U16326 (N_16326,N_4797,N_1961);
xor U16327 (N_16327,N_8046,N_372);
nand U16328 (N_16328,N_1232,N_778);
nand U16329 (N_16329,N_883,N_7986);
and U16330 (N_16330,N_1363,N_9955);
and U16331 (N_16331,N_371,N_8445);
nand U16332 (N_16332,N_5777,N_7652);
nand U16333 (N_16333,N_6102,N_8433);
nand U16334 (N_16334,N_2943,N_3632);
or U16335 (N_16335,N_434,N_8874);
nand U16336 (N_16336,N_7776,N_2052);
nand U16337 (N_16337,N_2140,N_4961);
and U16338 (N_16338,N_4200,N_2753);
and U16339 (N_16339,N_8032,N_7163);
or U16340 (N_16340,N_1275,N_7239);
or U16341 (N_16341,N_5499,N_3385);
nor U16342 (N_16342,N_3612,N_1552);
xor U16343 (N_16343,N_3720,N_2388);
xor U16344 (N_16344,N_6975,N_366);
or U16345 (N_16345,N_9683,N_661);
nand U16346 (N_16346,N_7653,N_8754);
nand U16347 (N_16347,N_5095,N_3947);
or U16348 (N_16348,N_9383,N_758);
nand U16349 (N_16349,N_255,N_4240);
xnor U16350 (N_16350,N_9751,N_3504);
and U16351 (N_16351,N_7978,N_2832);
xnor U16352 (N_16352,N_8235,N_3846);
nand U16353 (N_16353,N_1102,N_688);
and U16354 (N_16354,N_1393,N_8308);
xnor U16355 (N_16355,N_3230,N_2431);
or U16356 (N_16356,N_6108,N_8766);
and U16357 (N_16357,N_2643,N_5394);
xnor U16358 (N_16358,N_6751,N_7103);
nand U16359 (N_16359,N_9687,N_1861);
nor U16360 (N_16360,N_1649,N_4086);
nand U16361 (N_16361,N_8237,N_1883);
nor U16362 (N_16362,N_1856,N_7093);
nand U16363 (N_16363,N_6010,N_5746);
xnor U16364 (N_16364,N_9108,N_17);
or U16365 (N_16365,N_8753,N_3164);
nor U16366 (N_16366,N_7565,N_3086);
nor U16367 (N_16367,N_5597,N_1079);
nand U16368 (N_16368,N_11,N_7905);
nor U16369 (N_16369,N_7588,N_5903);
nand U16370 (N_16370,N_6280,N_2513);
or U16371 (N_16371,N_8956,N_7895);
xor U16372 (N_16372,N_7111,N_7978);
nor U16373 (N_16373,N_2247,N_1773);
and U16374 (N_16374,N_7303,N_3242);
and U16375 (N_16375,N_7892,N_1871);
and U16376 (N_16376,N_4102,N_3680);
nand U16377 (N_16377,N_2059,N_8791);
xnor U16378 (N_16378,N_5354,N_3258);
or U16379 (N_16379,N_2004,N_6112);
and U16380 (N_16380,N_194,N_6760);
or U16381 (N_16381,N_4390,N_6179);
or U16382 (N_16382,N_151,N_282);
or U16383 (N_16383,N_2410,N_5911);
xor U16384 (N_16384,N_605,N_6276);
nor U16385 (N_16385,N_9048,N_3988);
and U16386 (N_16386,N_394,N_3098);
and U16387 (N_16387,N_7728,N_5523);
xor U16388 (N_16388,N_2694,N_6455);
nor U16389 (N_16389,N_4363,N_2937);
nor U16390 (N_16390,N_735,N_7589);
and U16391 (N_16391,N_8302,N_3261);
or U16392 (N_16392,N_2567,N_7426);
xnor U16393 (N_16393,N_3999,N_8990);
xor U16394 (N_16394,N_2781,N_103);
and U16395 (N_16395,N_6252,N_8154);
or U16396 (N_16396,N_4370,N_4116);
xnor U16397 (N_16397,N_3114,N_5871);
nand U16398 (N_16398,N_4720,N_6766);
and U16399 (N_16399,N_649,N_4962);
or U16400 (N_16400,N_4011,N_8154);
nor U16401 (N_16401,N_423,N_6699);
or U16402 (N_16402,N_4859,N_5763);
and U16403 (N_16403,N_4504,N_1574);
xor U16404 (N_16404,N_9592,N_2112);
and U16405 (N_16405,N_2918,N_4317);
and U16406 (N_16406,N_5459,N_9450);
and U16407 (N_16407,N_3122,N_6756);
xor U16408 (N_16408,N_1775,N_3421);
or U16409 (N_16409,N_6770,N_7280);
xnor U16410 (N_16410,N_2255,N_2663);
nand U16411 (N_16411,N_6702,N_930);
and U16412 (N_16412,N_9930,N_8501);
or U16413 (N_16413,N_1969,N_8958);
nor U16414 (N_16414,N_2686,N_1535);
or U16415 (N_16415,N_7663,N_9370);
nand U16416 (N_16416,N_2517,N_3679);
and U16417 (N_16417,N_9694,N_6773);
xnor U16418 (N_16418,N_3356,N_3004);
xor U16419 (N_16419,N_20,N_7235);
or U16420 (N_16420,N_6114,N_9498);
xor U16421 (N_16421,N_7193,N_3985);
xor U16422 (N_16422,N_5758,N_51);
and U16423 (N_16423,N_8135,N_8989);
nor U16424 (N_16424,N_5308,N_5607);
nand U16425 (N_16425,N_2471,N_1929);
or U16426 (N_16426,N_4224,N_674);
or U16427 (N_16427,N_167,N_7427);
and U16428 (N_16428,N_5672,N_1799);
or U16429 (N_16429,N_2901,N_8083);
or U16430 (N_16430,N_6402,N_8030);
nor U16431 (N_16431,N_6741,N_9750);
or U16432 (N_16432,N_1246,N_590);
xnor U16433 (N_16433,N_1005,N_3165);
nor U16434 (N_16434,N_2456,N_5976);
nand U16435 (N_16435,N_6700,N_2525);
nand U16436 (N_16436,N_7243,N_1481);
nand U16437 (N_16437,N_9330,N_9092);
and U16438 (N_16438,N_5431,N_383);
nand U16439 (N_16439,N_1522,N_6861);
nor U16440 (N_16440,N_1179,N_6807);
nand U16441 (N_16441,N_1513,N_8797);
nor U16442 (N_16442,N_75,N_1410);
nor U16443 (N_16443,N_697,N_5618);
and U16444 (N_16444,N_4841,N_5691);
and U16445 (N_16445,N_5854,N_2337);
nand U16446 (N_16446,N_8683,N_144);
nor U16447 (N_16447,N_8835,N_9755);
or U16448 (N_16448,N_2403,N_1631);
xnor U16449 (N_16449,N_5684,N_7261);
and U16450 (N_16450,N_3113,N_1208);
xnor U16451 (N_16451,N_611,N_6097);
nand U16452 (N_16452,N_7773,N_4112);
and U16453 (N_16453,N_9098,N_4866);
nand U16454 (N_16454,N_6986,N_743);
nor U16455 (N_16455,N_216,N_5576);
nand U16456 (N_16456,N_6094,N_8800);
or U16457 (N_16457,N_1553,N_9178);
xnor U16458 (N_16458,N_3378,N_4945);
nor U16459 (N_16459,N_882,N_2647);
or U16460 (N_16460,N_9973,N_6938);
nor U16461 (N_16461,N_6548,N_2425);
nand U16462 (N_16462,N_8761,N_7374);
or U16463 (N_16463,N_43,N_2616);
nand U16464 (N_16464,N_1816,N_4235);
or U16465 (N_16465,N_7177,N_1843);
and U16466 (N_16466,N_1997,N_7122);
xnor U16467 (N_16467,N_8097,N_4381);
or U16468 (N_16468,N_2271,N_1518);
nand U16469 (N_16469,N_4977,N_2459);
or U16470 (N_16470,N_5992,N_6578);
xnor U16471 (N_16471,N_8958,N_6641);
nor U16472 (N_16472,N_7201,N_8212);
nand U16473 (N_16473,N_7629,N_3318);
nor U16474 (N_16474,N_9236,N_8012);
or U16475 (N_16475,N_7004,N_8145);
and U16476 (N_16476,N_5813,N_357);
xnor U16477 (N_16477,N_6260,N_9475);
xor U16478 (N_16478,N_4751,N_4689);
nor U16479 (N_16479,N_7515,N_9281);
nor U16480 (N_16480,N_7099,N_9344);
or U16481 (N_16481,N_8041,N_2942);
or U16482 (N_16482,N_5013,N_3573);
nand U16483 (N_16483,N_872,N_994);
nor U16484 (N_16484,N_6363,N_2054);
or U16485 (N_16485,N_7178,N_5738);
or U16486 (N_16486,N_516,N_787);
and U16487 (N_16487,N_5564,N_167);
nand U16488 (N_16488,N_6745,N_4839);
nand U16489 (N_16489,N_803,N_327);
nand U16490 (N_16490,N_9692,N_5253);
and U16491 (N_16491,N_2172,N_8269);
xor U16492 (N_16492,N_4874,N_2003);
or U16493 (N_16493,N_7693,N_8510);
nand U16494 (N_16494,N_6702,N_3939);
and U16495 (N_16495,N_1932,N_6945);
xnor U16496 (N_16496,N_5206,N_7835);
nor U16497 (N_16497,N_9011,N_2037);
nor U16498 (N_16498,N_5157,N_4806);
and U16499 (N_16499,N_2773,N_7292);
and U16500 (N_16500,N_2985,N_319);
and U16501 (N_16501,N_2762,N_2445);
nand U16502 (N_16502,N_8649,N_1638);
or U16503 (N_16503,N_7685,N_3244);
or U16504 (N_16504,N_5661,N_1512);
nor U16505 (N_16505,N_5604,N_4633);
or U16506 (N_16506,N_3502,N_3753);
or U16507 (N_16507,N_1091,N_353);
and U16508 (N_16508,N_336,N_4222);
xor U16509 (N_16509,N_5441,N_7295);
nor U16510 (N_16510,N_5612,N_1891);
or U16511 (N_16511,N_1924,N_2164);
nor U16512 (N_16512,N_2304,N_2719);
or U16513 (N_16513,N_7346,N_1091);
or U16514 (N_16514,N_4467,N_8165);
xnor U16515 (N_16515,N_3697,N_9604);
nor U16516 (N_16516,N_9548,N_2667);
nor U16517 (N_16517,N_902,N_4971);
nor U16518 (N_16518,N_7005,N_1308);
nor U16519 (N_16519,N_6332,N_344);
or U16520 (N_16520,N_7960,N_9577);
or U16521 (N_16521,N_8350,N_3346);
or U16522 (N_16522,N_9770,N_2999);
and U16523 (N_16523,N_756,N_4957);
nand U16524 (N_16524,N_2309,N_166);
and U16525 (N_16525,N_9193,N_6884);
and U16526 (N_16526,N_8670,N_90);
nor U16527 (N_16527,N_8602,N_2511);
nor U16528 (N_16528,N_649,N_5947);
xor U16529 (N_16529,N_5144,N_3078);
nor U16530 (N_16530,N_5962,N_5386);
nor U16531 (N_16531,N_9395,N_998);
and U16532 (N_16532,N_1071,N_1660);
xor U16533 (N_16533,N_3343,N_223);
xnor U16534 (N_16534,N_8516,N_393);
xnor U16535 (N_16535,N_8779,N_3406);
and U16536 (N_16536,N_541,N_211);
nand U16537 (N_16537,N_313,N_7760);
xor U16538 (N_16538,N_2072,N_4183);
or U16539 (N_16539,N_1644,N_3157);
xnor U16540 (N_16540,N_3843,N_5292);
and U16541 (N_16541,N_1599,N_523);
xor U16542 (N_16542,N_9722,N_1816);
nor U16543 (N_16543,N_5892,N_9507);
or U16544 (N_16544,N_5611,N_5580);
and U16545 (N_16545,N_4338,N_6249);
nor U16546 (N_16546,N_8775,N_8065);
nand U16547 (N_16547,N_6086,N_3099);
and U16548 (N_16548,N_9795,N_4835);
or U16549 (N_16549,N_646,N_6726);
and U16550 (N_16550,N_3535,N_3337);
xor U16551 (N_16551,N_13,N_4680);
xnor U16552 (N_16552,N_2262,N_907);
or U16553 (N_16553,N_380,N_4927);
nor U16554 (N_16554,N_7136,N_4191);
and U16555 (N_16555,N_783,N_5253);
and U16556 (N_16556,N_3409,N_5827);
nand U16557 (N_16557,N_2609,N_8348);
and U16558 (N_16558,N_929,N_8729);
and U16559 (N_16559,N_2655,N_9226);
and U16560 (N_16560,N_9857,N_6305);
or U16561 (N_16561,N_5752,N_8349);
nor U16562 (N_16562,N_1648,N_4349);
or U16563 (N_16563,N_8284,N_8961);
and U16564 (N_16564,N_9439,N_2350);
xnor U16565 (N_16565,N_8938,N_5604);
nor U16566 (N_16566,N_2834,N_9601);
and U16567 (N_16567,N_4028,N_3149);
xor U16568 (N_16568,N_128,N_6709);
or U16569 (N_16569,N_9454,N_92);
or U16570 (N_16570,N_9787,N_2888);
or U16571 (N_16571,N_3093,N_7358);
xor U16572 (N_16572,N_6802,N_8304);
and U16573 (N_16573,N_5902,N_2829);
nor U16574 (N_16574,N_5957,N_5423);
xnor U16575 (N_16575,N_2123,N_2598);
and U16576 (N_16576,N_8423,N_7359);
and U16577 (N_16577,N_3646,N_3598);
and U16578 (N_16578,N_3334,N_9761);
and U16579 (N_16579,N_4926,N_6855);
xor U16580 (N_16580,N_2258,N_785);
xnor U16581 (N_16581,N_3922,N_8656);
xor U16582 (N_16582,N_4303,N_5743);
nor U16583 (N_16583,N_4832,N_1191);
xnor U16584 (N_16584,N_3960,N_4478);
nor U16585 (N_16585,N_9722,N_5038);
xor U16586 (N_16586,N_1863,N_7198);
nand U16587 (N_16587,N_9941,N_1668);
and U16588 (N_16588,N_1180,N_7215);
and U16589 (N_16589,N_1434,N_3493);
or U16590 (N_16590,N_9220,N_4618);
nand U16591 (N_16591,N_145,N_1177);
xor U16592 (N_16592,N_4273,N_1006);
nand U16593 (N_16593,N_4650,N_6288);
nand U16594 (N_16594,N_3322,N_6631);
and U16595 (N_16595,N_7023,N_5811);
and U16596 (N_16596,N_9221,N_3668);
and U16597 (N_16597,N_32,N_3994);
and U16598 (N_16598,N_2581,N_776);
nor U16599 (N_16599,N_8576,N_5);
and U16600 (N_16600,N_673,N_1745);
and U16601 (N_16601,N_884,N_9487);
and U16602 (N_16602,N_4050,N_2766);
nor U16603 (N_16603,N_5821,N_1524);
xor U16604 (N_16604,N_2588,N_742);
nor U16605 (N_16605,N_6009,N_510);
or U16606 (N_16606,N_1656,N_3172);
nor U16607 (N_16607,N_7910,N_9992);
or U16608 (N_16608,N_8928,N_1711);
and U16609 (N_16609,N_7815,N_8881);
and U16610 (N_16610,N_4568,N_6556);
xnor U16611 (N_16611,N_1411,N_297);
nor U16612 (N_16612,N_352,N_7492);
xnor U16613 (N_16613,N_2512,N_7613);
nand U16614 (N_16614,N_2333,N_1343);
or U16615 (N_16615,N_7406,N_4973);
xor U16616 (N_16616,N_2248,N_2096);
nand U16617 (N_16617,N_3480,N_4023);
and U16618 (N_16618,N_8758,N_7507);
or U16619 (N_16619,N_1488,N_5733);
xnor U16620 (N_16620,N_7660,N_6189);
nand U16621 (N_16621,N_4430,N_5368);
nand U16622 (N_16622,N_6644,N_8477);
xnor U16623 (N_16623,N_626,N_7848);
nor U16624 (N_16624,N_3837,N_6649);
xor U16625 (N_16625,N_5026,N_5281);
nor U16626 (N_16626,N_2249,N_4788);
nand U16627 (N_16627,N_5942,N_9198);
nor U16628 (N_16628,N_3214,N_504);
xnor U16629 (N_16629,N_1300,N_496);
and U16630 (N_16630,N_2863,N_9379);
and U16631 (N_16631,N_9306,N_5379);
and U16632 (N_16632,N_2895,N_1066);
or U16633 (N_16633,N_2220,N_7780);
nand U16634 (N_16634,N_8343,N_1389);
nor U16635 (N_16635,N_3937,N_6859);
xnor U16636 (N_16636,N_9978,N_4819);
or U16637 (N_16637,N_6970,N_1113);
xor U16638 (N_16638,N_2208,N_7647);
nand U16639 (N_16639,N_4393,N_7314);
nand U16640 (N_16640,N_5680,N_9252);
and U16641 (N_16641,N_1368,N_4634);
or U16642 (N_16642,N_274,N_1943);
nor U16643 (N_16643,N_1903,N_3168);
nand U16644 (N_16644,N_5722,N_3301);
nand U16645 (N_16645,N_8319,N_8133);
nor U16646 (N_16646,N_3776,N_1671);
or U16647 (N_16647,N_9233,N_1568);
nand U16648 (N_16648,N_7203,N_3072);
xor U16649 (N_16649,N_2013,N_5843);
or U16650 (N_16650,N_6339,N_892);
or U16651 (N_16651,N_8993,N_8421);
nor U16652 (N_16652,N_4308,N_7750);
nor U16653 (N_16653,N_3004,N_3598);
xor U16654 (N_16654,N_5579,N_4314);
nor U16655 (N_16655,N_7574,N_1218);
xnor U16656 (N_16656,N_9503,N_8548);
nand U16657 (N_16657,N_8007,N_3313);
xnor U16658 (N_16658,N_1777,N_4517);
or U16659 (N_16659,N_4648,N_2461);
or U16660 (N_16660,N_9255,N_8488);
or U16661 (N_16661,N_9180,N_6491);
nand U16662 (N_16662,N_1257,N_5888);
or U16663 (N_16663,N_26,N_8061);
nand U16664 (N_16664,N_579,N_3904);
or U16665 (N_16665,N_3232,N_6859);
or U16666 (N_16666,N_8969,N_8558);
and U16667 (N_16667,N_6137,N_3916);
xnor U16668 (N_16668,N_6659,N_3059);
nor U16669 (N_16669,N_4589,N_8072);
nand U16670 (N_16670,N_1931,N_6860);
and U16671 (N_16671,N_8503,N_2058);
or U16672 (N_16672,N_6532,N_1728);
or U16673 (N_16673,N_9318,N_6370);
xor U16674 (N_16674,N_9287,N_1786);
or U16675 (N_16675,N_4234,N_727);
xor U16676 (N_16676,N_1003,N_8315);
nor U16677 (N_16677,N_4065,N_5166);
nand U16678 (N_16678,N_8308,N_3762);
nor U16679 (N_16679,N_1978,N_1943);
and U16680 (N_16680,N_6707,N_3492);
and U16681 (N_16681,N_8028,N_1158);
and U16682 (N_16682,N_5455,N_586);
xor U16683 (N_16683,N_9553,N_2284);
xnor U16684 (N_16684,N_9211,N_4752);
or U16685 (N_16685,N_7417,N_2470);
or U16686 (N_16686,N_97,N_7708);
xor U16687 (N_16687,N_4762,N_2683);
nand U16688 (N_16688,N_2554,N_7279);
xnor U16689 (N_16689,N_3953,N_4280);
and U16690 (N_16690,N_9549,N_2447);
xor U16691 (N_16691,N_9980,N_1103);
xor U16692 (N_16692,N_2174,N_2335);
nand U16693 (N_16693,N_9922,N_9403);
xnor U16694 (N_16694,N_8337,N_8784);
nor U16695 (N_16695,N_5820,N_353);
or U16696 (N_16696,N_992,N_3463);
and U16697 (N_16697,N_7073,N_384);
xor U16698 (N_16698,N_224,N_7028);
nand U16699 (N_16699,N_2389,N_3083);
xor U16700 (N_16700,N_5118,N_390);
nand U16701 (N_16701,N_6357,N_4044);
nand U16702 (N_16702,N_9435,N_1163);
nand U16703 (N_16703,N_9216,N_7797);
or U16704 (N_16704,N_2012,N_7387);
nand U16705 (N_16705,N_9895,N_168);
or U16706 (N_16706,N_2597,N_1409);
xnor U16707 (N_16707,N_7742,N_5302);
nand U16708 (N_16708,N_6091,N_4935);
nand U16709 (N_16709,N_8164,N_1690);
and U16710 (N_16710,N_6972,N_420);
nand U16711 (N_16711,N_616,N_924);
nor U16712 (N_16712,N_4685,N_9751);
or U16713 (N_16713,N_8547,N_3887);
xnor U16714 (N_16714,N_8627,N_9094);
nor U16715 (N_16715,N_7578,N_98);
nand U16716 (N_16716,N_8049,N_7341);
nand U16717 (N_16717,N_5219,N_7415);
xor U16718 (N_16718,N_5829,N_6799);
xnor U16719 (N_16719,N_7986,N_7454);
nand U16720 (N_16720,N_1759,N_240);
or U16721 (N_16721,N_2270,N_9373);
nor U16722 (N_16722,N_7602,N_4728);
nor U16723 (N_16723,N_5310,N_5109);
and U16724 (N_16724,N_1323,N_9242);
xor U16725 (N_16725,N_2071,N_8801);
nor U16726 (N_16726,N_4853,N_8822);
or U16727 (N_16727,N_4742,N_9262);
xnor U16728 (N_16728,N_6432,N_4490);
or U16729 (N_16729,N_246,N_5943);
nor U16730 (N_16730,N_5171,N_89);
nand U16731 (N_16731,N_1568,N_7441);
and U16732 (N_16732,N_1257,N_5856);
xor U16733 (N_16733,N_8438,N_2688);
or U16734 (N_16734,N_9035,N_4169);
xnor U16735 (N_16735,N_8471,N_8617);
nor U16736 (N_16736,N_6506,N_5236);
xor U16737 (N_16737,N_6834,N_5674);
nand U16738 (N_16738,N_2494,N_7469);
xnor U16739 (N_16739,N_7369,N_4676);
or U16740 (N_16740,N_4334,N_2198);
nand U16741 (N_16741,N_6335,N_6399);
or U16742 (N_16742,N_6923,N_1403);
nor U16743 (N_16743,N_6120,N_5325);
and U16744 (N_16744,N_2095,N_7030);
and U16745 (N_16745,N_4996,N_5567);
or U16746 (N_16746,N_1325,N_4270);
and U16747 (N_16747,N_6520,N_542);
or U16748 (N_16748,N_3619,N_1265);
xor U16749 (N_16749,N_5575,N_7357);
nor U16750 (N_16750,N_3725,N_1947);
xor U16751 (N_16751,N_4083,N_5388);
nor U16752 (N_16752,N_9214,N_8728);
nand U16753 (N_16753,N_3221,N_4576);
nor U16754 (N_16754,N_9375,N_490);
nor U16755 (N_16755,N_3448,N_5242);
xor U16756 (N_16756,N_7516,N_2896);
nor U16757 (N_16757,N_1486,N_8130);
and U16758 (N_16758,N_8916,N_5508);
or U16759 (N_16759,N_4221,N_7401);
nand U16760 (N_16760,N_1885,N_5136);
xor U16761 (N_16761,N_9165,N_6885);
nor U16762 (N_16762,N_2369,N_2060);
nand U16763 (N_16763,N_4990,N_6265);
and U16764 (N_16764,N_8239,N_8229);
and U16765 (N_16765,N_3771,N_4686);
xnor U16766 (N_16766,N_7794,N_4916);
xnor U16767 (N_16767,N_4341,N_2561);
or U16768 (N_16768,N_615,N_5951);
and U16769 (N_16769,N_2897,N_8844);
nand U16770 (N_16770,N_2625,N_6824);
nand U16771 (N_16771,N_7537,N_5650);
nand U16772 (N_16772,N_9083,N_1278);
xor U16773 (N_16773,N_7014,N_1470);
and U16774 (N_16774,N_3688,N_4061);
and U16775 (N_16775,N_6533,N_3066);
or U16776 (N_16776,N_797,N_5813);
nand U16777 (N_16777,N_9751,N_9090);
or U16778 (N_16778,N_3417,N_6902);
and U16779 (N_16779,N_2335,N_8105);
xnor U16780 (N_16780,N_2472,N_9678);
xnor U16781 (N_16781,N_5278,N_6081);
nor U16782 (N_16782,N_5831,N_7643);
or U16783 (N_16783,N_4845,N_2711);
xor U16784 (N_16784,N_8754,N_290);
nor U16785 (N_16785,N_1564,N_9161);
or U16786 (N_16786,N_3853,N_6485);
nor U16787 (N_16787,N_4310,N_4002);
nor U16788 (N_16788,N_2852,N_4458);
nand U16789 (N_16789,N_6912,N_1721);
and U16790 (N_16790,N_7642,N_7367);
nor U16791 (N_16791,N_6160,N_2249);
nor U16792 (N_16792,N_4743,N_3328);
xor U16793 (N_16793,N_5799,N_8751);
xnor U16794 (N_16794,N_1020,N_9243);
or U16795 (N_16795,N_415,N_8083);
or U16796 (N_16796,N_2582,N_2537);
nand U16797 (N_16797,N_4449,N_1924);
nor U16798 (N_16798,N_5845,N_6012);
and U16799 (N_16799,N_9110,N_1181);
nand U16800 (N_16800,N_4232,N_8070);
nor U16801 (N_16801,N_5529,N_4089);
and U16802 (N_16802,N_7789,N_7748);
nor U16803 (N_16803,N_2476,N_1075);
xnor U16804 (N_16804,N_432,N_8729);
nand U16805 (N_16805,N_1559,N_1278);
nand U16806 (N_16806,N_4936,N_8417);
xnor U16807 (N_16807,N_7351,N_291);
or U16808 (N_16808,N_9275,N_8836);
or U16809 (N_16809,N_2650,N_8268);
nor U16810 (N_16810,N_1326,N_9661);
xor U16811 (N_16811,N_7197,N_157);
nand U16812 (N_16812,N_3639,N_5216);
xor U16813 (N_16813,N_6147,N_7196);
xor U16814 (N_16814,N_631,N_3431);
xor U16815 (N_16815,N_4138,N_2431);
xor U16816 (N_16816,N_2045,N_8239);
and U16817 (N_16817,N_280,N_3968);
and U16818 (N_16818,N_8956,N_2822);
or U16819 (N_16819,N_7438,N_3784);
xor U16820 (N_16820,N_1113,N_8590);
nor U16821 (N_16821,N_3114,N_6777);
nand U16822 (N_16822,N_6288,N_7425);
xor U16823 (N_16823,N_1886,N_7036);
nand U16824 (N_16824,N_1582,N_2359);
and U16825 (N_16825,N_2296,N_8322);
nand U16826 (N_16826,N_9826,N_9288);
xor U16827 (N_16827,N_622,N_4018);
nor U16828 (N_16828,N_8594,N_4861);
and U16829 (N_16829,N_2440,N_6104);
xor U16830 (N_16830,N_5853,N_7859);
or U16831 (N_16831,N_2342,N_4985);
or U16832 (N_16832,N_8529,N_2565);
and U16833 (N_16833,N_5192,N_4924);
and U16834 (N_16834,N_1360,N_7052);
nand U16835 (N_16835,N_4215,N_9966);
and U16836 (N_16836,N_442,N_3676);
and U16837 (N_16837,N_9336,N_6929);
and U16838 (N_16838,N_9387,N_9611);
nand U16839 (N_16839,N_5102,N_5429);
xor U16840 (N_16840,N_3786,N_8462);
nor U16841 (N_16841,N_6148,N_4202);
or U16842 (N_16842,N_2777,N_2486);
nand U16843 (N_16843,N_2877,N_2305);
or U16844 (N_16844,N_9891,N_7460);
nand U16845 (N_16845,N_5551,N_6260);
or U16846 (N_16846,N_5114,N_1108);
nand U16847 (N_16847,N_2667,N_3913);
xnor U16848 (N_16848,N_9508,N_1342);
nand U16849 (N_16849,N_85,N_3691);
xor U16850 (N_16850,N_9935,N_1897);
nand U16851 (N_16851,N_4538,N_9741);
or U16852 (N_16852,N_8611,N_466);
xor U16853 (N_16853,N_2505,N_8483);
xnor U16854 (N_16854,N_6583,N_5477);
xnor U16855 (N_16855,N_8385,N_8745);
nand U16856 (N_16856,N_1983,N_3538);
or U16857 (N_16857,N_5286,N_1262);
nand U16858 (N_16858,N_3872,N_1514);
and U16859 (N_16859,N_5736,N_6604);
or U16860 (N_16860,N_5469,N_7644);
nor U16861 (N_16861,N_3693,N_4322);
xnor U16862 (N_16862,N_5197,N_6967);
or U16863 (N_16863,N_6934,N_7870);
and U16864 (N_16864,N_9238,N_1211);
nand U16865 (N_16865,N_7429,N_2896);
and U16866 (N_16866,N_7065,N_6821);
or U16867 (N_16867,N_3157,N_3328);
and U16868 (N_16868,N_7566,N_3184);
or U16869 (N_16869,N_9778,N_9689);
nand U16870 (N_16870,N_7324,N_2962);
nor U16871 (N_16871,N_8663,N_27);
and U16872 (N_16872,N_6597,N_6140);
nand U16873 (N_16873,N_1904,N_9823);
nor U16874 (N_16874,N_1415,N_9905);
or U16875 (N_16875,N_640,N_4478);
or U16876 (N_16876,N_1989,N_3746);
nor U16877 (N_16877,N_8864,N_8596);
or U16878 (N_16878,N_584,N_2786);
or U16879 (N_16879,N_6422,N_7807);
and U16880 (N_16880,N_7487,N_2858);
and U16881 (N_16881,N_169,N_7657);
xor U16882 (N_16882,N_4233,N_3416);
and U16883 (N_16883,N_428,N_2944);
xor U16884 (N_16884,N_4071,N_1237);
nand U16885 (N_16885,N_6065,N_2906);
xor U16886 (N_16886,N_7574,N_433);
and U16887 (N_16887,N_520,N_6777);
nand U16888 (N_16888,N_9070,N_7403);
nand U16889 (N_16889,N_8823,N_1817);
nand U16890 (N_16890,N_5735,N_8562);
or U16891 (N_16891,N_4372,N_3537);
nor U16892 (N_16892,N_7863,N_205);
xor U16893 (N_16893,N_3301,N_3484);
nor U16894 (N_16894,N_3312,N_2026);
nor U16895 (N_16895,N_2679,N_4253);
xor U16896 (N_16896,N_6493,N_6727);
xnor U16897 (N_16897,N_5146,N_6055);
nor U16898 (N_16898,N_6002,N_6800);
nor U16899 (N_16899,N_774,N_9142);
xor U16900 (N_16900,N_5357,N_1698);
nand U16901 (N_16901,N_9665,N_2944);
nand U16902 (N_16902,N_4133,N_4760);
or U16903 (N_16903,N_5047,N_2830);
nor U16904 (N_16904,N_6879,N_4603);
nand U16905 (N_16905,N_1087,N_7884);
or U16906 (N_16906,N_6217,N_8992);
and U16907 (N_16907,N_4037,N_26);
nand U16908 (N_16908,N_303,N_3126);
nor U16909 (N_16909,N_2925,N_3458);
and U16910 (N_16910,N_2749,N_9426);
nor U16911 (N_16911,N_7073,N_7876);
xor U16912 (N_16912,N_1696,N_5540);
nand U16913 (N_16913,N_3476,N_2902);
nor U16914 (N_16914,N_4374,N_6534);
nor U16915 (N_16915,N_8228,N_4622);
nand U16916 (N_16916,N_7553,N_7175);
nand U16917 (N_16917,N_1378,N_7926);
and U16918 (N_16918,N_9762,N_3164);
nor U16919 (N_16919,N_678,N_1881);
xnor U16920 (N_16920,N_9416,N_2718);
xnor U16921 (N_16921,N_1592,N_9994);
and U16922 (N_16922,N_693,N_475);
nor U16923 (N_16923,N_4075,N_7584);
or U16924 (N_16924,N_5161,N_2309);
or U16925 (N_16925,N_2417,N_9528);
xnor U16926 (N_16926,N_7787,N_6811);
and U16927 (N_16927,N_4051,N_2290);
nor U16928 (N_16928,N_8746,N_3530);
xor U16929 (N_16929,N_5339,N_4746);
xnor U16930 (N_16930,N_251,N_486);
and U16931 (N_16931,N_3697,N_7844);
nor U16932 (N_16932,N_134,N_1095);
nand U16933 (N_16933,N_4338,N_3074);
xnor U16934 (N_16934,N_5860,N_6772);
nor U16935 (N_16935,N_2404,N_6009);
and U16936 (N_16936,N_3686,N_8375);
or U16937 (N_16937,N_532,N_2315);
or U16938 (N_16938,N_4379,N_6140);
nor U16939 (N_16939,N_1017,N_3211);
xnor U16940 (N_16940,N_453,N_8335);
nand U16941 (N_16941,N_2267,N_1568);
and U16942 (N_16942,N_2617,N_5435);
xnor U16943 (N_16943,N_6861,N_3407);
and U16944 (N_16944,N_567,N_9357);
or U16945 (N_16945,N_4853,N_6602);
nand U16946 (N_16946,N_6286,N_2343);
xor U16947 (N_16947,N_6929,N_9905);
or U16948 (N_16948,N_951,N_5526);
and U16949 (N_16949,N_366,N_1442);
nand U16950 (N_16950,N_6551,N_7071);
or U16951 (N_16951,N_3299,N_3461);
nand U16952 (N_16952,N_4809,N_3007);
and U16953 (N_16953,N_7449,N_6501);
or U16954 (N_16954,N_7939,N_205);
nor U16955 (N_16955,N_8214,N_9024);
and U16956 (N_16956,N_9993,N_1442);
nor U16957 (N_16957,N_2436,N_5803);
and U16958 (N_16958,N_2619,N_529);
and U16959 (N_16959,N_7731,N_1912);
xnor U16960 (N_16960,N_9391,N_6139);
nand U16961 (N_16961,N_3852,N_5292);
nand U16962 (N_16962,N_5382,N_8883);
xnor U16963 (N_16963,N_5887,N_7652);
and U16964 (N_16964,N_1199,N_7909);
or U16965 (N_16965,N_7643,N_7602);
nor U16966 (N_16966,N_9095,N_6349);
or U16967 (N_16967,N_3811,N_6155);
nand U16968 (N_16968,N_5949,N_8443);
or U16969 (N_16969,N_1675,N_2285);
or U16970 (N_16970,N_4385,N_3006);
nor U16971 (N_16971,N_2248,N_8058);
and U16972 (N_16972,N_4040,N_9904);
xnor U16973 (N_16973,N_8326,N_9446);
nor U16974 (N_16974,N_26,N_1385);
or U16975 (N_16975,N_2159,N_7587);
nor U16976 (N_16976,N_368,N_7741);
and U16977 (N_16977,N_5071,N_9940);
nand U16978 (N_16978,N_3934,N_996);
and U16979 (N_16979,N_6267,N_3295);
and U16980 (N_16980,N_9572,N_4917);
nor U16981 (N_16981,N_4164,N_1300);
or U16982 (N_16982,N_3358,N_4031);
xor U16983 (N_16983,N_5737,N_6447);
or U16984 (N_16984,N_4151,N_9034);
xor U16985 (N_16985,N_9936,N_5242);
xnor U16986 (N_16986,N_225,N_563);
or U16987 (N_16987,N_7183,N_4776);
or U16988 (N_16988,N_7369,N_1403);
nor U16989 (N_16989,N_4859,N_6234);
and U16990 (N_16990,N_4529,N_9453);
nand U16991 (N_16991,N_6746,N_1978);
or U16992 (N_16992,N_8895,N_160);
or U16993 (N_16993,N_5505,N_5806);
or U16994 (N_16994,N_1391,N_3400);
xnor U16995 (N_16995,N_2945,N_9706);
or U16996 (N_16996,N_5780,N_4055);
nor U16997 (N_16997,N_9531,N_6809);
and U16998 (N_16998,N_5346,N_7820);
and U16999 (N_16999,N_6644,N_1306);
xor U17000 (N_17000,N_2678,N_237);
nor U17001 (N_17001,N_8422,N_2365);
xnor U17002 (N_17002,N_8341,N_3315);
nand U17003 (N_17003,N_3828,N_8664);
xor U17004 (N_17004,N_3507,N_4679);
and U17005 (N_17005,N_5979,N_4648);
xor U17006 (N_17006,N_2407,N_8376);
nor U17007 (N_17007,N_3500,N_8347);
and U17008 (N_17008,N_5768,N_221);
and U17009 (N_17009,N_5241,N_522);
and U17010 (N_17010,N_6610,N_2485);
and U17011 (N_17011,N_8429,N_5118);
nor U17012 (N_17012,N_3366,N_865);
nor U17013 (N_17013,N_2083,N_8021);
or U17014 (N_17014,N_8387,N_501);
nor U17015 (N_17015,N_5654,N_3710);
nor U17016 (N_17016,N_581,N_297);
and U17017 (N_17017,N_3301,N_4413);
or U17018 (N_17018,N_7009,N_7570);
or U17019 (N_17019,N_3997,N_8839);
nand U17020 (N_17020,N_3133,N_3393);
and U17021 (N_17021,N_7619,N_2290);
or U17022 (N_17022,N_1263,N_8535);
xnor U17023 (N_17023,N_1869,N_4450);
or U17024 (N_17024,N_9499,N_1645);
or U17025 (N_17025,N_9863,N_2335);
nor U17026 (N_17026,N_7959,N_2563);
or U17027 (N_17027,N_6164,N_4439);
nand U17028 (N_17028,N_5837,N_1401);
or U17029 (N_17029,N_9668,N_4498);
and U17030 (N_17030,N_4199,N_3816);
xnor U17031 (N_17031,N_4055,N_4297);
nand U17032 (N_17032,N_1306,N_395);
xor U17033 (N_17033,N_8945,N_9560);
xor U17034 (N_17034,N_7273,N_7904);
and U17035 (N_17035,N_4023,N_8987);
xor U17036 (N_17036,N_9537,N_440);
or U17037 (N_17037,N_8397,N_7542);
xor U17038 (N_17038,N_2456,N_3231);
and U17039 (N_17039,N_8465,N_5906);
nor U17040 (N_17040,N_1291,N_1176);
or U17041 (N_17041,N_6491,N_3685);
xor U17042 (N_17042,N_3678,N_2623);
and U17043 (N_17043,N_4006,N_715);
nor U17044 (N_17044,N_7343,N_4908);
xnor U17045 (N_17045,N_1203,N_5909);
or U17046 (N_17046,N_8998,N_8191);
xnor U17047 (N_17047,N_6234,N_4630);
xor U17048 (N_17048,N_1820,N_3685);
and U17049 (N_17049,N_9550,N_5065);
or U17050 (N_17050,N_6767,N_2860);
xnor U17051 (N_17051,N_3248,N_6486);
nand U17052 (N_17052,N_7295,N_9715);
nor U17053 (N_17053,N_6330,N_8036);
nor U17054 (N_17054,N_6549,N_9159);
nand U17055 (N_17055,N_7784,N_36);
or U17056 (N_17056,N_4122,N_7230);
and U17057 (N_17057,N_3779,N_9001);
nor U17058 (N_17058,N_5667,N_3091);
nand U17059 (N_17059,N_4280,N_6472);
nor U17060 (N_17060,N_1468,N_8287);
or U17061 (N_17061,N_4175,N_3726);
nand U17062 (N_17062,N_4930,N_7876);
nor U17063 (N_17063,N_3749,N_9553);
nand U17064 (N_17064,N_8771,N_5264);
nand U17065 (N_17065,N_5130,N_4231);
xnor U17066 (N_17066,N_9549,N_9807);
nand U17067 (N_17067,N_5313,N_4057);
nand U17068 (N_17068,N_4136,N_524);
nand U17069 (N_17069,N_7101,N_3501);
or U17070 (N_17070,N_4617,N_2675);
or U17071 (N_17071,N_7654,N_3477);
and U17072 (N_17072,N_8798,N_4718);
nor U17073 (N_17073,N_1835,N_1103);
nor U17074 (N_17074,N_2949,N_3380);
and U17075 (N_17075,N_9383,N_8346);
and U17076 (N_17076,N_2674,N_4937);
and U17077 (N_17077,N_4558,N_6535);
xor U17078 (N_17078,N_8695,N_9624);
or U17079 (N_17079,N_2675,N_7750);
xnor U17080 (N_17080,N_390,N_922);
or U17081 (N_17081,N_8266,N_9191);
nor U17082 (N_17082,N_8753,N_6201);
or U17083 (N_17083,N_3177,N_1512);
or U17084 (N_17084,N_2556,N_8645);
nor U17085 (N_17085,N_1519,N_146);
xnor U17086 (N_17086,N_7691,N_6203);
nor U17087 (N_17087,N_6434,N_1757);
nand U17088 (N_17088,N_6110,N_9637);
nand U17089 (N_17089,N_4344,N_8482);
and U17090 (N_17090,N_1188,N_5624);
or U17091 (N_17091,N_6615,N_4431);
and U17092 (N_17092,N_975,N_1720);
nand U17093 (N_17093,N_469,N_5942);
nand U17094 (N_17094,N_2315,N_1878);
and U17095 (N_17095,N_2861,N_2426);
xnor U17096 (N_17096,N_968,N_1216);
or U17097 (N_17097,N_720,N_6683);
xor U17098 (N_17098,N_3507,N_79);
or U17099 (N_17099,N_7273,N_4157);
xor U17100 (N_17100,N_9286,N_2934);
nand U17101 (N_17101,N_6000,N_6508);
xor U17102 (N_17102,N_6959,N_7665);
and U17103 (N_17103,N_6872,N_4749);
or U17104 (N_17104,N_6625,N_5200);
or U17105 (N_17105,N_7408,N_7587);
or U17106 (N_17106,N_646,N_4708);
xnor U17107 (N_17107,N_8306,N_4968);
or U17108 (N_17108,N_8243,N_8869);
nand U17109 (N_17109,N_7776,N_8698);
nand U17110 (N_17110,N_5328,N_609);
and U17111 (N_17111,N_9052,N_3038);
nor U17112 (N_17112,N_8957,N_8912);
nand U17113 (N_17113,N_5729,N_3599);
nand U17114 (N_17114,N_8957,N_1441);
xnor U17115 (N_17115,N_7285,N_3312);
nand U17116 (N_17116,N_2689,N_7133);
nand U17117 (N_17117,N_9314,N_4639);
nand U17118 (N_17118,N_171,N_3784);
and U17119 (N_17119,N_862,N_5848);
and U17120 (N_17120,N_4115,N_4705);
nor U17121 (N_17121,N_8757,N_9032);
nand U17122 (N_17122,N_4529,N_7381);
xnor U17123 (N_17123,N_7301,N_3892);
xor U17124 (N_17124,N_9101,N_6008);
or U17125 (N_17125,N_8406,N_7459);
xor U17126 (N_17126,N_3586,N_4959);
or U17127 (N_17127,N_9259,N_9153);
or U17128 (N_17128,N_7250,N_645);
nor U17129 (N_17129,N_5754,N_1901);
or U17130 (N_17130,N_9641,N_5475);
nand U17131 (N_17131,N_2333,N_9955);
xnor U17132 (N_17132,N_1289,N_7030);
xor U17133 (N_17133,N_1563,N_5536);
and U17134 (N_17134,N_1166,N_2390);
or U17135 (N_17135,N_4832,N_5385);
xnor U17136 (N_17136,N_8135,N_6917);
or U17137 (N_17137,N_4526,N_5689);
xnor U17138 (N_17138,N_2220,N_2127);
nand U17139 (N_17139,N_1101,N_827);
nor U17140 (N_17140,N_7039,N_5122);
nor U17141 (N_17141,N_483,N_5280);
xor U17142 (N_17142,N_4389,N_1118);
or U17143 (N_17143,N_6340,N_1311);
and U17144 (N_17144,N_7743,N_9358);
nor U17145 (N_17145,N_1388,N_3961);
nand U17146 (N_17146,N_4259,N_7207);
nor U17147 (N_17147,N_1849,N_1834);
and U17148 (N_17148,N_4401,N_8562);
or U17149 (N_17149,N_7804,N_8486);
and U17150 (N_17150,N_5112,N_3832);
or U17151 (N_17151,N_1587,N_7210);
xor U17152 (N_17152,N_8536,N_8524);
nor U17153 (N_17153,N_3171,N_6735);
nor U17154 (N_17154,N_8288,N_1271);
or U17155 (N_17155,N_1298,N_158);
or U17156 (N_17156,N_9089,N_3826);
nand U17157 (N_17157,N_9039,N_6899);
xnor U17158 (N_17158,N_2751,N_2044);
nor U17159 (N_17159,N_1152,N_6072);
or U17160 (N_17160,N_2765,N_6481);
nand U17161 (N_17161,N_1880,N_2708);
and U17162 (N_17162,N_5062,N_3771);
nand U17163 (N_17163,N_9713,N_7524);
xor U17164 (N_17164,N_5767,N_6052);
or U17165 (N_17165,N_1165,N_5714);
nor U17166 (N_17166,N_6914,N_3873);
or U17167 (N_17167,N_8571,N_3344);
nor U17168 (N_17168,N_1756,N_4541);
nand U17169 (N_17169,N_4123,N_7067);
nor U17170 (N_17170,N_475,N_9663);
and U17171 (N_17171,N_8508,N_7886);
nor U17172 (N_17172,N_6660,N_6761);
and U17173 (N_17173,N_9004,N_9475);
or U17174 (N_17174,N_2285,N_5212);
nor U17175 (N_17175,N_9641,N_3831);
nor U17176 (N_17176,N_7094,N_3565);
xnor U17177 (N_17177,N_9751,N_7682);
nand U17178 (N_17178,N_1831,N_4401);
nor U17179 (N_17179,N_9483,N_4480);
xor U17180 (N_17180,N_9655,N_4983);
nand U17181 (N_17181,N_1322,N_9497);
nor U17182 (N_17182,N_7148,N_2405);
xor U17183 (N_17183,N_9524,N_5944);
xnor U17184 (N_17184,N_6410,N_1257);
or U17185 (N_17185,N_6,N_6195);
and U17186 (N_17186,N_8725,N_8461);
nand U17187 (N_17187,N_1964,N_7994);
nand U17188 (N_17188,N_6300,N_1359);
and U17189 (N_17189,N_3664,N_5691);
nand U17190 (N_17190,N_3581,N_4262);
xnor U17191 (N_17191,N_3348,N_4481);
or U17192 (N_17192,N_5118,N_7954);
and U17193 (N_17193,N_9532,N_6000);
and U17194 (N_17194,N_1109,N_5828);
and U17195 (N_17195,N_8872,N_4664);
or U17196 (N_17196,N_5475,N_7911);
and U17197 (N_17197,N_4079,N_6933);
xor U17198 (N_17198,N_1770,N_3785);
xnor U17199 (N_17199,N_5843,N_1036);
or U17200 (N_17200,N_6111,N_7139);
nor U17201 (N_17201,N_4382,N_537);
nand U17202 (N_17202,N_5586,N_4322);
xnor U17203 (N_17203,N_9928,N_4731);
and U17204 (N_17204,N_9546,N_6925);
nand U17205 (N_17205,N_5177,N_5965);
nor U17206 (N_17206,N_7987,N_1192);
nor U17207 (N_17207,N_2390,N_7617);
nor U17208 (N_17208,N_8370,N_4954);
nand U17209 (N_17209,N_8012,N_3221);
nor U17210 (N_17210,N_7808,N_2823);
or U17211 (N_17211,N_2610,N_362);
and U17212 (N_17212,N_4652,N_2470);
nor U17213 (N_17213,N_8530,N_6608);
nand U17214 (N_17214,N_2775,N_7026);
nor U17215 (N_17215,N_3811,N_4982);
nor U17216 (N_17216,N_2924,N_2727);
and U17217 (N_17217,N_2873,N_4119);
xnor U17218 (N_17218,N_3236,N_7505);
xnor U17219 (N_17219,N_8400,N_776);
or U17220 (N_17220,N_7198,N_5609);
or U17221 (N_17221,N_899,N_8597);
and U17222 (N_17222,N_1433,N_2590);
or U17223 (N_17223,N_9253,N_186);
and U17224 (N_17224,N_8761,N_4779);
and U17225 (N_17225,N_5412,N_7409);
or U17226 (N_17226,N_8894,N_2273);
or U17227 (N_17227,N_1147,N_3787);
and U17228 (N_17228,N_9063,N_5920);
and U17229 (N_17229,N_9252,N_104);
nand U17230 (N_17230,N_6931,N_4769);
nor U17231 (N_17231,N_1798,N_6379);
xnor U17232 (N_17232,N_4021,N_5540);
or U17233 (N_17233,N_5645,N_4048);
nand U17234 (N_17234,N_928,N_7264);
xnor U17235 (N_17235,N_5282,N_2503);
nand U17236 (N_17236,N_5937,N_8622);
nand U17237 (N_17237,N_5382,N_4885);
or U17238 (N_17238,N_3865,N_1436);
nor U17239 (N_17239,N_6794,N_9720);
xor U17240 (N_17240,N_2885,N_6128);
nand U17241 (N_17241,N_701,N_6514);
and U17242 (N_17242,N_788,N_7039);
or U17243 (N_17243,N_8872,N_183);
or U17244 (N_17244,N_1192,N_7365);
nor U17245 (N_17245,N_3351,N_8713);
xor U17246 (N_17246,N_3335,N_4405);
or U17247 (N_17247,N_168,N_1994);
and U17248 (N_17248,N_8793,N_7460);
nor U17249 (N_17249,N_7906,N_2055);
and U17250 (N_17250,N_159,N_8170);
and U17251 (N_17251,N_9029,N_6677);
and U17252 (N_17252,N_1705,N_3254);
nand U17253 (N_17253,N_4969,N_8107);
or U17254 (N_17254,N_6275,N_5509);
nand U17255 (N_17255,N_7818,N_7991);
xnor U17256 (N_17256,N_2609,N_6137);
xnor U17257 (N_17257,N_9355,N_8621);
and U17258 (N_17258,N_9616,N_9873);
nand U17259 (N_17259,N_2461,N_6642);
xnor U17260 (N_17260,N_5126,N_4091);
or U17261 (N_17261,N_9481,N_6395);
nor U17262 (N_17262,N_7019,N_9585);
or U17263 (N_17263,N_238,N_2203);
nor U17264 (N_17264,N_361,N_2361);
or U17265 (N_17265,N_1798,N_2030);
and U17266 (N_17266,N_25,N_2521);
nand U17267 (N_17267,N_2548,N_9503);
or U17268 (N_17268,N_4403,N_8572);
nor U17269 (N_17269,N_4009,N_6832);
nand U17270 (N_17270,N_4362,N_7321);
nor U17271 (N_17271,N_4226,N_7898);
xnor U17272 (N_17272,N_3290,N_6890);
xnor U17273 (N_17273,N_2760,N_7071);
xor U17274 (N_17274,N_633,N_1329);
nor U17275 (N_17275,N_4957,N_2791);
xor U17276 (N_17276,N_739,N_6084);
and U17277 (N_17277,N_3391,N_9687);
xor U17278 (N_17278,N_5082,N_818);
nor U17279 (N_17279,N_7730,N_7638);
or U17280 (N_17280,N_2058,N_2030);
nand U17281 (N_17281,N_1509,N_8467);
nor U17282 (N_17282,N_7851,N_5391);
nor U17283 (N_17283,N_2184,N_6624);
nor U17284 (N_17284,N_2806,N_9263);
or U17285 (N_17285,N_8607,N_2896);
nor U17286 (N_17286,N_1074,N_7527);
or U17287 (N_17287,N_6296,N_7146);
and U17288 (N_17288,N_8704,N_8737);
nand U17289 (N_17289,N_1432,N_9144);
or U17290 (N_17290,N_2290,N_7741);
nor U17291 (N_17291,N_4365,N_6988);
nor U17292 (N_17292,N_6765,N_5361);
or U17293 (N_17293,N_308,N_6672);
nand U17294 (N_17294,N_2912,N_529);
nand U17295 (N_17295,N_5169,N_8119);
and U17296 (N_17296,N_5730,N_5153);
or U17297 (N_17297,N_1101,N_1662);
nand U17298 (N_17298,N_3620,N_7610);
nor U17299 (N_17299,N_786,N_310);
nand U17300 (N_17300,N_333,N_3168);
and U17301 (N_17301,N_6660,N_1468);
and U17302 (N_17302,N_6278,N_7634);
nand U17303 (N_17303,N_8233,N_8903);
or U17304 (N_17304,N_5457,N_6404);
nand U17305 (N_17305,N_3870,N_4938);
xnor U17306 (N_17306,N_3788,N_8161);
or U17307 (N_17307,N_8949,N_3090);
or U17308 (N_17308,N_1077,N_9174);
or U17309 (N_17309,N_8644,N_799);
nand U17310 (N_17310,N_3347,N_5994);
or U17311 (N_17311,N_7647,N_555);
nor U17312 (N_17312,N_6096,N_1508);
and U17313 (N_17313,N_148,N_9114);
and U17314 (N_17314,N_4469,N_4654);
nor U17315 (N_17315,N_8964,N_3953);
and U17316 (N_17316,N_714,N_8886);
or U17317 (N_17317,N_1910,N_4032);
nor U17318 (N_17318,N_8365,N_4071);
nand U17319 (N_17319,N_3010,N_3413);
nor U17320 (N_17320,N_7646,N_7540);
xnor U17321 (N_17321,N_2961,N_4022);
or U17322 (N_17322,N_1420,N_8612);
xor U17323 (N_17323,N_1408,N_3725);
or U17324 (N_17324,N_1071,N_4567);
nand U17325 (N_17325,N_1744,N_3964);
xnor U17326 (N_17326,N_6113,N_7042);
or U17327 (N_17327,N_3148,N_2037);
and U17328 (N_17328,N_5339,N_3891);
xnor U17329 (N_17329,N_1611,N_4922);
nor U17330 (N_17330,N_9394,N_2660);
nor U17331 (N_17331,N_2292,N_9938);
nor U17332 (N_17332,N_661,N_6370);
nor U17333 (N_17333,N_7078,N_589);
nand U17334 (N_17334,N_9734,N_3216);
or U17335 (N_17335,N_3398,N_1126);
nand U17336 (N_17336,N_6593,N_8380);
or U17337 (N_17337,N_6075,N_463);
or U17338 (N_17338,N_256,N_3497);
or U17339 (N_17339,N_5054,N_5696);
and U17340 (N_17340,N_2871,N_5917);
nand U17341 (N_17341,N_2309,N_7544);
nor U17342 (N_17342,N_9093,N_420);
and U17343 (N_17343,N_2397,N_9838);
xnor U17344 (N_17344,N_7483,N_8942);
or U17345 (N_17345,N_7190,N_1576);
nor U17346 (N_17346,N_4597,N_891);
nand U17347 (N_17347,N_8808,N_4707);
nand U17348 (N_17348,N_6500,N_5720);
xor U17349 (N_17349,N_6651,N_2061);
and U17350 (N_17350,N_5578,N_8468);
nor U17351 (N_17351,N_9528,N_6860);
xor U17352 (N_17352,N_9425,N_9567);
and U17353 (N_17353,N_8061,N_8945);
and U17354 (N_17354,N_179,N_2949);
or U17355 (N_17355,N_910,N_5577);
nor U17356 (N_17356,N_3616,N_6970);
or U17357 (N_17357,N_8092,N_4951);
nor U17358 (N_17358,N_4544,N_3395);
nand U17359 (N_17359,N_5664,N_6001);
nand U17360 (N_17360,N_579,N_7126);
and U17361 (N_17361,N_9547,N_1465);
nor U17362 (N_17362,N_6195,N_2491);
and U17363 (N_17363,N_4406,N_7184);
and U17364 (N_17364,N_7751,N_6110);
nor U17365 (N_17365,N_9295,N_8810);
nor U17366 (N_17366,N_6510,N_6713);
and U17367 (N_17367,N_6725,N_6351);
nand U17368 (N_17368,N_4940,N_3433);
xor U17369 (N_17369,N_3028,N_70);
xnor U17370 (N_17370,N_1255,N_8740);
nor U17371 (N_17371,N_7781,N_206);
nand U17372 (N_17372,N_8068,N_4411);
and U17373 (N_17373,N_4465,N_2815);
xor U17374 (N_17374,N_3854,N_2197);
xnor U17375 (N_17375,N_1490,N_7721);
or U17376 (N_17376,N_9390,N_8835);
and U17377 (N_17377,N_6761,N_183);
nand U17378 (N_17378,N_6031,N_3725);
xor U17379 (N_17379,N_3075,N_4186);
nor U17380 (N_17380,N_654,N_8321);
or U17381 (N_17381,N_6761,N_4311);
or U17382 (N_17382,N_3050,N_6554);
nor U17383 (N_17383,N_5291,N_3315);
or U17384 (N_17384,N_4794,N_6613);
nand U17385 (N_17385,N_2488,N_3532);
nor U17386 (N_17386,N_9483,N_7197);
xnor U17387 (N_17387,N_5644,N_8521);
nor U17388 (N_17388,N_981,N_8576);
and U17389 (N_17389,N_9404,N_2424);
nor U17390 (N_17390,N_5766,N_4068);
or U17391 (N_17391,N_3712,N_6003);
or U17392 (N_17392,N_3885,N_7917);
xor U17393 (N_17393,N_5223,N_6246);
or U17394 (N_17394,N_6794,N_8440);
and U17395 (N_17395,N_1176,N_2952);
nand U17396 (N_17396,N_2813,N_4631);
xor U17397 (N_17397,N_1485,N_129);
nand U17398 (N_17398,N_1050,N_4665);
xor U17399 (N_17399,N_1372,N_9646);
or U17400 (N_17400,N_2121,N_9640);
nor U17401 (N_17401,N_499,N_6901);
xnor U17402 (N_17402,N_1652,N_5784);
and U17403 (N_17403,N_9318,N_6253);
nor U17404 (N_17404,N_2431,N_6146);
nand U17405 (N_17405,N_1721,N_9549);
nand U17406 (N_17406,N_6314,N_4890);
nand U17407 (N_17407,N_8097,N_3782);
or U17408 (N_17408,N_8133,N_8643);
and U17409 (N_17409,N_3235,N_8435);
and U17410 (N_17410,N_9998,N_6317);
and U17411 (N_17411,N_7307,N_5401);
nor U17412 (N_17412,N_424,N_896);
nand U17413 (N_17413,N_1571,N_5156);
and U17414 (N_17414,N_4495,N_63);
nor U17415 (N_17415,N_4881,N_9724);
or U17416 (N_17416,N_8132,N_87);
nand U17417 (N_17417,N_1349,N_9226);
nor U17418 (N_17418,N_8361,N_7271);
and U17419 (N_17419,N_1208,N_9050);
nand U17420 (N_17420,N_3716,N_7978);
or U17421 (N_17421,N_72,N_1864);
nand U17422 (N_17422,N_9650,N_8971);
nor U17423 (N_17423,N_5415,N_8390);
nand U17424 (N_17424,N_2990,N_1987);
or U17425 (N_17425,N_5172,N_2203);
xnor U17426 (N_17426,N_3180,N_2146);
xor U17427 (N_17427,N_6820,N_9328);
nor U17428 (N_17428,N_1908,N_7061);
nand U17429 (N_17429,N_719,N_8543);
and U17430 (N_17430,N_727,N_6406);
nor U17431 (N_17431,N_4643,N_4224);
nand U17432 (N_17432,N_7625,N_5661);
xnor U17433 (N_17433,N_3392,N_3693);
and U17434 (N_17434,N_1622,N_7472);
xnor U17435 (N_17435,N_2033,N_2612);
nand U17436 (N_17436,N_453,N_120);
or U17437 (N_17437,N_9510,N_9790);
xor U17438 (N_17438,N_6871,N_1539);
xnor U17439 (N_17439,N_4364,N_6180);
xnor U17440 (N_17440,N_5684,N_8241);
nor U17441 (N_17441,N_4321,N_6231);
nor U17442 (N_17442,N_1852,N_4457);
and U17443 (N_17443,N_3120,N_5132);
xnor U17444 (N_17444,N_4734,N_1618);
or U17445 (N_17445,N_6036,N_9606);
nand U17446 (N_17446,N_5598,N_3529);
nor U17447 (N_17447,N_3054,N_4974);
or U17448 (N_17448,N_7883,N_5104);
or U17449 (N_17449,N_8400,N_9099);
and U17450 (N_17450,N_2182,N_6996);
nand U17451 (N_17451,N_8449,N_4078);
and U17452 (N_17452,N_5229,N_9459);
xor U17453 (N_17453,N_9693,N_7750);
and U17454 (N_17454,N_1887,N_8152);
xor U17455 (N_17455,N_4346,N_2277);
nor U17456 (N_17456,N_5045,N_3971);
xnor U17457 (N_17457,N_7673,N_7074);
or U17458 (N_17458,N_6661,N_9996);
xor U17459 (N_17459,N_1415,N_2036);
xnor U17460 (N_17460,N_8082,N_6985);
nor U17461 (N_17461,N_4529,N_5960);
nand U17462 (N_17462,N_451,N_9660);
nor U17463 (N_17463,N_1852,N_3160);
or U17464 (N_17464,N_5561,N_5300);
and U17465 (N_17465,N_5785,N_1069);
xor U17466 (N_17466,N_2542,N_9967);
and U17467 (N_17467,N_3045,N_7110);
or U17468 (N_17468,N_5711,N_7936);
xnor U17469 (N_17469,N_8175,N_5580);
nand U17470 (N_17470,N_8381,N_1134);
or U17471 (N_17471,N_4715,N_4713);
nand U17472 (N_17472,N_2853,N_2826);
nor U17473 (N_17473,N_5819,N_6402);
nor U17474 (N_17474,N_19,N_783);
xor U17475 (N_17475,N_4217,N_5599);
xor U17476 (N_17476,N_4471,N_8190);
and U17477 (N_17477,N_4260,N_4964);
and U17478 (N_17478,N_5211,N_3455);
nor U17479 (N_17479,N_1810,N_7771);
xnor U17480 (N_17480,N_6878,N_9739);
nor U17481 (N_17481,N_1225,N_9654);
xnor U17482 (N_17482,N_6774,N_2029);
and U17483 (N_17483,N_7033,N_71);
xor U17484 (N_17484,N_8322,N_889);
and U17485 (N_17485,N_7417,N_1195);
nand U17486 (N_17486,N_3874,N_9396);
or U17487 (N_17487,N_823,N_7887);
or U17488 (N_17488,N_3763,N_5809);
nand U17489 (N_17489,N_2012,N_6399);
xor U17490 (N_17490,N_4035,N_4529);
xnor U17491 (N_17491,N_3645,N_951);
and U17492 (N_17492,N_6196,N_9269);
xnor U17493 (N_17493,N_9973,N_7151);
xnor U17494 (N_17494,N_587,N_1966);
xnor U17495 (N_17495,N_1372,N_8722);
nor U17496 (N_17496,N_7592,N_4980);
xor U17497 (N_17497,N_6615,N_3787);
nand U17498 (N_17498,N_2456,N_6321);
and U17499 (N_17499,N_8806,N_9418);
nor U17500 (N_17500,N_2544,N_9173);
nand U17501 (N_17501,N_1036,N_744);
nand U17502 (N_17502,N_5062,N_1150);
xnor U17503 (N_17503,N_1216,N_5201);
nand U17504 (N_17504,N_3566,N_9213);
nand U17505 (N_17505,N_847,N_8895);
or U17506 (N_17506,N_7494,N_2662);
nand U17507 (N_17507,N_4812,N_726);
nand U17508 (N_17508,N_502,N_1670);
nand U17509 (N_17509,N_5616,N_1291);
nor U17510 (N_17510,N_8114,N_4381);
or U17511 (N_17511,N_7578,N_8674);
nor U17512 (N_17512,N_2259,N_4742);
nor U17513 (N_17513,N_1975,N_1304);
xnor U17514 (N_17514,N_927,N_78);
xor U17515 (N_17515,N_7509,N_1373);
xor U17516 (N_17516,N_41,N_5489);
or U17517 (N_17517,N_2253,N_6086);
or U17518 (N_17518,N_1830,N_4687);
nor U17519 (N_17519,N_882,N_9600);
nor U17520 (N_17520,N_9126,N_2629);
and U17521 (N_17521,N_4313,N_2072);
and U17522 (N_17522,N_5687,N_4637);
and U17523 (N_17523,N_672,N_276);
nor U17524 (N_17524,N_2845,N_9709);
and U17525 (N_17525,N_9558,N_4205);
nand U17526 (N_17526,N_6772,N_6617);
and U17527 (N_17527,N_5592,N_2292);
nor U17528 (N_17528,N_7860,N_9817);
or U17529 (N_17529,N_2862,N_6105);
and U17530 (N_17530,N_1931,N_6609);
nand U17531 (N_17531,N_7216,N_823);
or U17532 (N_17532,N_8256,N_2598);
or U17533 (N_17533,N_5019,N_4290);
nand U17534 (N_17534,N_238,N_8080);
nand U17535 (N_17535,N_1072,N_1550);
nand U17536 (N_17536,N_4953,N_5691);
nor U17537 (N_17537,N_3822,N_6054);
or U17538 (N_17538,N_2876,N_457);
or U17539 (N_17539,N_1154,N_8349);
nand U17540 (N_17540,N_2236,N_8149);
or U17541 (N_17541,N_8795,N_5166);
xor U17542 (N_17542,N_9062,N_9824);
nor U17543 (N_17543,N_4602,N_3852);
and U17544 (N_17544,N_1062,N_5061);
nand U17545 (N_17545,N_8504,N_1902);
xnor U17546 (N_17546,N_2488,N_1192);
xnor U17547 (N_17547,N_462,N_7024);
nor U17548 (N_17548,N_1793,N_5254);
and U17549 (N_17549,N_5834,N_7807);
xnor U17550 (N_17550,N_5520,N_8840);
xor U17551 (N_17551,N_6208,N_2452);
nand U17552 (N_17552,N_5517,N_3675);
and U17553 (N_17553,N_8545,N_5864);
nand U17554 (N_17554,N_8253,N_649);
and U17555 (N_17555,N_2433,N_5872);
nor U17556 (N_17556,N_4968,N_4881);
and U17557 (N_17557,N_6540,N_3785);
and U17558 (N_17558,N_5312,N_9017);
nor U17559 (N_17559,N_4398,N_3711);
xnor U17560 (N_17560,N_7709,N_2568);
nand U17561 (N_17561,N_5072,N_1471);
nand U17562 (N_17562,N_1020,N_8875);
nand U17563 (N_17563,N_2558,N_4024);
or U17564 (N_17564,N_9835,N_6535);
or U17565 (N_17565,N_5278,N_4865);
xor U17566 (N_17566,N_34,N_401);
nand U17567 (N_17567,N_5598,N_7969);
nand U17568 (N_17568,N_4031,N_665);
nor U17569 (N_17569,N_4981,N_6853);
nand U17570 (N_17570,N_5295,N_3287);
xor U17571 (N_17571,N_9659,N_7782);
and U17572 (N_17572,N_138,N_4901);
nand U17573 (N_17573,N_4198,N_7500);
or U17574 (N_17574,N_6745,N_2291);
nand U17575 (N_17575,N_9563,N_3286);
xnor U17576 (N_17576,N_7290,N_6653);
nand U17577 (N_17577,N_4912,N_2702);
xor U17578 (N_17578,N_8892,N_7399);
nand U17579 (N_17579,N_6587,N_6209);
or U17580 (N_17580,N_1999,N_95);
and U17581 (N_17581,N_6134,N_8423);
and U17582 (N_17582,N_9325,N_7486);
nor U17583 (N_17583,N_8839,N_1240);
nor U17584 (N_17584,N_2182,N_5880);
nor U17585 (N_17585,N_4101,N_7867);
or U17586 (N_17586,N_3449,N_4154);
or U17587 (N_17587,N_225,N_4334);
and U17588 (N_17588,N_3289,N_2116);
xor U17589 (N_17589,N_8426,N_6690);
or U17590 (N_17590,N_5960,N_1364);
nand U17591 (N_17591,N_1081,N_1091);
and U17592 (N_17592,N_8354,N_5971);
xnor U17593 (N_17593,N_4322,N_3962);
nor U17594 (N_17594,N_3681,N_7426);
nor U17595 (N_17595,N_3334,N_6709);
nor U17596 (N_17596,N_1194,N_4931);
and U17597 (N_17597,N_4848,N_2584);
xnor U17598 (N_17598,N_8922,N_2855);
nor U17599 (N_17599,N_839,N_2525);
nor U17600 (N_17600,N_6413,N_8519);
or U17601 (N_17601,N_5965,N_1958);
or U17602 (N_17602,N_8137,N_8088);
nor U17603 (N_17603,N_9920,N_1277);
nor U17604 (N_17604,N_8410,N_3068);
nor U17605 (N_17605,N_4922,N_9375);
or U17606 (N_17606,N_3304,N_6814);
or U17607 (N_17607,N_7885,N_7348);
nor U17608 (N_17608,N_2557,N_2341);
nand U17609 (N_17609,N_3636,N_4880);
xnor U17610 (N_17610,N_5338,N_512);
nor U17611 (N_17611,N_9814,N_3717);
nor U17612 (N_17612,N_7281,N_9367);
nor U17613 (N_17613,N_2794,N_9170);
or U17614 (N_17614,N_2594,N_8996);
nand U17615 (N_17615,N_8428,N_252);
nand U17616 (N_17616,N_5692,N_2870);
and U17617 (N_17617,N_548,N_5249);
and U17618 (N_17618,N_1103,N_1726);
or U17619 (N_17619,N_9697,N_8258);
or U17620 (N_17620,N_7156,N_8848);
xnor U17621 (N_17621,N_592,N_5360);
xor U17622 (N_17622,N_3787,N_6424);
nor U17623 (N_17623,N_8749,N_3394);
xnor U17624 (N_17624,N_2645,N_8915);
and U17625 (N_17625,N_7206,N_4022);
xnor U17626 (N_17626,N_5766,N_7943);
xnor U17627 (N_17627,N_6137,N_9180);
and U17628 (N_17628,N_2084,N_8503);
nand U17629 (N_17629,N_1797,N_1388);
nand U17630 (N_17630,N_6524,N_1812);
nor U17631 (N_17631,N_9987,N_8025);
nand U17632 (N_17632,N_9937,N_3812);
xor U17633 (N_17633,N_8162,N_4886);
xnor U17634 (N_17634,N_6144,N_9474);
xor U17635 (N_17635,N_2156,N_3457);
and U17636 (N_17636,N_9296,N_4547);
nor U17637 (N_17637,N_7628,N_9736);
xor U17638 (N_17638,N_5629,N_3539);
or U17639 (N_17639,N_4668,N_7391);
nand U17640 (N_17640,N_3175,N_940);
nor U17641 (N_17641,N_5186,N_7320);
xnor U17642 (N_17642,N_6745,N_880);
xor U17643 (N_17643,N_16,N_2187);
or U17644 (N_17644,N_4064,N_667);
xnor U17645 (N_17645,N_1090,N_2178);
and U17646 (N_17646,N_24,N_2487);
nor U17647 (N_17647,N_25,N_5230);
and U17648 (N_17648,N_5688,N_8403);
or U17649 (N_17649,N_1322,N_8866);
nor U17650 (N_17650,N_6951,N_9919);
and U17651 (N_17651,N_6008,N_1912);
nor U17652 (N_17652,N_6215,N_6556);
nand U17653 (N_17653,N_2146,N_881);
and U17654 (N_17654,N_7107,N_6511);
nand U17655 (N_17655,N_5779,N_501);
nor U17656 (N_17656,N_8145,N_8399);
and U17657 (N_17657,N_3842,N_533);
xor U17658 (N_17658,N_8382,N_7872);
and U17659 (N_17659,N_250,N_3773);
nor U17660 (N_17660,N_9063,N_7187);
or U17661 (N_17661,N_186,N_4548);
and U17662 (N_17662,N_5811,N_4295);
xor U17663 (N_17663,N_5473,N_4670);
nand U17664 (N_17664,N_5043,N_3415);
xnor U17665 (N_17665,N_3185,N_7912);
xor U17666 (N_17666,N_6708,N_8850);
xnor U17667 (N_17667,N_8291,N_6266);
nand U17668 (N_17668,N_4283,N_4756);
or U17669 (N_17669,N_3794,N_5262);
nand U17670 (N_17670,N_8505,N_5589);
and U17671 (N_17671,N_1595,N_5963);
nor U17672 (N_17672,N_821,N_8544);
or U17673 (N_17673,N_4945,N_8752);
and U17674 (N_17674,N_7122,N_9086);
or U17675 (N_17675,N_3924,N_3159);
and U17676 (N_17676,N_7936,N_1102);
xor U17677 (N_17677,N_4757,N_6344);
or U17678 (N_17678,N_3896,N_1338);
nand U17679 (N_17679,N_8452,N_7);
xor U17680 (N_17680,N_4442,N_1987);
nand U17681 (N_17681,N_9451,N_5961);
nor U17682 (N_17682,N_4188,N_1972);
and U17683 (N_17683,N_2792,N_2639);
and U17684 (N_17684,N_8920,N_7136);
nor U17685 (N_17685,N_6159,N_1836);
xor U17686 (N_17686,N_2226,N_3383);
or U17687 (N_17687,N_5723,N_3231);
and U17688 (N_17688,N_482,N_8440);
or U17689 (N_17689,N_1746,N_7689);
nand U17690 (N_17690,N_3356,N_7960);
or U17691 (N_17691,N_5530,N_1044);
nor U17692 (N_17692,N_7969,N_2638);
nand U17693 (N_17693,N_261,N_4186);
nor U17694 (N_17694,N_4690,N_5305);
nand U17695 (N_17695,N_6185,N_2020);
and U17696 (N_17696,N_979,N_2448);
or U17697 (N_17697,N_5425,N_8885);
nor U17698 (N_17698,N_8997,N_3286);
and U17699 (N_17699,N_4892,N_3910);
nor U17700 (N_17700,N_8161,N_9299);
nand U17701 (N_17701,N_3391,N_3181);
and U17702 (N_17702,N_4283,N_1045);
or U17703 (N_17703,N_1477,N_5509);
and U17704 (N_17704,N_5408,N_4552);
nand U17705 (N_17705,N_1459,N_3190);
xnor U17706 (N_17706,N_7228,N_3329);
nor U17707 (N_17707,N_8358,N_4267);
xnor U17708 (N_17708,N_2534,N_3769);
or U17709 (N_17709,N_2616,N_2435);
or U17710 (N_17710,N_301,N_7323);
nor U17711 (N_17711,N_746,N_6384);
nand U17712 (N_17712,N_2713,N_8391);
or U17713 (N_17713,N_500,N_6226);
nor U17714 (N_17714,N_7735,N_916);
nand U17715 (N_17715,N_7223,N_3059);
nor U17716 (N_17716,N_828,N_3319);
nand U17717 (N_17717,N_1978,N_1077);
nor U17718 (N_17718,N_9129,N_6661);
and U17719 (N_17719,N_4865,N_5490);
xnor U17720 (N_17720,N_9516,N_1401);
nand U17721 (N_17721,N_6526,N_7372);
and U17722 (N_17722,N_3871,N_6769);
nor U17723 (N_17723,N_8628,N_4214);
and U17724 (N_17724,N_5754,N_8384);
nand U17725 (N_17725,N_8561,N_3528);
or U17726 (N_17726,N_4241,N_2427);
and U17727 (N_17727,N_7830,N_5522);
nand U17728 (N_17728,N_4269,N_9268);
nand U17729 (N_17729,N_6933,N_6807);
or U17730 (N_17730,N_5018,N_6381);
or U17731 (N_17731,N_1423,N_2609);
nor U17732 (N_17732,N_3117,N_6118);
or U17733 (N_17733,N_6327,N_8505);
nor U17734 (N_17734,N_9426,N_8077);
xor U17735 (N_17735,N_9232,N_5917);
and U17736 (N_17736,N_9701,N_2831);
xor U17737 (N_17737,N_5952,N_8358);
nand U17738 (N_17738,N_9725,N_3683);
or U17739 (N_17739,N_6028,N_7025);
nor U17740 (N_17740,N_3333,N_7271);
nor U17741 (N_17741,N_3896,N_4604);
and U17742 (N_17742,N_5775,N_2546);
or U17743 (N_17743,N_3192,N_1150);
xnor U17744 (N_17744,N_4352,N_3570);
xor U17745 (N_17745,N_9381,N_593);
and U17746 (N_17746,N_1510,N_4343);
nor U17747 (N_17747,N_5364,N_3959);
nand U17748 (N_17748,N_6145,N_8873);
and U17749 (N_17749,N_4503,N_4026);
and U17750 (N_17750,N_4564,N_9127);
xnor U17751 (N_17751,N_4901,N_6049);
nor U17752 (N_17752,N_1953,N_5393);
or U17753 (N_17753,N_134,N_1311);
nand U17754 (N_17754,N_51,N_9202);
or U17755 (N_17755,N_9403,N_9466);
or U17756 (N_17756,N_3962,N_9237);
nand U17757 (N_17757,N_439,N_741);
and U17758 (N_17758,N_4083,N_7796);
nand U17759 (N_17759,N_6603,N_2483);
and U17760 (N_17760,N_8564,N_4522);
xnor U17761 (N_17761,N_8196,N_5820);
xnor U17762 (N_17762,N_6637,N_6221);
or U17763 (N_17763,N_3908,N_213);
xor U17764 (N_17764,N_5656,N_6438);
and U17765 (N_17765,N_3138,N_2573);
nor U17766 (N_17766,N_4806,N_1707);
xnor U17767 (N_17767,N_6530,N_3978);
xor U17768 (N_17768,N_9010,N_58);
nand U17769 (N_17769,N_7562,N_9515);
nor U17770 (N_17770,N_3019,N_2011);
xnor U17771 (N_17771,N_9744,N_4608);
xor U17772 (N_17772,N_7740,N_9383);
xor U17773 (N_17773,N_9873,N_8511);
and U17774 (N_17774,N_3007,N_5075);
nand U17775 (N_17775,N_1502,N_7190);
nand U17776 (N_17776,N_812,N_4218);
nand U17777 (N_17777,N_3039,N_51);
xor U17778 (N_17778,N_1095,N_6324);
xnor U17779 (N_17779,N_8870,N_1853);
and U17780 (N_17780,N_2011,N_5034);
xor U17781 (N_17781,N_1461,N_5663);
and U17782 (N_17782,N_5150,N_8973);
and U17783 (N_17783,N_8060,N_6495);
xor U17784 (N_17784,N_3843,N_7346);
xnor U17785 (N_17785,N_3035,N_7598);
nand U17786 (N_17786,N_7490,N_5116);
nand U17787 (N_17787,N_2685,N_5889);
nand U17788 (N_17788,N_6423,N_2830);
nand U17789 (N_17789,N_6995,N_7655);
xor U17790 (N_17790,N_2430,N_9630);
nor U17791 (N_17791,N_5185,N_8009);
nand U17792 (N_17792,N_8407,N_4844);
and U17793 (N_17793,N_3606,N_4931);
and U17794 (N_17794,N_6394,N_4595);
nand U17795 (N_17795,N_7180,N_6853);
xor U17796 (N_17796,N_5917,N_766);
or U17797 (N_17797,N_6957,N_5325);
and U17798 (N_17798,N_1265,N_5184);
and U17799 (N_17799,N_6632,N_9348);
or U17800 (N_17800,N_145,N_7616);
or U17801 (N_17801,N_2120,N_558);
nor U17802 (N_17802,N_6225,N_2778);
nand U17803 (N_17803,N_7936,N_1004);
or U17804 (N_17804,N_3655,N_4055);
xor U17805 (N_17805,N_1022,N_7663);
and U17806 (N_17806,N_3696,N_9669);
nand U17807 (N_17807,N_3212,N_777);
or U17808 (N_17808,N_8626,N_9431);
and U17809 (N_17809,N_8045,N_7161);
nand U17810 (N_17810,N_5920,N_5870);
nor U17811 (N_17811,N_3602,N_2828);
or U17812 (N_17812,N_5959,N_7810);
nor U17813 (N_17813,N_6152,N_7211);
or U17814 (N_17814,N_5495,N_7403);
xor U17815 (N_17815,N_5073,N_7891);
or U17816 (N_17816,N_5778,N_3955);
or U17817 (N_17817,N_85,N_8008);
nand U17818 (N_17818,N_394,N_9719);
nor U17819 (N_17819,N_1839,N_7917);
nor U17820 (N_17820,N_6013,N_745);
xnor U17821 (N_17821,N_5144,N_6314);
xnor U17822 (N_17822,N_2193,N_4121);
nand U17823 (N_17823,N_2918,N_8991);
xor U17824 (N_17824,N_8806,N_2899);
nand U17825 (N_17825,N_4929,N_333);
and U17826 (N_17826,N_4132,N_323);
nor U17827 (N_17827,N_7385,N_4897);
nand U17828 (N_17828,N_7379,N_9425);
or U17829 (N_17829,N_3480,N_3883);
and U17830 (N_17830,N_4250,N_2624);
nand U17831 (N_17831,N_6424,N_8934);
nor U17832 (N_17832,N_9437,N_7484);
and U17833 (N_17833,N_5123,N_8815);
xnor U17834 (N_17834,N_8326,N_7556);
xor U17835 (N_17835,N_5589,N_5582);
or U17836 (N_17836,N_7075,N_8543);
nand U17837 (N_17837,N_729,N_823);
xor U17838 (N_17838,N_886,N_178);
and U17839 (N_17839,N_6196,N_1643);
and U17840 (N_17840,N_4405,N_2265);
nor U17841 (N_17841,N_2352,N_9435);
and U17842 (N_17842,N_8095,N_4107);
nand U17843 (N_17843,N_1567,N_5986);
xnor U17844 (N_17844,N_8959,N_9002);
xor U17845 (N_17845,N_7561,N_2913);
and U17846 (N_17846,N_6532,N_6379);
xor U17847 (N_17847,N_4869,N_7429);
xor U17848 (N_17848,N_6366,N_2969);
xnor U17849 (N_17849,N_7208,N_1604);
nand U17850 (N_17850,N_4551,N_6990);
and U17851 (N_17851,N_5911,N_9225);
nor U17852 (N_17852,N_1386,N_4648);
or U17853 (N_17853,N_3885,N_6260);
and U17854 (N_17854,N_8735,N_4430);
or U17855 (N_17855,N_3165,N_3191);
xnor U17856 (N_17856,N_8311,N_2503);
nor U17857 (N_17857,N_4874,N_6727);
and U17858 (N_17858,N_4189,N_1973);
nor U17859 (N_17859,N_4174,N_8396);
and U17860 (N_17860,N_4217,N_5429);
and U17861 (N_17861,N_3235,N_3916);
or U17862 (N_17862,N_3314,N_7898);
and U17863 (N_17863,N_4329,N_9318);
and U17864 (N_17864,N_9184,N_5249);
xnor U17865 (N_17865,N_2532,N_9768);
and U17866 (N_17866,N_2316,N_4022);
nor U17867 (N_17867,N_1306,N_3670);
or U17868 (N_17868,N_2359,N_3990);
nand U17869 (N_17869,N_329,N_4899);
xor U17870 (N_17870,N_5507,N_2232);
and U17871 (N_17871,N_9162,N_3299);
nand U17872 (N_17872,N_6690,N_7365);
xor U17873 (N_17873,N_1172,N_300);
and U17874 (N_17874,N_8313,N_6753);
nor U17875 (N_17875,N_3829,N_9000);
nand U17876 (N_17876,N_2143,N_7594);
nand U17877 (N_17877,N_1485,N_1978);
or U17878 (N_17878,N_2334,N_9408);
or U17879 (N_17879,N_4878,N_2013);
and U17880 (N_17880,N_7028,N_7687);
xor U17881 (N_17881,N_5964,N_934);
nand U17882 (N_17882,N_8846,N_8005);
nand U17883 (N_17883,N_358,N_4933);
nor U17884 (N_17884,N_4237,N_4790);
nand U17885 (N_17885,N_5165,N_8128);
and U17886 (N_17886,N_9988,N_8636);
or U17887 (N_17887,N_1462,N_2083);
nor U17888 (N_17888,N_7200,N_9556);
or U17889 (N_17889,N_4965,N_6794);
and U17890 (N_17890,N_4254,N_6896);
nand U17891 (N_17891,N_2223,N_4538);
nand U17892 (N_17892,N_9059,N_9510);
nor U17893 (N_17893,N_3049,N_5369);
and U17894 (N_17894,N_6706,N_1714);
xor U17895 (N_17895,N_7058,N_9295);
nor U17896 (N_17896,N_1246,N_7153);
xor U17897 (N_17897,N_4925,N_8203);
nor U17898 (N_17898,N_7795,N_8664);
nand U17899 (N_17899,N_3864,N_564);
nand U17900 (N_17900,N_4281,N_9190);
or U17901 (N_17901,N_2083,N_7614);
and U17902 (N_17902,N_6828,N_7186);
or U17903 (N_17903,N_948,N_6814);
nor U17904 (N_17904,N_5417,N_6366);
nor U17905 (N_17905,N_6130,N_9755);
or U17906 (N_17906,N_4479,N_3194);
nand U17907 (N_17907,N_3376,N_3997);
nand U17908 (N_17908,N_2453,N_9918);
nor U17909 (N_17909,N_2700,N_4159);
and U17910 (N_17910,N_4420,N_7979);
or U17911 (N_17911,N_8419,N_5803);
nor U17912 (N_17912,N_6478,N_9731);
or U17913 (N_17913,N_6857,N_4056);
xor U17914 (N_17914,N_3963,N_4692);
or U17915 (N_17915,N_8601,N_9157);
nand U17916 (N_17916,N_1299,N_8190);
nand U17917 (N_17917,N_4854,N_5845);
or U17918 (N_17918,N_3493,N_1202);
nor U17919 (N_17919,N_8708,N_5931);
nor U17920 (N_17920,N_2920,N_7475);
nand U17921 (N_17921,N_1143,N_1242);
or U17922 (N_17922,N_3712,N_1303);
and U17923 (N_17923,N_5454,N_5397);
and U17924 (N_17924,N_5184,N_4813);
and U17925 (N_17925,N_1116,N_8620);
or U17926 (N_17926,N_3582,N_7796);
and U17927 (N_17927,N_6830,N_3373);
and U17928 (N_17928,N_4520,N_7365);
nand U17929 (N_17929,N_1927,N_2190);
and U17930 (N_17930,N_1762,N_12);
nand U17931 (N_17931,N_5881,N_1957);
nand U17932 (N_17932,N_6788,N_5728);
nand U17933 (N_17933,N_7385,N_9962);
nor U17934 (N_17934,N_8857,N_8979);
or U17935 (N_17935,N_8981,N_5268);
xor U17936 (N_17936,N_7539,N_9254);
xor U17937 (N_17937,N_8827,N_7172);
xor U17938 (N_17938,N_4319,N_8218);
nor U17939 (N_17939,N_4590,N_5094);
xor U17940 (N_17940,N_4602,N_986);
or U17941 (N_17941,N_5135,N_1590);
nor U17942 (N_17942,N_7645,N_6893);
or U17943 (N_17943,N_4454,N_1743);
and U17944 (N_17944,N_8588,N_9942);
nor U17945 (N_17945,N_2280,N_5247);
xor U17946 (N_17946,N_930,N_1941);
or U17947 (N_17947,N_3339,N_2609);
xor U17948 (N_17948,N_4939,N_4798);
and U17949 (N_17949,N_7564,N_8632);
or U17950 (N_17950,N_5289,N_292);
or U17951 (N_17951,N_7992,N_765);
or U17952 (N_17952,N_4893,N_1603);
nand U17953 (N_17953,N_7727,N_6690);
or U17954 (N_17954,N_7116,N_3370);
or U17955 (N_17955,N_878,N_5592);
nor U17956 (N_17956,N_852,N_582);
nand U17957 (N_17957,N_70,N_2496);
nor U17958 (N_17958,N_6549,N_3793);
and U17959 (N_17959,N_5359,N_5170);
nand U17960 (N_17960,N_6152,N_1271);
or U17961 (N_17961,N_8314,N_9198);
nor U17962 (N_17962,N_812,N_106);
xor U17963 (N_17963,N_9716,N_8295);
and U17964 (N_17964,N_8947,N_6746);
and U17965 (N_17965,N_9426,N_5408);
nor U17966 (N_17966,N_5502,N_1469);
nor U17967 (N_17967,N_3223,N_3786);
xnor U17968 (N_17968,N_354,N_1297);
or U17969 (N_17969,N_5493,N_3400);
xnor U17970 (N_17970,N_5667,N_5612);
xor U17971 (N_17971,N_2019,N_6343);
nand U17972 (N_17972,N_4670,N_4235);
and U17973 (N_17973,N_2134,N_4358);
xor U17974 (N_17974,N_5790,N_5706);
nand U17975 (N_17975,N_6089,N_1536);
xor U17976 (N_17976,N_4557,N_5331);
and U17977 (N_17977,N_828,N_7824);
nor U17978 (N_17978,N_9282,N_5111);
and U17979 (N_17979,N_5552,N_1979);
or U17980 (N_17980,N_9691,N_3419);
nand U17981 (N_17981,N_1367,N_4013);
xnor U17982 (N_17982,N_9135,N_2695);
xnor U17983 (N_17983,N_6563,N_9014);
xor U17984 (N_17984,N_4749,N_2883);
nand U17985 (N_17985,N_3360,N_9760);
nand U17986 (N_17986,N_7787,N_6564);
nand U17987 (N_17987,N_6408,N_9898);
nor U17988 (N_17988,N_4564,N_9932);
xnor U17989 (N_17989,N_1253,N_7598);
or U17990 (N_17990,N_7947,N_554);
nor U17991 (N_17991,N_8449,N_1687);
nor U17992 (N_17992,N_88,N_2214);
nand U17993 (N_17993,N_7353,N_9145);
nand U17994 (N_17994,N_3336,N_2283);
and U17995 (N_17995,N_4006,N_3754);
and U17996 (N_17996,N_5546,N_1046);
nand U17997 (N_17997,N_9894,N_3005);
and U17998 (N_17998,N_5858,N_471);
nor U17999 (N_17999,N_5884,N_8509);
nor U18000 (N_18000,N_6288,N_8520);
nand U18001 (N_18001,N_4394,N_6609);
or U18002 (N_18002,N_6700,N_1981);
nor U18003 (N_18003,N_9528,N_6337);
and U18004 (N_18004,N_8096,N_7251);
or U18005 (N_18005,N_5485,N_8737);
nand U18006 (N_18006,N_465,N_5300);
nor U18007 (N_18007,N_4323,N_982);
and U18008 (N_18008,N_8260,N_7008);
and U18009 (N_18009,N_1129,N_8028);
xor U18010 (N_18010,N_4800,N_2678);
and U18011 (N_18011,N_3358,N_9259);
nor U18012 (N_18012,N_4081,N_8633);
or U18013 (N_18013,N_1459,N_5005);
nor U18014 (N_18014,N_9900,N_5456);
and U18015 (N_18015,N_3325,N_2090);
nand U18016 (N_18016,N_8434,N_9365);
and U18017 (N_18017,N_9145,N_7617);
or U18018 (N_18018,N_603,N_4503);
or U18019 (N_18019,N_9912,N_7277);
xnor U18020 (N_18020,N_1882,N_4922);
nor U18021 (N_18021,N_8232,N_787);
or U18022 (N_18022,N_8909,N_8326);
nor U18023 (N_18023,N_2978,N_9965);
and U18024 (N_18024,N_4013,N_7911);
or U18025 (N_18025,N_4205,N_3804);
nor U18026 (N_18026,N_8806,N_2354);
or U18027 (N_18027,N_4122,N_4514);
and U18028 (N_18028,N_4382,N_2248);
and U18029 (N_18029,N_5411,N_4960);
xnor U18030 (N_18030,N_1940,N_4667);
nor U18031 (N_18031,N_8911,N_353);
and U18032 (N_18032,N_919,N_7711);
nand U18033 (N_18033,N_9788,N_3986);
xnor U18034 (N_18034,N_2232,N_1021);
or U18035 (N_18035,N_5067,N_1428);
or U18036 (N_18036,N_8806,N_3765);
and U18037 (N_18037,N_7378,N_9715);
nor U18038 (N_18038,N_6273,N_3487);
or U18039 (N_18039,N_1794,N_839);
nand U18040 (N_18040,N_5118,N_5348);
nor U18041 (N_18041,N_2003,N_3164);
nor U18042 (N_18042,N_80,N_3690);
or U18043 (N_18043,N_7198,N_3864);
nor U18044 (N_18044,N_2665,N_9838);
nand U18045 (N_18045,N_9958,N_1324);
nand U18046 (N_18046,N_6962,N_7709);
or U18047 (N_18047,N_4689,N_5929);
or U18048 (N_18048,N_4322,N_2034);
nor U18049 (N_18049,N_5305,N_96);
or U18050 (N_18050,N_6983,N_618);
xnor U18051 (N_18051,N_9549,N_6288);
nand U18052 (N_18052,N_749,N_5707);
or U18053 (N_18053,N_4604,N_6759);
and U18054 (N_18054,N_8853,N_2637);
nand U18055 (N_18055,N_6740,N_7985);
nand U18056 (N_18056,N_1921,N_5771);
xor U18057 (N_18057,N_3135,N_3335);
and U18058 (N_18058,N_5378,N_4597);
or U18059 (N_18059,N_6083,N_5086);
and U18060 (N_18060,N_9822,N_7792);
or U18061 (N_18061,N_9573,N_2905);
nand U18062 (N_18062,N_9309,N_4525);
nor U18063 (N_18063,N_1540,N_9610);
or U18064 (N_18064,N_2075,N_8226);
or U18065 (N_18065,N_928,N_2856);
and U18066 (N_18066,N_8461,N_5036);
nand U18067 (N_18067,N_7733,N_2663);
and U18068 (N_18068,N_7295,N_2317);
nor U18069 (N_18069,N_8652,N_9392);
nand U18070 (N_18070,N_2525,N_6894);
nor U18071 (N_18071,N_2045,N_9114);
nand U18072 (N_18072,N_5697,N_3528);
or U18073 (N_18073,N_6964,N_4985);
nand U18074 (N_18074,N_2731,N_9731);
nor U18075 (N_18075,N_1868,N_7777);
nor U18076 (N_18076,N_840,N_7704);
xnor U18077 (N_18077,N_1633,N_9958);
nand U18078 (N_18078,N_2306,N_9146);
nor U18079 (N_18079,N_8373,N_2361);
or U18080 (N_18080,N_3226,N_331);
xor U18081 (N_18081,N_3518,N_9255);
nand U18082 (N_18082,N_9445,N_2968);
xor U18083 (N_18083,N_6569,N_1411);
nand U18084 (N_18084,N_452,N_2010);
nand U18085 (N_18085,N_5615,N_7959);
nand U18086 (N_18086,N_4986,N_1293);
and U18087 (N_18087,N_2556,N_1037);
nand U18088 (N_18088,N_3595,N_7066);
or U18089 (N_18089,N_1050,N_2197);
or U18090 (N_18090,N_9204,N_2101);
nand U18091 (N_18091,N_7257,N_3863);
or U18092 (N_18092,N_2541,N_8932);
and U18093 (N_18093,N_735,N_8103);
and U18094 (N_18094,N_4658,N_1464);
and U18095 (N_18095,N_5321,N_9155);
and U18096 (N_18096,N_7969,N_8061);
xnor U18097 (N_18097,N_4536,N_5137);
nand U18098 (N_18098,N_6469,N_4741);
nand U18099 (N_18099,N_8485,N_806);
nand U18100 (N_18100,N_1022,N_8824);
xnor U18101 (N_18101,N_1475,N_8589);
and U18102 (N_18102,N_4186,N_5785);
nor U18103 (N_18103,N_2011,N_815);
or U18104 (N_18104,N_4748,N_4613);
nand U18105 (N_18105,N_6278,N_1469);
nor U18106 (N_18106,N_4974,N_4037);
nand U18107 (N_18107,N_890,N_4525);
or U18108 (N_18108,N_1998,N_9896);
nand U18109 (N_18109,N_7188,N_6811);
nand U18110 (N_18110,N_2288,N_2423);
and U18111 (N_18111,N_5542,N_3554);
or U18112 (N_18112,N_7638,N_4458);
nor U18113 (N_18113,N_9906,N_6851);
xor U18114 (N_18114,N_6504,N_8446);
xnor U18115 (N_18115,N_557,N_1991);
or U18116 (N_18116,N_2896,N_2977);
or U18117 (N_18117,N_835,N_3391);
xor U18118 (N_18118,N_524,N_4753);
and U18119 (N_18119,N_2378,N_3550);
and U18120 (N_18120,N_9882,N_8961);
nand U18121 (N_18121,N_9146,N_2966);
and U18122 (N_18122,N_1786,N_8677);
nor U18123 (N_18123,N_3261,N_1816);
or U18124 (N_18124,N_7865,N_5972);
nand U18125 (N_18125,N_3699,N_6712);
or U18126 (N_18126,N_1567,N_1264);
nor U18127 (N_18127,N_4772,N_8070);
xor U18128 (N_18128,N_7556,N_3906);
or U18129 (N_18129,N_1025,N_6482);
and U18130 (N_18130,N_4967,N_732);
or U18131 (N_18131,N_1820,N_5993);
and U18132 (N_18132,N_2315,N_5959);
nand U18133 (N_18133,N_5020,N_772);
nand U18134 (N_18134,N_5285,N_2575);
xnor U18135 (N_18135,N_2182,N_9282);
or U18136 (N_18136,N_1024,N_5914);
xor U18137 (N_18137,N_8292,N_2052);
or U18138 (N_18138,N_6894,N_2274);
nor U18139 (N_18139,N_8777,N_193);
xor U18140 (N_18140,N_6614,N_5734);
xor U18141 (N_18141,N_4519,N_5723);
or U18142 (N_18142,N_8046,N_2555);
xnor U18143 (N_18143,N_402,N_9725);
and U18144 (N_18144,N_1658,N_8613);
xor U18145 (N_18145,N_6695,N_3877);
nor U18146 (N_18146,N_1210,N_9122);
and U18147 (N_18147,N_7466,N_1149);
and U18148 (N_18148,N_5159,N_8565);
nor U18149 (N_18149,N_6002,N_3742);
nor U18150 (N_18150,N_8366,N_6175);
and U18151 (N_18151,N_7502,N_6285);
or U18152 (N_18152,N_5539,N_6122);
xor U18153 (N_18153,N_5632,N_7102);
nor U18154 (N_18154,N_1587,N_7147);
or U18155 (N_18155,N_3334,N_439);
nand U18156 (N_18156,N_908,N_9668);
xor U18157 (N_18157,N_1573,N_3166);
xor U18158 (N_18158,N_6492,N_7955);
xnor U18159 (N_18159,N_3291,N_9444);
nor U18160 (N_18160,N_25,N_3597);
or U18161 (N_18161,N_8501,N_6670);
xnor U18162 (N_18162,N_9330,N_8460);
nor U18163 (N_18163,N_4044,N_6400);
nand U18164 (N_18164,N_1346,N_8919);
and U18165 (N_18165,N_2159,N_9225);
or U18166 (N_18166,N_9524,N_8545);
nand U18167 (N_18167,N_1084,N_3115);
xnor U18168 (N_18168,N_471,N_5054);
nor U18169 (N_18169,N_2480,N_2051);
xnor U18170 (N_18170,N_6450,N_5425);
nor U18171 (N_18171,N_5065,N_5078);
nor U18172 (N_18172,N_4260,N_3874);
nand U18173 (N_18173,N_2805,N_4907);
and U18174 (N_18174,N_83,N_7260);
or U18175 (N_18175,N_4535,N_2917);
and U18176 (N_18176,N_520,N_1664);
nor U18177 (N_18177,N_6138,N_8953);
or U18178 (N_18178,N_3230,N_5672);
and U18179 (N_18179,N_5756,N_5122);
or U18180 (N_18180,N_6968,N_2131);
xnor U18181 (N_18181,N_8824,N_7820);
nand U18182 (N_18182,N_2274,N_9905);
xnor U18183 (N_18183,N_2239,N_8751);
nand U18184 (N_18184,N_9817,N_7415);
nand U18185 (N_18185,N_9722,N_8185);
nor U18186 (N_18186,N_6137,N_2674);
nor U18187 (N_18187,N_3455,N_3004);
or U18188 (N_18188,N_1704,N_3022);
and U18189 (N_18189,N_7234,N_1124);
xnor U18190 (N_18190,N_2700,N_6853);
nor U18191 (N_18191,N_9434,N_6438);
nand U18192 (N_18192,N_7359,N_1530);
and U18193 (N_18193,N_5866,N_5567);
and U18194 (N_18194,N_2851,N_4278);
xnor U18195 (N_18195,N_5464,N_915);
or U18196 (N_18196,N_267,N_86);
and U18197 (N_18197,N_9556,N_1008);
and U18198 (N_18198,N_5153,N_8960);
nor U18199 (N_18199,N_6329,N_1034);
nor U18200 (N_18200,N_9179,N_3477);
or U18201 (N_18201,N_6374,N_7333);
nor U18202 (N_18202,N_1174,N_8410);
and U18203 (N_18203,N_2581,N_2295);
nor U18204 (N_18204,N_2924,N_8701);
xnor U18205 (N_18205,N_9952,N_1061);
or U18206 (N_18206,N_3299,N_5725);
xnor U18207 (N_18207,N_8692,N_5287);
or U18208 (N_18208,N_5911,N_9252);
or U18209 (N_18209,N_1714,N_4415);
nand U18210 (N_18210,N_8765,N_6826);
or U18211 (N_18211,N_7747,N_9670);
nor U18212 (N_18212,N_6060,N_9855);
or U18213 (N_18213,N_4481,N_2437);
nor U18214 (N_18214,N_5853,N_156);
nand U18215 (N_18215,N_525,N_9476);
and U18216 (N_18216,N_9590,N_6673);
nand U18217 (N_18217,N_2174,N_6970);
xor U18218 (N_18218,N_8760,N_7724);
or U18219 (N_18219,N_5385,N_679);
or U18220 (N_18220,N_2323,N_4681);
or U18221 (N_18221,N_3120,N_4760);
nand U18222 (N_18222,N_2677,N_1963);
xor U18223 (N_18223,N_8888,N_3196);
nor U18224 (N_18224,N_3302,N_7116);
and U18225 (N_18225,N_2656,N_6880);
and U18226 (N_18226,N_3128,N_5982);
xor U18227 (N_18227,N_92,N_356);
nand U18228 (N_18228,N_7139,N_4031);
or U18229 (N_18229,N_1941,N_9951);
xor U18230 (N_18230,N_1780,N_1314);
nand U18231 (N_18231,N_9464,N_9667);
or U18232 (N_18232,N_6866,N_948);
or U18233 (N_18233,N_3601,N_3223);
xor U18234 (N_18234,N_9616,N_5209);
nor U18235 (N_18235,N_1135,N_2977);
or U18236 (N_18236,N_715,N_2911);
and U18237 (N_18237,N_3207,N_6336);
or U18238 (N_18238,N_7668,N_2030);
nor U18239 (N_18239,N_7636,N_6570);
nand U18240 (N_18240,N_3170,N_1053);
xnor U18241 (N_18241,N_8031,N_7558);
xnor U18242 (N_18242,N_2363,N_8630);
xnor U18243 (N_18243,N_6593,N_6229);
and U18244 (N_18244,N_8878,N_2995);
nand U18245 (N_18245,N_2198,N_3089);
xor U18246 (N_18246,N_73,N_4664);
and U18247 (N_18247,N_3532,N_9273);
nand U18248 (N_18248,N_9009,N_4220);
and U18249 (N_18249,N_8941,N_7088);
nand U18250 (N_18250,N_5448,N_2792);
or U18251 (N_18251,N_5250,N_549);
nor U18252 (N_18252,N_2409,N_3812);
nand U18253 (N_18253,N_1392,N_7068);
and U18254 (N_18254,N_8832,N_8212);
or U18255 (N_18255,N_1985,N_7709);
or U18256 (N_18256,N_7492,N_7227);
nand U18257 (N_18257,N_1113,N_3640);
or U18258 (N_18258,N_9634,N_3858);
nand U18259 (N_18259,N_9718,N_5196);
or U18260 (N_18260,N_2167,N_9918);
nand U18261 (N_18261,N_1753,N_6567);
and U18262 (N_18262,N_7491,N_8079);
and U18263 (N_18263,N_4867,N_6434);
nor U18264 (N_18264,N_4201,N_5275);
nor U18265 (N_18265,N_1814,N_8986);
or U18266 (N_18266,N_8729,N_3825);
and U18267 (N_18267,N_7209,N_4452);
nand U18268 (N_18268,N_733,N_7220);
and U18269 (N_18269,N_306,N_5088);
xor U18270 (N_18270,N_4857,N_2737);
nand U18271 (N_18271,N_8781,N_4356);
xnor U18272 (N_18272,N_9482,N_1987);
and U18273 (N_18273,N_8427,N_8235);
nor U18274 (N_18274,N_1819,N_1766);
or U18275 (N_18275,N_229,N_698);
nand U18276 (N_18276,N_4664,N_9833);
nand U18277 (N_18277,N_5284,N_9467);
xnor U18278 (N_18278,N_9265,N_6728);
nand U18279 (N_18279,N_9494,N_7461);
or U18280 (N_18280,N_5823,N_7605);
or U18281 (N_18281,N_6666,N_2750);
xnor U18282 (N_18282,N_4288,N_4743);
nor U18283 (N_18283,N_7045,N_494);
nand U18284 (N_18284,N_2356,N_4789);
xnor U18285 (N_18285,N_9090,N_5614);
nor U18286 (N_18286,N_2694,N_1738);
and U18287 (N_18287,N_8047,N_2405);
nand U18288 (N_18288,N_7750,N_6816);
nor U18289 (N_18289,N_4774,N_1953);
xor U18290 (N_18290,N_3643,N_1228);
xor U18291 (N_18291,N_2354,N_9822);
nand U18292 (N_18292,N_6737,N_8020);
nor U18293 (N_18293,N_345,N_1168);
nand U18294 (N_18294,N_7575,N_9282);
and U18295 (N_18295,N_3663,N_5377);
nand U18296 (N_18296,N_2765,N_1747);
nand U18297 (N_18297,N_3234,N_293);
nor U18298 (N_18298,N_8163,N_2608);
xnor U18299 (N_18299,N_5100,N_7612);
or U18300 (N_18300,N_6460,N_3415);
xor U18301 (N_18301,N_9564,N_5139);
nand U18302 (N_18302,N_3216,N_6368);
or U18303 (N_18303,N_142,N_5923);
or U18304 (N_18304,N_9461,N_902);
nor U18305 (N_18305,N_492,N_1336);
xnor U18306 (N_18306,N_9863,N_7561);
nor U18307 (N_18307,N_7091,N_9943);
or U18308 (N_18308,N_8620,N_6669);
nand U18309 (N_18309,N_4259,N_8556);
xnor U18310 (N_18310,N_9972,N_7201);
xor U18311 (N_18311,N_9,N_3856);
xnor U18312 (N_18312,N_2540,N_8754);
or U18313 (N_18313,N_6744,N_6579);
or U18314 (N_18314,N_3995,N_9927);
xor U18315 (N_18315,N_7862,N_4332);
nand U18316 (N_18316,N_3133,N_4689);
and U18317 (N_18317,N_126,N_9778);
and U18318 (N_18318,N_2163,N_8123);
nor U18319 (N_18319,N_9550,N_8541);
or U18320 (N_18320,N_5412,N_6991);
and U18321 (N_18321,N_5643,N_320);
nand U18322 (N_18322,N_6596,N_705);
nor U18323 (N_18323,N_8202,N_178);
nand U18324 (N_18324,N_1694,N_8109);
nand U18325 (N_18325,N_2131,N_6043);
and U18326 (N_18326,N_8579,N_6684);
or U18327 (N_18327,N_3179,N_7712);
or U18328 (N_18328,N_1429,N_8087);
or U18329 (N_18329,N_769,N_6649);
nor U18330 (N_18330,N_6740,N_2402);
nand U18331 (N_18331,N_1198,N_1394);
or U18332 (N_18332,N_2358,N_1864);
and U18333 (N_18333,N_3170,N_8117);
xnor U18334 (N_18334,N_5805,N_6908);
nor U18335 (N_18335,N_9540,N_1245);
and U18336 (N_18336,N_6698,N_9283);
nor U18337 (N_18337,N_7535,N_4258);
nor U18338 (N_18338,N_1096,N_5419);
nand U18339 (N_18339,N_800,N_5928);
or U18340 (N_18340,N_1378,N_1893);
nor U18341 (N_18341,N_3217,N_1861);
nor U18342 (N_18342,N_285,N_9536);
and U18343 (N_18343,N_2968,N_1042);
nand U18344 (N_18344,N_4704,N_615);
and U18345 (N_18345,N_1077,N_8170);
and U18346 (N_18346,N_8358,N_3134);
or U18347 (N_18347,N_5925,N_4651);
xnor U18348 (N_18348,N_8627,N_4064);
nand U18349 (N_18349,N_5213,N_830);
and U18350 (N_18350,N_2847,N_7474);
nor U18351 (N_18351,N_3754,N_1903);
and U18352 (N_18352,N_4573,N_3814);
xor U18353 (N_18353,N_1989,N_4300);
xnor U18354 (N_18354,N_5699,N_4680);
and U18355 (N_18355,N_8922,N_9569);
xnor U18356 (N_18356,N_9274,N_2235);
nand U18357 (N_18357,N_2872,N_141);
xnor U18358 (N_18358,N_3206,N_4015);
nor U18359 (N_18359,N_6150,N_9633);
nor U18360 (N_18360,N_2000,N_5789);
nand U18361 (N_18361,N_1173,N_7379);
nand U18362 (N_18362,N_2601,N_2757);
or U18363 (N_18363,N_6896,N_3537);
or U18364 (N_18364,N_5760,N_3579);
nand U18365 (N_18365,N_5805,N_7730);
and U18366 (N_18366,N_2248,N_1484);
and U18367 (N_18367,N_7857,N_9509);
nand U18368 (N_18368,N_6985,N_973);
and U18369 (N_18369,N_2877,N_3160);
and U18370 (N_18370,N_8253,N_5291);
nand U18371 (N_18371,N_6416,N_809);
nor U18372 (N_18372,N_211,N_3868);
nor U18373 (N_18373,N_2544,N_4104);
nor U18374 (N_18374,N_5545,N_2430);
xor U18375 (N_18375,N_4648,N_2922);
nor U18376 (N_18376,N_1286,N_4833);
or U18377 (N_18377,N_1267,N_906);
nor U18378 (N_18378,N_3139,N_8405);
xor U18379 (N_18379,N_4245,N_2508);
or U18380 (N_18380,N_1488,N_361);
or U18381 (N_18381,N_8118,N_2304);
or U18382 (N_18382,N_5528,N_8001);
nor U18383 (N_18383,N_3648,N_6916);
nor U18384 (N_18384,N_9519,N_3198);
nand U18385 (N_18385,N_9400,N_477);
and U18386 (N_18386,N_6888,N_9865);
or U18387 (N_18387,N_5160,N_4609);
nor U18388 (N_18388,N_565,N_5165);
nor U18389 (N_18389,N_7387,N_1807);
and U18390 (N_18390,N_4986,N_9385);
nand U18391 (N_18391,N_2072,N_3461);
nor U18392 (N_18392,N_6933,N_6432);
or U18393 (N_18393,N_3872,N_4823);
nand U18394 (N_18394,N_136,N_864);
xor U18395 (N_18395,N_5770,N_9589);
nor U18396 (N_18396,N_5359,N_5596);
nor U18397 (N_18397,N_6879,N_9131);
or U18398 (N_18398,N_4028,N_8642);
xor U18399 (N_18399,N_5970,N_9165);
or U18400 (N_18400,N_2107,N_3642);
and U18401 (N_18401,N_6134,N_2019);
and U18402 (N_18402,N_8560,N_6477);
xnor U18403 (N_18403,N_7563,N_9540);
nand U18404 (N_18404,N_4723,N_6321);
and U18405 (N_18405,N_7598,N_7734);
nand U18406 (N_18406,N_829,N_2948);
nor U18407 (N_18407,N_5675,N_1959);
and U18408 (N_18408,N_6385,N_2459);
or U18409 (N_18409,N_3143,N_6666);
and U18410 (N_18410,N_5532,N_9903);
xor U18411 (N_18411,N_9591,N_617);
nor U18412 (N_18412,N_5338,N_4604);
and U18413 (N_18413,N_7071,N_2639);
nand U18414 (N_18414,N_6041,N_16);
nor U18415 (N_18415,N_2097,N_6539);
or U18416 (N_18416,N_8057,N_828);
xnor U18417 (N_18417,N_430,N_4411);
nor U18418 (N_18418,N_1422,N_21);
xnor U18419 (N_18419,N_3060,N_535);
nor U18420 (N_18420,N_3508,N_4765);
nand U18421 (N_18421,N_5424,N_3261);
or U18422 (N_18422,N_6912,N_9874);
and U18423 (N_18423,N_2020,N_2228);
and U18424 (N_18424,N_7587,N_7578);
or U18425 (N_18425,N_7081,N_6878);
and U18426 (N_18426,N_8896,N_9809);
xnor U18427 (N_18427,N_6615,N_290);
nor U18428 (N_18428,N_1021,N_7089);
or U18429 (N_18429,N_7167,N_2045);
or U18430 (N_18430,N_5325,N_1101);
nor U18431 (N_18431,N_1117,N_8092);
or U18432 (N_18432,N_9834,N_6098);
nand U18433 (N_18433,N_7611,N_3143);
or U18434 (N_18434,N_4767,N_7152);
xor U18435 (N_18435,N_8891,N_1161);
and U18436 (N_18436,N_8599,N_6866);
nand U18437 (N_18437,N_5355,N_1615);
nand U18438 (N_18438,N_658,N_9120);
nor U18439 (N_18439,N_4663,N_9147);
and U18440 (N_18440,N_8607,N_1485);
nor U18441 (N_18441,N_747,N_478);
or U18442 (N_18442,N_1892,N_3995);
nor U18443 (N_18443,N_734,N_1790);
nand U18444 (N_18444,N_8958,N_3237);
xnor U18445 (N_18445,N_4297,N_7069);
nor U18446 (N_18446,N_7318,N_5217);
or U18447 (N_18447,N_1756,N_5935);
or U18448 (N_18448,N_1818,N_5290);
and U18449 (N_18449,N_5206,N_8701);
and U18450 (N_18450,N_980,N_3022);
or U18451 (N_18451,N_5333,N_5339);
or U18452 (N_18452,N_3784,N_2874);
nor U18453 (N_18453,N_5933,N_3248);
or U18454 (N_18454,N_5087,N_2454);
or U18455 (N_18455,N_4764,N_3443);
nand U18456 (N_18456,N_4649,N_7362);
and U18457 (N_18457,N_8134,N_9984);
nor U18458 (N_18458,N_69,N_8225);
or U18459 (N_18459,N_1969,N_8521);
or U18460 (N_18460,N_8868,N_7508);
and U18461 (N_18461,N_8574,N_1728);
nand U18462 (N_18462,N_1021,N_5395);
nand U18463 (N_18463,N_4215,N_6347);
nand U18464 (N_18464,N_8940,N_7610);
nand U18465 (N_18465,N_8708,N_239);
nand U18466 (N_18466,N_3832,N_9935);
nor U18467 (N_18467,N_575,N_7043);
nand U18468 (N_18468,N_2798,N_1128);
and U18469 (N_18469,N_5204,N_7564);
and U18470 (N_18470,N_113,N_7039);
or U18471 (N_18471,N_7191,N_7301);
xor U18472 (N_18472,N_8171,N_526);
nand U18473 (N_18473,N_1939,N_2057);
and U18474 (N_18474,N_7432,N_1030);
nand U18475 (N_18475,N_8185,N_9372);
nand U18476 (N_18476,N_669,N_9737);
and U18477 (N_18477,N_5318,N_9951);
nor U18478 (N_18478,N_9699,N_9337);
or U18479 (N_18479,N_625,N_7630);
nor U18480 (N_18480,N_9423,N_7352);
xnor U18481 (N_18481,N_504,N_9350);
nand U18482 (N_18482,N_5712,N_1852);
nor U18483 (N_18483,N_6677,N_8896);
or U18484 (N_18484,N_5334,N_5512);
or U18485 (N_18485,N_1062,N_923);
or U18486 (N_18486,N_7838,N_5086);
or U18487 (N_18487,N_1166,N_4086);
and U18488 (N_18488,N_3708,N_3660);
nor U18489 (N_18489,N_6799,N_3844);
or U18490 (N_18490,N_1721,N_7566);
and U18491 (N_18491,N_7068,N_944);
and U18492 (N_18492,N_7787,N_6699);
or U18493 (N_18493,N_3210,N_9562);
nand U18494 (N_18494,N_3543,N_2166);
nand U18495 (N_18495,N_3940,N_2317);
or U18496 (N_18496,N_7137,N_5437);
xor U18497 (N_18497,N_4390,N_7790);
and U18498 (N_18498,N_8465,N_8694);
nor U18499 (N_18499,N_9375,N_9856);
xnor U18500 (N_18500,N_1104,N_9828);
or U18501 (N_18501,N_1005,N_2794);
nand U18502 (N_18502,N_2052,N_1655);
and U18503 (N_18503,N_4129,N_8316);
nor U18504 (N_18504,N_4012,N_6732);
or U18505 (N_18505,N_5468,N_6760);
xnor U18506 (N_18506,N_1443,N_167);
xor U18507 (N_18507,N_7575,N_1701);
and U18508 (N_18508,N_5029,N_1785);
or U18509 (N_18509,N_2171,N_4004);
or U18510 (N_18510,N_7609,N_1544);
xor U18511 (N_18511,N_1423,N_4861);
xor U18512 (N_18512,N_8581,N_1511);
and U18513 (N_18513,N_9138,N_6573);
or U18514 (N_18514,N_17,N_8444);
xor U18515 (N_18515,N_3267,N_6675);
nand U18516 (N_18516,N_2708,N_1103);
nand U18517 (N_18517,N_5610,N_1434);
xor U18518 (N_18518,N_6125,N_9354);
nor U18519 (N_18519,N_4063,N_1482);
or U18520 (N_18520,N_1163,N_7389);
nand U18521 (N_18521,N_318,N_806);
xnor U18522 (N_18522,N_7359,N_3008);
and U18523 (N_18523,N_2986,N_967);
nor U18524 (N_18524,N_6615,N_9083);
or U18525 (N_18525,N_4101,N_6573);
and U18526 (N_18526,N_5161,N_7968);
nand U18527 (N_18527,N_8956,N_788);
nand U18528 (N_18528,N_8250,N_5379);
xor U18529 (N_18529,N_8625,N_3813);
nor U18530 (N_18530,N_4402,N_8866);
nor U18531 (N_18531,N_4526,N_329);
nand U18532 (N_18532,N_9402,N_9744);
nand U18533 (N_18533,N_5968,N_7075);
nor U18534 (N_18534,N_6761,N_1933);
and U18535 (N_18535,N_7913,N_1468);
nand U18536 (N_18536,N_9960,N_2689);
nor U18537 (N_18537,N_6983,N_2597);
and U18538 (N_18538,N_7303,N_6348);
xor U18539 (N_18539,N_4021,N_6713);
nand U18540 (N_18540,N_4615,N_7829);
and U18541 (N_18541,N_3835,N_6289);
xor U18542 (N_18542,N_3935,N_8719);
nand U18543 (N_18543,N_6372,N_9820);
and U18544 (N_18544,N_915,N_6160);
nand U18545 (N_18545,N_1671,N_8932);
xnor U18546 (N_18546,N_6731,N_5958);
or U18547 (N_18547,N_1685,N_1202);
and U18548 (N_18548,N_9370,N_5038);
nor U18549 (N_18549,N_8235,N_7024);
nor U18550 (N_18550,N_9095,N_2248);
nand U18551 (N_18551,N_9465,N_7543);
or U18552 (N_18552,N_2740,N_1844);
and U18553 (N_18553,N_5988,N_1618);
nand U18554 (N_18554,N_7382,N_7172);
or U18555 (N_18555,N_1539,N_3185);
and U18556 (N_18556,N_2110,N_8954);
or U18557 (N_18557,N_4179,N_5652);
nor U18558 (N_18558,N_2398,N_3344);
nor U18559 (N_18559,N_7885,N_5774);
xor U18560 (N_18560,N_1364,N_7423);
xnor U18561 (N_18561,N_8400,N_5553);
nor U18562 (N_18562,N_2635,N_2121);
or U18563 (N_18563,N_1449,N_4406);
xor U18564 (N_18564,N_8714,N_8125);
xnor U18565 (N_18565,N_4870,N_8212);
nand U18566 (N_18566,N_6260,N_3112);
xnor U18567 (N_18567,N_289,N_5341);
or U18568 (N_18568,N_8992,N_2816);
nor U18569 (N_18569,N_6535,N_9047);
and U18570 (N_18570,N_568,N_4053);
nand U18571 (N_18571,N_3776,N_1734);
or U18572 (N_18572,N_827,N_213);
and U18573 (N_18573,N_8315,N_4628);
nand U18574 (N_18574,N_7994,N_9242);
xnor U18575 (N_18575,N_3909,N_6716);
nand U18576 (N_18576,N_8847,N_3830);
or U18577 (N_18577,N_1884,N_64);
nand U18578 (N_18578,N_1383,N_7704);
and U18579 (N_18579,N_8923,N_6832);
nor U18580 (N_18580,N_1813,N_5556);
or U18581 (N_18581,N_9497,N_4966);
nor U18582 (N_18582,N_7611,N_6949);
and U18583 (N_18583,N_8811,N_4535);
and U18584 (N_18584,N_1486,N_331);
nor U18585 (N_18585,N_121,N_5839);
nand U18586 (N_18586,N_7368,N_2070);
or U18587 (N_18587,N_5486,N_2793);
and U18588 (N_18588,N_9874,N_773);
and U18589 (N_18589,N_2251,N_9228);
or U18590 (N_18590,N_2292,N_9507);
xnor U18591 (N_18591,N_8056,N_6537);
nand U18592 (N_18592,N_1577,N_6807);
and U18593 (N_18593,N_9676,N_6377);
or U18594 (N_18594,N_3058,N_443);
xnor U18595 (N_18595,N_8292,N_3814);
or U18596 (N_18596,N_9989,N_4830);
or U18597 (N_18597,N_2034,N_2997);
xor U18598 (N_18598,N_9563,N_6091);
nor U18599 (N_18599,N_6488,N_8792);
and U18600 (N_18600,N_5758,N_9370);
nand U18601 (N_18601,N_4180,N_6376);
nand U18602 (N_18602,N_6693,N_975);
nand U18603 (N_18603,N_1560,N_4622);
xor U18604 (N_18604,N_1391,N_3706);
nand U18605 (N_18605,N_8276,N_3264);
nor U18606 (N_18606,N_1397,N_4123);
nand U18607 (N_18607,N_636,N_3494);
nor U18608 (N_18608,N_6800,N_3097);
or U18609 (N_18609,N_9391,N_8555);
nand U18610 (N_18610,N_3714,N_6923);
nor U18611 (N_18611,N_2491,N_8905);
or U18612 (N_18612,N_7425,N_4686);
nor U18613 (N_18613,N_5546,N_977);
or U18614 (N_18614,N_9889,N_4444);
nor U18615 (N_18615,N_1260,N_4975);
xnor U18616 (N_18616,N_2383,N_1053);
and U18617 (N_18617,N_5056,N_879);
xor U18618 (N_18618,N_9488,N_4068);
or U18619 (N_18619,N_9151,N_7059);
xor U18620 (N_18620,N_1675,N_2527);
or U18621 (N_18621,N_7867,N_7217);
and U18622 (N_18622,N_8735,N_4112);
nand U18623 (N_18623,N_7024,N_8794);
xnor U18624 (N_18624,N_3875,N_1081);
or U18625 (N_18625,N_6157,N_1516);
or U18626 (N_18626,N_3761,N_2986);
and U18627 (N_18627,N_4223,N_6246);
or U18628 (N_18628,N_7460,N_849);
and U18629 (N_18629,N_9343,N_2469);
or U18630 (N_18630,N_7854,N_4376);
nor U18631 (N_18631,N_4693,N_2806);
nand U18632 (N_18632,N_8867,N_4112);
xnor U18633 (N_18633,N_9805,N_4819);
or U18634 (N_18634,N_4631,N_1947);
nand U18635 (N_18635,N_9399,N_990);
nor U18636 (N_18636,N_7616,N_6211);
xnor U18637 (N_18637,N_1268,N_8055);
or U18638 (N_18638,N_2250,N_3572);
or U18639 (N_18639,N_6646,N_6955);
xnor U18640 (N_18640,N_275,N_1544);
nor U18641 (N_18641,N_9714,N_1916);
nand U18642 (N_18642,N_3886,N_8173);
or U18643 (N_18643,N_4870,N_4431);
or U18644 (N_18644,N_7317,N_7808);
nor U18645 (N_18645,N_2756,N_7286);
or U18646 (N_18646,N_4402,N_4113);
and U18647 (N_18647,N_5345,N_2792);
and U18648 (N_18648,N_2184,N_103);
xnor U18649 (N_18649,N_655,N_6687);
nand U18650 (N_18650,N_4317,N_5050);
and U18651 (N_18651,N_7782,N_348);
or U18652 (N_18652,N_1267,N_9858);
and U18653 (N_18653,N_9116,N_3228);
nand U18654 (N_18654,N_8602,N_6622);
nand U18655 (N_18655,N_246,N_6511);
and U18656 (N_18656,N_9969,N_6159);
nand U18657 (N_18657,N_6481,N_1015);
and U18658 (N_18658,N_4310,N_6927);
xor U18659 (N_18659,N_1807,N_7126);
xnor U18660 (N_18660,N_8519,N_5537);
nand U18661 (N_18661,N_9671,N_2728);
nor U18662 (N_18662,N_3195,N_6963);
and U18663 (N_18663,N_3705,N_7738);
nand U18664 (N_18664,N_1857,N_7259);
and U18665 (N_18665,N_971,N_1175);
xnor U18666 (N_18666,N_6552,N_1693);
xnor U18667 (N_18667,N_5495,N_5372);
xnor U18668 (N_18668,N_3751,N_7656);
nor U18669 (N_18669,N_9223,N_603);
xnor U18670 (N_18670,N_4404,N_9251);
xnor U18671 (N_18671,N_5034,N_9458);
nor U18672 (N_18672,N_7839,N_5215);
nor U18673 (N_18673,N_5559,N_5482);
or U18674 (N_18674,N_642,N_7739);
or U18675 (N_18675,N_1158,N_9648);
xnor U18676 (N_18676,N_4023,N_7935);
or U18677 (N_18677,N_4259,N_4384);
xnor U18678 (N_18678,N_7523,N_6835);
xnor U18679 (N_18679,N_4562,N_2915);
xnor U18680 (N_18680,N_952,N_9028);
nand U18681 (N_18681,N_3796,N_7112);
xor U18682 (N_18682,N_4502,N_9251);
or U18683 (N_18683,N_6020,N_9051);
and U18684 (N_18684,N_3467,N_6456);
nor U18685 (N_18685,N_7951,N_4149);
and U18686 (N_18686,N_1059,N_9235);
and U18687 (N_18687,N_7223,N_4080);
nand U18688 (N_18688,N_7630,N_5202);
nand U18689 (N_18689,N_1997,N_2423);
xnor U18690 (N_18690,N_5437,N_1396);
xnor U18691 (N_18691,N_84,N_5987);
and U18692 (N_18692,N_5106,N_2837);
or U18693 (N_18693,N_5011,N_8913);
xor U18694 (N_18694,N_1864,N_2444);
xnor U18695 (N_18695,N_9822,N_6639);
and U18696 (N_18696,N_5641,N_6275);
xnor U18697 (N_18697,N_3038,N_1482);
and U18698 (N_18698,N_7801,N_6070);
nor U18699 (N_18699,N_4812,N_9660);
nand U18700 (N_18700,N_200,N_6996);
xor U18701 (N_18701,N_7335,N_6979);
xnor U18702 (N_18702,N_2143,N_8109);
nor U18703 (N_18703,N_7592,N_400);
xnor U18704 (N_18704,N_46,N_4582);
or U18705 (N_18705,N_1170,N_7171);
xor U18706 (N_18706,N_276,N_8781);
or U18707 (N_18707,N_6002,N_3483);
or U18708 (N_18708,N_5122,N_3227);
nand U18709 (N_18709,N_8963,N_4126);
or U18710 (N_18710,N_440,N_4501);
nor U18711 (N_18711,N_1213,N_7263);
xor U18712 (N_18712,N_359,N_5915);
nand U18713 (N_18713,N_4484,N_793);
and U18714 (N_18714,N_1707,N_8033);
and U18715 (N_18715,N_1746,N_6787);
xor U18716 (N_18716,N_5441,N_607);
and U18717 (N_18717,N_4643,N_4677);
nand U18718 (N_18718,N_696,N_8372);
and U18719 (N_18719,N_9109,N_4318);
and U18720 (N_18720,N_2411,N_4999);
nand U18721 (N_18721,N_4912,N_8080);
or U18722 (N_18722,N_6374,N_7185);
or U18723 (N_18723,N_6990,N_9862);
or U18724 (N_18724,N_8166,N_9164);
or U18725 (N_18725,N_6888,N_5304);
xnor U18726 (N_18726,N_1282,N_4078);
xnor U18727 (N_18727,N_6886,N_7186);
nor U18728 (N_18728,N_6930,N_6993);
xnor U18729 (N_18729,N_8474,N_2922);
nor U18730 (N_18730,N_4611,N_4017);
and U18731 (N_18731,N_3820,N_7927);
nand U18732 (N_18732,N_9058,N_8353);
nor U18733 (N_18733,N_6738,N_7274);
and U18734 (N_18734,N_556,N_8700);
nand U18735 (N_18735,N_7769,N_8566);
nor U18736 (N_18736,N_745,N_5898);
and U18737 (N_18737,N_4412,N_2627);
xor U18738 (N_18738,N_4185,N_15);
nor U18739 (N_18739,N_1340,N_6504);
nor U18740 (N_18740,N_9327,N_2527);
or U18741 (N_18741,N_1382,N_2987);
nor U18742 (N_18742,N_8710,N_6703);
nand U18743 (N_18743,N_7356,N_8815);
xnor U18744 (N_18744,N_6920,N_2408);
nor U18745 (N_18745,N_3018,N_3026);
or U18746 (N_18746,N_6948,N_6848);
nor U18747 (N_18747,N_7111,N_4273);
nand U18748 (N_18748,N_1406,N_4645);
nor U18749 (N_18749,N_5805,N_3988);
nand U18750 (N_18750,N_5336,N_6490);
and U18751 (N_18751,N_7797,N_6407);
and U18752 (N_18752,N_3319,N_8895);
nand U18753 (N_18753,N_4284,N_3003);
or U18754 (N_18754,N_6311,N_2781);
nor U18755 (N_18755,N_1186,N_9610);
nand U18756 (N_18756,N_1749,N_190);
or U18757 (N_18757,N_2791,N_2345);
xnor U18758 (N_18758,N_8490,N_8002);
xor U18759 (N_18759,N_8172,N_2515);
xnor U18760 (N_18760,N_3552,N_7706);
or U18761 (N_18761,N_1691,N_7849);
and U18762 (N_18762,N_1175,N_4085);
nor U18763 (N_18763,N_9404,N_3141);
nor U18764 (N_18764,N_7323,N_3638);
xnor U18765 (N_18765,N_4480,N_5076);
or U18766 (N_18766,N_1201,N_6891);
nand U18767 (N_18767,N_423,N_223);
and U18768 (N_18768,N_6176,N_1416);
and U18769 (N_18769,N_9716,N_507);
xnor U18770 (N_18770,N_393,N_2190);
or U18771 (N_18771,N_6325,N_9577);
nand U18772 (N_18772,N_2847,N_9352);
nor U18773 (N_18773,N_5126,N_1914);
or U18774 (N_18774,N_4688,N_9113);
and U18775 (N_18775,N_3075,N_6533);
nor U18776 (N_18776,N_4678,N_501);
xnor U18777 (N_18777,N_8037,N_7061);
or U18778 (N_18778,N_3264,N_5778);
nor U18779 (N_18779,N_7586,N_4384);
and U18780 (N_18780,N_4760,N_3843);
nand U18781 (N_18781,N_577,N_2923);
xnor U18782 (N_18782,N_3062,N_4423);
or U18783 (N_18783,N_5533,N_2594);
or U18784 (N_18784,N_3049,N_2534);
and U18785 (N_18785,N_3581,N_5884);
nor U18786 (N_18786,N_6486,N_7312);
and U18787 (N_18787,N_9180,N_3686);
nor U18788 (N_18788,N_6935,N_6291);
nor U18789 (N_18789,N_6421,N_3594);
nand U18790 (N_18790,N_7490,N_3688);
or U18791 (N_18791,N_5238,N_9721);
or U18792 (N_18792,N_8327,N_1718);
nor U18793 (N_18793,N_1023,N_5741);
xor U18794 (N_18794,N_5339,N_347);
nand U18795 (N_18795,N_6834,N_2500);
nand U18796 (N_18796,N_4430,N_1173);
nor U18797 (N_18797,N_5663,N_5746);
nand U18798 (N_18798,N_5264,N_7293);
and U18799 (N_18799,N_2325,N_1505);
nand U18800 (N_18800,N_6635,N_9038);
nand U18801 (N_18801,N_6221,N_462);
xor U18802 (N_18802,N_2404,N_1556);
or U18803 (N_18803,N_7974,N_3424);
nand U18804 (N_18804,N_9242,N_1545);
nand U18805 (N_18805,N_6290,N_7384);
and U18806 (N_18806,N_6776,N_3033);
xnor U18807 (N_18807,N_6417,N_6439);
nor U18808 (N_18808,N_791,N_4141);
or U18809 (N_18809,N_5211,N_4168);
nor U18810 (N_18810,N_8234,N_21);
and U18811 (N_18811,N_3393,N_9543);
nor U18812 (N_18812,N_2725,N_4247);
or U18813 (N_18813,N_5464,N_266);
or U18814 (N_18814,N_9250,N_1315);
nor U18815 (N_18815,N_142,N_9857);
xnor U18816 (N_18816,N_4844,N_386);
or U18817 (N_18817,N_9444,N_8790);
xor U18818 (N_18818,N_521,N_4494);
nor U18819 (N_18819,N_7869,N_676);
nor U18820 (N_18820,N_1314,N_6614);
or U18821 (N_18821,N_7913,N_3893);
and U18822 (N_18822,N_821,N_1511);
xor U18823 (N_18823,N_1887,N_3167);
nor U18824 (N_18824,N_2511,N_1895);
or U18825 (N_18825,N_163,N_2924);
and U18826 (N_18826,N_3677,N_6581);
xnor U18827 (N_18827,N_8037,N_4394);
and U18828 (N_18828,N_8473,N_9882);
and U18829 (N_18829,N_3503,N_8911);
nor U18830 (N_18830,N_2917,N_6910);
or U18831 (N_18831,N_4522,N_4516);
and U18832 (N_18832,N_3341,N_324);
nor U18833 (N_18833,N_1168,N_8411);
nand U18834 (N_18834,N_4924,N_8077);
and U18835 (N_18835,N_719,N_2659);
nand U18836 (N_18836,N_7815,N_7126);
or U18837 (N_18837,N_9145,N_9234);
or U18838 (N_18838,N_6693,N_3824);
and U18839 (N_18839,N_6456,N_687);
nand U18840 (N_18840,N_5912,N_9851);
nor U18841 (N_18841,N_3858,N_3245);
nand U18842 (N_18842,N_958,N_5735);
and U18843 (N_18843,N_966,N_3952);
or U18844 (N_18844,N_7192,N_689);
nand U18845 (N_18845,N_3207,N_2271);
nor U18846 (N_18846,N_9744,N_4766);
nand U18847 (N_18847,N_5387,N_9948);
and U18848 (N_18848,N_7860,N_2522);
or U18849 (N_18849,N_7611,N_6450);
nor U18850 (N_18850,N_4062,N_5172);
nor U18851 (N_18851,N_2842,N_6145);
nand U18852 (N_18852,N_2196,N_4289);
xnor U18853 (N_18853,N_1521,N_7003);
xor U18854 (N_18854,N_2901,N_3923);
nor U18855 (N_18855,N_9909,N_2405);
xor U18856 (N_18856,N_2628,N_2476);
or U18857 (N_18857,N_5820,N_9819);
xnor U18858 (N_18858,N_9509,N_8374);
xor U18859 (N_18859,N_5359,N_6560);
xor U18860 (N_18860,N_3771,N_9746);
nand U18861 (N_18861,N_7081,N_2407);
or U18862 (N_18862,N_3143,N_4968);
nor U18863 (N_18863,N_3575,N_3956);
nor U18864 (N_18864,N_6650,N_6937);
xor U18865 (N_18865,N_2707,N_2804);
xnor U18866 (N_18866,N_2861,N_2386);
xor U18867 (N_18867,N_4928,N_6462);
nor U18868 (N_18868,N_1303,N_1137);
or U18869 (N_18869,N_1382,N_8553);
xor U18870 (N_18870,N_9478,N_3082);
or U18871 (N_18871,N_1051,N_8707);
nand U18872 (N_18872,N_3337,N_957);
nor U18873 (N_18873,N_7888,N_9075);
nand U18874 (N_18874,N_4850,N_3965);
xor U18875 (N_18875,N_5813,N_1731);
or U18876 (N_18876,N_7996,N_720);
or U18877 (N_18877,N_8176,N_5649);
nand U18878 (N_18878,N_8398,N_7523);
or U18879 (N_18879,N_4273,N_4157);
or U18880 (N_18880,N_2662,N_1089);
nand U18881 (N_18881,N_4044,N_6810);
and U18882 (N_18882,N_6307,N_7345);
nand U18883 (N_18883,N_3708,N_3015);
xnor U18884 (N_18884,N_9233,N_3755);
nand U18885 (N_18885,N_1688,N_8910);
xor U18886 (N_18886,N_1576,N_3404);
nor U18887 (N_18887,N_6865,N_4479);
nor U18888 (N_18888,N_6894,N_8468);
nor U18889 (N_18889,N_6404,N_7000);
xnor U18890 (N_18890,N_339,N_7641);
nor U18891 (N_18891,N_2472,N_1895);
nor U18892 (N_18892,N_4080,N_9919);
nand U18893 (N_18893,N_2903,N_1184);
or U18894 (N_18894,N_5749,N_2744);
or U18895 (N_18895,N_2300,N_8869);
nand U18896 (N_18896,N_6342,N_8121);
or U18897 (N_18897,N_7053,N_159);
nor U18898 (N_18898,N_2154,N_3874);
xnor U18899 (N_18899,N_6645,N_7102);
nand U18900 (N_18900,N_1796,N_7498);
or U18901 (N_18901,N_9508,N_6133);
or U18902 (N_18902,N_8418,N_3415);
and U18903 (N_18903,N_2995,N_6193);
xor U18904 (N_18904,N_3394,N_7676);
xor U18905 (N_18905,N_5726,N_2815);
nand U18906 (N_18906,N_1295,N_3232);
xor U18907 (N_18907,N_703,N_5679);
or U18908 (N_18908,N_8171,N_4041);
and U18909 (N_18909,N_6511,N_9398);
xor U18910 (N_18910,N_7641,N_7100);
and U18911 (N_18911,N_6539,N_945);
or U18912 (N_18912,N_5859,N_8464);
nor U18913 (N_18913,N_7527,N_2549);
or U18914 (N_18914,N_8621,N_7957);
or U18915 (N_18915,N_1074,N_4898);
or U18916 (N_18916,N_6671,N_8899);
and U18917 (N_18917,N_9817,N_208);
xnor U18918 (N_18918,N_973,N_2026);
and U18919 (N_18919,N_6596,N_765);
xor U18920 (N_18920,N_7824,N_2766);
and U18921 (N_18921,N_7853,N_5945);
or U18922 (N_18922,N_9576,N_7966);
and U18923 (N_18923,N_1217,N_2335);
nand U18924 (N_18924,N_8753,N_9619);
nor U18925 (N_18925,N_7801,N_514);
and U18926 (N_18926,N_5301,N_5172);
xnor U18927 (N_18927,N_2794,N_1089);
or U18928 (N_18928,N_6154,N_8124);
and U18929 (N_18929,N_994,N_5738);
and U18930 (N_18930,N_7622,N_1307);
and U18931 (N_18931,N_5588,N_4780);
and U18932 (N_18932,N_5064,N_7114);
nand U18933 (N_18933,N_2841,N_7604);
xnor U18934 (N_18934,N_6887,N_6755);
or U18935 (N_18935,N_8920,N_9699);
xor U18936 (N_18936,N_8810,N_5500);
nor U18937 (N_18937,N_8140,N_5232);
or U18938 (N_18938,N_3218,N_7968);
xnor U18939 (N_18939,N_7258,N_9029);
nor U18940 (N_18940,N_2165,N_9512);
nand U18941 (N_18941,N_4698,N_6513);
nand U18942 (N_18942,N_43,N_1079);
nor U18943 (N_18943,N_2097,N_6917);
or U18944 (N_18944,N_5430,N_6617);
xnor U18945 (N_18945,N_4187,N_2094);
nand U18946 (N_18946,N_9792,N_8681);
or U18947 (N_18947,N_6602,N_1873);
xor U18948 (N_18948,N_8407,N_8186);
or U18949 (N_18949,N_9185,N_8275);
or U18950 (N_18950,N_4954,N_6639);
or U18951 (N_18951,N_6130,N_7863);
or U18952 (N_18952,N_291,N_2639);
or U18953 (N_18953,N_68,N_7977);
xnor U18954 (N_18954,N_2209,N_6511);
and U18955 (N_18955,N_8189,N_3897);
nor U18956 (N_18956,N_3173,N_8470);
and U18957 (N_18957,N_4420,N_5781);
nor U18958 (N_18958,N_1841,N_6832);
nor U18959 (N_18959,N_5509,N_652);
xor U18960 (N_18960,N_1055,N_519);
nand U18961 (N_18961,N_7676,N_9470);
and U18962 (N_18962,N_3372,N_1537);
xnor U18963 (N_18963,N_5446,N_9419);
and U18964 (N_18964,N_3478,N_4993);
xnor U18965 (N_18965,N_9660,N_2864);
nor U18966 (N_18966,N_317,N_484);
nand U18967 (N_18967,N_2369,N_954);
nand U18968 (N_18968,N_164,N_2962);
nand U18969 (N_18969,N_4886,N_2862);
xor U18970 (N_18970,N_1983,N_5534);
xnor U18971 (N_18971,N_7095,N_42);
and U18972 (N_18972,N_6249,N_357);
and U18973 (N_18973,N_5896,N_9090);
or U18974 (N_18974,N_4402,N_8562);
nor U18975 (N_18975,N_9063,N_9813);
or U18976 (N_18976,N_378,N_7232);
nand U18977 (N_18977,N_2835,N_516);
or U18978 (N_18978,N_5017,N_3024);
and U18979 (N_18979,N_2929,N_7713);
nand U18980 (N_18980,N_8621,N_8708);
nor U18981 (N_18981,N_3395,N_8822);
nor U18982 (N_18982,N_204,N_5516);
and U18983 (N_18983,N_1011,N_9188);
xor U18984 (N_18984,N_3056,N_3644);
and U18985 (N_18985,N_5607,N_3111);
xnor U18986 (N_18986,N_6931,N_5599);
nor U18987 (N_18987,N_2542,N_9203);
nand U18988 (N_18988,N_7725,N_2499);
nand U18989 (N_18989,N_2882,N_5468);
or U18990 (N_18990,N_4504,N_6787);
nor U18991 (N_18991,N_219,N_1527);
and U18992 (N_18992,N_9537,N_3534);
or U18993 (N_18993,N_7332,N_2777);
or U18994 (N_18994,N_1974,N_1372);
or U18995 (N_18995,N_6870,N_9810);
nor U18996 (N_18996,N_8165,N_1720);
and U18997 (N_18997,N_3532,N_7376);
and U18998 (N_18998,N_6671,N_1542);
xnor U18999 (N_18999,N_7173,N_636);
or U19000 (N_19000,N_846,N_9281);
xor U19001 (N_19001,N_3881,N_5082);
or U19002 (N_19002,N_3074,N_3857);
or U19003 (N_19003,N_3896,N_1121);
or U19004 (N_19004,N_3759,N_862);
xor U19005 (N_19005,N_6700,N_4279);
nor U19006 (N_19006,N_6637,N_3426);
xnor U19007 (N_19007,N_6303,N_1268);
and U19008 (N_19008,N_6811,N_9986);
xor U19009 (N_19009,N_9941,N_6113);
or U19010 (N_19010,N_4402,N_3826);
xor U19011 (N_19011,N_6048,N_9843);
or U19012 (N_19012,N_9374,N_4399);
xnor U19013 (N_19013,N_2746,N_2912);
or U19014 (N_19014,N_2051,N_6742);
nor U19015 (N_19015,N_7522,N_4257);
nand U19016 (N_19016,N_5052,N_7487);
xor U19017 (N_19017,N_5118,N_3659);
nor U19018 (N_19018,N_9864,N_3860);
xnor U19019 (N_19019,N_9049,N_1585);
and U19020 (N_19020,N_2469,N_5795);
nand U19021 (N_19021,N_5587,N_8316);
nor U19022 (N_19022,N_9008,N_4684);
nand U19023 (N_19023,N_1450,N_5139);
or U19024 (N_19024,N_3975,N_9097);
nor U19025 (N_19025,N_1239,N_2454);
or U19026 (N_19026,N_9242,N_195);
nand U19027 (N_19027,N_8491,N_8155);
xor U19028 (N_19028,N_9817,N_8921);
nand U19029 (N_19029,N_2468,N_3000);
xor U19030 (N_19030,N_1962,N_1006);
nor U19031 (N_19031,N_7598,N_5506);
nor U19032 (N_19032,N_9443,N_1580);
xnor U19033 (N_19033,N_1118,N_1722);
and U19034 (N_19034,N_9281,N_487);
nor U19035 (N_19035,N_3693,N_1451);
nand U19036 (N_19036,N_1204,N_4709);
or U19037 (N_19037,N_9035,N_2544);
xnor U19038 (N_19038,N_3448,N_1195);
nand U19039 (N_19039,N_9736,N_9611);
nand U19040 (N_19040,N_5470,N_5123);
xnor U19041 (N_19041,N_286,N_5819);
xor U19042 (N_19042,N_1115,N_3782);
xnor U19043 (N_19043,N_8460,N_9850);
and U19044 (N_19044,N_3741,N_2505);
nand U19045 (N_19045,N_7027,N_4920);
xor U19046 (N_19046,N_2248,N_1935);
and U19047 (N_19047,N_6501,N_1075);
or U19048 (N_19048,N_8783,N_6659);
nand U19049 (N_19049,N_4122,N_7163);
or U19050 (N_19050,N_3016,N_5160);
or U19051 (N_19051,N_8312,N_7343);
and U19052 (N_19052,N_6466,N_8270);
nor U19053 (N_19053,N_6570,N_4924);
nor U19054 (N_19054,N_4653,N_284);
nor U19055 (N_19055,N_7569,N_9395);
nand U19056 (N_19056,N_7657,N_4694);
and U19057 (N_19057,N_5712,N_8945);
nand U19058 (N_19058,N_2895,N_23);
and U19059 (N_19059,N_9355,N_6191);
nor U19060 (N_19060,N_8478,N_8492);
nand U19061 (N_19061,N_92,N_3580);
xor U19062 (N_19062,N_1086,N_9288);
and U19063 (N_19063,N_8243,N_4745);
xnor U19064 (N_19064,N_5794,N_7004);
nor U19065 (N_19065,N_6243,N_9591);
xnor U19066 (N_19066,N_2694,N_9152);
and U19067 (N_19067,N_2567,N_6926);
nor U19068 (N_19068,N_735,N_8926);
xor U19069 (N_19069,N_5958,N_2198);
xor U19070 (N_19070,N_6112,N_3071);
and U19071 (N_19071,N_4514,N_3623);
nor U19072 (N_19072,N_5217,N_98);
xnor U19073 (N_19073,N_6326,N_5838);
nor U19074 (N_19074,N_4979,N_9839);
nand U19075 (N_19075,N_9697,N_951);
xnor U19076 (N_19076,N_2756,N_8176);
nor U19077 (N_19077,N_4295,N_8128);
nor U19078 (N_19078,N_3458,N_3410);
xnor U19079 (N_19079,N_3849,N_3711);
and U19080 (N_19080,N_4044,N_2309);
xnor U19081 (N_19081,N_8577,N_766);
and U19082 (N_19082,N_3947,N_1769);
or U19083 (N_19083,N_9049,N_6534);
and U19084 (N_19084,N_6270,N_7869);
or U19085 (N_19085,N_8390,N_8018);
nor U19086 (N_19086,N_5141,N_1684);
and U19087 (N_19087,N_5126,N_9382);
or U19088 (N_19088,N_6373,N_7373);
nand U19089 (N_19089,N_5992,N_9214);
and U19090 (N_19090,N_6236,N_7075);
xor U19091 (N_19091,N_2522,N_5917);
and U19092 (N_19092,N_2845,N_4454);
nand U19093 (N_19093,N_5382,N_9653);
nor U19094 (N_19094,N_9632,N_6687);
nand U19095 (N_19095,N_8930,N_2743);
xor U19096 (N_19096,N_3980,N_61);
xnor U19097 (N_19097,N_861,N_8838);
or U19098 (N_19098,N_506,N_3538);
xor U19099 (N_19099,N_3782,N_8907);
xnor U19100 (N_19100,N_528,N_1614);
xnor U19101 (N_19101,N_6377,N_3111);
nor U19102 (N_19102,N_4310,N_996);
or U19103 (N_19103,N_9489,N_4625);
and U19104 (N_19104,N_4663,N_1292);
xor U19105 (N_19105,N_2954,N_4634);
and U19106 (N_19106,N_3749,N_3648);
or U19107 (N_19107,N_4738,N_620);
and U19108 (N_19108,N_1112,N_6626);
nor U19109 (N_19109,N_3128,N_5655);
and U19110 (N_19110,N_1809,N_8535);
nor U19111 (N_19111,N_9568,N_9319);
nor U19112 (N_19112,N_3210,N_2219);
xor U19113 (N_19113,N_7200,N_1850);
or U19114 (N_19114,N_2600,N_9830);
or U19115 (N_19115,N_4403,N_5090);
nand U19116 (N_19116,N_8488,N_3679);
and U19117 (N_19117,N_3225,N_8511);
and U19118 (N_19118,N_4199,N_2574);
xor U19119 (N_19119,N_5850,N_1714);
nor U19120 (N_19120,N_8995,N_6632);
and U19121 (N_19121,N_5568,N_4756);
or U19122 (N_19122,N_803,N_8687);
nand U19123 (N_19123,N_2711,N_6237);
and U19124 (N_19124,N_7001,N_5580);
xor U19125 (N_19125,N_8805,N_4741);
and U19126 (N_19126,N_2565,N_6640);
nor U19127 (N_19127,N_2205,N_2519);
or U19128 (N_19128,N_7739,N_8460);
and U19129 (N_19129,N_9953,N_2707);
nor U19130 (N_19130,N_7133,N_5108);
xor U19131 (N_19131,N_9395,N_7666);
and U19132 (N_19132,N_6796,N_8852);
xor U19133 (N_19133,N_3176,N_2584);
nor U19134 (N_19134,N_2799,N_8080);
nand U19135 (N_19135,N_9780,N_1470);
or U19136 (N_19136,N_5282,N_5001);
and U19137 (N_19137,N_7733,N_6185);
nand U19138 (N_19138,N_5895,N_6176);
or U19139 (N_19139,N_7089,N_1828);
xnor U19140 (N_19140,N_4277,N_8716);
or U19141 (N_19141,N_328,N_5945);
nand U19142 (N_19142,N_1366,N_5677);
or U19143 (N_19143,N_5172,N_4180);
nand U19144 (N_19144,N_9995,N_6475);
xnor U19145 (N_19145,N_5534,N_817);
xnor U19146 (N_19146,N_3170,N_3270);
xnor U19147 (N_19147,N_5618,N_5530);
and U19148 (N_19148,N_105,N_7464);
or U19149 (N_19149,N_7601,N_4677);
nand U19150 (N_19150,N_9175,N_4223);
nand U19151 (N_19151,N_5871,N_8764);
xor U19152 (N_19152,N_6400,N_3122);
and U19153 (N_19153,N_1835,N_6158);
nand U19154 (N_19154,N_6161,N_4303);
or U19155 (N_19155,N_8001,N_2788);
and U19156 (N_19156,N_5323,N_3887);
or U19157 (N_19157,N_4724,N_3089);
or U19158 (N_19158,N_2428,N_2855);
nor U19159 (N_19159,N_4451,N_2769);
or U19160 (N_19160,N_5994,N_4035);
xnor U19161 (N_19161,N_1727,N_7249);
or U19162 (N_19162,N_1733,N_1942);
and U19163 (N_19163,N_2680,N_617);
or U19164 (N_19164,N_8867,N_681);
xnor U19165 (N_19165,N_4551,N_443);
nor U19166 (N_19166,N_4885,N_4676);
xnor U19167 (N_19167,N_9008,N_209);
nor U19168 (N_19168,N_8600,N_3799);
and U19169 (N_19169,N_5771,N_5591);
nor U19170 (N_19170,N_3112,N_3673);
and U19171 (N_19171,N_5678,N_4680);
and U19172 (N_19172,N_8610,N_8764);
nor U19173 (N_19173,N_2295,N_1114);
xnor U19174 (N_19174,N_1554,N_4825);
nand U19175 (N_19175,N_7816,N_2606);
xor U19176 (N_19176,N_8879,N_5458);
and U19177 (N_19177,N_4324,N_2802);
xor U19178 (N_19178,N_2996,N_6743);
nor U19179 (N_19179,N_8467,N_9367);
and U19180 (N_19180,N_9935,N_3523);
nand U19181 (N_19181,N_962,N_2928);
nand U19182 (N_19182,N_7273,N_9874);
nor U19183 (N_19183,N_2920,N_6683);
nand U19184 (N_19184,N_8327,N_1861);
nor U19185 (N_19185,N_8390,N_6771);
xor U19186 (N_19186,N_9398,N_6217);
and U19187 (N_19187,N_4921,N_4871);
and U19188 (N_19188,N_6454,N_958);
and U19189 (N_19189,N_8742,N_1897);
nor U19190 (N_19190,N_1721,N_634);
nor U19191 (N_19191,N_2414,N_7771);
nor U19192 (N_19192,N_8740,N_3540);
xor U19193 (N_19193,N_1335,N_1394);
and U19194 (N_19194,N_6577,N_7918);
nor U19195 (N_19195,N_2946,N_9373);
or U19196 (N_19196,N_2145,N_1918);
and U19197 (N_19197,N_2892,N_7732);
nor U19198 (N_19198,N_8350,N_5214);
nand U19199 (N_19199,N_1586,N_2412);
and U19200 (N_19200,N_9442,N_8169);
nand U19201 (N_19201,N_8948,N_2425);
xnor U19202 (N_19202,N_3319,N_1244);
nand U19203 (N_19203,N_1575,N_1053);
nand U19204 (N_19204,N_4026,N_2305);
and U19205 (N_19205,N_8707,N_5269);
nand U19206 (N_19206,N_5278,N_9080);
xnor U19207 (N_19207,N_7640,N_1029);
xnor U19208 (N_19208,N_4067,N_2613);
and U19209 (N_19209,N_9297,N_5247);
xor U19210 (N_19210,N_186,N_4991);
and U19211 (N_19211,N_8517,N_334);
or U19212 (N_19212,N_3305,N_3494);
xor U19213 (N_19213,N_6136,N_2193);
and U19214 (N_19214,N_7608,N_8381);
and U19215 (N_19215,N_6188,N_6994);
xnor U19216 (N_19216,N_8547,N_4961);
xor U19217 (N_19217,N_9034,N_8271);
xor U19218 (N_19218,N_8929,N_2655);
nor U19219 (N_19219,N_3203,N_7376);
and U19220 (N_19220,N_8263,N_6261);
xnor U19221 (N_19221,N_4252,N_3139);
and U19222 (N_19222,N_1225,N_9033);
nand U19223 (N_19223,N_7414,N_3381);
or U19224 (N_19224,N_9226,N_2819);
and U19225 (N_19225,N_5525,N_3858);
xor U19226 (N_19226,N_6869,N_2307);
or U19227 (N_19227,N_6256,N_1328);
nand U19228 (N_19228,N_1649,N_1122);
or U19229 (N_19229,N_2616,N_869);
xnor U19230 (N_19230,N_2712,N_8302);
or U19231 (N_19231,N_2592,N_6568);
nor U19232 (N_19232,N_9745,N_5424);
xor U19233 (N_19233,N_6267,N_7680);
xor U19234 (N_19234,N_3473,N_3088);
nand U19235 (N_19235,N_3227,N_4360);
nor U19236 (N_19236,N_4025,N_8886);
nor U19237 (N_19237,N_7678,N_7707);
nand U19238 (N_19238,N_7641,N_1423);
nand U19239 (N_19239,N_3215,N_6150);
nor U19240 (N_19240,N_2565,N_3340);
xor U19241 (N_19241,N_8807,N_236);
nor U19242 (N_19242,N_4366,N_5213);
and U19243 (N_19243,N_3796,N_601);
nand U19244 (N_19244,N_5465,N_1412);
and U19245 (N_19245,N_2700,N_4948);
nand U19246 (N_19246,N_6705,N_8636);
and U19247 (N_19247,N_7523,N_6695);
xor U19248 (N_19248,N_3602,N_2803);
nand U19249 (N_19249,N_2676,N_311);
and U19250 (N_19250,N_7957,N_9621);
nand U19251 (N_19251,N_2693,N_5421);
nor U19252 (N_19252,N_479,N_7500);
or U19253 (N_19253,N_4976,N_7466);
nor U19254 (N_19254,N_5410,N_8447);
xnor U19255 (N_19255,N_6472,N_6246);
xnor U19256 (N_19256,N_6900,N_6313);
or U19257 (N_19257,N_8838,N_4459);
or U19258 (N_19258,N_3267,N_4495);
or U19259 (N_19259,N_2188,N_5620);
nor U19260 (N_19260,N_5232,N_6744);
or U19261 (N_19261,N_9048,N_5298);
or U19262 (N_19262,N_2171,N_4686);
nand U19263 (N_19263,N_2127,N_9431);
xnor U19264 (N_19264,N_9668,N_2809);
or U19265 (N_19265,N_4253,N_3728);
and U19266 (N_19266,N_51,N_7338);
nand U19267 (N_19267,N_2652,N_8582);
nor U19268 (N_19268,N_5410,N_1492);
nand U19269 (N_19269,N_2385,N_2584);
or U19270 (N_19270,N_1125,N_6349);
and U19271 (N_19271,N_8818,N_5527);
nand U19272 (N_19272,N_3539,N_1651);
or U19273 (N_19273,N_3736,N_6359);
and U19274 (N_19274,N_3478,N_8244);
nor U19275 (N_19275,N_3003,N_5875);
nor U19276 (N_19276,N_2056,N_7037);
nor U19277 (N_19277,N_9190,N_2215);
nand U19278 (N_19278,N_7128,N_9452);
xor U19279 (N_19279,N_9148,N_6969);
and U19280 (N_19280,N_5362,N_5928);
nor U19281 (N_19281,N_1118,N_6491);
or U19282 (N_19282,N_5350,N_622);
and U19283 (N_19283,N_4008,N_1636);
or U19284 (N_19284,N_878,N_7161);
nor U19285 (N_19285,N_2578,N_5328);
xor U19286 (N_19286,N_9981,N_7361);
or U19287 (N_19287,N_6362,N_2937);
xor U19288 (N_19288,N_9207,N_2822);
or U19289 (N_19289,N_4244,N_855);
nand U19290 (N_19290,N_5251,N_9829);
and U19291 (N_19291,N_8192,N_6159);
and U19292 (N_19292,N_2253,N_2208);
nand U19293 (N_19293,N_4632,N_6276);
and U19294 (N_19294,N_7416,N_4589);
nor U19295 (N_19295,N_2595,N_64);
nand U19296 (N_19296,N_2078,N_9732);
or U19297 (N_19297,N_8450,N_4661);
or U19298 (N_19298,N_2321,N_6176);
nand U19299 (N_19299,N_6753,N_2906);
nor U19300 (N_19300,N_4242,N_6997);
or U19301 (N_19301,N_5619,N_6672);
xnor U19302 (N_19302,N_3755,N_3723);
and U19303 (N_19303,N_5546,N_6411);
nor U19304 (N_19304,N_5834,N_9218);
xor U19305 (N_19305,N_6931,N_583);
nand U19306 (N_19306,N_7404,N_1744);
and U19307 (N_19307,N_2013,N_8458);
or U19308 (N_19308,N_8545,N_140);
xor U19309 (N_19309,N_5790,N_6376);
or U19310 (N_19310,N_4873,N_6383);
and U19311 (N_19311,N_6573,N_3675);
or U19312 (N_19312,N_4809,N_518);
or U19313 (N_19313,N_7636,N_155);
and U19314 (N_19314,N_6341,N_1983);
xnor U19315 (N_19315,N_4968,N_1781);
nand U19316 (N_19316,N_4793,N_6833);
or U19317 (N_19317,N_6715,N_4109);
nor U19318 (N_19318,N_3264,N_1610);
nor U19319 (N_19319,N_1975,N_1942);
nand U19320 (N_19320,N_9402,N_9334);
or U19321 (N_19321,N_5,N_8697);
or U19322 (N_19322,N_6262,N_8949);
nand U19323 (N_19323,N_905,N_4350);
nor U19324 (N_19324,N_5827,N_100);
nand U19325 (N_19325,N_3574,N_7233);
xor U19326 (N_19326,N_731,N_3051);
nand U19327 (N_19327,N_3281,N_1674);
nand U19328 (N_19328,N_7675,N_930);
and U19329 (N_19329,N_8690,N_49);
and U19330 (N_19330,N_5083,N_9259);
and U19331 (N_19331,N_1610,N_9659);
nor U19332 (N_19332,N_8339,N_9856);
or U19333 (N_19333,N_946,N_6157);
or U19334 (N_19334,N_5863,N_1956);
xnor U19335 (N_19335,N_5307,N_3836);
xor U19336 (N_19336,N_9274,N_4753);
and U19337 (N_19337,N_2533,N_5775);
and U19338 (N_19338,N_2601,N_8069);
and U19339 (N_19339,N_3199,N_8708);
nand U19340 (N_19340,N_8373,N_8397);
xor U19341 (N_19341,N_2289,N_5863);
nand U19342 (N_19342,N_7802,N_9472);
nand U19343 (N_19343,N_2,N_4348);
nor U19344 (N_19344,N_8299,N_657);
or U19345 (N_19345,N_3340,N_278);
nand U19346 (N_19346,N_744,N_7471);
nor U19347 (N_19347,N_7478,N_2577);
xnor U19348 (N_19348,N_9321,N_4957);
or U19349 (N_19349,N_6117,N_2484);
nand U19350 (N_19350,N_8291,N_5584);
xnor U19351 (N_19351,N_5441,N_574);
nor U19352 (N_19352,N_9837,N_7166);
xnor U19353 (N_19353,N_6194,N_8232);
and U19354 (N_19354,N_1793,N_2380);
nor U19355 (N_19355,N_1404,N_6728);
nand U19356 (N_19356,N_7233,N_4525);
or U19357 (N_19357,N_3803,N_201);
nor U19358 (N_19358,N_2955,N_5544);
and U19359 (N_19359,N_1052,N_4498);
nor U19360 (N_19360,N_7811,N_9382);
and U19361 (N_19361,N_7155,N_7178);
nor U19362 (N_19362,N_1640,N_5531);
nor U19363 (N_19363,N_9059,N_9894);
and U19364 (N_19364,N_9183,N_2060);
nor U19365 (N_19365,N_2464,N_5918);
and U19366 (N_19366,N_7390,N_4681);
or U19367 (N_19367,N_2866,N_8076);
xnor U19368 (N_19368,N_2157,N_5061);
nor U19369 (N_19369,N_3883,N_8188);
xnor U19370 (N_19370,N_1158,N_7645);
or U19371 (N_19371,N_8975,N_443);
and U19372 (N_19372,N_2247,N_2959);
and U19373 (N_19373,N_9538,N_2596);
nand U19374 (N_19374,N_1421,N_3794);
nand U19375 (N_19375,N_1720,N_6541);
nor U19376 (N_19376,N_8036,N_4800);
and U19377 (N_19377,N_8374,N_2076);
nand U19378 (N_19378,N_8759,N_5529);
nor U19379 (N_19379,N_494,N_6373);
nand U19380 (N_19380,N_5156,N_7155);
and U19381 (N_19381,N_9898,N_4631);
and U19382 (N_19382,N_3884,N_3181);
and U19383 (N_19383,N_2493,N_7935);
nand U19384 (N_19384,N_2254,N_9078);
nand U19385 (N_19385,N_6999,N_8215);
or U19386 (N_19386,N_7134,N_8755);
xor U19387 (N_19387,N_3703,N_6628);
and U19388 (N_19388,N_1648,N_4955);
nand U19389 (N_19389,N_3180,N_3451);
and U19390 (N_19390,N_2260,N_192);
nor U19391 (N_19391,N_5507,N_2769);
and U19392 (N_19392,N_6800,N_4720);
and U19393 (N_19393,N_2184,N_1028);
or U19394 (N_19394,N_5430,N_3088);
xnor U19395 (N_19395,N_3517,N_1415);
nor U19396 (N_19396,N_845,N_1767);
nand U19397 (N_19397,N_1851,N_1241);
xnor U19398 (N_19398,N_1554,N_4783);
nor U19399 (N_19399,N_1271,N_9774);
nor U19400 (N_19400,N_4636,N_4586);
nor U19401 (N_19401,N_6293,N_141);
and U19402 (N_19402,N_3405,N_712);
nor U19403 (N_19403,N_6741,N_2651);
nor U19404 (N_19404,N_3904,N_4234);
nand U19405 (N_19405,N_8313,N_1550);
nand U19406 (N_19406,N_3583,N_1072);
and U19407 (N_19407,N_1005,N_4160);
and U19408 (N_19408,N_4504,N_8997);
nand U19409 (N_19409,N_8102,N_7625);
and U19410 (N_19410,N_3435,N_6103);
or U19411 (N_19411,N_178,N_2738);
or U19412 (N_19412,N_5151,N_6470);
nand U19413 (N_19413,N_5038,N_7712);
nand U19414 (N_19414,N_9081,N_1724);
xor U19415 (N_19415,N_4377,N_637);
and U19416 (N_19416,N_4409,N_1629);
or U19417 (N_19417,N_4718,N_1433);
nand U19418 (N_19418,N_7287,N_5068);
nor U19419 (N_19419,N_4898,N_5250);
nor U19420 (N_19420,N_2541,N_5369);
xnor U19421 (N_19421,N_8710,N_9100);
nor U19422 (N_19422,N_2068,N_5481);
xor U19423 (N_19423,N_4066,N_9221);
nand U19424 (N_19424,N_852,N_5772);
xnor U19425 (N_19425,N_5247,N_176);
nand U19426 (N_19426,N_4925,N_4409);
or U19427 (N_19427,N_6479,N_4851);
nor U19428 (N_19428,N_3035,N_5613);
and U19429 (N_19429,N_2377,N_9069);
nor U19430 (N_19430,N_1764,N_1274);
or U19431 (N_19431,N_1337,N_821);
and U19432 (N_19432,N_2370,N_1254);
nand U19433 (N_19433,N_9595,N_3097);
nand U19434 (N_19434,N_9999,N_55);
nor U19435 (N_19435,N_1222,N_6683);
nor U19436 (N_19436,N_3982,N_6213);
or U19437 (N_19437,N_7464,N_1097);
xnor U19438 (N_19438,N_7593,N_350);
or U19439 (N_19439,N_3804,N_1208);
xor U19440 (N_19440,N_6210,N_7896);
nor U19441 (N_19441,N_1398,N_705);
nor U19442 (N_19442,N_5987,N_746);
or U19443 (N_19443,N_2803,N_642);
xnor U19444 (N_19444,N_2895,N_5163);
xor U19445 (N_19445,N_7632,N_9693);
or U19446 (N_19446,N_1015,N_6740);
nand U19447 (N_19447,N_7194,N_2350);
nand U19448 (N_19448,N_6187,N_8298);
nor U19449 (N_19449,N_1754,N_9476);
nor U19450 (N_19450,N_635,N_8996);
and U19451 (N_19451,N_9237,N_802);
nor U19452 (N_19452,N_114,N_1320);
and U19453 (N_19453,N_586,N_2144);
nor U19454 (N_19454,N_9534,N_7692);
and U19455 (N_19455,N_7734,N_1327);
nand U19456 (N_19456,N_6324,N_2599);
xor U19457 (N_19457,N_8475,N_3397);
nor U19458 (N_19458,N_2397,N_3784);
nor U19459 (N_19459,N_1282,N_1853);
nor U19460 (N_19460,N_5191,N_4745);
nor U19461 (N_19461,N_4324,N_4739);
nand U19462 (N_19462,N_8105,N_9172);
nand U19463 (N_19463,N_7222,N_282);
or U19464 (N_19464,N_1058,N_8066);
xor U19465 (N_19465,N_9503,N_7521);
xor U19466 (N_19466,N_2815,N_8137);
nand U19467 (N_19467,N_918,N_8945);
nand U19468 (N_19468,N_3786,N_6997);
or U19469 (N_19469,N_1041,N_5961);
nor U19470 (N_19470,N_2019,N_9098);
xnor U19471 (N_19471,N_2288,N_5386);
and U19472 (N_19472,N_5129,N_3151);
or U19473 (N_19473,N_2728,N_5039);
nand U19474 (N_19474,N_6059,N_9400);
nand U19475 (N_19475,N_3489,N_9573);
xor U19476 (N_19476,N_7981,N_8585);
nor U19477 (N_19477,N_6218,N_4957);
xor U19478 (N_19478,N_8560,N_7581);
nand U19479 (N_19479,N_7003,N_1184);
xnor U19480 (N_19480,N_4110,N_5144);
and U19481 (N_19481,N_6231,N_2729);
and U19482 (N_19482,N_3422,N_6266);
and U19483 (N_19483,N_1128,N_9113);
nor U19484 (N_19484,N_6664,N_566);
nor U19485 (N_19485,N_690,N_6609);
and U19486 (N_19486,N_1504,N_5487);
or U19487 (N_19487,N_3521,N_9006);
xor U19488 (N_19488,N_1854,N_9023);
or U19489 (N_19489,N_8919,N_6353);
nand U19490 (N_19490,N_1440,N_1077);
or U19491 (N_19491,N_3120,N_6417);
or U19492 (N_19492,N_7448,N_5692);
or U19493 (N_19493,N_6369,N_763);
and U19494 (N_19494,N_1872,N_577);
or U19495 (N_19495,N_2524,N_3726);
nor U19496 (N_19496,N_8970,N_7260);
nor U19497 (N_19497,N_9905,N_9676);
nor U19498 (N_19498,N_2016,N_4734);
and U19499 (N_19499,N_9823,N_4268);
xnor U19500 (N_19500,N_2579,N_7774);
or U19501 (N_19501,N_1228,N_1488);
xor U19502 (N_19502,N_3891,N_2636);
nand U19503 (N_19503,N_5934,N_4300);
nor U19504 (N_19504,N_8538,N_3707);
xor U19505 (N_19505,N_8788,N_7226);
nand U19506 (N_19506,N_7225,N_9867);
nor U19507 (N_19507,N_2910,N_1810);
nand U19508 (N_19508,N_9026,N_2487);
or U19509 (N_19509,N_9495,N_2420);
xor U19510 (N_19510,N_2699,N_4144);
nor U19511 (N_19511,N_34,N_671);
nor U19512 (N_19512,N_6456,N_9963);
nor U19513 (N_19513,N_5755,N_8397);
nand U19514 (N_19514,N_9919,N_3180);
nand U19515 (N_19515,N_6294,N_1204);
nand U19516 (N_19516,N_7973,N_8474);
xnor U19517 (N_19517,N_4876,N_4573);
nand U19518 (N_19518,N_4177,N_6913);
nand U19519 (N_19519,N_5709,N_4224);
and U19520 (N_19520,N_1489,N_2591);
xnor U19521 (N_19521,N_2194,N_2669);
nor U19522 (N_19522,N_492,N_9661);
nor U19523 (N_19523,N_6704,N_1008);
nor U19524 (N_19524,N_9175,N_9319);
nor U19525 (N_19525,N_3301,N_1768);
and U19526 (N_19526,N_3523,N_1675);
nand U19527 (N_19527,N_3428,N_5959);
nand U19528 (N_19528,N_3981,N_2352);
and U19529 (N_19529,N_8615,N_2967);
nand U19530 (N_19530,N_5123,N_6183);
xnor U19531 (N_19531,N_6113,N_4351);
or U19532 (N_19532,N_5281,N_1223);
nor U19533 (N_19533,N_6968,N_941);
nand U19534 (N_19534,N_1429,N_2173);
and U19535 (N_19535,N_8897,N_1873);
and U19536 (N_19536,N_849,N_6968);
or U19537 (N_19537,N_5862,N_4133);
nand U19538 (N_19538,N_9078,N_9010);
nand U19539 (N_19539,N_746,N_5514);
nor U19540 (N_19540,N_7870,N_7355);
and U19541 (N_19541,N_1193,N_2937);
or U19542 (N_19542,N_5761,N_6037);
and U19543 (N_19543,N_6418,N_7042);
and U19544 (N_19544,N_2285,N_1552);
xor U19545 (N_19545,N_4192,N_3186);
or U19546 (N_19546,N_7728,N_5379);
or U19547 (N_19547,N_772,N_6109);
and U19548 (N_19548,N_8993,N_159);
nor U19549 (N_19549,N_2744,N_4717);
xor U19550 (N_19550,N_6233,N_9624);
nand U19551 (N_19551,N_4551,N_2410);
nor U19552 (N_19552,N_7190,N_6748);
nor U19553 (N_19553,N_3151,N_2060);
and U19554 (N_19554,N_3673,N_1497);
xor U19555 (N_19555,N_5747,N_4971);
xor U19556 (N_19556,N_89,N_9373);
nor U19557 (N_19557,N_5791,N_8425);
nor U19558 (N_19558,N_8203,N_8012);
nor U19559 (N_19559,N_9508,N_6199);
nor U19560 (N_19560,N_2528,N_8588);
nand U19561 (N_19561,N_3071,N_6026);
or U19562 (N_19562,N_8731,N_2267);
xor U19563 (N_19563,N_4205,N_7880);
nand U19564 (N_19564,N_226,N_5847);
and U19565 (N_19565,N_2364,N_1765);
nor U19566 (N_19566,N_8558,N_5326);
or U19567 (N_19567,N_1767,N_6465);
and U19568 (N_19568,N_5460,N_6380);
and U19569 (N_19569,N_6896,N_1284);
or U19570 (N_19570,N_1188,N_4727);
nand U19571 (N_19571,N_9722,N_6602);
or U19572 (N_19572,N_9069,N_9663);
and U19573 (N_19573,N_7709,N_3649);
nor U19574 (N_19574,N_7084,N_4755);
and U19575 (N_19575,N_3120,N_5775);
and U19576 (N_19576,N_7768,N_5463);
or U19577 (N_19577,N_7827,N_2934);
nand U19578 (N_19578,N_3197,N_2968);
nand U19579 (N_19579,N_7352,N_1538);
or U19580 (N_19580,N_8580,N_1277);
or U19581 (N_19581,N_1838,N_9039);
or U19582 (N_19582,N_558,N_9594);
nand U19583 (N_19583,N_3520,N_9699);
nor U19584 (N_19584,N_5999,N_5575);
nor U19585 (N_19585,N_2287,N_4124);
xor U19586 (N_19586,N_5674,N_5420);
or U19587 (N_19587,N_8180,N_8710);
nor U19588 (N_19588,N_2152,N_5808);
xor U19589 (N_19589,N_8602,N_8018);
or U19590 (N_19590,N_9038,N_7775);
nand U19591 (N_19591,N_4945,N_8294);
nor U19592 (N_19592,N_5741,N_3070);
xnor U19593 (N_19593,N_3832,N_4958);
xnor U19594 (N_19594,N_5385,N_9556);
and U19595 (N_19595,N_1600,N_2261);
xnor U19596 (N_19596,N_1502,N_1975);
nor U19597 (N_19597,N_2758,N_9870);
or U19598 (N_19598,N_1171,N_8949);
or U19599 (N_19599,N_5579,N_7093);
nor U19600 (N_19600,N_3868,N_6505);
nand U19601 (N_19601,N_1883,N_2579);
xnor U19602 (N_19602,N_9138,N_1056);
xor U19603 (N_19603,N_7468,N_4874);
nor U19604 (N_19604,N_1847,N_2598);
or U19605 (N_19605,N_6704,N_1731);
nor U19606 (N_19606,N_6401,N_4773);
or U19607 (N_19607,N_418,N_1726);
nor U19608 (N_19608,N_9890,N_9445);
nand U19609 (N_19609,N_7990,N_1206);
nand U19610 (N_19610,N_4784,N_5602);
and U19611 (N_19611,N_7747,N_8508);
xnor U19612 (N_19612,N_9894,N_2858);
nor U19613 (N_19613,N_7710,N_9062);
and U19614 (N_19614,N_3858,N_8799);
nand U19615 (N_19615,N_3520,N_8844);
nor U19616 (N_19616,N_8059,N_3324);
xor U19617 (N_19617,N_261,N_7683);
or U19618 (N_19618,N_3524,N_5515);
and U19619 (N_19619,N_7695,N_816);
nand U19620 (N_19620,N_2139,N_6749);
xnor U19621 (N_19621,N_4933,N_6844);
nor U19622 (N_19622,N_3379,N_5089);
or U19623 (N_19623,N_5330,N_7479);
nor U19624 (N_19624,N_5934,N_4784);
xor U19625 (N_19625,N_3383,N_3982);
xnor U19626 (N_19626,N_1053,N_685);
nor U19627 (N_19627,N_3136,N_8339);
nand U19628 (N_19628,N_3402,N_4224);
nor U19629 (N_19629,N_3691,N_7454);
or U19630 (N_19630,N_1846,N_8860);
xnor U19631 (N_19631,N_5283,N_8435);
or U19632 (N_19632,N_9109,N_2780);
nor U19633 (N_19633,N_5755,N_2355);
or U19634 (N_19634,N_4679,N_3712);
nand U19635 (N_19635,N_462,N_4989);
nand U19636 (N_19636,N_5179,N_3501);
and U19637 (N_19637,N_1820,N_4137);
and U19638 (N_19638,N_6048,N_5659);
and U19639 (N_19639,N_3389,N_5476);
and U19640 (N_19640,N_8357,N_7169);
nor U19641 (N_19641,N_7273,N_8642);
nand U19642 (N_19642,N_5229,N_5559);
xnor U19643 (N_19643,N_3402,N_2134);
or U19644 (N_19644,N_7338,N_6398);
or U19645 (N_19645,N_4027,N_222);
xor U19646 (N_19646,N_4505,N_9730);
nand U19647 (N_19647,N_1474,N_1713);
nor U19648 (N_19648,N_9928,N_9483);
or U19649 (N_19649,N_7710,N_103);
and U19650 (N_19650,N_1732,N_3581);
and U19651 (N_19651,N_2362,N_553);
nand U19652 (N_19652,N_2885,N_5359);
nand U19653 (N_19653,N_2326,N_7997);
nor U19654 (N_19654,N_1963,N_178);
nand U19655 (N_19655,N_9603,N_3118);
xnor U19656 (N_19656,N_7154,N_9882);
nand U19657 (N_19657,N_9329,N_1030);
xnor U19658 (N_19658,N_4088,N_6059);
xor U19659 (N_19659,N_2885,N_3151);
xor U19660 (N_19660,N_8196,N_4725);
nor U19661 (N_19661,N_7729,N_2645);
and U19662 (N_19662,N_1578,N_2046);
nand U19663 (N_19663,N_7503,N_2045);
nor U19664 (N_19664,N_8540,N_2933);
xor U19665 (N_19665,N_7105,N_5785);
and U19666 (N_19666,N_7672,N_8661);
or U19667 (N_19667,N_2149,N_9668);
nand U19668 (N_19668,N_8084,N_597);
nand U19669 (N_19669,N_730,N_45);
or U19670 (N_19670,N_1963,N_1427);
and U19671 (N_19671,N_9649,N_1358);
xor U19672 (N_19672,N_4047,N_6217);
nor U19673 (N_19673,N_7231,N_6417);
xor U19674 (N_19674,N_3690,N_9106);
xnor U19675 (N_19675,N_5305,N_44);
nand U19676 (N_19676,N_8327,N_7037);
and U19677 (N_19677,N_3021,N_9559);
nor U19678 (N_19678,N_7855,N_9982);
nor U19679 (N_19679,N_1819,N_9278);
and U19680 (N_19680,N_3749,N_9646);
xor U19681 (N_19681,N_6950,N_755);
and U19682 (N_19682,N_8308,N_411);
or U19683 (N_19683,N_530,N_9360);
xor U19684 (N_19684,N_2694,N_9513);
and U19685 (N_19685,N_9766,N_599);
and U19686 (N_19686,N_8712,N_422);
nand U19687 (N_19687,N_8159,N_2271);
and U19688 (N_19688,N_3872,N_5957);
and U19689 (N_19689,N_5860,N_4036);
nor U19690 (N_19690,N_142,N_6743);
or U19691 (N_19691,N_6588,N_2504);
and U19692 (N_19692,N_7907,N_2123);
xor U19693 (N_19693,N_3053,N_7721);
or U19694 (N_19694,N_5810,N_1585);
or U19695 (N_19695,N_7608,N_6699);
xor U19696 (N_19696,N_5873,N_7267);
nand U19697 (N_19697,N_8516,N_6487);
nor U19698 (N_19698,N_4751,N_3104);
and U19699 (N_19699,N_6409,N_9384);
nor U19700 (N_19700,N_3815,N_9562);
xor U19701 (N_19701,N_4625,N_4395);
or U19702 (N_19702,N_6827,N_298);
xor U19703 (N_19703,N_5862,N_1563);
xor U19704 (N_19704,N_4795,N_1386);
nand U19705 (N_19705,N_8373,N_5410);
nor U19706 (N_19706,N_3282,N_7423);
nor U19707 (N_19707,N_6336,N_1480);
or U19708 (N_19708,N_8333,N_9250);
nor U19709 (N_19709,N_2143,N_3248);
or U19710 (N_19710,N_6028,N_9513);
or U19711 (N_19711,N_9444,N_4686);
nor U19712 (N_19712,N_2274,N_208);
and U19713 (N_19713,N_7040,N_5039);
xnor U19714 (N_19714,N_888,N_8891);
nand U19715 (N_19715,N_816,N_8178);
nor U19716 (N_19716,N_9803,N_1994);
or U19717 (N_19717,N_9826,N_9515);
nand U19718 (N_19718,N_6717,N_952);
nand U19719 (N_19719,N_5903,N_2881);
or U19720 (N_19720,N_4087,N_3981);
or U19721 (N_19721,N_588,N_4812);
nor U19722 (N_19722,N_2677,N_9998);
nand U19723 (N_19723,N_8120,N_5483);
or U19724 (N_19724,N_5536,N_8061);
and U19725 (N_19725,N_7662,N_399);
or U19726 (N_19726,N_8845,N_692);
nor U19727 (N_19727,N_1473,N_311);
or U19728 (N_19728,N_1507,N_6113);
xnor U19729 (N_19729,N_8767,N_9801);
or U19730 (N_19730,N_8314,N_8653);
xor U19731 (N_19731,N_7568,N_874);
or U19732 (N_19732,N_5575,N_76);
xor U19733 (N_19733,N_3894,N_7146);
nor U19734 (N_19734,N_109,N_5280);
or U19735 (N_19735,N_1321,N_7658);
nor U19736 (N_19736,N_5389,N_4019);
nand U19737 (N_19737,N_1567,N_1040);
or U19738 (N_19738,N_4175,N_8863);
xor U19739 (N_19739,N_2169,N_600);
and U19740 (N_19740,N_9033,N_6055);
nor U19741 (N_19741,N_8183,N_5476);
nor U19742 (N_19742,N_8223,N_2144);
and U19743 (N_19743,N_210,N_9385);
nor U19744 (N_19744,N_3223,N_4011);
nand U19745 (N_19745,N_3948,N_4402);
or U19746 (N_19746,N_9105,N_5958);
or U19747 (N_19747,N_5728,N_6330);
nor U19748 (N_19748,N_6385,N_920);
and U19749 (N_19749,N_5065,N_86);
nand U19750 (N_19750,N_9240,N_7448);
nand U19751 (N_19751,N_9704,N_5525);
and U19752 (N_19752,N_9669,N_6877);
nor U19753 (N_19753,N_6437,N_7232);
xnor U19754 (N_19754,N_2265,N_4464);
and U19755 (N_19755,N_8705,N_5973);
xnor U19756 (N_19756,N_3083,N_1588);
nor U19757 (N_19757,N_3944,N_2304);
and U19758 (N_19758,N_3801,N_9690);
and U19759 (N_19759,N_6262,N_7911);
and U19760 (N_19760,N_2080,N_6625);
and U19761 (N_19761,N_6337,N_2253);
or U19762 (N_19762,N_6075,N_3454);
or U19763 (N_19763,N_4187,N_1005);
and U19764 (N_19764,N_5768,N_617);
xor U19765 (N_19765,N_8030,N_4050);
or U19766 (N_19766,N_4624,N_5538);
nor U19767 (N_19767,N_1070,N_2471);
nand U19768 (N_19768,N_7737,N_887);
and U19769 (N_19769,N_1436,N_3342);
nor U19770 (N_19770,N_3398,N_7557);
nand U19771 (N_19771,N_4113,N_9613);
or U19772 (N_19772,N_7134,N_6446);
or U19773 (N_19773,N_2513,N_9514);
nand U19774 (N_19774,N_2694,N_8366);
and U19775 (N_19775,N_9384,N_2108);
xnor U19776 (N_19776,N_6712,N_3947);
nor U19777 (N_19777,N_8034,N_6345);
or U19778 (N_19778,N_3999,N_9988);
or U19779 (N_19779,N_9018,N_41);
and U19780 (N_19780,N_3378,N_6914);
nor U19781 (N_19781,N_6741,N_2673);
nor U19782 (N_19782,N_8596,N_9586);
xnor U19783 (N_19783,N_2191,N_2179);
and U19784 (N_19784,N_2869,N_866);
xnor U19785 (N_19785,N_9900,N_1340);
nand U19786 (N_19786,N_293,N_7480);
nand U19787 (N_19787,N_9548,N_2890);
nand U19788 (N_19788,N_3470,N_4517);
nor U19789 (N_19789,N_4327,N_1509);
nor U19790 (N_19790,N_4701,N_7050);
or U19791 (N_19791,N_9157,N_9643);
nand U19792 (N_19792,N_1871,N_7628);
xnor U19793 (N_19793,N_8230,N_93);
nand U19794 (N_19794,N_8729,N_5256);
nor U19795 (N_19795,N_3810,N_1673);
or U19796 (N_19796,N_8220,N_434);
nor U19797 (N_19797,N_1482,N_6190);
nand U19798 (N_19798,N_8151,N_5755);
nand U19799 (N_19799,N_4801,N_7612);
nor U19800 (N_19800,N_4881,N_2974);
xnor U19801 (N_19801,N_4513,N_882);
nand U19802 (N_19802,N_2241,N_3622);
xnor U19803 (N_19803,N_4797,N_3271);
nor U19804 (N_19804,N_9791,N_6600);
or U19805 (N_19805,N_8275,N_9630);
and U19806 (N_19806,N_1017,N_2983);
nand U19807 (N_19807,N_9474,N_8781);
nand U19808 (N_19808,N_4327,N_7611);
nand U19809 (N_19809,N_3318,N_7535);
and U19810 (N_19810,N_6024,N_3113);
nand U19811 (N_19811,N_4586,N_936);
and U19812 (N_19812,N_3995,N_4785);
nor U19813 (N_19813,N_4419,N_7773);
or U19814 (N_19814,N_1305,N_9512);
xor U19815 (N_19815,N_2035,N_253);
xor U19816 (N_19816,N_9296,N_4871);
nand U19817 (N_19817,N_8805,N_6343);
xnor U19818 (N_19818,N_8257,N_9903);
or U19819 (N_19819,N_3369,N_6307);
nor U19820 (N_19820,N_2681,N_8164);
nand U19821 (N_19821,N_8850,N_2438);
xnor U19822 (N_19822,N_536,N_9268);
xor U19823 (N_19823,N_579,N_7117);
nor U19824 (N_19824,N_180,N_8587);
nor U19825 (N_19825,N_459,N_5949);
nand U19826 (N_19826,N_8590,N_8820);
nand U19827 (N_19827,N_5521,N_8868);
xor U19828 (N_19828,N_6915,N_7058);
and U19829 (N_19829,N_8552,N_4928);
nand U19830 (N_19830,N_5439,N_2839);
and U19831 (N_19831,N_2463,N_4671);
and U19832 (N_19832,N_8619,N_4015);
or U19833 (N_19833,N_3259,N_7851);
xor U19834 (N_19834,N_5219,N_8604);
nor U19835 (N_19835,N_3410,N_4418);
or U19836 (N_19836,N_7266,N_7892);
or U19837 (N_19837,N_6724,N_840);
and U19838 (N_19838,N_1328,N_5700);
nor U19839 (N_19839,N_4311,N_9606);
xor U19840 (N_19840,N_4290,N_9117);
and U19841 (N_19841,N_474,N_6643);
and U19842 (N_19842,N_7956,N_8885);
xor U19843 (N_19843,N_2976,N_9870);
xor U19844 (N_19844,N_8398,N_3331);
nand U19845 (N_19845,N_8908,N_7892);
nand U19846 (N_19846,N_3994,N_9940);
and U19847 (N_19847,N_4043,N_2011);
or U19848 (N_19848,N_5952,N_9766);
and U19849 (N_19849,N_1572,N_2934);
nand U19850 (N_19850,N_5844,N_4164);
and U19851 (N_19851,N_9992,N_9453);
nor U19852 (N_19852,N_8196,N_9208);
nor U19853 (N_19853,N_6244,N_9739);
xor U19854 (N_19854,N_6482,N_4718);
nand U19855 (N_19855,N_2005,N_312);
nand U19856 (N_19856,N_642,N_2537);
nand U19857 (N_19857,N_6524,N_1166);
and U19858 (N_19858,N_6547,N_7842);
and U19859 (N_19859,N_8299,N_2446);
or U19860 (N_19860,N_9061,N_136);
nor U19861 (N_19861,N_1003,N_3526);
nand U19862 (N_19862,N_3845,N_6923);
xor U19863 (N_19863,N_2479,N_1994);
or U19864 (N_19864,N_7899,N_402);
nand U19865 (N_19865,N_7925,N_8322);
or U19866 (N_19866,N_2835,N_8902);
nand U19867 (N_19867,N_2574,N_7357);
xnor U19868 (N_19868,N_2004,N_8273);
or U19869 (N_19869,N_3049,N_6034);
xor U19870 (N_19870,N_4515,N_1815);
and U19871 (N_19871,N_1313,N_8658);
xnor U19872 (N_19872,N_4114,N_1305);
and U19873 (N_19873,N_9583,N_8440);
or U19874 (N_19874,N_8452,N_7539);
xnor U19875 (N_19875,N_6326,N_3120);
or U19876 (N_19876,N_4387,N_8746);
or U19877 (N_19877,N_6246,N_8204);
or U19878 (N_19878,N_180,N_7112);
or U19879 (N_19879,N_511,N_7667);
nand U19880 (N_19880,N_7309,N_5879);
or U19881 (N_19881,N_7196,N_6735);
xor U19882 (N_19882,N_3698,N_7055);
nor U19883 (N_19883,N_2148,N_5039);
nand U19884 (N_19884,N_8247,N_3012);
xnor U19885 (N_19885,N_2208,N_7738);
or U19886 (N_19886,N_2345,N_557);
and U19887 (N_19887,N_4952,N_3510);
nor U19888 (N_19888,N_3157,N_7543);
or U19889 (N_19889,N_862,N_7849);
and U19890 (N_19890,N_2730,N_738);
and U19891 (N_19891,N_3863,N_2178);
and U19892 (N_19892,N_8672,N_5542);
or U19893 (N_19893,N_2992,N_9932);
nand U19894 (N_19894,N_1888,N_4711);
and U19895 (N_19895,N_3301,N_9159);
or U19896 (N_19896,N_2155,N_7074);
nor U19897 (N_19897,N_1076,N_5762);
or U19898 (N_19898,N_2168,N_2051);
xnor U19899 (N_19899,N_2208,N_7871);
nor U19900 (N_19900,N_4757,N_2906);
or U19901 (N_19901,N_7859,N_9022);
xnor U19902 (N_19902,N_1850,N_3733);
or U19903 (N_19903,N_8055,N_5989);
or U19904 (N_19904,N_2223,N_4663);
and U19905 (N_19905,N_5871,N_8148);
or U19906 (N_19906,N_2819,N_1141);
or U19907 (N_19907,N_8522,N_6850);
xor U19908 (N_19908,N_9564,N_1854);
nor U19909 (N_19909,N_9791,N_7897);
xnor U19910 (N_19910,N_6857,N_2006);
nand U19911 (N_19911,N_8166,N_6768);
xor U19912 (N_19912,N_1954,N_590);
nor U19913 (N_19913,N_2412,N_7398);
nand U19914 (N_19914,N_1987,N_8658);
and U19915 (N_19915,N_6313,N_678);
or U19916 (N_19916,N_55,N_1617);
xor U19917 (N_19917,N_3586,N_1077);
or U19918 (N_19918,N_9693,N_4136);
nand U19919 (N_19919,N_2024,N_346);
and U19920 (N_19920,N_1479,N_8149);
nand U19921 (N_19921,N_1920,N_9260);
xnor U19922 (N_19922,N_8731,N_5402);
or U19923 (N_19923,N_1330,N_6528);
xnor U19924 (N_19924,N_4044,N_6713);
nand U19925 (N_19925,N_4424,N_698);
xnor U19926 (N_19926,N_3819,N_9866);
nand U19927 (N_19927,N_1858,N_2589);
nand U19928 (N_19928,N_2880,N_6516);
nand U19929 (N_19929,N_1120,N_5688);
nand U19930 (N_19930,N_758,N_969);
or U19931 (N_19931,N_4252,N_8880);
nor U19932 (N_19932,N_5885,N_8143);
xnor U19933 (N_19933,N_5181,N_8906);
nor U19934 (N_19934,N_5137,N_4995);
and U19935 (N_19935,N_9877,N_5777);
or U19936 (N_19936,N_9658,N_1693);
xnor U19937 (N_19937,N_2875,N_8264);
and U19938 (N_19938,N_6905,N_5533);
xor U19939 (N_19939,N_7522,N_6749);
or U19940 (N_19940,N_5780,N_6509);
xor U19941 (N_19941,N_2736,N_2253);
nand U19942 (N_19942,N_4644,N_5213);
nor U19943 (N_19943,N_2768,N_9428);
nand U19944 (N_19944,N_2826,N_7100);
and U19945 (N_19945,N_5005,N_9837);
and U19946 (N_19946,N_2473,N_5318);
nand U19947 (N_19947,N_8986,N_2708);
and U19948 (N_19948,N_7043,N_7737);
xnor U19949 (N_19949,N_216,N_9578);
nand U19950 (N_19950,N_1094,N_217);
and U19951 (N_19951,N_5482,N_3645);
nor U19952 (N_19952,N_1074,N_9521);
nor U19953 (N_19953,N_3204,N_2346);
and U19954 (N_19954,N_2538,N_8117);
nand U19955 (N_19955,N_9144,N_2883);
and U19956 (N_19956,N_7493,N_6537);
and U19957 (N_19957,N_6355,N_1358);
nor U19958 (N_19958,N_5592,N_4101);
nor U19959 (N_19959,N_8936,N_917);
xnor U19960 (N_19960,N_657,N_8135);
xor U19961 (N_19961,N_615,N_8539);
xnor U19962 (N_19962,N_4413,N_299);
and U19963 (N_19963,N_504,N_8919);
nand U19964 (N_19964,N_1238,N_6820);
nand U19965 (N_19965,N_9790,N_3932);
nand U19966 (N_19966,N_7799,N_9205);
xnor U19967 (N_19967,N_8321,N_1885);
nor U19968 (N_19968,N_1096,N_143);
nand U19969 (N_19969,N_3575,N_3544);
nand U19970 (N_19970,N_9060,N_1786);
xor U19971 (N_19971,N_3734,N_5102);
or U19972 (N_19972,N_4683,N_5510);
xnor U19973 (N_19973,N_519,N_4512);
nand U19974 (N_19974,N_1133,N_3962);
nor U19975 (N_19975,N_7080,N_6450);
nor U19976 (N_19976,N_7504,N_8860);
xnor U19977 (N_19977,N_1959,N_3239);
nand U19978 (N_19978,N_3909,N_4202);
nor U19979 (N_19979,N_2324,N_8470);
and U19980 (N_19980,N_956,N_5389);
xor U19981 (N_19981,N_3021,N_487);
nor U19982 (N_19982,N_8393,N_6457);
and U19983 (N_19983,N_2194,N_7751);
nand U19984 (N_19984,N_9819,N_9970);
xnor U19985 (N_19985,N_5675,N_2858);
xnor U19986 (N_19986,N_932,N_4707);
nor U19987 (N_19987,N_3268,N_7891);
nor U19988 (N_19988,N_8683,N_6837);
nand U19989 (N_19989,N_9257,N_6887);
nand U19990 (N_19990,N_9493,N_3750);
xnor U19991 (N_19991,N_7944,N_5407);
or U19992 (N_19992,N_1407,N_6640);
and U19993 (N_19993,N_673,N_6982);
nand U19994 (N_19994,N_476,N_3587);
nand U19995 (N_19995,N_5788,N_2759);
or U19996 (N_19996,N_8790,N_262);
xor U19997 (N_19997,N_9196,N_6083);
or U19998 (N_19998,N_191,N_5745);
nor U19999 (N_19999,N_9245,N_2741);
nor U20000 (N_20000,N_18348,N_11096);
xor U20001 (N_20001,N_11117,N_11597);
nand U20002 (N_20002,N_10873,N_15007);
nor U20003 (N_20003,N_13799,N_12862);
or U20004 (N_20004,N_17517,N_17534);
and U20005 (N_20005,N_13015,N_16025);
xor U20006 (N_20006,N_12219,N_17109);
xor U20007 (N_20007,N_16780,N_15998);
xor U20008 (N_20008,N_16123,N_16702);
and U20009 (N_20009,N_16656,N_13155);
nor U20010 (N_20010,N_11312,N_12799);
nand U20011 (N_20011,N_10839,N_17758);
xor U20012 (N_20012,N_12641,N_18469);
nand U20013 (N_20013,N_13259,N_18909);
or U20014 (N_20014,N_13136,N_15666);
xor U20015 (N_20015,N_11976,N_12541);
xor U20016 (N_20016,N_19600,N_13875);
or U20017 (N_20017,N_13785,N_11079);
nand U20018 (N_20018,N_19464,N_12877);
nor U20019 (N_20019,N_17288,N_17639);
or U20020 (N_20020,N_16544,N_18533);
nand U20021 (N_20021,N_10180,N_15641);
and U20022 (N_20022,N_17623,N_16849);
or U20023 (N_20023,N_10610,N_10804);
and U20024 (N_20024,N_18174,N_19495);
xor U20025 (N_20025,N_19681,N_17078);
nor U20026 (N_20026,N_11755,N_11456);
nor U20027 (N_20027,N_10893,N_19684);
and U20028 (N_20028,N_10015,N_18952);
nand U20029 (N_20029,N_16081,N_10755);
or U20030 (N_20030,N_13534,N_16237);
and U20031 (N_20031,N_11325,N_13682);
xor U20032 (N_20032,N_19667,N_11113);
nor U20033 (N_20033,N_18302,N_11251);
nand U20034 (N_20034,N_13152,N_17310);
nand U20035 (N_20035,N_16838,N_16916);
or U20036 (N_20036,N_11141,N_15076);
or U20037 (N_20037,N_17342,N_15225);
and U20038 (N_20038,N_16685,N_11630);
and U20039 (N_20039,N_14393,N_13648);
or U20040 (N_20040,N_18216,N_15442);
and U20041 (N_20041,N_16418,N_11169);
nand U20042 (N_20042,N_11135,N_16731);
and U20043 (N_20043,N_15813,N_12720);
nor U20044 (N_20044,N_15157,N_10390);
xor U20045 (N_20045,N_13229,N_13522);
nand U20046 (N_20046,N_13450,N_15968);
nor U20047 (N_20047,N_14345,N_14563);
nor U20048 (N_20048,N_11443,N_16568);
xnor U20049 (N_20049,N_10957,N_15170);
or U20050 (N_20050,N_16890,N_18268);
nand U20051 (N_20051,N_11640,N_19620);
xor U20052 (N_20052,N_14484,N_11722);
or U20053 (N_20053,N_12557,N_13565);
nor U20054 (N_20054,N_13180,N_16172);
and U20055 (N_20055,N_18892,N_17742);
and U20056 (N_20056,N_18221,N_10356);
or U20057 (N_20057,N_11713,N_10846);
xnor U20058 (N_20058,N_17678,N_16255);
and U20059 (N_20059,N_13214,N_10993);
nand U20060 (N_20060,N_12568,N_17111);
nand U20061 (N_20061,N_10684,N_16018);
or U20062 (N_20062,N_11925,N_10441);
nor U20063 (N_20063,N_17622,N_10262);
nor U20064 (N_20064,N_17782,N_14387);
xnor U20065 (N_20065,N_16091,N_12684);
nand U20066 (N_20066,N_17512,N_18518);
nand U20067 (N_20067,N_15067,N_15193);
and U20068 (N_20068,N_15546,N_19624);
xor U20069 (N_20069,N_18482,N_13325);
xor U20070 (N_20070,N_10157,N_17492);
nand U20071 (N_20071,N_13745,N_10489);
xnor U20072 (N_20072,N_11863,N_12719);
and U20073 (N_20073,N_17659,N_13810);
and U20074 (N_20074,N_12352,N_18078);
nand U20075 (N_20075,N_10773,N_19007);
nor U20076 (N_20076,N_15000,N_16120);
nor U20077 (N_20077,N_18609,N_19457);
nor U20078 (N_20078,N_14213,N_11812);
or U20079 (N_20079,N_13000,N_18716);
nand U20080 (N_20080,N_15733,N_17168);
xor U20081 (N_20081,N_18391,N_17754);
or U20082 (N_20082,N_14756,N_10927);
nor U20083 (N_20083,N_14182,N_13542);
nor U20084 (N_20084,N_16115,N_12965);
or U20085 (N_20085,N_13725,N_14299);
or U20086 (N_20086,N_17529,N_16695);
nor U20087 (N_20087,N_19991,N_15343);
xor U20088 (N_20088,N_17525,N_12394);
and U20089 (N_20089,N_10621,N_14933);
and U20090 (N_20090,N_19721,N_17508);
nor U20091 (N_20091,N_12346,N_14144);
nor U20092 (N_20092,N_12001,N_18882);
nor U20093 (N_20093,N_10806,N_14335);
nand U20094 (N_20094,N_17478,N_13270);
and U20095 (N_20095,N_19739,N_11192);
xnor U20096 (N_20096,N_12879,N_12115);
nor U20097 (N_20097,N_14186,N_16814);
xnor U20098 (N_20098,N_16016,N_17069);
nor U20099 (N_20099,N_18126,N_16183);
nand U20100 (N_20100,N_11709,N_15751);
nor U20101 (N_20101,N_14128,N_10584);
and U20102 (N_20102,N_11446,N_16066);
nor U20103 (N_20103,N_12212,N_11508);
nor U20104 (N_20104,N_17079,N_19527);
nor U20105 (N_20105,N_17992,N_10860);
nand U20106 (N_20106,N_19585,N_18015);
xnor U20107 (N_20107,N_10506,N_10371);
and U20108 (N_20108,N_11944,N_10599);
xnor U20109 (N_20109,N_13528,N_19259);
nand U20110 (N_20110,N_15959,N_15856);
nor U20111 (N_20111,N_15415,N_12844);
xnor U20112 (N_20112,N_16156,N_11786);
nand U20113 (N_20113,N_13075,N_16096);
and U20114 (N_20114,N_16426,N_18683);
or U20115 (N_20115,N_19572,N_16068);
nand U20116 (N_20116,N_18874,N_19673);
or U20117 (N_20117,N_13198,N_13660);
or U20118 (N_20118,N_13492,N_16285);
xor U20119 (N_20119,N_19175,N_17337);
xnor U20120 (N_20120,N_17942,N_15297);
or U20121 (N_20121,N_12493,N_12163);
and U20122 (N_20122,N_14917,N_11857);
or U20123 (N_20123,N_19346,N_11780);
xor U20124 (N_20124,N_13949,N_12886);
nand U20125 (N_20125,N_13477,N_18331);
nand U20126 (N_20126,N_13192,N_14012);
nand U20127 (N_20127,N_19305,N_17896);
xor U20128 (N_20128,N_18919,N_10534);
nor U20129 (N_20129,N_13590,N_13472);
nor U20130 (N_20130,N_19955,N_19845);
and U20131 (N_20131,N_19756,N_14413);
nor U20132 (N_20132,N_14321,N_17422);
or U20133 (N_20133,N_17663,N_17156);
or U20134 (N_20134,N_19635,N_12967);
xnor U20135 (N_20135,N_11165,N_18059);
and U20136 (N_20136,N_15347,N_13438);
nand U20137 (N_20137,N_19246,N_18612);
xnor U20138 (N_20138,N_13020,N_12790);
nand U20139 (N_20139,N_12581,N_16798);
xnor U20140 (N_20140,N_18572,N_11178);
xnor U20141 (N_20141,N_14377,N_10131);
or U20142 (N_20142,N_16396,N_13564);
or U20143 (N_20143,N_17825,N_14284);
xor U20144 (N_20144,N_17693,N_19767);
nand U20145 (N_20145,N_19191,N_18012);
and U20146 (N_20146,N_11629,N_15576);
nand U20147 (N_20147,N_10124,N_12591);
nor U20148 (N_20148,N_19248,N_10077);
xnor U20149 (N_20149,N_14202,N_12389);
nor U20150 (N_20150,N_16268,N_18681);
and U20151 (N_20151,N_13604,N_10510);
xor U20152 (N_20152,N_15953,N_19717);
nand U20153 (N_20153,N_14098,N_16319);
or U20154 (N_20154,N_12547,N_10593);
xnor U20155 (N_20155,N_13372,N_17047);
nor U20156 (N_20156,N_11054,N_11573);
nand U20157 (N_20157,N_12985,N_16423);
or U20158 (N_20158,N_12653,N_13251);
and U20159 (N_20159,N_15381,N_17554);
nand U20160 (N_20160,N_15747,N_10564);
nor U20161 (N_20161,N_11952,N_16637);
and U20162 (N_20162,N_17088,N_12702);
nand U20163 (N_20163,N_16110,N_17443);
xnor U20164 (N_20164,N_19378,N_15251);
nand U20165 (N_20165,N_12495,N_18862);
or U20166 (N_20166,N_16470,N_11444);
nor U20167 (N_20167,N_18594,N_13841);
or U20168 (N_20168,N_13097,N_15571);
xor U20169 (N_20169,N_13333,N_14034);
xnor U20170 (N_20170,N_13529,N_18364);
or U20171 (N_20171,N_18337,N_12302);
nand U20172 (N_20172,N_18301,N_18604);
or U20173 (N_20173,N_13811,N_17154);
nand U20174 (N_20174,N_19576,N_16905);
xnor U20175 (N_20175,N_15500,N_16379);
or U20176 (N_20176,N_15321,N_13719);
nand U20177 (N_20177,N_14625,N_19461);
nor U20178 (N_20178,N_14600,N_16769);
or U20179 (N_20179,N_14216,N_17868);
xor U20180 (N_20180,N_15861,N_17461);
xor U20181 (N_20181,N_12096,N_19700);
nand U20182 (N_20182,N_18185,N_17619);
nor U20183 (N_20183,N_17062,N_14386);
or U20184 (N_20184,N_15783,N_13771);
or U20185 (N_20185,N_10772,N_18349);
xnor U20186 (N_20186,N_19167,N_13614);
nand U20187 (N_20187,N_16730,N_13615);
nand U20188 (N_20188,N_14181,N_10398);
nor U20189 (N_20189,N_13688,N_11663);
or U20190 (N_20190,N_15665,N_15431);
nor U20191 (N_20191,N_16304,N_15308);
nand U20192 (N_20192,N_12100,N_18929);
xor U20193 (N_20193,N_15525,N_19370);
and U20194 (N_20194,N_14928,N_11208);
or U20195 (N_20195,N_16220,N_15020);
and U20196 (N_20196,N_16185,N_12957);
xnor U20197 (N_20197,N_12535,N_15531);
or U20198 (N_20198,N_16491,N_12255);
or U20199 (N_20199,N_17832,N_16811);
or U20200 (N_20200,N_11384,N_19606);
and U20201 (N_20201,N_14565,N_15178);
nor U20202 (N_20202,N_18066,N_19902);
nand U20203 (N_20203,N_11343,N_16532);
nand U20204 (N_20204,N_10914,N_11739);
or U20205 (N_20205,N_12709,N_13824);
and U20206 (N_20206,N_11701,N_13717);
or U20207 (N_20207,N_19713,N_14220);
xor U20208 (N_20208,N_17008,N_16466);
nand U20209 (N_20209,N_18369,N_17700);
nor U20210 (N_20210,N_13007,N_13910);
or U20211 (N_20211,N_19610,N_16837);
nand U20212 (N_20212,N_12567,N_19813);
and U20213 (N_20213,N_19937,N_17287);
nor U20214 (N_20214,N_18426,N_13686);
xnor U20215 (N_20215,N_15978,N_13267);
nand U20216 (N_20216,N_17155,N_16474);
xor U20217 (N_20217,N_16817,N_12978);
xnor U20218 (N_20218,N_17974,N_12672);
xnor U20219 (N_20219,N_17230,N_16233);
and U20220 (N_20220,N_12640,N_14866);
or U20221 (N_20221,N_13040,N_13311);
nand U20222 (N_20222,N_10774,N_14308);
xor U20223 (N_20223,N_19117,N_12652);
xnor U20224 (N_20224,N_17209,N_18471);
or U20225 (N_20225,N_12201,N_16772);
and U20226 (N_20226,N_17875,N_17394);
nand U20227 (N_20227,N_19692,N_11134);
xor U20228 (N_20228,N_11289,N_13758);
or U20229 (N_20229,N_11085,N_14215);
nor U20230 (N_20230,N_18827,N_16948);
or U20231 (N_20231,N_11903,N_14588);
nand U20232 (N_20232,N_17851,N_17914);
xor U20233 (N_20233,N_17420,N_16103);
or U20234 (N_20234,N_18585,N_11557);
and U20235 (N_20235,N_15030,N_13399);
and U20236 (N_20236,N_12408,N_14319);
and U20237 (N_20237,N_16661,N_13840);
nor U20238 (N_20238,N_16313,N_11961);
or U20239 (N_20239,N_16572,N_10276);
nor U20240 (N_20240,N_13948,N_12998);
xnor U20241 (N_20241,N_11570,N_19106);
or U20242 (N_20242,N_11898,N_17296);
xnor U20243 (N_20243,N_12503,N_14719);
and U20244 (N_20244,N_11265,N_10147);
nand U20245 (N_20245,N_19404,N_15836);
and U20246 (N_20246,N_10940,N_11045);
nor U20247 (N_20247,N_13306,N_12164);
xnor U20248 (N_20248,N_16075,N_18635);
or U20249 (N_20249,N_12611,N_17481);
and U20250 (N_20250,N_17816,N_18641);
nand U20251 (N_20251,N_11324,N_11746);
or U20252 (N_20252,N_12135,N_16445);
nand U20253 (N_20253,N_11617,N_18982);
nor U20254 (N_20254,N_12062,N_18229);
xor U20255 (N_20255,N_12023,N_19124);
xnor U20256 (N_20256,N_14639,N_11571);
nor U20257 (N_20257,N_16259,N_14373);
nand U20258 (N_20258,N_19967,N_15638);
or U20259 (N_20259,N_11291,N_14615);
xor U20260 (N_20260,N_16834,N_16528);
xnor U20261 (N_20261,N_10938,N_11679);
xor U20262 (N_20262,N_11853,N_19649);
nand U20263 (N_20263,N_19321,N_18991);
or U20264 (N_20264,N_18043,N_12177);
nand U20265 (N_20265,N_11787,N_19381);
nor U20266 (N_20266,N_10508,N_13035);
and U20267 (N_20267,N_18409,N_18806);
or U20268 (N_20268,N_11523,N_14947);
and U20269 (N_20269,N_10532,N_18860);
or U20270 (N_20270,N_17737,N_12933);
nand U20271 (N_20271,N_18577,N_14322);
and U20272 (N_20272,N_18355,N_19060);
and U20273 (N_20273,N_13713,N_11299);
xor U20274 (N_20274,N_15167,N_18670);
nand U20275 (N_20275,N_17289,N_12361);
or U20276 (N_20276,N_13759,N_15675);
nor U20277 (N_20277,N_13307,N_15444);
xnor U20278 (N_20278,N_16196,N_19774);
nor U20279 (N_20279,N_16274,N_17925);
xnor U20280 (N_20280,N_18009,N_13865);
nand U20281 (N_20281,N_13550,N_19494);
nor U20282 (N_20282,N_12003,N_19376);
or U20283 (N_20283,N_15328,N_17530);
or U20284 (N_20284,N_18508,N_10876);
xnor U20285 (N_20285,N_10010,N_15952);
or U20286 (N_20286,N_12384,N_18879);
nand U20287 (N_20287,N_12937,N_19749);
nand U20288 (N_20288,N_19256,N_15687);
or U20289 (N_20289,N_11751,N_17785);
nand U20290 (N_20290,N_11146,N_18237);
and U20291 (N_20291,N_13796,N_10465);
and U20292 (N_20292,N_19625,N_19389);
or U20293 (N_20293,N_12808,N_13117);
or U20294 (N_20294,N_18274,N_13332);
nand U20295 (N_20295,N_19838,N_10429);
or U20296 (N_20296,N_11757,N_16188);
and U20297 (N_20297,N_15649,N_11792);
xor U20298 (N_20298,N_18852,N_12550);
or U20299 (N_20299,N_19819,N_10819);
nor U20300 (N_20300,N_15758,N_17355);
and U20301 (N_20301,N_11409,N_19946);
nand U20302 (N_20302,N_18651,N_11161);
and U20303 (N_20303,N_10812,N_14232);
nor U20304 (N_20304,N_11652,N_13278);
or U20305 (N_20305,N_18343,N_13519);
xnor U20306 (N_20306,N_17876,N_15117);
nor U20307 (N_20307,N_14158,N_13437);
xor U20308 (N_20308,N_18354,N_10394);
nor U20309 (N_20309,N_17564,N_14618);
nand U20310 (N_20310,N_17203,N_19997);
nand U20311 (N_20311,N_11465,N_12359);
and U20312 (N_20312,N_15651,N_18721);
nor U20313 (N_20313,N_18724,N_19951);
xor U20314 (N_20314,N_16339,N_12121);
nor U20315 (N_20315,N_12678,N_10255);
xor U20316 (N_20316,N_19851,N_11164);
or U20317 (N_20317,N_14962,N_10655);
nor U20318 (N_20318,N_19848,N_12109);
nand U20319 (N_20319,N_12191,N_15173);
nand U20320 (N_20320,N_16720,N_17953);
nor U20321 (N_20321,N_19471,N_18578);
and U20322 (N_20322,N_19932,N_11318);
xor U20323 (N_20323,N_10225,N_17674);
xor U20324 (N_20324,N_13303,N_12610);
xor U20325 (N_20325,N_19898,N_10918);
nor U20326 (N_20326,N_16264,N_15974);
xor U20327 (N_20327,N_17810,N_16836);
and U20328 (N_20328,N_15942,N_13718);
nor U20329 (N_20329,N_14260,N_10889);
nor U20330 (N_20330,N_10607,N_15116);
nor U20331 (N_20331,N_11087,N_10330);
nand U20332 (N_20332,N_16971,N_13668);
xnor U20333 (N_20333,N_15603,N_18096);
nor U20334 (N_20334,N_14069,N_16210);
xnor U20335 (N_20335,N_18989,N_12617);
or U20336 (N_20336,N_13181,N_19919);
xor U20337 (N_20337,N_18456,N_15830);
or U20338 (N_20338,N_19714,N_17715);
or U20339 (N_20339,N_10336,N_14318);
nor U20340 (N_20340,N_14786,N_16616);
nand U20341 (N_20341,N_16606,N_13247);
nand U20342 (N_20342,N_18685,N_16988);
nor U20343 (N_20343,N_12355,N_18050);
nor U20344 (N_20344,N_14400,N_14461);
xor U20345 (N_20345,N_19662,N_17378);
or U20346 (N_20346,N_14129,N_18633);
nand U20347 (N_20347,N_17753,N_11267);
and U20348 (N_20348,N_19509,N_19515);
nand U20349 (N_20349,N_12662,N_19458);
or U20350 (N_20350,N_15795,N_18452);
xor U20351 (N_20351,N_10998,N_14463);
nand U20352 (N_20352,N_10971,N_10058);
or U20353 (N_20353,N_16239,N_11985);
and U20354 (N_20354,N_18472,N_19672);
and U20355 (N_20355,N_12217,N_13200);
and U20356 (N_20356,N_14651,N_10982);
and U20357 (N_20357,N_16547,N_13358);
and U20358 (N_20358,N_12913,N_11461);
nor U20359 (N_20359,N_12485,N_18479);
nand U20360 (N_20360,N_19901,N_17035);
or U20361 (N_20361,N_18037,N_10039);
nand U20362 (N_20362,N_18584,N_13381);
and U20363 (N_20363,N_14860,N_18839);
and U20364 (N_20364,N_12880,N_14407);
or U20365 (N_20365,N_19785,N_18918);
and U20366 (N_20366,N_15997,N_11960);
or U20367 (N_20367,N_13780,N_14388);
or U20368 (N_20368,N_19675,N_18175);
nand U20369 (N_20369,N_18754,N_10220);
nor U20370 (N_20370,N_13254,N_14988);
and U20371 (N_20371,N_17829,N_18876);
and U20372 (N_20372,N_11368,N_12386);
nor U20373 (N_20373,N_15163,N_16759);
nand U20374 (N_20374,N_12296,N_16002);
or U20375 (N_20375,N_13849,N_13257);
or U20376 (N_20376,N_19472,N_18884);
nor U20377 (N_20377,N_19094,N_17057);
xnor U20378 (N_20378,N_12129,N_12940);
and U20379 (N_20379,N_14027,N_19922);
and U20380 (N_20380,N_11704,N_13154);
or U20381 (N_20381,N_18280,N_10376);
xnor U20382 (N_20382,N_12894,N_13894);
and U20383 (N_20383,N_17618,N_16394);
nand U20384 (N_20384,N_16820,N_16309);
or U20385 (N_20385,N_14164,N_19534);
nor U20386 (N_20386,N_14320,N_18778);
and U20387 (N_20387,N_10838,N_15661);
or U20388 (N_20388,N_12342,N_12939);
nand U20389 (N_20389,N_17637,N_14834);
xor U20390 (N_20390,N_14939,N_12156);
nand U20391 (N_20391,N_10603,N_16051);
nand U20392 (N_20392,N_16789,N_12083);
xnor U20393 (N_20393,N_18696,N_16258);
xor U20394 (N_20394,N_19799,N_17255);
or U20395 (N_20395,N_16131,N_10906);
xnor U20396 (N_20396,N_13500,N_10503);
nand U20397 (N_20397,N_12787,N_14520);
and U20398 (N_20398,N_13856,N_13217);
nor U20399 (N_20399,N_16711,N_16086);
and U20400 (N_20400,N_16871,N_10259);
nand U20401 (N_20401,N_18486,N_18614);
and U20402 (N_20402,N_16974,N_17240);
xnor U20403 (N_20403,N_14113,N_14776);
xor U20404 (N_20404,N_16013,N_10862);
nor U20405 (N_20405,N_16543,N_18453);
nor U20406 (N_20406,N_14586,N_14147);
xor U20407 (N_20407,N_11849,N_14751);
and U20408 (N_20408,N_10654,N_18883);
xnor U20409 (N_20409,N_18130,N_19917);
xnor U20410 (N_20410,N_10581,N_19956);
nand U20411 (N_20411,N_11483,N_16956);
xnor U20412 (N_20412,N_17595,N_14442);
or U20413 (N_20413,N_12968,N_14847);
nor U20414 (N_20414,N_15736,N_15038);
or U20415 (N_20415,N_18109,N_12513);
and U20416 (N_20416,N_17706,N_11627);
and U20417 (N_20417,N_12859,N_14088);
or U20418 (N_20418,N_10252,N_11071);
nand U20419 (N_20419,N_19658,N_14122);
nor U20420 (N_20420,N_13541,N_13232);
xor U20421 (N_20421,N_18141,N_18911);
xor U20422 (N_20422,N_11088,N_17976);
xor U20423 (N_20423,N_18138,N_14294);
nor U20424 (N_20424,N_16742,N_15074);
and U20425 (N_20425,N_16099,N_18468);
xnor U20426 (N_20426,N_18525,N_12802);
or U20427 (N_20427,N_13825,N_18782);
xor U20428 (N_20428,N_15555,N_11850);
nand U20429 (N_20429,N_17024,N_18484);
or U20430 (N_20430,N_16435,N_10929);
nor U20431 (N_20431,N_13631,N_10278);
nand U20432 (N_20432,N_10248,N_19407);
nor U20433 (N_20433,N_11973,N_11750);
xor U20434 (N_20434,N_11864,N_14076);
xor U20435 (N_20435,N_19545,N_19828);
or U20436 (N_20436,N_11065,N_11184);
nor U20437 (N_20437,N_15684,N_17537);
nand U20438 (N_20438,N_14398,N_19857);
or U20439 (N_20439,N_18671,N_13048);
nor U20440 (N_20440,N_16773,N_17684);
and U20441 (N_20441,N_15288,N_13034);
xnor U20442 (N_20442,N_12736,N_18285);
or U20443 (N_20443,N_15897,N_15222);
xnor U20444 (N_20444,N_18407,N_19390);
nor U20445 (N_20445,N_11730,N_13954);
or U20446 (N_20446,N_18213,N_10386);
or U20447 (N_20447,N_15887,N_10176);
or U20448 (N_20448,N_14217,N_19603);
xor U20449 (N_20449,N_19019,N_16372);
or U20450 (N_20450,N_19299,N_14993);
nor U20451 (N_20451,N_15370,N_13553);
xnor U20452 (N_20452,N_19514,N_13683);
or U20453 (N_20453,N_11800,N_16340);
nand U20454 (N_20454,N_13657,N_10751);
nand U20455 (N_20455,N_16852,N_10139);
nor U20456 (N_20456,N_12604,N_19221);
nor U20457 (N_20457,N_15791,N_16190);
xnor U20458 (N_20458,N_17189,N_12464);
and U20459 (N_20459,N_15544,N_14051);
nor U20460 (N_20460,N_10163,N_16082);
xnor U20461 (N_20461,N_10817,N_17726);
and U20462 (N_20462,N_16888,N_19100);
and U20463 (N_20463,N_12722,N_12596);
nand U20464 (N_20464,N_18664,N_14663);
or U20465 (N_20465,N_16935,N_18586);
and U20466 (N_20466,N_19274,N_17464);
xnor U20467 (N_20467,N_12800,N_19004);
nor U20468 (N_20468,N_19992,N_16316);
or U20469 (N_20469,N_14392,N_14270);
nor U20470 (N_20470,N_17695,N_12087);
and U20471 (N_20471,N_16984,N_16270);
nor U20472 (N_20472,N_18809,N_14914);
xnor U20473 (N_20473,N_18458,N_11945);
nand U20474 (N_20474,N_14857,N_17335);
and U20475 (N_20475,N_12784,N_19417);
and U20476 (N_20476,N_16132,N_19482);
or U20477 (N_20477,N_17015,N_14077);
and U20478 (N_20478,N_13546,N_14667);
xnor U20479 (N_20479,N_11260,N_12403);
nand U20480 (N_20480,N_14328,N_11575);
nor U20481 (N_20481,N_17356,N_16221);
and U20482 (N_20482,N_12282,N_14513);
nand U20483 (N_20483,N_11190,N_16252);
and U20484 (N_20484,N_12264,N_18908);
and U20485 (N_20485,N_13554,N_15459);
nand U20486 (N_20486,N_14883,N_12947);
and U20487 (N_20487,N_12078,N_14647);
nand U20488 (N_20488,N_18854,N_15709);
nand U20489 (N_20489,N_16095,N_10208);
nor U20490 (N_20490,N_13208,N_18904);
or U20491 (N_20491,N_14560,N_11379);
xnor U20492 (N_20492,N_13953,N_18785);
or U20493 (N_20493,N_12921,N_12585);
nand U20494 (N_20494,N_19978,N_11315);
or U20495 (N_20495,N_18548,N_12252);
nor U20496 (N_20496,N_14677,N_18972);
xnor U20497 (N_20497,N_16549,N_18397);
or U20498 (N_20498,N_14058,N_18385);
or U20499 (N_20499,N_17581,N_16301);
xnor U20500 (N_20500,N_19598,N_13363);
xor U20501 (N_20501,N_15581,N_16669);
nand U20502 (N_20502,N_12960,N_13858);
nor U20503 (N_20503,N_12836,N_17000);
xor U20504 (N_20504,N_19772,N_16964);
xnor U20505 (N_20505,N_10688,N_12487);
nand U20506 (N_20506,N_14790,N_17366);
nand U20507 (N_20507,N_19318,N_14376);
nor U20508 (N_20508,N_11900,N_11901);
nor U20509 (N_20509,N_10200,N_15694);
xor U20510 (N_20510,N_17719,N_18087);
nor U20511 (N_20511,N_12256,N_12423);
and U20512 (N_20512,N_19863,N_19449);
nand U20513 (N_20513,N_12673,N_18921);
nor U20514 (N_20514,N_10788,N_19434);
or U20515 (N_20515,N_19121,N_18928);
nand U20516 (N_20516,N_17865,N_18741);
and U20517 (N_20517,N_16144,N_16037);
or U20518 (N_20518,N_10114,N_12607);
or U20519 (N_20519,N_14124,N_17767);
or U20520 (N_20520,N_11340,N_13494);
and U20521 (N_20521,N_14330,N_10350);
or U20522 (N_20522,N_11290,N_14292);
nand U20523 (N_20523,N_18366,N_18736);
and U20524 (N_20524,N_13666,N_15467);
xnor U20525 (N_20525,N_15380,N_13999);
and U20526 (N_20526,N_15138,N_11525);
xnor U20527 (N_20527,N_10953,N_17463);
or U20528 (N_20528,N_15750,N_12152);
nand U20529 (N_20529,N_19493,N_19086);
and U20530 (N_20530,N_13701,N_17727);
nor U20531 (N_20531,N_17460,N_19268);
and U20532 (N_20532,N_14490,N_18687);
and U20533 (N_20533,N_19786,N_15787);
and U20534 (N_20534,N_17169,N_11577);
xor U20535 (N_20535,N_12949,N_13893);
nor U20536 (N_20536,N_12024,N_10351);
xor U20537 (N_20537,N_19832,N_16804);
nor U20538 (N_20538,N_16214,N_19688);
xor U20539 (N_20539,N_13587,N_11455);
nand U20540 (N_20540,N_18746,N_19050);
and U20541 (N_20541,N_19241,N_16589);
nand U20542 (N_20542,N_17406,N_10340);
nand U20543 (N_20543,N_17361,N_15833);
or U20544 (N_20544,N_11632,N_15913);
xor U20545 (N_20545,N_10909,N_13371);
nor U20546 (N_20546,N_15517,N_10308);
nand U20547 (N_20547,N_16179,N_17036);
nor U20548 (N_20548,N_14643,N_18916);
nand U20549 (N_20549,N_12624,N_14753);
or U20550 (N_20550,N_18187,N_17430);
nand U20551 (N_20551,N_10695,N_13431);
nor U20552 (N_20552,N_14635,N_12339);
nor U20553 (N_20553,N_17037,N_18532);
xnor U20554 (N_20554,N_16879,N_18230);
nor U20555 (N_20555,N_10515,N_13389);
nor U20556 (N_20556,N_16858,N_14946);
or U20557 (N_20557,N_11127,N_10861);
or U20558 (N_20558,N_19961,N_18017);
nand U20559 (N_20559,N_11582,N_18372);
or U20560 (N_20560,N_19797,N_16565);
nand U20561 (N_20561,N_12349,N_14465);
nor U20562 (N_20562,N_13377,N_16665);
and U20563 (N_20563,N_14264,N_10310);
or U20564 (N_20564,N_17772,N_19454);
and U20565 (N_20565,N_17970,N_16999);
nand U20566 (N_20566,N_13105,N_10930);
nand U20567 (N_20567,N_17377,N_15976);
or U20568 (N_20568,N_18753,N_15411);
nor U20569 (N_20569,N_15994,N_14218);
nand U20570 (N_20570,N_17065,N_13226);
xnor U20571 (N_20571,N_15731,N_14084);
xor U20572 (N_20572,N_19187,N_17012);
and U20573 (N_20573,N_14976,N_14549);
nor U20574 (N_20574,N_11781,N_12701);
nand U20575 (N_20575,N_11152,N_12814);
nand U20576 (N_20576,N_15725,N_17649);
or U20577 (N_20577,N_10721,N_11584);
nor U20578 (N_20578,N_16581,N_15105);
nand U20579 (N_20579,N_19513,N_15711);
nor U20580 (N_20580,N_15695,N_15653);
nand U20581 (N_20581,N_16518,N_18142);
and U20582 (N_20582,N_16440,N_11707);
xnor U20583 (N_20583,N_14943,N_19815);
or U20584 (N_20584,N_15153,N_18703);
or U20585 (N_20585,N_11258,N_16447);
xor U20586 (N_20586,N_13364,N_15377);
or U20587 (N_20587,N_15062,N_18234);
or U20588 (N_20588,N_13687,N_13121);
xnor U20589 (N_20589,N_18235,N_17667);
xnor U20590 (N_20590,N_16217,N_19846);
and U20591 (N_20591,N_11837,N_19265);
or U20592 (N_20592,N_18106,N_13184);
and U20593 (N_20593,N_11489,N_11090);
nor U20594 (N_20594,N_17094,N_17756);
nor U20595 (N_20595,N_18330,N_11026);
xnor U20596 (N_20596,N_13765,N_12283);
nand U20597 (N_20597,N_11606,N_14668);
nand U20598 (N_20598,N_18328,N_17298);
xor U20599 (N_20599,N_10573,N_18654);
xnor U20600 (N_20600,N_14234,N_18069);
and U20601 (N_20601,N_15093,N_19689);
and U20602 (N_20602,N_13862,N_18675);
nand U20603 (N_20603,N_12057,N_14496);
or U20604 (N_20604,N_10140,N_17257);
nor U20605 (N_20605,N_14835,N_10912);
nor U20606 (N_20606,N_15604,N_17668);
and U20607 (N_20607,N_15068,N_19000);
nor U20608 (N_20608,N_16453,N_12856);
nor U20609 (N_20609,N_14474,N_14431);
and U20610 (N_20610,N_10438,N_12443);
xnor U20611 (N_20611,N_14825,N_19157);
or U20612 (N_20612,N_10545,N_14604);
and U20613 (N_20613,N_14481,N_16228);
nor U20614 (N_20614,N_13463,N_14033);
and U20615 (N_20615,N_18920,N_16882);
or U20616 (N_20616,N_14223,N_16015);
nor U20617 (N_20617,N_13400,N_12973);
nor U20618 (N_20618,N_10104,N_18261);
nand U20619 (N_20619,N_18521,N_12488);
nor U20620 (N_20620,N_17138,N_13816);
and U20621 (N_20621,N_13053,N_12074);
nor U20622 (N_20622,N_14009,N_18367);
nand U20623 (N_20623,N_14907,N_16560);
nand U20624 (N_20624,N_11041,N_17265);
nand U20625 (N_20625,N_18254,N_11555);
xnor U20626 (N_20626,N_15757,N_13467);
and U20627 (N_20627,N_13293,N_15362);
and U20628 (N_20628,N_14466,N_18303);
and U20629 (N_20629,N_13628,N_17453);
nand U20630 (N_20630,N_18528,N_11330);
or U20631 (N_20631,N_11078,N_19706);
or U20632 (N_20632,N_14080,N_17780);
nand U20633 (N_20633,N_11230,N_14529);
xnor U20634 (N_20634,N_10379,N_10955);
xnor U20635 (N_20635,N_18042,N_16357);
and U20636 (N_20636,N_10537,N_11328);
or U20637 (N_20637,N_15676,N_16812);
or U20638 (N_20638,N_14878,N_13063);
and U20639 (N_20639,N_15645,N_15671);
nand U20640 (N_20640,N_13694,N_16178);
and U20641 (N_20641,N_13056,N_18131);
or U20642 (N_20642,N_14152,N_13113);
or U20643 (N_20643,N_19076,N_10093);
or U20644 (N_20644,N_14055,N_16652);
nor U20645 (N_20645,N_17899,N_18810);
nand U20646 (N_20646,N_11259,N_18733);
or U20647 (N_20647,N_17547,N_15748);
and U20648 (N_20648,N_16280,N_13932);
nor U20649 (N_20649,N_17916,N_10285);
or U20650 (N_20650,N_19468,N_17446);
xor U20651 (N_20651,N_10574,N_15706);
and U20652 (N_20652,N_15151,N_10224);
xor U20653 (N_20653,N_13933,N_15699);
nor U20654 (N_20654,N_16562,N_18722);
or U20655 (N_20655,N_12499,N_10052);
xor U20656 (N_20656,N_12143,N_13070);
nand U20657 (N_20657,N_17596,N_11556);
or U20658 (N_20658,N_15989,N_15796);
or U20659 (N_20659,N_16147,N_10756);
and U20660 (N_20660,N_15189,N_13741);
nor U20661 (N_20661,N_10109,N_18710);
and U20662 (N_20662,N_19609,N_13350);
xnor U20663 (N_20663,N_18922,N_13961);
xnor U20664 (N_20664,N_17820,N_17256);
xnor U20665 (N_20665,N_10703,N_19567);
xnor U20666 (N_20666,N_11975,N_14743);
nand U20667 (N_20667,N_18262,N_12376);
xor U20668 (N_20668,N_16061,N_12025);
xor U20669 (N_20669,N_19808,N_19727);
or U20670 (N_20670,N_12006,N_18208);
and U20671 (N_20671,N_14272,N_15497);
nor U20672 (N_20672,N_17385,N_13183);
or U20673 (N_20673,N_19111,N_12297);
nor U20674 (N_20674,N_11426,N_12295);
nor U20675 (N_20675,N_18896,N_15739);
nor U20676 (N_20676,N_14775,N_12054);
or U20677 (N_20677,N_11899,N_14121);
or U20678 (N_20678,N_17149,N_14780);
or U20679 (N_20679,N_17631,N_16557);
xnor U20680 (N_20680,N_16083,N_18542);
xnor U20681 (N_20681,N_11689,N_19487);
xor U20682 (N_20682,N_15246,N_16593);
nand U20683 (N_20683,N_11044,N_11093);
nand U20684 (N_20684,N_19842,N_19962);
nor U20685 (N_20685,N_17329,N_15501);
nand U20686 (N_20686,N_10651,N_16939);
xor U20687 (N_20687,N_14265,N_19555);
xnor U20688 (N_20688,N_19806,N_18063);
and U20689 (N_20689,N_11687,N_12857);
and U20690 (N_20690,N_13890,N_12766);
xor U20691 (N_20691,N_19271,N_17073);
or U20692 (N_20692,N_10118,N_13148);
and U20693 (N_20693,N_19260,N_13561);
nor U20694 (N_20694,N_16204,N_12315);
or U20695 (N_20695,N_16602,N_11529);
nor U20696 (N_20696,N_11370,N_12867);
or U20697 (N_20697,N_19016,N_18764);
or U20698 (N_20698,N_10578,N_16722);
nor U20699 (N_20699,N_17511,N_17175);
and U20700 (N_20700,N_17243,N_17885);
nand U20701 (N_20701,N_15802,N_15097);
or U20702 (N_20702,N_13588,N_11672);
xnor U20703 (N_20703,N_12579,N_13611);
nor U20704 (N_20704,N_15550,N_14471);
and U20705 (N_20705,N_12052,N_18197);
or U20706 (N_20706,N_12105,N_15294);
or U20707 (N_20707,N_12042,N_14531);
nor U20708 (N_20708,N_13511,N_11929);
and U20709 (N_20709,N_16413,N_12823);
and U20710 (N_20710,N_15600,N_16021);
and U20711 (N_20711,N_13654,N_18190);
or U20712 (N_20712,N_16114,N_14488);
nand U20713 (N_20713,N_18600,N_19745);
nand U20714 (N_20714,N_19730,N_14521);
xor U20715 (N_20715,N_11189,N_17043);
nand U20716 (N_20716,N_13794,N_12243);
and U20717 (N_20717,N_12885,N_15658);
nor U20718 (N_20718,N_13599,N_16643);
nand U20719 (N_20719,N_18449,N_14443);
xnor U20720 (N_20720,N_18728,N_19194);
nor U20721 (N_20721,N_15866,N_10222);
nor U20722 (N_20722,N_13379,N_19385);
nand U20723 (N_20723,N_13557,N_10900);
and U20724 (N_20724,N_17895,N_14979);
and U20725 (N_20725,N_12077,N_11433);
and U20726 (N_20726,N_18501,N_19112);
nor U20727 (N_20727,N_10094,N_19161);
nor U20728 (N_20728,N_19904,N_17862);
xnor U20729 (N_20729,N_17826,N_15708);
or U20730 (N_20730,N_16963,N_10363);
nor U20731 (N_20731,N_13280,N_10837);
or U20732 (N_20732,N_13475,N_17325);
xnor U20733 (N_20733,N_11292,N_15395);
and U20734 (N_20734,N_18519,N_16787);
and U20735 (N_20735,N_19452,N_16671);
xnor U20736 (N_20736,N_16551,N_15504);
or U20737 (N_20737,N_19431,N_15019);
or U20738 (N_20738,N_15724,N_11940);
and U20739 (N_20739,N_11472,N_19960);
or U20740 (N_20740,N_13126,N_13812);
or U20741 (N_20741,N_17379,N_17658);
nand U20742 (N_20742,N_15557,N_18094);
and U20743 (N_20743,N_14394,N_16523);
nand U20744 (N_20744,N_17709,N_17686);
xor U20745 (N_20745,N_19477,N_11873);
xor U20746 (N_20746,N_13174,N_13527);
or U20747 (N_20747,N_11377,N_17309);
nor U20748 (N_20748,N_10550,N_16932);
nand U20749 (N_20749,N_19219,N_18300);
or U20750 (N_20750,N_11421,N_14766);
and U20751 (N_20751,N_13285,N_14797);
or U20752 (N_20752,N_13055,N_17603);
and U20753 (N_20753,N_17994,N_19450);
or U20754 (N_20754,N_13861,N_17219);
nor U20755 (N_20755,N_12491,N_15874);
nand U20756 (N_20756,N_16628,N_18321);
and U20757 (N_20757,N_13574,N_12711);
nand U20758 (N_20758,N_18742,N_15420);
or U20759 (N_20759,N_16124,N_15090);
nand U20760 (N_20760,N_19342,N_13420);
or U20761 (N_20761,N_10085,N_12817);
or U20762 (N_20762,N_10009,N_18476);
nor U20763 (N_20763,N_11840,N_10711);
nor U20764 (N_20764,N_16979,N_11760);
xnor U20765 (N_20765,N_10969,N_10619);
nor U20766 (N_20766,N_19938,N_19605);
xnor U20767 (N_20767,N_17045,N_17085);
xnor U20768 (N_20768,N_12614,N_15851);
nand U20769 (N_20769,N_10349,N_19329);
and U20770 (N_20770,N_19532,N_17142);
or U20771 (N_20771,N_19811,N_14469);
nand U20772 (N_20772,N_10805,N_14703);
or U20773 (N_20773,N_12745,N_15607);
nand U20774 (N_20774,N_18562,N_17343);
nand U20775 (N_20775,N_17053,N_11788);
xor U20776 (N_20776,N_16128,N_17427);
and U20777 (N_20777,N_14354,N_12108);
nand U20778 (N_20778,N_11852,N_19678);
xor U20779 (N_20779,N_13792,N_14408);
nor U20780 (N_20780,N_19027,N_18709);
and U20781 (N_20781,N_16201,N_14117);
or U20782 (N_20782,N_14470,N_16738);
or U20783 (N_20783,N_19465,N_18099);
nand U20784 (N_20784,N_13915,N_13296);
and U20785 (N_20785,N_13501,N_10195);
nand U20786 (N_20786,N_14519,N_18248);
nor U20787 (N_20787,N_18073,N_13715);
xor U20788 (N_20788,N_14083,N_13595);
or U20789 (N_20789,N_11737,N_14656);
nand U20790 (N_20790,N_11890,N_16077);
nand U20791 (N_20791,N_11649,N_15311);
nand U20792 (N_20792,N_13854,N_13456);
xnor U20793 (N_20793,N_19456,N_19039);
or U20794 (N_20794,N_11070,N_14018);
nor U20795 (N_20795,N_11022,N_18666);
and U20796 (N_20796,N_10364,N_12696);
and U20797 (N_20797,N_11938,N_10003);
or U20798 (N_20798,N_18446,N_11868);
xor U20799 (N_20799,N_12822,N_18289);
and U20800 (N_20800,N_18531,N_15502);
xnor U20801 (N_20801,N_10101,N_12277);
nand U20802 (N_20802,N_16863,N_15633);
nand U20803 (N_20803,N_16150,N_19950);
or U20804 (N_20804,N_10137,N_12562);
and U20805 (N_20805,N_19959,N_10347);
nor U20806 (N_20806,N_19198,N_12110);
xor U20807 (N_20807,N_12291,N_17951);
and U20808 (N_20808,N_15002,N_19551);
xnor U20809 (N_20809,N_14696,N_12863);
nand U20810 (N_20810,N_15084,N_15013);
nand U20811 (N_20811,N_14814,N_14017);
nand U20812 (N_20812,N_10030,N_12132);
and U20813 (N_20813,N_19866,N_14103);
or U20814 (N_20814,N_15200,N_16111);
xnor U20815 (N_20815,N_13696,N_12433);
nand U20816 (N_20816,N_17192,N_17212);
nand U20817 (N_20817,N_15896,N_16914);
xor U20818 (N_20818,N_17692,N_11793);
xnor U20819 (N_20819,N_19234,N_16501);
nand U20820 (N_20820,N_15564,N_15061);
or U20821 (N_20821,N_19170,N_16674);
and U20822 (N_20822,N_12457,N_19484);
and U20823 (N_20823,N_18359,N_18569);
and U20824 (N_20824,N_16736,N_11979);
or U20825 (N_20825,N_10372,N_16521);
nand U20826 (N_20826,N_16520,N_10521);
or U20827 (N_20827,N_10402,N_10728);
or U20828 (N_20828,N_14090,N_19723);
xor U20829 (N_20829,N_19447,N_17578);
nor U20830 (N_20830,N_16017,N_15313);
or U20831 (N_20831,N_10939,N_18105);
and U20832 (N_20832,N_16815,N_12040);
or U20833 (N_20833,N_12775,N_13790);
or U20834 (N_20834,N_18793,N_18377);
nand U20835 (N_20835,N_18250,N_16928);
nor U20836 (N_20836,N_10082,N_15578);
nor U20837 (N_20837,N_13109,N_13436);
nor U20838 (N_20838,N_18825,N_14682);
or U20839 (N_20839,N_12236,N_13223);
nor U20840 (N_20840,N_12914,N_10617);
and U20841 (N_20841,N_13434,N_18252);
xnor U20842 (N_20842,N_17839,N_13926);
nand U20843 (N_20843,N_12837,N_18020);
or U20844 (N_20844,N_16945,N_10182);
xor U20845 (N_20845,N_18751,N_13986);
and U20846 (N_20846,N_17389,N_18749);
nand U20847 (N_20847,N_13442,N_10870);
nor U20848 (N_20848,N_19831,N_15280);
xor U20849 (N_20849,N_19653,N_19397);
and U20850 (N_20850,N_15229,N_12801);
xnor U20851 (N_20851,N_11228,N_11311);
or U20852 (N_20852,N_17740,N_15925);
nor U20853 (N_20853,N_10132,N_15456);
nand U20854 (N_20854,N_12750,N_16566);
nor U20855 (N_20855,N_19693,N_15884);
and U20856 (N_20856,N_19650,N_14068);
xor U20857 (N_20857,N_16390,N_12715);
or U20858 (N_20858,N_19270,N_11670);
or U20859 (N_20859,N_18832,N_18512);
nor U20860 (N_20860,N_19971,N_16385);
xnor U20861 (N_20861,N_16384,N_14889);
xnor U20862 (N_20862,N_12203,N_17952);
nand U20863 (N_20863,N_15883,N_17735);
nand U20864 (N_20864,N_17769,N_17315);
nor U20865 (N_20865,N_10242,N_10303);
nand U20866 (N_20866,N_14168,N_17878);
or U20867 (N_20867,N_19120,N_10383);
or U20868 (N_20868,N_11566,N_15838);
or U20869 (N_20869,N_16824,N_13453);
or U20870 (N_20870,N_11802,N_11109);
or U20871 (N_20871,N_11631,N_17893);
or U20872 (N_20872,N_15639,N_18869);
nand U20873 (N_20873,N_15806,N_17158);
nor U20874 (N_20874,N_11838,N_10282);
and U20875 (N_20875,N_15800,N_16653);
nor U20876 (N_20876,N_14823,N_18658);
nand U20877 (N_20877,N_12168,N_11522);
and U20878 (N_20878,N_14153,N_15114);
or U20879 (N_20879,N_13081,N_17400);
and U20880 (N_20880,N_19057,N_12575);
and U20881 (N_20881,N_11677,N_13324);
nor U20882 (N_20882,N_17147,N_15785);
or U20883 (N_20883,N_18979,N_10338);
nand U20884 (N_20884,N_16299,N_19258);
and U20885 (N_20885,N_18924,N_14454);
or U20886 (N_20886,N_18259,N_19871);
or U20887 (N_20887,N_12971,N_12180);
nor U20888 (N_20888,N_17063,N_13271);
xor U20889 (N_20889,N_15334,N_16020);
and U20890 (N_20890,N_19580,N_12334);
nand U20891 (N_20891,N_17569,N_13766);
nand U20892 (N_20892,N_11487,N_13883);
xor U20893 (N_20893,N_15967,N_19463);
xnor U20894 (N_20894,N_14874,N_17474);
or U20895 (N_20895,N_18006,N_18556);
nor U20896 (N_20896,N_14198,N_11692);
or U20897 (N_20897,N_13253,N_14449);
xnor U20898 (N_20898,N_12118,N_12543);
nand U20899 (N_20899,N_12520,N_10525);
nand U20900 (N_20900,N_15601,N_18786);
or U20901 (N_20901,N_10606,N_12450);
nor U20902 (N_20902,N_19704,N_18726);
and U20903 (N_20903,N_10726,N_11829);
nor U20904 (N_20904,N_13268,N_17591);
nand U20905 (N_20905,N_15848,N_13680);
xnor U20906 (N_20906,N_16625,N_19097);
nand U20907 (N_20907,N_10044,N_11182);
nand U20908 (N_20908,N_14028,N_12634);
xnor U20909 (N_20909,N_14902,N_12944);
nor U20910 (N_20910,N_18159,N_17943);
nor U20911 (N_20911,N_19896,N_10706);
nand U20912 (N_20912,N_18291,N_15469);
xor U20913 (N_20913,N_19566,N_16163);
and U20914 (N_20914,N_12991,N_18700);
nor U20915 (N_20915,N_12743,N_10397);
nand U20916 (N_20916,N_12514,N_13098);
nand U20917 (N_20917,N_15130,N_11462);
xnor U20918 (N_20918,N_18402,N_14106);
xor U20919 (N_20919,N_15915,N_15050);
nor U20920 (N_20920,N_13985,N_12628);
xor U20921 (N_20921,N_12651,N_14371);
nand U20922 (N_20922,N_18606,N_15143);
and U20923 (N_20923,N_15702,N_18002);
and U20924 (N_20924,N_17297,N_13735);
xor U20925 (N_20925,N_17485,N_10190);
or U20926 (N_20926,N_11641,N_18619);
xnor U20927 (N_20927,N_16057,N_16472);
xnor U20928 (N_20928,N_16718,N_11481);
nor U20929 (N_20929,N_15843,N_12563);
xor U20930 (N_20930,N_12521,N_16659);
nand U20931 (N_20931,N_15947,N_15327);
xor U20932 (N_20932,N_12727,N_11610);
nor U20933 (N_20933,N_11493,N_11814);
xor U20934 (N_20934,N_11005,N_12552);
nor U20935 (N_20935,N_13620,N_13598);
or U20936 (N_20936,N_12470,N_15141);
nand U20937 (N_20937,N_13722,N_19497);
or U20938 (N_20938,N_12287,N_19856);
xor U20939 (N_20939,N_12644,N_19733);
xor U20940 (N_20940,N_17223,N_13791);
nand U20941 (N_20941,N_15971,N_12395);
xnor U20942 (N_20942,N_16553,N_18384);
or U20943 (N_20943,N_15098,N_16310);
or U20944 (N_20944,N_18317,N_11568);
nand U20945 (N_20945,N_12390,N_14538);
nor U20946 (N_20946,N_16667,N_10586);
nor U20947 (N_20947,N_10964,N_14527);
or U20948 (N_20948,N_16266,N_14486);
or U20949 (N_20949,N_11219,N_11789);
nand U20950 (N_20950,N_16182,N_11154);
or U20951 (N_20951,N_15816,N_19781);
and U20952 (N_20952,N_10797,N_13967);
nor U20953 (N_20953,N_13721,N_13752);
and U20954 (N_20954,N_11778,N_10113);
nand U20955 (N_20955,N_17761,N_18643);
nand U20956 (N_20956,N_11333,N_18655);
nand U20957 (N_20957,N_12911,N_17750);
and U20958 (N_20958,N_11338,N_17208);
nand U20959 (N_20959,N_10999,N_11372);
nand U20960 (N_20960,N_10116,N_11972);
nand U20961 (N_20961,N_16107,N_11067);
nand U20962 (N_20962,N_15439,N_12032);
and U20963 (N_20963,N_13651,N_13288);
nand U20964 (N_20964,N_18206,N_17590);
xnor U20965 (N_20965,N_14050,N_14462);
and U20966 (N_20966,N_14110,N_14433);
nor U20967 (N_20967,N_12178,N_17732);
or U20968 (N_20968,N_18808,N_13592);
nand U20969 (N_20969,N_14777,N_12028);
or U20970 (N_20970,N_19127,N_17921);
and U20971 (N_20971,N_10801,N_10354);
and U20972 (N_20972,N_11224,N_17654);
nand U20973 (N_20973,N_14922,N_10766);
nand U20974 (N_20974,N_15282,N_13928);
nor U20975 (N_20975,N_11799,N_13107);
and U20976 (N_20976,N_13709,N_12215);
xor U20977 (N_20977,N_14816,N_12262);
and U20978 (N_20978,N_17447,N_14989);
nor U20979 (N_20979,N_14035,N_19143);
xor U20980 (N_20980,N_17206,N_17960);
or U20981 (N_20981,N_14846,N_16230);
or U20982 (N_20982,N_19707,N_12343);
or U20983 (N_20983,N_17589,N_15175);
nor U20984 (N_20984,N_12528,N_11309);
nor U20985 (N_20985,N_19795,N_11831);
and U20986 (N_20986,N_11614,N_13909);
and U20987 (N_20987,N_18824,N_11346);
xnor U20988 (N_20988,N_12927,N_15774);
xnor U20989 (N_20989,N_13300,N_10328);
nand U20990 (N_20990,N_17253,N_12088);
or U20991 (N_20991,N_13900,N_14064);
nor U20992 (N_20992,N_13488,N_10119);
and U20993 (N_20993,N_14426,N_11550);
nand U20994 (N_20994,N_14590,N_11836);
and U20995 (N_20995,N_15202,N_16832);
nor U20996 (N_20996,N_10373,N_12222);
and U20997 (N_20997,N_17001,N_17666);
and U20998 (N_20998,N_15124,N_17891);
and U20999 (N_20999,N_10989,N_17075);
nand U21000 (N_21000,N_17842,N_14997);
or U21001 (N_21001,N_11254,N_15199);
xnor U21002 (N_21002,N_18413,N_14545);
nand U21003 (N_21003,N_10341,N_16165);
or U21004 (N_21004,N_18582,N_17655);
nand U21005 (N_21005,N_18495,N_17180);
nand U21006 (N_21006,N_19333,N_17981);
xor U21007 (N_21007,N_18956,N_15622);
and U21008 (N_21008,N_17457,N_15372);
or U21009 (N_21009,N_13760,N_12337);
nand U21010 (N_21010,N_14238,N_13165);
nor U21011 (N_21011,N_11782,N_15149);
nor U21012 (N_21012,N_16823,N_13864);
xnor U21013 (N_21013,N_13134,N_12293);
nand U21014 (N_21014,N_10990,N_17587);
or U21015 (N_21015,N_19581,N_14812);
nor U21016 (N_21016,N_12330,N_17087);
nand U21017 (N_21017,N_10829,N_12454);
nand U21018 (N_21018,N_11454,N_19179);
xnor U21019 (N_21019,N_18125,N_10261);
nor U21020 (N_21020,N_14646,N_15409);
or U21021 (N_21021,N_13860,N_18680);
nand U21022 (N_21022,N_14702,N_15119);
or U21023 (N_21023,N_19595,N_14092);
nand U21024 (N_21024,N_19539,N_19384);
nand U21025 (N_21025,N_10378,N_10423);
xnor U21026 (N_21026,N_19929,N_15669);
or U21027 (N_21027,N_11683,N_19419);
xnor U21028 (N_21028,N_12600,N_18613);
or U21029 (N_21029,N_18238,N_13918);
and U21030 (N_21030,N_12734,N_18357);
nand U21031 (N_21031,N_11142,N_18318);
nand U21032 (N_21032,N_15535,N_18155);
nor U21033 (N_21033,N_19829,N_15433);
xnor U21034 (N_21034,N_19753,N_14107);
xnor U21035 (N_21035,N_17330,N_15964);
nor U21036 (N_21036,N_10549,N_19920);
nor U21037 (N_21037,N_11907,N_17369);
and U21038 (N_21038,N_13584,N_13163);
or U21039 (N_21039,N_19348,N_13408);
and U21040 (N_21040,N_14209,N_17060);
nor U21041 (N_21041,N_16484,N_14119);
or U21042 (N_21042,N_18387,N_12809);
or U21043 (N_21043,N_12265,N_10274);
and U21044 (N_21044,N_14898,N_12982);
or U21045 (N_21045,N_15759,N_18797);
nand U21046 (N_21046,N_14525,N_12713);
and U21047 (N_21047,N_12932,N_14798);
and U21048 (N_21048,N_19490,N_19957);
and U21049 (N_21049,N_12375,N_19180);
or U21050 (N_21050,N_16098,N_13207);
and U21051 (N_21051,N_14840,N_11204);
nor U21052 (N_21052,N_15465,N_12496);
or U21053 (N_21053,N_15730,N_19425);
and U21054 (N_21054,N_18552,N_15357);
nor U21055 (N_21055,N_12595,N_15919);
or U21056 (N_21056,N_13065,N_19945);
nor U21057 (N_21057,N_17290,N_15212);
or U21058 (N_21058,N_17239,N_10904);
nor U21059 (N_21059,N_15021,N_14712);
nor U21060 (N_21060,N_19291,N_10732);
xor U21061 (N_21061,N_13882,N_11374);
xor U21062 (N_21062,N_12492,N_14448);
and U21063 (N_21063,N_18507,N_18296);
and U21064 (N_21064,N_11809,N_15491);
xor U21065 (N_21065,N_17908,N_13945);
or U21066 (N_21066,N_10466,N_11255);
nor U21067 (N_21067,N_11441,N_10512);
xnor U21068 (N_21068,N_16349,N_12587);
nand U21069 (N_21069,N_19220,N_16439);
nor U21070 (N_21070,N_14888,N_13401);
and U21071 (N_21071,N_13979,N_10495);
and U21072 (N_21072,N_19686,N_15176);
and U21073 (N_21073,N_14197,N_11813);
and U21074 (N_21074,N_19056,N_11741);
xor U21075 (N_21075,N_11125,N_18958);
nand U21076 (N_21076,N_14190,N_10555);
nor U21077 (N_21077,N_12017,N_17806);
xor U21078 (N_21078,N_16424,N_13199);
nand U21079 (N_21079,N_18396,N_12570);
xnor U21080 (N_21080,N_17751,N_16597);
nor U21081 (N_21081,N_13244,N_15426);
and U21082 (N_21082,N_16276,N_11098);
and U21083 (N_21083,N_15755,N_11080);
nand U21084 (N_21084,N_12340,N_16240);
nand U21085 (N_21085,N_14315,N_12553);
nand U21086 (N_21086,N_15317,N_17033);
nand U21087 (N_21087,N_15900,N_13495);
nor U21088 (N_21088,N_10670,N_11223);
or U21089 (N_21089,N_11160,N_13060);
and U21090 (N_21090,N_15008,N_18489);
nand U21091 (N_21091,N_17638,N_17927);
nand U21092 (N_21092,N_16208,N_12693);
nand U21093 (N_21093,N_17070,N_12064);
nand U21094 (N_21094,N_15272,N_19072);
and U21095 (N_21095,N_18417,N_11790);
xnor U21096 (N_21096,N_12011,N_11362);
nand U21097 (N_21097,N_14805,N_10145);
nor U21098 (N_21098,N_15955,N_12586);
nor U21099 (N_21099,N_11430,N_14199);
nand U21100 (N_21100,N_14801,N_18004);
xnor U21101 (N_21101,N_19469,N_11645);
and U21102 (N_21102,N_14528,N_12504);
and U21103 (N_21103,N_17375,N_17258);
and U21104 (N_21104,N_18711,N_14355);
nor U21105 (N_21105,N_15112,N_15752);
xnor U21106 (N_21106,N_17945,N_16854);
and U21107 (N_21107,N_18022,N_19430);
nor U21108 (N_21108,N_12429,N_13545);
nand U21109 (N_21109,N_12771,N_15850);
and U21110 (N_21110,N_19351,N_10269);
nor U21111 (N_21111,N_13242,N_10004);
nand U21112 (N_21112,N_13366,N_10243);
nand U21113 (N_21113,N_13009,N_10088);
xnor U21114 (N_21114,N_11053,N_14932);
or U21115 (N_21115,N_12288,N_15972);
or U21116 (N_21116,N_16273,N_18857);
and U21117 (N_21117,N_14870,N_18947);
and U21118 (N_21118,N_10295,N_18147);
xor U21119 (N_21119,N_14277,N_19188);
nand U21120 (N_21120,N_10068,N_12812);
xor U21121 (N_21121,N_16704,N_12756);
or U21122 (N_21122,N_14967,N_19549);
nand U21123 (N_21123,N_10959,N_16918);
or U21124 (N_21124,N_10442,N_13407);
or U21125 (N_21125,N_10592,N_14654);
nand U21126 (N_21126,N_16158,N_19612);
or U21127 (N_21127,N_11235,N_11013);
xor U21128 (N_21128,N_18425,N_12564);
and U21129 (N_21129,N_11266,N_16368);
nor U21130 (N_21130,N_15852,N_15488);
xnor U21131 (N_21131,N_17196,N_14587);
nor U21132 (N_21132,N_10374,N_19979);
xor U21133 (N_21133,N_13433,N_11989);
and U21134 (N_21134,N_15428,N_13147);
and U21135 (N_21135,N_19926,N_14439);
or U21136 (N_21136,N_18558,N_15305);
xor U21137 (N_21137,N_13062,N_19063);
xnor U21138 (N_21138,N_16864,N_16038);
nor U21139 (N_21139,N_16464,N_10631);
or U21140 (N_21140,N_12854,N_12622);
xnor U21141 (N_21141,N_17246,N_14958);
xnor U21142 (N_21142,N_19405,N_19987);
or U21143 (N_21143,N_17635,N_12391);
xor U21144 (N_21144,N_18821,N_12953);
and U21145 (N_21145,N_12137,N_11504);
and U21146 (N_21146,N_17926,N_10883);
and U21147 (N_21147,N_10601,N_16113);
xor U21148 (N_21148,N_19729,N_17585);
nand U21149 (N_21149,N_13162,N_17479);
or U21150 (N_21150,N_11216,N_19794);
xnor U21151 (N_21151,N_11887,N_10777);
xnor U21152 (N_21152,N_15876,N_18623);
nand U21153 (N_21153,N_10036,N_13836);
nor U21154 (N_21154,N_16913,N_15400);
xnor U21155 (N_21155,N_13146,N_19032);
xnor U21156 (N_21156,N_12261,N_17054);
xor U21157 (N_21157,N_13465,N_15940);
nor U21158 (N_21158,N_11811,N_10840);
nor U21159 (N_21159,N_16796,N_16042);
nor U21160 (N_21160,N_13656,N_18172);
nor U21161 (N_21161,N_12393,N_11407);
nor U21162 (N_21162,N_19391,N_11636);
or U21163 (N_21163,N_15853,N_16347);
nand U21164 (N_21164,N_16055,N_13755);
or U21165 (N_21165,N_11186,N_12908);
and U21166 (N_21166,N_16640,N_19466);
and U21167 (N_21167,N_17228,N_13418);
xor U21168 (N_21168,N_18290,N_19975);
and U21169 (N_21169,N_15873,N_11229);
and U21170 (N_21170,N_12285,N_14807);
nor U21171 (N_21171,N_11680,N_10741);
nand U21172 (N_21172,N_14741,N_17650);
nor U21173 (N_21173,N_14923,N_16459);
nand U21174 (N_21174,N_14862,N_15954);
nor U21175 (N_21175,N_18305,N_14085);
nor U21176 (N_21176,N_17171,N_18981);
nor U21177 (N_21177,N_13305,N_13091);
nor U21178 (N_21178,N_18788,N_10820);
or U21179 (N_21179,N_15446,N_14288);
or U21180 (N_21180,N_13817,N_17106);
xnor U21181 (N_21181,N_11999,N_12667);
or U21182 (N_21182,N_17515,N_10098);
or U21183 (N_21183,N_14203,N_17932);
and U21184 (N_21184,N_17353,N_18511);
or U21185 (N_21185,N_14438,N_15085);
nor U21186 (N_21186,N_16967,N_11870);
xor U21187 (N_21187,N_16910,N_14767);
or U21188 (N_21188,N_11765,N_12056);
nor U21189 (N_21189,N_10211,N_18392);
nor U21190 (N_21190,N_10445,N_18645);
nor U21191 (N_21191,N_17440,N_13962);
nand U21192 (N_21192,N_11553,N_13748);
xnor U21193 (N_21193,N_12676,N_16923);
nor U21194 (N_21194,N_18970,N_16633);
nor U21195 (N_21195,N_13877,N_12260);
nand U21196 (N_21196,N_17656,N_11173);
or U21197 (N_21197,N_16028,N_11644);
and U21198 (N_21198,N_17433,N_11076);
nor U21199 (N_21199,N_11921,N_19711);
and U21200 (N_21200,N_12910,N_12758);
and U21201 (N_21201,N_17077,N_15223);
or U21202 (N_21202,N_15691,N_13446);
xor U21203 (N_21203,N_15110,N_15962);
or U21204 (N_21204,N_11510,N_19085);
nand U21205 (N_21205,N_16326,N_12976);
xor U21206 (N_21206,N_14422,N_18477);
and U21207 (N_21207,N_18079,N_14427);
xor U21208 (N_21208,N_19183,N_12781);
nor U21209 (N_21209,N_10240,N_14885);
xor U21210 (N_21210,N_18844,N_13337);
nand U21211 (N_21211,N_15721,N_18376);
xor U21212 (N_21212,N_11196,N_11138);
or U21213 (N_21213,N_16897,N_16036);
xor U21214 (N_21214,N_13914,N_17049);
nor U21215 (N_21215,N_16613,N_19066);
nand U21216 (N_21216,N_14214,N_14059);
and U21217 (N_21217,N_12904,N_13272);
or U21218 (N_21218,N_14305,N_10161);
and U21219 (N_21219,N_12245,N_16479);
and U21220 (N_21220,N_14498,N_17278);
xnor U21221 (N_21221,N_16421,N_19905);
nor U21222 (N_21222,N_15594,N_18730);
or U21223 (N_21223,N_19630,N_15855);
xor U21224 (N_21224,N_14022,N_13421);
nand U21225 (N_21225,N_10697,N_19702);
xnor U21226 (N_21226,N_17584,N_17733);
or U21227 (N_21227,N_18973,N_17473);
xor U21228 (N_21228,N_19195,N_11322);
or U21229 (N_21229,N_13398,N_18082);
nor U21230 (N_21230,N_19986,N_15772);
or U21231 (N_21231,N_19377,N_16635);
nor U21232 (N_21232,N_17601,N_12643);
and U21233 (N_21233,N_18129,N_13537);
nand U21234 (N_21234,N_13349,N_14493);
nand U21235 (N_21235,N_10203,N_10835);
xnor U21236 (N_21236,N_13857,N_12278);
and U21237 (N_21237,N_18568,N_16683);
xor U21238 (N_21238,N_12612,N_15430);
or U21239 (N_21239,N_14791,N_15591);
and U21240 (N_21240,N_10527,N_12901);
xor U21241 (N_21241,N_13886,N_11894);
nand U21242 (N_21242,N_10931,N_19839);
nor U21243 (N_21243,N_10460,N_14133);
or U21244 (N_21244,N_19403,N_15150);
or U21245 (N_21245,N_19070,N_17126);
and U21246 (N_21246,N_16962,N_12832);
or U21247 (N_21247,N_15567,N_10757);
or U21248 (N_21248,N_13583,N_13763);
xor U21249 (N_21249,N_10128,N_14067);
xor U21250 (N_21250,N_12353,N_12534);
nand U21251 (N_21251,N_17099,N_19893);
nor U21252 (N_21252,N_19825,N_16995);
nor U21253 (N_21253,N_10042,N_13298);
and U21254 (N_21254,N_12237,N_10117);
nand U21255 (N_21255,N_15011,N_18723);
nor U21256 (N_21256,N_13089,N_16203);
nand U21257 (N_21257,N_17602,N_15807);
nand U21258 (N_21258,N_18524,N_10944);
xnor U21259 (N_21259,N_17124,N_10141);
or U21260 (N_21260,N_10212,N_11668);
nor U21261 (N_21261,N_16346,N_13170);
and U21262 (N_21262,N_16211,N_17718);
nand U21263 (N_21263,N_11287,N_12107);
xnor U21264 (N_21264,N_18608,N_19990);
xnor U21265 (N_21265,N_16893,N_14060);
or U21266 (N_21266,N_15338,N_11293);
xor U21267 (N_21267,N_18410,N_14918);
or U21268 (N_21268,N_18470,N_13279);
nor U21269 (N_21269,N_10355,N_11682);
or U21270 (N_21270,N_10563,N_14428);
nor U21271 (N_21271,N_13524,N_10616);
or U21272 (N_21272,N_15689,N_11665);
or U21273 (N_21273,N_19200,N_19522);
nor U21274 (N_21274,N_19483,N_18474);
nand U21275 (N_21275,N_14551,N_17134);
and U21276 (N_21276,N_17405,N_18388);
or U21277 (N_21277,N_11867,N_11791);
nand U21278 (N_21278,N_16247,N_13315);
and U21279 (N_21279,N_14236,N_19123);
nor U21280 (N_21280,N_13188,N_12924);
or U21281 (N_21281,N_16000,N_10591);
nand U21282 (N_21282,N_15582,N_11639);
xnor U21283 (N_21283,N_15756,N_13536);
or U21284 (N_21284,N_10698,N_11367);
and U21285 (N_21285,N_18632,N_18900);
xor U21286 (N_21286,N_11547,N_17140);
nand U21287 (N_21287,N_13635,N_14996);
and U21288 (N_21288,N_12465,N_16614);
and U21289 (N_21289,N_18747,N_18035);
or U21290 (N_21290,N_19359,N_14640);
xor U21291 (N_21291,N_10784,N_19185);
and U21292 (N_21292,N_14253,N_14010);
and U21293 (N_21293,N_17809,N_15556);
nor U21294 (N_21294,N_10375,N_12099);
nor U21295 (N_21295,N_18277,N_11452);
xor U21296 (N_21296,N_12321,N_13818);
nor U21297 (N_21297,N_14162,N_14011);
nor U21298 (N_21298,N_17388,N_11968);
or U21299 (N_21299,N_14919,N_13025);
nor U21300 (N_21300,N_10045,N_12498);
and U21301 (N_21301,N_16035,N_14810);
or U21302 (N_21302,N_13095,N_17010);
nor U21303 (N_21303,N_19656,N_16734);
nor U21304 (N_21304,N_10286,N_14003);
or U21305 (N_21305,N_12716,N_18861);
nand U21306 (N_21306,N_12445,N_17991);
xnor U21307 (N_21307,N_12753,N_11986);
nor U21308 (N_21308,N_11980,N_10808);
nand U21309 (N_21309,N_16034,N_12170);
nand U21310 (N_21310,N_19849,N_10744);
xnor U21311 (N_21311,N_17912,N_17200);
nor U21312 (N_21312,N_18432,N_18720);
nor U21313 (N_21313,N_14611,N_12344);
xor U21314 (N_21314,N_10752,N_16826);
nor U21315 (N_21315,N_17358,N_15770);
nand U21316 (N_21316,N_11402,N_18429);
or U21317 (N_21317,N_12182,N_11264);
nand U21318 (N_21318,N_16985,N_10856);
xnor U21319 (N_21319,N_17516,N_14367);
or U21320 (N_21320,N_13677,N_15107);
xnor U21321 (N_21321,N_11391,N_13964);
nor U21322 (N_21322,N_16256,N_16699);
nor U21323 (N_21323,N_16574,N_13634);
nand U21324 (N_21324,N_10887,N_15179);
nand U21325 (N_21325,N_16148,N_15667);
or U21326 (N_21326,N_15902,N_18734);
nor U21327 (N_21327,N_19861,N_12209);
nor U21328 (N_21328,N_11082,N_10313);
or U21329 (N_21329,N_12228,N_12983);
xor U21330 (N_21330,N_15626,N_18881);
xnor U21331 (N_21331,N_13768,N_14118);
nand U21332 (N_21332,N_12469,N_15236);
nand U21333 (N_21333,N_15198,N_12958);
nand U21334 (N_21334,N_12675,N_17861);
nor U21335 (N_21335,N_12510,N_11822);
nor U21336 (N_21336,N_10622,N_13404);
nor U21337 (N_21337,N_19557,N_11591);
nor U21338 (N_21338,N_17833,N_15254);
or U21339 (N_21339,N_13636,N_11674);
or U21340 (N_21340,N_13977,N_10410);
nand U21341 (N_21341,N_18255,N_12645);
xnor U21342 (N_21342,N_10761,N_16359);
and U21343 (N_21343,N_15505,N_10517);
and U21344 (N_21344,N_13940,N_17198);
and U21345 (N_21345,N_10097,N_11499);
or U21346 (N_21346,N_18890,N_15966);
nor U21347 (N_21347,N_10187,N_14310);
nand U21348 (N_21348,N_18784,N_12120);
xnor U21349 (N_21349,N_13767,N_15930);
nand U21350 (N_21350,N_14313,N_18865);
nor U21351 (N_21351,N_14567,N_18766);
or U21352 (N_21352,N_10590,N_14109);
or U21353 (N_21353,N_17025,N_16631);
or U21354 (N_21354,N_11734,N_15437);
nand U21355 (N_21355,N_11011,N_12621);
nand U21356 (N_21356,N_12379,N_19096);
or U21357 (N_21357,N_12358,N_12242);
nand U21358 (N_21358,N_11997,N_14201);
xor U21359 (N_21359,N_13345,N_15165);
nand U21360 (N_21360,N_18729,N_15936);
or U21361 (N_21361,N_14206,N_15337);
and U21362 (N_21362,N_10288,N_13204);
xor U21363 (N_21363,N_18946,N_16033);
xor U21364 (N_21364,N_19837,N_14352);
nor U21365 (N_21365,N_12089,N_18657);
or U21366 (N_21366,N_11304,N_11594);
or U21367 (N_21367,N_15162,N_13228);
xnor U21368 (N_21368,N_11122,N_19983);
nand U21369 (N_21369,N_13924,N_10035);
nor U21370 (N_21370,N_14659,N_12179);
and U21371 (N_21371,N_14554,N_15844);
and U21372 (N_21372,N_16442,N_18090);
xnor U21373 (N_21373,N_12724,N_10556);
nand U21374 (N_21374,N_17598,N_14023);
nand U21375 (N_21375,N_11545,N_19590);
xor U21376 (N_21376,N_18813,N_13787);
nand U21377 (N_21377,N_10648,N_18757);
nand U21378 (N_21378,N_18327,N_15048);
nand U21379 (N_21379,N_15878,N_12942);
nand U21380 (N_21380,N_10618,N_10281);
nand U21381 (N_21381,N_16235,N_19791);
and U21382 (N_21382,N_14562,N_13827);
xnor U21383 (N_21383,N_17482,N_15637);
or U21384 (N_21384,N_17103,N_17264);
nand U21385 (N_21385,N_16603,N_13960);
nor U21386 (N_21386,N_15242,N_14750);
and U21387 (N_21387,N_12373,N_13459);
or U21388 (N_21388,N_14555,N_18350);
and U21389 (N_21389,N_19212,N_18395);
or U21390 (N_21390,N_14437,N_14574);
or U21391 (N_21391,N_15132,N_11551);
and U21392 (N_21392,N_10685,N_15668);
and U21393 (N_21393,N_14634,N_13800);
or U21394 (N_21394,N_18284,N_12703);
nor U21395 (N_21395,N_19597,N_16351);
nand U21396 (N_21396,N_17177,N_16777);
xnor U21397 (N_21397,N_15466,N_19663);
and U21398 (N_21398,N_16212,N_17271);
nand U21399 (N_21399,N_14856,N_16496);
nor U21400 (N_21400,N_12356,N_18581);
nand U21401 (N_21401,N_18158,N_13161);
xnor U21402 (N_21402,N_15120,N_18678);
or U21403 (N_21403,N_18618,N_16584);
nor U21404 (N_21404,N_12681,N_10911);
nand U21405 (N_21405,N_10213,N_11126);
nor U21406 (N_21406,N_16709,N_14705);
nand U21407 (N_21407,N_15605,N_15365);
nor U21408 (N_21408,N_14233,N_12210);
xor U21409 (N_21409,N_12831,N_14057);
nor U21410 (N_21410,N_16943,N_16074);
and U21411 (N_21411,N_11618,N_13392);
nand U21412 (N_21412,N_17691,N_18435);
or U21413 (N_21413,N_16411,N_13714);
and U21414 (N_21414,N_13784,N_11773);
nor U21415 (N_21415,N_15429,N_12422);
and U21416 (N_21416,N_13243,N_11288);
nand U21417 (N_21417,N_18036,N_16771);
and U21418 (N_21418,N_14041,N_10523);
or U21419 (N_21419,N_12076,N_12313);
nor U21420 (N_21420,N_12699,N_11991);
nand U21421 (N_21421,N_12259,N_10902);
nand U21422 (N_21422,N_16318,N_10177);
xnor U21423 (N_21423,N_14395,N_17902);
and U21424 (N_21424,N_15113,N_19504);
nand U21425 (N_21425,N_18602,N_17459);
nor U21426 (N_21426,N_10916,N_16537);
nor U21427 (N_21427,N_19278,N_14338);
or U21428 (N_21428,N_19092,N_10960);
and U21429 (N_21429,N_19314,N_10570);
or U21430 (N_21430,N_11847,N_14237);
or U21431 (N_21431,N_11992,N_18771);
and U21432 (N_21432,N_13050,N_11604);
nor U21433 (N_21433,N_19892,N_12852);
and U21434 (N_21434,N_18665,N_15186);
nor U21435 (N_21435,N_13675,N_11981);
nor U21436 (N_21436,N_18592,N_17132);
nand U21437 (N_21437,N_15054,N_15980);
or U21438 (N_21438,N_19858,N_15451);
and U21439 (N_21439,N_18817,N_18231);
or U21440 (N_21440,N_19146,N_14375);
nor U21441 (N_21441,N_11738,N_12525);
and U21442 (N_21442,N_18944,N_14446);
or U21443 (N_21443,N_18163,N_10933);
xor U21444 (N_21444,N_16444,N_16576);
nand U21445 (N_21445,N_11210,N_11399);
nor U21446 (N_21446,N_17538,N_18240);
xnor U21447 (N_21447,N_16610,N_19237);
nand U21448 (N_21448,N_14189,N_19230);
and U21449 (N_21449,N_12819,N_11807);
nand U21450 (N_21450,N_13085,N_18748);
nor U21451 (N_21451,N_10054,N_10418);
nor U21452 (N_21452,N_18038,N_14046);
or U21453 (N_21453,N_12655,N_18182);
or U21454 (N_21454,N_19697,N_14301);
and U21455 (N_21455,N_19172,N_14275);
or U21456 (N_21456,N_15233,N_17887);
nand U21457 (N_21457,N_16073,N_12866);
or U21458 (N_21458,N_15401,N_14244);
nor U21459 (N_21459,N_18269,N_11167);
or U21460 (N_21460,N_18487,N_16004);
or U21461 (N_21461,N_15562,N_16499);
or U21462 (N_21462,N_15355,N_13454);
and U21463 (N_21463,N_19214,N_14670);
and U21464 (N_21464,N_17938,N_11025);
xnor U21465 (N_21465,N_13998,N_17266);
xnor U21466 (N_21466,N_17661,N_13250);
and U21467 (N_21467,N_11892,N_18845);
and U21468 (N_21468,N_10667,N_10589);
and U21469 (N_21469,N_12606,N_16207);
xnor U21470 (N_21470,N_10370,N_19570);
nor U21471 (N_21471,N_15819,N_18917);
nand U21472 (N_21472,N_10484,N_16517);
xnor U21473 (N_21473,N_11716,N_16611);
nand U21474 (N_21474,N_12685,N_16801);
and U21475 (N_21475,N_12155,N_13936);
nand U21476 (N_21476,N_18217,N_17815);
nand U21477 (N_21477,N_14954,N_15879);
nand U21478 (N_21478,N_11027,N_13045);
nand U21479 (N_21479,N_13430,N_17763);
nor U21480 (N_21480,N_10620,N_17116);
and U21481 (N_21481,N_14717,N_14624);
or U21482 (N_21482,N_16334,N_17592);
nor U21483 (N_21483,N_12627,N_18627);
nand U21484 (N_21484,N_19189,N_13213);
xnor U21485 (N_21485,N_19972,N_18258);
xor U21486 (N_21486,N_11467,N_14440);
or U21487 (N_21487,N_12690,N_19976);
nand U21488 (N_21488,N_15828,N_12647);
nor U21489 (N_21489,N_12162,N_14978);
nor U21490 (N_21490,N_18193,N_17660);
nand U21491 (N_21491,N_15087,N_19501);
and U21492 (N_21492,N_13297,N_17627);
xor U21493 (N_21493,N_15782,N_10314);
nand U21494 (N_21494,N_12338,N_16802);
nand U21495 (N_21495,N_11345,N_16164);
or U21496 (N_21496,N_10810,N_10291);
nor U21497 (N_21497,N_10783,N_11099);
and U21498 (N_21498,N_13346,N_10737);
or U21499 (N_21499,N_11419,N_19473);
nor U21500 (N_21500,N_19470,N_17313);
nor U21501 (N_21501,N_15487,N_16728);
xor U21502 (N_21502,N_10888,N_11804);
or U21503 (N_21503,N_15530,N_18939);
and U21504 (N_21504,N_15423,N_14269);
or U21505 (N_21505,N_11653,N_15049);
xor U21506 (N_21506,N_11239,N_16154);
xor U21507 (N_21507,N_17983,N_10451);
xor U21508 (N_21508,N_16953,N_19889);
or U21509 (N_21509,N_10565,N_16381);
nor U21510 (N_21510,N_14409,N_17486);
or U21511 (N_21511,N_15478,N_14752);
nor U21512 (N_21512,N_16112,N_17509);
and U21513 (N_21513,N_17066,N_16510);
nor U21514 (N_21514,N_18335,N_12539);
nand U21515 (N_21515,N_12909,N_10597);
nand U21516 (N_21516,N_18557,N_15108);
xnor U21517 (N_21517,N_13172,N_14881);
nor U21518 (N_21518,N_15393,N_11841);
nand U21519 (N_21519,N_10947,N_17605);
xnor U21520 (N_21520,N_12306,N_18007);
nor U21521 (N_21521,N_14208,N_12656);
nor U21522 (N_21522,N_12566,N_16775);
and U21523 (N_21523,N_19757,N_16788);
and U21524 (N_21524,N_15864,N_17971);
nand U21525 (N_21525,N_16335,N_18430);
nor U21526 (N_21526,N_10319,N_13245);
and U21527 (N_21527,N_15285,N_13351);
nand U21528 (N_21528,N_12466,N_15867);
nor U21529 (N_21529,N_11360,N_10600);
xnor U21530 (N_21530,N_13724,N_10787);
nor U21531 (N_21531,N_11064,N_13276);
and U21532 (N_21532,N_19141,N_11712);
and U21533 (N_21533,N_17966,N_16678);
nand U21534 (N_21534,N_11369,N_19554);
nor U21535 (N_21535,N_14141,N_17996);
and U21536 (N_21536,N_10604,N_13004);
nand U21537 (N_21537,N_14219,N_19406);
or U21538 (N_21538,N_13708,N_17819);
xnor U21539 (N_21539,N_13341,N_13769);
and U21540 (N_21540,N_17676,N_18781);
nor U21541 (N_21541,N_11602,N_16700);
nor U21542 (N_21542,N_17466,N_12091);
and U21543 (N_21543,N_16719,N_15539);
xor U21544 (N_21544,N_19276,N_19238);
or U21545 (N_21545,N_15793,N_16232);
and U21546 (N_21546,N_14734,N_14053);
nor U21547 (N_21547,N_10168,N_16666);
and U21548 (N_21548,N_19282,N_16476);
or U21549 (N_21549,N_13706,N_19525);
or U21550 (N_21550,N_18373,N_17071);
or U21551 (N_21551,N_16320,N_17818);
nand U21552 (N_21552,N_10580,N_11151);
nor U21553 (N_21553,N_12962,N_14001);
nand U21554 (N_21554,N_14772,N_13602);
or U21555 (N_21555,N_10219,N_12227);
nand U21556 (N_21556,N_16867,N_16540);
xor U21557 (N_21557,N_19726,N_15029);
and U21558 (N_21558,N_13082,N_15948);
and U21559 (N_21559,N_19251,N_10845);
xnor U21560 (N_21560,N_12704,N_11213);
nor U21561 (N_21561,N_17234,N_17382);
nor U21562 (N_21562,N_13445,N_14854);
nand U21563 (N_21563,N_15729,N_11609);
nor U21564 (N_21564,N_10380,N_14537);
nor U21565 (N_21565,N_16238,N_15982);
and U21566 (N_21566,N_16215,N_12213);
or U21567 (N_21567,N_19499,N_10234);
xnor U21568 (N_21568,N_14550,N_15006);
and U21569 (N_21569,N_19716,N_17122);
nand U21570 (N_21570,N_18121,N_18656);
nand U21571 (N_21571,N_15156,N_11763);
and U21572 (N_21572,N_15449,N_15841);
xnor U21573 (N_21573,N_16676,N_16177);
and U21574 (N_21574,N_11263,N_17331);
nand U21575 (N_21575,N_11574,N_11939);
nand U21576 (N_21576,N_12281,N_14804);
or U21577 (N_21577,N_11042,N_17897);
nor U21578 (N_21578,N_14316,N_16843);
nor U21579 (N_21579,N_15713,N_18110);
and U21580 (N_21580,N_13872,N_16272);
or U21581 (N_21581,N_14472,N_10477);
nor U21582 (N_21582,N_12805,N_10585);
nor U21583 (N_21583,N_12174,N_12882);
or U21584 (N_21584,N_16361,N_10668);
and U21585 (N_21585,N_10815,N_14207);
xnor U21586 (N_21586,N_15743,N_13021);
and U21587 (N_21587,N_13597,N_11392);
or U21588 (N_21588,N_14901,N_16291);
nand U21589 (N_21589,N_16287,N_17852);
nor U21590 (N_21590,N_19074,N_17323);
nand U21591 (N_21591,N_14855,N_10175);
nand U21592 (N_21592,N_17964,N_11006);
nor U21593 (N_21593,N_13641,N_10566);
and U21594 (N_21594,N_12888,N_10579);
nand U21595 (N_21595,N_14730,N_19888);
nor U21596 (N_21596,N_15394,N_13464);
and U21597 (N_21597,N_15960,N_16929);
or U21598 (N_21598,N_19852,N_19118);
nand U21599 (N_21599,N_14283,N_19427);
and U21600 (N_21600,N_12399,N_14307);
nor U21601 (N_21601,N_13556,N_12951);
nand U21602 (N_21602,N_10133,N_13403);
xor U21603 (N_21603,N_11073,N_17958);
nand U21604 (N_21604,N_15696,N_19272);
nor U21605 (N_21605,N_14477,N_19289);
or U21606 (N_21606,N_10384,N_14000);
xor U21607 (N_21607,N_16044,N_14740);
nand U21608 (N_21608,N_15537,N_10230);
and U21609 (N_21609,N_18406,N_19091);
and U21610 (N_21610,N_14539,N_17428);
and U21611 (N_21611,N_16441,N_10426);
and U21612 (N_21612,N_13068,N_19847);
nor U21613 (N_21613,N_13086,N_17095);
and U21614 (N_21614,N_19508,N_18597);
nand U21615 (N_21615,N_11048,N_10750);
or U21616 (N_21616,N_12072,N_15230);
nor U21617 (N_21617,N_15672,N_18517);
or U21618 (N_21618,N_18499,N_19244);
or U21619 (N_21619,N_12194,N_14745);
xnor U21620 (N_21620,N_16024,N_14547);
xnor U21621 (N_21621,N_16399,N_10954);
nor U21622 (N_21622,N_15847,N_10669);
xnor U21623 (N_21623,N_12246,N_12461);
nand U21624 (N_21624,N_17350,N_15425);
nand U21625 (N_21625,N_15999,N_12707);
nor U21626 (N_21626,N_15082,N_12840);
and U21627 (N_21627,N_18974,N_14553);
nor U21628 (N_21628,N_18777,N_18829);
nand U21629 (N_21629,N_12994,N_10053);
or U21630 (N_21630,N_11725,N_11996);
xnor U21631 (N_21631,N_13103,N_14598);
and U21632 (N_21632,N_18814,N_11412);
nor U21633 (N_21633,N_18662,N_19535);
nand U21634 (N_21634,N_11950,N_12728);
xnor U21635 (N_21635,N_14130,N_17760);
and U21636 (N_21636,N_18307,N_14722);
nand U21637 (N_21637,N_18715,N_11656);
and U21638 (N_21638,N_18242,N_18324);
and U21639 (N_21639,N_14839,N_14627);
nor U21640 (N_21640,N_13058,N_14254);
nor U21641 (N_21641,N_17411,N_12095);
xor U21642 (N_21642,N_19742,N_11112);
nor U21643 (N_21643,N_17005,N_18072);
xor U21644 (N_21644,N_15700,N_19245);
and U21645 (N_21645,N_12872,N_10081);
nor U21646 (N_21646,N_14768,N_14412);
or U21647 (N_21647,N_11596,N_13375);
nand U21648 (N_21648,N_11350,N_11519);
nand U21649 (N_21649,N_16407,N_12318);
and U21650 (N_21650,N_19966,N_16331);
xnor U21651 (N_21651,N_10306,N_17267);
and U21652 (N_21652,N_14803,N_14779);
nor U21653 (N_21653,N_15197,N_17724);
nor U21654 (N_21654,N_15677,N_19269);
and U21655 (N_21655,N_14955,N_10046);
nor U21656 (N_21656,N_10360,N_16707);
nand U21657 (N_21657,N_12414,N_14278);
nand U21658 (N_21658,N_10401,N_12773);
nor U21659 (N_21659,N_18054,N_19528);
or U21660 (N_21660,N_11019,N_14302);
and U21661 (N_21661,N_18737,N_15493);
nand U21662 (N_21662,N_14255,N_17600);
or U21663 (N_21663,N_14366,N_12920);
nand U21664 (N_21664,N_11449,N_15484);
nor U21665 (N_21665,N_19036,N_17766);
or U21666 (N_21666,N_17531,N_17173);
or U21667 (N_21667,N_16139,N_11995);
xor U21668 (N_21668,N_16556,N_11909);
and U21669 (N_21669,N_11232,N_12441);
nor U21670 (N_21670,N_19295,N_15326);
nand U21671 (N_21671,N_15560,N_18763);
nor U21672 (N_21672,N_14249,N_14380);
or U21673 (N_21673,N_13621,N_11015);
xor U21674 (N_21674,N_11881,N_17711);
and U21675 (N_21675,N_15253,N_18381);
nor U21676 (N_21676,N_18419,N_11546);
nand U21677 (N_21677,N_13129,N_10789);
and U21678 (N_21678,N_17729,N_12049);
or U21679 (N_21679,N_17513,N_16776);
or U21680 (N_21680,N_15265,N_12198);
nand U21681 (N_21681,N_10758,N_15389);
and U21682 (N_21682,N_19530,N_17448);
and U21683 (N_21683,N_19778,N_13968);
xnor U21684 (N_21684,N_14578,N_18118);
and U21685 (N_21685,N_12876,N_17195);
and U21686 (N_21686,N_14853,N_18767);
nor U21687 (N_21687,N_17067,N_12141);
or U21688 (N_21688,N_19533,N_11830);
or U21689 (N_21689,N_12124,N_16376);
nand U21690 (N_21690,N_10024,N_18503);
nand U21691 (N_21691,N_15390,N_16019);
nand U21692 (N_21692,N_15612,N_12650);
nor U21693 (N_21693,N_15906,N_17359);
nor U21694 (N_21694,N_17866,N_14771);
or U21695 (N_21695,N_17847,N_16594);
nand U21696 (N_21696,N_13770,N_17414);
nor U21697 (N_21697,N_19055,N_11388);
or U21698 (N_21698,N_12668,N_11225);
nand U21699 (N_21699,N_19240,N_12332);
xor U21700 (N_21700,N_11565,N_19441);
xor U21701 (N_21701,N_15259,N_14605);
or U21702 (N_21702,N_17830,N_12397);
xor U21703 (N_21703,N_10923,N_16170);
xnor U21704 (N_21704,N_10038,N_13156);
nand U21705 (N_21705,N_15686,N_14735);
or U21706 (N_21706,N_12544,N_11035);
nor U21707 (N_21707,N_16857,N_12786);
nand U21708 (N_21708,N_11404,N_13108);
and U21709 (N_21709,N_14196,N_10318);
and U21710 (N_21710,N_17977,N_17628);
nand U21711 (N_21711,N_15507,N_15518);
nor U21712 (N_21712,N_14262,N_11097);
xnor U21713 (N_21713,N_13622,N_11524);
nor U21714 (N_21714,N_18031,N_16369);
or U21715 (N_21715,N_17384,N_13653);
xor U21716 (N_21716,N_12744,N_12046);
or U21717 (N_21717,N_18759,N_15243);
nand U21718 (N_21718,N_15361,N_11031);
xnor U21719 (N_21719,N_17698,N_15569);
xor U21720 (N_21720,N_15631,N_16432);
and U21721 (N_21721,N_14075,N_14744);
and U21722 (N_21722,N_10440,N_11319);
and U21723 (N_21723,N_15211,N_16585);
or U21724 (N_21724,N_10880,N_19725);
nor U21725 (N_21725,N_19209,N_15398);
nor U21726 (N_21726,N_17320,N_13262);
nand U21727 (N_21727,N_13471,N_14773);
nand U21728 (N_21728,N_15831,N_17302);
and U21729 (N_21729,N_12597,N_14341);
and U21730 (N_21730,N_15623,N_17800);
xor U21731 (N_21731,N_11056,N_10056);
nand U21732 (N_21732,N_14617,N_16800);
nand U21733 (N_21733,N_14827,N_10468);
nor U21734 (N_21734,N_18420,N_13907);
or U21735 (N_21735,N_10143,N_13044);
or U21736 (N_21736,N_19666,N_14890);
xnor U21737 (N_21737,N_15358,N_10025);
or U21738 (N_21738,N_16946,N_19517);
xor U21739 (N_21739,N_11711,N_18752);
nand U21740 (N_21740,N_10069,N_13441);
nand U21741 (N_21741,N_16583,N_11998);
nand U21742 (N_21742,N_10002,N_11498);
nor U21743 (N_21743,N_17573,N_10575);
nor U21744 (N_21744,N_10739,N_15744);
and U21745 (N_21745,N_11171,N_15330);
and U21746 (N_21746,N_15943,N_15296);
xnor U21747 (N_21747,N_14384,N_17634);
or U21748 (N_21748,N_12327,N_19330);
nor U21749 (N_21749,N_12269,N_10475);
xnor U21750 (N_21750,N_18351,N_11527);
xor U21751 (N_21751,N_13302,N_11003);
nor U21752 (N_21752,N_10780,N_18800);
nand U21753 (N_21753,N_11851,N_19660);
xor U21754 (N_21754,N_14054,N_16875);
and U21755 (N_21755,N_11243,N_17788);
nand U21756 (N_21756,N_17864,N_17609);
xor U21757 (N_21757,N_18247,N_16485);
and U21758 (N_21758,N_13922,N_13625);
nor U21759 (N_21759,N_11994,N_16306);
xnor U21760 (N_21760,N_16991,N_19052);
and U21761 (N_21761,N_18547,N_17425);
or U21762 (N_21762,N_14418,N_10080);
nand U21763 (N_21763,N_11257,N_10718);
and U21764 (N_21764,N_12858,N_11891);
nor U21765 (N_21765,N_14820,N_19343);
xnor U21766 (N_21766,N_13726,N_15977);
nor U21767 (N_21767,N_10062,N_18626);
nor U21768 (N_21768,N_17362,N_19051);
xor U21769 (N_21769,N_11132,N_10544);
or U21770 (N_21770,N_13670,N_16636);
xor U21771 (N_21771,N_10461,N_16161);
and U21772 (N_21772,N_15040,N_13734);
xor U21773 (N_21773,N_16527,N_16886);
and U21774 (N_21774,N_16822,N_10345);
nor U21775 (N_21775,N_12782,N_19903);
nor U21776 (N_21776,N_19281,N_10925);
and U21777 (N_21777,N_16619,N_17812);
xor U21778 (N_21778,N_13432,N_15654);
and U21779 (N_21779,N_18765,N_15599);
nor U21780 (N_21780,N_12410,N_11970);
nor U21781 (N_21781,N_19519,N_14056);
and U21782 (N_21782,N_16513,N_10502);
nor U21783 (N_21783,N_13153,N_14559);
nor U21784 (N_21784,N_13523,N_13419);
or U21785 (N_21785,N_15278,N_16415);
and U21786 (N_21786,N_17873,N_15984);
nor U21787 (N_21787,N_13241,N_14374);
nor U21788 (N_21788,N_15086,N_15995);
xor U21789 (N_21789,N_11153,N_13385);
nand U21790 (N_21790,N_11466,N_11058);
xor U21791 (N_21791,N_17989,N_11270);
nor U21792 (N_21792,N_14014,N_11017);
or U21793 (N_21793,N_13314,N_11277);
nor U21794 (N_21794,N_16093,N_16168);
nand U21795 (N_21795,N_16053,N_15123);
nand U21796 (N_21796,N_16069,N_17506);
or U21797 (N_21797,N_12774,N_18196);
nand U21798 (N_21798,N_10948,N_10174);
or U21799 (N_21799,N_14621,N_16388);
and U21800 (N_21800,N_19743,N_18272);
nand U21801 (N_21801,N_18593,N_14637);
or U21802 (N_21802,N_14620,N_16166);
nand U21803 (N_21803,N_13644,N_10666);
xnor U21804 (N_21804,N_17567,N_17276);
xor U21805 (N_21805,N_12123,N_12325);
nand U21806 (N_21806,N_10473,N_13563);
nand U21807 (N_21807,N_14327,N_13917);
nor U21808 (N_21808,N_14006,N_16380);
xnor U21809 (N_21809,N_14042,N_14995);
or U21810 (N_21810,N_11470,N_10120);
nor U21811 (N_21811,N_13662,N_13159);
xnor U21812 (N_21812,N_14984,N_16874);
xor U21813 (N_21813,N_12157,N_14838);
nand U21814 (N_21814,N_11124,N_16752);
or U21815 (N_21815,N_13874,N_15227);
xor U21816 (N_21816,N_14813,N_14980);
and U21817 (N_21817,N_10640,N_10331);
or U21818 (N_21818,N_18731,N_18846);
xor U21819 (N_21819,N_12185,N_17252);
nor U21820 (N_21820,N_16064,N_10991);
nor U21821 (N_21821,N_16898,N_17295);
nand U21822 (N_21822,N_15514,N_18631);
and U21823 (N_21823,N_18293,N_13972);
or U21824 (N_21824,N_13566,N_17827);
xnor U21825 (N_21825,N_17042,N_10122);
nor U21826 (N_21826,N_14864,N_14836);
or U21827 (N_21827,N_15727,N_18145);
and U21828 (N_21828,N_13397,N_13190);
nor U21829 (N_21829,N_14623,N_18915);
nand U21830 (N_21830,N_18993,N_14381);
xor U21831 (N_21831,N_11954,N_18133);
or U21832 (N_21832,N_17941,N_14817);
nand U21833 (N_21833,N_17734,N_17980);
or U21834 (N_21834,N_13076,N_10628);
nand U21835 (N_21835,N_16404,N_10704);
nand U21836 (N_21836,N_14081,N_10480);
nor U21837 (N_21837,N_16715,N_17114);
and U21838 (N_21838,N_15593,N_19017);
nand U21839 (N_21839,N_17268,N_17487);
nand U21840 (N_21840,N_12658,N_19943);
nand U21841 (N_21841,N_17998,N_17642);
nand U21842 (N_21842,N_11422,N_19186);
or U21843 (N_21843,N_17436,N_10095);
or U21844 (N_21844,N_16949,N_18286);
xor U21845 (N_21845,N_16436,N_11694);
and U21846 (N_21846,N_12848,N_13120);
or U21847 (N_21847,N_10454,N_10542);
nand U21848 (N_21848,N_10705,N_15875);
xor U21849 (N_21849,N_10090,N_18122);
or U21850 (N_21850,N_14348,N_14732);
or U21851 (N_21851,N_16364,N_13265);
or U21852 (N_21852,N_13695,N_13852);
xnor U21853 (N_21853,N_15701,N_13078);
or U21854 (N_21854,N_14657,N_12075);
or U21855 (N_21855,N_14796,N_14191);
or U21856 (N_21856,N_15927,N_11854);
nor U21857 (N_21857,N_13947,N_15269);
or U21858 (N_21858,N_11619,N_19026);
xnor U21859 (N_21859,N_18624,N_10083);
or U21860 (N_21860,N_12268,N_19288);
and U21861 (N_21861,N_18092,N_11072);
and U21862 (N_21862,N_12741,N_15164);
nand U21863 (N_21863,N_13720,N_19552);
or U21864 (N_21864,N_10293,N_16588);
xnor U21865 (N_21865,N_18804,N_19354);
nor U21866 (N_21866,N_18156,N_10073);
or U21867 (N_21867,N_18676,N_17056);
nand U21868 (N_21868,N_14573,N_13658);
nor U21869 (N_21869,N_10871,N_16504);
xnor U21870 (N_21870,N_17179,N_19083);
nand U21871 (N_21871,N_11416,N_15910);
or U21872 (N_21872,N_15693,N_15129);
nand U21873 (N_21873,N_16373,N_12406);
nand U21874 (N_21874,N_15513,N_10032);
xor U21875 (N_21875,N_16542,N_17536);
xor U21876 (N_21876,N_16841,N_16079);
nand U21877 (N_21877,N_14990,N_14593);
xor U21878 (N_21878,N_11785,N_19361);
nor U21879 (N_21879,N_13230,N_10197);
or U21880 (N_21880,N_15935,N_18761);
nor U21881 (N_21881,N_15716,N_16071);
and U21882 (N_21882,N_15951,N_18758);
nor U21883 (N_21883,N_14724,N_17606);
nor U21884 (N_21884,N_15240,N_12605);
nor U21885 (N_21885,N_18112,N_17299);
and U21886 (N_21886,N_10358,N_12158);
nor U21887 (N_21887,N_16765,N_15970);
xor U21888 (N_21888,N_18162,N_13911);
nand U21889 (N_21889,N_12590,N_12446);
nand U21890 (N_21890,N_11356,N_10740);
or U21891 (N_21891,N_11561,N_19098);
nor U21892 (N_21892,N_10493,N_17210);
nor U21893 (N_21893,N_11403,N_10407);
and U21894 (N_21894,N_13212,N_17022);
xnor U21895 (N_21895,N_11326,N_14336);
nand U21896 (N_21896,N_16878,N_18473);
or U21897 (N_21897,N_17855,N_10699);
xnor U21898 (N_21898,N_13402,N_14421);
and U21899 (N_21899,N_12192,N_11188);
nand U21900 (N_21900,N_19239,N_11176);
xor U21901 (N_21901,N_17032,N_19058);
xor U21902 (N_21902,N_16813,N_17170);
nand U21903 (N_21903,N_14959,N_16774);
nand U21904 (N_21904,N_19569,N_10736);
nand U21905 (N_21905,N_15973,N_12847);
nand U21906 (N_21906,N_19506,N_13173);
nor U21907 (N_21907,N_16175,N_10193);
or U21908 (N_21908,N_14078,N_15091);
and U21909 (N_21909,N_19380,N_10636);
nand U21910 (N_21910,N_15161,N_12828);
and U21911 (N_21911,N_11115,N_10327);
nor U21912 (N_21912,N_10854,N_15480);
nand U21913 (N_21913,N_15009,N_11835);
nand U21914 (N_21914,N_13388,N_19084);
xor U21915 (N_21915,N_12345,N_11828);
xnor U21916 (N_21916,N_13423,N_14349);
xor U21917 (N_21917,N_15185,N_13513);
and U21918 (N_21918,N_19616,N_10678);
nor U21919 (N_21919,N_14580,N_12654);
or U21920 (N_21920,N_19547,N_17260);
nand U21921 (N_21921,N_14015,N_18677);
or U21922 (N_21922,N_10594,N_13624);
nand U21923 (N_21923,N_17275,N_12833);
and U21924 (N_21924,N_17381,N_14974);
xnor U21925 (N_21925,N_11034,N_11203);
nand U21926 (N_21926,N_12763,N_13301);
nand U21927 (N_21927,N_14570,N_10491);
or U21928 (N_21928,N_13730,N_18137);
xnor U21929 (N_21929,N_12524,N_15837);
nand U21930 (N_21930,N_19503,N_15842);
and U21931 (N_21931,N_13642,N_18294);
or U21932 (N_21932,N_18443,N_17340);
nand U21933 (N_21933,N_11420,N_13289);
xnor U21934 (N_21934,N_19982,N_15147);
xnor U21935 (N_21935,N_17148,N_13252);
xor U21936 (N_21936,N_11028,N_13370);
nand U21937 (N_21937,N_11247,N_13885);
nor U21938 (N_21938,N_13762,N_14306);
and U21939 (N_21939,N_12166,N_11622);
or U21940 (N_21940,N_13069,N_11349);
nor U21941 (N_21941,N_11039,N_12008);
or U21942 (N_21942,N_16104,N_13084);
nand U21943 (N_21943,N_19550,N_19150);
nand U21944 (N_21944,N_16577,N_18527);
or U21945 (N_21945,N_18978,N_19444);
nand U21946 (N_21946,N_15273,N_14379);
nand U21947 (N_21947,N_19701,N_12030);
nor U21948 (N_21948,N_15249,N_18198);
or U21949 (N_21949,N_15422,N_13264);
or U21950 (N_21950,N_17799,N_17577);
xor U21951 (N_21951,N_17821,N_10689);
xor U21952 (N_21952,N_13981,N_14557);
nor U21953 (N_21953,N_19336,N_11690);
nor U21954 (N_21954,N_10496,N_10949);
or U21955 (N_21955,N_19601,N_14267);
or U21956 (N_21956,N_15712,N_18379);
or U21957 (N_21957,N_14868,N_19228);
or U21958 (N_21958,N_17096,N_19182);
nor U21959 (N_21959,N_16859,N_11654);
nor U21960 (N_21960,N_19885,N_19911);
or U21961 (N_21961,N_11536,N_16282);
nand U21962 (N_21962,N_17565,N_18549);
nor U21963 (N_21963,N_13194,N_12161);
nand U21964 (N_21964,N_17327,N_11634);
and U21965 (N_21965,N_11810,N_15310);
and U21966 (N_21966,N_18322,N_17130);
or U21967 (N_21967,N_18084,N_11513);
xor U21968 (N_21968,N_12915,N_10467);
or U21969 (N_21969,N_18480,N_16764);
and U21970 (N_21970,N_11199,N_12748);
nand U21971 (N_21971,N_14865,N_12421);
xnor U21972 (N_21972,N_15461,N_12821);
and U21973 (N_21973,N_15545,N_15903);
nand U21974 (N_21974,N_18033,N_11492);
or U21975 (N_21975,N_16400,N_13698);
xor U21976 (N_21976,N_19192,N_11832);
nand U21977 (N_21977,N_13041,N_14867);
or U21978 (N_21978,N_16405,N_11191);
nand U21979 (N_21979,N_12239,N_14683);
xor U21980 (N_21980,N_18931,N_14626);
xnor U21981 (N_21981,N_11475,N_16944);
and U21982 (N_21982,N_18400,N_19443);
nor U21983 (N_21983,N_11608,N_19005);
or U21984 (N_21984,N_14193,N_14787);
and U21985 (N_21985,N_11579,N_12907);
xor U21986 (N_21986,N_15771,N_12226);
xnor U21987 (N_21987,N_19108,N_10027);
or U21988 (N_21988,N_14729,N_10952);
xor U21989 (N_21989,N_16632,N_12471);
nand U21990 (N_21990,N_13630,N_17221);
nor U21991 (N_21991,N_19779,N_15554);
or U21992 (N_21992,N_16677,N_10290);
or U21993 (N_21993,N_11534,N_11089);
xor U21994 (N_21994,N_11520,N_15778);
or U21995 (N_21995,N_16003,N_11537);
nand U21996 (N_21996,N_10087,N_15267);
nor U21997 (N_21997,N_11331,N_19876);
nor U21998 (N_21998,N_11445,N_13530);
or U21999 (N_21999,N_10221,N_17713);
nand U22000 (N_22000,N_13246,N_16591);
or U22001 (N_22001,N_12299,N_19890);
nor U22002 (N_22002,N_10292,N_16726);
or U22003 (N_22003,N_13124,N_16713);
and U22004 (N_22004,N_18646,N_17396);
and U22005 (N_22005,N_17201,N_19067);
xor U22006 (N_22006,N_17670,N_17050);
and U22007 (N_22007,N_15565,N_16828);
xor U22008 (N_22008,N_11378,N_12258);
xor U22009 (N_22009,N_14503,N_15707);
nand U22010 (N_22010,N_12697,N_10981);
nand U22011 (N_22011,N_14210,N_12768);
and U22012 (N_22012,N_12674,N_14714);
or U22013 (N_22013,N_16146,N_10112);
nand U22014 (N_22014,N_17471,N_15003);
xnor U22015 (N_22015,N_17997,N_12813);
xnor U22016 (N_22016,N_17093,N_17755);
nor U22017 (N_22017,N_17261,N_14613);
xor U22018 (N_22018,N_16332,N_11514);
nand U22019 (N_22019,N_11389,N_11007);
xnor U22020 (N_22020,N_18485,N_17794);
xnor U22021 (N_22021,N_10206,N_15344);
or U22022 (N_22022,N_15718,N_15858);
nor U22023 (N_22023,N_18561,N_14571);
xor U22024 (N_22024,N_19491,N_15059);
xor U22025 (N_22025,N_19433,N_18894);
nand U22026 (N_22026,N_11706,N_14420);
nand U22027 (N_22027,N_11748,N_16300);
xor U22028 (N_22028,N_11040,N_18431);
and U22029 (N_22029,N_18789,N_14876);
nor U22030 (N_22030,N_14899,N_18075);
xor U22031 (N_22031,N_10392,N_13508);
and U22032 (N_22032,N_13140,N_15399);
and U22033 (N_22033,N_11626,N_12234);
xor U22034 (N_22034,N_17284,N_18515);
xor U22035 (N_22035,N_18251,N_16621);
nor U22036 (N_22036,N_10450,N_13380);
and U22037 (N_22037,N_14572,N_10533);
nand U22038 (N_22038,N_10171,N_14505);
nor U22039 (N_22039,N_19327,N_12070);
nor U22040 (N_22040,N_15023,N_13499);
or U22041 (N_22041,N_12140,N_17318);
nor U22042 (N_22042,N_10149,N_12906);
xnor U22043 (N_22043,N_13506,N_16134);
xor U22044 (N_22044,N_11227,N_15624);
nand U22045 (N_22045,N_17949,N_17334);
xor U22046 (N_22046,N_16976,N_18298);
nand U22047 (N_22047,N_13663,N_10419);
xnor U22048 (N_22048,N_18836,N_12061);
nor U22049 (N_22049,N_18575,N_12427);
or U22050 (N_22050,N_16660,N_19518);
nand U22051 (N_22051,N_14402,N_14543);
and U22052 (N_22052,N_11729,N_15256);
and U22053 (N_22053,N_16127,N_17038);
or U22054 (N_22054,N_16167,N_14205);
nor U22055 (N_22055,N_10444,N_19334);
nor U22056 (N_22056,N_12546,N_11775);
nand U22057 (N_22057,N_15803,N_11103);
nor U22058 (N_22058,N_14697,N_19082);
or U22059 (N_22059,N_15804,N_13016);
nor U22060 (N_22060,N_11428,N_14518);
and U22061 (N_22061,N_12021,N_11496);
or U22062 (N_22062,N_18823,N_19989);
and U22063 (N_22063,N_19300,N_13685);
nand U22064 (N_22064,N_12897,N_17283);
nor U22065 (N_22065,N_17115,N_13205);
and U22066 (N_22066,N_11662,N_16348);
or U22067 (N_22067,N_17416,N_19860);
or U22068 (N_22068,N_19283,N_16883);
nor U22069 (N_22069,N_15126,N_18136);
xnor U22070 (N_22070,N_19040,N_12896);
or U22071 (N_22071,N_16983,N_19207);
or U22072 (N_22072,N_11049,N_18260);
nor U22073 (N_22073,N_18966,N_19498);
xnor U22074 (N_22074,N_19538,N_10717);
and U22075 (N_22075,N_15454,N_16026);
or U22076 (N_22076,N_13567,N_16126);
and U22077 (N_22077,N_16555,N_16686);
nand U22078 (N_22078,N_18984,N_13476);
nand U22079 (N_22079,N_11876,N_13125);
nand U22080 (N_22080,N_16992,N_15780);
nor U22081 (N_22081,N_11030,N_12679);
and U22082 (N_22082,N_13931,N_16249);
nand U22083 (N_22083,N_12451,N_12144);
or U22084 (N_22084,N_16756,N_17497);
xnor U22085 (N_22085,N_12922,N_12438);
or U22086 (N_22086,N_19626,N_12772);
nor U22087 (N_22087,N_11502,N_17965);
and U22088 (N_22088,N_19574,N_13059);
xnor U22089 (N_22089,N_14523,N_10803);
or U22090 (N_22090,N_10320,N_13919);
xor U22091 (N_22091,N_19320,N_11511);
and U22092 (N_22092,N_17871,N_10111);
and U22093 (N_22093,N_10624,N_19516);
xnor U22094 (N_22094,N_12103,N_13591);
and U22095 (N_22095,N_10707,N_14687);
xor U22096 (N_22096,N_16793,N_15350);
nor U22097 (N_22097,N_16586,N_13376);
nand U22098 (N_22098,N_15849,N_16533);
nor U22099 (N_22099,N_13593,N_19822);
and U22100 (N_22100,N_10850,N_16023);
nand U22101 (N_22101,N_13806,N_16260);
nand U22102 (N_22102,N_13387,N_13815);
xor U22103 (N_22103,N_19211,N_19640);
nor U22104 (N_22104,N_13983,N_16303);
or U22105 (N_22105,N_15958,N_15295);
xnor U22106 (N_22106,N_17404,N_14222);
or U22107 (N_22107,N_17371,N_10387);
nor U22108 (N_22108,N_12257,N_10153);
nand U22109 (N_22109,N_15106,N_19199);
nand U22110 (N_22110,N_16362,N_17162);
xor U22111 (N_22111,N_14690,N_14886);
nand U22112 (N_22112,N_14485,N_14297);
and U22113 (N_22113,N_18770,N_18001);
nor U22114 (N_22114,N_10385,N_10266);
nor U22115 (N_22115,N_15450,N_11366);
and U22116 (N_22116,N_18841,N_11275);
xnor U22117 (N_22117,N_17616,N_14473);
and U22118 (N_22118,N_10538,N_14300);
xnor U22119 (N_22119,N_18949,N_15457);
xor U22120 (N_22120,N_18383,N_12267);
xor U22121 (N_22121,N_18103,N_14991);
or U22122 (N_22122,N_17792,N_14875);
nand U22123 (N_22123,N_14904,N_14383);
xnor U22124 (N_22124,N_11477,N_11942);
and U22125 (N_22125,N_12963,N_13168);
or U22126 (N_22126,N_18579,N_13348);
nand U22127 (N_22127,N_12875,N_10779);
or U22128 (N_22128,N_16157,N_15237);
or U22129 (N_22129,N_16244,N_11815);
nand U22130 (N_22130,N_10997,N_15753);
xor U22131 (N_22131,N_15118,N_11095);
or U22132 (N_22132,N_14720,N_15314);
xnor U22133 (N_22133,N_16512,N_17708);
and U22134 (N_22134,N_19371,N_19136);
nor U22135 (N_22135,N_10890,N_14091);
xnor U22136 (N_22136,N_14960,N_15826);
xnor U22137 (N_22137,N_14733,N_12425);
xor U22138 (N_22138,N_14609,N_14887);
and U22139 (N_22139,N_13878,N_18165);
nand U22140 (N_22140,N_14094,N_16092);
nand U22141 (N_22141,N_13618,N_11684);
xor U22142 (N_22142,N_13992,N_19059);
and U22143 (N_22143,N_17743,N_13692);
nor U22144 (N_22144,N_15408,N_14784);
nor U22145 (N_22145,N_14212,N_12623);
nor U22146 (N_22146,N_15070,N_19235);
nor U22147 (N_22147,N_19266,N_17640);
or U22148 (N_22148,N_16365,N_11018);
and U22149 (N_22149,N_15540,N_12303);
xor U22150 (N_22150,N_12970,N_10742);
xor U22151 (N_22151,N_10935,N_11480);
and U22152 (N_22152,N_15047,N_16105);
and U22153 (N_22153,N_14287,N_18088);
xnor U22154 (N_22154,N_13873,N_14718);
or U22155 (N_22155,N_11347,N_17621);
nor U22156 (N_22156,N_19210,N_15289);
nor U22157 (N_22157,N_15558,N_13410);
xnor U22158 (N_22158,N_10260,N_11215);
nand U22159 (N_22159,N_18467,N_16468);
nor U22160 (N_22160,N_13328,N_14504);
or U22161 (N_22161,N_16729,N_16925);
nor U22162 (N_22162,N_12573,N_16250);
nand U22163 (N_22163,N_11675,N_10478);
or U22164 (N_22164,N_15405,N_10643);
xnor U22165 (N_22165,N_12494,N_13551);
and U22166 (N_22166,N_18649,N_19526);
nor U22167 (N_22167,N_16785,N_11300);
nand U22168 (N_22168,N_13549,N_19936);
nor U22169 (N_22169,N_16012,N_19171);
nor U22170 (N_22170,N_13316,N_13227);
nand U22171 (N_22171,N_12435,N_18025);
xnor U22172 (N_22172,N_11724,N_16451);
and U22173 (N_22173,N_10078,N_12377);
nor U22174 (N_22174,N_14691,N_16181);
nor U22175 (N_22175,N_11761,N_15066);
nor U22176 (N_22176,N_15137,N_14755);
or U22177 (N_22177,N_15939,N_19315);
and U22178 (N_22178,N_16032,N_17336);
nand U22179 (N_22179,N_17712,N_13266);
xnor U22180 (N_22180,N_12126,N_13613);
nor U22181 (N_22181,N_12874,N_16419);
and U22182 (N_22182,N_10614,N_10734);
and U22183 (N_22183,N_15436,N_19766);
xor U22184 (N_22184,N_18313,N_15168);
nor U22185 (N_22185,N_19227,N_18363);
or U22186 (N_22186,N_11393,N_11337);
and U22187 (N_22187,N_10437,N_11468);
nand U22188 (N_22188,N_11408,N_14086);
xnor U22189 (N_22189,N_16600,N_13132);
nor U22190 (N_22190,N_17857,N_16664);
nor U22191 (N_22191,N_16350,N_15052);
xnor U22192 (N_22192,N_16314,N_19409);
xnor U22193 (N_22193,N_18504,N_18576);
nand U22194 (N_22194,N_10435,N_19771);
nor U22195 (N_22195,N_12116,N_16488);
and U22196 (N_22196,N_17365,N_11953);
nor U22197 (N_22197,N_13356,N_13503);
and U22198 (N_22198,N_15373,N_11784);
nand U22199 (N_22199,N_15092,N_16969);
nor U22200 (N_22200,N_19250,N_13114);
nor U22201 (N_22201,N_17438,N_15155);
xor U22202 (N_22202,N_16356,N_18864);
nand U22203 (N_22203,N_17410,N_17817);
and U22204 (N_22204,N_15805,N_19718);
and U22205 (N_22205,N_17345,N_15660);
nand U22206 (N_22206,N_18872,N_16406);
or U22207 (N_22207,N_10650,N_18886);
xnor U22208 (N_22208,N_10476,N_10309);
or U22209 (N_22209,N_16030,N_13520);
nand U22210 (N_22210,N_14036,N_11987);
and U22211 (N_22211,N_17141,N_10422);
and U22212 (N_22212,N_17434,N_13485);
nand U22213 (N_22213,N_11302,N_15463);
or U22214 (N_22214,N_10071,N_16343);
nand U22215 (N_22215,N_18529,N_10019);
and U22216 (N_22216,N_13390,N_11697);
nor U22217 (N_22217,N_12601,N_16792);
nor U22218 (N_22218,N_15863,N_18980);
nor U22219 (N_22219,N_18113,N_10464);
nand U22220 (N_22220,N_18820,N_10362);
xor U22221 (N_22221,N_18693,N_16408);
or U22222 (N_22222,N_12825,N_17363);
and U22223 (N_22223,N_10016,N_17636);
nor U22224 (N_22224,N_18718,N_10265);
and U22225 (N_22225,N_15549,N_16737);
xor U22226 (N_22226,N_14416,N_14879);
xnor U22227 (N_22227,N_16187,N_12434);
and U22228 (N_22228,N_12378,N_11172);
xor U22229 (N_22229,N_19145,N_19341);
nand U22230 (N_22230,N_14983,N_16579);
and U22231 (N_22231,N_18257,N_11990);
nand U22232 (N_22232,N_15026,N_16198);
or U22233 (N_22233,N_13049,N_16712);
xnor U22234 (N_22234,N_13673,N_14425);
or U22235 (N_22235,N_18843,N_17633);
nand U22236 (N_22236,N_19345,N_15928);
xnor U22237 (N_22237,N_19677,N_17556);
xor U22238 (N_22238,N_16539,N_15171);
or U22239 (N_22239,N_11016,N_12670);
or U22240 (N_22240,N_15892,N_19037);
or U22241 (N_22241,N_16856,N_15481);
nor U22242 (N_22242,N_13443,N_10995);
nor U22243 (N_22243,N_19331,N_13921);
and U22244 (N_22244,N_14762,N_16904);
and U22245 (N_22245,N_17617,N_19413);
xnor U22246 (N_22246,N_14536,N_10239);
or U22247 (N_22247,N_18365,N_10479);
nand U22248 (N_22248,N_17883,N_11984);
or U22249 (N_22249,N_16009,N_19476);
and U22250 (N_22250,N_15416,N_19296);
nand U22251 (N_22251,N_14592,N_10729);
or U22252 (N_22252,N_15914,N_11296);
and U22253 (N_22253,N_15215,N_13010);
or U22254 (N_22254,N_11883,N_19874);
nor U22255 (N_22255,N_14859,N_13210);
nor U22256 (N_22256,N_14329,N_10731);
nand U22257 (N_22257,N_12700,N_15044);
nand U22258 (N_22258,N_18340,N_11238);
or U22259 (N_22259,N_16398,N_16942);
nand U22260 (N_22260,N_10156,N_17836);
and U22261 (N_22261,N_14114,N_14506);
and U22262 (N_22262,N_18160,N_17136);
nand U22263 (N_22263,N_18466,N_13218);
or U22264 (N_22264,N_14630,N_18684);
nor U22265 (N_22265,N_18541,N_16174);
nor U22266 (N_22266,N_18601,N_13655);
nor U22267 (N_22267,N_12864,N_15205);
and U22268 (N_22268,N_19878,N_11658);
or U22269 (N_22269,N_11611,N_10996);
or U22270 (N_22270,N_16041,N_17098);
nand U22271 (N_22271,N_15060,N_19275);
xnor U22272 (N_22272,N_19071,N_16231);
nor U22273 (N_22273,N_14929,N_12324);
nor U22274 (N_22274,N_13737,N_13989);
nor U22275 (N_22275,N_16022,N_19840);
xnor U22276 (N_22276,N_10217,N_18447);
nand U22277 (N_22277,N_10023,N_19028);
nand U22278 (N_22278,N_19833,N_14230);
or U22279 (N_22279,N_18411,N_10814);
and U22280 (N_22280,N_14160,N_19790);
nor U22281 (N_22281,N_11365,N_18053);
xnor U22282 (N_22282,N_12954,N_14312);
nor U22283 (N_22283,N_19104,N_19204);
nand U22284 (N_22284,N_18885,N_18617);
or U22285 (N_22285,N_19631,N_18960);
nor U22286 (N_22286,N_14564,N_13802);
or U22287 (N_22287,N_12902,N_10504);
and U22288 (N_22288,N_16831,N_11114);
nand U22289 (N_22289,N_11307,N_17128);
nand U22290 (N_22290,N_13281,N_16516);
or U22291 (N_22291,N_18132,N_10126);
nor U22292 (N_22292,N_16043,N_15885);
and U22293 (N_22293,N_17541,N_11194);
xor U22294 (N_22294,N_17972,N_15880);
nor U22295 (N_22295,N_18076,N_11193);
nor U22296 (N_22296,N_10937,N_13937);
or U22297 (N_22297,N_10400,N_10433);
nor U22298 (N_22298,N_14873,N_18016);
or U22299 (N_22299,N_18024,N_13822);
nand U22300 (N_22300,N_17779,N_13955);
xnor U22301 (N_22301,N_19788,N_14822);
nor U22302 (N_22302,N_14391,N_17939);
or U22303 (N_22303,N_16329,N_14969);
and U22304 (N_22304,N_19206,N_16446);
xnor U22305 (N_22305,N_15956,N_12613);
and U22306 (N_22306,N_13906,N_13449);
xnor U22307 (N_22307,N_15058,N_12574);
nor U22308 (N_22308,N_12216,N_14713);
nor U22309 (N_22309,N_16143,N_18098);
and U22310 (N_22310,N_18488,N_13312);
nor U22311 (N_22311,N_13674,N_16253);
nor U22312 (N_22312,N_15452,N_11310);
xnor U22313 (N_22313,N_18448,N_10637);
nand U22314 (N_22314,N_18115,N_16770);
and U22315 (N_22315,N_11805,N_11558);
nand U22316 (N_22316,N_14013,N_13286);
or U22317 (N_22317,N_10672,N_16494);
and U22318 (N_22318,N_16596,N_18990);
or U22319 (N_22319,N_10047,N_17144);
and U22320 (N_22320,N_17539,N_18403);
or U22321 (N_22321,N_18907,N_18074);
xnor U22322 (N_22322,N_18830,N_15990);
nand U22323 (N_22323,N_16431,N_15628);
nand U22324 (N_22324,N_12733,N_13067);
nor U22325 (N_22325,N_10519,N_16762);
xnor U22326 (N_22326,N_10361,N_15388);
or U22327 (N_22327,N_16672,N_15652);
and U22328 (N_22328,N_18554,N_12797);
xor U22329 (N_22329,N_11635,N_12987);
nor U22330 (N_22330,N_19760,N_12452);
xnor U22331 (N_22331,N_14986,N_17262);
xor U22332 (N_22332,N_11047,N_15499);
and U22333 (N_22333,N_15479,N_13935);
nor U22334 (N_22334,N_14089,N_19316);
nor U22335 (N_22335,N_16267,N_17514);
and U22336 (N_22336,N_19368,N_18045);
or U22337 (N_22337,N_11495,N_10326);
xor U22338 (N_22338,N_18976,N_11659);
and U22339 (N_22339,N_12737,N_15606);
nand U22340 (N_22340,N_19589,N_19641);
or U22341 (N_22341,N_18225,N_12505);
or U22342 (N_22342,N_12986,N_10936);
xnor U22343 (N_22343,N_19637,N_17947);
xor U22344 (N_22344,N_10879,N_16571);
and U22345 (N_22345,N_18889,N_16060);
or U22346 (N_22346,N_19416,N_11896);
nand U22347 (N_22347,N_12871,N_13236);
and U22348 (N_22348,N_18834,N_12069);
nand U22349 (N_22349,N_16443,N_19584);
xor U22350 (N_22350,N_17091,N_19755);
and U22351 (N_22351,N_10836,N_18667);
nand U22352 (N_22352,N_10509,N_13845);
or U22353 (N_22353,N_14849,N_17856);
nand U22354 (N_22354,N_14851,N_17263);
xor U22355 (N_22355,N_16478,N_14195);
nand U22356 (N_22356,N_13100,N_13850);
xnor U22357 (N_22357,N_19215,N_19474);
or U22358 (N_22358,N_18179,N_13950);
xnor U22359 (N_22359,N_13386,N_18342);
or U22360 (N_22360,N_10214,N_11919);
and U22361 (N_22361,N_12430,N_10110);
xor U22362 (N_22362,N_19399,N_14257);
nand U22363 (N_22363,N_11400,N_10709);
and U22364 (N_22364,N_10055,N_11878);
or U22365 (N_22365,N_17904,N_19352);
or U22366 (N_22366,N_14692,N_17907);
xor U22367 (N_22367,N_10229,N_19741);
and U22368 (N_22368,N_11373,N_10531);
xnor U22369 (N_22369,N_17489,N_18567);
or U22370 (N_22370,N_10639,N_11036);
nand U22371 (N_22371,N_16135,N_12240);
or U22372 (N_22372,N_13260,N_14858);
and U22373 (N_22373,N_12220,N_18333);
or U22374 (N_22374,N_16321,N_10001);
xor U22375 (N_22375,N_10681,N_19854);
and U22376 (N_22376,N_12235,N_14240);
xnor U22377 (N_22377,N_15596,N_17648);
and U22378 (N_22378,N_19617,N_16679);
nor U22379 (N_22379,N_16279,N_16137);
or U22380 (N_22380,N_11148,N_18969);
and U22381 (N_22381,N_15889,N_16982);
nand U22382 (N_22382,N_18346,N_17920);
or U22383 (N_22383,N_13150,N_10529);
nand U22384 (N_22384,N_19284,N_14628);
nor U22385 (N_22385,N_15538,N_11497);
nor U22386 (N_22386,N_13224,N_10950);
and U22387 (N_22387,N_12320,N_10311);
xor U22388 (N_22388,N_14994,N_16508);
or U22389 (N_22389,N_12413,N_14669);
xor U22390 (N_22390,N_11043,N_15490);
and U22391 (N_22391,N_10162,N_19231);
xnor U22392 (N_22392,N_11532,N_18948);
and U22393 (N_22393,N_17890,N_13052);
xor U22394 (N_22394,N_10226,N_14666);
nand U22395 (N_22395,N_15975,N_11717);
or U22396 (N_22396,N_14184,N_11971);
and U22397 (N_22397,N_10768,N_12148);
nor U22398 (N_22398,N_10223,N_13178);
nand U22399 (N_22399,N_15125,N_11988);
nor U22400 (N_22400,N_10228,N_12551);
and U22401 (N_22401,N_16056,N_16101);
xnor U22402 (N_22402,N_19095,N_15829);
xnor U22403 (N_22403,N_11226,N_13292);
nand U22404 (N_22404,N_13576,N_14576);
nand U22405 (N_22405,N_10623,N_18611);
xor U22406 (N_22406,N_11162,N_16825);
or U22407 (N_22407,N_10634,N_12031);
or U22408 (N_22408,N_19537,N_14148);
xnor U22409 (N_22409,N_14681,N_18543);
nor U22410 (N_22410,N_14495,N_13971);
and U22411 (N_22411,N_11175,N_11474);
nand U22412 (N_22412,N_15472,N_14863);
or U22413 (N_22413,N_18727,N_10884);
nor U22414 (N_22414,N_17395,N_13368);
nor U22415 (N_22415,N_18483,N_14285);
nor U22416 (N_22416,N_10872,N_16839);
nand U22417 (N_22417,N_19020,N_14458);
nand U22418 (N_22418,N_12497,N_10494);
xor U22419 (N_22419,N_10488,N_13927);
xor U22420 (N_22420,N_11313,N_12263);
and U22421 (N_22421,N_11702,N_14709);
nor U22422 (N_22422,N_18380,N_18897);
xor U22423 (N_22423,N_13448,N_14378);
nor U22424 (N_22424,N_16430,N_15949);
nand U22425 (N_22425,N_15453,N_13608);
and U22426 (N_22426,N_15329,N_10011);
nand U22427 (N_22427,N_19439,N_12730);
nand U22428 (N_22428,N_18596,N_15245);
xnor U22429 (N_22429,N_13128,N_19685);
and U22430 (N_22430,N_14645,N_11084);
and U22431 (N_22431,N_16286,N_16690);
nor U22432 (N_22432,N_16269,N_13532);
and U22433 (N_22433,N_19079,N_17164);
xor U22434 (N_22434,N_14005,N_16994);
nand U22435 (N_22435,N_13884,N_12889);
xor U22436 (N_22436,N_13439,N_14809);
nand U22437 (N_22437,N_18893,N_10381);
or U22438 (N_22438,N_18961,N_17084);
and U22439 (N_22439,N_12455,N_13209);
nor U22440 (N_22440,N_15073,N_15375);
nand U22441 (N_22441,N_11250,N_10406);
nor U22442 (N_22442,N_19252,N_14806);
and U22443 (N_22443,N_12090,N_11866);
and U22444 (N_22444,N_19643,N_19132);
and U22445 (N_22445,N_18699,N_18178);
xnor U22446 (N_22446,N_12992,N_11323);
nor U22447 (N_22447,N_14293,N_16248);
or U22448 (N_22448,N_10679,N_13700);
xnor U22449 (N_22449,N_19573,N_12698);
or U22450 (N_22450,N_13299,N_13690);
nand U22451 (N_22451,N_13773,N_18954);
or U22452 (N_22452,N_15824,N_16750);
xnor U22453 (N_22453,N_10878,N_16725);
or U22454 (N_22454,N_17752,N_18743);
or U22455 (N_22455,N_15663,N_14792);
or U22456 (N_22456,N_17294,N_17776);
or U22457 (N_22457,N_15566,N_19824);
nor U22458 (N_22458,N_10905,N_10079);
xnor U22459 (N_22459,N_15714,N_19999);
nor U22460 (N_22460,N_13219,N_10733);
and U22461 (N_22461,N_17739,N_13665);
nand U22462 (N_22462,N_14211,N_10548);
xnor U22463 (N_22463,N_15728,N_13888);
and U22464 (N_22464,N_10924,N_16422);
and U22465 (N_22465,N_18526,N_16218);
and U22466 (N_22466,N_11796,N_13001);
xnor U22467 (N_22467,N_19613,N_17967);
and U22468 (N_22468,N_13022,N_11957);
or U22469 (N_22469,N_17946,N_12592);
nor U22470 (N_22470,N_19780,N_15522);
and U22471 (N_22471,N_16723,N_19930);
or U22472 (N_22472,N_18776,N_11206);
or U22473 (N_22473,N_14500,N_17316);
xnor U22474 (N_22474,N_14019,N_13211);
xnor U22475 (N_22475,N_16265,N_15226);
xor U22476 (N_22476,N_15548,N_11721);
nor U22477 (N_22477,N_17915,N_12629);
or U22478 (N_22478,N_11714,N_15122);
nor U22479 (N_22479,N_10427,N_11010);
nor U22480 (N_22480,N_12187,N_11978);
or U22481 (N_22481,N_18440,N_12388);
and U22482 (N_22482,N_18513,N_12839);
xnor U22483 (N_22483,N_13581,N_14694);
or U22484 (N_22484,N_14680,N_18436);
or U22485 (N_22485,N_17843,N_12119);
or U22486 (N_22486,N_12632,N_19629);
nor U22487 (N_22487,N_19344,N_13319);
or U22488 (N_22488,N_11107,N_12034);
and U22489 (N_22489,N_16216,N_10065);
nand U22490 (N_22490,N_16546,N_14204);
nand U22491 (N_22491,N_12584,N_13789);
nor U22492 (N_22492,N_10164,N_18394);
or U22493 (N_22493,N_17133,N_15798);
and U22494 (N_22494,N_12146,N_15145);
nand U22495 (N_22495,N_19623,N_15217);
xnor U22496 (N_22496,N_12368,N_15801);
nor U22497 (N_22497,N_10776,N_14795);
nor U22498 (N_22498,N_12080,N_16721);
nor U22499 (N_22499,N_12609,N_10486);
and U22500 (N_22500,N_19582,N_15909);
nor U22501 (N_22501,N_12448,N_15926);
or U22502 (N_22502,N_11646,N_14653);
nor U22503 (N_22503,N_19116,N_10499);
xor U22504 (N_22504,N_14579,N_11252);
and U22505 (N_22505,N_11541,N_18802);
nand U22506 (N_22506,N_14514,N_19561);
nand U22507 (N_22507,N_17429,N_18719);
xnor U22508 (N_22508,N_12310,N_13750);
nand U22509 (N_22509,N_10770,N_11074);
nor U22510 (N_22510,N_14176,N_16159);
nand U22511 (N_22511,N_12721,N_16261);
nor U22512 (N_22512,N_15737,N_14794);
or U22513 (N_22513,N_18345,N_18164);
xor U22514 (N_22514,N_17014,N_14248);
nand U22515 (N_22515,N_18873,N_16500);
or U22516 (N_22516,N_15077,N_19940);
nand U22517 (N_22517,N_10304,N_16011);
xor U22518 (N_22518,N_10665,N_14456);
xor U22519 (N_22519,N_19158,N_10786);
or U22520 (N_22520,N_18863,N_12780);
xnor U22521 (N_22521,N_10941,N_15559);
nor U22522 (N_22522,N_11100,N_16755);
nor U22523 (N_22523,N_15611,N_11281);
xor U22524 (N_22524,N_18510,N_16067);
xnor U22525 (N_22525,N_17630,N_16457);
or U22526 (N_22526,N_10986,N_18570);
or U22527 (N_22527,N_13002,N_11387);
xor U22528 (N_22528,N_19748,N_14108);
nor U22529 (N_22529,N_12598,N_13908);
nand U22530 (N_22530,N_11414,N_12999);
or U22531 (N_22531,N_11569,N_18465);
xnor U22532 (N_22532,N_12104,N_10632);
nand U22533 (N_22533,N_14757,N_15035);
nor U22534 (N_22534,N_10298,N_18204);
and U22535 (N_22535,N_19835,N_13428);
and U22536 (N_22536,N_14365,N_12444);
and U22537 (N_22537,N_12659,N_11177);
nor U22538 (N_22538,N_10701,N_10723);
or U22539 (N_22539,N_12946,N_13474);
nand U22540 (N_22540,N_14159,N_19621);
nor U22541 (N_22541,N_18428,N_19249);
nand U22542 (N_22542,N_14728,N_17064);
nor U22543 (N_22543,N_12000,N_16973);
and U22544 (N_22544,N_15498,N_11217);
nand U22545 (N_22545,N_16085,N_13426);
nand U22546 (N_22546,N_18630,N_11842);
or U22547 (N_22547,N_15625,N_13177);
nand U22548 (N_22548,N_14120,N_11965);
and U22549 (N_22549,N_13879,N_14517);
and U22550 (N_22550,N_11678,N_16536);
nand U22551 (N_22551,N_10965,N_15872);
nand U22552 (N_22552,N_15862,N_12788);
nand U22553 (N_22553,N_16489,N_10972);
or U22554 (N_22554,N_11158,N_16745);
nand U22555 (N_22555,N_14475,N_11506);
nand U22556 (N_22556,N_10881,N_16753);
nand U22557 (N_22557,N_16189,N_11720);
nand U22558 (N_22558,N_19724,N_10551);
nand U22559 (N_22559,N_15524,N_16978);
and U22560 (N_22560,N_12511,N_10676);
nor U22561 (N_22561,N_10061,N_18673);
nand U22562 (N_22562,N_19054,N_16324);
xor U22563 (N_22563,N_16673,N_15495);
xnor U22564 (N_22564,N_16389,N_19412);
or U22565 (N_22565,N_11418,N_10287);
xor U22566 (N_22566,N_18856,N_18595);
xor U22567 (N_22567,N_13013,N_11240);
nand U22568 (N_22568,N_15216,N_11844);
nand U22569 (N_22569,N_11752,N_16692);
and U22570 (N_22570,N_19969,N_17236);
and U22571 (N_22571,N_16007,N_12582);
xnor U22572 (N_22572,N_13552,N_17213);
nand U22573 (N_22573,N_19372,N_19218);
nor U22574 (N_22574,N_10798,N_13521);
or U22575 (N_22575,N_14143,N_19396);
nor U22576 (N_22576,N_13347,N_14911);
nand U22577 (N_22577,N_16887,N_11833);
or U22578 (N_22578,N_19290,N_19884);
xnor U22579 (N_22579,N_15275,N_10834);
nand U22580 (N_22580,N_15306,N_15407);
nand U22581 (N_22581,N_11218,N_11106);
nand U22582 (N_22582,N_11004,N_17317);
and U22583 (N_22583,N_18692,N_11123);
or U22584 (N_22584,N_10921,N_18774);
or U22585 (N_22585,N_13798,N_11771);
or U22586 (N_22586,N_18878,N_18047);
and U22587 (N_22587,N_11271,N_18588);
and U22588 (N_22588,N_17526,N_19025);
nor U22589 (N_22589,N_13043,N_14241);
nand U22590 (N_22590,N_16884,N_16981);
nor U22591 (N_22591,N_19261,N_11598);
xnor U22592 (N_22592,N_16724,N_15268);
nor U22593 (N_22593,N_17510,N_14636);
nor U22594 (N_22594,N_17026,N_15018);
or U22595 (N_22595,N_15904,N_12975);
xor U22596 (N_22596,N_19286,N_19812);
or U22597 (N_22597,N_17407,N_13413);
nor U22598 (N_22598,N_12221,N_19297);
nand U22599 (N_22599,N_19225,N_11948);
or U22600 (N_22600,N_11882,N_14861);
nand U22601 (N_22601,N_12312,N_16710);
nor U22602 (N_22602,N_11581,N_12167);
xor U22603 (N_22603,N_18114,N_13047);
xor U22604 (N_22604,N_12746,N_10675);
xnor U22605 (N_22605,N_16414,N_11200);
nand U22606 (N_22606,N_15427,N_17194);
or U22607 (N_22607,N_14273,N_17424);
nor U22608 (N_22608,N_14045,N_13196);
xnor U22609 (N_22609,N_17187,N_11187);
nor U22610 (N_22610,N_12599,N_13460);
and U22611 (N_22611,N_12050,N_12964);
nand U22612 (N_22612,N_13057,N_14693);
or U22613 (N_22613,N_19139,N_14177);
nand U22614 (N_22614,N_13871,N_12238);
or U22615 (N_22615,N_17191,N_11517);
and U22616 (N_22616,N_14268,N_19349);
or U22617 (N_22617,N_18523,N_14556);
or U22618 (N_22618,N_15353,N_17575);
and U22619 (N_22619,N_13405,N_16561);
xor U22620 (N_22620,N_19565,N_14638);
xor U22621 (N_22621,N_17040,N_14137);
nand U22622 (N_22622,N_10511,N_14649);
xnor U22623 (N_22623,N_15834,N_10702);
or U22624 (N_22624,N_19928,N_15266);
or U22625 (N_22625,N_11233,N_19263);
nand U22626 (N_22626,N_10530,N_19575);
or U22627 (N_22627,N_19728,N_19887);
or U22628 (N_22628,N_15037,N_16846);
or U22629 (N_22629,N_11476,N_12807);
xor U22630 (N_22630,N_12638,N_17651);
or U22631 (N_22631,N_13491,N_14793);
or U22632 (N_22632,N_17620,N_12489);
nor U22633 (N_22633,N_16768,N_11601);
nand U22634 (N_22634,N_15031,N_12428);
nor U22635 (N_22635,N_16495,N_14678);
or U22636 (N_22636,N_19872,N_18923);
nand U22637 (N_22637,N_18971,N_10368);
xor U22638 (N_22638,N_10227,N_10720);
or U22639 (N_22639,N_16386,N_12059);
nor U22640 (N_22640,N_11317,N_19277);
and U22641 (N_22641,N_10017,N_17500);
xor U22642 (N_22642,N_16186,N_11482);
xnor U22643 (N_22643,N_13051,N_17841);
nor U22644 (N_22644,N_12677,N_10917);
nor U22645 (N_22645,N_17370,N_14583);
nor U22646 (N_22646,N_16977,N_15683);
xnor U22647 (N_22647,N_10658,N_18427);
or U22648 (N_22648,N_18891,N_13623);
and U22649 (N_22649,N_10868,N_19313);
and U22650 (N_22650,N_11062,N_19614);
nand U22651 (N_22651,N_13991,N_17522);
nand U22652 (N_22652,N_16001,N_13775);
xor U22653 (N_22653,N_12483,N_16703);
nand U22654 (N_22654,N_10572,N_11501);
xnor U22655 (N_22655,N_13248,N_19373);
or U22656 (N_22656,N_14228,N_18520);
nor U22657 (N_22657,N_18338,N_16866);
or U22658 (N_22658,N_10130,N_18034);
and U22659 (N_22659,N_16469,N_12625);
xnor U22660 (N_22660,N_18505,N_14841);
and U22661 (N_22661,N_10859,N_18308);
and U22662 (N_22662,N_10403,N_19011);
xor U22663 (N_22663,N_15690,N_13037);
xnor U22664 (N_22664,N_18143,N_12777);
nor U22665 (N_22665,N_11332,N_10920);
nand U22666 (N_22666,N_17030,N_14975);
xor U22667 (N_22667,N_19176,N_15740);
and U22668 (N_22668,N_14415,N_15042);
and U22669 (N_22669,N_18535,N_15792);
nor U22670 (N_22670,N_15208,N_10411);
or U22671 (N_22671,N_19365,N_15053);
nand U22672 (N_22672,N_10724,N_13157);
xor U22673 (N_22673,N_12765,N_16604);
or U22674 (N_22674,N_11916,N_16031);
xnor U22675 (N_22675,N_19952,N_18932);
or U22676 (N_22676,N_16184,N_16292);
nand U22677 (N_22677,N_12002,N_18704);
xor U22678 (N_22678,N_14259,N_11354);
xor U22679 (N_22679,N_13334,N_15749);
or U22680 (N_22680,N_15644,N_17705);
nor U22681 (N_22681,N_13797,N_18399);
and U22682 (N_22682,N_15016,N_17572);
nand U22683 (N_22683,N_15932,N_17697);
nand U22684 (N_22684,N_14908,N_16366);
and U22685 (N_22685,N_13957,N_18358);
or U22686 (N_22686,N_17957,N_10696);
and U22687 (N_22687,N_19034,N_14030);
nand U22688 (N_22688,N_17561,N_14397);
and U22689 (N_22689,N_10858,N_11845);
and U22690 (N_22690,N_11818,N_13963);
nand U22691 (N_22691,N_17034,N_18146);
or U22692 (N_22692,N_18039,N_17901);
nor U22693 (N_22693,N_12527,N_15931);
nand U22694 (N_22694,N_13805,N_19941);
xor U22695 (N_22695,N_10980,N_10339);
and U22696 (N_22696,N_17139,N_16534);
and U22697 (N_22697,N_16241,N_11101);
and U22698 (N_22698,N_14953,N_16298);
xor U22699 (N_22699,N_17055,N_19953);
and U22700 (N_22700,N_12136,N_12169);
xnor U22701 (N_22701,N_16741,N_11032);
nand U22702 (N_22702,N_11283,N_13216);
or U22703 (N_22703,N_13367,N_16986);
nand U22704 (N_22704,N_19426,N_18933);
or U22705 (N_22705,N_14173,N_16327);
or U22706 (N_22706,N_13510,N_15349);
or U22707 (N_22707,N_15656,N_18459);
xor U22708 (N_22708,N_15572,N_11066);
nor U22709 (N_22709,N_15194,N_18668);
and U22710 (N_22710,N_14765,N_18188);
and U22711 (N_22711,N_12183,N_12890);
or U22712 (N_22712,N_13017,N_17376);
xor U22713 (N_22713,N_17104,N_13362);
or U22714 (N_22714,N_11912,N_19980);
and U22715 (N_22715,N_19834,N_19319);
or U22716 (N_22716,N_18171,N_14452);
and U22717 (N_22717,N_18311,N_15781);
nor U22718 (N_22718,N_18170,N_14819);
xor U22719 (N_22719,N_12815,N_18833);
and U22720 (N_22720,N_14698,N_15014);
or U22721 (N_22721,N_16193,N_18647);
nor U22722 (N_22722,N_17696,N_16290);
xor U22723 (N_22723,N_10943,N_16229);
xor U22724 (N_22724,N_14382,N_17570);
or U22725 (N_22725,N_19909,N_18220);
xor U22726 (N_22726,N_11143,N_15678);
nor U22727 (N_22727,N_18516,N_18013);
and U22728 (N_22728,N_19168,N_18352);
xor U22729 (N_22729,N_19531,N_18975);
or U22730 (N_22730,N_11666,N_16382);
xnor U22731 (N_22731,N_11308,N_18559);
xnor U22732 (N_22732,N_11884,N_16538);
nand U22733 (N_22733,N_14451,N_10108);
nand U22734 (N_22734,N_10968,N_19543);
xnor U22735 (N_22735,N_15934,N_15351);
nor U22736 (N_22736,N_14403,N_17802);
xnor U22737 (N_22737,N_12289,N_11638);
or U22738 (N_22738,N_14944,N_19411);
nand U22739 (N_22739,N_17120,N_12615);
nand U22740 (N_22740,N_17689,N_16281);
or U22741 (N_22741,N_12319,N_18414);
nor U22742 (N_22742,N_17900,N_10189);
nand U22743 (N_22743,N_14530,N_12453);
xnor U22744 (N_22744,N_13603,N_12079);
nor U22745 (N_22745,N_10609,N_10983);
nor U22746 (N_22746,N_14024,N_15777);
and U22747 (N_22747,N_13518,N_15590);
nand U22748 (N_22748,N_18545,N_11633);
or U22749 (N_22749,N_13739,N_10482);
and U22750 (N_22750,N_14047,N_10802);
xor U22751 (N_22751,N_18887,N_15650);
nand U22752 (N_22752,N_10497,N_17373);
nand U22753 (N_22753,N_15209,N_18690);
or U22754 (N_22754,N_11137,N_14595);
or U22755 (N_22755,N_10680,N_19254);
or U22756 (N_22756,N_18177,N_10553);
or U22757 (N_22757,N_12200,N_18326);
nand U22758 (N_22758,N_10317,N_13572);
or U22759 (N_22759,N_14347,N_12952);
nand U22760 (N_22760,N_10254,N_17118);
nor U22761 (N_22761,N_17944,N_14764);
or U22762 (N_22762,N_17403,N_14389);
nand U22763 (N_22763,N_19560,N_19201);
nor U22764 (N_22764,N_13416,N_14964);
and U22765 (N_22765,N_10867,N_11276);
and U22766 (N_22766,N_10425,N_12838);
nand U22767 (N_22767,N_18564,N_11375);
or U22768 (N_22768,N_13061,N_15195);
or U22769 (N_22769,N_14945,N_19731);
nor U22770 (N_22770,N_13585,N_15496);
xnor U22771 (N_22771,N_17254,N_16754);
or U22772 (N_22772,N_15083,N_17906);
and U22773 (N_22773,N_17804,N_19394);
nand U22774 (N_22774,N_19853,N_18375);
nor U22775 (N_22775,N_12657,N_14783);
nand U22776 (N_22776,N_15647,N_11657);
and U22777 (N_22777,N_16779,N_16926);
nand U22778 (N_22778,N_13425,N_16647);
and U22779 (N_22779,N_19155,N_19505);
nor U22780 (N_22780,N_14280,N_13473);
and U22781 (N_22781,N_12895,N_17227);
and U22782 (N_22782,N_19796,N_14464);
and U22783 (N_22783,N_14884,N_10365);
nand U22784 (N_22784,N_10823,N_10271);
nand U22785 (N_22785,N_12010,N_12593);
nand U22786 (N_22786,N_12512,N_17245);
and U22787 (N_22787,N_15846,N_15356);
and U22788 (N_22788,N_14188,N_17688);
and U22789 (N_22789,N_16307,N_15767);
xnor U22790 (N_22790,N_18622,N_16449);
xor U22791 (N_22791,N_11727,N_16564);
nor U22792 (N_22792,N_11484,N_11505);
nor U22793 (N_22793,N_14073,N_15414);
xnor U22794 (N_22794,N_14951,N_16900);
and U22795 (N_22795,N_10181,N_19836);
nor U22796 (N_22796,N_10932,N_16818);
xnor U22797 (N_22797,N_10738,N_10105);
nand U22798 (N_22798,N_11756,N_12459);
xor U22799 (N_22799,N_14123,N_17993);
nand U22800 (N_22800,N_12751,N_19793);
xor U22801 (N_22801,N_17959,N_19639);
nand U22802 (N_22802,N_16781,N_10765);
nand U22803 (N_22803,N_11587,N_17061);
or U22804 (N_22804,N_11795,N_12841);
and U22805 (N_22805,N_19599,N_12305);
nand U22806 (N_22806,N_15286,N_14040);
or U22807 (N_22807,N_18014,N_18987);
nand U22808 (N_22808,N_13036,N_11548);
and U22809 (N_22809,N_19906,N_10746);
nand U22810 (N_22810,N_14699,N_10979);
xor U22811 (N_22811,N_14977,N_13843);
nor U22812 (N_22812,N_18253,N_19558);
or U22813 (N_22813,N_18739,N_14940);
or U22814 (N_22814,N_11559,N_18745);
nor U22815 (N_22815,N_18438,N_17360);
or U22816 (N_22816,N_14938,N_12794);
nor U22817 (N_22817,N_10178,N_11108);
xnor U22818 (N_22818,N_18955,N_19883);
or U22819 (N_22819,N_16355,N_10719);
nand U22820 (N_22820,N_15010,N_15486);
xor U22821 (N_22821,N_18226,N_15523);
nor U22822 (N_22822,N_10851,N_14843);
nand U22823 (N_22823,N_12608,N_16054);
nor U22824 (N_22824,N_15528,N_15890);
nor U22825 (N_22825,N_14482,N_10251);
nand U22826 (N_22826,N_10716,N_14601);
nor U22827 (N_22827,N_19694,N_19507);
and U22828 (N_22828,N_13384,N_15174);
xnor U22829 (N_22829,N_16575,N_15845);
nor U22830 (N_22830,N_14569,N_14641);
and U22831 (N_22831,N_10656,N_10662);
xnor U22832 (N_22832,N_19475,N_10405);
xnor U22833 (N_22833,N_12202,N_16100);
or U22834 (N_22834,N_15432,N_12868);
nor U22835 (N_22835,N_14134,N_10985);
and U22836 (N_22836,N_13973,N_19043);
xnor U22837 (N_22837,N_17112,N_18494);
nor U22838 (N_22838,N_10472,N_13469);
nand U22839 (N_22839,N_19633,N_19078);
nor U22840 (N_22840,N_18740,N_13342);
xnor U22841 (N_22841,N_19129,N_14616);
nand U22842 (N_22842,N_16277,N_10974);
nor U22843 (N_22843,N_18270,N_19758);
and U22844 (N_22844,N_19489,N_12472);
xnor U22845 (N_22845,N_16511,N_12383);
xor U22846 (N_22846,N_15218,N_10436);
or U22847 (N_22847,N_11102,N_17197);
nor U22848 (N_22848,N_15397,N_19977);
nand U22849 (N_22849,N_10185,N_16251);
xor U22850 (N_22850,N_11179,N_17146);
xor U22851 (N_22851,N_17757,N_11212);
and U22852 (N_22852,N_17233,N_16938);
and U22853 (N_22853,N_16749,N_12501);
nand U22854 (N_22854,N_15588,N_15629);
xnor U22855 (N_22855,N_15115,N_16951);
xor U22856 (N_22856,N_17105,N_14758);
or U22857 (N_22857,N_19042,N_14541);
and U22858 (N_22858,N_19279,N_19089);
xnor U22859 (N_22859,N_13137,N_13558);
and U22860 (N_22860,N_18048,N_13943);
nand U22861 (N_22861,N_10369,N_12139);
nand U22862 (N_22862,N_11486,N_10869);
xor U22863 (N_22863,N_16058,N_11660);
or U22864 (N_22864,N_13969,N_11643);
nor U22865 (N_22865,N_15899,N_14921);
xor U22866 (N_22866,N_19451,N_12806);
nand U22867 (N_22867,N_17282,N_13335);
or U22868 (N_22868,N_15621,N_15882);
and U22869 (N_22869,N_14276,N_18183);
xor U22870 (N_22870,N_14065,N_17913);
nor U22871 (N_22871,N_12055,N_19787);
nand U22872 (N_22872,N_13946,N_17580);
nor U22873 (N_22873,N_18461,N_18023);
xnor U22874 (N_22874,N_12094,N_17722);
nor U22875 (N_22875,N_13892,N_11607);
nand U22876 (N_22876,N_15136,N_14594);
and U22877 (N_22877,N_19973,N_12015);
nand U22878 (N_22878,N_11969,N_16961);
xor U22879 (N_22879,N_18218,N_11783);
nor U22880 (N_22880,N_18775,N_18959);
and U22881 (N_22881,N_19226,N_16194);
nand U22882 (N_22882,N_17272,N_14370);
nand U22883 (N_22883,N_12648,N_12005);
nand U22884 (N_22884,N_17044,N_11413);
xnor U22885 (N_22885,N_18095,N_13111);
xnor U22886 (N_22886,N_16311,N_11136);
nor U22887 (N_22887,N_16682,N_16412);
nor U22888 (N_22888,N_11181,N_11865);
or U22889 (N_22889,N_18423,N_10754);
nand U22890 (N_22890,N_14778,N_17220);
xnor U22891 (N_22891,N_17731,N_15768);
or U22892 (N_22892,N_10267,N_13831);
xnor U22893 (N_22893,N_14597,N_17922);
and U22894 (N_22894,N_19912,N_18663);
nand U22895 (N_22895,N_14848,N_16224);
nor U22896 (N_22896,N_13273,N_13483);
and U22897 (N_22897,N_19064,N_11671);
xnor U22898 (N_22898,N_18434,N_19744);
nor U22899 (N_22899,N_15471,N_16807);
and U22900 (N_22900,N_11459,N_16502);
and U22901 (N_22901,N_16880,N_10767);
xor U22902 (N_22902,N_18599,N_10207);
nand U22903 (N_22903,N_18202,N_10253);
xnor U22904 (N_22904,N_17717,N_10280);
and U22905 (N_22905,N_10434,N_15584);
xnor U22906 (N_22906,N_12073,N_12691);
xor U22907 (N_22907,N_12616,N_19326);
or U22908 (N_22908,N_19479,N_15859);
xor U22909 (N_22909,N_19915,N_17614);
or U22910 (N_22910,N_10000,N_16162);
and U22911 (N_22911,N_13412,N_12380);
or U22912 (N_22912,N_17390,N_15985);
nand U22913 (N_22913,N_10694,N_19041);
or U22914 (N_22914,N_14479,N_12835);
nor U22915 (N_22915,N_18157,N_11029);
nand U22916 (N_22916,N_10246,N_12759);
and U22917 (N_22917,N_17006,N_18735);
or U22918 (N_22918,N_13728,N_17307);
and U22919 (N_22919,N_16746,N_12424);
nor U22920 (N_22920,N_16454,N_12385);
nor U22921 (N_22921,N_18334,N_17923);
xnor U22922 (N_22922,N_16623,N_10043);
and U22923 (N_22923,N_10831,N_13703);
and U22924 (N_22924,N_17019,N_13233);
and U22925 (N_22925,N_18246,N_12480);
nor U22926 (N_22926,N_17242,N_16076);
nand U22927 (N_22927,N_19850,N_14842);
xor U22928 (N_22928,N_19002,N_14135);
xnor U22929 (N_22929,N_17586,N_13920);
or U22930 (N_22930,N_16615,N_18941);
xnor U22931 (N_22931,N_17167,N_10915);
or U22932 (N_22932,N_16102,N_16121);
xor U22933 (N_22933,N_17559,N_19012);
nor U22934 (N_22934,N_10852,N_13740);
and U22935 (N_22935,N_18682,N_10066);
and U22936 (N_22936,N_16827,N_10833);
nor U22937 (N_22937,N_10352,N_14150);
and U22938 (N_22938,N_11719,N_19392);
nand U22939 (N_22939,N_19035,N_15104);
and U22940 (N_22940,N_14968,N_13225);
and U22941 (N_22941,N_19809,N_19592);
and U22942 (N_22942,N_13197,N_13415);
nand U22943 (N_22943,N_18514,N_18091);
and U22944 (N_22944,N_16747,N_18266);
nor U22945 (N_22945,N_15166,N_16315);
xor U22946 (N_22946,N_19003,N_13659);
and U22947 (N_22947,N_12572,N_13507);
nor U22948 (N_22948,N_19247,N_14032);
xor U22949 (N_22949,N_17181,N_15443);
xor U22950 (N_22950,N_10413,N_14546);
and U22951 (N_22951,N_14163,N_17332);
or U22952 (N_22952,N_14102,N_11911);
nor U22953 (N_22953,N_19364,N_12456);
nand U22954 (N_22954,N_11024,N_10414);
nor U22955 (N_22955,N_13716,N_18107);
nor U22956 (N_22956,N_14715,N_16689);
xnor U22957 (N_22957,N_19024,N_16283);
and U22958 (N_22958,N_15775,N_17499);
nor U22959 (N_22959,N_17226,N_16850);
nor U22960 (N_22960,N_11928,N_13074);
nor U22961 (N_22961,N_10184,N_18906);
nor U22962 (N_22962,N_16757,N_15941);
nand U22963 (N_22963,N_18818,N_17721);
and U22964 (N_22964,N_10642,N_17007);
nand U22965 (N_22965,N_10233,N_19224);
and U22966 (N_22966,N_13612,N_15788);
xor U22967 (N_22967,N_15907,N_16567);
nand U22968 (N_22968,N_19622,N_19886);
and U22969 (N_22969,N_15547,N_13832);
or U22970 (N_22970,N_17029,N_14930);
xnor U22971 (N_22971,N_18135,N_10853);
or U22972 (N_22972,N_16639,N_16213);
nand U22973 (N_22973,N_18930,N_17653);
xnor U22974 (N_22974,N_18853,N_14071);
and U22975 (N_22975,N_15376,N_13925);
or U22976 (N_22976,N_16595,N_14061);
nand U22977 (N_22977,N_12639,N_13667);
nor U22978 (N_22978,N_17527,N_10778);
or U22979 (N_22979,N_16242,N_14952);
or U22980 (N_22980,N_15627,N_17484);
nand U22981 (N_22981,N_10416,N_18139);
xor U22982 (N_22982,N_12516,N_15648);
nand U22983 (N_22983,N_19671,N_13804);
nor U22984 (N_22984,N_10334,N_12160);
nand U22985 (N_22985,N_19442,N_19038);
or U22986 (N_22986,N_15598,N_18983);
nor U22987 (N_22987,N_19562,N_19045);
and U22988 (N_22988,N_12329,N_13761);
nand U22989 (N_22989,N_19921,N_19665);
and U22990 (N_22990,N_12231,N_11121);
xor U22991 (N_22991,N_19792,N_17188);
or U22992 (N_22992,N_19009,N_19437);
xnor U22993 (N_22993,N_16119,N_15857);
or U22994 (N_22994,N_11358,N_12311);
and U22995 (N_22995,N_15812,N_15585);
or U22996 (N_22996,N_12502,N_13570);
nand U22997 (N_22997,N_14581,N_18058);
xnor U22998 (N_22998,N_16341,N_16727);
or U22999 (N_22999,N_17535,N_18634);
nor U23000 (N_23000,N_10346,N_17532);
nand U23001 (N_23001,N_18867,N_17612);
xor U23002 (N_23002,N_19657,N_12175);
or U23003 (N_23003,N_11221,N_17041);
xnor U23004 (N_23004,N_12292,N_10167);
nor U23005 (N_23005,N_17795,N_11937);
nand U23006 (N_23006,N_17675,N_19607);
or U23007 (N_23007,N_12669,N_14242);
nand U23008 (N_23008,N_12290,N_17787);
nor U23009 (N_23009,N_17247,N_10150);
or U23010 (N_23010,N_18245,N_18672);
nand U23011 (N_23011,N_16014,N_12884);
nor U23012 (N_23012,N_13976,N_17110);
nor U23013 (N_23013,N_17549,N_11278);
nor U23014 (N_23014,N_19916,N_15201);
nand U23015 (N_23015,N_12903,N_18000);
nand U23016 (N_23016,N_19362,N_17347);
nand U23017 (N_23017,N_19093,N_14404);
nand U23018 (N_23018,N_11105,N_18299);
and U23019 (N_23019,N_12517,N_11469);
and U23020 (N_23020,N_10305,N_19081);
nand U23021 (N_23021,N_18184,N_16607);
nor U23022 (N_23022,N_19236,N_18457);
or U23023 (N_23023,N_11155,N_12478);
and U23024 (N_23024,N_17777,N_19137);
and U23025 (N_23025,N_18008,N_18962);
and U23026 (N_23026,N_13360,N_14043);
nand U23027 (N_23027,N_15937,N_18464);
or U23028 (N_23028,N_18826,N_14742);
nand U23029 (N_23029,N_15839,N_11920);
xnor U23030 (N_23030,N_15366,N_12618);
xor U23031 (N_23031,N_16293,N_16225);
and U23032 (N_23032,N_10048,N_11754);
xor U23033 (N_23033,N_14558,N_18493);
xnor U23034 (N_23034,N_13382,N_17540);
nor U23035 (N_23035,N_19410,N_17292);
and U23036 (N_23036,N_11860,N_17470);
xor U23037 (N_23037,N_12229,N_15655);
xor U23038 (N_23038,N_17898,N_13304);
nand U23039 (N_23039,N_13353,N_10963);
and U23040 (N_23040,N_10064,N_12683);
nor U23041 (N_23041,N_10855,N_17193);
and U23042 (N_23042,N_14115,N_14501);
xnor U23043 (N_23043,N_18263,N_12926);
xnor U23044 (N_23044,N_19651,N_12637);
and U23045 (N_23045,N_18610,N_13038);
nor U23046 (N_23046,N_15187,N_15983);
nor U23047 (N_23047,N_12147,N_18101);
nor U23048 (N_23048,N_15794,N_17933);
nor U23049 (N_23049,N_11605,N_13317);
and U23050 (N_23050,N_13330,N_16947);
or U23051 (N_23051,N_16354,N_19602);
xor U23052 (N_23052,N_12646,N_11061);
nand U23053 (N_23053,N_11708,N_10848);
and U23054 (N_23054,N_19386,N_19596);
nand U23055 (N_23055,N_15697,N_12308);
or U23056 (N_23056,N_10994,N_14332);
or U23057 (N_23057,N_16008,N_19467);
and U23058 (N_23058,N_18319,N_12558);
nor U23059 (N_23059,N_19985,N_15991);
nand U23060 (N_23060,N_19939,N_11768);
and U23061 (N_23061,N_17599,N_14896);
nand U23062 (N_23062,N_16149,N_13018);
nor U23063 (N_23063,N_18779,N_11731);
xor U23064 (N_23064,N_15996,N_11357);
nand U23065 (N_23065,N_13118,N_19869);
nor U23066 (N_23066,N_19807,N_16125);
xor U23067 (N_23067,N_15503,N_10895);
or U23068 (N_23068,N_13215,N_11593);
and U23069 (N_23069,N_10992,N_18868);
nor U23070 (N_23070,N_10559,N_19868);
nand U23071 (N_23071,N_18762,N_15412);
and U23072 (N_23072,N_19719,N_15417);
or U23073 (N_23073,N_13842,N_16305);
xnor U23074 (N_23074,N_10041,N_12396);
nand U23075 (N_23075,N_12208,N_17845);
or U23076 (N_23076,N_19587,N_18421);
xor U23077 (N_23077,N_15325,N_16455);
and U23078 (N_23078,N_17338,N_17680);
and U23079 (N_23079,N_19113,N_18374);
or U23080 (N_23080,N_19138,N_15483);
nor U23081 (N_23081,N_17613,N_16705);
and U23082 (N_23082,N_11655,N_12153);
xnor U23083 (N_23083,N_13099,N_10159);
nand U23084 (N_23084,N_18040,N_12134);
nor U23085 (N_23085,N_10962,N_14723);
nor U23086 (N_23086,N_14072,N_15160);
or U23087 (N_23087,N_13606,N_17346);
or U23088 (N_23088,N_14281,N_16751);
and U23089 (N_23089,N_11348,N_19882);
nand U23090 (N_23090,N_14390,N_12917);
nor U23091 (N_23091,N_19696,N_14295);
xnor U23092 (N_23092,N_13793,N_17483);
or U23093 (N_23093,N_19636,N_14603);
nand U23094 (N_23094,N_13135,N_19529);
nand U23095 (N_23095,N_19801,N_12834);
nor U23096 (N_23096,N_15617,N_19047);
xor U23097 (N_23097,N_10424,N_15921);
xor U23098 (N_23098,N_16047,N_13679);
and U23099 (N_23099,N_19735,N_12230);
or U23100 (N_23100,N_19648,N_12779);
or U23101 (N_23101,N_13294,N_16199);
and U23102 (N_23102,N_16482,N_14127);
nand U23103 (N_23103,N_11767,N_12131);
nor U23104 (N_23104,N_17207,N_14987);
xnor U23105 (N_23105,N_17837,N_10913);
or U23106 (N_23106,N_18997,N_14731);
nand U23107 (N_23107,N_17730,N_11383);
xor U23108 (N_23108,N_16840,N_15929);
xnor U23109 (N_23109,N_17322,N_11543);
and U23110 (N_23110,N_14915,N_19880);
nand U23111 (N_23111,N_13729,N_17468);
nor U23112 (N_23112,N_10528,N_12224);
nand U23113 (N_23113,N_10420,N_18361);
or U23114 (N_23114,N_18083,N_18370);
and U23115 (N_23115,N_13096,N_12666);
or U23116 (N_23116,N_18018,N_10302);
xor U23117 (N_23117,N_17879,N_12044);
nand U23118 (N_23118,N_19229,N_18451);
nor U23119 (N_23119,N_10382,N_11145);
nand U23120 (N_23120,N_11119,N_12928);
or U23121 (N_23121,N_16450,N_12309);
xnor U23122 (N_23122,N_11241,N_11211);
nor U23123 (N_23123,N_18638,N_15933);
nand U23124 (N_23124,N_13782,N_13470);
nor U23125 (N_23125,N_13956,N_15614);
or U23126 (N_23126,N_11458,N_17415);
and U23127 (N_23127,N_11057,N_14818);
or U23128 (N_23128,N_15250,N_16490);
nand U23129 (N_23129,N_12555,N_17546);
xnor U23130 (N_23130,N_15860,N_18148);
xnor U23131 (N_23131,N_17786,N_10428);
or U23132 (N_23132,N_11077,N_11827);
xor U23133 (N_23133,N_15190,N_10155);
nand U23134 (N_23134,N_12029,N_12067);
and U23135 (N_23135,N_19382,N_11923);
or U23136 (N_23136,N_10615,N_11460);
nand U23137 (N_23137,N_15877,N_15553);
and U23138 (N_23138,N_17472,N_12371);
nor U23139 (N_23139,N_10885,N_13435);
and U23140 (N_23140,N_17100,N_18271);
nor U23141 (N_23141,N_13637,N_17892);
and U23142 (N_23142,N_15304,N_10514);
nand U23143 (N_23143,N_19759,N_18999);
xor U23144 (N_23144,N_16714,N_13889);
or U23145 (N_23145,N_19996,N_10138);
nor U23146 (N_23146,N_18386,N_16191);
nand U23147 (N_23147,N_11432,N_16851);
xor U23148 (N_23148,N_10160,N_17184);
xor U23149 (N_23149,N_13422,N_10432);
or U23150 (N_23150,N_19130,N_15299);
nand U23151 (N_23151,N_15364,N_19015);
nor U23152 (N_23152,N_14711,N_10760);
nor U23153 (N_23153,N_15247,N_18967);
or U23154 (N_23154,N_11542,N_17749);
nor U23155 (N_23155,N_14224,N_18783);
xor U23156 (N_23156,N_16173,N_12811);
nor U23157 (N_23157,N_10526,N_14097);
and U23158 (N_23158,N_13578,N_11274);
xor U23159 (N_23159,N_16483,N_10459);
or U23160 (N_23160,N_18870,N_17341);
or U23161 (N_23161,N_17979,N_19014);
xor U23162 (N_23162,N_18123,N_12974);
nand U23163 (N_23163,N_12150,N_11766);
xnor U23164 (N_23164,N_19208,N_17723);
or U23165 (N_23165,N_14296,N_17305);
or U23166 (N_23166,N_18194,N_17807);
or U23167 (N_23167,N_19075,N_12117);
or U23168 (N_23168,N_18060,N_19010);
nand U23169 (N_23169,N_11563,N_13354);
and U23170 (N_23170,N_14665,N_15257);
nor U23171 (N_23171,N_14256,N_17677);
or U23172 (N_23172,N_18437,N_10674);
or U23173 (N_23173,N_19773,N_17593);
nand U23174 (N_23174,N_13970,N_16784);
nor U23175 (N_23175,N_16410,N_13573);
nand U23176 (N_23176,N_18416,N_17183);
xnor U23177 (N_23177,N_13809,N_17764);
or U23178 (N_23178,N_15134,N_18855);
and U23179 (N_23179,N_19722,N_18439);
xor U23180 (N_23180,N_14476,N_17685);
and U23181 (N_23181,N_12778,N_15301);
and U23182 (N_23182,N_17903,N_19485);
nand U23183 (N_23183,N_15359,N_14356);
and U23184 (N_23184,N_13738,N_13596);
and U23185 (N_23185,N_17259,N_10204);
or U23186 (N_23186,N_19800,N_17127);
or U23187 (N_23187,N_14789,N_10958);
or U23188 (N_23188,N_12357,N_16308);
nand U23189 (N_23189,N_10393,N_15568);
xor U23190 (N_23190,N_15080,N_17123);
nor U23191 (N_23191,N_18714,N_17690);
nor U23192 (N_23192,N_17687,N_10849);
and U23193 (N_23193,N_16192,N_11507);
nand U23194 (N_23194,N_13179,N_14450);
and U23195 (N_23195,N_15264,N_19823);
nor U23196 (N_23196,N_10172,N_16649);
and U23197 (N_23197,N_19115,N_13544);
or U23198 (N_23198,N_11236,N_15815);
and U23199 (N_23199,N_19335,N_13042);
nand U23200 (N_23200,N_17823,N_11564);
xor U23201 (N_23201,N_15835,N_13916);
nand U23202 (N_23202,N_12193,N_17458);
nor U23203 (N_23203,N_17021,N_19029);
or U23204 (N_23204,N_14052,N_11398);
xnor U23205 (N_23205,N_15680,N_14664);
and U23206 (N_23206,N_19705,N_14271);
or U23207 (N_23207,N_13605,N_13395);
or U23208 (N_23208,N_12989,N_11749);
xnor U23209 (N_23209,N_18848,N_15101);
and U23210 (N_23210,N_12106,N_10791);
or U23211 (N_23211,N_16681,N_13710);
or U23212 (N_23212,N_14869,N_15063);
nor U23213 (N_23213,N_19680,N_13149);
nor U23214 (N_23214,N_16842,N_18200);
nand U23215 (N_23215,N_19763,N_15679);
and U23216 (N_23216,N_14192,N_11693);
or U23217 (N_23217,N_17311,N_19301);
nand U23218 (N_23218,N_13080,N_16330);
and U23219 (N_23219,N_12796,N_13699);
or U23220 (N_23220,N_14432,N_18192);
nand U23221 (N_23221,N_15529,N_12577);
nand U23222 (N_23222,N_17834,N_11298);
xnor U23223 (N_23223,N_17626,N_10283);
nand U23224 (N_23224,N_17576,N_16409);
or U23225 (N_23225,N_10192,N_12580);
or U23226 (N_23226,N_11676,N_13176);
nand U23227 (N_23227,N_11874,N_18660);
and U23228 (N_23228,N_10391,N_14802);
and U23229 (N_23229,N_14891,N_18026);
and U23230 (N_23230,N_12058,N_15992);
xor U23231 (N_23231,N_11417,N_13643);
xnor U23232 (N_23232,N_15320,N_13365);
nor U23233 (N_23233,N_16487,N_15511);
nand U23234 (N_23234,N_10469,N_16475);
nor U23235 (N_23235,N_16959,N_19375);
xor U23236 (N_23236,N_17046,N_10942);
nor U23237 (N_23237,N_19571,N_16428);
and U23238 (N_23238,N_19216,N_16323);
nor U23239 (N_23239,N_13589,N_19894);
and U23240 (N_23240,N_10007,N_16397);
and U23241 (N_23241,N_14800,N_10154);
nand U23242 (N_23242,N_18124,N_11435);
nor U23243 (N_23243,N_10901,N_10324);
xnor U23244 (N_23244,N_18998,N_18371);
or U23245 (N_23245,N_12887,N_17797);
or U23246 (N_23246,N_19169,N_14187);
xnor U23247 (N_23247,N_13575,N_13106);
nand U23248 (N_23248,N_10270,N_15302);
and U23249 (N_23249,N_10457,N_14029);
and U23250 (N_23250,N_15231,N_19298);
or U23251 (N_23251,N_12138,N_15438);
nor U23252 (N_23252,N_17973,N_18988);
and U23253 (N_23253,N_12442,N_12317);
and U23254 (N_23254,N_12578,N_12251);
or U23255 (N_23255,N_17386,N_11144);
xnor U23256 (N_23256,N_14808,N_15741);
xor U23257 (N_23257,N_11180,N_19339);
nor U23258 (N_23258,N_15300,N_10485);
or U23259 (N_23259,N_15219,N_17699);
nand U23260 (N_23260,N_14845,N_14025);
nor U23261 (N_23261,N_13231,N_14589);
nor U23262 (N_23262,N_19511,N_19654);
and U23263 (N_23263,N_17520,N_18256);
or U23264 (N_23264,N_16467,N_15986);
or U23265 (N_23265,N_17249,N_11918);
xnor U23266 (N_23266,N_15239,N_18460);
xnor U23267 (N_23267,N_17961,N_13749);
xnor U23268 (N_23268,N_15657,N_14445);
xor U23269 (N_23269,N_13515,N_13203);
nor U23270 (N_23270,N_19775,N_18097);
nor U23271 (N_23271,N_11875,N_10775);
xnor U23272 (N_23272,N_17286,N_11877);
xor U23273 (N_23273,N_12426,N_12849);
and U23274 (N_23274,N_14399,N_19750);
or U23275 (N_23275,N_17645,N_15131);
or U23276 (N_23276,N_11509,N_16655);
and U23277 (N_23277,N_14837,N_17089);
or U23278 (N_23278,N_10209,N_10961);
or U23279 (N_23279,N_10092,N_15763);
nor U23280 (N_23280,N_16524,N_18140);
xor U23281 (N_23281,N_14363,N_10951);
and U23282 (N_23282,N_14566,N_10956);
nor U23283 (N_23283,N_19126,N_18995);
xnor U23284 (N_23284,N_17009,N_12082);
nand U23285 (N_23285,N_18796,N_12542);
xor U23286 (N_23286,N_10037,N_17491);
or U23287 (N_23287,N_14701,N_19102);
or U23288 (N_23288,N_11735,N_19135);
and U23289 (N_23289,N_18161,N_13026);
nor U23290 (N_23290,N_16402,N_18659);
xor U23291 (N_23291,N_11759,N_10026);
nand U23292 (N_23292,N_11503,N_14290);
nor U23293 (N_23293,N_12705,N_13490);
and U23294 (N_23294,N_16582,N_15924);
or U23295 (N_23295,N_11201,N_19232);
and U23296 (N_23296,N_17746,N_19031);
and U23297 (N_23297,N_18325,N_18424);
nor U23298 (N_23298,N_18295,N_18985);
and U23299 (N_23299,N_12929,N_11163);
nand U23300 (N_23300,N_11628,N_14916);
xor U23301 (N_23301,N_11624,N_11910);
xnor U23302 (N_23302,N_13166,N_10554);
nor U23303 (N_23303,N_14309,N_16877);
xnor U23304 (N_23304,N_19424,N_13844);
nor U23305 (N_23305,N_15765,N_15293);
nand U23306 (N_23306,N_12048,N_18149);
nand U23307 (N_23307,N_11246,N_17710);
nand U23308 (N_23308,N_15111,N_14478);
or U23309 (N_23309,N_19415,N_17917);
and U23310 (N_23310,N_10321,N_14494);
and U23311 (N_23311,N_12019,N_19827);
and U23312 (N_23312,N_18953,N_18316);
xor U23313 (N_23313,N_10977,N_16937);
nand U23314 (N_23314,N_17160,N_14892);
xor U23315 (N_23315,N_10816,N_14629);
or U23316 (N_23316,N_14746,N_15244);
and U23317 (N_23317,N_13966,N_18794);
nor U23318 (N_23318,N_18498,N_13652);
xnor U23319 (N_23319,N_14512,N_10661);
or U23320 (N_23320,N_18732,N_17665);
or U23321 (N_23321,N_14172,N_19156);
xnor U23322 (N_23322,N_13071,N_15332);
or U23323 (N_23323,N_11648,N_18628);
nor U23324 (N_23324,N_15685,N_18492);
nor U23325 (N_23325,N_10826,N_15148);
or U23326 (N_23326,N_18032,N_15284);
and U23327 (N_23327,N_14710,N_15309);
and U23328 (N_23328,N_19934,N_17495);
nor U23329 (N_23329,N_19563,N_16902);
nand U23330 (N_23330,N_13776,N_15988);
or U23331 (N_23331,N_19710,N_12013);
and U23332 (N_23332,N_11963,N_14156);
xor U23333 (N_23333,N_18344,N_17159);
nand U23334 (N_23334,N_17934,N_13468);
xor U23335 (N_23335,N_14096,N_10215);
nand U23336 (N_23336,N_10987,N_19107);
and U23337 (N_23337,N_19746,N_17781);
and U23338 (N_23338,N_17304,N_13930);
xor U23339 (N_23339,N_12695,N_13829);
nand U23340 (N_23340,N_12462,N_19736);
nor U23341 (N_23341,N_12785,N_11352);
and U23342 (N_23342,N_13639,N_11589);
or U23343 (N_23343,N_11861,N_19193);
nand U23344 (N_23344,N_15809,N_12101);
or U23345 (N_23345,N_19080,N_16106);
nand U23346 (N_23346,N_11450,N_10576);
and U23347 (N_23347,N_15742,N_17174);
and U23348 (N_23348,N_11777,N_18150);
nand U23349 (N_23349,N_14007,N_14331);
nand U23350 (N_23350,N_13127,N_19818);
and U23351 (N_23351,N_12035,N_16688);
nand U23352 (N_23352,N_10735,N_19770);
xnor U23353 (N_23353,N_16919,N_14985);
nand U23354 (N_23354,N_18755,N_14132);
nand U23355 (N_23355,N_16909,N_12098);
xor U23356 (N_23356,N_12367,N_14304);
xor U23357 (N_23357,N_17594,N_18880);
xnor U23358 (N_23358,N_15075,N_16766);
xnor U23359 (N_23359,N_17129,N_17931);
and U23360 (N_23360,N_19683,N_18209);
and U23361 (N_23361,N_13982,N_11879);
and U23362 (N_23362,N_19303,N_17306);
nor U23363 (N_23363,N_15823,N_16980);
nor U23364 (N_23364,N_18615,N_19900);
or U23365 (N_23365,N_17357,N_10297);
or U23366 (N_23366,N_17280,N_19594);
xor U23367 (N_23367,N_12620,N_16005);
nand U23368 (N_23368,N_10543,N_19993);
or U23369 (N_23369,N_16140,N_19428);
xor U23370 (N_23370,N_15342,N_13424);
and U23371 (N_23371,N_13974,N_16039);
and U23372 (N_23372,N_10898,N_14414);
nand U23373 (N_23373,N_16941,N_18799);
nor U23374 (N_23374,N_18566,N_12036);
nand U23375 (N_23375,N_19777,N_17566);
nor U23376 (N_23376,N_14303,N_10560);
or U23377 (N_23377,N_18281,N_18694);
and U23378 (N_23378,N_11150,N_19958);
nor U23379 (N_23379,N_13133,N_17551);
nand U23380 (N_23380,N_18029,N_18574);
xor U23381 (N_23381,N_16791,N_16927);
or U23382 (N_23382,N_12918,N_11086);
nand U23383 (N_23383,N_14893,N_11261);
xor U23384 (N_23384,N_19023,N_10463);
nor U23385 (N_23385,N_10677,N_11202);
xor U23386 (N_23386,N_18067,N_11733);
and U23387 (N_23387,N_15379,N_12301);
nand U23388 (N_23388,N_17229,N_15005);
and U23389 (N_23389,N_12016,N_17354);
xnor U23390 (N_23390,N_16799,N_17445);
and U23391 (N_23391,N_18550,N_10664);
nor U23392 (N_23392,N_11926,N_16861);
xor U23393 (N_23393,N_14872,N_17402);
xnor U23394 (N_23394,N_14346,N_18378);
nor U23395 (N_23395,N_11491,N_19309);
nor U23396 (N_23396,N_15277,N_14706);
nor U23397 (N_23397,N_11248,N_12824);
nor U23398 (N_23398,N_15886,N_12731);
xor U23399 (N_23399,N_15825,N_16289);
and U23400 (N_23400,N_16294,N_14358);
or U23401 (N_23401,N_15870,N_14971);
or U23402 (N_23402,N_16933,N_14459);
nor U23403 (N_23403,N_11824,N_11974);
or U23404 (N_23404,N_13723,N_18708);
xor U23405 (N_23405,N_18168,N_10121);
nand U23406 (N_23406,N_19332,N_19181);
nand U23407 (N_23407,N_17269,N_13110);
nand U23408 (N_23408,N_14763,N_12097);
nand U23409 (N_23409,N_18927,N_14145);
xnor U23410 (N_23410,N_12195,N_15574);
nand U23411 (N_23411,N_19981,N_17562);
nand U23412 (N_23412,N_14508,N_15383);
nor U23413 (N_23413,N_12266,N_19148);
or U23414 (N_23414,N_12738,N_14736);
or U23415 (N_23415,N_12941,N_11560);
and U23416 (N_23416,N_13160,N_17300);
nand U23417 (N_23417,N_14749,N_15619);
or U23418 (N_23418,N_11620,N_19128);
or U23419 (N_23419,N_11578,N_16288);
nand U23420 (N_23420,N_17610,N_18847);
xnor U23421 (N_23421,N_17714,N_17835);
nand U23422 (N_23422,N_14101,N_18189);
xor U23423 (N_23423,N_16873,N_12418);
nor U23424 (N_23424,N_12893,N_10946);
and U23425 (N_23425,N_17119,N_12810);
or U23426 (N_23426,N_13427,N_13807);
nor U23427 (N_23427,N_13757,N_19682);
nand U23428 (N_23428,N_10687,N_18222);
and U23429 (N_23429,N_15573,N_19213);
or U23430 (N_23430,N_10455,N_16869);
nand U23431 (N_23431,N_16601,N_12664);
nor U23432 (N_23432,N_10377,N_10481);
and U23433 (N_23433,N_15868,N_11774);
xor U23434 (N_23434,N_15784,N_16629);
nand U23435 (N_23435,N_15543,N_16894);
and U23436 (N_23436,N_12630,N_10647);
and U23437 (N_23437,N_18205,N_11843);
or U23438 (N_23438,N_19280,N_16296);
and U23439 (N_23439,N_19166,N_10218);
nand U23440 (N_23440,N_10782,N_12112);
xnor U23441 (N_23441,N_19159,N_16609);
or U23442 (N_23442,N_11242,N_15561);
and U23443 (N_23443,N_15177,N_19374);
or U23444 (N_23444,N_18807,N_11977);
or U23445 (N_23445,N_12458,N_15025);
nor U23446 (N_23446,N_12851,N_19350);
and U23447 (N_23447,N_14444,N_16958);
xor U23448 (N_23448,N_13626,N_17672);
or U23449 (N_23449,N_16395,N_19690);
xor U23450 (N_23450,N_11249,N_12706);
or U23451 (N_23451,N_11051,N_15911);
xor U23452 (N_23452,N_11406,N_11859);
or U23453 (N_23453,N_14695,N_19062);
and U23454 (N_23454,N_16903,N_18249);
and U23455 (N_23455,N_17869,N_15532);
xor U23456 (N_23456,N_19435,N_13676);
and U23457 (N_23457,N_10690,N_10013);
and U23458 (N_23458,N_12792,N_13193);
xor U23459 (N_23459,N_19769,N_15281);
or U23460 (N_23460,N_12740,N_13310);
nor U23461 (N_23461,N_16322,N_15688);
or U23462 (N_23462,N_13661,N_16377);
or U23463 (N_23463,N_14674,N_17204);
xor U23464 (N_23464,N_12569,N_15799);
and U23465 (N_23465,N_11902,N_10100);
nor U23466 (N_23466,N_13414,N_16891);
nor U23467 (N_23467,N_13975,N_13011);
xor U23468 (N_23468,N_12047,N_10743);
and U23469 (N_23469,N_16920,N_18356);
nor U23470 (N_23470,N_17380,N_18522);
xor U23471 (N_23471,N_11052,N_17137);
nand U23472 (N_23472,N_18837,N_18842);
nand U23473 (N_23473,N_11515,N_13594);
and U23474 (N_23474,N_13142,N_15790);
and U23475 (N_23475,N_13343,N_12791);
xnor U23476 (N_23476,N_18273,N_15682);
nor U23477 (N_23477,N_18041,N_19125);
nor U23478 (N_23478,N_15441,N_11463);
nor U23479 (N_23479,N_18462,N_19203);
nor U23480 (N_23480,N_16855,N_13327);
nand U23481 (N_23481,N_12762,N_14136);
xnor U23482 (N_23482,N_14405,N_12412);
xor U23483 (N_23483,N_10644,N_18652);
nor U23484 (N_23484,N_17762,N_18790);
nand U23485 (N_23485,N_15618,N_10329);
xor U23486 (N_23486,N_18992,N_10301);
or U23487 (N_23487,N_18943,N_15262);
nand U23488 (N_23488,N_13457,N_11897);
nor U23489 (N_23489,N_12761,N_10874);
nor U23490 (N_23490,N_18965,N_14385);
nand U23491 (N_23491,N_18475,N_18210);
and U23492 (N_23492,N_18553,N_13980);
or U23493 (N_23493,N_18224,N_16908);
nand U23494 (N_23494,N_13394,N_12912);
xor U23495 (N_23495,N_13863,N_17018);
nor U23496 (N_23496,N_11612,N_17048);
nand U23497 (N_23497,N_10123,N_12735);
xnor U23498 (N_23498,N_17624,N_16558);
nor U23499 (N_23499,N_19393,N_14157);
nand U23500 (N_23500,N_14721,N_15462);
and U23501 (N_23501,N_15064,N_11396);
and U23502 (N_23502,N_15348,N_16987);
nand U23503 (N_23503,N_12540,N_14142);
nand U23504 (N_23504,N_13638,N_16151);
and U23505 (N_23505,N_17241,N_14251);
nor U23506 (N_23506,N_14619,N_10638);
nand U23507 (N_23507,N_13480,N_12286);
and U23508 (N_23508,N_13447,N_12767);
xnor U23509 (N_23509,N_16427,N_19954);
nor U23510 (N_23510,N_10250,N_17308);
or U23511 (N_23511,N_18587,N_10605);
nand U23512 (N_23512,N_15634,N_10809);
or U23513 (N_23513,N_11390,N_12665);
xor U23514 (N_23514,N_16425,N_10241);
nor U23515 (N_23515,N_11269,N_15905);
and U23516 (N_23516,N_18275,N_15705);
and U23517 (N_23517,N_17016,N_19273);
nand U23518 (N_23518,N_16155,N_13357);
xor U23519 (N_23519,N_10877,N_11440);
or U23520 (N_23520,N_10072,N_12275);
nand U23521 (N_23521,N_13378,N_11758);
xnor U23522 (N_23522,N_13006,N_16740);
or U23523 (N_23523,N_11149,N_13867);
xor U23524 (N_23524,N_16403,N_16302);
nor U23525 (N_23525,N_12154,N_14509);
xnor U23526 (N_23526,N_17462,N_12420);
nor U23527 (N_23527,N_11993,N_16748);
and U23528 (N_23528,N_19998,N_10142);
and U23529 (N_23529,N_17152,N_18181);
or U23530 (N_23530,N_19317,N_11688);
nand U23531 (N_23531,N_19400,N_18214);
or U23532 (N_23532,N_12254,N_17962);
or U23533 (N_23533,N_16153,N_13221);
nor U23534 (N_23534,N_17999,N_17344);
nor U23535 (N_23535,N_11436,N_15109);
xor U23536 (N_23536,N_15368,N_14175);
or U23537 (N_23537,N_10715,N_10060);
xnor U23538 (N_23538,N_18100,N_11650);
and U23539 (N_23539,N_13323,N_14125);
or U23540 (N_23540,N_11858,N_19312);
and U23541 (N_23541,N_10359,N_14048);
nand U23542 (N_23542,N_15274,N_19401);
nor U23543 (N_23543,N_12545,N_12956);
xor U23544 (N_23544,N_11371,N_15516);
and U23545 (N_23545,N_16580,N_18227);
xor U23546 (N_23546,N_14235,N_14243);
nor U23547 (N_23547,N_16358,N_10641);
and U23548 (N_23548,N_15180,N_13913);
nor U23549 (N_23549,N_17771,N_13008);
and U23550 (N_23550,N_10051,N_12977);
xor U23551 (N_23551,N_19131,N_18850);
nor U23552 (N_23552,N_19162,N_15640);
or U23553 (N_23553,N_14737,N_12993);
xor U23554 (N_23554,N_16257,N_14585);
or U23555 (N_23555,N_11038,N_17418);
xor U23556 (N_23556,N_15474,N_13835);
nand U23557 (N_23557,N_15738,N_15587);
or U23558 (N_23558,N_15279,N_10894);
or U23559 (N_23559,N_10712,N_14112);
and U23560 (N_23560,N_18639,N_17910);
and U23561 (N_23561,N_11753,N_16393);
or U23562 (N_23562,N_15527,N_14522);
xor U23563 (N_23563,N_17399,N_16072);
nand U23564 (N_23564,N_19520,N_14020);
nand U23565 (N_23565,N_18404,N_10535);
or U23566 (N_23566,N_17441,N_15595);
or U23567 (N_23567,N_16284,N_15536);
nand U23568 (N_23568,N_14229,N_17372);
xnor U23569 (N_23569,N_12861,N_14250);
xor U23570 (N_23570,N_17768,N_16940);
and U23571 (N_23571,N_10692,N_14655);
and U23572 (N_23572,N_13897,N_14291);
nor U23573 (N_23573,N_16006,N_14935);
nor U23574 (N_23574,N_14483,N_15821);
xor U23575 (N_23575,N_12548,N_11342);
and U23576 (N_23576,N_12749,N_16063);
and U23577 (N_23577,N_17858,N_13984);
xor U23578 (N_23578,N_14524,N_12350);
nand U23579 (N_23579,N_18405,N_12523);
nor U23580 (N_23580,N_16797,N_15854);
nand U23581 (N_23581,N_18490,N_11198);
or U23582 (N_23582,N_19588,N_15410);
xor U23583 (N_23583,N_19659,N_19738);
nand U23584 (N_23584,N_15234,N_15912);
xnor U23585 (N_23585,N_14909,N_10926);
xor U23586 (N_23586,N_15506,N_15404);
nor U23587 (N_23587,N_16227,N_13012);
or U23588 (N_23588,N_19687,N_16297);
xor U23589 (N_23589,N_19949,N_11059);
nor U23590 (N_23590,N_19205,N_19360);
xnor U23591 (N_23591,N_12972,N_18996);
nand U23592 (N_23592,N_17608,N_17321);
and U23593 (N_23593,N_13329,N_18697);
nor U23594 (N_23594,N_16090,N_19285);
nor U23595 (N_23595,N_11872,N_19460);
xor U23596 (N_23596,N_11415,N_17387);
and U23597 (N_23597,N_17533,N_19153);
xnor U23598 (N_23598,N_10612,N_14263);
nand U23599 (N_23599,N_17681,N_15969);
nand U23600 (N_23600,N_13514,N_13072);
xnor U23601 (N_23601,N_10316,N_18798);
xor U23602 (N_23602,N_14185,N_10152);
nor U23603 (N_23603,N_14298,N_12130);
nor U23604 (N_23604,N_11473,N_17560);
nor U23605 (N_23605,N_17528,N_15918);
nor U23606 (N_23606,N_14972,N_12351);
or U23607 (N_23607,N_12033,N_19611);
or U23608 (N_23608,N_19897,N_13754);
nand U23609 (N_23609,N_16535,N_13031);
nor U23610 (N_23610,N_16416,N_18169);
nand U23611 (N_23611,N_10388,N_13409);
xnor U23612 (N_23612,N_12830,N_14499);
nor U23613 (N_23613,N_19925,N_15761);
nor U23614 (N_23614,N_10296,N_11431);
and U23615 (N_23615,N_18756,N_11411);
nor U23616 (N_23616,N_12687,N_16522);
and U23617 (N_23617,N_14038,N_13396);
xor U23618 (N_23618,N_16917,N_15027);
nand U23619 (N_23619,N_10875,N_17791);
and U23620 (N_23620,N_15012,N_12484);
nand U23621 (N_23621,N_11327,N_17488);
nand U23622 (N_23622,N_12284,N_14648);
xnor U23623 (N_23623,N_19163,N_19347);
xnor U23624 (N_23624,N_17770,N_10568);
nand U23625 (N_23625,N_19149,N_11905);
and U23626 (N_23626,N_18244,N_18166);
xnor U23627 (N_23627,N_10307,N_11359);
xor U23628 (N_23628,N_13130,N_19521);
and U23629 (N_23629,N_11932,N_15945);
nor U23630 (N_23630,N_10332,N_15662);
or U23631 (N_23631,N_18010,N_15276);
or U23632 (N_23632,N_12936,N_16052);
nor U23633 (N_23633,N_12795,N_19821);
and U23634 (N_23634,N_18573,N_13112);
nor U23635 (N_23635,N_11397,N_19783);
or U23636 (N_23636,N_18877,N_15213);
or U23637 (N_23637,N_17741,N_12043);
and U23638 (N_23638,N_13669,N_15646);
nor U23639 (N_23639,N_12752,N_15402);
nor U23640 (N_23640,N_15303,N_15298);
nand U23641 (N_23641,N_12294,N_14026);
and U23642 (N_23642,N_12742,N_14599);
and U23643 (N_23643,N_16080,N_18805);
xor U23644 (N_23644,N_16197,N_16448);
xnor U23645 (N_23645,N_16634,N_18068);
nand U23646 (N_23646,N_14359,N_12688);
or U23647 (N_23647,N_13988,N_11567);
nand U23648 (N_23648,N_18506,N_19500);
xnor U23649 (N_23649,N_17849,N_19293);
and U23650 (N_23650,N_12565,N_12407);
and U23651 (N_23651,N_12084,N_17143);
nand U23652 (N_23652,N_13440,N_10389);
xnor U23653 (N_23653,N_18056,N_12900);
or U23654 (N_23654,N_16830,N_10333);
and U23655 (N_23655,N_14782,N_16767);
nor U23656 (N_23656,N_19432,N_17250);
xor U23657 (N_23657,N_11490,N_15963);
or U23658 (N_23658,N_13201,N_17646);
nand U23659 (N_23659,N_16912,N_15036);
and U23660 (N_23660,N_13014,N_15760);
nand U23661 (N_23661,N_16899,N_14515);
xnor U23662 (N_23662,N_17417,N_17274);
xor U23663 (N_23663,N_11301,N_19830);
nand U23664 (N_23664,N_10235,N_13064);
nor U23665 (N_23665,N_14247,N_15894);
nor U23666 (N_23666,N_19353,N_14852);
nor U23667 (N_23667,N_11913,N_13054);
or U23668 (N_23668,N_17928,N_12474);
nor U23669 (N_23669,N_10125,N_17392);
and U23670 (N_23670,N_17775,N_13756);
or U23671 (N_23671,N_14149,N_17455);
nand U23672 (N_23672,N_16965,N_12692);
nand U23673 (N_23673,N_13847,N_17774);
nand U23674 (N_23674,N_12409,N_14227);
xnor U23675 (N_23675,N_10249,N_17796);
and U23676 (N_23676,N_15732,N_15403);
and U23677 (N_23677,N_13821,N_18831);
xnor U23678 (N_23678,N_14161,N_16129);
xnor U23679 (N_23679,N_13338,N_16458);
or U23680 (N_23680,N_16195,N_17725);
and U23681 (N_23681,N_17669,N_18283);
nor U23682 (N_23682,N_18679,N_13647);
and U23683 (N_23683,N_12554,N_10312);
or U23684 (N_23684,N_16803,N_11745);
nand U23685 (N_23685,N_11736,N_18086);
nor U23686 (N_23686,N_17521,N_10470);
nand U23687 (N_23687,N_18389,N_12845);
and U23688 (N_23688,N_13959,N_10165);
and U23689 (N_23689,N_13141,N_11245);
xnor U23690 (N_23690,N_16654,N_19963);
nand U23691 (N_23691,N_13191,N_19496);
and U23692 (N_23692,N_17863,N_17936);
nand U23693 (N_23693,N_17157,N_19546);
nor U23694 (N_23694,N_14239,N_16808);
or U23695 (N_23695,N_16507,N_15895);
xnor U23696 (N_23696,N_17273,N_16889);
and U23697 (N_23697,N_10827,N_17456);
nor U23698 (N_23698,N_10452,N_13853);
nand U23699 (N_23699,N_19018,N_12279);
xor U23700 (N_23700,N_18243,N_14044);
nand U23701 (N_23701,N_19670,N_18412);
xnor U23702 (N_23702,N_14905,N_16046);
nor U23703 (N_23703,N_15447,N_18019);
nand U23704 (N_23704,N_19021,N_10818);
and U23705 (N_23705,N_18772,N_12916);
nor U23706 (N_23706,N_16966,N_19445);
or U23707 (N_23707,N_16141,N_12850);
xor U23708 (N_23708,N_10771,N_11572);
xor U23709 (N_23709,N_10863,N_14166);
nand U23710 (N_23710,N_14231,N_11237);
nand U23711 (N_23711,N_15069,N_12818);
xor U23712 (N_23712,N_19302,N_16970);
and U23713 (N_23713,N_15703,N_13369);
nand U23714 (N_23714,N_17632,N_10813);
nand U23715 (N_23715,N_19324,N_19988);
xor U23716 (N_23716,N_16657,N_16907);
nor U23717 (N_23717,N_18895,N_18705);
xor U23718 (N_23718,N_12816,N_13517);
nand U23719 (N_23719,N_15232,N_12300);
or U23720 (N_23720,N_17398,N_13235);
nand U23721 (N_23721,N_19875,N_11131);
xnor U23722 (N_23722,N_15315,N_17423);
xor U23723 (N_23723,N_11457,N_17190);
nor U23724 (N_23724,N_14815,N_11447);
and U23725 (N_23725,N_14727,N_18278);
or U23726 (N_23726,N_15034,N_14225);
nor U23727 (N_23727,N_13115,N_17431);
nor U23728 (N_23728,N_18701,N_16829);
nand U23729 (N_23729,N_12415,N_11334);
nor U23730 (N_23730,N_15214,N_16206);
or U23731 (N_23731,N_16708,N_19540);
nor U23732 (N_23732,N_11580,N_11718);
nand U23733 (N_23733,N_17886,N_13361);
nand U23734 (N_23734,N_15957,N_16160);
nand U23735 (N_23735,N_13186,N_19879);
and U23736 (N_23736,N_12273,N_12370);
and U23737 (N_23737,N_10693,N_10825);
xnor U23738 (N_23738,N_17574,N_17314);
nand U23739 (N_23739,N_16570,N_11935);
nand U23740 (N_23740,N_16717,N_13234);
xor U23741 (N_23741,N_12417,N_13533);
nand U23742 (N_23742,N_15140,N_13929);
nand U23743 (N_23743,N_16694,N_13326);
and U23744 (N_23744,N_14266,N_15950);
nand U23745 (N_23745,N_16684,N_18003);
nor U23746 (N_23746,N_12086,N_12004);
nand U23747 (N_23747,N_14351,N_12642);
or U23748 (N_23748,N_19363,N_19395);
and U23749 (N_23749,N_10844,N_16040);
or U23750 (N_23750,N_12798,N_19147);
nand U23751 (N_23751,N_12479,N_10018);
and U23752 (N_23752,N_11673,N_14534);
nor U23753 (N_23753,N_12726,N_13498);
nand U23754 (N_23754,N_14342,N_19099);
or U23755 (N_23755,N_17496,N_15152);
nand U23756 (N_23756,N_13287,N_16993);
or U23757 (N_23757,N_16328,N_11183);
nand U23758 (N_23758,N_11889,N_13820);
xnor U23759 (N_23759,N_15779,N_14087);
nand U23760 (N_23760,N_10598,N_15142);
or U23761 (N_23761,N_17086,N_16957);
or U23762 (N_23762,N_15128,N_18950);
or U23763 (N_23763,N_14532,N_10976);
or U23764 (N_23764,N_19154,N_11637);
nor U23765 (N_23765,N_13502,N_17867);
nand U23766 (N_23766,N_12486,N_19798);
and U23767 (N_23767,N_17153,N_14575);
and U23768 (N_23768,N_15210,N_16529);
nor U23769 (N_23769,N_13237,N_14612);
xor U23770 (N_23770,N_11691,N_19655);
xnor U23771 (N_23771,N_17859,N_13144);
or U23772 (N_23772,N_10448,N_12754);
or U23773 (N_23773,N_16383,N_17449);
xnor U23774 (N_23774,N_16592,N_15726);
and U23775 (N_23775,N_18945,N_12190);
and U23776 (N_23776,N_16795,N_16246);
or U23777 (N_23777,N_17437,N_11120);
and U23778 (N_23778,N_11531,N_15635);
and U23779 (N_23779,N_16950,N_12440);
and U23780 (N_23780,N_17679,N_19895);
xor U23781 (N_23781,N_13990,N_19140);
xnor U23782 (N_23782,N_19160,N_12571);
or U23783 (N_23783,N_19065,N_19638);
nand U23784 (N_23784,N_11294,N_10487);
xnor U23785 (N_23785,N_14049,N_19030);
nor U23786 (N_23786,N_12663,N_12271);
and U23787 (N_23787,N_17172,N_13093);
or U23788 (N_23788,N_17454,N_19740);
xnor U23789 (N_23789,N_12793,N_10430);
nand U23790 (N_23790,N_17814,N_16437);
nor U23791 (N_23791,N_12943,N_10063);
xor U23792 (N_23792,N_13478,N_15592);
nand U23793 (N_23793,N_12027,N_17716);
nand U23794 (N_23794,N_17135,N_17694);
nand U23795 (N_23795,N_19964,N_18442);
nand U23796 (N_23796,N_19647,N_14973);
and U23797 (N_23797,N_14774,N_17854);
and U23798 (N_23798,N_12509,N_15476);
nor U23799 (N_23799,N_17884,N_18539);
and U23800 (N_23800,N_11214,N_13461);
or U23801 (N_23801,N_10483,N_10412);
xor U23802 (N_23802,N_11621,N_16806);
nor U23803 (N_23803,N_18544,N_12304);
nand U23804 (N_23804,N_13783,N_11353);
nand U23805 (N_23805,N_19480,N_18583);
xor U23806 (N_23806,N_17558,N_14372);
xor U23807 (N_23807,N_19803,N_11314);
and U23808 (N_23808,N_12012,N_12171);
xor U23809 (N_23809,N_11819,N_13577);
nor U23810 (N_23810,N_10049,N_12113);
and U23811 (N_23811,N_16352,N_13151);
or U23812 (N_23812,N_10399,N_13240);
nor U23813 (N_23813,N_10671,N_16701);
xor U23814 (N_23814,N_11769,N_12588);
nand U23815 (N_23815,N_11743,N_15055);
and U23816 (N_23816,N_19379,N_13496);
xnor U23817 (N_23817,N_13255,N_10273);
and U23818 (N_23818,N_14455,N_12460);
nor U23819 (N_23819,N_12873,N_15865);
nand U23820 (N_23820,N_17121,N_19873);
or U23821 (N_23821,N_18942,N_10127);
or U23822 (N_23822,N_13579,N_18713);
and U23823 (N_23823,N_18580,N_13681);
or U23824 (N_23824,N_15135,N_15363);
or U23825 (N_23825,N_19308,N_17248);
xor U23826 (N_23826,N_13239,N_11305);
nor U23827 (N_23827,N_19222,N_17789);
and U23828 (N_23828,N_12111,N_12930);
xnor U23829 (N_23829,N_19931,N_13993);
nand U23830 (N_23830,N_19676,N_15203);
or U23831 (N_23831,N_11386,N_16670);
or U23832 (N_23832,N_14568,N_12843);
nand U23833 (N_23833,N_14460,N_18080);
nor U23834 (N_23834,N_11615,N_15613);
nor U23835 (N_23835,N_18738,N_19751);
xor U23836 (N_23836,N_13023,N_17107);
nand U23837 (N_23837,N_13869,N_15494);
xor U23838 (N_23838,N_15261,N_11540);
nand U23839 (N_23839,N_16835,N_10627);
xnor U23840 (N_23840,N_14912,N_18590);
nor U23841 (N_23841,N_13222,N_16545);
nand U23842 (N_23842,N_16375,N_15632);
nand U23843 (N_23843,N_19645,N_13355);
and U23844 (N_23844,N_18211,N_17702);
nor U23845 (N_23845,N_16465,N_12437);
nor U23846 (N_23846,N_13487,N_10626);
and U23847 (N_23847,N_13092,N_15776);
xnor U23848 (N_23848,N_12603,N_11395);
and U23849 (N_23849,N_12560,N_14360);
or U23850 (N_23850,N_14410,N_17131);
nor U23851 (N_23851,N_15473,N_10151);
nor U23852 (N_23852,N_19233,N_18603);
nand U23853 (N_23853,N_10562,N_13102);
nand U23854 (N_23854,N_12199,N_14334);
or U23855 (N_23855,N_15102,N_16401);
or U23856 (N_23856,N_18120,N_19810);
and U23857 (N_23857,N_19855,N_16732);
nand U23858 (N_23858,N_17364,N_19642);
nor U23859 (N_23859,N_12298,N_10357);
or U23860 (N_23860,N_18108,N_16598);
xor U23861 (N_23861,N_13291,N_18212);
and U23862 (N_23862,N_13548,N_13019);
nand U23863 (N_23863,N_12196,N_14689);
nor U23864 (N_23864,N_12186,N_10967);
xor U23865 (N_23865,N_12820,N_19765);
nand U23866 (N_23866,N_12060,N_19402);
nand U23867 (N_23867,N_14906,N_11033);
or U23868 (N_23868,N_18046,N_19661);
nand U23869 (N_23869,N_17480,N_15692);
xor U23870 (N_23870,N_15392,N_18691);
nand U23871 (N_23871,N_15158,N_16563);
or U23872 (N_23872,N_18937,N_18925);
nor U23873 (N_23873,N_11341,N_16638);
or U23874 (N_23874,N_13261,N_19965);
xnor U23875 (N_23875,N_15374,N_13505);
xor U23876 (N_23876,N_14821,N_17391);
xnor U23877 (N_23877,N_15224,N_17778);
nor U23878 (N_23878,N_16805,N_19151);
xnor U23879 (N_23879,N_19618,N_12468);
and U23880 (N_23880,N_15993,N_11895);
or U23881 (N_23881,N_18201,N_10745);
nand U23882 (N_23882,N_12341,N_14138);
nor U23883 (N_23883,N_10541,N_12253);
xnor U23884 (N_23884,N_11091,N_13830);
xor U23885 (N_23885,N_18102,N_15015);
nor U23886 (N_23886,N_15072,N_13033);
nor U23887 (N_23887,N_18064,N_11008);
nor U23888 (N_23888,N_19942,N_17783);
and U23889 (N_23889,N_15789,N_12732);
and U23890 (N_23890,N_14561,N_15322);
nor U23891 (N_23891,N_11234,N_19006);
and U23892 (N_23892,N_13649,N_11279);
nand U23893 (N_23893,N_13540,N_19184);
nor U23894 (N_23894,N_18057,N_15608);
nor U23895 (N_23895,N_18239,N_15916);
nor U23896 (N_23896,N_10415,N_12436);
or U23897 (N_23897,N_12165,N_16205);
and U23898 (N_23898,N_15745,N_14982);
nand U23899 (N_23899,N_10431,N_17291);
and U23900 (N_23900,N_11364,N_15192);
and U23901 (N_23901,N_10762,N_12860);
and U23902 (N_23902,N_19478,N_11437);
nor U23903 (N_23903,N_14642,N_11933);
or U23904 (N_23904,N_18292,N_14788);
nand U23905 (N_23905,N_12764,N_11046);
xnor U23906 (N_23906,N_15367,N_15181);
or U23907 (N_23907,N_13839,N_10029);
nand U23908 (N_23908,N_15920,N_11770);
xnor U23909 (N_23909,N_11834,N_18840);
and U23910 (N_23910,N_18027,N_16084);
and U23911 (N_23911,N_18968,N_18605);
and U23912 (N_23912,N_13753,N_17870);
and U23913 (N_23913,N_10842,N_13139);
nor U23914 (N_23914,N_17765,N_10781);
and U23915 (N_23915,N_10625,N_14258);
or U23916 (N_23916,N_11423,N_12363);
nor U23917 (N_23917,N_15206,N_10857);
nor U23918 (N_23918,N_15169,N_10864);
and U23919 (N_23919,N_15468,N_17218);
or U23920 (N_23920,N_11023,N_16514);
or U23921 (N_23921,N_13079,N_11856);
nor U23922 (N_23922,N_17285,N_15888);
nor U23923 (N_23923,N_17215,N_19615);
and U23924 (N_23924,N_16848,N_12583);
or U23925 (N_23925,N_17568,N_17518);
nand U23926 (N_23926,N_16675,N_16819);
xnor U23927 (N_23927,N_10070,N_11539);
or U23928 (N_23928,N_13336,N_13848);
and U23929 (N_23929,N_16761,N_11914);
and U23930 (N_23930,N_12923,N_18104);
or U23931 (N_23931,N_10725,N_14021);
nor U23932 (N_23932,N_13764,N_15384);
or U23933 (N_23933,N_13417,N_10830);
and U23934 (N_23934,N_15575,N_17205);
and U23935 (N_23935,N_16599,N_17773);
nand U23936 (N_23936,N_11156,N_13455);
and U23937 (N_23937,N_10264,N_13876);
nor U23938 (N_23938,N_12919,N_17301);
xnor U23939 (N_23939,N_19899,N_11094);
and U23940 (N_23940,N_11801,N_10682);
nor U23941 (N_23941,N_16778,N_13838);
or U23942 (N_23942,N_12522,N_19816);
or U23943 (N_23943,N_16998,N_12022);
nand U23944 (N_23944,N_10074,N_14903);
nor U23945 (N_23945,N_10611,N_14577);
xor U23946 (N_23946,N_11951,N_15570);
nor U23947 (N_23947,N_14652,N_19202);
nand U23948 (N_23948,N_18496,N_11803);
nand U23949 (N_23949,N_19995,N_19323);
and U23950 (N_23950,N_14066,N_15354);
nor U23951 (N_23951,N_18310,N_10807);
xor U23952 (N_23952,N_10396,N_12865);
xnor U23953 (N_23953,N_11001,N_14070);
and U23954 (N_23954,N_10794,N_18901);
xnor U23955 (N_23955,N_14676,N_14895);
nand U23956 (N_23956,N_12045,N_17831);
xor U23957 (N_23957,N_17080,N_11405);
and U23958 (N_23958,N_14406,N_14140);
xnor U23959 (N_23959,N_17072,N_12869);
xor U23960 (N_23960,N_15681,N_15586);
xor U23961 (N_23961,N_14829,N_15965);
and U23962 (N_23962,N_10325,N_18049);
and U23963 (N_23963,N_17542,N_16456);
and U23964 (N_23964,N_16870,N_15099);
or U23965 (N_23965,N_13742,N_18698);
or U23966 (N_23966,N_14708,N_12729);
nand U23967 (N_23967,N_13891,N_14700);
xnor U23968 (N_23968,N_10536,N_17151);
and U23969 (N_23969,N_13169,N_11647);
and U23970 (N_23970,N_11253,N_12392);
nand U23971 (N_23971,N_10067,N_12348);
nand U23972 (N_23972,N_11906,N_14434);
xor U23973 (N_23973,N_13819,N_13029);
or U23974 (N_23974,N_12769,N_13339);
and U23975 (N_23975,N_11185,N_15307);
xnor U23976 (N_23976,N_10492,N_17401);
nand U23977 (N_23977,N_17367,N_16136);
nand U23978 (N_23978,N_13189,N_16530);
nand U23979 (N_23979,N_16809,N_12537);
nand U23980 (N_23980,N_13571,N_18191);
xor U23981 (N_23981,N_10453,N_11282);
nor U23982 (N_23982,N_12411,N_12589);
xnor U23983 (N_23983,N_10903,N_10201);
xnor U23984 (N_23984,N_16975,N_13123);
xor U23985 (N_23985,N_15360,N_16972);
nor U23986 (N_23986,N_16065,N_11516);
xnor U23987 (N_23987,N_14684,N_11037);
or U23988 (N_23988,N_17543,N_14183);
xor U23989 (N_23989,N_10686,N_18304);
or U23990 (N_23990,N_11381,N_14880);
xnor U23991 (N_23991,N_18152,N_12250);
xor U23992 (N_23992,N_15065,N_16463);
nand U23993 (N_23993,N_10978,N_11744);
xnor U23994 (N_23994,N_12948,N_15283);
and U23995 (N_23995,N_17986,N_10516);
or U23996 (N_23996,N_11351,N_17068);
xnor U23997 (N_23997,N_15893,N_12328);
nor U23998 (N_23998,N_17312,N_15033);
and U23999 (N_23999,N_12529,N_12481);
or U24000 (N_24000,N_10179,N_17662);
nand U24001 (N_24001,N_12419,N_12660);
xnor U24002 (N_24002,N_18702,N_10730);
nand U24003 (N_24003,N_10588,N_18398);
or U24004 (N_24004,N_18912,N_11922);
xnor U24005 (N_24005,N_17011,N_16865);
nor U24006 (N_24006,N_12531,N_11376);
nor U24007 (N_24007,N_12718,N_14920);
or U24008 (N_24008,N_15735,N_12482);
nor U24009 (N_24009,N_14317,N_19608);
xnor U24010 (N_24010,N_18936,N_16548);
nand U24011 (N_24011,N_13145,N_16954);
xnor U24012 (N_24012,N_13206,N_18433);
xor U24013 (N_24013,N_16275,N_19257);
nand U24014 (N_24014,N_15196,N_17224);
xor U24015 (N_24015,N_15340,N_15139);
or U24016 (N_24016,N_18555,N_16706);
xnor U24017 (N_24017,N_12404,N_13479);
nor U24018 (N_24018,N_10828,N_16627);
nand U24019 (N_24019,N_18625,N_11321);
xor U24020 (N_24020,N_12274,N_18061);
or U24021 (N_24021,N_15028,N_13318);
nor U24022 (N_24022,N_14453,N_16934);
nor U24023 (N_24023,N_10567,N_17877);
and U24024 (N_24024,N_17222,N_17108);
xor U24025 (N_24025,N_16344,N_19924);
xor U24026 (N_24026,N_19804,N_14350);
nor U24027 (N_24027,N_13678,N_17277);
or U24028 (N_24028,N_17150,N_13617);
or U24029 (N_24029,N_15184,N_18838);
nor U24030 (N_24030,N_19604,N_13952);
and U24031 (N_24031,N_17948,N_11355);
nand U24032 (N_24032,N_14167,N_13555);
and U24033 (N_24033,N_10540,N_15827);
and U24034 (N_24034,N_14423,N_17647);
nand U24035 (N_24035,N_15908,N_16996);
nand U24036 (N_24036,N_15734,N_14126);
nor U24037 (N_24037,N_15088,N_14116);
nand U24038 (N_24038,N_11295,N_13778);
nor U24039 (N_24039,N_18871,N_15923);
nor U24040 (N_24040,N_16845,N_18636);
or U24041 (N_24041,N_18497,N_18071);
nand U24042 (N_24042,N_11425,N_12686);
and U24043 (N_24043,N_11207,N_19008);
and U24044 (N_24044,N_17176,N_14016);
nand U24045 (N_24045,N_17117,N_12387);
and U24046 (N_24046,N_11272,N_10700);
nor U24047 (N_24047,N_13923,N_12218);
nor U24048 (N_24048,N_15045,N_19436);
nand U24049 (N_24049,N_13122,N_18339);
or U24050 (N_24050,N_15512,N_17442);
and U24051 (N_24051,N_19196,N_13462);
nor U24052 (N_24052,N_19556,N_17163);
nand U24053 (N_24053,N_13030,N_16438);
nand U24054 (N_24054,N_12594,N_16658);
xnor U24055 (N_24055,N_11772,N_12366);
xor U24056 (N_24056,N_18215,N_10050);
or U24057 (N_24057,N_14039,N_11055);
xnor U24058 (N_24058,N_16371,N_11600);
and U24059 (N_24059,N_10417,N_16363);
nand U24060 (N_24060,N_14830,N_17744);
nand U24061 (N_24061,N_14548,N_16254);
and U24062 (N_24062,N_12247,N_10421);
or U24063 (N_24063,N_12081,N_16219);
and U24064 (N_24064,N_15385,N_15551);
or U24065 (N_24065,N_14748,N_12214);
nor U24066 (N_24066,N_17553,N_11764);
or U24067 (N_24067,N_17251,N_13320);
nor U24068 (N_24068,N_12439,N_17017);
and U24069 (N_24069,N_19090,N_14824);
nand U24070 (N_24070,N_12980,N_17929);
nand U24071 (N_24071,N_14591,N_12899);
xnor U24072 (N_24072,N_16847,N_14671);
and U24073 (N_24073,N_10633,N_14492);
or U24074 (N_24074,N_17237,N_14832);
nand U24075 (N_24075,N_18089,N_15448);
or U24076 (N_24076,N_13866,N_18070);
and U24077 (N_24077,N_14826,N_17813);
and U24078 (N_24078,N_16461,N_18913);
or U24079 (N_24079,N_19814,N_13958);
xnor U24080 (N_24080,N_10166,N_18279);
or U24081 (N_24081,N_18811,N_10005);
nand U24082 (N_24082,N_17439,N_10458);
nor U24083 (N_24083,N_16760,N_13138);
and U24084 (N_24084,N_12549,N_18689);
and U24085 (N_24085,N_15577,N_18648);
xnor U24086 (N_24086,N_17326,N_13087);
nand U24087 (N_24087,N_11485,N_18309);
xor U24088 (N_24088,N_13600,N_17178);
nand U24089 (N_24089,N_15434,N_13580);
nor U24090 (N_24090,N_13393,N_12467);
nor U24091 (N_24091,N_15946,N_12671);
or U24092 (N_24092,N_11244,N_15620);
or U24093 (N_24093,N_13309,N_15418);
and U24094 (N_24094,N_19712,N_14644);
nor U24095 (N_24095,N_12189,N_13175);
nor U24096 (N_24096,N_10232,N_13331);
or U24097 (N_24097,N_14154,N_11715);
or U24098 (N_24098,N_18315,N_11394);
nand U24099 (N_24099,N_18267,N_12694);
nor U24100 (N_24100,N_14633,N_19695);
nand U24101 (N_24101,N_14079,N_12803);
nand U24102 (N_24102,N_18819,N_14900);
nor U24103 (N_24103,N_14194,N_18415);
nor U24104 (N_24104,N_11817,N_16117);
and U24105 (N_24105,N_19109,N_14871);
or U24106 (N_24106,N_11958,N_13938);
xor U24107 (N_24107,N_13539,N_16245);
nor U24108 (N_24108,N_11442,N_15191);
or U24109 (N_24109,N_14093,N_12561);
and U24110 (N_24110,N_15489,N_16662);
nor U24111 (N_24111,N_16336,N_19948);
nand U24112 (N_24112,N_11075,N_10608);
or U24113 (N_24113,N_13295,N_18450);
or U24114 (N_24114,N_18368,N_17303);
or U24115 (N_24115,N_17413,N_15869);
or U24116 (N_24116,N_16989,N_19708);
xor U24117 (N_24117,N_19698,N_11982);
xor U24118 (N_24118,N_19174,N_10170);
nor U24119 (N_24119,N_12382,N_13987);
or U24120 (N_24120,N_16116,N_11385);
or U24121 (N_24121,N_13321,N_18347);
or U24122 (N_24122,N_10749,N_11157);
and U24123 (N_24123,N_14662,N_18241);
or U24124 (N_24124,N_16906,N_14610);
nor U24125 (N_24125,N_14171,N_10513);
nor U24126 (N_24126,N_10764,N_12322);
and U24127 (N_24127,N_14441,N_15440);
nand U24128 (N_24128,N_16590,N_10342);
xnor U24129 (N_24129,N_19310,N_10076);
nand U24130 (N_24130,N_11339,N_19322);
nor U24131 (N_24131,N_17828,N_12369);
nand U24132 (N_24132,N_17968,N_10135);
and U24133 (N_24133,N_11956,N_12829);
or U24134 (N_24134,N_10490,N_15435);
nand U24135 (N_24135,N_18154,N_18653);
nand U24136 (N_24136,N_12878,N_15475);
xnor U24137 (N_24137,N_11586,N_15144);
nand U24138 (N_24138,N_15396,N_13978);
xnor U24139 (N_24139,N_12934,N_19927);
nand U24140 (N_24140,N_12473,N_17683);
nor U24141 (N_24141,N_14675,N_15981);
and U24142 (N_24142,N_16138,N_17319);
xnor U24143 (N_24143,N_12961,N_18780);
nor U24144 (N_24144,N_10196,N_18560);
and U24145 (N_24145,N_13088,N_16262);
and U24146 (N_24146,N_16552,N_18898);
and U24147 (N_24147,N_19088,N_10395);
and U24148 (N_24148,N_17894,N_12725);
nand U24149 (N_24149,N_10272,N_12127);
and U24150 (N_24150,N_14686,N_11410);
and U24151 (N_24151,N_15817,N_12532);
and U24152 (N_24152,N_18589,N_14467);
and U24153 (N_24153,N_16353,N_10337);
nand U24154 (N_24154,N_17426,N_10443);
or U24155 (N_24155,N_11209,N_17507);
xnor U24156 (N_24156,N_15127,N_15248);
nor U24157 (N_24157,N_17202,N_18276);
or U24158 (N_24158,N_10034,N_12333);
nand U24159 (N_24159,N_18607,N_17664);
or U24160 (N_24160,N_11306,N_17058);
xor U24161 (N_24161,N_17083,N_16872);
nand U24162 (N_24162,N_10792,N_16650);
and U24163 (N_24163,N_13032,N_10583);
nand U24164 (N_24164,N_12959,N_15922);
xnor U24165 (N_24165,N_16896,N_11139);
and U24166 (N_24166,N_10134,N_15022);
nand U24167 (N_24167,N_15238,N_19388);
nand U24168 (N_24168,N_15081,N_11747);
nand U24169 (N_24169,N_14799,N_16931);
xnor U24170 (N_24170,N_18478,N_14170);
or U24171 (N_24171,N_13834,N_16997);
nor U24172 (N_24172,N_16417,N_14963);
nor U24173 (N_24173,N_15255,N_19709);
nor U24174 (N_24174,N_12405,N_13607);
or U24175 (N_24175,N_13359,N_11488);
and U24176 (N_24176,N_12649,N_19619);
or U24177 (N_24177,N_18288,N_19267);
nand U24178 (N_24178,N_16118,N_13691);
xnor U24179 (N_24179,N_10021,N_19541);
and U24180 (N_24180,N_10040,N_12063);
nand U24181 (N_24181,N_17882,N_14169);
nand U24182 (N_24182,N_11908,N_14289);
nor U24183 (N_24183,N_18787,N_12374);
or U24184 (N_24184,N_19453,N_11081);
xnor U24185 (N_24185,N_18620,N_18044);
and U24186 (N_24186,N_19935,N_16620);
and U24187 (N_24187,N_19776,N_18167);
or U24188 (N_24188,N_16687,N_10800);
and U24189 (N_24189,N_17519,N_17349);
or U24190 (N_24190,N_15898,N_10299);
xnor U24191 (N_24191,N_11316,N_14966);
nor U24192 (N_24192,N_18695,N_15324);
nor U24193 (N_24193,N_11931,N_10824);
or U24194 (N_24194,N_19524,N_15509);
nor U24195 (N_24195,N_18875,N_12176);
or U24196 (N_24196,N_17759,N_10158);
and U24197 (N_24197,N_18674,N_12398);
and U24198 (N_24198,N_18591,N_17161);
nor U24199 (N_24199,N_18914,N_13308);
and U24200 (N_24200,N_17673,N_16569);
or U24201 (N_24201,N_19061,N_11642);
and U24202 (N_24202,N_10507,N_12249);
nor U24203 (N_24203,N_10447,N_11616);
xor U24204 (N_24204,N_19105,N_19119);
and U24205 (N_24205,N_17225,N_12712);
or U24206 (N_24206,N_16833,N_11424);
or U24207 (N_24207,N_19974,N_10710);
xor U24208 (N_24208,N_19734,N_13672);
xnor U24209 (N_24209,N_11941,N_19918);
and U24210 (N_24210,N_12633,N_18849);
nand U24211 (N_24211,N_13131,N_16094);
or U24212 (N_24212,N_19559,N_12508);
nand U24213 (N_24213,N_18228,N_18551);
nor U24214 (N_24214,N_19087,N_11779);
nand U24215 (N_24215,N_14468,N_11862);
xor U24216 (N_24216,N_14411,N_14526);
xnor U24217 (N_24217,N_17409,N_10102);
or U24218 (N_24218,N_13859,N_15520);
nor U24219 (N_24219,N_17383,N_19492);
nor U24220 (N_24220,N_10934,N_12602);
or U24221 (N_24221,N_13944,N_10446);
nand U24222 (N_24222,N_11623,N_14031);
nor U24223 (N_24223,N_13610,N_19292);
nor U24224 (N_24224,N_10988,N_13322);
nand U24225 (N_24225,N_17216,N_17597);
and U24226 (N_24226,N_14279,N_19944);
xnor U24227 (N_24227,N_17501,N_17995);
and U24228 (N_24228,N_10790,N_19049);
and U24229 (N_24229,N_18312,N_11521);
nand U24230 (N_24230,N_12881,N_16790);
nor U24231 (N_24231,N_14396,N_15881);
and U24232 (N_24232,N_16169,N_12714);
or U24233 (N_24233,N_18768,N_19881);
or U24234 (N_24234,N_18791,N_14924);
and U24235 (N_24235,N_13702,N_19459);
nor U24236 (N_24236,N_13504,N_10546);
xor U24237 (N_24237,N_19053,N_11471);
and U24238 (N_24238,N_14507,N_17552);
nand U24239 (N_24239,N_17408,N_18329);
or U24240 (N_24240,N_13535,N_19578);
nand U24241 (N_24241,N_13851,N_11438);
and U24242 (N_24242,N_10084,N_12789);
or U24243 (N_24243,N_17625,N_19583);
and U24244 (N_24244,N_14325,N_16333);
nor U24245 (N_24245,N_14368,N_19307);
nor U24246 (N_24246,N_17412,N_10714);
nand U24247 (N_24247,N_16145,N_13616);
nor U24248 (N_24248,N_12336,N_17582);
nand U24249 (N_24249,N_18051,N_10146);
nand U24250 (N_24250,N_12331,N_17846);
nand U24251 (N_24251,N_19646,N_13559);
xnor U24252 (N_24252,N_14343,N_10928);
or U24253 (N_24253,N_10663,N_10769);
nor U24254 (N_24254,N_10922,N_12360);
nor U24255 (N_24255,N_11798,N_11599);
and U24256 (N_24256,N_11434,N_10263);
or U24257 (N_24257,N_10708,N_12400);
and U24258 (N_24258,N_10343,N_11195);
xor U24259 (N_24259,N_16360,N_10673);
or U24260 (N_24260,N_19844,N_11955);
or U24261 (N_24261,N_16029,N_14179);
nand U24262 (N_24262,N_11871,N_16651);
xnor U24263 (N_24263,N_12184,N_11888);
or U24264 (N_24264,N_11936,N_10462);
and U24265 (N_24265,N_15391,N_17728);
nor U24266 (N_24266,N_13444,N_15056);
or U24267 (N_24267,N_11686,N_11915);
nor U24268 (N_24268,N_14489,N_19553);
and U24269 (N_24269,N_15818,N_13258);
nand U24270 (N_24270,N_14339,N_17611);
nor U24271 (N_24271,N_18717,N_15580);
and U24272 (N_24272,N_15017,N_13899);
nand U24273 (N_24273,N_12530,N_16097);
nor U24274 (N_24274,N_12776,N_16744);
nand U24275 (N_24275,N_12233,N_16892);
nand U24276 (N_24276,N_12151,N_13965);
xor U24277 (N_24277,N_11742,N_15630);
or U24278 (N_24278,N_17969,N_19644);
or U24279 (N_24279,N_12891,N_19548);
and U24280 (N_24280,N_10498,N_19843);
nand U24281 (N_24281,N_16541,N_18537);
or U24282 (N_24282,N_13512,N_14516);
nand U24283 (N_24283,N_11439,N_10315);
or U24284 (N_24284,N_10144,N_11014);
xor U24285 (N_24285,N_11382,N_13880);
nand U24286 (N_24286,N_13912,N_19864);
or U24287 (N_24287,N_13727,N_11917);
and U24288 (N_24288,N_14759,N_11846);
xnor U24289 (N_24289,N_16783,N_18534);
nand U24290 (N_24290,N_13786,N_10344);
or U24291 (N_24291,N_11667,N_18232);
nor U24292 (N_24292,N_15822,N_16180);
xnor U24293 (N_24293,N_19914,N_10882);
nor U24294 (N_24294,N_14831,N_19429);
xnor U24295 (N_24295,N_16370,N_18536);
or U24296 (N_24296,N_19046,N_12827);
nand U24297 (N_24297,N_19789,N_18081);
and U24298 (N_24298,N_17940,N_15460);
or U24299 (N_24299,N_13601,N_11943);
nor U24300 (N_24300,N_10892,N_16503);
xnor U24301 (N_24301,N_17475,N_15722);
nor U24302 (N_24302,N_10148,N_18021);
and U24303 (N_24303,N_12747,N_13881);
nor U24304 (N_24304,N_13547,N_15071);
nand U24305 (N_24305,N_16010,N_13340);
nor U24306 (N_24306,N_18816,N_17811);
xnor U24307 (N_24307,N_14510,N_11464);
xnor U24308 (N_24308,N_17978,N_18866);
nor U24309 (N_24309,N_18011,N_16049);
and U24310 (N_24310,N_18463,N_15263);
xnor U24311 (N_24311,N_12990,N_10086);
nand U24312 (N_24312,N_14221,N_18706);
nor U24313 (N_24313,N_18195,N_14095);
and U24314 (N_24314,N_18669,N_11698);
nand U24315 (N_24315,N_13481,N_18390);
and U24316 (N_24316,N_12997,N_12232);
or U24317 (N_24317,N_16059,N_16648);
nand U24318 (N_24318,N_11820,N_19134);
xor U24319 (N_24319,N_12323,N_11664);
or U24320 (N_24320,N_12225,N_10059);
xnor U24321 (N_24321,N_11603,N_16915);
nor U24322 (N_24322,N_10191,N_16078);
nand U24323 (N_24323,N_11130,N_13609);
or U24324 (N_24324,N_13238,N_18815);
nand U24325 (N_24325,N_11528,N_12533);
and U24326 (N_24326,N_10474,N_10727);
and U24327 (N_24327,N_10832,N_10456);
xnor U24328 (N_24328,N_16027,N_17090);
and U24329 (N_24329,N_13028,N_16587);
nor U24330 (N_24330,N_18725,N_11806);
or U24331 (N_24331,N_14544,N_10183);
nand U24332 (N_24332,N_15871,N_15319);
and U24333 (N_24333,N_12068,N_19133);
xnor U24334 (N_24334,N_13374,N_12449);
and U24335 (N_24335,N_15477,N_10202);
nor U24336 (N_24336,N_11512,N_14502);
nand U24337 (N_24337,N_13777,N_13629);
xor U24338 (N_24338,N_15287,N_12739);
nand U24339 (N_24339,N_19747,N_11966);
xor U24340 (N_24340,N_16223,N_10106);
nor U24341 (N_24341,N_17822,N_18332);
nand U24342 (N_24342,N_12354,N_10279);
xor U24343 (N_24343,N_16295,N_10984);
and U24344 (N_24344,N_16922,N_19369);
xnor U24345 (N_24345,N_19142,N_15519);
xnor U24346 (N_24346,N_12996,N_17145);
nor U24347 (N_24347,N_12883,N_13027);
or U24348 (N_24348,N_19679,N_10186);
nand U24349 (N_24349,N_14165,N_15043);
and U24350 (N_24350,N_13003,N_14361);
xor U24351 (N_24351,N_16853,N_18085);
xor U24352 (N_24352,N_10966,N_10899);
xor U24353 (N_24353,N_19579,N_18934);
xor U24354 (N_24354,N_11964,N_13633);
nand U24355 (N_24355,N_14631,N_13171);
xnor U24356 (N_24356,N_13904,N_16862);
nor U24357 (N_24357,N_13083,N_17235);
and U24358 (N_24358,N_17950,N_17435);
and U24359 (N_24359,N_11669,N_10793);
xor U24360 (N_24360,N_17082,N_14535);
nand U24361 (N_24361,N_17477,N_19820);
and U24362 (N_24362,N_19013,N_11401);
nor U24363 (N_24363,N_13451,N_13995);
nor U24364 (N_24364,N_13274,N_10256);
and U24365 (N_24365,N_16234,N_18077);
or U24366 (N_24366,N_14333,N_13808);
nor U24367 (N_24367,N_12981,N_19243);
nor U24368 (N_24368,N_11967,N_16122);
xnor U24369 (N_24369,N_16990,N_10587);
nand U24370 (N_24370,N_15515,N_11021);
and U24371 (N_24371,N_13901,N_17504);
xnor U24372 (N_24372,N_19255,N_19802);
and U24373 (N_24373,N_17476,N_17682);
nand U24374 (N_24374,N_16881,N_19420);
nor U24375 (N_24375,N_18336,N_15318);
nand U24376 (N_24376,N_18571,N_10353);
and U24377 (N_24377,N_15424,N_17990);
nor U24378 (N_24378,N_17270,N_18957);
nand U24379 (N_24379,N_15133,N_11002);
xnor U24380 (N_24380,N_17081,N_11794);
nand U24381 (N_24381,N_13313,N_19762);
xnor U24382 (N_24382,N_13795,N_14850);
and U24383 (N_24383,N_18938,N_17588);
and U24384 (N_24384,N_18236,N_10811);
and U24385 (N_24385,N_13516,N_11063);
nand U24386 (N_24386,N_11050,N_14606);
and U24387 (N_24387,N_16317,N_11776);
nand U24388 (N_24388,N_10520,N_13525);
nor U24389 (N_24389,N_13195,N_16733);
nand U24390 (N_24390,N_16821,N_13746);
nor U24391 (N_24391,N_14607,N_10245);
nand U24392 (N_24392,N_15762,N_15352);
nand U24393 (N_24393,N_14949,N_19340);
nand U24394 (N_24394,N_18792,N_14429);
xor U24395 (N_24395,N_19367,N_10652);
nand U24396 (N_24396,N_15154,N_17745);
xor U24397 (N_24397,N_16758,N_12477);
nor U24398 (N_24398,N_18926,N_15220);
and U24399 (N_24399,N_18637,N_14970);
xnor U24400 (N_24400,N_12757,N_15378);
nand U24401 (N_24401,N_10763,N_15485);
or U24402 (N_24402,N_19761,N_15292);
xnor U24403 (N_24403,N_10449,N_17031);
xnor U24404 (N_24404,N_14608,N_15492);
nor U24405 (N_24405,N_19968,N_12717);
and U24406 (N_24406,N_16312,N_15001);
nor U24407 (N_24407,N_16876,N_15172);
nor U24408 (N_24408,N_15636,N_11554);
or U24409 (N_24409,N_12826,N_16087);
xnor U24410 (N_24410,N_13814,N_14961);
nor U24411 (N_24411,N_14582,N_10323);
nand U24412 (N_24412,N_17450,N_12431);
xnor U24413 (N_24413,N_10657,N_13373);
nand U24414 (N_24414,N_11685,N_14100);
xor U24415 (N_24415,N_19448,N_12870);
nand U24416 (N_24416,N_14650,N_14716);
xnor U24417 (N_24417,N_14739,N_15235);
nor U24418 (N_24418,N_11297,N_10367);
and U24419 (N_24419,N_10683,N_14139);
or U24420 (N_24420,N_11429,N_17293);
or U24421 (N_24421,N_10275,N_14596);
xnor U24422 (N_24422,N_14658,N_14008);
nor U24423 (N_24423,N_19440,N_15270);
nand U24424 (N_24424,N_13101,N_11128);
nor U24425 (N_24425,N_19737,N_14760);
or U24426 (N_24426,N_11174,N_11336);
xor U24427 (N_24427,N_10031,N_13493);
and U24428 (N_24428,N_17351,N_18393);
nand U24429 (N_24429,N_14956,N_19387);
and U24430 (N_24430,N_17838,N_13801);
or U24431 (N_24431,N_10645,N_13697);
nor U24432 (N_24432,N_15610,N_15046);
xor U24433 (N_24433,N_13828,N_19754);
nor U24434 (N_24434,N_16739,N_17955);
nor U24435 (N_24435,N_16624,N_13143);
nor U24436 (N_24436,N_15664,N_18127);
or U24437 (N_24437,N_19699,N_14063);
xnor U24438 (N_24438,N_13689,N_15508);
nor U24439 (N_24439,N_17738,N_19177);
and U24440 (N_24440,N_15840,N_19859);
nor U24441 (N_24441,N_10188,N_19110);
nand U24442 (N_24442,N_12760,N_18153);
nand U24443 (N_24443,N_12372,N_17452);
nand U24444 (N_24444,N_16050,N_13526);
nand U24445 (N_24445,N_17028,N_10722);
xnor U24446 (N_24446,N_19674,N_11949);
xnor U24447 (N_24447,N_18502,N_11268);
nor U24448 (N_24448,N_16617,N_10759);
or U24449 (N_24449,N_14622,N_19564);
or U24450 (N_24450,N_17720,N_17505);
or U24451 (N_24451,N_11448,N_11273);
nand U24452 (N_24452,N_15719,N_13482);
nand U24453 (N_24453,N_11220,N_17808);
nand U24454 (N_24454,N_10505,N_13073);
or U24455 (N_24455,N_14511,N_11893);
nor U24456 (N_24456,N_16429,N_16550);
nand U24457 (N_24457,N_11699,N_18828);
and U24458 (N_24458,N_14769,N_17736);
and U24459 (N_24459,N_14401,N_16525);
and U24460 (N_24460,N_12066,N_17165);
nand U24461 (N_24461,N_19306,N_10500);
or U24462 (N_24462,N_11588,N_16481);
or U24463 (N_24463,N_10237,N_11726);
xnor U24464 (N_24464,N_14491,N_15754);
nand U24465 (N_24465,N_10582,N_16338);
or U24466 (N_24466,N_13903,N_14099);
nor U24467 (N_24467,N_15583,N_15820);
and U24468 (N_24468,N_18207,N_16420);
xor U24469 (N_24469,N_12401,N_17975);
or U24470 (N_24470,N_12507,N_11934);
or U24471 (N_24471,N_18052,N_10897);
nor U24472 (N_24472,N_12093,N_12037);
xnor U24473 (N_24473,N_14178,N_11592);
or U24474 (N_24474,N_19217,N_13705);
nand U24475 (N_24475,N_12272,N_17824);
and U24476 (N_24476,N_19264,N_17937);
nand U24477 (N_24477,N_19462,N_15291);
xor U24478 (N_24478,N_18144,N_13736);
and U24479 (N_24479,N_14180,N_19627);
nor U24480 (N_24480,N_15901,N_14761);
nor U24481 (N_24481,N_19069,N_10020);
and U24482 (N_24482,N_18986,N_15715);
or U24483 (N_24483,N_16452,N_18905);
and U24484 (N_24484,N_12280,N_11451);
and U24485 (N_24485,N_16387,N_11924);
or U24486 (N_24486,N_13747,N_13290);
nand U24487 (N_24487,N_12969,N_11885);
nand U24488 (N_24488,N_11808,N_16236);
and U24489 (N_24489,N_18801,N_15333);
nand U24490 (N_24490,N_18509,N_10748);
or U24491 (N_24491,N_12770,N_19994);
or U24492 (N_24492,N_16062,N_14833);
or U24493 (N_24493,N_16142,N_10199);
xnor U24494 (N_24494,N_13344,N_10847);
nor U24495 (N_24495,N_19294,N_16505);
and U24496 (N_24496,N_17703,N_12142);
xnor U24497 (N_24497,N_15039,N_19356);
xor U24498 (N_24498,N_10973,N_18065);
or U24499 (N_24499,N_19668,N_17524);
nand U24500 (N_24500,N_11168,N_17747);
nand U24501 (N_24501,N_15421,N_19103);
nor U24502 (N_24502,N_13024,N_15051);
nor U24503 (N_24503,N_19287,N_16641);
nor U24504 (N_24504,N_13902,N_17545);
xnor U24505 (N_24505,N_19438,N_15979);
nor U24506 (N_24506,N_18910,N_13743);
nand U24507 (N_24507,N_11710,N_14602);
or U24508 (N_24508,N_14323,N_19408);
nand U24509 (N_24509,N_15609,N_10569);
xor U24510 (N_24510,N_19383,N_10198);
and U24511 (N_24511,N_19910,N_14965);
and U24512 (N_24512,N_18621,N_12039);
nand U24513 (N_24513,N_11695,N_19664);
nor U24514 (N_24514,N_14369,N_13569);
and U24515 (N_24515,N_14754,N_14146);
and U24516 (N_24516,N_19720,N_14661);
nor U24517 (N_24517,N_15917,N_15944);
and U24518 (N_24518,N_11930,N_17469);
xnor U24519 (N_24519,N_15183,N_16960);
or U24520 (N_24520,N_18362,N_13833);
or U24521 (N_24521,N_13704,N_15290);
xnor U24522 (N_24522,N_12755,N_11140);
nand U24523 (N_24523,N_12014,N_13429);
nand U24524 (N_24524,N_10409,N_12979);
or U24525 (N_24525,N_10945,N_11848);
xor U24526 (N_24526,N_16480,N_17963);
nor U24527 (N_24527,N_14131,N_18481);
and U24528 (N_24528,N_17102,N_19907);
and U24529 (N_24529,N_12938,N_14937);
nand U24530 (N_24530,N_16618,N_12051);
nor U24531 (N_24531,N_16526,N_18422);
and U24532 (N_24532,N_10841,N_17604);
and U24533 (N_24533,N_17707,N_15938);
nand U24534 (N_24534,N_17840,N_12172);
or U24535 (N_24535,N_13895,N_16509);
or U24536 (N_24536,N_16573,N_10602);
or U24537 (N_24537,N_13627,N_14430);
or U24538 (N_24538,N_19173,N_19328);
nor U24539 (N_24539,N_17954,N_12631);
nor U24540 (N_24540,N_11231,N_10103);
nor U24541 (N_24541,N_12966,N_12925);
nor U24542 (N_24542,N_14770,N_15769);
or U24543 (N_24543,N_12526,N_10522);
and U24544 (N_24544,N_17231,N_12905);
nor U24545 (N_24545,N_15723,N_12018);
nor U24546 (N_24546,N_11762,N_10613);
or U24547 (N_24547,N_14614,N_16952);
or U24548 (N_24548,N_10552,N_11880);
nor U24549 (N_24549,N_18282,N_11533);
xnor U24550 (N_24550,N_14785,N_18851);
or U24551 (N_24551,N_12475,N_14913);
nor U24552 (N_24552,N_16901,N_19568);
or U24553 (N_24553,N_12197,N_13744);
xor U24554 (N_24554,N_17232,N_18360);
xor U24555 (N_24555,N_16226,N_14326);
nand U24556 (N_24556,N_17544,N_19033);
and U24557 (N_24557,N_19865,N_18134);
or U24558 (N_24558,N_11453,N_15252);
nand U24559 (N_24559,N_12307,N_15615);
nand U24560 (N_24560,N_18963,N_17935);
xor U24561 (N_24561,N_18859,N_14688);
or U24562 (N_24562,N_13167,N_10539);
and U24563 (N_24563,N_17571,N_12125);
nor U24564 (N_24564,N_13942,N_15533);
or U24565 (N_24565,N_10057,N_14282);
and U24566 (N_24566,N_12842,N_14105);
nor U24567 (N_24567,N_14941,N_16070);
nor U24568 (N_24568,N_13645,N_17211);
or U24569 (N_24569,N_11732,N_17803);
and U24570 (N_24570,N_12619,N_12365);
or U24571 (N_24571,N_17027,N_11012);
or U24572 (N_24572,N_10865,N_19669);
or U24573 (N_24573,N_17185,N_19652);
nand U24574 (N_24574,N_19512,N_19523);
and U24575 (N_24575,N_10524,N_10886);
xor U24576 (N_24576,N_10169,N_13452);
and U24577 (N_24577,N_16930,N_16794);
and U24578 (N_24578,N_16911,N_15670);
nand U24579 (N_24579,N_13774,N_19593);
or U24580 (N_24580,N_18686,N_18180);
nor U24581 (N_24581,N_16696,N_11613);
and U24582 (N_24582,N_17059,N_14457);
xnor U24583 (N_24583,N_17930,N_18382);
nor U24584 (N_24584,N_11116,N_11170);
nand U24585 (N_24585,N_15717,N_12133);
or U24586 (N_24586,N_10799,N_14781);
nand U24587 (N_24587,N_11335,N_13813);
nor U24588 (N_24588,N_13090,N_10629);
nor U24589 (N_24589,N_16222,N_19421);
or U24590 (N_24590,N_14357,N_12855);
xnor U24591 (N_24591,N_11723,N_10908);
or U24592 (N_24592,N_13711,N_16271);
nor U24593 (N_24593,N_13531,N_17076);
nand U24594 (N_24594,N_12432,N_17324);
nor U24595 (N_24595,N_15616,N_12009);
nor U24596 (N_24596,N_15260,N_10501);
nor U24597 (N_24597,N_11320,N_14925);
or U24598 (N_24598,N_19703,N_13905);
and U24599 (N_24599,N_13632,N_11681);
nor U24600 (N_24600,N_15095,N_14882);
nand U24601 (N_24601,N_11797,N_15079);
or U24602 (N_24602,N_16844,N_19510);
nor U24603 (N_24603,N_17281,N_18028);
nand U24604 (N_24604,N_11661,N_15808);
or U24605 (N_24605,N_15207,N_16698);
and U24606 (N_24606,N_11535,N_15382);
or U24607 (N_24607,N_14337,N_17872);
or U24608 (N_24608,N_13586,N_17003);
or U24609 (N_24609,N_12206,N_13997);
nand U24610 (N_24610,N_11083,N_12041);
nor U24611 (N_24611,N_19044,N_14037);
xnor U24612 (N_24612,N_19481,N_17352);
or U24613 (N_24613,N_10257,N_18858);
xor U24614 (N_24614,N_13560,N_11478);
nand U24615 (N_24615,N_11060,N_12364);
nand U24616 (N_24616,N_11549,N_12463);
nand U24617 (N_24617,N_19486,N_14897);
and U24618 (N_24618,N_14314,N_16433);
and U24619 (N_24619,N_10660,N_18233);
nand U24620 (N_24620,N_11284,N_16434);
xnor U24621 (N_24621,N_12710,N_19178);
nand U24622 (N_24622,N_18444,N_16936);
and U24623 (N_24623,N_19122,N_13182);
nor U24624 (N_24624,N_18644,N_14480);
nand U24625 (N_24625,N_15413,N_13568);
nand U24626 (N_24626,N_17494,N_16486);
or U24627 (N_24627,N_13391,N_16782);
xor U24628 (N_24628,N_11703,N_17984);
nor U24629 (N_24629,N_10557,N_15659);
xnor U24630 (N_24630,N_18565,N_17657);
or U24631 (N_24631,N_11823,N_11286);
xnor U24632 (N_24632,N_19414,N_16612);
and U24633 (N_24633,N_17550,N_10713);
and U24634 (N_24634,N_12490,N_13772);
or U24635 (N_24635,N_16392,N_19764);
nand U24636 (N_24636,N_11166,N_13870);
nor U24637 (N_24637,N_11740,N_17548);
nor U24638 (N_24638,N_12680,N_15271);
nand U24639 (N_24639,N_19357,N_18902);
nand U24640 (N_24640,N_18530,N_15182);
and U24641 (N_24641,N_11361,N_13263);
nor U24642 (N_24642,N_10115,N_13256);
or U24643 (N_24643,N_16626,N_14261);
nand U24644 (N_24644,N_12538,N_16735);
or U24645 (N_24645,N_11825,N_11092);
and U24646 (N_24646,N_12519,N_14584);
nand U24647 (N_24647,N_17748,N_11068);
nor U24648 (N_24648,N_19577,N_18903);
and U24649 (N_24649,N_10096,N_16209);
and U24650 (N_24650,N_11983,N_18062);
nand U24651 (N_24651,N_18117,N_14340);
nand U24652 (N_24652,N_14155,N_12381);
nor U24653 (N_24653,N_17004,N_18320);
and U24654 (N_24654,N_19970,N_19223);
nor U24655 (N_24655,N_18306,N_11518);
nand U24656 (N_24656,N_10659,N_14226);
and U24657 (N_24657,N_16691,N_16337);
nand U24658 (N_24658,N_17051,N_10439);
or U24659 (N_24659,N_17368,N_12159);
nor U24660 (N_24660,N_15710,N_14725);
and U24661 (N_24661,N_17850,N_17790);
xor U24662 (N_24662,N_18812,N_12335);
or U24663 (N_24663,N_14111,N_15746);
xor U24664 (N_24664,N_11947,N_15589);
nand U24665 (N_24665,N_17374,N_12447);
nor U24666 (N_24666,N_13939,N_10919);
xor U24667 (N_24667,N_18977,N_17498);
or U24668 (N_24668,N_10099,N_12518);
or U24669 (N_24669,N_14632,N_19536);
or U24670 (N_24670,N_12248,N_17186);
and U24671 (N_24671,N_11886,N_18994);
xnor U24672 (N_24672,N_16786,N_12128);
or U24673 (N_24673,N_10289,N_16342);
xor U24674 (N_24674,N_10596,N_17874);
xor U24675 (N_24675,N_14246,N_17502);
nor U24676 (N_24676,N_14672,N_15674);
or U24677 (N_24677,N_18199,N_19628);
and U24678 (N_24678,N_11544,N_13005);
and U24679 (N_24679,N_17432,N_11839);
and U24680 (N_24680,N_18445,N_10173);
nand U24681 (N_24681,N_15221,N_14704);
and U24682 (N_24682,N_15146,N_11576);
and U24683 (N_24683,N_17909,N_14344);
and U24684 (N_24684,N_11696,N_14200);
nand U24685 (N_24685,N_13489,N_14252);
nand U24686 (N_24686,N_14487,N_16089);
nor U24687 (N_24687,N_15094,N_13094);
xor U24688 (N_24688,N_15386,N_19068);
and U24689 (N_24689,N_14151,N_17523);
or U24690 (N_24690,N_11590,N_13846);
and U24691 (N_24691,N_17805,N_16462);
nand U24692 (N_24692,N_15720,N_10236);
or U24693 (N_24693,N_18119,N_10348);
xor U24694 (N_24694,N_17801,N_18176);
and U24695 (N_24695,N_14497,N_12626);
nor U24696 (N_24696,N_16493,N_17467);
nor U24697 (N_24697,N_11000,N_12326);
xnor U24698 (N_24698,N_18055,N_17919);
or U24699 (N_24699,N_11009,N_13887);
and U24700 (N_24700,N_15335,N_18323);
xor U24701 (N_24701,N_14998,N_14673);
or U24702 (N_24702,N_12783,N_19908);
xnor U24703 (N_24703,N_17652,N_18116);
and U24704 (N_24704,N_11927,N_12149);
and U24705 (N_24705,N_12316,N_17023);
nand U24706 (N_24706,N_17888,N_13671);
nor U24707 (N_24707,N_10300,N_19634);
or U24708 (N_24708,N_16921,N_12362);
nand U24709 (N_24709,N_10571,N_16895);
xor U24710 (N_24710,N_18803,N_10649);
nor U24711 (N_24711,N_11494,N_10896);
nor U24712 (N_24712,N_17493,N_11104);
or U24713 (N_24713,N_10866,N_10089);
and U24714 (N_24714,N_15089,N_10033);
or U24715 (N_24715,N_16133,N_17798);
and U24716 (N_24716,N_16697,N_14417);
nand U24717 (N_24717,N_17166,N_17339);
or U24718 (N_24718,N_18418,N_11700);
xor U24719 (N_24719,N_16743,N_15510);
or U24720 (N_24720,N_18899,N_16885);
and U24721 (N_24721,N_14910,N_12173);
nor U24722 (N_24722,N_14533,N_12988);
nand U24723 (N_24723,N_19455,N_17853);
xor U24724 (N_24724,N_19632,N_15642);
or U24725 (N_24725,N_11147,N_16608);
xnor U24726 (N_24726,N_19691,N_14877);
nor U24727 (N_24727,N_18773,N_18186);
or U24728 (N_24728,N_19077,N_18964);
nand U24729 (N_24729,N_14245,N_15534);
and U24730 (N_24730,N_13283,N_17348);
or U24731 (N_24731,N_16391,N_15563);
and U24732 (N_24732,N_12092,N_19877);
or U24733 (N_24733,N_19114,N_10785);
and U24734 (N_24734,N_13803,N_11110);
nand U24735 (N_24735,N_17039,N_14062);
nand U24736 (N_24736,N_17214,N_18454);
nand U24737 (N_24737,N_18111,N_13855);
and U24738 (N_24738,N_16644,N_12007);
nor U24739 (N_24739,N_12270,N_13202);
or U24740 (N_24740,N_16868,N_12689);
and U24741 (N_24741,N_10595,N_12661);
nor U24742 (N_24742,N_10277,N_15797);
nor U24743 (N_24743,N_16477,N_12020);
xor U24744 (N_24744,N_11285,N_11526);
and U24745 (N_24745,N_18265,N_11904);
xor U24746 (N_24746,N_12476,N_12122);
nand U24747 (N_24747,N_17444,N_19732);
xnor U24748 (N_24748,N_18287,N_19366);
nor U24749 (N_24749,N_12556,N_13275);
or U24750 (N_24750,N_14286,N_16243);
or U24751 (N_24751,N_13779,N_17988);
nor U24752 (N_24752,N_11855,N_13383);
and U24753 (N_24753,N_14362,N_13684);
or U24754 (N_24754,N_14999,N_17641);
nor U24755 (N_24755,N_12515,N_15331);
nand U24756 (N_24756,N_17918,N_14552);
xor U24757 (N_24757,N_10471,N_11427);
nor U24758 (N_24758,N_15579,N_15346);
and U24759 (N_24759,N_16630,N_13277);
nor U24760 (N_24760,N_15103,N_12205);
and U24761 (N_24761,N_18128,N_11959);
nor U24762 (N_24762,N_19891,N_15121);
or U24763 (N_24763,N_15773,N_19826);
nor U24764 (N_24764,N_15024,N_17643);
or U24765 (N_24765,N_10231,N_14936);
xnor U24766 (N_24766,N_15464,N_10129);
nor U24767 (N_24767,N_15832,N_15078);
and U24768 (N_24768,N_10294,N_11380);
nor U24769 (N_24769,N_17397,N_10075);
nand U24770 (N_24770,N_15470,N_16473);
and U24771 (N_24771,N_16325,N_13934);
and U24772 (N_24772,N_17419,N_15766);
or U24773 (N_24773,N_14435,N_11262);
nor U24774 (N_24774,N_14981,N_11946);
xnor U24775 (N_24775,N_11705,N_12935);
xor U24776 (N_24776,N_15258,N_19784);
xnor U24777 (N_24777,N_13158,N_14002);
nor U24778 (N_24778,N_15786,N_12102);
or U24779 (N_24779,N_15814,N_12635);
or U24780 (N_24780,N_17579,N_16088);
nand U24781 (N_24781,N_18491,N_16605);
and U24782 (N_24782,N_13823,N_12241);
xnor U24783 (N_24783,N_18616,N_13282);
nand U24784 (N_24784,N_18441,N_19446);
xnor U24785 (N_24785,N_11826,N_15961);
nor U24786 (N_24786,N_19101,N_10284);
nor U24787 (N_24787,N_19190,N_17555);
and U24788 (N_24788,N_15406,N_12682);
nor U24789 (N_24789,N_14950,N_13732);
nor U24790 (N_24790,N_17956,N_18707);
or U24791 (N_24791,N_17490,N_17503);
nand U24792 (N_24792,N_13116,N_18750);
or U24793 (N_24793,N_17113,N_10975);
nor U24794 (N_24794,N_17393,N_14447);
or U24795 (N_24795,N_18640,N_18835);
nor U24796 (N_24796,N_13582,N_17451);
xnor U24797 (N_24797,N_18353,N_17052);
nor U24798 (N_24798,N_18219,N_10107);
nand U24799 (N_24799,N_19358,N_10008);
nand U24800 (N_24800,N_18223,N_17182);
xor U24801 (N_24801,N_11129,N_11020);
and U24802 (N_24802,N_10335,N_19325);
or U24803 (N_24803,N_10821,N_12804);
and U24804 (N_24804,N_18546,N_10014);
and U24805 (N_24805,N_13066,N_15057);
and U24806 (N_24806,N_12536,N_19418);
nand U24807 (N_24807,N_15987,N_12416);
or U24808 (N_24808,N_10028,N_19073);
nor U24809 (N_24809,N_12576,N_16519);
xnor U24810 (N_24810,N_18951,N_19805);
and U24811 (N_24811,N_19867,N_17092);
xnor U24812 (N_24812,N_17002,N_13486);
and U24813 (N_24813,N_15419,N_12276);
xor U24814 (N_24814,N_10891,N_19752);
and U24815 (N_24815,N_14419,N_14992);
or U24816 (N_24816,N_11303,N_18888);
xnor U24817 (N_24817,N_17101,N_12945);
nand U24818 (N_24818,N_11562,N_14931);
and U24819 (N_24819,N_15241,N_11222);
and U24820 (N_24820,N_14004,N_16716);
nand U24821 (N_24821,N_12114,N_11205);
and U24822 (N_24822,N_13619,N_19152);
nor U24823 (N_24823,N_19398,N_13733);
xor U24824 (N_24824,N_10366,N_17793);
nand U24825 (N_24825,N_10577,N_18598);
or U24826 (N_24826,N_13712,N_13284);
or U24827 (N_24827,N_18297,N_11500);
nand U24828 (N_24828,N_17671,N_16955);
or U24829 (N_24829,N_15526,N_17704);
nor U24830 (N_24830,N_18030,N_10518);
and U24831 (N_24831,N_16109,N_18822);
xor U24832 (N_24832,N_15339,N_17644);
nor U24833 (N_24833,N_16968,N_14957);
xnor U24834 (N_24834,N_19502,N_16374);
and U24835 (N_24835,N_16130,N_16471);
nor U24836 (N_24836,N_13185,N_17615);
or U24837 (N_24837,N_19586,N_18712);
xnor U24838 (N_24838,N_13046,N_17629);
and U24839 (N_24839,N_17020,N_16176);
nand U24840 (N_24840,N_11583,N_19311);
nor U24841 (N_24841,N_13562,N_12708);
and U24842 (N_24842,N_18264,N_16200);
nand U24843 (N_24843,N_13039,N_12211);
nand U24844 (N_24844,N_18688,N_16492);
and U24845 (N_24845,N_15041,N_19001);
and U24846 (N_24846,N_13352,N_12500);
nand U24847 (N_24847,N_19984,N_19197);
nand U24848 (N_24848,N_18563,N_18935);
nor U24849 (N_24849,N_19262,N_11197);
and U24850 (N_24850,N_16860,N_13538);
or U24851 (N_24851,N_13646,N_18151);
nand U24852 (N_24852,N_14424,N_13994);
xor U24853 (N_24853,N_13406,N_16263);
xor U24854 (N_24854,N_19355,N_10210);
nand U24855 (N_24855,N_10194,N_10561);
and U24856 (N_24856,N_14747,N_11869);
or U24857 (N_24857,N_16152,N_11552);
and U24858 (N_24858,N_12053,N_13220);
xnor U24859 (N_24859,N_14274,N_12026);
nand U24860 (N_24860,N_15341,N_14364);
nor U24861 (N_24861,N_13868,N_19933);
and U24862 (N_24862,N_14542,N_16810);
nand U24863 (N_24863,N_10630,N_10322);
or U24864 (N_24864,N_18744,N_19542);
nand U24865 (N_24865,N_14685,N_10910);
and U24866 (N_24866,N_12402,N_16693);
xnor U24867 (N_24867,N_10747,N_16345);
and U24868 (N_24868,N_16642,N_17985);
xor U24869 (N_24869,N_10796,N_17421);
or U24870 (N_24870,N_12931,N_15673);
nand U24871 (N_24871,N_18314,N_13249);
nand U24872 (N_24872,N_16559,N_17125);
nor U24873 (N_24873,N_13269,N_17328);
nand U24874 (N_24874,N_17784,N_18455);
and U24875 (N_24875,N_19422,N_15764);
nor U24876 (N_24876,N_11133,N_18769);
xnor U24877 (N_24877,N_16645,N_17465);
and U24878 (N_24878,N_11821,N_11625);
nor U24879 (N_24879,N_14436,N_14934);
or U24880 (N_24880,N_14707,N_16506);
nand U24881 (N_24881,N_11256,N_12188);
xor U24882 (N_24882,N_13497,N_13896);
or U24883 (N_24883,N_10907,N_19862);
or U24884 (N_24884,N_12207,N_15810);
or U24885 (N_24885,N_12984,N_19591);
nor U24886 (N_24886,N_13826,N_16680);
or U24887 (N_24887,N_15387,N_19337);
nor U24888 (N_24888,N_12898,N_12636);
xor U24889 (N_24889,N_17333,N_10558);
and U24890 (N_24890,N_17982,N_17905);
nand U24891 (N_24891,N_15316,N_13898);
or U24892 (N_24892,N_10091,N_16378);
nor U24893 (N_24893,N_13781,N_16278);
nor U24894 (N_24894,N_14828,N_18760);
and U24895 (N_24895,N_15455,N_19022);
nand U24896 (N_24896,N_14174,N_19164);
and U24897 (N_24897,N_11344,N_16924);
nand U24898 (N_24898,N_12145,N_16515);
nand U24899 (N_24899,N_15704,N_15602);
xor U24900 (N_24900,N_15643,N_15032);
nor U24901 (N_24901,N_14082,N_10408);
xor U24902 (N_24902,N_10753,N_12314);
or U24903 (N_24903,N_19768,N_16763);
or U24904 (N_24904,N_10022,N_17557);
and U24905 (N_24905,N_17881,N_17880);
xor U24906 (N_24906,N_12065,N_18661);
nand U24907 (N_24907,N_16663,N_16045);
or U24908 (N_24908,N_19423,N_10006);
or U24909 (N_24909,N_15891,N_16202);
nand U24910 (N_24910,N_10404,N_10258);
xor U24911 (N_24911,N_12038,N_10843);
and U24912 (N_24912,N_11118,N_13640);
xnor U24913 (N_24913,N_14074,N_16622);
xor U24914 (N_24914,N_14540,N_15597);
xor U24915 (N_24915,N_16108,N_14811);
nand U24916 (N_24916,N_12204,N_16531);
nor U24917 (N_24917,N_19544,N_17244);
or U24918 (N_24918,N_18203,N_11280);
or U24919 (N_24919,N_15345,N_17074);
and U24920 (N_24920,N_11159,N_13187);
and U24921 (N_24921,N_15371,N_19253);
and U24922 (N_24922,N_19338,N_11585);
nand U24923 (N_24923,N_17844,N_13104);
and U24924 (N_24924,N_17701,N_17889);
and U24925 (N_24925,N_12085,N_17217);
or U24926 (N_24926,N_18093,N_18005);
xnor U24927 (N_24927,N_19782,N_14948);
and U24928 (N_24928,N_14726,N_18629);
nand U24929 (N_24929,N_16497,N_10012);
nand U24930 (N_24930,N_13837,N_16816);
nor U24931 (N_24931,N_13650,N_12853);
or U24932 (N_24932,N_18540,N_18642);
and U24933 (N_24933,N_16048,N_19242);
xor U24934 (N_24934,N_16578,N_10244);
nand U24935 (N_24935,N_13466,N_11728);
nand U24936 (N_24936,N_16554,N_13996);
xor U24937 (N_24937,N_13951,N_13543);
nor U24938 (N_24938,N_14660,N_17279);
nor U24939 (N_24939,N_11069,N_18408);
xnor U24940 (N_24940,N_15458,N_11479);
or U24941 (N_24941,N_18401,N_15541);
xnor U24942 (N_24942,N_17238,N_10547);
nor U24943 (N_24943,N_19304,N_11111);
and U24944 (N_24944,N_18173,N_19913);
or U24945 (N_24945,N_10216,N_11329);
nor U24946 (N_24946,N_10822,N_10970);
nor U24947 (N_24947,N_15228,N_16646);
nand U24948 (N_24948,N_10691,N_14894);
xnor U24949 (N_24949,N_10646,N_11816);
nand U24950 (N_24950,N_13509,N_19144);
and U24951 (N_24951,N_12506,N_18795);
nand U24952 (N_24952,N_13664,N_17924);
and U24953 (N_24953,N_13751,N_13077);
nand U24954 (N_24954,N_13788,N_14311);
nor U24955 (N_24955,N_17563,N_13707);
xor U24956 (N_24956,N_16367,N_15482);
nand U24957 (N_24957,N_19488,N_14942);
xnor U24958 (N_24958,N_14927,N_17607);
xor U24959 (N_24959,N_16668,N_12995);
nand U24960 (N_24960,N_10795,N_15336);
and U24961 (N_24961,N_11530,N_12846);
xnor U24962 (N_24962,N_17097,N_19841);
nand U24963 (N_24963,N_13693,N_18940);
or U24964 (N_24964,N_17860,N_12950);
xor U24965 (N_24965,N_15188,N_15004);
nand U24966 (N_24966,N_14679,N_13164);
nor U24967 (N_24967,N_12244,N_15096);
xnor U24968 (N_24968,N_11651,N_10268);
and U24969 (N_24969,N_19947,N_12071);
xor U24970 (N_24970,N_15552,N_17848);
or U24971 (N_24971,N_11962,N_15369);
nand U24972 (N_24972,N_15521,N_17199);
xnor U24973 (N_24973,N_14926,N_12223);
nand U24974 (N_24974,N_18341,N_12723);
nor U24975 (N_24975,N_15159,N_15100);
nand U24976 (N_24976,N_19870,N_15312);
nor U24977 (N_24977,N_13119,N_16171);
or U24978 (N_24978,N_19715,N_11538);
nand U24979 (N_24979,N_19165,N_14738);
xnor U24980 (N_24980,N_10247,N_19048);
nor U24981 (N_24981,N_10238,N_15323);
and U24982 (N_24982,N_14353,N_19817);
nand U24983 (N_24983,N_10205,N_13411);
xor U24984 (N_24984,N_17583,N_12892);
and U24985 (N_24985,N_11363,N_13458);
xnor U24986 (N_24986,N_10653,N_15698);
xor U24987 (N_24987,N_13731,N_10635);
or U24988 (N_24988,N_10136,N_17013);
xor U24989 (N_24989,N_19923,N_16498);
nor U24990 (N_24990,N_13941,N_13484);
and U24991 (N_24991,N_15542,N_18650);
nand U24992 (N_24992,N_14324,N_17911);
xor U24993 (N_24993,N_15445,N_12955);
or U24994 (N_24994,N_12347,N_11595);
or U24995 (N_24995,N_15204,N_15811);
xor U24996 (N_24996,N_12181,N_14844);
and U24997 (N_24997,N_16460,N_18538);
or U24998 (N_24998,N_17987,N_12559);
and U24999 (N_24999,N_14104,N_18500);
or U25000 (N_25000,N_16705,N_12792);
nor U25001 (N_25001,N_12646,N_11436);
xor U25002 (N_25002,N_18312,N_15129);
nand U25003 (N_25003,N_15184,N_12337);
nand U25004 (N_25004,N_11538,N_14449);
and U25005 (N_25005,N_14244,N_12784);
nand U25006 (N_25006,N_10018,N_12280);
nor U25007 (N_25007,N_17478,N_18592);
or U25008 (N_25008,N_12846,N_12789);
xnor U25009 (N_25009,N_15660,N_14580);
xor U25010 (N_25010,N_19835,N_12737);
or U25011 (N_25011,N_10817,N_13390);
xor U25012 (N_25012,N_16902,N_11498);
nor U25013 (N_25013,N_19856,N_12291);
xor U25014 (N_25014,N_16987,N_14175);
nand U25015 (N_25015,N_19012,N_11720);
or U25016 (N_25016,N_16404,N_17979);
and U25017 (N_25017,N_18521,N_10452);
and U25018 (N_25018,N_16210,N_18568);
or U25019 (N_25019,N_16302,N_11825);
nand U25020 (N_25020,N_11883,N_16950);
and U25021 (N_25021,N_10881,N_18117);
or U25022 (N_25022,N_15310,N_14318);
nand U25023 (N_25023,N_15448,N_12922);
nor U25024 (N_25024,N_14082,N_10474);
and U25025 (N_25025,N_15379,N_16811);
nand U25026 (N_25026,N_12676,N_18966);
and U25027 (N_25027,N_17363,N_15514);
or U25028 (N_25028,N_12258,N_14102);
or U25029 (N_25029,N_15685,N_18160);
and U25030 (N_25030,N_18711,N_17147);
and U25031 (N_25031,N_15088,N_18461);
xnor U25032 (N_25032,N_10254,N_14919);
or U25033 (N_25033,N_11131,N_19407);
nand U25034 (N_25034,N_11460,N_19712);
nor U25035 (N_25035,N_10843,N_19389);
xor U25036 (N_25036,N_18418,N_10634);
xor U25037 (N_25037,N_18496,N_18119);
or U25038 (N_25038,N_18102,N_19803);
nand U25039 (N_25039,N_17835,N_11232);
and U25040 (N_25040,N_15792,N_17032);
or U25041 (N_25041,N_19448,N_17603);
and U25042 (N_25042,N_11560,N_17328);
nand U25043 (N_25043,N_16842,N_14413);
or U25044 (N_25044,N_18767,N_16593);
nor U25045 (N_25045,N_16434,N_14702);
or U25046 (N_25046,N_10467,N_14444);
xor U25047 (N_25047,N_10445,N_16304);
or U25048 (N_25048,N_19556,N_12808);
nor U25049 (N_25049,N_16803,N_15643);
nor U25050 (N_25050,N_12557,N_12963);
xnor U25051 (N_25051,N_13080,N_14758);
and U25052 (N_25052,N_15373,N_10050);
and U25053 (N_25053,N_10644,N_18126);
nor U25054 (N_25054,N_10206,N_11360);
nand U25055 (N_25055,N_15086,N_19464);
xor U25056 (N_25056,N_18803,N_10437);
nand U25057 (N_25057,N_19237,N_14967);
or U25058 (N_25058,N_12038,N_15155);
nand U25059 (N_25059,N_19094,N_19363);
xor U25060 (N_25060,N_19416,N_10944);
nor U25061 (N_25061,N_13593,N_16862);
xnor U25062 (N_25062,N_12414,N_11702);
xor U25063 (N_25063,N_16179,N_15370);
nand U25064 (N_25064,N_11246,N_12937);
nor U25065 (N_25065,N_13087,N_12361);
xor U25066 (N_25066,N_10672,N_18364);
and U25067 (N_25067,N_12503,N_17198);
xnor U25068 (N_25068,N_17544,N_19472);
or U25069 (N_25069,N_18026,N_15001);
and U25070 (N_25070,N_16205,N_12870);
and U25071 (N_25071,N_13520,N_16010);
xor U25072 (N_25072,N_15189,N_10291);
or U25073 (N_25073,N_12550,N_10041);
or U25074 (N_25074,N_19111,N_14805);
nor U25075 (N_25075,N_18249,N_11404);
nor U25076 (N_25076,N_18412,N_13676);
nor U25077 (N_25077,N_11880,N_15789);
nand U25078 (N_25078,N_11959,N_11277);
nor U25079 (N_25079,N_11713,N_17539);
xnor U25080 (N_25080,N_10383,N_17349);
or U25081 (N_25081,N_19194,N_19864);
and U25082 (N_25082,N_18032,N_14827);
or U25083 (N_25083,N_10136,N_16059);
nor U25084 (N_25084,N_14092,N_12630);
or U25085 (N_25085,N_16747,N_14218);
nand U25086 (N_25086,N_16881,N_12056);
xnor U25087 (N_25087,N_17783,N_11355);
xnor U25088 (N_25088,N_12521,N_16740);
xnor U25089 (N_25089,N_15015,N_11580);
nor U25090 (N_25090,N_10202,N_12350);
nand U25091 (N_25091,N_13161,N_18006);
or U25092 (N_25092,N_18127,N_11036);
or U25093 (N_25093,N_10820,N_19560);
or U25094 (N_25094,N_10013,N_19985);
xor U25095 (N_25095,N_12465,N_12859);
or U25096 (N_25096,N_19441,N_12440);
xor U25097 (N_25097,N_12254,N_18941);
nor U25098 (N_25098,N_12944,N_14350);
and U25099 (N_25099,N_18664,N_17714);
nand U25100 (N_25100,N_16652,N_17640);
and U25101 (N_25101,N_13278,N_17284);
or U25102 (N_25102,N_15280,N_11645);
nand U25103 (N_25103,N_14674,N_13153);
xnor U25104 (N_25104,N_18979,N_16042);
xor U25105 (N_25105,N_13092,N_16605);
xor U25106 (N_25106,N_18862,N_17041);
nand U25107 (N_25107,N_17535,N_15949);
or U25108 (N_25108,N_17645,N_13106);
and U25109 (N_25109,N_14710,N_19080);
nand U25110 (N_25110,N_10755,N_11113);
or U25111 (N_25111,N_19023,N_19839);
and U25112 (N_25112,N_18603,N_16019);
xor U25113 (N_25113,N_16879,N_12406);
nand U25114 (N_25114,N_16572,N_18930);
and U25115 (N_25115,N_12614,N_16875);
xor U25116 (N_25116,N_18533,N_15200);
nor U25117 (N_25117,N_10133,N_18186);
or U25118 (N_25118,N_11582,N_11660);
and U25119 (N_25119,N_11541,N_11359);
xor U25120 (N_25120,N_10727,N_16186);
and U25121 (N_25121,N_11637,N_11877);
nor U25122 (N_25122,N_10443,N_19542);
xnor U25123 (N_25123,N_12973,N_17928);
nand U25124 (N_25124,N_17592,N_16577);
nand U25125 (N_25125,N_10569,N_11623);
nor U25126 (N_25126,N_13896,N_19995);
and U25127 (N_25127,N_13270,N_15748);
nor U25128 (N_25128,N_12009,N_10965);
nand U25129 (N_25129,N_19027,N_19281);
nand U25130 (N_25130,N_13082,N_12128);
xor U25131 (N_25131,N_10484,N_11223);
and U25132 (N_25132,N_11481,N_19617);
nor U25133 (N_25133,N_18206,N_13499);
nor U25134 (N_25134,N_12982,N_12364);
and U25135 (N_25135,N_19001,N_17254);
or U25136 (N_25136,N_17521,N_17498);
and U25137 (N_25137,N_13333,N_13558);
nor U25138 (N_25138,N_18437,N_15762);
and U25139 (N_25139,N_10766,N_12420);
nand U25140 (N_25140,N_13952,N_16529);
xnor U25141 (N_25141,N_19518,N_12673);
nand U25142 (N_25142,N_17113,N_19959);
xor U25143 (N_25143,N_15227,N_14374);
and U25144 (N_25144,N_16156,N_14847);
nor U25145 (N_25145,N_13677,N_12951);
and U25146 (N_25146,N_16079,N_10277);
nor U25147 (N_25147,N_12708,N_17905);
and U25148 (N_25148,N_16742,N_18285);
nand U25149 (N_25149,N_17717,N_18944);
or U25150 (N_25150,N_14181,N_18583);
nand U25151 (N_25151,N_13263,N_14313);
nor U25152 (N_25152,N_15144,N_19720);
nor U25153 (N_25153,N_11607,N_13703);
nor U25154 (N_25154,N_17245,N_10614);
and U25155 (N_25155,N_13413,N_18214);
nor U25156 (N_25156,N_15299,N_10808);
and U25157 (N_25157,N_16328,N_18068);
or U25158 (N_25158,N_14791,N_13732);
nand U25159 (N_25159,N_13081,N_15923);
and U25160 (N_25160,N_14253,N_14521);
nor U25161 (N_25161,N_12866,N_14697);
and U25162 (N_25162,N_16097,N_18087);
nand U25163 (N_25163,N_15807,N_17627);
or U25164 (N_25164,N_12472,N_19561);
nor U25165 (N_25165,N_11922,N_13480);
nor U25166 (N_25166,N_13393,N_15551);
nand U25167 (N_25167,N_15399,N_18196);
and U25168 (N_25168,N_10286,N_12189);
and U25169 (N_25169,N_10804,N_13202);
nand U25170 (N_25170,N_17408,N_14247);
and U25171 (N_25171,N_18787,N_15488);
nor U25172 (N_25172,N_10597,N_10390);
nand U25173 (N_25173,N_15961,N_12556);
xnor U25174 (N_25174,N_10977,N_15935);
xor U25175 (N_25175,N_19242,N_16340);
and U25176 (N_25176,N_10318,N_15509);
and U25177 (N_25177,N_11704,N_12973);
xor U25178 (N_25178,N_13779,N_12894);
and U25179 (N_25179,N_19259,N_15305);
and U25180 (N_25180,N_15482,N_13977);
nor U25181 (N_25181,N_14563,N_10757);
xor U25182 (N_25182,N_10344,N_18225);
and U25183 (N_25183,N_10275,N_14869);
or U25184 (N_25184,N_11253,N_18629);
nand U25185 (N_25185,N_10882,N_18922);
nand U25186 (N_25186,N_13533,N_18280);
and U25187 (N_25187,N_18351,N_14295);
or U25188 (N_25188,N_12336,N_16820);
xor U25189 (N_25189,N_19563,N_19248);
nand U25190 (N_25190,N_10771,N_12138);
nand U25191 (N_25191,N_19701,N_12076);
xor U25192 (N_25192,N_19596,N_15355);
nand U25193 (N_25193,N_18822,N_12907);
and U25194 (N_25194,N_11422,N_19909);
or U25195 (N_25195,N_15737,N_12549);
nor U25196 (N_25196,N_14990,N_13720);
and U25197 (N_25197,N_10724,N_15109);
nand U25198 (N_25198,N_10951,N_11868);
nand U25199 (N_25199,N_18321,N_10586);
nor U25200 (N_25200,N_10388,N_13469);
xnor U25201 (N_25201,N_18730,N_18711);
nor U25202 (N_25202,N_10915,N_17088);
nand U25203 (N_25203,N_10549,N_19210);
nand U25204 (N_25204,N_13173,N_19028);
xor U25205 (N_25205,N_15858,N_16380);
nand U25206 (N_25206,N_11134,N_11440);
xnor U25207 (N_25207,N_16307,N_13404);
nor U25208 (N_25208,N_16398,N_17705);
and U25209 (N_25209,N_13664,N_10769);
or U25210 (N_25210,N_18120,N_17010);
xnor U25211 (N_25211,N_11847,N_19104);
and U25212 (N_25212,N_14945,N_14486);
or U25213 (N_25213,N_19764,N_18391);
nand U25214 (N_25214,N_10016,N_10418);
or U25215 (N_25215,N_13617,N_19204);
and U25216 (N_25216,N_12465,N_15664);
xnor U25217 (N_25217,N_10031,N_13972);
nor U25218 (N_25218,N_15713,N_15808);
or U25219 (N_25219,N_18960,N_15634);
and U25220 (N_25220,N_17217,N_17837);
and U25221 (N_25221,N_16837,N_14905);
and U25222 (N_25222,N_18709,N_10881);
or U25223 (N_25223,N_18891,N_13076);
or U25224 (N_25224,N_12533,N_17721);
nor U25225 (N_25225,N_13215,N_18562);
or U25226 (N_25226,N_10606,N_18397);
xnor U25227 (N_25227,N_15531,N_13953);
xnor U25228 (N_25228,N_16897,N_19905);
xor U25229 (N_25229,N_18353,N_19544);
nand U25230 (N_25230,N_18826,N_12931);
xor U25231 (N_25231,N_15000,N_17429);
xnor U25232 (N_25232,N_11879,N_12885);
nand U25233 (N_25233,N_14715,N_15320);
or U25234 (N_25234,N_13579,N_19317);
and U25235 (N_25235,N_19529,N_15706);
nand U25236 (N_25236,N_11718,N_13183);
xnor U25237 (N_25237,N_12569,N_16463);
xnor U25238 (N_25238,N_19235,N_14192);
xor U25239 (N_25239,N_14146,N_13356);
or U25240 (N_25240,N_18370,N_19915);
nand U25241 (N_25241,N_15251,N_13287);
and U25242 (N_25242,N_12199,N_19883);
nor U25243 (N_25243,N_19327,N_17008);
nand U25244 (N_25244,N_12518,N_16290);
xor U25245 (N_25245,N_11457,N_19985);
and U25246 (N_25246,N_14279,N_16749);
nand U25247 (N_25247,N_14014,N_16696);
and U25248 (N_25248,N_18752,N_15736);
nand U25249 (N_25249,N_13019,N_15486);
nor U25250 (N_25250,N_11552,N_18894);
and U25251 (N_25251,N_15362,N_13022);
xnor U25252 (N_25252,N_13711,N_17856);
nand U25253 (N_25253,N_10689,N_15511);
and U25254 (N_25254,N_19111,N_19890);
and U25255 (N_25255,N_12879,N_16660);
and U25256 (N_25256,N_19006,N_13870);
or U25257 (N_25257,N_19963,N_10369);
nor U25258 (N_25258,N_12175,N_19673);
xnor U25259 (N_25259,N_19170,N_16411);
and U25260 (N_25260,N_10154,N_11760);
nor U25261 (N_25261,N_14115,N_10243);
or U25262 (N_25262,N_18564,N_10114);
nand U25263 (N_25263,N_14796,N_17467);
and U25264 (N_25264,N_18493,N_13924);
nor U25265 (N_25265,N_12175,N_12185);
nor U25266 (N_25266,N_18732,N_12950);
or U25267 (N_25267,N_17971,N_19588);
nand U25268 (N_25268,N_13897,N_14314);
nand U25269 (N_25269,N_18672,N_11855);
xor U25270 (N_25270,N_13264,N_12096);
or U25271 (N_25271,N_16128,N_16691);
nand U25272 (N_25272,N_11211,N_12583);
xor U25273 (N_25273,N_13731,N_17351);
xor U25274 (N_25274,N_12999,N_13274);
xor U25275 (N_25275,N_19987,N_13312);
nor U25276 (N_25276,N_18672,N_19155);
and U25277 (N_25277,N_16779,N_16026);
nand U25278 (N_25278,N_19901,N_18249);
xnor U25279 (N_25279,N_10604,N_13677);
nor U25280 (N_25280,N_13818,N_12982);
and U25281 (N_25281,N_15927,N_14362);
nor U25282 (N_25282,N_12214,N_19433);
or U25283 (N_25283,N_19672,N_12789);
xor U25284 (N_25284,N_18169,N_11908);
nand U25285 (N_25285,N_14376,N_16452);
nor U25286 (N_25286,N_11548,N_19867);
nand U25287 (N_25287,N_17502,N_16987);
xnor U25288 (N_25288,N_13214,N_11514);
nor U25289 (N_25289,N_10897,N_15238);
xnor U25290 (N_25290,N_18566,N_16535);
and U25291 (N_25291,N_11178,N_19637);
or U25292 (N_25292,N_11281,N_19870);
and U25293 (N_25293,N_14635,N_16916);
or U25294 (N_25294,N_16502,N_10898);
nor U25295 (N_25295,N_11435,N_12992);
xnor U25296 (N_25296,N_17481,N_19524);
nor U25297 (N_25297,N_10499,N_18503);
or U25298 (N_25298,N_16299,N_13248);
nor U25299 (N_25299,N_16341,N_16402);
and U25300 (N_25300,N_15682,N_11571);
or U25301 (N_25301,N_17436,N_19079);
nor U25302 (N_25302,N_10129,N_15726);
nand U25303 (N_25303,N_17432,N_16080);
and U25304 (N_25304,N_11969,N_16533);
xnor U25305 (N_25305,N_16520,N_16921);
nand U25306 (N_25306,N_15012,N_13717);
nand U25307 (N_25307,N_14302,N_10569);
xnor U25308 (N_25308,N_19484,N_13570);
and U25309 (N_25309,N_13577,N_15424);
and U25310 (N_25310,N_19130,N_14272);
xnor U25311 (N_25311,N_18266,N_10017);
nor U25312 (N_25312,N_18400,N_13942);
and U25313 (N_25313,N_15246,N_16459);
xnor U25314 (N_25314,N_18273,N_10677);
xor U25315 (N_25315,N_11043,N_15924);
or U25316 (N_25316,N_17120,N_11478);
or U25317 (N_25317,N_18668,N_18516);
nor U25318 (N_25318,N_19594,N_15516);
nor U25319 (N_25319,N_11208,N_16680);
and U25320 (N_25320,N_16041,N_16632);
nor U25321 (N_25321,N_13313,N_18792);
nand U25322 (N_25322,N_11977,N_12822);
xnor U25323 (N_25323,N_12596,N_19531);
and U25324 (N_25324,N_15176,N_10191);
and U25325 (N_25325,N_11627,N_16850);
nor U25326 (N_25326,N_15782,N_12639);
nor U25327 (N_25327,N_11644,N_18411);
xnor U25328 (N_25328,N_14381,N_16214);
nor U25329 (N_25329,N_11589,N_16479);
and U25330 (N_25330,N_18578,N_18478);
and U25331 (N_25331,N_12849,N_19117);
nor U25332 (N_25332,N_11589,N_17662);
or U25333 (N_25333,N_18928,N_18614);
and U25334 (N_25334,N_14159,N_15828);
nand U25335 (N_25335,N_11054,N_19045);
xor U25336 (N_25336,N_12363,N_11704);
xor U25337 (N_25337,N_19105,N_15435);
nand U25338 (N_25338,N_18191,N_18085);
nand U25339 (N_25339,N_16619,N_18756);
nand U25340 (N_25340,N_12988,N_15749);
nand U25341 (N_25341,N_11370,N_12360);
nand U25342 (N_25342,N_15877,N_14116);
nor U25343 (N_25343,N_13401,N_12193);
and U25344 (N_25344,N_11809,N_18325);
or U25345 (N_25345,N_10159,N_12735);
nor U25346 (N_25346,N_15866,N_17779);
nand U25347 (N_25347,N_19898,N_17936);
nand U25348 (N_25348,N_11438,N_13388);
xor U25349 (N_25349,N_14761,N_14557);
nor U25350 (N_25350,N_19598,N_15307);
or U25351 (N_25351,N_16015,N_19052);
nand U25352 (N_25352,N_12222,N_13441);
and U25353 (N_25353,N_14759,N_11095);
nor U25354 (N_25354,N_19220,N_16666);
xor U25355 (N_25355,N_13462,N_13848);
or U25356 (N_25356,N_10904,N_12816);
and U25357 (N_25357,N_12596,N_18866);
or U25358 (N_25358,N_11459,N_19256);
or U25359 (N_25359,N_19503,N_12775);
nor U25360 (N_25360,N_13633,N_14028);
or U25361 (N_25361,N_14634,N_15153);
xor U25362 (N_25362,N_11016,N_18304);
xor U25363 (N_25363,N_15863,N_12175);
nor U25364 (N_25364,N_17471,N_16026);
and U25365 (N_25365,N_12949,N_13812);
and U25366 (N_25366,N_16627,N_14745);
xnor U25367 (N_25367,N_19839,N_16195);
and U25368 (N_25368,N_18736,N_13672);
xnor U25369 (N_25369,N_14872,N_18995);
xor U25370 (N_25370,N_13822,N_15811);
nand U25371 (N_25371,N_13561,N_13309);
or U25372 (N_25372,N_10088,N_18638);
xnor U25373 (N_25373,N_12847,N_16881);
nor U25374 (N_25374,N_15736,N_16010);
or U25375 (N_25375,N_18930,N_19480);
and U25376 (N_25376,N_10784,N_10697);
xnor U25377 (N_25377,N_13857,N_10122);
nand U25378 (N_25378,N_10066,N_15765);
and U25379 (N_25379,N_19240,N_12385);
or U25380 (N_25380,N_14458,N_13587);
nor U25381 (N_25381,N_16626,N_18931);
nor U25382 (N_25382,N_10216,N_18628);
or U25383 (N_25383,N_11845,N_19385);
nand U25384 (N_25384,N_15211,N_13648);
xor U25385 (N_25385,N_10570,N_18877);
or U25386 (N_25386,N_11601,N_19122);
nand U25387 (N_25387,N_16536,N_16191);
or U25388 (N_25388,N_15435,N_18988);
nand U25389 (N_25389,N_11566,N_11850);
xor U25390 (N_25390,N_10202,N_15944);
nand U25391 (N_25391,N_18986,N_11829);
or U25392 (N_25392,N_19004,N_17437);
and U25393 (N_25393,N_10049,N_15653);
nand U25394 (N_25394,N_11094,N_18227);
nand U25395 (N_25395,N_16961,N_18379);
xnor U25396 (N_25396,N_17900,N_19222);
nand U25397 (N_25397,N_19548,N_16252);
nand U25398 (N_25398,N_16988,N_19871);
nor U25399 (N_25399,N_14283,N_17681);
or U25400 (N_25400,N_11975,N_17119);
nor U25401 (N_25401,N_16704,N_16323);
nand U25402 (N_25402,N_19501,N_18857);
nor U25403 (N_25403,N_16861,N_15872);
nand U25404 (N_25404,N_12648,N_18536);
nor U25405 (N_25405,N_16935,N_15679);
nand U25406 (N_25406,N_13244,N_14682);
or U25407 (N_25407,N_19697,N_10704);
nor U25408 (N_25408,N_15713,N_14926);
or U25409 (N_25409,N_19800,N_11257);
xor U25410 (N_25410,N_18395,N_13112);
xor U25411 (N_25411,N_10944,N_16272);
and U25412 (N_25412,N_13725,N_16517);
and U25413 (N_25413,N_18890,N_10071);
or U25414 (N_25414,N_15692,N_18121);
nor U25415 (N_25415,N_17703,N_12007);
nand U25416 (N_25416,N_11283,N_12974);
nor U25417 (N_25417,N_17599,N_14383);
nor U25418 (N_25418,N_10046,N_13733);
or U25419 (N_25419,N_10119,N_15576);
and U25420 (N_25420,N_18721,N_10771);
and U25421 (N_25421,N_16182,N_12335);
and U25422 (N_25422,N_13426,N_11526);
nand U25423 (N_25423,N_18230,N_19044);
xor U25424 (N_25424,N_18696,N_14504);
nand U25425 (N_25425,N_19213,N_16719);
and U25426 (N_25426,N_12224,N_17573);
or U25427 (N_25427,N_11881,N_14006);
xnor U25428 (N_25428,N_18503,N_14203);
xnor U25429 (N_25429,N_19133,N_15742);
nand U25430 (N_25430,N_17358,N_16442);
nor U25431 (N_25431,N_11195,N_11569);
nand U25432 (N_25432,N_14483,N_11550);
nor U25433 (N_25433,N_17260,N_18383);
xnor U25434 (N_25434,N_11974,N_16316);
nor U25435 (N_25435,N_15527,N_19376);
nand U25436 (N_25436,N_12410,N_12000);
xnor U25437 (N_25437,N_11856,N_10174);
xnor U25438 (N_25438,N_12737,N_13596);
nor U25439 (N_25439,N_13608,N_13422);
or U25440 (N_25440,N_15068,N_14018);
nand U25441 (N_25441,N_10839,N_18179);
and U25442 (N_25442,N_17476,N_14685);
or U25443 (N_25443,N_16465,N_13880);
nor U25444 (N_25444,N_13109,N_15398);
nor U25445 (N_25445,N_19102,N_17822);
and U25446 (N_25446,N_17538,N_13834);
and U25447 (N_25447,N_18819,N_15772);
xor U25448 (N_25448,N_10127,N_11319);
or U25449 (N_25449,N_11967,N_13911);
or U25450 (N_25450,N_18683,N_10631);
or U25451 (N_25451,N_16835,N_13415);
xnor U25452 (N_25452,N_14388,N_19569);
nor U25453 (N_25453,N_12967,N_12998);
nor U25454 (N_25454,N_12433,N_10101);
nor U25455 (N_25455,N_12377,N_15278);
nand U25456 (N_25456,N_14440,N_10577);
and U25457 (N_25457,N_14786,N_16359);
xor U25458 (N_25458,N_14391,N_11932);
nor U25459 (N_25459,N_13976,N_12429);
xor U25460 (N_25460,N_18495,N_10439);
or U25461 (N_25461,N_14325,N_14018);
or U25462 (N_25462,N_14780,N_11438);
xor U25463 (N_25463,N_13352,N_18197);
or U25464 (N_25464,N_18635,N_10733);
nor U25465 (N_25465,N_19500,N_19296);
xnor U25466 (N_25466,N_19222,N_10960);
xor U25467 (N_25467,N_17142,N_13667);
and U25468 (N_25468,N_13527,N_16869);
nand U25469 (N_25469,N_17780,N_18250);
nand U25470 (N_25470,N_18253,N_15567);
nand U25471 (N_25471,N_12084,N_18912);
or U25472 (N_25472,N_14681,N_13094);
nor U25473 (N_25473,N_17039,N_14209);
and U25474 (N_25474,N_14452,N_12239);
and U25475 (N_25475,N_19669,N_12912);
nor U25476 (N_25476,N_13873,N_17140);
or U25477 (N_25477,N_12020,N_17941);
xnor U25478 (N_25478,N_17743,N_15353);
nor U25479 (N_25479,N_14672,N_15638);
or U25480 (N_25480,N_17842,N_15198);
and U25481 (N_25481,N_11509,N_19153);
and U25482 (N_25482,N_16674,N_10154);
xnor U25483 (N_25483,N_18750,N_18967);
nor U25484 (N_25484,N_12133,N_10692);
and U25485 (N_25485,N_18008,N_12864);
or U25486 (N_25486,N_10789,N_11948);
and U25487 (N_25487,N_15105,N_13556);
xnor U25488 (N_25488,N_17371,N_15128);
nand U25489 (N_25489,N_11656,N_18355);
nor U25490 (N_25490,N_17668,N_19027);
nor U25491 (N_25491,N_12219,N_18261);
nand U25492 (N_25492,N_18662,N_18722);
nand U25493 (N_25493,N_11469,N_16619);
nand U25494 (N_25494,N_19546,N_16652);
nor U25495 (N_25495,N_12980,N_14777);
xnor U25496 (N_25496,N_18128,N_19646);
nor U25497 (N_25497,N_18788,N_19291);
and U25498 (N_25498,N_17241,N_10565);
xnor U25499 (N_25499,N_15517,N_15109);
or U25500 (N_25500,N_19950,N_10173);
nor U25501 (N_25501,N_11672,N_19531);
or U25502 (N_25502,N_19025,N_15912);
nand U25503 (N_25503,N_14218,N_18624);
nand U25504 (N_25504,N_13922,N_17836);
nand U25505 (N_25505,N_19202,N_10300);
xnor U25506 (N_25506,N_13364,N_14075);
and U25507 (N_25507,N_13382,N_15176);
xor U25508 (N_25508,N_18925,N_15735);
nand U25509 (N_25509,N_14960,N_13576);
and U25510 (N_25510,N_17123,N_15161);
nand U25511 (N_25511,N_15349,N_12106);
and U25512 (N_25512,N_16766,N_12602);
and U25513 (N_25513,N_11210,N_19942);
nor U25514 (N_25514,N_16229,N_15577);
and U25515 (N_25515,N_13338,N_18148);
and U25516 (N_25516,N_14542,N_16843);
and U25517 (N_25517,N_19885,N_16048);
and U25518 (N_25518,N_15590,N_12383);
and U25519 (N_25519,N_16649,N_12343);
nand U25520 (N_25520,N_14412,N_13793);
xnor U25521 (N_25521,N_17026,N_12580);
and U25522 (N_25522,N_15305,N_17444);
or U25523 (N_25523,N_19587,N_13275);
or U25524 (N_25524,N_10200,N_13907);
nor U25525 (N_25525,N_15932,N_15006);
nand U25526 (N_25526,N_18344,N_17466);
xnor U25527 (N_25527,N_11024,N_15472);
or U25528 (N_25528,N_12819,N_17354);
xnor U25529 (N_25529,N_11744,N_16965);
nand U25530 (N_25530,N_11955,N_12136);
nand U25531 (N_25531,N_18116,N_12381);
xnor U25532 (N_25532,N_12149,N_17348);
and U25533 (N_25533,N_15172,N_18420);
and U25534 (N_25534,N_18055,N_17401);
nor U25535 (N_25535,N_15577,N_12325);
and U25536 (N_25536,N_14952,N_15248);
nor U25537 (N_25537,N_14309,N_15750);
nor U25538 (N_25538,N_15192,N_12052);
nand U25539 (N_25539,N_11213,N_19386);
xnor U25540 (N_25540,N_13067,N_14212);
and U25541 (N_25541,N_17839,N_19430);
nor U25542 (N_25542,N_14076,N_11552);
nand U25543 (N_25543,N_13967,N_16622);
xor U25544 (N_25544,N_18499,N_15212);
xnor U25545 (N_25545,N_19406,N_10959);
and U25546 (N_25546,N_19913,N_16401);
and U25547 (N_25547,N_16240,N_14972);
nor U25548 (N_25548,N_18580,N_10542);
and U25549 (N_25549,N_18732,N_17571);
nor U25550 (N_25550,N_10782,N_17328);
nand U25551 (N_25551,N_19672,N_15121);
xor U25552 (N_25552,N_19857,N_15912);
nand U25553 (N_25553,N_19240,N_19580);
and U25554 (N_25554,N_11476,N_11226);
nand U25555 (N_25555,N_15527,N_13521);
or U25556 (N_25556,N_19660,N_18328);
nor U25557 (N_25557,N_17174,N_11070);
xnor U25558 (N_25558,N_15754,N_11460);
nor U25559 (N_25559,N_12133,N_12165);
and U25560 (N_25560,N_19182,N_17051);
nand U25561 (N_25561,N_18475,N_13682);
xor U25562 (N_25562,N_11670,N_10997);
nor U25563 (N_25563,N_19114,N_15356);
or U25564 (N_25564,N_14085,N_13026);
and U25565 (N_25565,N_15807,N_11891);
or U25566 (N_25566,N_17439,N_16838);
and U25567 (N_25567,N_16299,N_18951);
nand U25568 (N_25568,N_10588,N_11598);
nand U25569 (N_25569,N_11568,N_11637);
and U25570 (N_25570,N_15563,N_15990);
nand U25571 (N_25571,N_13889,N_10729);
xor U25572 (N_25572,N_13483,N_10217);
xor U25573 (N_25573,N_17712,N_19329);
xnor U25574 (N_25574,N_19850,N_12432);
xor U25575 (N_25575,N_19845,N_10862);
and U25576 (N_25576,N_10010,N_12559);
nand U25577 (N_25577,N_13908,N_18129);
nand U25578 (N_25578,N_12275,N_15271);
or U25579 (N_25579,N_12224,N_12300);
and U25580 (N_25580,N_11603,N_16061);
nand U25581 (N_25581,N_18151,N_15793);
xnor U25582 (N_25582,N_17629,N_16747);
nor U25583 (N_25583,N_18098,N_12022);
nor U25584 (N_25584,N_10906,N_16291);
or U25585 (N_25585,N_17522,N_13884);
nand U25586 (N_25586,N_14018,N_14009);
nand U25587 (N_25587,N_11960,N_18134);
nand U25588 (N_25588,N_17709,N_13986);
xnor U25589 (N_25589,N_19916,N_19175);
nor U25590 (N_25590,N_17705,N_10072);
or U25591 (N_25591,N_10647,N_18079);
nand U25592 (N_25592,N_10844,N_10888);
xnor U25593 (N_25593,N_10147,N_14565);
nor U25594 (N_25594,N_14798,N_10983);
xnor U25595 (N_25595,N_16663,N_13114);
nor U25596 (N_25596,N_13316,N_10421);
and U25597 (N_25597,N_14595,N_19672);
nor U25598 (N_25598,N_13962,N_18982);
nand U25599 (N_25599,N_13836,N_15800);
or U25600 (N_25600,N_10668,N_13706);
nand U25601 (N_25601,N_16798,N_13074);
xor U25602 (N_25602,N_12732,N_11316);
xnor U25603 (N_25603,N_12665,N_12201);
nor U25604 (N_25604,N_15989,N_14873);
or U25605 (N_25605,N_10874,N_10760);
nand U25606 (N_25606,N_12508,N_12211);
nor U25607 (N_25607,N_17196,N_17921);
nor U25608 (N_25608,N_14014,N_19515);
nand U25609 (N_25609,N_18235,N_19857);
nor U25610 (N_25610,N_11202,N_11039);
and U25611 (N_25611,N_12365,N_18352);
nor U25612 (N_25612,N_14185,N_13428);
or U25613 (N_25613,N_17189,N_17500);
xnor U25614 (N_25614,N_11654,N_12640);
or U25615 (N_25615,N_19672,N_19873);
xnor U25616 (N_25616,N_17774,N_12090);
nor U25617 (N_25617,N_18603,N_12445);
nor U25618 (N_25618,N_12672,N_13767);
nor U25619 (N_25619,N_11753,N_19079);
or U25620 (N_25620,N_15030,N_12695);
xnor U25621 (N_25621,N_13508,N_17687);
or U25622 (N_25622,N_12361,N_18165);
or U25623 (N_25623,N_16753,N_18826);
xnor U25624 (N_25624,N_14793,N_12620);
nor U25625 (N_25625,N_13767,N_16044);
nor U25626 (N_25626,N_16537,N_14629);
nor U25627 (N_25627,N_11734,N_18629);
and U25628 (N_25628,N_18232,N_14656);
nor U25629 (N_25629,N_16636,N_12566);
or U25630 (N_25630,N_19824,N_12755);
or U25631 (N_25631,N_18991,N_14668);
xnor U25632 (N_25632,N_13145,N_11281);
and U25633 (N_25633,N_18418,N_13941);
or U25634 (N_25634,N_13112,N_19911);
nor U25635 (N_25635,N_14201,N_11617);
xor U25636 (N_25636,N_10713,N_12877);
nor U25637 (N_25637,N_12505,N_10502);
xnor U25638 (N_25638,N_19276,N_13090);
xor U25639 (N_25639,N_19659,N_12736);
nand U25640 (N_25640,N_13826,N_10611);
nor U25641 (N_25641,N_18708,N_14074);
nand U25642 (N_25642,N_17533,N_13647);
and U25643 (N_25643,N_17292,N_11406);
nand U25644 (N_25644,N_18491,N_14058);
nor U25645 (N_25645,N_16864,N_19564);
and U25646 (N_25646,N_10268,N_15012);
or U25647 (N_25647,N_10113,N_11646);
nand U25648 (N_25648,N_19289,N_18825);
or U25649 (N_25649,N_10834,N_15077);
xnor U25650 (N_25650,N_13216,N_17567);
or U25651 (N_25651,N_18636,N_15477);
and U25652 (N_25652,N_15246,N_10051);
xnor U25653 (N_25653,N_18638,N_11733);
nand U25654 (N_25654,N_14357,N_17113);
nor U25655 (N_25655,N_17709,N_12193);
xor U25656 (N_25656,N_11732,N_13676);
nand U25657 (N_25657,N_14322,N_17612);
and U25658 (N_25658,N_19402,N_15631);
or U25659 (N_25659,N_15807,N_17770);
xnor U25660 (N_25660,N_12973,N_12468);
or U25661 (N_25661,N_19669,N_12229);
xnor U25662 (N_25662,N_10873,N_19068);
nor U25663 (N_25663,N_11766,N_10163);
xnor U25664 (N_25664,N_16052,N_19640);
nor U25665 (N_25665,N_18132,N_14922);
nor U25666 (N_25666,N_13370,N_15382);
nor U25667 (N_25667,N_14879,N_11746);
or U25668 (N_25668,N_14151,N_16647);
or U25669 (N_25669,N_12845,N_19563);
nor U25670 (N_25670,N_19541,N_11636);
and U25671 (N_25671,N_11822,N_10834);
nor U25672 (N_25672,N_18928,N_18558);
xnor U25673 (N_25673,N_15001,N_12343);
nor U25674 (N_25674,N_15074,N_11746);
and U25675 (N_25675,N_17652,N_19009);
nand U25676 (N_25676,N_16568,N_14906);
and U25677 (N_25677,N_16182,N_19336);
and U25678 (N_25678,N_10132,N_15329);
nand U25679 (N_25679,N_10422,N_10376);
xnor U25680 (N_25680,N_17523,N_13449);
nor U25681 (N_25681,N_18620,N_19224);
nor U25682 (N_25682,N_19593,N_12836);
and U25683 (N_25683,N_16013,N_10324);
nor U25684 (N_25684,N_12353,N_17013);
or U25685 (N_25685,N_19820,N_12146);
and U25686 (N_25686,N_14554,N_12641);
xor U25687 (N_25687,N_17058,N_16717);
or U25688 (N_25688,N_16203,N_10092);
and U25689 (N_25689,N_15122,N_13305);
nand U25690 (N_25690,N_14914,N_14421);
or U25691 (N_25691,N_12015,N_10254);
and U25692 (N_25692,N_17173,N_17152);
nand U25693 (N_25693,N_18318,N_10473);
nor U25694 (N_25694,N_18926,N_18541);
or U25695 (N_25695,N_18535,N_18155);
nor U25696 (N_25696,N_11569,N_11570);
nand U25697 (N_25697,N_14343,N_11073);
nand U25698 (N_25698,N_10877,N_12254);
or U25699 (N_25699,N_16267,N_15758);
and U25700 (N_25700,N_10531,N_10893);
or U25701 (N_25701,N_12828,N_17212);
or U25702 (N_25702,N_16304,N_14293);
or U25703 (N_25703,N_15812,N_18763);
or U25704 (N_25704,N_11209,N_17227);
nand U25705 (N_25705,N_11759,N_12180);
and U25706 (N_25706,N_11688,N_16899);
nor U25707 (N_25707,N_19809,N_13319);
nor U25708 (N_25708,N_13325,N_12359);
nand U25709 (N_25709,N_15491,N_14151);
xnor U25710 (N_25710,N_15140,N_13173);
and U25711 (N_25711,N_10578,N_14561);
or U25712 (N_25712,N_18449,N_11147);
and U25713 (N_25713,N_12338,N_11992);
xnor U25714 (N_25714,N_11111,N_11507);
and U25715 (N_25715,N_14923,N_11054);
and U25716 (N_25716,N_13049,N_19009);
nor U25717 (N_25717,N_18611,N_12136);
and U25718 (N_25718,N_13889,N_17748);
nand U25719 (N_25719,N_14147,N_10450);
nor U25720 (N_25720,N_19410,N_10792);
xor U25721 (N_25721,N_10004,N_10257);
and U25722 (N_25722,N_10278,N_17921);
or U25723 (N_25723,N_10272,N_18789);
nand U25724 (N_25724,N_13535,N_19780);
or U25725 (N_25725,N_16978,N_18874);
xnor U25726 (N_25726,N_16424,N_15077);
xor U25727 (N_25727,N_12082,N_11744);
or U25728 (N_25728,N_13946,N_12947);
or U25729 (N_25729,N_13902,N_16116);
and U25730 (N_25730,N_14272,N_19620);
xor U25731 (N_25731,N_15503,N_10038);
nor U25732 (N_25732,N_17900,N_14400);
nand U25733 (N_25733,N_11358,N_18867);
nand U25734 (N_25734,N_15833,N_12939);
nor U25735 (N_25735,N_16065,N_14679);
nand U25736 (N_25736,N_11993,N_16749);
nor U25737 (N_25737,N_14663,N_15761);
or U25738 (N_25738,N_15632,N_18377);
and U25739 (N_25739,N_14331,N_10727);
nand U25740 (N_25740,N_19234,N_14855);
nor U25741 (N_25741,N_12332,N_10578);
and U25742 (N_25742,N_10482,N_13751);
xnor U25743 (N_25743,N_10494,N_10631);
or U25744 (N_25744,N_15437,N_16922);
nor U25745 (N_25745,N_17629,N_12667);
nor U25746 (N_25746,N_17665,N_18030);
nor U25747 (N_25747,N_19558,N_11131);
nor U25748 (N_25748,N_15213,N_10674);
nor U25749 (N_25749,N_18658,N_17814);
or U25750 (N_25750,N_16906,N_10240);
xor U25751 (N_25751,N_10329,N_16396);
xor U25752 (N_25752,N_10230,N_12425);
nor U25753 (N_25753,N_15322,N_17826);
nor U25754 (N_25754,N_13200,N_12451);
xnor U25755 (N_25755,N_14436,N_15092);
nor U25756 (N_25756,N_15903,N_16124);
nor U25757 (N_25757,N_18846,N_13545);
nor U25758 (N_25758,N_11583,N_11082);
nand U25759 (N_25759,N_14457,N_12790);
nor U25760 (N_25760,N_11324,N_18299);
nor U25761 (N_25761,N_12510,N_13854);
xor U25762 (N_25762,N_18230,N_14814);
and U25763 (N_25763,N_19978,N_10065);
xor U25764 (N_25764,N_15059,N_13110);
or U25765 (N_25765,N_16226,N_11496);
and U25766 (N_25766,N_12786,N_10791);
xor U25767 (N_25767,N_17228,N_17431);
nand U25768 (N_25768,N_19438,N_10048);
xnor U25769 (N_25769,N_14747,N_19523);
nor U25770 (N_25770,N_17961,N_16006);
or U25771 (N_25771,N_12899,N_10926);
and U25772 (N_25772,N_19200,N_12105);
nor U25773 (N_25773,N_15663,N_14905);
nand U25774 (N_25774,N_10231,N_17796);
nand U25775 (N_25775,N_17251,N_13294);
xnor U25776 (N_25776,N_10851,N_13444);
nand U25777 (N_25777,N_15851,N_10385);
xor U25778 (N_25778,N_19621,N_12809);
xnor U25779 (N_25779,N_15532,N_10981);
nand U25780 (N_25780,N_11378,N_18181);
and U25781 (N_25781,N_11350,N_14607);
or U25782 (N_25782,N_11862,N_13014);
xor U25783 (N_25783,N_10617,N_14760);
nor U25784 (N_25784,N_10806,N_15000);
nor U25785 (N_25785,N_13378,N_10962);
or U25786 (N_25786,N_12692,N_14712);
or U25787 (N_25787,N_16755,N_10611);
nand U25788 (N_25788,N_16418,N_13071);
nand U25789 (N_25789,N_11620,N_17596);
or U25790 (N_25790,N_19727,N_15740);
and U25791 (N_25791,N_17580,N_18837);
nor U25792 (N_25792,N_15347,N_13362);
xnor U25793 (N_25793,N_17162,N_19576);
xor U25794 (N_25794,N_12947,N_13762);
or U25795 (N_25795,N_13275,N_10981);
or U25796 (N_25796,N_10246,N_16885);
xnor U25797 (N_25797,N_19067,N_17856);
xnor U25798 (N_25798,N_13089,N_14645);
and U25799 (N_25799,N_19834,N_15660);
xnor U25800 (N_25800,N_14879,N_19956);
nand U25801 (N_25801,N_14111,N_17220);
and U25802 (N_25802,N_11997,N_15580);
xor U25803 (N_25803,N_11337,N_19383);
or U25804 (N_25804,N_12081,N_12671);
xnor U25805 (N_25805,N_16695,N_13592);
nand U25806 (N_25806,N_11920,N_11739);
nor U25807 (N_25807,N_11906,N_19298);
or U25808 (N_25808,N_18996,N_14558);
nand U25809 (N_25809,N_17159,N_18368);
nand U25810 (N_25810,N_12929,N_10280);
and U25811 (N_25811,N_10320,N_10625);
nor U25812 (N_25812,N_14708,N_10913);
xor U25813 (N_25813,N_10485,N_17811);
or U25814 (N_25814,N_11579,N_14900);
nor U25815 (N_25815,N_17966,N_17407);
nor U25816 (N_25816,N_10199,N_19783);
nand U25817 (N_25817,N_17580,N_10497);
nor U25818 (N_25818,N_14651,N_11849);
or U25819 (N_25819,N_13496,N_16191);
nand U25820 (N_25820,N_12730,N_19371);
nand U25821 (N_25821,N_14608,N_16882);
xnor U25822 (N_25822,N_16987,N_10445);
or U25823 (N_25823,N_18865,N_14306);
or U25824 (N_25824,N_16111,N_19443);
and U25825 (N_25825,N_17211,N_13385);
or U25826 (N_25826,N_18766,N_16788);
and U25827 (N_25827,N_15313,N_10243);
and U25828 (N_25828,N_18580,N_18392);
nor U25829 (N_25829,N_10092,N_10193);
and U25830 (N_25830,N_14422,N_17984);
and U25831 (N_25831,N_15010,N_17095);
nor U25832 (N_25832,N_13746,N_10917);
nor U25833 (N_25833,N_11054,N_16168);
or U25834 (N_25834,N_13810,N_17276);
and U25835 (N_25835,N_15599,N_15312);
xnor U25836 (N_25836,N_12040,N_10711);
nand U25837 (N_25837,N_17033,N_10867);
xor U25838 (N_25838,N_18857,N_17888);
nor U25839 (N_25839,N_19438,N_14018);
nor U25840 (N_25840,N_11698,N_12278);
xor U25841 (N_25841,N_12854,N_19755);
nand U25842 (N_25842,N_13861,N_19199);
and U25843 (N_25843,N_11206,N_18597);
xor U25844 (N_25844,N_17701,N_16598);
xor U25845 (N_25845,N_18562,N_13084);
xnor U25846 (N_25846,N_15677,N_10058);
nor U25847 (N_25847,N_19353,N_15521);
nand U25848 (N_25848,N_18154,N_15312);
xnor U25849 (N_25849,N_15455,N_13844);
or U25850 (N_25850,N_10359,N_11666);
and U25851 (N_25851,N_12024,N_11390);
xor U25852 (N_25852,N_14527,N_11210);
or U25853 (N_25853,N_14770,N_15351);
nand U25854 (N_25854,N_10539,N_12002);
and U25855 (N_25855,N_13639,N_17311);
and U25856 (N_25856,N_11945,N_11057);
nor U25857 (N_25857,N_13526,N_11398);
xor U25858 (N_25858,N_16014,N_15135);
or U25859 (N_25859,N_17115,N_17723);
or U25860 (N_25860,N_16092,N_15056);
nand U25861 (N_25861,N_13623,N_16683);
nand U25862 (N_25862,N_19760,N_10128);
xnor U25863 (N_25863,N_16251,N_13788);
and U25864 (N_25864,N_10071,N_14769);
or U25865 (N_25865,N_11896,N_17475);
xnor U25866 (N_25866,N_14325,N_14264);
nand U25867 (N_25867,N_10275,N_17194);
or U25868 (N_25868,N_15173,N_13589);
nor U25869 (N_25869,N_16280,N_12902);
nand U25870 (N_25870,N_15622,N_16136);
xnor U25871 (N_25871,N_10129,N_17629);
or U25872 (N_25872,N_14600,N_10579);
nor U25873 (N_25873,N_13383,N_16715);
nand U25874 (N_25874,N_15881,N_15627);
nand U25875 (N_25875,N_15068,N_15717);
and U25876 (N_25876,N_17436,N_12776);
xnor U25877 (N_25877,N_15532,N_11463);
nor U25878 (N_25878,N_14236,N_18501);
xnor U25879 (N_25879,N_16502,N_17815);
xnor U25880 (N_25880,N_12402,N_17543);
and U25881 (N_25881,N_16606,N_10276);
xor U25882 (N_25882,N_16832,N_10942);
xor U25883 (N_25883,N_10713,N_19782);
xnor U25884 (N_25884,N_13311,N_11253);
nor U25885 (N_25885,N_19261,N_12598);
xnor U25886 (N_25886,N_18365,N_13600);
or U25887 (N_25887,N_14390,N_18206);
xnor U25888 (N_25888,N_13090,N_13213);
and U25889 (N_25889,N_17103,N_18265);
nand U25890 (N_25890,N_11441,N_13798);
or U25891 (N_25891,N_14246,N_13439);
and U25892 (N_25892,N_13552,N_19650);
and U25893 (N_25893,N_13995,N_14538);
nor U25894 (N_25894,N_16844,N_15286);
and U25895 (N_25895,N_15856,N_13602);
or U25896 (N_25896,N_16210,N_11195);
nand U25897 (N_25897,N_19656,N_12600);
xor U25898 (N_25898,N_10817,N_11706);
nor U25899 (N_25899,N_14169,N_17818);
nor U25900 (N_25900,N_19594,N_14995);
xnor U25901 (N_25901,N_11454,N_10239);
and U25902 (N_25902,N_11269,N_19572);
nand U25903 (N_25903,N_16754,N_17653);
xor U25904 (N_25904,N_13559,N_19988);
nand U25905 (N_25905,N_11656,N_15265);
and U25906 (N_25906,N_10066,N_14675);
xor U25907 (N_25907,N_16731,N_11665);
or U25908 (N_25908,N_13191,N_11538);
nand U25909 (N_25909,N_15270,N_13791);
and U25910 (N_25910,N_11647,N_19696);
nor U25911 (N_25911,N_17208,N_18707);
nand U25912 (N_25912,N_11005,N_12089);
xnor U25913 (N_25913,N_19845,N_16507);
and U25914 (N_25914,N_14276,N_13107);
and U25915 (N_25915,N_11288,N_12943);
or U25916 (N_25916,N_15866,N_17650);
and U25917 (N_25917,N_14281,N_15842);
and U25918 (N_25918,N_18010,N_11900);
or U25919 (N_25919,N_13754,N_19679);
or U25920 (N_25920,N_13195,N_16037);
and U25921 (N_25921,N_19326,N_16301);
xor U25922 (N_25922,N_11797,N_15479);
nand U25923 (N_25923,N_10008,N_16691);
and U25924 (N_25924,N_18245,N_17901);
xnor U25925 (N_25925,N_14581,N_18775);
and U25926 (N_25926,N_15003,N_16716);
xnor U25927 (N_25927,N_18524,N_15445);
nand U25928 (N_25928,N_10033,N_12378);
nor U25929 (N_25929,N_17751,N_13829);
nor U25930 (N_25930,N_11887,N_14353);
or U25931 (N_25931,N_10994,N_15446);
nor U25932 (N_25932,N_15336,N_13844);
nand U25933 (N_25933,N_15938,N_13439);
nand U25934 (N_25934,N_11992,N_17700);
xnor U25935 (N_25935,N_15800,N_17788);
nand U25936 (N_25936,N_13827,N_13578);
nand U25937 (N_25937,N_19019,N_19462);
and U25938 (N_25938,N_19020,N_18709);
xor U25939 (N_25939,N_10258,N_19643);
or U25940 (N_25940,N_16512,N_10763);
nand U25941 (N_25941,N_12713,N_15290);
nand U25942 (N_25942,N_10254,N_16216);
and U25943 (N_25943,N_15835,N_11730);
and U25944 (N_25944,N_14096,N_10138);
and U25945 (N_25945,N_17242,N_17682);
nor U25946 (N_25946,N_19118,N_10934);
nand U25947 (N_25947,N_17417,N_17695);
xnor U25948 (N_25948,N_16273,N_17252);
or U25949 (N_25949,N_14589,N_16994);
nand U25950 (N_25950,N_13303,N_10759);
nand U25951 (N_25951,N_11178,N_19082);
xor U25952 (N_25952,N_16872,N_12363);
xnor U25953 (N_25953,N_12583,N_17437);
or U25954 (N_25954,N_11380,N_14684);
xor U25955 (N_25955,N_19617,N_18848);
nand U25956 (N_25956,N_19765,N_16813);
and U25957 (N_25957,N_18474,N_16204);
nor U25958 (N_25958,N_10812,N_11689);
nand U25959 (N_25959,N_17382,N_14878);
and U25960 (N_25960,N_18328,N_13705);
and U25961 (N_25961,N_19296,N_17550);
nor U25962 (N_25962,N_15490,N_15456);
nor U25963 (N_25963,N_11900,N_16909);
and U25964 (N_25964,N_18218,N_17804);
xnor U25965 (N_25965,N_13475,N_17583);
nor U25966 (N_25966,N_11583,N_10104);
xor U25967 (N_25967,N_12932,N_10799);
nor U25968 (N_25968,N_16895,N_12740);
nor U25969 (N_25969,N_19982,N_11687);
and U25970 (N_25970,N_10389,N_10199);
nand U25971 (N_25971,N_19712,N_11636);
nor U25972 (N_25972,N_10554,N_11450);
and U25973 (N_25973,N_15684,N_17723);
and U25974 (N_25974,N_16036,N_11887);
xor U25975 (N_25975,N_15480,N_16490);
nand U25976 (N_25976,N_17961,N_16102);
and U25977 (N_25977,N_17690,N_11978);
or U25978 (N_25978,N_15633,N_12978);
or U25979 (N_25979,N_16530,N_18723);
nand U25980 (N_25980,N_15671,N_18447);
or U25981 (N_25981,N_16920,N_11810);
or U25982 (N_25982,N_11227,N_16758);
nand U25983 (N_25983,N_11104,N_15502);
and U25984 (N_25984,N_18363,N_16742);
nor U25985 (N_25985,N_18661,N_18258);
and U25986 (N_25986,N_13430,N_12874);
nand U25987 (N_25987,N_16880,N_10339);
or U25988 (N_25988,N_18254,N_14857);
and U25989 (N_25989,N_10961,N_18206);
xnor U25990 (N_25990,N_12670,N_17673);
and U25991 (N_25991,N_18963,N_15981);
or U25992 (N_25992,N_19404,N_18435);
or U25993 (N_25993,N_15415,N_19700);
nor U25994 (N_25994,N_16272,N_17885);
nand U25995 (N_25995,N_12073,N_12033);
or U25996 (N_25996,N_16043,N_15749);
xnor U25997 (N_25997,N_11960,N_13836);
xnor U25998 (N_25998,N_18158,N_16943);
nor U25999 (N_25999,N_18624,N_14551);
xnor U26000 (N_26000,N_10829,N_10869);
xnor U26001 (N_26001,N_18443,N_13781);
and U26002 (N_26002,N_17542,N_11839);
nor U26003 (N_26003,N_15145,N_18201);
and U26004 (N_26004,N_10985,N_14841);
or U26005 (N_26005,N_10770,N_14209);
nand U26006 (N_26006,N_17859,N_10535);
nor U26007 (N_26007,N_15502,N_16128);
xor U26008 (N_26008,N_16137,N_15659);
xor U26009 (N_26009,N_13160,N_15398);
xor U26010 (N_26010,N_19131,N_19968);
or U26011 (N_26011,N_17383,N_16474);
nor U26012 (N_26012,N_17973,N_18257);
and U26013 (N_26013,N_14281,N_11918);
or U26014 (N_26014,N_10236,N_16511);
or U26015 (N_26015,N_12388,N_11568);
nor U26016 (N_26016,N_13551,N_10275);
or U26017 (N_26017,N_10284,N_12912);
nand U26018 (N_26018,N_15292,N_18969);
xnor U26019 (N_26019,N_16466,N_16894);
xnor U26020 (N_26020,N_13025,N_13145);
nand U26021 (N_26021,N_19968,N_13613);
or U26022 (N_26022,N_14740,N_13636);
and U26023 (N_26023,N_12483,N_10898);
nand U26024 (N_26024,N_14459,N_18852);
and U26025 (N_26025,N_10275,N_15749);
nand U26026 (N_26026,N_11610,N_15009);
nor U26027 (N_26027,N_15504,N_14701);
nor U26028 (N_26028,N_11151,N_17532);
or U26029 (N_26029,N_11253,N_10789);
nand U26030 (N_26030,N_11792,N_10922);
nor U26031 (N_26031,N_10853,N_14321);
or U26032 (N_26032,N_13461,N_16454);
and U26033 (N_26033,N_11466,N_11347);
xnor U26034 (N_26034,N_11513,N_13144);
nand U26035 (N_26035,N_10812,N_15258);
xor U26036 (N_26036,N_11934,N_17072);
nor U26037 (N_26037,N_19891,N_18612);
nand U26038 (N_26038,N_13462,N_19083);
nor U26039 (N_26039,N_13796,N_15965);
and U26040 (N_26040,N_14812,N_11366);
nor U26041 (N_26041,N_15124,N_17274);
nor U26042 (N_26042,N_16387,N_13391);
nand U26043 (N_26043,N_14104,N_12532);
xor U26044 (N_26044,N_18782,N_15852);
and U26045 (N_26045,N_13185,N_19444);
and U26046 (N_26046,N_19369,N_12517);
nand U26047 (N_26047,N_13616,N_13722);
xor U26048 (N_26048,N_10091,N_12729);
nand U26049 (N_26049,N_13319,N_12340);
or U26050 (N_26050,N_10007,N_11773);
and U26051 (N_26051,N_17724,N_14840);
or U26052 (N_26052,N_19500,N_19130);
nand U26053 (N_26053,N_13948,N_17703);
nor U26054 (N_26054,N_14165,N_10297);
and U26055 (N_26055,N_16906,N_18311);
and U26056 (N_26056,N_18606,N_13268);
nand U26057 (N_26057,N_15228,N_10034);
or U26058 (N_26058,N_14100,N_13189);
nand U26059 (N_26059,N_19877,N_15950);
and U26060 (N_26060,N_14194,N_14578);
and U26061 (N_26061,N_19084,N_17273);
nor U26062 (N_26062,N_10931,N_10096);
or U26063 (N_26063,N_16100,N_12136);
nor U26064 (N_26064,N_12068,N_15155);
and U26065 (N_26065,N_12596,N_12398);
nor U26066 (N_26066,N_11879,N_18831);
xnor U26067 (N_26067,N_11797,N_15095);
and U26068 (N_26068,N_18433,N_10005);
nand U26069 (N_26069,N_17406,N_19681);
nand U26070 (N_26070,N_10012,N_11986);
or U26071 (N_26071,N_19025,N_12537);
xor U26072 (N_26072,N_10877,N_16376);
nor U26073 (N_26073,N_17038,N_11748);
or U26074 (N_26074,N_12300,N_16753);
or U26075 (N_26075,N_14076,N_16497);
nand U26076 (N_26076,N_16167,N_13424);
nand U26077 (N_26077,N_17980,N_12971);
nor U26078 (N_26078,N_12860,N_11603);
nor U26079 (N_26079,N_16946,N_12463);
or U26080 (N_26080,N_16126,N_12930);
nand U26081 (N_26081,N_16053,N_14425);
nor U26082 (N_26082,N_19872,N_17039);
or U26083 (N_26083,N_12313,N_10126);
nand U26084 (N_26084,N_16973,N_11293);
nor U26085 (N_26085,N_19988,N_15810);
nor U26086 (N_26086,N_16785,N_14311);
xnor U26087 (N_26087,N_10337,N_11613);
nand U26088 (N_26088,N_14218,N_18605);
nor U26089 (N_26089,N_11998,N_13743);
and U26090 (N_26090,N_10448,N_12262);
nor U26091 (N_26091,N_13330,N_13064);
xnor U26092 (N_26092,N_13493,N_18898);
or U26093 (N_26093,N_18958,N_12365);
xnor U26094 (N_26094,N_17654,N_16604);
nor U26095 (N_26095,N_17990,N_16110);
and U26096 (N_26096,N_19941,N_18604);
nand U26097 (N_26097,N_12686,N_18866);
xor U26098 (N_26098,N_12340,N_12556);
nand U26099 (N_26099,N_18659,N_14902);
xor U26100 (N_26100,N_14644,N_10954);
and U26101 (N_26101,N_13529,N_13356);
xnor U26102 (N_26102,N_13680,N_10812);
nor U26103 (N_26103,N_16544,N_13197);
and U26104 (N_26104,N_16632,N_10441);
xor U26105 (N_26105,N_12253,N_12708);
nand U26106 (N_26106,N_15309,N_15756);
and U26107 (N_26107,N_10762,N_15794);
xnor U26108 (N_26108,N_17186,N_10768);
and U26109 (N_26109,N_13307,N_16979);
and U26110 (N_26110,N_19988,N_19548);
nor U26111 (N_26111,N_18614,N_14575);
xnor U26112 (N_26112,N_17129,N_14963);
and U26113 (N_26113,N_11128,N_18419);
xor U26114 (N_26114,N_10487,N_18975);
or U26115 (N_26115,N_16550,N_15492);
xnor U26116 (N_26116,N_19488,N_12890);
xnor U26117 (N_26117,N_15174,N_11268);
nor U26118 (N_26118,N_14037,N_10299);
or U26119 (N_26119,N_16393,N_10547);
nand U26120 (N_26120,N_14878,N_13633);
nor U26121 (N_26121,N_17194,N_19704);
xor U26122 (N_26122,N_13314,N_17148);
nor U26123 (N_26123,N_13232,N_14754);
nand U26124 (N_26124,N_16491,N_15542);
and U26125 (N_26125,N_17686,N_17736);
xnor U26126 (N_26126,N_16172,N_15452);
nor U26127 (N_26127,N_13975,N_13799);
and U26128 (N_26128,N_13833,N_14574);
and U26129 (N_26129,N_16777,N_17201);
or U26130 (N_26130,N_16628,N_10778);
and U26131 (N_26131,N_10872,N_10378);
and U26132 (N_26132,N_11730,N_16621);
or U26133 (N_26133,N_14887,N_10578);
xor U26134 (N_26134,N_15984,N_18293);
or U26135 (N_26135,N_18185,N_17270);
nand U26136 (N_26136,N_16826,N_19027);
nor U26137 (N_26137,N_18932,N_13911);
or U26138 (N_26138,N_14371,N_13199);
nor U26139 (N_26139,N_16864,N_12986);
nor U26140 (N_26140,N_16486,N_15306);
nand U26141 (N_26141,N_13070,N_19046);
nor U26142 (N_26142,N_17621,N_17684);
nand U26143 (N_26143,N_13868,N_12034);
nand U26144 (N_26144,N_11123,N_16040);
nor U26145 (N_26145,N_14622,N_12447);
nor U26146 (N_26146,N_16864,N_10147);
xor U26147 (N_26147,N_18853,N_13773);
nand U26148 (N_26148,N_16267,N_19967);
nor U26149 (N_26149,N_13168,N_19524);
and U26150 (N_26150,N_19065,N_13850);
and U26151 (N_26151,N_17509,N_19203);
xor U26152 (N_26152,N_18597,N_14938);
or U26153 (N_26153,N_16568,N_15571);
nand U26154 (N_26154,N_14439,N_18039);
or U26155 (N_26155,N_15791,N_15001);
nand U26156 (N_26156,N_11647,N_15624);
nand U26157 (N_26157,N_17758,N_15973);
nand U26158 (N_26158,N_15302,N_13188);
nor U26159 (N_26159,N_11028,N_17568);
nor U26160 (N_26160,N_18457,N_12549);
or U26161 (N_26161,N_12651,N_12300);
nor U26162 (N_26162,N_13101,N_17429);
and U26163 (N_26163,N_12800,N_12602);
and U26164 (N_26164,N_13672,N_14458);
or U26165 (N_26165,N_10042,N_14902);
nor U26166 (N_26166,N_13468,N_12655);
or U26167 (N_26167,N_14581,N_17264);
or U26168 (N_26168,N_19987,N_13781);
xor U26169 (N_26169,N_15800,N_14154);
nor U26170 (N_26170,N_19218,N_13199);
xor U26171 (N_26171,N_17993,N_15412);
or U26172 (N_26172,N_13035,N_10442);
nor U26173 (N_26173,N_14011,N_14466);
nor U26174 (N_26174,N_18584,N_14002);
nor U26175 (N_26175,N_17014,N_15543);
nor U26176 (N_26176,N_12096,N_13509);
or U26177 (N_26177,N_19497,N_10975);
xor U26178 (N_26178,N_13273,N_18397);
and U26179 (N_26179,N_10703,N_18289);
and U26180 (N_26180,N_16696,N_18340);
xor U26181 (N_26181,N_14806,N_13750);
nor U26182 (N_26182,N_17505,N_10088);
and U26183 (N_26183,N_15222,N_15442);
nor U26184 (N_26184,N_12973,N_17913);
and U26185 (N_26185,N_19455,N_18163);
xnor U26186 (N_26186,N_14268,N_13113);
nand U26187 (N_26187,N_15996,N_14831);
or U26188 (N_26188,N_19052,N_18995);
or U26189 (N_26189,N_14415,N_16033);
nor U26190 (N_26190,N_15642,N_11916);
or U26191 (N_26191,N_10457,N_19961);
nand U26192 (N_26192,N_15116,N_12525);
and U26193 (N_26193,N_18345,N_15097);
and U26194 (N_26194,N_19752,N_10244);
xnor U26195 (N_26195,N_12255,N_15865);
and U26196 (N_26196,N_19149,N_15156);
or U26197 (N_26197,N_14623,N_15940);
and U26198 (N_26198,N_17738,N_10120);
nor U26199 (N_26199,N_19867,N_17501);
nand U26200 (N_26200,N_17060,N_13771);
nor U26201 (N_26201,N_14632,N_12119);
xnor U26202 (N_26202,N_16944,N_10003);
nand U26203 (N_26203,N_13581,N_18602);
nand U26204 (N_26204,N_19650,N_11598);
and U26205 (N_26205,N_14714,N_17794);
or U26206 (N_26206,N_16814,N_17504);
and U26207 (N_26207,N_13604,N_12946);
and U26208 (N_26208,N_12841,N_16106);
xor U26209 (N_26209,N_17098,N_19060);
or U26210 (N_26210,N_13690,N_18895);
xnor U26211 (N_26211,N_10876,N_10766);
nor U26212 (N_26212,N_10531,N_17592);
and U26213 (N_26213,N_14936,N_18682);
xor U26214 (N_26214,N_12865,N_12423);
or U26215 (N_26215,N_13744,N_10830);
nand U26216 (N_26216,N_18047,N_18367);
nand U26217 (N_26217,N_17791,N_19864);
or U26218 (N_26218,N_14914,N_11543);
or U26219 (N_26219,N_14453,N_18247);
nand U26220 (N_26220,N_11935,N_13745);
and U26221 (N_26221,N_10303,N_10215);
xor U26222 (N_26222,N_15621,N_13167);
or U26223 (N_26223,N_11166,N_17274);
nor U26224 (N_26224,N_18591,N_15294);
xor U26225 (N_26225,N_11689,N_17276);
nor U26226 (N_26226,N_15920,N_16693);
nor U26227 (N_26227,N_17081,N_11323);
nor U26228 (N_26228,N_11018,N_10821);
and U26229 (N_26229,N_19833,N_13519);
nor U26230 (N_26230,N_15312,N_12096);
nand U26231 (N_26231,N_15981,N_19337);
nand U26232 (N_26232,N_12740,N_19545);
nand U26233 (N_26233,N_17535,N_14726);
or U26234 (N_26234,N_13196,N_13182);
nor U26235 (N_26235,N_19460,N_18407);
xor U26236 (N_26236,N_11086,N_14688);
nor U26237 (N_26237,N_10388,N_19066);
and U26238 (N_26238,N_14916,N_18046);
or U26239 (N_26239,N_17855,N_18250);
nor U26240 (N_26240,N_10307,N_18755);
or U26241 (N_26241,N_17891,N_15750);
and U26242 (N_26242,N_14294,N_14171);
xor U26243 (N_26243,N_18164,N_13251);
or U26244 (N_26244,N_13571,N_15193);
xnor U26245 (N_26245,N_17568,N_18374);
nor U26246 (N_26246,N_12635,N_10104);
xnor U26247 (N_26247,N_18057,N_16318);
or U26248 (N_26248,N_18139,N_15483);
nor U26249 (N_26249,N_15174,N_16839);
nor U26250 (N_26250,N_12961,N_13286);
or U26251 (N_26251,N_12387,N_13935);
and U26252 (N_26252,N_13975,N_12750);
xnor U26253 (N_26253,N_10881,N_16354);
nor U26254 (N_26254,N_17881,N_14822);
and U26255 (N_26255,N_13330,N_11654);
or U26256 (N_26256,N_10119,N_10849);
nand U26257 (N_26257,N_10164,N_14547);
nor U26258 (N_26258,N_11286,N_13523);
xor U26259 (N_26259,N_11258,N_10227);
nand U26260 (N_26260,N_15634,N_19545);
or U26261 (N_26261,N_16679,N_19840);
and U26262 (N_26262,N_13556,N_15957);
nor U26263 (N_26263,N_14004,N_10982);
nand U26264 (N_26264,N_12799,N_10169);
nand U26265 (N_26265,N_14937,N_17330);
xnor U26266 (N_26266,N_15161,N_16840);
and U26267 (N_26267,N_12520,N_10873);
nor U26268 (N_26268,N_16142,N_17770);
xnor U26269 (N_26269,N_10477,N_13850);
and U26270 (N_26270,N_17791,N_14828);
or U26271 (N_26271,N_10851,N_13726);
nor U26272 (N_26272,N_14199,N_10218);
and U26273 (N_26273,N_13405,N_19631);
nand U26274 (N_26274,N_12879,N_13014);
nand U26275 (N_26275,N_16318,N_19190);
or U26276 (N_26276,N_14270,N_10143);
xnor U26277 (N_26277,N_18029,N_14359);
nor U26278 (N_26278,N_14203,N_17941);
xnor U26279 (N_26279,N_11139,N_18616);
and U26280 (N_26280,N_17171,N_12640);
xor U26281 (N_26281,N_10551,N_19501);
or U26282 (N_26282,N_14226,N_18669);
xor U26283 (N_26283,N_19113,N_11156);
nand U26284 (N_26284,N_10465,N_16446);
nand U26285 (N_26285,N_18749,N_14773);
nor U26286 (N_26286,N_14101,N_15314);
nand U26287 (N_26287,N_12178,N_18512);
and U26288 (N_26288,N_13256,N_14642);
nand U26289 (N_26289,N_19070,N_11310);
or U26290 (N_26290,N_18140,N_18768);
nand U26291 (N_26291,N_16874,N_16968);
or U26292 (N_26292,N_12418,N_18435);
and U26293 (N_26293,N_18189,N_12650);
or U26294 (N_26294,N_15921,N_11730);
and U26295 (N_26295,N_14828,N_17106);
and U26296 (N_26296,N_10141,N_13762);
and U26297 (N_26297,N_14929,N_12054);
xnor U26298 (N_26298,N_14507,N_10943);
xor U26299 (N_26299,N_10651,N_13411);
nor U26300 (N_26300,N_10052,N_13603);
or U26301 (N_26301,N_12580,N_13201);
and U26302 (N_26302,N_14780,N_11385);
xor U26303 (N_26303,N_19950,N_18532);
xnor U26304 (N_26304,N_18686,N_14184);
nand U26305 (N_26305,N_18489,N_10609);
nor U26306 (N_26306,N_11678,N_12392);
or U26307 (N_26307,N_10639,N_13198);
xor U26308 (N_26308,N_13213,N_14421);
xor U26309 (N_26309,N_11459,N_18039);
nor U26310 (N_26310,N_18310,N_18183);
or U26311 (N_26311,N_13969,N_11532);
or U26312 (N_26312,N_14229,N_13670);
nand U26313 (N_26313,N_12112,N_10559);
xnor U26314 (N_26314,N_13630,N_19987);
and U26315 (N_26315,N_15468,N_18818);
nand U26316 (N_26316,N_18789,N_13743);
and U26317 (N_26317,N_17567,N_12046);
nor U26318 (N_26318,N_13982,N_10317);
xnor U26319 (N_26319,N_14128,N_16591);
nor U26320 (N_26320,N_16652,N_13088);
nor U26321 (N_26321,N_15917,N_10324);
or U26322 (N_26322,N_14732,N_10109);
or U26323 (N_26323,N_13698,N_13080);
or U26324 (N_26324,N_10096,N_13834);
or U26325 (N_26325,N_16242,N_13228);
or U26326 (N_26326,N_19429,N_13392);
or U26327 (N_26327,N_15002,N_10875);
nand U26328 (N_26328,N_13914,N_17125);
xor U26329 (N_26329,N_12043,N_11832);
and U26330 (N_26330,N_17119,N_12018);
xor U26331 (N_26331,N_17294,N_15634);
nor U26332 (N_26332,N_10316,N_15751);
nor U26333 (N_26333,N_15010,N_16971);
nor U26334 (N_26334,N_19373,N_10932);
nor U26335 (N_26335,N_17894,N_13349);
xnor U26336 (N_26336,N_15099,N_12794);
nand U26337 (N_26337,N_11920,N_12507);
xor U26338 (N_26338,N_12822,N_12334);
xnor U26339 (N_26339,N_12878,N_12439);
or U26340 (N_26340,N_14891,N_16946);
xnor U26341 (N_26341,N_12687,N_18417);
xor U26342 (N_26342,N_11330,N_12052);
nor U26343 (N_26343,N_13782,N_11718);
xor U26344 (N_26344,N_17072,N_13731);
xnor U26345 (N_26345,N_18571,N_12058);
or U26346 (N_26346,N_12353,N_11580);
or U26347 (N_26347,N_15717,N_15463);
nor U26348 (N_26348,N_18913,N_14659);
and U26349 (N_26349,N_12531,N_12297);
nand U26350 (N_26350,N_13918,N_15593);
or U26351 (N_26351,N_11135,N_12930);
nor U26352 (N_26352,N_12082,N_11610);
xor U26353 (N_26353,N_15229,N_13190);
and U26354 (N_26354,N_13991,N_15954);
nand U26355 (N_26355,N_16288,N_14016);
nor U26356 (N_26356,N_10306,N_16446);
nor U26357 (N_26357,N_17289,N_11073);
nor U26358 (N_26358,N_11715,N_10419);
nor U26359 (N_26359,N_19034,N_15042);
and U26360 (N_26360,N_14600,N_19505);
nand U26361 (N_26361,N_10365,N_11132);
xnor U26362 (N_26362,N_18214,N_14250);
or U26363 (N_26363,N_17311,N_18243);
nor U26364 (N_26364,N_17746,N_12142);
and U26365 (N_26365,N_12744,N_18337);
nor U26366 (N_26366,N_16674,N_16593);
nand U26367 (N_26367,N_11677,N_15902);
nor U26368 (N_26368,N_10259,N_16776);
and U26369 (N_26369,N_15330,N_16126);
nand U26370 (N_26370,N_11797,N_10034);
nor U26371 (N_26371,N_12715,N_17501);
xor U26372 (N_26372,N_17335,N_12614);
nor U26373 (N_26373,N_16171,N_14976);
and U26374 (N_26374,N_14311,N_12707);
xor U26375 (N_26375,N_10564,N_14582);
xor U26376 (N_26376,N_17811,N_10928);
nand U26377 (N_26377,N_19203,N_12121);
xor U26378 (N_26378,N_10466,N_13729);
or U26379 (N_26379,N_11719,N_12933);
or U26380 (N_26380,N_17033,N_15697);
xor U26381 (N_26381,N_11804,N_19354);
and U26382 (N_26382,N_19132,N_17685);
and U26383 (N_26383,N_16936,N_19189);
nand U26384 (N_26384,N_10746,N_14052);
nor U26385 (N_26385,N_16974,N_18375);
and U26386 (N_26386,N_10320,N_18701);
nand U26387 (N_26387,N_18819,N_18140);
or U26388 (N_26388,N_14088,N_15206);
nor U26389 (N_26389,N_19792,N_12526);
nor U26390 (N_26390,N_18662,N_16461);
nor U26391 (N_26391,N_18153,N_17449);
xnor U26392 (N_26392,N_17660,N_18401);
xor U26393 (N_26393,N_15203,N_18259);
nand U26394 (N_26394,N_15890,N_19487);
nor U26395 (N_26395,N_18106,N_19666);
nor U26396 (N_26396,N_15513,N_11789);
nor U26397 (N_26397,N_13917,N_14158);
xor U26398 (N_26398,N_17817,N_14503);
or U26399 (N_26399,N_17354,N_16255);
xor U26400 (N_26400,N_15556,N_18028);
nor U26401 (N_26401,N_16245,N_14152);
and U26402 (N_26402,N_17318,N_11063);
nand U26403 (N_26403,N_15093,N_11775);
or U26404 (N_26404,N_15645,N_12944);
or U26405 (N_26405,N_17610,N_17188);
xnor U26406 (N_26406,N_16678,N_15622);
xor U26407 (N_26407,N_17471,N_11653);
or U26408 (N_26408,N_12026,N_12003);
or U26409 (N_26409,N_19196,N_11383);
xor U26410 (N_26410,N_10696,N_17391);
nand U26411 (N_26411,N_19172,N_15382);
and U26412 (N_26412,N_13691,N_19012);
nor U26413 (N_26413,N_11676,N_19830);
and U26414 (N_26414,N_19103,N_19554);
or U26415 (N_26415,N_12732,N_13367);
nand U26416 (N_26416,N_19470,N_17787);
xor U26417 (N_26417,N_14383,N_18347);
and U26418 (N_26418,N_17337,N_11818);
or U26419 (N_26419,N_11175,N_15789);
nor U26420 (N_26420,N_13087,N_15385);
nor U26421 (N_26421,N_14838,N_11942);
nor U26422 (N_26422,N_14088,N_15165);
xor U26423 (N_26423,N_17961,N_10440);
nand U26424 (N_26424,N_13819,N_17402);
and U26425 (N_26425,N_10346,N_13071);
or U26426 (N_26426,N_16104,N_14075);
nand U26427 (N_26427,N_19609,N_17641);
or U26428 (N_26428,N_13802,N_12318);
nor U26429 (N_26429,N_10735,N_14534);
and U26430 (N_26430,N_17769,N_11393);
and U26431 (N_26431,N_19477,N_10079);
and U26432 (N_26432,N_13362,N_12233);
xor U26433 (N_26433,N_17847,N_18826);
nor U26434 (N_26434,N_10074,N_11752);
and U26435 (N_26435,N_10995,N_13630);
xnor U26436 (N_26436,N_14404,N_14659);
xor U26437 (N_26437,N_12554,N_12828);
and U26438 (N_26438,N_12992,N_11019);
or U26439 (N_26439,N_13596,N_11767);
nand U26440 (N_26440,N_15807,N_17595);
nand U26441 (N_26441,N_13979,N_14162);
nand U26442 (N_26442,N_12269,N_12225);
and U26443 (N_26443,N_16607,N_15300);
or U26444 (N_26444,N_12487,N_12527);
nand U26445 (N_26445,N_15480,N_10021);
and U26446 (N_26446,N_15543,N_14995);
nand U26447 (N_26447,N_11533,N_14535);
nor U26448 (N_26448,N_12536,N_16826);
and U26449 (N_26449,N_18096,N_12513);
or U26450 (N_26450,N_15098,N_18730);
nor U26451 (N_26451,N_16376,N_19953);
or U26452 (N_26452,N_17344,N_19720);
or U26453 (N_26453,N_15163,N_13291);
and U26454 (N_26454,N_11787,N_10140);
and U26455 (N_26455,N_12356,N_15950);
xnor U26456 (N_26456,N_13479,N_11257);
nor U26457 (N_26457,N_12066,N_12289);
xnor U26458 (N_26458,N_15242,N_14845);
nor U26459 (N_26459,N_14735,N_12927);
or U26460 (N_26460,N_16158,N_10669);
and U26461 (N_26461,N_12722,N_16928);
nor U26462 (N_26462,N_10441,N_17078);
nor U26463 (N_26463,N_10373,N_15389);
xor U26464 (N_26464,N_17582,N_15587);
or U26465 (N_26465,N_16468,N_11318);
nor U26466 (N_26466,N_15679,N_10317);
nand U26467 (N_26467,N_12735,N_19027);
nand U26468 (N_26468,N_13495,N_15657);
and U26469 (N_26469,N_19062,N_16074);
or U26470 (N_26470,N_14282,N_12740);
nand U26471 (N_26471,N_19091,N_10425);
nand U26472 (N_26472,N_13644,N_11529);
or U26473 (N_26473,N_19014,N_17258);
nand U26474 (N_26474,N_19935,N_18429);
and U26475 (N_26475,N_17896,N_12419);
xnor U26476 (N_26476,N_12510,N_16990);
and U26477 (N_26477,N_18487,N_16316);
or U26478 (N_26478,N_14064,N_12975);
xnor U26479 (N_26479,N_10699,N_19563);
nor U26480 (N_26480,N_18194,N_18383);
nor U26481 (N_26481,N_16876,N_18449);
xor U26482 (N_26482,N_10700,N_16549);
xor U26483 (N_26483,N_19130,N_12805);
xnor U26484 (N_26484,N_16722,N_10391);
and U26485 (N_26485,N_10920,N_15586);
nand U26486 (N_26486,N_17881,N_13861);
nor U26487 (N_26487,N_11976,N_19778);
or U26488 (N_26488,N_14585,N_13373);
nor U26489 (N_26489,N_13108,N_10412);
xor U26490 (N_26490,N_11010,N_16474);
xnor U26491 (N_26491,N_15652,N_17930);
or U26492 (N_26492,N_19482,N_19194);
nor U26493 (N_26493,N_13373,N_15669);
and U26494 (N_26494,N_18037,N_16820);
or U26495 (N_26495,N_16219,N_17373);
nor U26496 (N_26496,N_12935,N_16234);
xnor U26497 (N_26497,N_18397,N_16010);
and U26498 (N_26498,N_19698,N_17154);
xnor U26499 (N_26499,N_19042,N_17817);
nand U26500 (N_26500,N_11548,N_13134);
nor U26501 (N_26501,N_16794,N_18673);
and U26502 (N_26502,N_11241,N_12301);
and U26503 (N_26503,N_17092,N_13453);
nand U26504 (N_26504,N_17425,N_10102);
nand U26505 (N_26505,N_15904,N_10137);
xnor U26506 (N_26506,N_16337,N_18606);
nand U26507 (N_26507,N_18115,N_18634);
nand U26508 (N_26508,N_10744,N_16150);
nand U26509 (N_26509,N_15188,N_16259);
xor U26510 (N_26510,N_11736,N_14293);
nor U26511 (N_26511,N_13432,N_16403);
or U26512 (N_26512,N_13313,N_10284);
nand U26513 (N_26513,N_12146,N_18956);
nor U26514 (N_26514,N_12818,N_13536);
xnor U26515 (N_26515,N_17630,N_16013);
and U26516 (N_26516,N_13105,N_19042);
or U26517 (N_26517,N_11854,N_14584);
and U26518 (N_26518,N_16638,N_17970);
and U26519 (N_26519,N_10381,N_17153);
nor U26520 (N_26520,N_12233,N_19734);
and U26521 (N_26521,N_17162,N_12402);
or U26522 (N_26522,N_14387,N_11612);
and U26523 (N_26523,N_11673,N_12639);
and U26524 (N_26524,N_12038,N_11926);
nand U26525 (N_26525,N_10213,N_11685);
nand U26526 (N_26526,N_15720,N_19283);
and U26527 (N_26527,N_19612,N_10261);
or U26528 (N_26528,N_14917,N_17832);
xor U26529 (N_26529,N_13030,N_11855);
nor U26530 (N_26530,N_14916,N_19429);
nand U26531 (N_26531,N_15308,N_12787);
nor U26532 (N_26532,N_14843,N_12094);
nor U26533 (N_26533,N_12472,N_15297);
or U26534 (N_26534,N_14999,N_18901);
nor U26535 (N_26535,N_18775,N_12508);
nor U26536 (N_26536,N_14737,N_15127);
and U26537 (N_26537,N_15826,N_18268);
nor U26538 (N_26538,N_11953,N_15370);
xor U26539 (N_26539,N_19779,N_12806);
nor U26540 (N_26540,N_10811,N_11023);
nor U26541 (N_26541,N_13390,N_17772);
nor U26542 (N_26542,N_14239,N_17403);
nor U26543 (N_26543,N_16524,N_17657);
nor U26544 (N_26544,N_15917,N_10665);
nor U26545 (N_26545,N_18624,N_12414);
xnor U26546 (N_26546,N_10819,N_19048);
nor U26547 (N_26547,N_18391,N_15030);
xor U26548 (N_26548,N_16955,N_17464);
or U26549 (N_26549,N_11049,N_19558);
xnor U26550 (N_26550,N_16664,N_10413);
nand U26551 (N_26551,N_11148,N_13031);
or U26552 (N_26552,N_10790,N_13008);
xnor U26553 (N_26553,N_16961,N_11764);
nand U26554 (N_26554,N_15845,N_11769);
or U26555 (N_26555,N_16548,N_14428);
nor U26556 (N_26556,N_11364,N_19613);
nand U26557 (N_26557,N_17537,N_10676);
xor U26558 (N_26558,N_15638,N_15681);
and U26559 (N_26559,N_19026,N_17363);
nor U26560 (N_26560,N_11919,N_12478);
and U26561 (N_26561,N_13145,N_17096);
nand U26562 (N_26562,N_17011,N_12314);
and U26563 (N_26563,N_14454,N_14248);
nand U26564 (N_26564,N_16884,N_14165);
and U26565 (N_26565,N_19789,N_13682);
and U26566 (N_26566,N_11216,N_14887);
nand U26567 (N_26567,N_10061,N_16878);
and U26568 (N_26568,N_19641,N_16205);
and U26569 (N_26569,N_14540,N_12766);
nand U26570 (N_26570,N_16255,N_14157);
nor U26571 (N_26571,N_13618,N_18309);
or U26572 (N_26572,N_13539,N_13672);
or U26573 (N_26573,N_18812,N_11308);
nand U26574 (N_26574,N_13286,N_19901);
xnor U26575 (N_26575,N_15406,N_16143);
nand U26576 (N_26576,N_16011,N_12589);
nand U26577 (N_26577,N_15218,N_10271);
and U26578 (N_26578,N_17783,N_15790);
nand U26579 (N_26579,N_19100,N_18769);
and U26580 (N_26580,N_12526,N_17479);
nand U26581 (N_26581,N_11692,N_18124);
nand U26582 (N_26582,N_11358,N_12768);
nor U26583 (N_26583,N_11822,N_18634);
or U26584 (N_26584,N_14099,N_19930);
and U26585 (N_26585,N_18666,N_12422);
or U26586 (N_26586,N_12972,N_16744);
xor U26587 (N_26587,N_13968,N_15024);
or U26588 (N_26588,N_19700,N_18823);
nand U26589 (N_26589,N_12138,N_18018);
and U26590 (N_26590,N_17891,N_17286);
and U26591 (N_26591,N_15759,N_19645);
or U26592 (N_26592,N_14697,N_13466);
nand U26593 (N_26593,N_16515,N_19118);
nor U26594 (N_26594,N_15772,N_14240);
xnor U26595 (N_26595,N_19083,N_13114);
and U26596 (N_26596,N_10844,N_11209);
or U26597 (N_26597,N_19876,N_16137);
nor U26598 (N_26598,N_14096,N_15180);
nand U26599 (N_26599,N_17161,N_12907);
nand U26600 (N_26600,N_19386,N_18800);
xor U26601 (N_26601,N_16292,N_11594);
and U26602 (N_26602,N_19004,N_17198);
nor U26603 (N_26603,N_14706,N_15342);
or U26604 (N_26604,N_17724,N_13855);
nor U26605 (N_26605,N_14831,N_12990);
nor U26606 (N_26606,N_19422,N_19836);
or U26607 (N_26607,N_10834,N_12029);
xnor U26608 (N_26608,N_14465,N_10121);
and U26609 (N_26609,N_10956,N_10714);
and U26610 (N_26610,N_16737,N_12876);
xor U26611 (N_26611,N_16610,N_18438);
nor U26612 (N_26612,N_16489,N_12272);
nand U26613 (N_26613,N_14656,N_17181);
or U26614 (N_26614,N_10723,N_11901);
nand U26615 (N_26615,N_13430,N_15716);
nor U26616 (N_26616,N_10384,N_10401);
or U26617 (N_26617,N_17872,N_10387);
or U26618 (N_26618,N_14876,N_11703);
xor U26619 (N_26619,N_15635,N_15707);
nor U26620 (N_26620,N_17326,N_11773);
xor U26621 (N_26621,N_17738,N_10919);
and U26622 (N_26622,N_11377,N_10714);
xor U26623 (N_26623,N_12594,N_16187);
xor U26624 (N_26624,N_16167,N_10803);
or U26625 (N_26625,N_13519,N_18503);
nor U26626 (N_26626,N_15938,N_17133);
and U26627 (N_26627,N_16045,N_18704);
nand U26628 (N_26628,N_19063,N_17757);
or U26629 (N_26629,N_15540,N_14836);
nand U26630 (N_26630,N_13812,N_15930);
nand U26631 (N_26631,N_12614,N_10330);
or U26632 (N_26632,N_15154,N_15169);
and U26633 (N_26633,N_11407,N_11128);
and U26634 (N_26634,N_19589,N_17280);
nand U26635 (N_26635,N_11173,N_15046);
and U26636 (N_26636,N_16770,N_19658);
and U26637 (N_26637,N_14326,N_16100);
nand U26638 (N_26638,N_10611,N_12170);
nor U26639 (N_26639,N_11277,N_16866);
nor U26640 (N_26640,N_11339,N_14812);
or U26641 (N_26641,N_12280,N_11402);
xor U26642 (N_26642,N_12599,N_13939);
and U26643 (N_26643,N_11130,N_15477);
nor U26644 (N_26644,N_19189,N_13403);
nor U26645 (N_26645,N_13690,N_14599);
xor U26646 (N_26646,N_12155,N_17906);
nor U26647 (N_26647,N_12404,N_13380);
xor U26648 (N_26648,N_16369,N_17941);
and U26649 (N_26649,N_15858,N_10232);
nor U26650 (N_26650,N_11941,N_16117);
nor U26651 (N_26651,N_13842,N_15042);
nor U26652 (N_26652,N_11331,N_11113);
nand U26653 (N_26653,N_11448,N_16188);
and U26654 (N_26654,N_14880,N_16656);
xor U26655 (N_26655,N_16520,N_14188);
nor U26656 (N_26656,N_13745,N_18559);
or U26657 (N_26657,N_12862,N_12938);
and U26658 (N_26658,N_15853,N_13869);
nand U26659 (N_26659,N_17403,N_13405);
or U26660 (N_26660,N_14811,N_19278);
nor U26661 (N_26661,N_13895,N_14846);
nor U26662 (N_26662,N_14774,N_19343);
nand U26663 (N_26663,N_13978,N_10527);
nand U26664 (N_26664,N_15844,N_17883);
or U26665 (N_26665,N_14887,N_19999);
or U26666 (N_26666,N_13063,N_13661);
xnor U26667 (N_26667,N_17215,N_15260);
or U26668 (N_26668,N_19576,N_15534);
xor U26669 (N_26669,N_12282,N_10678);
and U26670 (N_26670,N_17571,N_18195);
nor U26671 (N_26671,N_10470,N_12656);
nand U26672 (N_26672,N_10158,N_12586);
or U26673 (N_26673,N_12161,N_13725);
or U26674 (N_26674,N_17321,N_19752);
and U26675 (N_26675,N_13455,N_12592);
nand U26676 (N_26676,N_19529,N_14058);
nand U26677 (N_26677,N_15867,N_17268);
or U26678 (N_26678,N_12855,N_11297);
and U26679 (N_26679,N_19703,N_11902);
nor U26680 (N_26680,N_11728,N_17030);
and U26681 (N_26681,N_12422,N_14512);
or U26682 (N_26682,N_10215,N_10790);
nor U26683 (N_26683,N_13896,N_12847);
nor U26684 (N_26684,N_15140,N_17130);
nor U26685 (N_26685,N_13989,N_17035);
and U26686 (N_26686,N_11405,N_12689);
or U26687 (N_26687,N_14521,N_12618);
nand U26688 (N_26688,N_10645,N_12240);
or U26689 (N_26689,N_11160,N_19751);
nor U26690 (N_26690,N_12846,N_11285);
or U26691 (N_26691,N_16592,N_15667);
and U26692 (N_26692,N_17422,N_12005);
xor U26693 (N_26693,N_13259,N_19180);
or U26694 (N_26694,N_14720,N_16921);
nor U26695 (N_26695,N_11399,N_11605);
nor U26696 (N_26696,N_18878,N_17501);
and U26697 (N_26697,N_12197,N_17902);
xnor U26698 (N_26698,N_15181,N_15800);
nor U26699 (N_26699,N_19102,N_16982);
or U26700 (N_26700,N_14524,N_13180);
nor U26701 (N_26701,N_19472,N_19633);
and U26702 (N_26702,N_15880,N_13541);
nor U26703 (N_26703,N_11078,N_19327);
xor U26704 (N_26704,N_16655,N_19497);
nor U26705 (N_26705,N_19287,N_15257);
nand U26706 (N_26706,N_10396,N_12878);
xor U26707 (N_26707,N_15365,N_17731);
xnor U26708 (N_26708,N_18892,N_17158);
and U26709 (N_26709,N_11612,N_17931);
and U26710 (N_26710,N_16227,N_14657);
xor U26711 (N_26711,N_10065,N_11578);
xnor U26712 (N_26712,N_10043,N_10572);
or U26713 (N_26713,N_14019,N_15993);
and U26714 (N_26714,N_11687,N_16390);
and U26715 (N_26715,N_15633,N_13418);
or U26716 (N_26716,N_19874,N_17963);
and U26717 (N_26717,N_14458,N_17645);
or U26718 (N_26718,N_17970,N_11432);
or U26719 (N_26719,N_15819,N_15554);
and U26720 (N_26720,N_17673,N_16824);
xnor U26721 (N_26721,N_11397,N_10185);
nand U26722 (N_26722,N_16697,N_16555);
nand U26723 (N_26723,N_13112,N_16819);
or U26724 (N_26724,N_11881,N_17732);
nand U26725 (N_26725,N_16741,N_13984);
nand U26726 (N_26726,N_11973,N_18972);
nand U26727 (N_26727,N_14943,N_11855);
and U26728 (N_26728,N_10038,N_10855);
xnor U26729 (N_26729,N_15218,N_19951);
or U26730 (N_26730,N_17859,N_11419);
or U26731 (N_26731,N_11793,N_18907);
nor U26732 (N_26732,N_11323,N_12193);
and U26733 (N_26733,N_15079,N_15104);
nand U26734 (N_26734,N_13092,N_10509);
xnor U26735 (N_26735,N_12425,N_12296);
nor U26736 (N_26736,N_15622,N_15162);
xnor U26737 (N_26737,N_19316,N_15310);
nor U26738 (N_26738,N_19625,N_13076);
or U26739 (N_26739,N_17571,N_11255);
and U26740 (N_26740,N_16983,N_10401);
xnor U26741 (N_26741,N_17324,N_16375);
and U26742 (N_26742,N_17269,N_10003);
nand U26743 (N_26743,N_19611,N_15422);
or U26744 (N_26744,N_18769,N_18036);
or U26745 (N_26745,N_12486,N_15474);
nand U26746 (N_26746,N_11319,N_17836);
nor U26747 (N_26747,N_14918,N_18462);
or U26748 (N_26748,N_16679,N_14568);
and U26749 (N_26749,N_12828,N_16122);
or U26750 (N_26750,N_11948,N_14108);
or U26751 (N_26751,N_15767,N_10100);
and U26752 (N_26752,N_17587,N_19473);
xnor U26753 (N_26753,N_12574,N_10717);
nand U26754 (N_26754,N_19230,N_11783);
nor U26755 (N_26755,N_11655,N_11241);
nand U26756 (N_26756,N_17684,N_14163);
nor U26757 (N_26757,N_19571,N_18415);
and U26758 (N_26758,N_12522,N_13388);
nand U26759 (N_26759,N_16983,N_14463);
xnor U26760 (N_26760,N_10112,N_13251);
xnor U26761 (N_26761,N_10094,N_11357);
xnor U26762 (N_26762,N_17727,N_11751);
and U26763 (N_26763,N_13179,N_12988);
nor U26764 (N_26764,N_10247,N_14766);
or U26765 (N_26765,N_18565,N_11300);
or U26766 (N_26766,N_11058,N_10215);
xnor U26767 (N_26767,N_17010,N_16567);
or U26768 (N_26768,N_18355,N_15576);
and U26769 (N_26769,N_12446,N_13884);
or U26770 (N_26770,N_16384,N_19944);
and U26771 (N_26771,N_15955,N_15563);
xnor U26772 (N_26772,N_15363,N_18855);
nand U26773 (N_26773,N_15790,N_17876);
or U26774 (N_26774,N_13109,N_12988);
or U26775 (N_26775,N_12491,N_17821);
and U26776 (N_26776,N_13255,N_13389);
or U26777 (N_26777,N_16416,N_18095);
nor U26778 (N_26778,N_16923,N_17366);
nor U26779 (N_26779,N_13851,N_14782);
and U26780 (N_26780,N_16924,N_16410);
and U26781 (N_26781,N_12062,N_14662);
and U26782 (N_26782,N_18978,N_10227);
xnor U26783 (N_26783,N_13129,N_14136);
nand U26784 (N_26784,N_14707,N_17558);
nor U26785 (N_26785,N_18487,N_19063);
nand U26786 (N_26786,N_17177,N_15962);
nand U26787 (N_26787,N_14777,N_19855);
xor U26788 (N_26788,N_18283,N_19634);
xnor U26789 (N_26789,N_18854,N_19604);
xnor U26790 (N_26790,N_19710,N_18027);
nand U26791 (N_26791,N_10620,N_17082);
nor U26792 (N_26792,N_15818,N_17473);
and U26793 (N_26793,N_13817,N_10432);
and U26794 (N_26794,N_19841,N_12922);
or U26795 (N_26795,N_14019,N_15238);
nand U26796 (N_26796,N_15023,N_11646);
nand U26797 (N_26797,N_10553,N_19436);
xor U26798 (N_26798,N_10606,N_13279);
xor U26799 (N_26799,N_12593,N_15496);
xor U26800 (N_26800,N_12108,N_14148);
and U26801 (N_26801,N_10186,N_13805);
and U26802 (N_26802,N_15824,N_10801);
xnor U26803 (N_26803,N_17156,N_18609);
nor U26804 (N_26804,N_11516,N_16730);
or U26805 (N_26805,N_18914,N_10136);
and U26806 (N_26806,N_19833,N_17063);
nor U26807 (N_26807,N_18868,N_16243);
and U26808 (N_26808,N_14751,N_12141);
and U26809 (N_26809,N_14921,N_12563);
nand U26810 (N_26810,N_19451,N_15781);
nor U26811 (N_26811,N_18849,N_10517);
nand U26812 (N_26812,N_12186,N_19134);
nand U26813 (N_26813,N_15586,N_18314);
xor U26814 (N_26814,N_16733,N_14275);
and U26815 (N_26815,N_18537,N_13407);
nor U26816 (N_26816,N_18736,N_11737);
or U26817 (N_26817,N_12486,N_18065);
nor U26818 (N_26818,N_10781,N_16514);
nand U26819 (N_26819,N_14130,N_18546);
xor U26820 (N_26820,N_15884,N_14904);
nor U26821 (N_26821,N_16645,N_11666);
or U26822 (N_26822,N_17082,N_15183);
nand U26823 (N_26823,N_15423,N_19815);
nor U26824 (N_26824,N_12495,N_10725);
xor U26825 (N_26825,N_11255,N_17051);
nor U26826 (N_26826,N_12218,N_16687);
or U26827 (N_26827,N_16071,N_12279);
and U26828 (N_26828,N_13903,N_12731);
or U26829 (N_26829,N_18230,N_15729);
and U26830 (N_26830,N_18636,N_18154);
or U26831 (N_26831,N_11000,N_13927);
xor U26832 (N_26832,N_14781,N_13099);
or U26833 (N_26833,N_14584,N_12711);
nand U26834 (N_26834,N_19937,N_17292);
xor U26835 (N_26835,N_15273,N_19244);
and U26836 (N_26836,N_17283,N_16586);
or U26837 (N_26837,N_13187,N_17647);
and U26838 (N_26838,N_19116,N_12690);
nand U26839 (N_26839,N_18745,N_10519);
or U26840 (N_26840,N_17828,N_12049);
nand U26841 (N_26841,N_13632,N_12711);
and U26842 (N_26842,N_15205,N_19521);
nor U26843 (N_26843,N_15314,N_17763);
or U26844 (N_26844,N_18742,N_13012);
and U26845 (N_26845,N_18815,N_16734);
xnor U26846 (N_26846,N_10462,N_17842);
and U26847 (N_26847,N_14339,N_17564);
nand U26848 (N_26848,N_19191,N_19679);
nand U26849 (N_26849,N_17900,N_13059);
and U26850 (N_26850,N_14099,N_11962);
nor U26851 (N_26851,N_17001,N_15530);
nand U26852 (N_26852,N_13417,N_17266);
or U26853 (N_26853,N_12390,N_15149);
or U26854 (N_26854,N_18926,N_14577);
or U26855 (N_26855,N_11750,N_11567);
nor U26856 (N_26856,N_18545,N_17007);
or U26857 (N_26857,N_17914,N_15674);
and U26858 (N_26858,N_18711,N_14008);
or U26859 (N_26859,N_10663,N_10392);
and U26860 (N_26860,N_19888,N_10981);
nand U26861 (N_26861,N_10098,N_19402);
or U26862 (N_26862,N_12636,N_15606);
and U26863 (N_26863,N_14895,N_13098);
nand U26864 (N_26864,N_15678,N_13487);
nand U26865 (N_26865,N_10584,N_14166);
xor U26866 (N_26866,N_15312,N_13266);
and U26867 (N_26867,N_13059,N_17116);
nor U26868 (N_26868,N_18413,N_17475);
or U26869 (N_26869,N_15973,N_15367);
and U26870 (N_26870,N_18366,N_13411);
xor U26871 (N_26871,N_19633,N_19594);
xnor U26872 (N_26872,N_11535,N_11855);
and U26873 (N_26873,N_18481,N_19814);
and U26874 (N_26874,N_13700,N_11657);
or U26875 (N_26875,N_14855,N_16151);
nor U26876 (N_26876,N_10248,N_14997);
or U26877 (N_26877,N_16978,N_19461);
and U26878 (N_26878,N_17164,N_11640);
nor U26879 (N_26879,N_15790,N_11734);
and U26880 (N_26880,N_15005,N_13433);
nor U26881 (N_26881,N_15967,N_12248);
and U26882 (N_26882,N_19998,N_14633);
nand U26883 (N_26883,N_19403,N_18826);
nand U26884 (N_26884,N_19169,N_12491);
nand U26885 (N_26885,N_12548,N_14672);
or U26886 (N_26886,N_19935,N_11006);
nor U26887 (N_26887,N_12248,N_13418);
or U26888 (N_26888,N_12812,N_14302);
and U26889 (N_26889,N_18146,N_18532);
xnor U26890 (N_26890,N_17263,N_16257);
and U26891 (N_26891,N_16599,N_19451);
and U26892 (N_26892,N_19061,N_17850);
nand U26893 (N_26893,N_11513,N_11051);
xor U26894 (N_26894,N_12891,N_16941);
nor U26895 (N_26895,N_17528,N_16490);
xor U26896 (N_26896,N_16267,N_16419);
xor U26897 (N_26897,N_12184,N_16522);
or U26898 (N_26898,N_18629,N_19074);
xor U26899 (N_26899,N_18401,N_12498);
nor U26900 (N_26900,N_18131,N_15192);
or U26901 (N_26901,N_13227,N_19438);
and U26902 (N_26902,N_14646,N_10112);
nand U26903 (N_26903,N_11685,N_10306);
and U26904 (N_26904,N_14656,N_18771);
nand U26905 (N_26905,N_14967,N_14078);
and U26906 (N_26906,N_15048,N_15768);
xnor U26907 (N_26907,N_12298,N_13601);
and U26908 (N_26908,N_17614,N_12737);
nor U26909 (N_26909,N_17156,N_16664);
xor U26910 (N_26910,N_16201,N_14429);
xnor U26911 (N_26911,N_14932,N_18098);
nor U26912 (N_26912,N_10104,N_17944);
or U26913 (N_26913,N_12358,N_14743);
or U26914 (N_26914,N_13875,N_12965);
and U26915 (N_26915,N_10422,N_18269);
and U26916 (N_26916,N_17078,N_18287);
and U26917 (N_26917,N_11162,N_15699);
nand U26918 (N_26918,N_17169,N_17329);
nand U26919 (N_26919,N_11914,N_17669);
xnor U26920 (N_26920,N_16469,N_14453);
xnor U26921 (N_26921,N_18852,N_18025);
or U26922 (N_26922,N_15591,N_19781);
xnor U26923 (N_26923,N_13033,N_10703);
xnor U26924 (N_26924,N_19933,N_19111);
or U26925 (N_26925,N_15555,N_18520);
xor U26926 (N_26926,N_19171,N_19931);
nor U26927 (N_26927,N_15601,N_14687);
xor U26928 (N_26928,N_13118,N_17402);
nor U26929 (N_26929,N_19617,N_15467);
nor U26930 (N_26930,N_11241,N_13894);
nor U26931 (N_26931,N_15029,N_12802);
or U26932 (N_26932,N_15843,N_15276);
nand U26933 (N_26933,N_11546,N_14006);
xor U26934 (N_26934,N_17511,N_10587);
nor U26935 (N_26935,N_11152,N_15843);
and U26936 (N_26936,N_13221,N_11005);
xor U26937 (N_26937,N_10028,N_11231);
and U26938 (N_26938,N_13927,N_11466);
nand U26939 (N_26939,N_16717,N_13499);
nand U26940 (N_26940,N_13170,N_10170);
xnor U26941 (N_26941,N_15731,N_11738);
xnor U26942 (N_26942,N_19877,N_17241);
nor U26943 (N_26943,N_17312,N_12822);
and U26944 (N_26944,N_15531,N_15032);
xor U26945 (N_26945,N_18752,N_19609);
and U26946 (N_26946,N_19132,N_18498);
xor U26947 (N_26947,N_12642,N_19799);
and U26948 (N_26948,N_11387,N_10960);
xor U26949 (N_26949,N_12353,N_10163);
nand U26950 (N_26950,N_12786,N_18505);
or U26951 (N_26951,N_13615,N_16292);
nor U26952 (N_26952,N_11353,N_11973);
nand U26953 (N_26953,N_15063,N_13851);
and U26954 (N_26954,N_12802,N_17739);
nor U26955 (N_26955,N_14390,N_16238);
nand U26956 (N_26956,N_17247,N_16483);
and U26957 (N_26957,N_19716,N_14219);
nand U26958 (N_26958,N_14743,N_13973);
nand U26959 (N_26959,N_13143,N_16142);
or U26960 (N_26960,N_15953,N_16432);
and U26961 (N_26961,N_18752,N_15429);
and U26962 (N_26962,N_18190,N_14335);
or U26963 (N_26963,N_10960,N_14150);
nand U26964 (N_26964,N_10157,N_15777);
or U26965 (N_26965,N_13500,N_18610);
nand U26966 (N_26966,N_18228,N_13453);
and U26967 (N_26967,N_18927,N_11615);
and U26968 (N_26968,N_16889,N_19938);
nor U26969 (N_26969,N_10030,N_12341);
xor U26970 (N_26970,N_18280,N_12557);
nand U26971 (N_26971,N_15225,N_10265);
and U26972 (N_26972,N_19740,N_19817);
and U26973 (N_26973,N_13070,N_16015);
nand U26974 (N_26974,N_16364,N_19923);
or U26975 (N_26975,N_12566,N_15323);
xor U26976 (N_26976,N_14032,N_18172);
nor U26977 (N_26977,N_16235,N_13122);
xnor U26978 (N_26978,N_18096,N_13561);
nand U26979 (N_26979,N_13018,N_14715);
and U26980 (N_26980,N_10697,N_15621);
and U26981 (N_26981,N_17594,N_18564);
or U26982 (N_26982,N_16121,N_11321);
nand U26983 (N_26983,N_14255,N_18911);
nand U26984 (N_26984,N_18353,N_12550);
nand U26985 (N_26985,N_10339,N_15305);
nor U26986 (N_26986,N_14151,N_17121);
and U26987 (N_26987,N_18472,N_13444);
nor U26988 (N_26988,N_10118,N_18599);
nand U26989 (N_26989,N_11902,N_14427);
nor U26990 (N_26990,N_15855,N_17314);
xnor U26991 (N_26991,N_16689,N_11709);
nand U26992 (N_26992,N_18656,N_18359);
and U26993 (N_26993,N_14458,N_17304);
nor U26994 (N_26994,N_10128,N_19915);
or U26995 (N_26995,N_17709,N_12893);
nand U26996 (N_26996,N_15078,N_18107);
nor U26997 (N_26997,N_16668,N_10799);
nand U26998 (N_26998,N_10363,N_16211);
or U26999 (N_26999,N_13604,N_15146);
xnor U27000 (N_27000,N_19915,N_17669);
nor U27001 (N_27001,N_19703,N_10578);
or U27002 (N_27002,N_16575,N_12350);
nand U27003 (N_27003,N_13221,N_12748);
or U27004 (N_27004,N_13104,N_15729);
nand U27005 (N_27005,N_16010,N_19648);
and U27006 (N_27006,N_11908,N_19949);
xnor U27007 (N_27007,N_14227,N_16943);
xor U27008 (N_27008,N_13313,N_14324);
and U27009 (N_27009,N_15981,N_19959);
xor U27010 (N_27010,N_19194,N_12664);
xor U27011 (N_27011,N_13218,N_16057);
xor U27012 (N_27012,N_15070,N_14848);
nand U27013 (N_27013,N_14417,N_13433);
xor U27014 (N_27014,N_13198,N_15329);
xnor U27015 (N_27015,N_10702,N_18877);
nand U27016 (N_27016,N_14671,N_14208);
nand U27017 (N_27017,N_18163,N_12481);
nor U27018 (N_27018,N_19401,N_11666);
and U27019 (N_27019,N_13682,N_19257);
nor U27020 (N_27020,N_14627,N_13403);
xnor U27021 (N_27021,N_10118,N_11069);
or U27022 (N_27022,N_10325,N_19002);
and U27023 (N_27023,N_11681,N_15282);
xnor U27024 (N_27024,N_19930,N_15984);
xor U27025 (N_27025,N_16692,N_17776);
and U27026 (N_27026,N_14789,N_12621);
and U27027 (N_27027,N_10646,N_19963);
or U27028 (N_27028,N_10224,N_16966);
nor U27029 (N_27029,N_16867,N_12116);
nor U27030 (N_27030,N_11867,N_14331);
nand U27031 (N_27031,N_15495,N_12255);
or U27032 (N_27032,N_11247,N_12156);
xnor U27033 (N_27033,N_10607,N_10289);
nor U27034 (N_27034,N_13420,N_14304);
nor U27035 (N_27035,N_13905,N_16120);
or U27036 (N_27036,N_14514,N_16314);
xnor U27037 (N_27037,N_17858,N_16155);
or U27038 (N_27038,N_14121,N_12838);
and U27039 (N_27039,N_13360,N_13003);
and U27040 (N_27040,N_18265,N_13417);
nor U27041 (N_27041,N_15486,N_17140);
or U27042 (N_27042,N_10906,N_10201);
and U27043 (N_27043,N_13837,N_14208);
nand U27044 (N_27044,N_13283,N_18030);
nand U27045 (N_27045,N_17899,N_13746);
nor U27046 (N_27046,N_13811,N_13742);
or U27047 (N_27047,N_18156,N_18795);
or U27048 (N_27048,N_15887,N_17593);
and U27049 (N_27049,N_16568,N_18465);
and U27050 (N_27050,N_14508,N_19509);
and U27051 (N_27051,N_11634,N_14379);
nor U27052 (N_27052,N_13442,N_15726);
nor U27053 (N_27053,N_12941,N_10877);
nand U27054 (N_27054,N_10096,N_15187);
nor U27055 (N_27055,N_19269,N_12015);
nor U27056 (N_27056,N_15353,N_16866);
nand U27057 (N_27057,N_13254,N_16472);
xnor U27058 (N_27058,N_11177,N_15188);
nand U27059 (N_27059,N_15365,N_16628);
nor U27060 (N_27060,N_11262,N_13951);
and U27061 (N_27061,N_10375,N_18354);
and U27062 (N_27062,N_10642,N_11129);
and U27063 (N_27063,N_13699,N_16374);
nor U27064 (N_27064,N_13786,N_13778);
or U27065 (N_27065,N_10587,N_15042);
nand U27066 (N_27066,N_18148,N_10726);
nor U27067 (N_27067,N_18133,N_13862);
or U27068 (N_27068,N_10735,N_11945);
or U27069 (N_27069,N_16529,N_12978);
and U27070 (N_27070,N_19141,N_16061);
and U27071 (N_27071,N_15594,N_11175);
xnor U27072 (N_27072,N_16685,N_17674);
nand U27073 (N_27073,N_16804,N_16602);
and U27074 (N_27074,N_12412,N_16038);
and U27075 (N_27075,N_18646,N_10206);
or U27076 (N_27076,N_11469,N_13830);
or U27077 (N_27077,N_19469,N_12164);
xor U27078 (N_27078,N_12873,N_10150);
xnor U27079 (N_27079,N_14272,N_10526);
or U27080 (N_27080,N_19583,N_11049);
nand U27081 (N_27081,N_15983,N_15532);
nor U27082 (N_27082,N_13350,N_12529);
nor U27083 (N_27083,N_12128,N_15076);
nor U27084 (N_27084,N_14260,N_15613);
nor U27085 (N_27085,N_10051,N_12405);
nand U27086 (N_27086,N_17404,N_13933);
or U27087 (N_27087,N_16073,N_15802);
and U27088 (N_27088,N_14235,N_10251);
nor U27089 (N_27089,N_10500,N_17928);
and U27090 (N_27090,N_16347,N_11401);
xnor U27091 (N_27091,N_11570,N_11239);
nor U27092 (N_27092,N_17860,N_11722);
nand U27093 (N_27093,N_13817,N_15874);
nand U27094 (N_27094,N_10770,N_10356);
and U27095 (N_27095,N_18437,N_11507);
nand U27096 (N_27096,N_12227,N_17389);
and U27097 (N_27097,N_12005,N_16047);
xnor U27098 (N_27098,N_13331,N_15338);
nand U27099 (N_27099,N_15363,N_17556);
nand U27100 (N_27100,N_19321,N_17494);
or U27101 (N_27101,N_17653,N_15224);
xor U27102 (N_27102,N_13308,N_18407);
nor U27103 (N_27103,N_15284,N_14498);
or U27104 (N_27104,N_10432,N_13896);
nand U27105 (N_27105,N_13768,N_11738);
nor U27106 (N_27106,N_13069,N_18008);
xor U27107 (N_27107,N_14434,N_12067);
nand U27108 (N_27108,N_13821,N_12365);
and U27109 (N_27109,N_10310,N_17760);
nand U27110 (N_27110,N_10049,N_13461);
xnor U27111 (N_27111,N_15756,N_19240);
and U27112 (N_27112,N_12435,N_18244);
nor U27113 (N_27113,N_18615,N_11672);
xnor U27114 (N_27114,N_18967,N_17578);
or U27115 (N_27115,N_11474,N_13826);
xor U27116 (N_27116,N_14744,N_13390);
or U27117 (N_27117,N_17481,N_19897);
nor U27118 (N_27118,N_19971,N_12522);
xor U27119 (N_27119,N_11472,N_12216);
xor U27120 (N_27120,N_17392,N_10485);
nor U27121 (N_27121,N_18123,N_12279);
or U27122 (N_27122,N_15417,N_13525);
nor U27123 (N_27123,N_17430,N_18709);
nor U27124 (N_27124,N_15724,N_17430);
and U27125 (N_27125,N_14401,N_16464);
nor U27126 (N_27126,N_17045,N_15092);
xnor U27127 (N_27127,N_12463,N_10448);
and U27128 (N_27128,N_17820,N_13059);
nor U27129 (N_27129,N_12473,N_14457);
xor U27130 (N_27130,N_10004,N_12406);
and U27131 (N_27131,N_10208,N_12140);
xor U27132 (N_27132,N_11624,N_13598);
and U27133 (N_27133,N_10301,N_17121);
or U27134 (N_27134,N_16222,N_18627);
nand U27135 (N_27135,N_11487,N_18890);
nand U27136 (N_27136,N_11371,N_14522);
and U27137 (N_27137,N_17840,N_14814);
nor U27138 (N_27138,N_18063,N_13258);
nand U27139 (N_27139,N_18936,N_11660);
nand U27140 (N_27140,N_18391,N_14227);
xor U27141 (N_27141,N_18616,N_11398);
nand U27142 (N_27142,N_17087,N_14225);
nand U27143 (N_27143,N_14973,N_18361);
xnor U27144 (N_27144,N_19146,N_17552);
xnor U27145 (N_27145,N_13169,N_13683);
nand U27146 (N_27146,N_10742,N_10406);
xnor U27147 (N_27147,N_19106,N_16728);
nor U27148 (N_27148,N_12873,N_11650);
nand U27149 (N_27149,N_18194,N_11594);
nor U27150 (N_27150,N_13892,N_15700);
or U27151 (N_27151,N_15976,N_19430);
or U27152 (N_27152,N_15075,N_14380);
nand U27153 (N_27153,N_10638,N_15090);
nor U27154 (N_27154,N_19100,N_19206);
xor U27155 (N_27155,N_13509,N_10363);
nor U27156 (N_27156,N_14213,N_16186);
or U27157 (N_27157,N_17480,N_14085);
nand U27158 (N_27158,N_10127,N_11341);
nand U27159 (N_27159,N_11883,N_18519);
or U27160 (N_27160,N_13554,N_16864);
and U27161 (N_27161,N_19409,N_18690);
xor U27162 (N_27162,N_10471,N_14444);
and U27163 (N_27163,N_13868,N_11214);
nand U27164 (N_27164,N_14930,N_19957);
nand U27165 (N_27165,N_13697,N_17180);
and U27166 (N_27166,N_17190,N_10870);
nor U27167 (N_27167,N_16092,N_11709);
xnor U27168 (N_27168,N_17462,N_11631);
nor U27169 (N_27169,N_19628,N_19461);
nand U27170 (N_27170,N_10345,N_10005);
nor U27171 (N_27171,N_17074,N_19267);
nand U27172 (N_27172,N_10096,N_17071);
and U27173 (N_27173,N_19519,N_10830);
xor U27174 (N_27174,N_13898,N_13934);
or U27175 (N_27175,N_14347,N_13274);
nor U27176 (N_27176,N_18792,N_17885);
xnor U27177 (N_27177,N_17608,N_10075);
xor U27178 (N_27178,N_16332,N_13779);
nand U27179 (N_27179,N_13344,N_11168);
xnor U27180 (N_27180,N_18440,N_15363);
xnor U27181 (N_27181,N_12937,N_13314);
nor U27182 (N_27182,N_18207,N_11448);
and U27183 (N_27183,N_15757,N_11062);
xor U27184 (N_27184,N_11028,N_11983);
and U27185 (N_27185,N_11066,N_11642);
nand U27186 (N_27186,N_18966,N_15784);
and U27187 (N_27187,N_12423,N_17728);
xnor U27188 (N_27188,N_15817,N_16759);
and U27189 (N_27189,N_13358,N_11359);
xnor U27190 (N_27190,N_15647,N_17948);
and U27191 (N_27191,N_19961,N_12032);
xor U27192 (N_27192,N_18817,N_14074);
xnor U27193 (N_27193,N_11613,N_19527);
and U27194 (N_27194,N_18268,N_19391);
or U27195 (N_27195,N_18612,N_14613);
or U27196 (N_27196,N_16755,N_19622);
or U27197 (N_27197,N_15984,N_12709);
nor U27198 (N_27198,N_12149,N_14785);
xnor U27199 (N_27199,N_15665,N_15308);
nor U27200 (N_27200,N_13510,N_19606);
xor U27201 (N_27201,N_17460,N_11251);
xor U27202 (N_27202,N_19987,N_17982);
or U27203 (N_27203,N_15479,N_14636);
nand U27204 (N_27204,N_16639,N_10178);
xnor U27205 (N_27205,N_17501,N_19556);
or U27206 (N_27206,N_12035,N_14782);
or U27207 (N_27207,N_11267,N_17741);
nand U27208 (N_27208,N_18063,N_18039);
xnor U27209 (N_27209,N_19774,N_19487);
and U27210 (N_27210,N_17085,N_18531);
and U27211 (N_27211,N_14583,N_10689);
xor U27212 (N_27212,N_14548,N_13247);
nor U27213 (N_27213,N_10840,N_19603);
xor U27214 (N_27214,N_17943,N_10358);
nor U27215 (N_27215,N_10056,N_15118);
nand U27216 (N_27216,N_12414,N_17295);
or U27217 (N_27217,N_13871,N_14605);
xor U27218 (N_27218,N_15657,N_16000);
and U27219 (N_27219,N_10794,N_13723);
xnor U27220 (N_27220,N_18034,N_15494);
nand U27221 (N_27221,N_13886,N_15983);
nor U27222 (N_27222,N_16698,N_13829);
nand U27223 (N_27223,N_11254,N_12416);
nor U27224 (N_27224,N_18471,N_15830);
and U27225 (N_27225,N_12059,N_16511);
and U27226 (N_27226,N_17757,N_12199);
or U27227 (N_27227,N_17133,N_11505);
or U27228 (N_27228,N_18090,N_16680);
nand U27229 (N_27229,N_15732,N_19147);
nor U27230 (N_27230,N_15514,N_16672);
nor U27231 (N_27231,N_15144,N_12672);
nand U27232 (N_27232,N_12802,N_19957);
or U27233 (N_27233,N_18544,N_10376);
and U27234 (N_27234,N_16791,N_15457);
or U27235 (N_27235,N_17191,N_12326);
nor U27236 (N_27236,N_14813,N_15984);
xor U27237 (N_27237,N_13718,N_19780);
or U27238 (N_27238,N_19953,N_17579);
nand U27239 (N_27239,N_11053,N_13649);
and U27240 (N_27240,N_10239,N_14166);
nand U27241 (N_27241,N_12429,N_18789);
nor U27242 (N_27242,N_12251,N_15737);
or U27243 (N_27243,N_12141,N_19987);
and U27244 (N_27244,N_15026,N_12740);
or U27245 (N_27245,N_16375,N_14537);
or U27246 (N_27246,N_10919,N_16745);
xnor U27247 (N_27247,N_14226,N_15334);
or U27248 (N_27248,N_18601,N_19538);
nor U27249 (N_27249,N_10209,N_16362);
nand U27250 (N_27250,N_12078,N_15329);
xor U27251 (N_27251,N_12512,N_16656);
or U27252 (N_27252,N_18864,N_10545);
xor U27253 (N_27253,N_11746,N_14808);
or U27254 (N_27254,N_13722,N_17316);
or U27255 (N_27255,N_16070,N_13241);
nand U27256 (N_27256,N_17214,N_10430);
nor U27257 (N_27257,N_11991,N_13879);
and U27258 (N_27258,N_19063,N_19562);
and U27259 (N_27259,N_17209,N_19771);
nor U27260 (N_27260,N_17668,N_19679);
or U27261 (N_27261,N_11127,N_10524);
or U27262 (N_27262,N_12858,N_16446);
nor U27263 (N_27263,N_17189,N_16306);
and U27264 (N_27264,N_11610,N_17183);
nand U27265 (N_27265,N_12767,N_15748);
nor U27266 (N_27266,N_14473,N_15600);
or U27267 (N_27267,N_10789,N_12447);
xor U27268 (N_27268,N_17094,N_18242);
or U27269 (N_27269,N_16781,N_10042);
and U27270 (N_27270,N_18727,N_16946);
and U27271 (N_27271,N_11137,N_14803);
and U27272 (N_27272,N_15733,N_10752);
nor U27273 (N_27273,N_19363,N_19713);
xnor U27274 (N_27274,N_13522,N_15423);
nor U27275 (N_27275,N_10155,N_18019);
nand U27276 (N_27276,N_19924,N_18341);
nand U27277 (N_27277,N_11442,N_12584);
nor U27278 (N_27278,N_10383,N_14941);
nand U27279 (N_27279,N_12009,N_15470);
nor U27280 (N_27280,N_13644,N_14335);
or U27281 (N_27281,N_10753,N_19155);
or U27282 (N_27282,N_11582,N_12837);
nand U27283 (N_27283,N_10705,N_19245);
and U27284 (N_27284,N_16474,N_11361);
or U27285 (N_27285,N_14684,N_15632);
xor U27286 (N_27286,N_16326,N_12006);
nor U27287 (N_27287,N_19091,N_18024);
and U27288 (N_27288,N_19117,N_18589);
xnor U27289 (N_27289,N_16912,N_17762);
xnor U27290 (N_27290,N_12209,N_10349);
nor U27291 (N_27291,N_10502,N_12429);
xor U27292 (N_27292,N_19815,N_11944);
or U27293 (N_27293,N_19766,N_10113);
nand U27294 (N_27294,N_19472,N_15647);
xnor U27295 (N_27295,N_16525,N_17752);
and U27296 (N_27296,N_13638,N_15078);
xor U27297 (N_27297,N_14765,N_16400);
nand U27298 (N_27298,N_12123,N_10312);
and U27299 (N_27299,N_14141,N_12129);
and U27300 (N_27300,N_11217,N_18955);
nor U27301 (N_27301,N_15522,N_19209);
or U27302 (N_27302,N_16520,N_19301);
and U27303 (N_27303,N_12417,N_10327);
and U27304 (N_27304,N_15970,N_16554);
or U27305 (N_27305,N_12810,N_10383);
nor U27306 (N_27306,N_19895,N_11769);
nor U27307 (N_27307,N_13529,N_19794);
nand U27308 (N_27308,N_18637,N_19903);
nand U27309 (N_27309,N_10543,N_17084);
nor U27310 (N_27310,N_16666,N_16421);
xnor U27311 (N_27311,N_11521,N_12172);
or U27312 (N_27312,N_15116,N_15662);
or U27313 (N_27313,N_18209,N_14987);
and U27314 (N_27314,N_17043,N_13125);
nand U27315 (N_27315,N_18060,N_11405);
nand U27316 (N_27316,N_19255,N_10367);
and U27317 (N_27317,N_12681,N_12704);
and U27318 (N_27318,N_18734,N_16710);
nor U27319 (N_27319,N_15691,N_11560);
nand U27320 (N_27320,N_11713,N_17306);
nor U27321 (N_27321,N_13595,N_13786);
and U27322 (N_27322,N_19585,N_15074);
or U27323 (N_27323,N_16887,N_18291);
nor U27324 (N_27324,N_11223,N_13523);
or U27325 (N_27325,N_11239,N_11307);
nor U27326 (N_27326,N_16859,N_12216);
and U27327 (N_27327,N_13108,N_14228);
or U27328 (N_27328,N_17052,N_14298);
or U27329 (N_27329,N_11258,N_19836);
nand U27330 (N_27330,N_18371,N_14689);
xor U27331 (N_27331,N_12905,N_12593);
nand U27332 (N_27332,N_13405,N_19574);
or U27333 (N_27333,N_14508,N_13467);
or U27334 (N_27334,N_14587,N_17578);
and U27335 (N_27335,N_12960,N_12467);
xor U27336 (N_27336,N_18770,N_11211);
nor U27337 (N_27337,N_12302,N_16526);
and U27338 (N_27338,N_16958,N_11197);
nand U27339 (N_27339,N_14429,N_12092);
xnor U27340 (N_27340,N_10974,N_15745);
and U27341 (N_27341,N_14171,N_13371);
and U27342 (N_27342,N_12726,N_14489);
or U27343 (N_27343,N_17455,N_18363);
and U27344 (N_27344,N_11450,N_16192);
or U27345 (N_27345,N_18476,N_11034);
or U27346 (N_27346,N_10918,N_11022);
nor U27347 (N_27347,N_16740,N_12679);
or U27348 (N_27348,N_15519,N_14768);
xnor U27349 (N_27349,N_10003,N_15862);
or U27350 (N_27350,N_18227,N_18060);
and U27351 (N_27351,N_18347,N_10643);
nand U27352 (N_27352,N_11243,N_19198);
nor U27353 (N_27353,N_12096,N_11760);
xor U27354 (N_27354,N_17645,N_16006);
and U27355 (N_27355,N_15426,N_16070);
and U27356 (N_27356,N_12555,N_10597);
xnor U27357 (N_27357,N_18910,N_15912);
nor U27358 (N_27358,N_15186,N_17960);
or U27359 (N_27359,N_12607,N_11848);
and U27360 (N_27360,N_14810,N_10700);
nand U27361 (N_27361,N_15406,N_14903);
nand U27362 (N_27362,N_18661,N_14257);
xor U27363 (N_27363,N_18972,N_15823);
nand U27364 (N_27364,N_18482,N_14681);
nand U27365 (N_27365,N_14879,N_17569);
or U27366 (N_27366,N_15051,N_19937);
nand U27367 (N_27367,N_19357,N_18285);
xnor U27368 (N_27368,N_16304,N_17089);
nand U27369 (N_27369,N_19841,N_18308);
xnor U27370 (N_27370,N_19136,N_12814);
nand U27371 (N_27371,N_11434,N_15975);
nand U27372 (N_27372,N_14362,N_12646);
nand U27373 (N_27373,N_12495,N_16719);
or U27374 (N_27374,N_16604,N_13577);
or U27375 (N_27375,N_19353,N_11377);
xnor U27376 (N_27376,N_12517,N_16457);
or U27377 (N_27377,N_17203,N_12622);
and U27378 (N_27378,N_19926,N_12034);
or U27379 (N_27379,N_13318,N_15492);
and U27380 (N_27380,N_15967,N_10817);
and U27381 (N_27381,N_10371,N_13012);
nor U27382 (N_27382,N_11411,N_12324);
or U27383 (N_27383,N_14923,N_13204);
nor U27384 (N_27384,N_18649,N_16788);
or U27385 (N_27385,N_18063,N_14617);
xor U27386 (N_27386,N_11525,N_16284);
or U27387 (N_27387,N_11041,N_14828);
or U27388 (N_27388,N_12699,N_17869);
xnor U27389 (N_27389,N_17464,N_12913);
and U27390 (N_27390,N_18947,N_11128);
nor U27391 (N_27391,N_15417,N_13466);
and U27392 (N_27392,N_16481,N_16067);
xnor U27393 (N_27393,N_10392,N_17451);
and U27394 (N_27394,N_19591,N_11976);
or U27395 (N_27395,N_13938,N_19846);
xnor U27396 (N_27396,N_15174,N_14200);
xnor U27397 (N_27397,N_10560,N_18354);
nand U27398 (N_27398,N_16353,N_17824);
xor U27399 (N_27399,N_16284,N_10026);
nor U27400 (N_27400,N_12349,N_19984);
and U27401 (N_27401,N_13850,N_14044);
xnor U27402 (N_27402,N_12199,N_17803);
and U27403 (N_27403,N_19016,N_16518);
xor U27404 (N_27404,N_11531,N_10361);
nand U27405 (N_27405,N_11564,N_17203);
or U27406 (N_27406,N_11983,N_13928);
or U27407 (N_27407,N_19224,N_19388);
and U27408 (N_27408,N_18587,N_16826);
nor U27409 (N_27409,N_10184,N_12557);
xor U27410 (N_27410,N_19144,N_12158);
nor U27411 (N_27411,N_15739,N_13591);
xnor U27412 (N_27412,N_13099,N_14790);
or U27413 (N_27413,N_12163,N_18188);
or U27414 (N_27414,N_16998,N_17121);
or U27415 (N_27415,N_10864,N_15132);
or U27416 (N_27416,N_15336,N_18640);
nor U27417 (N_27417,N_13891,N_12269);
and U27418 (N_27418,N_11972,N_11534);
nand U27419 (N_27419,N_17429,N_11252);
nor U27420 (N_27420,N_12312,N_12003);
or U27421 (N_27421,N_18892,N_18495);
xnor U27422 (N_27422,N_12994,N_15813);
xor U27423 (N_27423,N_17201,N_14143);
and U27424 (N_27424,N_13301,N_11468);
or U27425 (N_27425,N_13748,N_14567);
xnor U27426 (N_27426,N_18358,N_19545);
and U27427 (N_27427,N_18724,N_12885);
nand U27428 (N_27428,N_16489,N_12562);
and U27429 (N_27429,N_13346,N_12251);
nor U27430 (N_27430,N_14723,N_12527);
nand U27431 (N_27431,N_12235,N_13972);
xnor U27432 (N_27432,N_17228,N_13206);
xnor U27433 (N_27433,N_14106,N_11859);
and U27434 (N_27434,N_10372,N_12028);
nand U27435 (N_27435,N_11203,N_16189);
or U27436 (N_27436,N_12404,N_13597);
nand U27437 (N_27437,N_13427,N_10446);
xnor U27438 (N_27438,N_19841,N_15844);
xor U27439 (N_27439,N_16667,N_18937);
and U27440 (N_27440,N_13922,N_10241);
and U27441 (N_27441,N_10162,N_10241);
xor U27442 (N_27442,N_19350,N_15702);
xnor U27443 (N_27443,N_18581,N_13925);
or U27444 (N_27444,N_12748,N_13521);
xnor U27445 (N_27445,N_13144,N_16447);
and U27446 (N_27446,N_11493,N_17552);
nand U27447 (N_27447,N_18705,N_15306);
or U27448 (N_27448,N_18191,N_18197);
or U27449 (N_27449,N_13642,N_16353);
or U27450 (N_27450,N_12747,N_12814);
and U27451 (N_27451,N_19443,N_13060);
xor U27452 (N_27452,N_10025,N_12111);
nand U27453 (N_27453,N_14369,N_15266);
and U27454 (N_27454,N_17794,N_16834);
or U27455 (N_27455,N_11784,N_13939);
nand U27456 (N_27456,N_16592,N_13109);
xor U27457 (N_27457,N_13156,N_13111);
and U27458 (N_27458,N_17744,N_13787);
or U27459 (N_27459,N_14676,N_11844);
and U27460 (N_27460,N_15293,N_19903);
xor U27461 (N_27461,N_14130,N_18980);
xor U27462 (N_27462,N_12411,N_15505);
nand U27463 (N_27463,N_14434,N_18215);
xnor U27464 (N_27464,N_19609,N_17970);
nor U27465 (N_27465,N_14814,N_16267);
nand U27466 (N_27466,N_18711,N_14040);
or U27467 (N_27467,N_12081,N_17396);
xor U27468 (N_27468,N_19564,N_16771);
or U27469 (N_27469,N_12972,N_12614);
nor U27470 (N_27470,N_11086,N_12294);
xor U27471 (N_27471,N_11128,N_13045);
nor U27472 (N_27472,N_16392,N_14213);
xor U27473 (N_27473,N_17769,N_18768);
xor U27474 (N_27474,N_18823,N_18941);
or U27475 (N_27475,N_13134,N_17271);
nor U27476 (N_27476,N_12739,N_17502);
and U27477 (N_27477,N_17135,N_19643);
xnor U27478 (N_27478,N_18531,N_16272);
nand U27479 (N_27479,N_11164,N_11026);
or U27480 (N_27480,N_16353,N_11701);
xnor U27481 (N_27481,N_10526,N_10364);
nor U27482 (N_27482,N_14990,N_15362);
nand U27483 (N_27483,N_16126,N_15348);
or U27484 (N_27484,N_10153,N_15345);
nand U27485 (N_27485,N_13445,N_10689);
and U27486 (N_27486,N_16040,N_18267);
and U27487 (N_27487,N_12833,N_15057);
nand U27488 (N_27488,N_13399,N_11514);
or U27489 (N_27489,N_16408,N_10094);
xnor U27490 (N_27490,N_18332,N_19087);
nand U27491 (N_27491,N_16291,N_14674);
and U27492 (N_27492,N_14981,N_15003);
and U27493 (N_27493,N_12569,N_17827);
nor U27494 (N_27494,N_12467,N_10357);
nand U27495 (N_27495,N_15534,N_15533);
and U27496 (N_27496,N_15130,N_16789);
nor U27497 (N_27497,N_16001,N_18316);
nand U27498 (N_27498,N_14017,N_12318);
and U27499 (N_27499,N_15115,N_14867);
xor U27500 (N_27500,N_15819,N_11650);
nor U27501 (N_27501,N_15634,N_19529);
and U27502 (N_27502,N_14696,N_15253);
xor U27503 (N_27503,N_19008,N_16744);
nor U27504 (N_27504,N_16814,N_15917);
nand U27505 (N_27505,N_16345,N_13446);
nor U27506 (N_27506,N_17156,N_17122);
nor U27507 (N_27507,N_13320,N_17600);
and U27508 (N_27508,N_15395,N_17531);
nand U27509 (N_27509,N_19459,N_14914);
nand U27510 (N_27510,N_18942,N_10476);
nor U27511 (N_27511,N_11032,N_13228);
or U27512 (N_27512,N_11257,N_16497);
nand U27513 (N_27513,N_10756,N_19071);
xnor U27514 (N_27514,N_16496,N_14047);
nand U27515 (N_27515,N_17796,N_11748);
nand U27516 (N_27516,N_19435,N_10081);
nand U27517 (N_27517,N_11821,N_14385);
nand U27518 (N_27518,N_16416,N_16728);
or U27519 (N_27519,N_18497,N_17236);
xor U27520 (N_27520,N_17394,N_10099);
nor U27521 (N_27521,N_16877,N_14951);
and U27522 (N_27522,N_11031,N_18601);
xor U27523 (N_27523,N_10627,N_12734);
nor U27524 (N_27524,N_18104,N_19318);
nand U27525 (N_27525,N_16168,N_16214);
or U27526 (N_27526,N_13993,N_19778);
nand U27527 (N_27527,N_15750,N_11512);
and U27528 (N_27528,N_10910,N_10155);
xor U27529 (N_27529,N_11232,N_19791);
nor U27530 (N_27530,N_11024,N_16092);
xor U27531 (N_27531,N_19705,N_18370);
and U27532 (N_27532,N_17346,N_14064);
xnor U27533 (N_27533,N_10523,N_13745);
nor U27534 (N_27534,N_17702,N_17187);
nor U27535 (N_27535,N_13778,N_12631);
or U27536 (N_27536,N_12146,N_17601);
nand U27537 (N_27537,N_19061,N_19983);
nand U27538 (N_27538,N_12943,N_10003);
nor U27539 (N_27539,N_13526,N_16714);
nand U27540 (N_27540,N_11432,N_19691);
nand U27541 (N_27541,N_16267,N_17002);
and U27542 (N_27542,N_12849,N_10690);
nor U27543 (N_27543,N_12438,N_10432);
nand U27544 (N_27544,N_15369,N_17973);
nand U27545 (N_27545,N_19737,N_15299);
nor U27546 (N_27546,N_10154,N_11144);
xor U27547 (N_27547,N_10465,N_10089);
nor U27548 (N_27548,N_15046,N_13815);
xnor U27549 (N_27549,N_12263,N_10729);
and U27550 (N_27550,N_10299,N_12979);
xnor U27551 (N_27551,N_13672,N_15354);
nand U27552 (N_27552,N_14802,N_13095);
xor U27553 (N_27553,N_19321,N_17141);
xnor U27554 (N_27554,N_19406,N_11327);
nand U27555 (N_27555,N_12320,N_16421);
nor U27556 (N_27556,N_13265,N_11203);
nand U27557 (N_27557,N_13705,N_11463);
nor U27558 (N_27558,N_15664,N_18150);
and U27559 (N_27559,N_16248,N_17857);
nor U27560 (N_27560,N_16042,N_13327);
or U27561 (N_27561,N_13159,N_11589);
nor U27562 (N_27562,N_12507,N_11989);
xnor U27563 (N_27563,N_15333,N_16235);
nand U27564 (N_27564,N_14656,N_18933);
or U27565 (N_27565,N_10145,N_11048);
nand U27566 (N_27566,N_11734,N_12342);
or U27567 (N_27567,N_13716,N_16317);
nand U27568 (N_27568,N_19630,N_14326);
and U27569 (N_27569,N_17821,N_14377);
nand U27570 (N_27570,N_16003,N_17725);
or U27571 (N_27571,N_13679,N_11030);
nand U27572 (N_27572,N_11347,N_10902);
xor U27573 (N_27573,N_15084,N_17506);
nand U27574 (N_27574,N_14581,N_19515);
or U27575 (N_27575,N_18953,N_16892);
nor U27576 (N_27576,N_18878,N_17293);
or U27577 (N_27577,N_13815,N_19522);
or U27578 (N_27578,N_14307,N_19441);
nor U27579 (N_27579,N_13747,N_13346);
nor U27580 (N_27580,N_19113,N_19195);
nand U27581 (N_27581,N_10005,N_15987);
xor U27582 (N_27582,N_13537,N_14325);
xnor U27583 (N_27583,N_19107,N_16544);
or U27584 (N_27584,N_11850,N_17104);
and U27585 (N_27585,N_19225,N_12390);
nor U27586 (N_27586,N_12124,N_12144);
and U27587 (N_27587,N_12466,N_12708);
xnor U27588 (N_27588,N_19672,N_15162);
or U27589 (N_27589,N_15643,N_10291);
xnor U27590 (N_27590,N_18975,N_10987);
xnor U27591 (N_27591,N_18990,N_12619);
and U27592 (N_27592,N_15349,N_15653);
xor U27593 (N_27593,N_19892,N_13996);
and U27594 (N_27594,N_18419,N_18070);
xor U27595 (N_27595,N_11851,N_11248);
xnor U27596 (N_27596,N_15956,N_11498);
or U27597 (N_27597,N_14593,N_12053);
nor U27598 (N_27598,N_11120,N_19927);
nor U27599 (N_27599,N_11858,N_17158);
or U27600 (N_27600,N_14197,N_15699);
nand U27601 (N_27601,N_12113,N_13467);
nand U27602 (N_27602,N_17554,N_15083);
nor U27603 (N_27603,N_11090,N_11728);
xnor U27604 (N_27604,N_11760,N_16956);
and U27605 (N_27605,N_17333,N_13791);
nand U27606 (N_27606,N_12863,N_16740);
nand U27607 (N_27607,N_12563,N_15150);
nor U27608 (N_27608,N_17655,N_13987);
xor U27609 (N_27609,N_14109,N_19369);
and U27610 (N_27610,N_17123,N_10742);
xor U27611 (N_27611,N_16642,N_16556);
and U27612 (N_27612,N_15508,N_15948);
nor U27613 (N_27613,N_13458,N_12071);
xnor U27614 (N_27614,N_10928,N_17637);
and U27615 (N_27615,N_15621,N_19705);
nand U27616 (N_27616,N_11645,N_17719);
nor U27617 (N_27617,N_13488,N_11342);
nand U27618 (N_27618,N_12367,N_14268);
xor U27619 (N_27619,N_10086,N_18905);
xnor U27620 (N_27620,N_15369,N_13803);
and U27621 (N_27621,N_15419,N_19179);
and U27622 (N_27622,N_17347,N_14471);
or U27623 (N_27623,N_18325,N_16819);
xor U27624 (N_27624,N_15749,N_18820);
and U27625 (N_27625,N_16203,N_14375);
or U27626 (N_27626,N_15368,N_19343);
nand U27627 (N_27627,N_13841,N_12295);
xor U27628 (N_27628,N_12753,N_13628);
and U27629 (N_27629,N_15198,N_19663);
nand U27630 (N_27630,N_18854,N_18478);
or U27631 (N_27631,N_13216,N_17004);
and U27632 (N_27632,N_15523,N_10839);
nand U27633 (N_27633,N_16137,N_16052);
or U27634 (N_27634,N_19162,N_13421);
and U27635 (N_27635,N_17010,N_14637);
and U27636 (N_27636,N_16628,N_11371);
nand U27637 (N_27637,N_14823,N_10483);
and U27638 (N_27638,N_11791,N_11937);
nand U27639 (N_27639,N_14403,N_12324);
and U27640 (N_27640,N_12355,N_12307);
nand U27641 (N_27641,N_12056,N_12448);
nand U27642 (N_27642,N_18099,N_16928);
nand U27643 (N_27643,N_15853,N_13190);
and U27644 (N_27644,N_19592,N_15925);
and U27645 (N_27645,N_11988,N_12325);
nor U27646 (N_27646,N_17930,N_15547);
or U27647 (N_27647,N_16425,N_18907);
nor U27648 (N_27648,N_17162,N_16590);
xnor U27649 (N_27649,N_19125,N_18510);
nand U27650 (N_27650,N_10887,N_18174);
nand U27651 (N_27651,N_11467,N_16820);
nor U27652 (N_27652,N_18132,N_15241);
xnor U27653 (N_27653,N_19012,N_17789);
xor U27654 (N_27654,N_14686,N_16682);
nor U27655 (N_27655,N_11164,N_11065);
or U27656 (N_27656,N_12841,N_12218);
nor U27657 (N_27657,N_19928,N_17120);
xor U27658 (N_27658,N_11619,N_11843);
nand U27659 (N_27659,N_18504,N_13260);
or U27660 (N_27660,N_19390,N_13497);
nor U27661 (N_27661,N_13833,N_12240);
or U27662 (N_27662,N_12864,N_12256);
xnor U27663 (N_27663,N_12119,N_11304);
xor U27664 (N_27664,N_17248,N_17636);
nor U27665 (N_27665,N_13625,N_12904);
nor U27666 (N_27666,N_12957,N_15896);
xnor U27667 (N_27667,N_14269,N_10573);
or U27668 (N_27668,N_19112,N_16524);
and U27669 (N_27669,N_12140,N_12988);
nand U27670 (N_27670,N_13048,N_15680);
and U27671 (N_27671,N_13160,N_11135);
nor U27672 (N_27672,N_15206,N_13996);
or U27673 (N_27673,N_13195,N_18218);
nor U27674 (N_27674,N_18712,N_10199);
nand U27675 (N_27675,N_10919,N_17665);
or U27676 (N_27676,N_13658,N_18640);
or U27677 (N_27677,N_13509,N_13024);
or U27678 (N_27678,N_18620,N_19149);
nand U27679 (N_27679,N_14710,N_13379);
or U27680 (N_27680,N_11738,N_16309);
nor U27681 (N_27681,N_16434,N_17761);
and U27682 (N_27682,N_11939,N_12355);
nor U27683 (N_27683,N_16554,N_14454);
nor U27684 (N_27684,N_17839,N_17208);
xnor U27685 (N_27685,N_11097,N_17910);
xor U27686 (N_27686,N_10936,N_11962);
xor U27687 (N_27687,N_18284,N_14395);
and U27688 (N_27688,N_10714,N_16088);
or U27689 (N_27689,N_18057,N_10988);
or U27690 (N_27690,N_15124,N_16140);
xnor U27691 (N_27691,N_16500,N_18047);
xnor U27692 (N_27692,N_19756,N_11619);
xor U27693 (N_27693,N_16713,N_18983);
nor U27694 (N_27694,N_12933,N_16892);
and U27695 (N_27695,N_13590,N_15795);
xnor U27696 (N_27696,N_12271,N_12766);
xnor U27697 (N_27697,N_14220,N_14525);
or U27698 (N_27698,N_19220,N_16129);
or U27699 (N_27699,N_14082,N_11309);
nor U27700 (N_27700,N_11185,N_13223);
and U27701 (N_27701,N_19682,N_16142);
and U27702 (N_27702,N_15394,N_12365);
xor U27703 (N_27703,N_11606,N_18759);
nand U27704 (N_27704,N_17015,N_14950);
nand U27705 (N_27705,N_12238,N_11124);
nand U27706 (N_27706,N_10075,N_19626);
nand U27707 (N_27707,N_13931,N_16877);
nor U27708 (N_27708,N_11635,N_10558);
xnor U27709 (N_27709,N_12289,N_19269);
nand U27710 (N_27710,N_19258,N_11155);
and U27711 (N_27711,N_10637,N_15007);
xor U27712 (N_27712,N_14196,N_17118);
nand U27713 (N_27713,N_15233,N_10882);
nor U27714 (N_27714,N_19858,N_14605);
xnor U27715 (N_27715,N_11460,N_18128);
xnor U27716 (N_27716,N_12775,N_11262);
and U27717 (N_27717,N_10588,N_11113);
xnor U27718 (N_27718,N_14211,N_12543);
and U27719 (N_27719,N_13454,N_12772);
and U27720 (N_27720,N_16313,N_17452);
or U27721 (N_27721,N_10715,N_17225);
nor U27722 (N_27722,N_18750,N_15646);
nand U27723 (N_27723,N_15782,N_16483);
xor U27724 (N_27724,N_18353,N_18454);
and U27725 (N_27725,N_14904,N_10294);
xor U27726 (N_27726,N_11353,N_13391);
xor U27727 (N_27727,N_10339,N_19086);
and U27728 (N_27728,N_10000,N_15369);
nor U27729 (N_27729,N_14873,N_10387);
or U27730 (N_27730,N_19134,N_13310);
nor U27731 (N_27731,N_16585,N_10306);
nand U27732 (N_27732,N_12826,N_14221);
xnor U27733 (N_27733,N_16345,N_16219);
nand U27734 (N_27734,N_17726,N_11113);
nand U27735 (N_27735,N_15535,N_17299);
xnor U27736 (N_27736,N_14674,N_19631);
xor U27737 (N_27737,N_11788,N_17982);
and U27738 (N_27738,N_10572,N_10615);
xor U27739 (N_27739,N_10244,N_12183);
or U27740 (N_27740,N_19481,N_18954);
nand U27741 (N_27741,N_16575,N_15590);
xnor U27742 (N_27742,N_12127,N_19199);
xnor U27743 (N_27743,N_19938,N_13913);
xnor U27744 (N_27744,N_17350,N_10622);
nand U27745 (N_27745,N_15007,N_11542);
nand U27746 (N_27746,N_15365,N_13977);
nor U27747 (N_27747,N_11323,N_14103);
nand U27748 (N_27748,N_14466,N_17009);
and U27749 (N_27749,N_15863,N_13559);
and U27750 (N_27750,N_18149,N_11311);
and U27751 (N_27751,N_11023,N_18904);
nor U27752 (N_27752,N_15146,N_16389);
nor U27753 (N_27753,N_16437,N_13131);
or U27754 (N_27754,N_18505,N_18573);
or U27755 (N_27755,N_15211,N_11964);
nand U27756 (N_27756,N_12930,N_18643);
nor U27757 (N_27757,N_15998,N_15068);
nor U27758 (N_27758,N_11386,N_13055);
or U27759 (N_27759,N_12736,N_13391);
or U27760 (N_27760,N_15086,N_17095);
nand U27761 (N_27761,N_17861,N_14180);
xor U27762 (N_27762,N_10551,N_18372);
or U27763 (N_27763,N_11630,N_10849);
or U27764 (N_27764,N_13362,N_14353);
and U27765 (N_27765,N_13069,N_16579);
nor U27766 (N_27766,N_17336,N_15118);
nand U27767 (N_27767,N_14223,N_15678);
nand U27768 (N_27768,N_11325,N_15181);
nor U27769 (N_27769,N_19524,N_12568);
and U27770 (N_27770,N_17629,N_18932);
and U27771 (N_27771,N_13943,N_11804);
nor U27772 (N_27772,N_16980,N_18702);
and U27773 (N_27773,N_17609,N_19938);
nand U27774 (N_27774,N_17630,N_17771);
nand U27775 (N_27775,N_12240,N_15267);
or U27776 (N_27776,N_11789,N_17364);
nand U27777 (N_27777,N_16153,N_19716);
xor U27778 (N_27778,N_10842,N_18804);
or U27779 (N_27779,N_18860,N_11638);
nor U27780 (N_27780,N_13257,N_17561);
nand U27781 (N_27781,N_15668,N_16695);
nor U27782 (N_27782,N_17006,N_14542);
or U27783 (N_27783,N_10610,N_18475);
and U27784 (N_27784,N_13845,N_10666);
xor U27785 (N_27785,N_19886,N_14787);
and U27786 (N_27786,N_14839,N_19663);
and U27787 (N_27787,N_10125,N_10228);
xor U27788 (N_27788,N_19560,N_15071);
or U27789 (N_27789,N_19817,N_13686);
nor U27790 (N_27790,N_14337,N_11264);
or U27791 (N_27791,N_14127,N_11961);
xor U27792 (N_27792,N_13244,N_18660);
nor U27793 (N_27793,N_15585,N_14178);
and U27794 (N_27794,N_13350,N_13598);
nor U27795 (N_27795,N_17842,N_19009);
nor U27796 (N_27796,N_10828,N_12225);
nand U27797 (N_27797,N_12013,N_18563);
nor U27798 (N_27798,N_18682,N_10074);
nor U27799 (N_27799,N_14584,N_17185);
and U27800 (N_27800,N_10354,N_18636);
and U27801 (N_27801,N_18140,N_15595);
xnor U27802 (N_27802,N_15136,N_11673);
nor U27803 (N_27803,N_14994,N_14624);
nor U27804 (N_27804,N_11718,N_18508);
and U27805 (N_27805,N_15209,N_19044);
nand U27806 (N_27806,N_12710,N_11548);
nand U27807 (N_27807,N_19152,N_12588);
nand U27808 (N_27808,N_18404,N_17678);
and U27809 (N_27809,N_13259,N_10579);
nor U27810 (N_27810,N_18537,N_19239);
and U27811 (N_27811,N_16220,N_10258);
xor U27812 (N_27812,N_19033,N_12217);
nor U27813 (N_27813,N_11749,N_13493);
nand U27814 (N_27814,N_17821,N_19014);
nand U27815 (N_27815,N_18805,N_12030);
nand U27816 (N_27816,N_15686,N_17917);
nor U27817 (N_27817,N_15112,N_19872);
nor U27818 (N_27818,N_18357,N_13593);
nor U27819 (N_27819,N_16926,N_15724);
nand U27820 (N_27820,N_11547,N_19952);
and U27821 (N_27821,N_15667,N_17629);
and U27822 (N_27822,N_10310,N_13281);
and U27823 (N_27823,N_19392,N_18709);
nor U27824 (N_27824,N_19757,N_16680);
nand U27825 (N_27825,N_13506,N_13437);
or U27826 (N_27826,N_14993,N_14263);
or U27827 (N_27827,N_16595,N_14480);
nand U27828 (N_27828,N_14755,N_10705);
and U27829 (N_27829,N_14115,N_19834);
and U27830 (N_27830,N_19102,N_17255);
or U27831 (N_27831,N_18859,N_18891);
xnor U27832 (N_27832,N_16981,N_15934);
and U27833 (N_27833,N_18451,N_17390);
nor U27834 (N_27834,N_13526,N_18891);
nor U27835 (N_27835,N_14353,N_13400);
or U27836 (N_27836,N_15588,N_12224);
or U27837 (N_27837,N_11046,N_10157);
xnor U27838 (N_27838,N_18654,N_16562);
and U27839 (N_27839,N_10485,N_19058);
xor U27840 (N_27840,N_15072,N_14054);
or U27841 (N_27841,N_13692,N_14677);
nand U27842 (N_27842,N_18405,N_16490);
or U27843 (N_27843,N_14077,N_11021);
nor U27844 (N_27844,N_14413,N_11185);
nand U27845 (N_27845,N_13998,N_10487);
or U27846 (N_27846,N_19922,N_10059);
or U27847 (N_27847,N_12440,N_11967);
or U27848 (N_27848,N_12345,N_19943);
and U27849 (N_27849,N_18731,N_10156);
nand U27850 (N_27850,N_16557,N_14013);
or U27851 (N_27851,N_13305,N_13552);
xnor U27852 (N_27852,N_15200,N_13478);
nor U27853 (N_27853,N_12212,N_16831);
nand U27854 (N_27854,N_18554,N_13107);
xnor U27855 (N_27855,N_11255,N_11459);
or U27856 (N_27856,N_15764,N_15913);
and U27857 (N_27857,N_17905,N_13205);
xor U27858 (N_27858,N_12822,N_10373);
and U27859 (N_27859,N_19943,N_12283);
nand U27860 (N_27860,N_13330,N_11936);
xor U27861 (N_27861,N_13550,N_14997);
or U27862 (N_27862,N_15741,N_19839);
xnor U27863 (N_27863,N_14937,N_11614);
xor U27864 (N_27864,N_13793,N_10793);
xor U27865 (N_27865,N_12234,N_13213);
nor U27866 (N_27866,N_10656,N_15676);
and U27867 (N_27867,N_15677,N_15821);
and U27868 (N_27868,N_13393,N_12597);
or U27869 (N_27869,N_10251,N_16054);
nand U27870 (N_27870,N_18664,N_13512);
and U27871 (N_27871,N_17897,N_10401);
nor U27872 (N_27872,N_12072,N_10131);
xor U27873 (N_27873,N_17535,N_17964);
nand U27874 (N_27874,N_14987,N_11235);
nor U27875 (N_27875,N_19432,N_18845);
nand U27876 (N_27876,N_15383,N_11697);
and U27877 (N_27877,N_16366,N_17909);
or U27878 (N_27878,N_11832,N_18141);
nor U27879 (N_27879,N_14865,N_19590);
and U27880 (N_27880,N_15361,N_10859);
or U27881 (N_27881,N_19505,N_15511);
xnor U27882 (N_27882,N_19852,N_12141);
or U27883 (N_27883,N_19424,N_19122);
xor U27884 (N_27884,N_10724,N_18435);
nand U27885 (N_27885,N_14653,N_17021);
nand U27886 (N_27886,N_13281,N_14106);
and U27887 (N_27887,N_11994,N_13848);
or U27888 (N_27888,N_10924,N_14878);
nor U27889 (N_27889,N_11920,N_11805);
or U27890 (N_27890,N_14065,N_18462);
and U27891 (N_27891,N_19174,N_15604);
and U27892 (N_27892,N_16486,N_15877);
or U27893 (N_27893,N_14656,N_12534);
or U27894 (N_27894,N_18307,N_12119);
nor U27895 (N_27895,N_14080,N_18346);
xor U27896 (N_27896,N_15717,N_19173);
and U27897 (N_27897,N_12055,N_13656);
xor U27898 (N_27898,N_13078,N_12471);
nand U27899 (N_27899,N_14509,N_15216);
or U27900 (N_27900,N_15998,N_15460);
or U27901 (N_27901,N_18644,N_13970);
and U27902 (N_27902,N_16512,N_17383);
nand U27903 (N_27903,N_14603,N_14421);
xnor U27904 (N_27904,N_15742,N_16494);
xnor U27905 (N_27905,N_10433,N_15120);
xor U27906 (N_27906,N_17788,N_12557);
and U27907 (N_27907,N_11325,N_18257);
or U27908 (N_27908,N_10365,N_19369);
nand U27909 (N_27909,N_10991,N_14491);
nor U27910 (N_27910,N_16143,N_15978);
xor U27911 (N_27911,N_11763,N_14969);
xor U27912 (N_27912,N_14988,N_15700);
and U27913 (N_27913,N_14971,N_10385);
nor U27914 (N_27914,N_14444,N_15432);
or U27915 (N_27915,N_12379,N_16673);
or U27916 (N_27916,N_14322,N_11927);
nand U27917 (N_27917,N_11862,N_12220);
and U27918 (N_27918,N_14465,N_11056);
nand U27919 (N_27919,N_10747,N_12962);
and U27920 (N_27920,N_13393,N_13960);
nand U27921 (N_27921,N_11198,N_18697);
or U27922 (N_27922,N_12673,N_13085);
nand U27923 (N_27923,N_17306,N_12765);
and U27924 (N_27924,N_13664,N_14749);
and U27925 (N_27925,N_11544,N_10050);
and U27926 (N_27926,N_14123,N_14885);
nor U27927 (N_27927,N_19350,N_12571);
or U27928 (N_27928,N_14526,N_17564);
nand U27929 (N_27929,N_17288,N_10446);
and U27930 (N_27930,N_11857,N_13032);
nor U27931 (N_27931,N_16040,N_17009);
and U27932 (N_27932,N_17639,N_11396);
or U27933 (N_27933,N_15313,N_11053);
nand U27934 (N_27934,N_19134,N_16094);
or U27935 (N_27935,N_10121,N_13992);
or U27936 (N_27936,N_18855,N_16158);
and U27937 (N_27937,N_18396,N_11952);
xor U27938 (N_27938,N_19596,N_10501);
and U27939 (N_27939,N_15812,N_17648);
nand U27940 (N_27940,N_11753,N_10812);
or U27941 (N_27941,N_11280,N_17481);
xor U27942 (N_27942,N_14957,N_17163);
nor U27943 (N_27943,N_13464,N_13503);
nand U27944 (N_27944,N_15030,N_13819);
xnor U27945 (N_27945,N_18759,N_10636);
or U27946 (N_27946,N_12085,N_12452);
nor U27947 (N_27947,N_18798,N_12779);
nand U27948 (N_27948,N_14053,N_14501);
xor U27949 (N_27949,N_14674,N_19909);
xnor U27950 (N_27950,N_10668,N_18424);
nand U27951 (N_27951,N_17227,N_12516);
and U27952 (N_27952,N_17617,N_15666);
nor U27953 (N_27953,N_11005,N_14371);
nand U27954 (N_27954,N_17015,N_10420);
and U27955 (N_27955,N_13813,N_10063);
xnor U27956 (N_27956,N_10340,N_15117);
xor U27957 (N_27957,N_10259,N_17497);
or U27958 (N_27958,N_13955,N_13203);
or U27959 (N_27959,N_10847,N_19020);
nand U27960 (N_27960,N_10897,N_12300);
xnor U27961 (N_27961,N_13129,N_17171);
nand U27962 (N_27962,N_19567,N_18228);
xnor U27963 (N_27963,N_16237,N_17404);
or U27964 (N_27964,N_12940,N_11392);
or U27965 (N_27965,N_14172,N_16903);
or U27966 (N_27966,N_12395,N_18522);
nand U27967 (N_27967,N_18286,N_17733);
or U27968 (N_27968,N_16387,N_12552);
nand U27969 (N_27969,N_14620,N_10318);
nor U27970 (N_27970,N_15195,N_19223);
xor U27971 (N_27971,N_10401,N_13092);
or U27972 (N_27972,N_10945,N_17869);
nand U27973 (N_27973,N_10563,N_10670);
nand U27974 (N_27974,N_10231,N_11416);
or U27975 (N_27975,N_18602,N_15385);
nor U27976 (N_27976,N_13382,N_11846);
xnor U27977 (N_27977,N_18205,N_18554);
xnor U27978 (N_27978,N_15434,N_19992);
and U27979 (N_27979,N_13276,N_16594);
and U27980 (N_27980,N_15914,N_13927);
nor U27981 (N_27981,N_19291,N_11319);
nand U27982 (N_27982,N_15832,N_11326);
and U27983 (N_27983,N_14795,N_18029);
or U27984 (N_27984,N_10084,N_18627);
xor U27985 (N_27985,N_10161,N_17460);
or U27986 (N_27986,N_11394,N_15934);
or U27987 (N_27987,N_10528,N_17334);
and U27988 (N_27988,N_17728,N_19437);
nand U27989 (N_27989,N_18157,N_16974);
nand U27990 (N_27990,N_13876,N_11058);
xor U27991 (N_27991,N_14716,N_10924);
nand U27992 (N_27992,N_14171,N_14052);
xnor U27993 (N_27993,N_16013,N_18104);
nand U27994 (N_27994,N_12672,N_14848);
nor U27995 (N_27995,N_10529,N_17318);
nand U27996 (N_27996,N_10624,N_13287);
nand U27997 (N_27997,N_18701,N_19885);
or U27998 (N_27998,N_18084,N_11233);
and U27999 (N_27999,N_10612,N_18184);
nand U28000 (N_28000,N_11976,N_17468);
and U28001 (N_28001,N_11919,N_12623);
nor U28002 (N_28002,N_10146,N_17412);
and U28003 (N_28003,N_15535,N_17883);
nand U28004 (N_28004,N_11146,N_16821);
and U28005 (N_28005,N_17886,N_12650);
nor U28006 (N_28006,N_11664,N_18048);
nor U28007 (N_28007,N_10049,N_15081);
nor U28008 (N_28008,N_12244,N_18769);
nor U28009 (N_28009,N_15981,N_16354);
xnor U28010 (N_28010,N_18122,N_15908);
nor U28011 (N_28011,N_12054,N_12747);
nor U28012 (N_28012,N_12315,N_18632);
or U28013 (N_28013,N_14846,N_18287);
and U28014 (N_28014,N_14094,N_14373);
xnor U28015 (N_28015,N_12931,N_13476);
xnor U28016 (N_28016,N_14765,N_15680);
nand U28017 (N_28017,N_12127,N_19081);
and U28018 (N_28018,N_17581,N_13817);
xor U28019 (N_28019,N_11571,N_19582);
nand U28020 (N_28020,N_14137,N_19366);
xor U28021 (N_28021,N_12625,N_17141);
or U28022 (N_28022,N_17360,N_16173);
or U28023 (N_28023,N_13339,N_13557);
nor U28024 (N_28024,N_17972,N_18541);
nand U28025 (N_28025,N_14537,N_14966);
or U28026 (N_28026,N_14698,N_11199);
xor U28027 (N_28027,N_10871,N_11984);
xnor U28028 (N_28028,N_16808,N_11420);
nand U28029 (N_28029,N_10006,N_19090);
nand U28030 (N_28030,N_17753,N_17853);
nand U28031 (N_28031,N_17744,N_14833);
nor U28032 (N_28032,N_12134,N_17410);
nand U28033 (N_28033,N_18938,N_14552);
and U28034 (N_28034,N_15689,N_17291);
xnor U28035 (N_28035,N_17922,N_11272);
or U28036 (N_28036,N_11229,N_16756);
and U28037 (N_28037,N_12080,N_15107);
xnor U28038 (N_28038,N_15359,N_19557);
nor U28039 (N_28039,N_12114,N_19031);
xor U28040 (N_28040,N_13329,N_10052);
or U28041 (N_28041,N_10963,N_19450);
or U28042 (N_28042,N_17827,N_19361);
nor U28043 (N_28043,N_17195,N_19717);
and U28044 (N_28044,N_10424,N_19969);
and U28045 (N_28045,N_19878,N_11216);
nand U28046 (N_28046,N_14093,N_17665);
nor U28047 (N_28047,N_14770,N_16399);
or U28048 (N_28048,N_13559,N_12816);
nor U28049 (N_28049,N_12496,N_16568);
xnor U28050 (N_28050,N_12694,N_15323);
or U28051 (N_28051,N_11357,N_14355);
and U28052 (N_28052,N_10572,N_10499);
xnor U28053 (N_28053,N_14813,N_13524);
xor U28054 (N_28054,N_12693,N_19103);
nand U28055 (N_28055,N_17066,N_12613);
nand U28056 (N_28056,N_13941,N_13219);
xnor U28057 (N_28057,N_10742,N_19729);
nor U28058 (N_28058,N_11911,N_12997);
or U28059 (N_28059,N_14637,N_11597);
xnor U28060 (N_28060,N_13592,N_15155);
xor U28061 (N_28061,N_10351,N_13119);
or U28062 (N_28062,N_12474,N_19541);
nand U28063 (N_28063,N_14423,N_12886);
nand U28064 (N_28064,N_19554,N_11855);
xor U28065 (N_28065,N_18990,N_15933);
xor U28066 (N_28066,N_15452,N_13706);
or U28067 (N_28067,N_19460,N_13574);
xnor U28068 (N_28068,N_15647,N_17535);
xnor U28069 (N_28069,N_13294,N_13614);
or U28070 (N_28070,N_13123,N_17642);
xnor U28071 (N_28071,N_15543,N_13190);
xor U28072 (N_28072,N_18265,N_16007);
xnor U28073 (N_28073,N_11149,N_18580);
or U28074 (N_28074,N_13580,N_11325);
or U28075 (N_28075,N_14301,N_19133);
and U28076 (N_28076,N_17387,N_17842);
nand U28077 (N_28077,N_16605,N_10419);
nand U28078 (N_28078,N_19065,N_12718);
nor U28079 (N_28079,N_16410,N_11884);
nand U28080 (N_28080,N_11941,N_15990);
xnor U28081 (N_28081,N_10596,N_10989);
or U28082 (N_28082,N_10259,N_15042);
and U28083 (N_28083,N_11260,N_17205);
xnor U28084 (N_28084,N_16337,N_17911);
nand U28085 (N_28085,N_18356,N_14148);
xor U28086 (N_28086,N_18733,N_15240);
nor U28087 (N_28087,N_12474,N_14666);
and U28088 (N_28088,N_12895,N_16087);
xnor U28089 (N_28089,N_16273,N_11025);
nand U28090 (N_28090,N_11505,N_14352);
and U28091 (N_28091,N_12612,N_15848);
nand U28092 (N_28092,N_12895,N_18130);
or U28093 (N_28093,N_15715,N_10223);
or U28094 (N_28094,N_11017,N_18253);
xor U28095 (N_28095,N_17971,N_18168);
xor U28096 (N_28096,N_16738,N_10269);
xor U28097 (N_28097,N_16364,N_12975);
nand U28098 (N_28098,N_15657,N_13901);
xor U28099 (N_28099,N_19513,N_17681);
or U28100 (N_28100,N_17200,N_14401);
nand U28101 (N_28101,N_17451,N_12038);
nor U28102 (N_28102,N_12080,N_17933);
and U28103 (N_28103,N_15082,N_15503);
and U28104 (N_28104,N_17430,N_16260);
or U28105 (N_28105,N_17714,N_15071);
and U28106 (N_28106,N_17256,N_11127);
nand U28107 (N_28107,N_13417,N_19227);
xor U28108 (N_28108,N_14121,N_16446);
and U28109 (N_28109,N_13650,N_19067);
or U28110 (N_28110,N_14489,N_14518);
nand U28111 (N_28111,N_12708,N_10206);
and U28112 (N_28112,N_14159,N_19875);
nand U28113 (N_28113,N_16682,N_15992);
and U28114 (N_28114,N_12973,N_17208);
and U28115 (N_28115,N_14717,N_16294);
xor U28116 (N_28116,N_12359,N_13379);
or U28117 (N_28117,N_14960,N_10985);
or U28118 (N_28118,N_16900,N_18050);
xnor U28119 (N_28119,N_15169,N_15959);
and U28120 (N_28120,N_16453,N_10075);
nand U28121 (N_28121,N_17467,N_13615);
and U28122 (N_28122,N_16930,N_12680);
nor U28123 (N_28123,N_15041,N_19111);
xor U28124 (N_28124,N_14604,N_15511);
xnor U28125 (N_28125,N_15200,N_16104);
nand U28126 (N_28126,N_18706,N_13383);
xor U28127 (N_28127,N_16802,N_19621);
nor U28128 (N_28128,N_15171,N_13659);
nand U28129 (N_28129,N_10620,N_13112);
or U28130 (N_28130,N_18848,N_17816);
xnor U28131 (N_28131,N_12675,N_10043);
and U28132 (N_28132,N_16397,N_17184);
nand U28133 (N_28133,N_10523,N_19747);
or U28134 (N_28134,N_11694,N_12284);
xnor U28135 (N_28135,N_15917,N_16995);
nand U28136 (N_28136,N_14409,N_14307);
nand U28137 (N_28137,N_11378,N_19245);
nand U28138 (N_28138,N_16052,N_17954);
nor U28139 (N_28139,N_13577,N_19763);
nand U28140 (N_28140,N_14396,N_10479);
nand U28141 (N_28141,N_17940,N_16372);
and U28142 (N_28142,N_14155,N_17014);
nor U28143 (N_28143,N_15233,N_15011);
nand U28144 (N_28144,N_16332,N_18301);
nand U28145 (N_28145,N_13158,N_17985);
or U28146 (N_28146,N_12693,N_10132);
and U28147 (N_28147,N_16904,N_16780);
xor U28148 (N_28148,N_13301,N_15630);
nor U28149 (N_28149,N_15907,N_17003);
nand U28150 (N_28150,N_15358,N_10605);
nand U28151 (N_28151,N_18890,N_11028);
or U28152 (N_28152,N_14501,N_19323);
nor U28153 (N_28153,N_15974,N_12058);
and U28154 (N_28154,N_18302,N_16535);
and U28155 (N_28155,N_18546,N_15805);
xor U28156 (N_28156,N_18687,N_15314);
nor U28157 (N_28157,N_19642,N_10667);
or U28158 (N_28158,N_16834,N_17687);
and U28159 (N_28159,N_19552,N_10806);
xnor U28160 (N_28160,N_19798,N_10997);
nand U28161 (N_28161,N_18595,N_10281);
nand U28162 (N_28162,N_15102,N_12811);
nand U28163 (N_28163,N_19943,N_14570);
or U28164 (N_28164,N_16090,N_13851);
nand U28165 (N_28165,N_11624,N_19514);
xor U28166 (N_28166,N_12772,N_17819);
or U28167 (N_28167,N_18004,N_16196);
nor U28168 (N_28168,N_16311,N_11934);
xor U28169 (N_28169,N_12396,N_19144);
and U28170 (N_28170,N_10259,N_15401);
nand U28171 (N_28171,N_12286,N_12970);
or U28172 (N_28172,N_14765,N_18782);
nor U28173 (N_28173,N_17479,N_10903);
and U28174 (N_28174,N_13026,N_10198);
and U28175 (N_28175,N_17068,N_10987);
nor U28176 (N_28176,N_18356,N_11872);
xor U28177 (N_28177,N_18886,N_11434);
nand U28178 (N_28178,N_17159,N_17653);
nor U28179 (N_28179,N_13976,N_18045);
nor U28180 (N_28180,N_19041,N_10060);
xnor U28181 (N_28181,N_13142,N_16201);
nor U28182 (N_28182,N_18131,N_16458);
xnor U28183 (N_28183,N_18182,N_16753);
nand U28184 (N_28184,N_19213,N_12340);
and U28185 (N_28185,N_18503,N_17588);
xor U28186 (N_28186,N_10577,N_13838);
or U28187 (N_28187,N_14144,N_13746);
and U28188 (N_28188,N_11642,N_18020);
and U28189 (N_28189,N_11650,N_12879);
or U28190 (N_28190,N_17561,N_18039);
and U28191 (N_28191,N_14016,N_11290);
or U28192 (N_28192,N_18459,N_10651);
xnor U28193 (N_28193,N_19850,N_13175);
nor U28194 (N_28194,N_11429,N_11855);
nand U28195 (N_28195,N_10621,N_17342);
or U28196 (N_28196,N_16808,N_12502);
or U28197 (N_28197,N_12782,N_10922);
nor U28198 (N_28198,N_17298,N_15907);
xor U28199 (N_28199,N_15508,N_13493);
xnor U28200 (N_28200,N_12326,N_16264);
nand U28201 (N_28201,N_19406,N_10950);
xor U28202 (N_28202,N_10453,N_15467);
nand U28203 (N_28203,N_13603,N_11066);
nand U28204 (N_28204,N_19873,N_11690);
nand U28205 (N_28205,N_10392,N_12802);
nor U28206 (N_28206,N_12353,N_14728);
or U28207 (N_28207,N_18628,N_16188);
nand U28208 (N_28208,N_17612,N_19588);
or U28209 (N_28209,N_13933,N_17851);
nand U28210 (N_28210,N_14096,N_16093);
nor U28211 (N_28211,N_12968,N_10827);
xor U28212 (N_28212,N_10285,N_15129);
and U28213 (N_28213,N_12925,N_19834);
xor U28214 (N_28214,N_13900,N_10908);
and U28215 (N_28215,N_11735,N_11176);
or U28216 (N_28216,N_18959,N_16434);
nor U28217 (N_28217,N_10939,N_17368);
nor U28218 (N_28218,N_13031,N_11092);
and U28219 (N_28219,N_15461,N_14845);
or U28220 (N_28220,N_13115,N_13964);
and U28221 (N_28221,N_13547,N_12297);
nand U28222 (N_28222,N_17917,N_18953);
nand U28223 (N_28223,N_12857,N_11118);
or U28224 (N_28224,N_15728,N_19060);
nor U28225 (N_28225,N_18748,N_12626);
and U28226 (N_28226,N_18820,N_17384);
nand U28227 (N_28227,N_18125,N_17386);
and U28228 (N_28228,N_19828,N_18125);
nor U28229 (N_28229,N_14594,N_18460);
nor U28230 (N_28230,N_18765,N_10384);
nor U28231 (N_28231,N_10390,N_13752);
xor U28232 (N_28232,N_10963,N_15082);
nor U28233 (N_28233,N_10294,N_15739);
xnor U28234 (N_28234,N_11824,N_12047);
nor U28235 (N_28235,N_11480,N_18646);
xor U28236 (N_28236,N_19450,N_16413);
nor U28237 (N_28237,N_18920,N_12661);
or U28238 (N_28238,N_17069,N_18198);
nand U28239 (N_28239,N_15441,N_15674);
and U28240 (N_28240,N_10386,N_14754);
nand U28241 (N_28241,N_10869,N_12607);
xor U28242 (N_28242,N_15446,N_11921);
nor U28243 (N_28243,N_18740,N_16135);
and U28244 (N_28244,N_17329,N_19842);
nand U28245 (N_28245,N_12530,N_12713);
nand U28246 (N_28246,N_17111,N_12891);
nor U28247 (N_28247,N_13434,N_16505);
nand U28248 (N_28248,N_16708,N_15617);
and U28249 (N_28249,N_15797,N_11789);
and U28250 (N_28250,N_17743,N_13470);
xor U28251 (N_28251,N_16577,N_18242);
or U28252 (N_28252,N_12796,N_15868);
or U28253 (N_28253,N_18482,N_13566);
or U28254 (N_28254,N_15403,N_10848);
nor U28255 (N_28255,N_18581,N_14856);
or U28256 (N_28256,N_18020,N_11353);
xor U28257 (N_28257,N_18179,N_14512);
nand U28258 (N_28258,N_14588,N_19187);
xor U28259 (N_28259,N_14925,N_15171);
or U28260 (N_28260,N_12988,N_14470);
nor U28261 (N_28261,N_13250,N_11372);
and U28262 (N_28262,N_16806,N_13959);
and U28263 (N_28263,N_19369,N_12127);
and U28264 (N_28264,N_12220,N_18615);
xnor U28265 (N_28265,N_14331,N_10182);
xnor U28266 (N_28266,N_10213,N_12999);
and U28267 (N_28267,N_11579,N_13820);
nand U28268 (N_28268,N_16234,N_12040);
or U28269 (N_28269,N_18760,N_14193);
xnor U28270 (N_28270,N_11721,N_19505);
or U28271 (N_28271,N_12644,N_15905);
nand U28272 (N_28272,N_12162,N_19123);
and U28273 (N_28273,N_17172,N_18289);
xor U28274 (N_28274,N_11861,N_10292);
xor U28275 (N_28275,N_15065,N_14204);
nor U28276 (N_28276,N_17701,N_12269);
xnor U28277 (N_28277,N_13654,N_11910);
or U28278 (N_28278,N_11521,N_10739);
nor U28279 (N_28279,N_14442,N_17643);
xor U28280 (N_28280,N_10047,N_10021);
xor U28281 (N_28281,N_17175,N_19650);
nor U28282 (N_28282,N_11177,N_14005);
and U28283 (N_28283,N_16872,N_11848);
and U28284 (N_28284,N_12680,N_12476);
xnor U28285 (N_28285,N_17954,N_18880);
and U28286 (N_28286,N_17535,N_17613);
nor U28287 (N_28287,N_11082,N_14654);
or U28288 (N_28288,N_10260,N_13421);
and U28289 (N_28289,N_11215,N_16082);
nor U28290 (N_28290,N_12833,N_13546);
and U28291 (N_28291,N_19944,N_11249);
nand U28292 (N_28292,N_17185,N_15106);
xnor U28293 (N_28293,N_15071,N_17847);
and U28294 (N_28294,N_18249,N_17819);
xnor U28295 (N_28295,N_18703,N_15073);
xnor U28296 (N_28296,N_17324,N_14680);
xor U28297 (N_28297,N_12637,N_13802);
and U28298 (N_28298,N_17277,N_11869);
nand U28299 (N_28299,N_16685,N_17335);
xnor U28300 (N_28300,N_16430,N_17421);
xor U28301 (N_28301,N_18474,N_17976);
xor U28302 (N_28302,N_11713,N_13544);
or U28303 (N_28303,N_19819,N_12967);
and U28304 (N_28304,N_14853,N_12422);
and U28305 (N_28305,N_10516,N_15790);
nor U28306 (N_28306,N_18787,N_13812);
or U28307 (N_28307,N_19475,N_14098);
and U28308 (N_28308,N_14266,N_16606);
nand U28309 (N_28309,N_17756,N_13325);
xor U28310 (N_28310,N_10823,N_15033);
nor U28311 (N_28311,N_12917,N_18629);
nand U28312 (N_28312,N_10476,N_16171);
or U28313 (N_28313,N_15044,N_12176);
or U28314 (N_28314,N_16140,N_10802);
xor U28315 (N_28315,N_16200,N_18456);
or U28316 (N_28316,N_18158,N_15558);
and U28317 (N_28317,N_11438,N_18170);
xor U28318 (N_28318,N_13468,N_13737);
xnor U28319 (N_28319,N_18313,N_18056);
xor U28320 (N_28320,N_15541,N_18462);
nor U28321 (N_28321,N_14023,N_13874);
or U28322 (N_28322,N_13736,N_18602);
and U28323 (N_28323,N_15082,N_10990);
nor U28324 (N_28324,N_10381,N_14221);
or U28325 (N_28325,N_17654,N_11820);
or U28326 (N_28326,N_10944,N_16498);
nand U28327 (N_28327,N_16182,N_18481);
or U28328 (N_28328,N_16219,N_13371);
xor U28329 (N_28329,N_10391,N_13619);
and U28330 (N_28330,N_17385,N_14130);
and U28331 (N_28331,N_12271,N_11822);
xor U28332 (N_28332,N_19007,N_18707);
or U28333 (N_28333,N_13369,N_16141);
nor U28334 (N_28334,N_17954,N_10794);
xor U28335 (N_28335,N_18149,N_13489);
and U28336 (N_28336,N_15701,N_15654);
nand U28337 (N_28337,N_10807,N_15853);
nor U28338 (N_28338,N_17820,N_15878);
xor U28339 (N_28339,N_10594,N_11447);
or U28340 (N_28340,N_17793,N_17002);
xor U28341 (N_28341,N_10557,N_13976);
and U28342 (N_28342,N_16558,N_19089);
or U28343 (N_28343,N_12988,N_15558);
or U28344 (N_28344,N_18154,N_14687);
nor U28345 (N_28345,N_19980,N_14255);
nor U28346 (N_28346,N_10625,N_17879);
nand U28347 (N_28347,N_18814,N_18282);
xnor U28348 (N_28348,N_14422,N_13471);
nor U28349 (N_28349,N_12928,N_18264);
nor U28350 (N_28350,N_12672,N_11987);
xnor U28351 (N_28351,N_14333,N_10430);
nor U28352 (N_28352,N_19148,N_12999);
nor U28353 (N_28353,N_19455,N_10838);
nand U28354 (N_28354,N_15582,N_11191);
and U28355 (N_28355,N_18489,N_19981);
xor U28356 (N_28356,N_19532,N_15049);
or U28357 (N_28357,N_10481,N_13068);
nand U28358 (N_28358,N_19443,N_11046);
xor U28359 (N_28359,N_19673,N_18850);
or U28360 (N_28360,N_16759,N_11066);
xor U28361 (N_28361,N_11989,N_10359);
or U28362 (N_28362,N_17841,N_16212);
nor U28363 (N_28363,N_14664,N_14584);
or U28364 (N_28364,N_12332,N_11988);
and U28365 (N_28365,N_19618,N_15746);
or U28366 (N_28366,N_14848,N_13311);
nand U28367 (N_28367,N_16961,N_17999);
xnor U28368 (N_28368,N_19132,N_17525);
nor U28369 (N_28369,N_13594,N_19628);
or U28370 (N_28370,N_12539,N_15258);
xnor U28371 (N_28371,N_11965,N_17314);
xor U28372 (N_28372,N_10772,N_14833);
and U28373 (N_28373,N_10423,N_12534);
xor U28374 (N_28374,N_19430,N_10685);
or U28375 (N_28375,N_14154,N_11557);
and U28376 (N_28376,N_13029,N_18840);
or U28377 (N_28377,N_10412,N_13704);
xnor U28378 (N_28378,N_13778,N_17617);
and U28379 (N_28379,N_11775,N_16938);
or U28380 (N_28380,N_16528,N_16135);
and U28381 (N_28381,N_16160,N_18500);
nand U28382 (N_28382,N_12817,N_15341);
nor U28383 (N_28383,N_17086,N_15852);
or U28384 (N_28384,N_16807,N_10151);
and U28385 (N_28385,N_12376,N_11375);
xor U28386 (N_28386,N_12791,N_11223);
or U28387 (N_28387,N_16004,N_11180);
nand U28388 (N_28388,N_10707,N_12379);
xnor U28389 (N_28389,N_14370,N_12533);
nor U28390 (N_28390,N_11304,N_14873);
nor U28391 (N_28391,N_10018,N_14605);
and U28392 (N_28392,N_16195,N_12758);
nand U28393 (N_28393,N_17502,N_17202);
and U28394 (N_28394,N_12890,N_16373);
nor U28395 (N_28395,N_10619,N_14654);
and U28396 (N_28396,N_14404,N_18529);
xor U28397 (N_28397,N_18890,N_15629);
xor U28398 (N_28398,N_13198,N_15841);
nand U28399 (N_28399,N_15437,N_10442);
nor U28400 (N_28400,N_16029,N_13473);
nand U28401 (N_28401,N_12667,N_10513);
xnor U28402 (N_28402,N_18952,N_13880);
xnor U28403 (N_28403,N_14905,N_14991);
or U28404 (N_28404,N_16230,N_15990);
nand U28405 (N_28405,N_18947,N_16636);
nor U28406 (N_28406,N_17541,N_19046);
or U28407 (N_28407,N_16221,N_16102);
or U28408 (N_28408,N_13975,N_17192);
and U28409 (N_28409,N_18175,N_10252);
xnor U28410 (N_28410,N_12230,N_10760);
or U28411 (N_28411,N_18855,N_12028);
nand U28412 (N_28412,N_12685,N_16028);
xor U28413 (N_28413,N_14960,N_13891);
and U28414 (N_28414,N_19415,N_11794);
nand U28415 (N_28415,N_11471,N_11439);
and U28416 (N_28416,N_10168,N_19561);
or U28417 (N_28417,N_12014,N_13290);
and U28418 (N_28418,N_11942,N_19512);
and U28419 (N_28419,N_14792,N_16466);
or U28420 (N_28420,N_18490,N_12680);
nor U28421 (N_28421,N_13272,N_12150);
xor U28422 (N_28422,N_16815,N_18535);
and U28423 (N_28423,N_12596,N_12303);
or U28424 (N_28424,N_18090,N_11184);
xnor U28425 (N_28425,N_13667,N_19537);
nor U28426 (N_28426,N_18682,N_16522);
xor U28427 (N_28427,N_11471,N_14481);
or U28428 (N_28428,N_17794,N_15898);
nor U28429 (N_28429,N_16392,N_14228);
or U28430 (N_28430,N_13279,N_14037);
and U28431 (N_28431,N_10031,N_14577);
xor U28432 (N_28432,N_18663,N_12835);
nor U28433 (N_28433,N_19314,N_17482);
and U28434 (N_28434,N_19176,N_14010);
nor U28435 (N_28435,N_10812,N_11920);
xor U28436 (N_28436,N_12483,N_19656);
or U28437 (N_28437,N_19120,N_15013);
and U28438 (N_28438,N_16092,N_12280);
or U28439 (N_28439,N_15459,N_15876);
or U28440 (N_28440,N_19437,N_14830);
nor U28441 (N_28441,N_10583,N_17792);
or U28442 (N_28442,N_17685,N_17256);
or U28443 (N_28443,N_11434,N_13158);
nor U28444 (N_28444,N_15018,N_15348);
xor U28445 (N_28445,N_11098,N_12260);
and U28446 (N_28446,N_12922,N_18474);
nand U28447 (N_28447,N_17891,N_19178);
or U28448 (N_28448,N_11585,N_10457);
and U28449 (N_28449,N_18148,N_13225);
xor U28450 (N_28450,N_11635,N_18499);
xor U28451 (N_28451,N_10732,N_19608);
nand U28452 (N_28452,N_15812,N_17164);
xor U28453 (N_28453,N_13251,N_12348);
and U28454 (N_28454,N_12212,N_14166);
and U28455 (N_28455,N_17323,N_15282);
and U28456 (N_28456,N_16094,N_16582);
xor U28457 (N_28457,N_19966,N_16198);
nor U28458 (N_28458,N_13720,N_10011);
xor U28459 (N_28459,N_15428,N_11176);
xnor U28460 (N_28460,N_19487,N_19881);
nand U28461 (N_28461,N_15587,N_11488);
and U28462 (N_28462,N_12591,N_11202);
or U28463 (N_28463,N_11379,N_12242);
and U28464 (N_28464,N_15238,N_10998);
nand U28465 (N_28465,N_19257,N_11334);
nand U28466 (N_28466,N_17294,N_12823);
xnor U28467 (N_28467,N_15485,N_13086);
xnor U28468 (N_28468,N_12954,N_14436);
and U28469 (N_28469,N_11710,N_17905);
and U28470 (N_28470,N_13704,N_15318);
nand U28471 (N_28471,N_13660,N_16149);
xnor U28472 (N_28472,N_17492,N_17681);
nor U28473 (N_28473,N_13326,N_17207);
or U28474 (N_28474,N_13958,N_14979);
and U28475 (N_28475,N_16563,N_17167);
nand U28476 (N_28476,N_11417,N_14970);
nand U28477 (N_28477,N_17164,N_17893);
xnor U28478 (N_28478,N_11566,N_14766);
nand U28479 (N_28479,N_15352,N_13298);
or U28480 (N_28480,N_10343,N_13185);
nor U28481 (N_28481,N_12657,N_11773);
and U28482 (N_28482,N_18185,N_13844);
and U28483 (N_28483,N_18860,N_14853);
or U28484 (N_28484,N_13755,N_11886);
and U28485 (N_28485,N_19756,N_15561);
and U28486 (N_28486,N_19965,N_16798);
and U28487 (N_28487,N_11184,N_16643);
and U28488 (N_28488,N_11335,N_19956);
nand U28489 (N_28489,N_11638,N_11731);
nor U28490 (N_28490,N_10188,N_13528);
nor U28491 (N_28491,N_18907,N_10841);
and U28492 (N_28492,N_16142,N_18970);
nand U28493 (N_28493,N_10013,N_16262);
or U28494 (N_28494,N_15404,N_16298);
or U28495 (N_28495,N_12258,N_11569);
nand U28496 (N_28496,N_15770,N_15526);
and U28497 (N_28497,N_15780,N_18632);
nand U28498 (N_28498,N_15258,N_19249);
nand U28499 (N_28499,N_14597,N_18935);
and U28500 (N_28500,N_11141,N_14327);
nor U28501 (N_28501,N_15389,N_17640);
and U28502 (N_28502,N_10277,N_18354);
xnor U28503 (N_28503,N_16983,N_11377);
nand U28504 (N_28504,N_12340,N_17431);
or U28505 (N_28505,N_19464,N_14971);
xor U28506 (N_28506,N_17506,N_19271);
and U28507 (N_28507,N_13011,N_11593);
xnor U28508 (N_28508,N_19266,N_19374);
xnor U28509 (N_28509,N_19399,N_14766);
xor U28510 (N_28510,N_19301,N_12208);
xnor U28511 (N_28511,N_16306,N_11678);
nand U28512 (N_28512,N_11651,N_19150);
nor U28513 (N_28513,N_12210,N_12163);
nor U28514 (N_28514,N_11879,N_15772);
nand U28515 (N_28515,N_15877,N_11016);
and U28516 (N_28516,N_15350,N_17081);
and U28517 (N_28517,N_10862,N_12825);
xnor U28518 (N_28518,N_14594,N_17721);
or U28519 (N_28519,N_19195,N_11345);
or U28520 (N_28520,N_15240,N_14270);
and U28521 (N_28521,N_11663,N_16094);
or U28522 (N_28522,N_14872,N_18124);
nand U28523 (N_28523,N_14461,N_14674);
nor U28524 (N_28524,N_17064,N_11198);
nand U28525 (N_28525,N_11612,N_17789);
and U28526 (N_28526,N_12400,N_11337);
and U28527 (N_28527,N_19114,N_17546);
nand U28528 (N_28528,N_17242,N_14305);
nand U28529 (N_28529,N_13960,N_10573);
xnor U28530 (N_28530,N_12870,N_17874);
nand U28531 (N_28531,N_10497,N_10391);
nand U28532 (N_28532,N_16449,N_16117);
xor U28533 (N_28533,N_10352,N_16589);
or U28534 (N_28534,N_15743,N_18165);
nand U28535 (N_28535,N_10140,N_16363);
nor U28536 (N_28536,N_18113,N_13032);
nor U28537 (N_28537,N_18355,N_10380);
or U28538 (N_28538,N_12523,N_14942);
nand U28539 (N_28539,N_12358,N_12396);
and U28540 (N_28540,N_19820,N_16227);
nand U28541 (N_28541,N_16420,N_16846);
xnor U28542 (N_28542,N_19177,N_11392);
nor U28543 (N_28543,N_13062,N_14918);
xor U28544 (N_28544,N_10328,N_13374);
and U28545 (N_28545,N_13327,N_17205);
xnor U28546 (N_28546,N_15479,N_15991);
nand U28547 (N_28547,N_10617,N_19634);
or U28548 (N_28548,N_12349,N_10538);
xor U28549 (N_28549,N_17816,N_16355);
nor U28550 (N_28550,N_14559,N_12392);
or U28551 (N_28551,N_15027,N_11702);
or U28552 (N_28552,N_19991,N_14770);
and U28553 (N_28553,N_10770,N_15450);
or U28554 (N_28554,N_15614,N_10680);
nor U28555 (N_28555,N_17228,N_18128);
xor U28556 (N_28556,N_15273,N_10612);
nor U28557 (N_28557,N_10310,N_19202);
xnor U28558 (N_28558,N_16216,N_13006);
and U28559 (N_28559,N_16158,N_16878);
nor U28560 (N_28560,N_13756,N_16191);
xnor U28561 (N_28561,N_16100,N_13873);
xor U28562 (N_28562,N_19084,N_16506);
xor U28563 (N_28563,N_10544,N_15390);
and U28564 (N_28564,N_19827,N_12318);
and U28565 (N_28565,N_19894,N_18394);
or U28566 (N_28566,N_10467,N_16622);
or U28567 (N_28567,N_16223,N_15120);
xnor U28568 (N_28568,N_13105,N_19774);
nand U28569 (N_28569,N_14134,N_14438);
xnor U28570 (N_28570,N_16511,N_12850);
nand U28571 (N_28571,N_14578,N_14689);
and U28572 (N_28572,N_13894,N_11535);
or U28573 (N_28573,N_18137,N_19046);
xnor U28574 (N_28574,N_18708,N_12008);
and U28575 (N_28575,N_10594,N_11518);
xor U28576 (N_28576,N_12532,N_15717);
and U28577 (N_28577,N_14913,N_11298);
nand U28578 (N_28578,N_10587,N_17353);
xnor U28579 (N_28579,N_19657,N_18808);
or U28580 (N_28580,N_15635,N_15617);
and U28581 (N_28581,N_10733,N_10947);
nand U28582 (N_28582,N_19670,N_19427);
xnor U28583 (N_28583,N_19633,N_10784);
xor U28584 (N_28584,N_10390,N_14814);
nand U28585 (N_28585,N_11981,N_18538);
nand U28586 (N_28586,N_10625,N_11519);
nor U28587 (N_28587,N_13931,N_16563);
or U28588 (N_28588,N_16487,N_17143);
xnor U28589 (N_28589,N_11963,N_13649);
and U28590 (N_28590,N_17861,N_13023);
xnor U28591 (N_28591,N_16944,N_10260);
and U28592 (N_28592,N_13682,N_12080);
and U28593 (N_28593,N_15496,N_17287);
nor U28594 (N_28594,N_18009,N_11079);
or U28595 (N_28595,N_18169,N_13479);
nor U28596 (N_28596,N_19815,N_11916);
nand U28597 (N_28597,N_12721,N_16853);
and U28598 (N_28598,N_14173,N_16681);
nor U28599 (N_28599,N_14016,N_17589);
nand U28600 (N_28600,N_12257,N_15651);
and U28601 (N_28601,N_13896,N_18797);
nor U28602 (N_28602,N_13861,N_17920);
or U28603 (N_28603,N_13400,N_19099);
or U28604 (N_28604,N_12593,N_19502);
nand U28605 (N_28605,N_19325,N_15461);
and U28606 (N_28606,N_19286,N_14584);
or U28607 (N_28607,N_17014,N_12542);
nor U28608 (N_28608,N_13541,N_14332);
xnor U28609 (N_28609,N_15459,N_14134);
nor U28610 (N_28610,N_11035,N_15521);
xnor U28611 (N_28611,N_12855,N_10404);
xor U28612 (N_28612,N_15449,N_15387);
nor U28613 (N_28613,N_13563,N_19361);
or U28614 (N_28614,N_15475,N_10056);
xor U28615 (N_28615,N_10371,N_10860);
xor U28616 (N_28616,N_11318,N_19779);
or U28617 (N_28617,N_11086,N_15516);
and U28618 (N_28618,N_19442,N_14923);
or U28619 (N_28619,N_10646,N_14746);
or U28620 (N_28620,N_15549,N_19537);
and U28621 (N_28621,N_19607,N_16024);
or U28622 (N_28622,N_12692,N_14076);
xnor U28623 (N_28623,N_19761,N_11825);
nor U28624 (N_28624,N_12181,N_18197);
xor U28625 (N_28625,N_19097,N_11357);
and U28626 (N_28626,N_16172,N_17033);
or U28627 (N_28627,N_13591,N_17929);
xnor U28628 (N_28628,N_15644,N_12332);
or U28629 (N_28629,N_18852,N_18961);
or U28630 (N_28630,N_13631,N_19927);
nand U28631 (N_28631,N_12085,N_11128);
nand U28632 (N_28632,N_16974,N_10294);
xnor U28633 (N_28633,N_15417,N_15554);
xor U28634 (N_28634,N_14754,N_17086);
nor U28635 (N_28635,N_14087,N_15713);
nand U28636 (N_28636,N_10963,N_15217);
or U28637 (N_28637,N_14578,N_16357);
and U28638 (N_28638,N_10910,N_13412);
and U28639 (N_28639,N_19517,N_18607);
and U28640 (N_28640,N_14627,N_16786);
or U28641 (N_28641,N_17122,N_17163);
nor U28642 (N_28642,N_11414,N_13206);
or U28643 (N_28643,N_12351,N_18192);
nor U28644 (N_28644,N_15763,N_14658);
or U28645 (N_28645,N_15503,N_13560);
xor U28646 (N_28646,N_16825,N_14094);
nand U28647 (N_28647,N_14828,N_17013);
and U28648 (N_28648,N_13403,N_14442);
or U28649 (N_28649,N_17846,N_13641);
and U28650 (N_28650,N_19303,N_15207);
nor U28651 (N_28651,N_18557,N_12871);
xnor U28652 (N_28652,N_11984,N_19127);
and U28653 (N_28653,N_17248,N_13180);
and U28654 (N_28654,N_15196,N_16764);
and U28655 (N_28655,N_14107,N_15469);
nand U28656 (N_28656,N_14077,N_19266);
nand U28657 (N_28657,N_17779,N_13019);
or U28658 (N_28658,N_14725,N_15663);
xor U28659 (N_28659,N_14173,N_14595);
or U28660 (N_28660,N_16871,N_10596);
or U28661 (N_28661,N_19211,N_19140);
nand U28662 (N_28662,N_13223,N_13217);
xor U28663 (N_28663,N_15003,N_15463);
or U28664 (N_28664,N_12018,N_16736);
nor U28665 (N_28665,N_14335,N_15964);
nor U28666 (N_28666,N_14378,N_12285);
or U28667 (N_28667,N_11673,N_10198);
and U28668 (N_28668,N_10791,N_18812);
nand U28669 (N_28669,N_13530,N_16758);
nand U28670 (N_28670,N_19087,N_19464);
nand U28671 (N_28671,N_17388,N_19128);
nor U28672 (N_28672,N_16707,N_18913);
and U28673 (N_28673,N_10311,N_17283);
nor U28674 (N_28674,N_18556,N_16638);
and U28675 (N_28675,N_14805,N_16046);
or U28676 (N_28676,N_11410,N_17932);
xor U28677 (N_28677,N_10738,N_13696);
nand U28678 (N_28678,N_16560,N_13257);
or U28679 (N_28679,N_10379,N_15707);
or U28680 (N_28680,N_12737,N_10708);
nor U28681 (N_28681,N_15141,N_14373);
nor U28682 (N_28682,N_18429,N_13352);
or U28683 (N_28683,N_14947,N_11943);
xor U28684 (N_28684,N_16774,N_19294);
xnor U28685 (N_28685,N_17277,N_19788);
or U28686 (N_28686,N_19960,N_13021);
xnor U28687 (N_28687,N_11955,N_15981);
nor U28688 (N_28688,N_13914,N_18075);
and U28689 (N_28689,N_10914,N_18125);
and U28690 (N_28690,N_10042,N_15650);
nand U28691 (N_28691,N_13762,N_16052);
xor U28692 (N_28692,N_13473,N_11564);
nand U28693 (N_28693,N_19968,N_16367);
and U28694 (N_28694,N_14065,N_17213);
xor U28695 (N_28695,N_11413,N_14145);
nor U28696 (N_28696,N_18925,N_17255);
and U28697 (N_28697,N_10578,N_16594);
xnor U28698 (N_28698,N_12833,N_18157);
xor U28699 (N_28699,N_12874,N_13419);
nand U28700 (N_28700,N_10027,N_15058);
and U28701 (N_28701,N_11545,N_12774);
and U28702 (N_28702,N_16672,N_15146);
and U28703 (N_28703,N_17525,N_12442);
nand U28704 (N_28704,N_11938,N_12470);
xnor U28705 (N_28705,N_13647,N_12048);
or U28706 (N_28706,N_15276,N_13689);
nand U28707 (N_28707,N_15724,N_10384);
xor U28708 (N_28708,N_15586,N_16545);
xnor U28709 (N_28709,N_17750,N_15097);
or U28710 (N_28710,N_19529,N_17265);
nor U28711 (N_28711,N_14706,N_14295);
nand U28712 (N_28712,N_16675,N_15498);
nand U28713 (N_28713,N_17539,N_15594);
and U28714 (N_28714,N_11883,N_12374);
xor U28715 (N_28715,N_11301,N_14797);
nor U28716 (N_28716,N_14656,N_14332);
nand U28717 (N_28717,N_18963,N_19939);
nor U28718 (N_28718,N_12472,N_11199);
xor U28719 (N_28719,N_12429,N_11631);
or U28720 (N_28720,N_19433,N_15771);
nor U28721 (N_28721,N_19604,N_15161);
xnor U28722 (N_28722,N_10266,N_19787);
nor U28723 (N_28723,N_18832,N_15281);
or U28724 (N_28724,N_19735,N_14770);
or U28725 (N_28725,N_10427,N_17360);
nand U28726 (N_28726,N_19310,N_11646);
xor U28727 (N_28727,N_12667,N_17625);
nor U28728 (N_28728,N_19754,N_18720);
xnor U28729 (N_28729,N_15884,N_17409);
or U28730 (N_28730,N_18402,N_13363);
and U28731 (N_28731,N_18938,N_17040);
and U28732 (N_28732,N_10804,N_17450);
or U28733 (N_28733,N_18681,N_10049);
and U28734 (N_28734,N_16508,N_13915);
nand U28735 (N_28735,N_13663,N_11999);
or U28736 (N_28736,N_17760,N_10372);
nor U28737 (N_28737,N_19269,N_14717);
nand U28738 (N_28738,N_13441,N_10629);
nor U28739 (N_28739,N_19423,N_10519);
xor U28740 (N_28740,N_13567,N_10717);
nand U28741 (N_28741,N_18286,N_17313);
nor U28742 (N_28742,N_18522,N_19343);
nand U28743 (N_28743,N_10237,N_15364);
nor U28744 (N_28744,N_13225,N_19957);
nor U28745 (N_28745,N_18572,N_17532);
nand U28746 (N_28746,N_11652,N_18117);
nand U28747 (N_28747,N_11871,N_16193);
or U28748 (N_28748,N_19209,N_12027);
nand U28749 (N_28749,N_17488,N_15774);
nand U28750 (N_28750,N_19318,N_18436);
nand U28751 (N_28751,N_15436,N_11079);
and U28752 (N_28752,N_17628,N_13461);
nand U28753 (N_28753,N_12401,N_17291);
xor U28754 (N_28754,N_15213,N_19930);
or U28755 (N_28755,N_19188,N_19992);
nand U28756 (N_28756,N_13768,N_16015);
nor U28757 (N_28757,N_11057,N_12195);
nand U28758 (N_28758,N_17793,N_11090);
or U28759 (N_28759,N_16249,N_18559);
nand U28760 (N_28760,N_17714,N_19645);
xor U28761 (N_28761,N_17599,N_10629);
xor U28762 (N_28762,N_14962,N_11630);
and U28763 (N_28763,N_12556,N_19402);
nand U28764 (N_28764,N_11777,N_18089);
nand U28765 (N_28765,N_15898,N_14515);
xor U28766 (N_28766,N_11880,N_12367);
nor U28767 (N_28767,N_14159,N_15220);
xnor U28768 (N_28768,N_16644,N_16565);
or U28769 (N_28769,N_16957,N_17984);
nor U28770 (N_28770,N_14832,N_13534);
nand U28771 (N_28771,N_14382,N_18818);
or U28772 (N_28772,N_14095,N_16396);
nand U28773 (N_28773,N_10638,N_16428);
nand U28774 (N_28774,N_10898,N_18560);
nand U28775 (N_28775,N_15624,N_14502);
or U28776 (N_28776,N_10189,N_19315);
xor U28777 (N_28777,N_14007,N_10837);
nand U28778 (N_28778,N_18292,N_10280);
nand U28779 (N_28779,N_14113,N_16878);
or U28780 (N_28780,N_17468,N_18997);
and U28781 (N_28781,N_18574,N_10599);
nand U28782 (N_28782,N_14699,N_12102);
and U28783 (N_28783,N_17438,N_13780);
xor U28784 (N_28784,N_11528,N_17192);
xor U28785 (N_28785,N_18029,N_13599);
and U28786 (N_28786,N_12408,N_18513);
or U28787 (N_28787,N_11201,N_11460);
or U28788 (N_28788,N_14787,N_16374);
nand U28789 (N_28789,N_17194,N_19265);
or U28790 (N_28790,N_11879,N_17493);
xor U28791 (N_28791,N_12447,N_17234);
or U28792 (N_28792,N_10729,N_16655);
nor U28793 (N_28793,N_10709,N_14205);
nand U28794 (N_28794,N_11546,N_16384);
or U28795 (N_28795,N_13574,N_15617);
or U28796 (N_28796,N_13419,N_15747);
and U28797 (N_28797,N_15432,N_18336);
nand U28798 (N_28798,N_15172,N_15867);
nand U28799 (N_28799,N_19853,N_17053);
xor U28800 (N_28800,N_10863,N_19253);
xnor U28801 (N_28801,N_13021,N_15711);
and U28802 (N_28802,N_14265,N_14141);
and U28803 (N_28803,N_14343,N_15174);
xnor U28804 (N_28804,N_11927,N_16309);
nor U28805 (N_28805,N_12805,N_14951);
and U28806 (N_28806,N_16959,N_13609);
and U28807 (N_28807,N_11714,N_16894);
and U28808 (N_28808,N_16991,N_17821);
nand U28809 (N_28809,N_15421,N_16245);
or U28810 (N_28810,N_16617,N_16370);
nor U28811 (N_28811,N_14132,N_17108);
and U28812 (N_28812,N_11606,N_19019);
nor U28813 (N_28813,N_19085,N_12172);
or U28814 (N_28814,N_17161,N_17995);
xor U28815 (N_28815,N_15519,N_19062);
nand U28816 (N_28816,N_16301,N_15410);
or U28817 (N_28817,N_12002,N_11391);
or U28818 (N_28818,N_14078,N_16216);
and U28819 (N_28819,N_14818,N_11106);
or U28820 (N_28820,N_10681,N_14501);
or U28821 (N_28821,N_19868,N_12711);
nand U28822 (N_28822,N_19167,N_17202);
and U28823 (N_28823,N_12178,N_11181);
xnor U28824 (N_28824,N_14509,N_18402);
nor U28825 (N_28825,N_14703,N_10304);
xor U28826 (N_28826,N_17429,N_10703);
xor U28827 (N_28827,N_18110,N_11666);
or U28828 (N_28828,N_19089,N_14252);
xor U28829 (N_28829,N_16739,N_11914);
and U28830 (N_28830,N_15436,N_16499);
nand U28831 (N_28831,N_16676,N_11008);
nor U28832 (N_28832,N_11060,N_13054);
nor U28833 (N_28833,N_17408,N_12319);
and U28834 (N_28834,N_14922,N_17191);
xnor U28835 (N_28835,N_11670,N_11029);
or U28836 (N_28836,N_10589,N_12544);
or U28837 (N_28837,N_17546,N_18205);
nor U28838 (N_28838,N_17637,N_11949);
or U28839 (N_28839,N_14416,N_13682);
nor U28840 (N_28840,N_14290,N_12828);
and U28841 (N_28841,N_14682,N_11896);
or U28842 (N_28842,N_16765,N_17949);
and U28843 (N_28843,N_12579,N_16755);
nor U28844 (N_28844,N_16652,N_12847);
or U28845 (N_28845,N_15656,N_13856);
nand U28846 (N_28846,N_14203,N_11358);
xnor U28847 (N_28847,N_13778,N_13922);
and U28848 (N_28848,N_13575,N_19588);
and U28849 (N_28849,N_15669,N_13266);
nor U28850 (N_28850,N_19390,N_10142);
and U28851 (N_28851,N_15259,N_10794);
nor U28852 (N_28852,N_11378,N_16434);
nand U28853 (N_28853,N_13562,N_12905);
nand U28854 (N_28854,N_11618,N_12008);
or U28855 (N_28855,N_15469,N_18618);
and U28856 (N_28856,N_19264,N_16341);
xor U28857 (N_28857,N_14442,N_12203);
nor U28858 (N_28858,N_12717,N_18740);
and U28859 (N_28859,N_19241,N_13849);
nand U28860 (N_28860,N_10787,N_18191);
nor U28861 (N_28861,N_10801,N_10221);
and U28862 (N_28862,N_11641,N_18750);
nor U28863 (N_28863,N_11736,N_14505);
or U28864 (N_28864,N_10049,N_18556);
xor U28865 (N_28865,N_17068,N_18544);
or U28866 (N_28866,N_15064,N_16626);
xnor U28867 (N_28867,N_17270,N_16433);
and U28868 (N_28868,N_10269,N_12725);
nor U28869 (N_28869,N_10708,N_18687);
and U28870 (N_28870,N_18272,N_13247);
xnor U28871 (N_28871,N_11143,N_13323);
xnor U28872 (N_28872,N_10617,N_14862);
xnor U28873 (N_28873,N_11059,N_11843);
and U28874 (N_28874,N_10814,N_10132);
nor U28875 (N_28875,N_17025,N_16814);
and U28876 (N_28876,N_18051,N_12346);
nand U28877 (N_28877,N_11952,N_13137);
xor U28878 (N_28878,N_19113,N_19231);
xor U28879 (N_28879,N_13928,N_10011);
or U28880 (N_28880,N_13667,N_11611);
or U28881 (N_28881,N_15686,N_17171);
nand U28882 (N_28882,N_16082,N_10699);
and U28883 (N_28883,N_13370,N_19990);
nand U28884 (N_28884,N_19277,N_19540);
nor U28885 (N_28885,N_11752,N_17506);
xor U28886 (N_28886,N_19662,N_12152);
xor U28887 (N_28887,N_16068,N_12295);
or U28888 (N_28888,N_12248,N_13856);
xnor U28889 (N_28889,N_13325,N_13798);
nor U28890 (N_28890,N_11242,N_11850);
xnor U28891 (N_28891,N_11752,N_14684);
or U28892 (N_28892,N_10225,N_19996);
or U28893 (N_28893,N_11419,N_17600);
and U28894 (N_28894,N_19973,N_10221);
or U28895 (N_28895,N_17957,N_13610);
or U28896 (N_28896,N_15026,N_17695);
and U28897 (N_28897,N_17279,N_11586);
xnor U28898 (N_28898,N_17023,N_10274);
nand U28899 (N_28899,N_12048,N_17449);
or U28900 (N_28900,N_11123,N_10476);
nor U28901 (N_28901,N_17105,N_11578);
or U28902 (N_28902,N_19890,N_14784);
nand U28903 (N_28903,N_18061,N_11376);
nor U28904 (N_28904,N_17010,N_19126);
xnor U28905 (N_28905,N_12547,N_15231);
nand U28906 (N_28906,N_14793,N_12638);
nor U28907 (N_28907,N_12379,N_17289);
or U28908 (N_28908,N_14527,N_15183);
nand U28909 (N_28909,N_12429,N_17556);
or U28910 (N_28910,N_12099,N_14790);
and U28911 (N_28911,N_10689,N_19694);
xnor U28912 (N_28912,N_14617,N_19468);
or U28913 (N_28913,N_11727,N_15274);
xnor U28914 (N_28914,N_11557,N_16475);
and U28915 (N_28915,N_14935,N_19614);
nor U28916 (N_28916,N_17505,N_16032);
xnor U28917 (N_28917,N_18236,N_10064);
or U28918 (N_28918,N_17379,N_11858);
nor U28919 (N_28919,N_14137,N_19330);
and U28920 (N_28920,N_11166,N_18367);
nor U28921 (N_28921,N_14421,N_13063);
xnor U28922 (N_28922,N_11368,N_16134);
nor U28923 (N_28923,N_19432,N_11241);
nand U28924 (N_28924,N_10859,N_12128);
and U28925 (N_28925,N_18055,N_15516);
nor U28926 (N_28926,N_11170,N_17211);
and U28927 (N_28927,N_14191,N_12584);
nand U28928 (N_28928,N_16577,N_18914);
or U28929 (N_28929,N_18147,N_19275);
and U28930 (N_28930,N_15507,N_19217);
nor U28931 (N_28931,N_19458,N_18812);
or U28932 (N_28932,N_15637,N_19155);
nand U28933 (N_28933,N_15546,N_11376);
and U28934 (N_28934,N_10690,N_13845);
and U28935 (N_28935,N_17429,N_16681);
nor U28936 (N_28936,N_15602,N_10363);
nor U28937 (N_28937,N_12418,N_15715);
xnor U28938 (N_28938,N_17060,N_13625);
xor U28939 (N_28939,N_14959,N_10351);
nor U28940 (N_28940,N_13128,N_13730);
nor U28941 (N_28941,N_10320,N_13376);
nand U28942 (N_28942,N_11435,N_14099);
xnor U28943 (N_28943,N_10904,N_18568);
and U28944 (N_28944,N_16586,N_10038);
nand U28945 (N_28945,N_12025,N_14700);
nand U28946 (N_28946,N_14328,N_14415);
nor U28947 (N_28947,N_17141,N_11341);
and U28948 (N_28948,N_18248,N_17903);
or U28949 (N_28949,N_14021,N_10298);
and U28950 (N_28950,N_14135,N_12168);
nand U28951 (N_28951,N_11182,N_16547);
nand U28952 (N_28952,N_13411,N_13099);
or U28953 (N_28953,N_11731,N_12509);
xor U28954 (N_28954,N_16512,N_12173);
nor U28955 (N_28955,N_10249,N_12954);
nor U28956 (N_28956,N_13841,N_10934);
nand U28957 (N_28957,N_17765,N_10502);
nor U28958 (N_28958,N_13655,N_15717);
or U28959 (N_28959,N_15688,N_16824);
or U28960 (N_28960,N_19598,N_19722);
or U28961 (N_28961,N_12764,N_18083);
nand U28962 (N_28962,N_16686,N_12080);
nand U28963 (N_28963,N_10476,N_11069);
nor U28964 (N_28964,N_11661,N_19956);
nand U28965 (N_28965,N_19627,N_12278);
nor U28966 (N_28966,N_18360,N_14751);
and U28967 (N_28967,N_11754,N_14608);
nand U28968 (N_28968,N_13387,N_13161);
nor U28969 (N_28969,N_10475,N_14309);
nand U28970 (N_28970,N_10091,N_16072);
nor U28971 (N_28971,N_18583,N_13892);
or U28972 (N_28972,N_12061,N_17776);
or U28973 (N_28973,N_19903,N_15631);
and U28974 (N_28974,N_13943,N_13248);
nand U28975 (N_28975,N_12948,N_17424);
nand U28976 (N_28976,N_16637,N_16379);
xnor U28977 (N_28977,N_12238,N_17814);
nor U28978 (N_28978,N_15483,N_12323);
xnor U28979 (N_28979,N_12656,N_14401);
nand U28980 (N_28980,N_17997,N_18482);
or U28981 (N_28981,N_16377,N_19756);
xor U28982 (N_28982,N_14278,N_11379);
xor U28983 (N_28983,N_10909,N_18904);
or U28984 (N_28984,N_12558,N_18298);
or U28985 (N_28985,N_17149,N_15281);
and U28986 (N_28986,N_10450,N_10129);
nor U28987 (N_28987,N_10757,N_13027);
and U28988 (N_28988,N_19542,N_17187);
xor U28989 (N_28989,N_15738,N_19270);
and U28990 (N_28990,N_13714,N_15238);
or U28991 (N_28991,N_12522,N_12787);
or U28992 (N_28992,N_16213,N_17496);
xnor U28993 (N_28993,N_15795,N_10760);
xnor U28994 (N_28994,N_19465,N_17568);
nand U28995 (N_28995,N_18955,N_12660);
xnor U28996 (N_28996,N_13256,N_15921);
xor U28997 (N_28997,N_19081,N_18661);
or U28998 (N_28998,N_11410,N_11008);
or U28999 (N_28999,N_15476,N_19231);
nor U29000 (N_29000,N_18289,N_10690);
nand U29001 (N_29001,N_17122,N_12162);
nand U29002 (N_29002,N_15332,N_19640);
or U29003 (N_29003,N_13737,N_16254);
and U29004 (N_29004,N_15258,N_19480);
or U29005 (N_29005,N_19844,N_12025);
xnor U29006 (N_29006,N_15220,N_12337);
or U29007 (N_29007,N_12716,N_14894);
and U29008 (N_29008,N_14441,N_19625);
xor U29009 (N_29009,N_13145,N_19504);
xor U29010 (N_29010,N_15875,N_12316);
or U29011 (N_29011,N_15442,N_13361);
nand U29012 (N_29012,N_18975,N_10968);
nor U29013 (N_29013,N_11805,N_11435);
nand U29014 (N_29014,N_19851,N_18906);
nand U29015 (N_29015,N_18989,N_18904);
xnor U29016 (N_29016,N_16217,N_14828);
nor U29017 (N_29017,N_13107,N_13827);
or U29018 (N_29018,N_14127,N_18811);
and U29019 (N_29019,N_13592,N_16974);
nor U29020 (N_29020,N_13363,N_17572);
or U29021 (N_29021,N_13984,N_15810);
nand U29022 (N_29022,N_13630,N_15363);
xor U29023 (N_29023,N_16228,N_16480);
xor U29024 (N_29024,N_10386,N_15515);
nand U29025 (N_29025,N_10930,N_10636);
and U29026 (N_29026,N_15102,N_15401);
or U29027 (N_29027,N_11356,N_10168);
nand U29028 (N_29028,N_12006,N_15169);
xnor U29029 (N_29029,N_15416,N_16537);
nand U29030 (N_29030,N_11812,N_15471);
xnor U29031 (N_29031,N_14028,N_10855);
nor U29032 (N_29032,N_19323,N_16786);
or U29033 (N_29033,N_17273,N_18558);
and U29034 (N_29034,N_19759,N_13737);
or U29035 (N_29035,N_13512,N_19032);
or U29036 (N_29036,N_11731,N_13154);
xor U29037 (N_29037,N_15724,N_17765);
nor U29038 (N_29038,N_18926,N_16057);
xnor U29039 (N_29039,N_19847,N_17207);
or U29040 (N_29040,N_13428,N_16192);
xor U29041 (N_29041,N_15861,N_14578);
or U29042 (N_29042,N_19647,N_11481);
and U29043 (N_29043,N_12280,N_14065);
nand U29044 (N_29044,N_13788,N_19019);
xor U29045 (N_29045,N_16177,N_11228);
xnor U29046 (N_29046,N_15859,N_17120);
and U29047 (N_29047,N_14803,N_19906);
xnor U29048 (N_29048,N_13105,N_17095);
and U29049 (N_29049,N_14783,N_15471);
or U29050 (N_29050,N_14306,N_19974);
nor U29051 (N_29051,N_14046,N_17101);
xnor U29052 (N_29052,N_14884,N_13892);
nor U29053 (N_29053,N_16261,N_13343);
nand U29054 (N_29054,N_16790,N_16141);
xor U29055 (N_29055,N_14096,N_17160);
nor U29056 (N_29056,N_14874,N_16309);
xnor U29057 (N_29057,N_10388,N_10883);
and U29058 (N_29058,N_15479,N_12183);
or U29059 (N_29059,N_15345,N_12951);
nor U29060 (N_29060,N_13373,N_15172);
nand U29061 (N_29061,N_17462,N_16607);
nand U29062 (N_29062,N_17986,N_15101);
or U29063 (N_29063,N_19218,N_13242);
nand U29064 (N_29064,N_18528,N_17785);
xor U29065 (N_29065,N_11987,N_16739);
and U29066 (N_29066,N_13212,N_13315);
nor U29067 (N_29067,N_13302,N_17541);
nor U29068 (N_29068,N_12099,N_12661);
and U29069 (N_29069,N_17761,N_16493);
xnor U29070 (N_29070,N_12135,N_10472);
or U29071 (N_29071,N_11165,N_19236);
and U29072 (N_29072,N_12978,N_15874);
and U29073 (N_29073,N_11112,N_17410);
nor U29074 (N_29074,N_17007,N_18341);
and U29075 (N_29075,N_10421,N_14848);
and U29076 (N_29076,N_17195,N_16969);
xnor U29077 (N_29077,N_11354,N_16896);
nand U29078 (N_29078,N_10876,N_13281);
nand U29079 (N_29079,N_18375,N_11730);
nand U29080 (N_29080,N_13635,N_17900);
and U29081 (N_29081,N_14786,N_15428);
or U29082 (N_29082,N_16331,N_15646);
xnor U29083 (N_29083,N_14623,N_14005);
or U29084 (N_29084,N_17079,N_17150);
and U29085 (N_29085,N_17187,N_19445);
xnor U29086 (N_29086,N_14908,N_11291);
nand U29087 (N_29087,N_11738,N_16569);
xnor U29088 (N_29088,N_14947,N_16123);
nand U29089 (N_29089,N_12322,N_15154);
or U29090 (N_29090,N_16084,N_11938);
xor U29091 (N_29091,N_10304,N_18938);
xnor U29092 (N_29092,N_18042,N_12651);
nor U29093 (N_29093,N_18456,N_14238);
nor U29094 (N_29094,N_11339,N_19637);
and U29095 (N_29095,N_14130,N_10487);
nor U29096 (N_29096,N_14974,N_16364);
nand U29097 (N_29097,N_19685,N_11185);
xnor U29098 (N_29098,N_10774,N_13224);
and U29099 (N_29099,N_13316,N_12779);
nand U29100 (N_29100,N_13336,N_17523);
and U29101 (N_29101,N_16699,N_13654);
nand U29102 (N_29102,N_19965,N_16345);
and U29103 (N_29103,N_19321,N_19192);
and U29104 (N_29104,N_19090,N_13487);
nor U29105 (N_29105,N_17681,N_10262);
nand U29106 (N_29106,N_14319,N_18452);
or U29107 (N_29107,N_19147,N_19721);
or U29108 (N_29108,N_19974,N_19411);
nand U29109 (N_29109,N_13974,N_12301);
and U29110 (N_29110,N_19322,N_17752);
xnor U29111 (N_29111,N_13274,N_14617);
or U29112 (N_29112,N_18025,N_19450);
and U29113 (N_29113,N_12530,N_11585);
nand U29114 (N_29114,N_13850,N_18514);
nand U29115 (N_29115,N_11203,N_11305);
nor U29116 (N_29116,N_14708,N_19121);
xor U29117 (N_29117,N_17135,N_10424);
nor U29118 (N_29118,N_19728,N_18349);
or U29119 (N_29119,N_13041,N_18462);
nor U29120 (N_29120,N_14058,N_19954);
and U29121 (N_29121,N_15291,N_12805);
nand U29122 (N_29122,N_12852,N_19322);
or U29123 (N_29123,N_10862,N_16797);
xnor U29124 (N_29124,N_11104,N_15988);
or U29125 (N_29125,N_16636,N_13762);
xor U29126 (N_29126,N_15901,N_19758);
nand U29127 (N_29127,N_18261,N_17887);
or U29128 (N_29128,N_19705,N_13416);
or U29129 (N_29129,N_13786,N_12289);
nor U29130 (N_29130,N_12382,N_11628);
nor U29131 (N_29131,N_15725,N_11991);
xor U29132 (N_29132,N_11313,N_13736);
nand U29133 (N_29133,N_11462,N_15399);
or U29134 (N_29134,N_13680,N_11390);
xnor U29135 (N_29135,N_15892,N_13837);
nand U29136 (N_29136,N_18333,N_16425);
nor U29137 (N_29137,N_19896,N_12444);
xnor U29138 (N_29138,N_10806,N_12591);
and U29139 (N_29139,N_16206,N_17288);
or U29140 (N_29140,N_15976,N_19065);
nand U29141 (N_29141,N_10832,N_17491);
nor U29142 (N_29142,N_19020,N_16009);
nor U29143 (N_29143,N_13164,N_16946);
xor U29144 (N_29144,N_11620,N_15245);
xnor U29145 (N_29145,N_12814,N_12217);
or U29146 (N_29146,N_19564,N_11198);
nand U29147 (N_29147,N_19144,N_18766);
and U29148 (N_29148,N_10874,N_17188);
nand U29149 (N_29149,N_19366,N_13307);
and U29150 (N_29150,N_13126,N_19097);
and U29151 (N_29151,N_10981,N_15474);
or U29152 (N_29152,N_19013,N_14840);
or U29153 (N_29153,N_17082,N_18076);
or U29154 (N_29154,N_17980,N_12678);
and U29155 (N_29155,N_14055,N_19829);
nand U29156 (N_29156,N_18592,N_17320);
xnor U29157 (N_29157,N_13857,N_18441);
nor U29158 (N_29158,N_19186,N_15245);
or U29159 (N_29159,N_10559,N_19821);
xnor U29160 (N_29160,N_11942,N_11673);
and U29161 (N_29161,N_16382,N_12433);
xnor U29162 (N_29162,N_12534,N_10821);
and U29163 (N_29163,N_17834,N_16009);
xnor U29164 (N_29164,N_12829,N_15567);
xnor U29165 (N_29165,N_12888,N_18542);
nor U29166 (N_29166,N_12203,N_15090);
or U29167 (N_29167,N_15292,N_12029);
nor U29168 (N_29168,N_12258,N_19061);
xnor U29169 (N_29169,N_11801,N_14107);
nor U29170 (N_29170,N_14444,N_15353);
nor U29171 (N_29171,N_11019,N_17398);
or U29172 (N_29172,N_17436,N_12519);
xnor U29173 (N_29173,N_14346,N_18739);
or U29174 (N_29174,N_15518,N_13218);
nor U29175 (N_29175,N_17153,N_10966);
or U29176 (N_29176,N_19612,N_10911);
or U29177 (N_29177,N_19454,N_16520);
nand U29178 (N_29178,N_10037,N_17531);
and U29179 (N_29179,N_13888,N_15489);
or U29180 (N_29180,N_12272,N_13789);
xor U29181 (N_29181,N_16465,N_12637);
xnor U29182 (N_29182,N_12129,N_17137);
or U29183 (N_29183,N_13511,N_19792);
nor U29184 (N_29184,N_14377,N_18557);
or U29185 (N_29185,N_10018,N_13652);
nor U29186 (N_29186,N_10530,N_10647);
nand U29187 (N_29187,N_18594,N_15644);
nor U29188 (N_29188,N_10847,N_19804);
or U29189 (N_29189,N_14189,N_12157);
or U29190 (N_29190,N_12945,N_14175);
nor U29191 (N_29191,N_13287,N_14299);
xor U29192 (N_29192,N_10696,N_15058);
or U29193 (N_29193,N_16960,N_11838);
or U29194 (N_29194,N_16790,N_16972);
or U29195 (N_29195,N_14757,N_18144);
or U29196 (N_29196,N_18274,N_10669);
or U29197 (N_29197,N_11180,N_12855);
and U29198 (N_29198,N_11730,N_12801);
and U29199 (N_29199,N_12974,N_17066);
or U29200 (N_29200,N_13815,N_15042);
xor U29201 (N_29201,N_14198,N_17858);
nand U29202 (N_29202,N_18656,N_16311);
nor U29203 (N_29203,N_17293,N_12993);
or U29204 (N_29204,N_15208,N_19825);
or U29205 (N_29205,N_13914,N_17332);
xnor U29206 (N_29206,N_10329,N_10738);
xnor U29207 (N_29207,N_19593,N_12745);
and U29208 (N_29208,N_17836,N_14480);
nor U29209 (N_29209,N_17045,N_18430);
nand U29210 (N_29210,N_19119,N_15800);
nor U29211 (N_29211,N_16616,N_17675);
or U29212 (N_29212,N_19148,N_10097);
nor U29213 (N_29213,N_10922,N_17034);
xor U29214 (N_29214,N_14300,N_14317);
nand U29215 (N_29215,N_10113,N_12280);
xor U29216 (N_29216,N_19460,N_15522);
xor U29217 (N_29217,N_18451,N_19898);
nand U29218 (N_29218,N_13246,N_12811);
and U29219 (N_29219,N_10108,N_13855);
xor U29220 (N_29220,N_14379,N_16078);
or U29221 (N_29221,N_14707,N_12345);
and U29222 (N_29222,N_18488,N_19283);
nand U29223 (N_29223,N_18470,N_11538);
or U29224 (N_29224,N_19803,N_14143);
nand U29225 (N_29225,N_19277,N_13629);
xnor U29226 (N_29226,N_10581,N_12523);
nand U29227 (N_29227,N_16065,N_14800);
and U29228 (N_29228,N_13752,N_14511);
and U29229 (N_29229,N_11330,N_13365);
xnor U29230 (N_29230,N_13044,N_12621);
or U29231 (N_29231,N_15982,N_13657);
nand U29232 (N_29232,N_15526,N_17838);
nor U29233 (N_29233,N_17132,N_17781);
and U29234 (N_29234,N_19890,N_12680);
xnor U29235 (N_29235,N_15700,N_13048);
and U29236 (N_29236,N_15640,N_19543);
nor U29237 (N_29237,N_10760,N_14137);
or U29238 (N_29238,N_16445,N_17347);
xnor U29239 (N_29239,N_18338,N_16106);
nor U29240 (N_29240,N_11130,N_14538);
and U29241 (N_29241,N_15501,N_13838);
nor U29242 (N_29242,N_15531,N_18801);
or U29243 (N_29243,N_10377,N_14464);
or U29244 (N_29244,N_12726,N_13073);
and U29245 (N_29245,N_18518,N_13446);
xnor U29246 (N_29246,N_16368,N_14733);
nor U29247 (N_29247,N_13157,N_12863);
and U29248 (N_29248,N_18550,N_11712);
or U29249 (N_29249,N_13392,N_13247);
nor U29250 (N_29250,N_16679,N_10012);
and U29251 (N_29251,N_14018,N_19870);
or U29252 (N_29252,N_14332,N_14200);
and U29253 (N_29253,N_19159,N_19308);
nand U29254 (N_29254,N_16287,N_14073);
or U29255 (N_29255,N_11410,N_11360);
xor U29256 (N_29256,N_11260,N_19498);
and U29257 (N_29257,N_10719,N_13467);
xor U29258 (N_29258,N_17122,N_13882);
nor U29259 (N_29259,N_10564,N_11026);
or U29260 (N_29260,N_16763,N_12256);
and U29261 (N_29261,N_18175,N_15912);
nor U29262 (N_29262,N_11042,N_12897);
xor U29263 (N_29263,N_17995,N_11494);
xor U29264 (N_29264,N_13482,N_18944);
and U29265 (N_29265,N_11099,N_11123);
xor U29266 (N_29266,N_18694,N_13326);
nor U29267 (N_29267,N_16719,N_16343);
or U29268 (N_29268,N_16759,N_15467);
nor U29269 (N_29269,N_13002,N_14419);
xor U29270 (N_29270,N_18811,N_16760);
xor U29271 (N_29271,N_11506,N_16378);
xnor U29272 (N_29272,N_14826,N_15792);
and U29273 (N_29273,N_17928,N_17997);
nand U29274 (N_29274,N_12802,N_10418);
and U29275 (N_29275,N_18362,N_16153);
nand U29276 (N_29276,N_12153,N_14324);
nor U29277 (N_29277,N_11390,N_11955);
or U29278 (N_29278,N_14212,N_10033);
xnor U29279 (N_29279,N_18968,N_14933);
nor U29280 (N_29280,N_19266,N_13736);
and U29281 (N_29281,N_14983,N_16222);
nor U29282 (N_29282,N_14742,N_11771);
nand U29283 (N_29283,N_12973,N_19821);
nand U29284 (N_29284,N_11980,N_14922);
xnor U29285 (N_29285,N_16031,N_11282);
or U29286 (N_29286,N_10565,N_14685);
or U29287 (N_29287,N_11592,N_10388);
nand U29288 (N_29288,N_16370,N_15736);
nand U29289 (N_29289,N_18796,N_14893);
xnor U29290 (N_29290,N_18927,N_14030);
nand U29291 (N_29291,N_15195,N_10732);
nand U29292 (N_29292,N_17427,N_18707);
nor U29293 (N_29293,N_14114,N_11628);
and U29294 (N_29294,N_13632,N_17865);
nand U29295 (N_29295,N_17025,N_17220);
and U29296 (N_29296,N_16173,N_15880);
or U29297 (N_29297,N_10148,N_14757);
nor U29298 (N_29298,N_11243,N_14884);
and U29299 (N_29299,N_16068,N_17625);
and U29300 (N_29300,N_17720,N_11081);
nand U29301 (N_29301,N_16696,N_10534);
nand U29302 (N_29302,N_13906,N_15069);
nor U29303 (N_29303,N_16961,N_16376);
and U29304 (N_29304,N_15979,N_10036);
and U29305 (N_29305,N_18075,N_15378);
and U29306 (N_29306,N_12149,N_18585);
xor U29307 (N_29307,N_13790,N_16712);
xnor U29308 (N_29308,N_15402,N_10645);
xnor U29309 (N_29309,N_14774,N_10355);
nand U29310 (N_29310,N_19377,N_17676);
nor U29311 (N_29311,N_17404,N_13574);
and U29312 (N_29312,N_18722,N_18090);
nand U29313 (N_29313,N_12315,N_15398);
xnor U29314 (N_29314,N_18185,N_13548);
xnor U29315 (N_29315,N_11310,N_15322);
xor U29316 (N_29316,N_15529,N_10361);
xnor U29317 (N_29317,N_13728,N_12940);
nor U29318 (N_29318,N_15821,N_16452);
and U29319 (N_29319,N_13542,N_19136);
nand U29320 (N_29320,N_19962,N_11355);
nand U29321 (N_29321,N_13673,N_19248);
or U29322 (N_29322,N_14070,N_16645);
nor U29323 (N_29323,N_12305,N_15621);
nand U29324 (N_29324,N_12846,N_14867);
nand U29325 (N_29325,N_14044,N_14573);
nand U29326 (N_29326,N_11440,N_12312);
and U29327 (N_29327,N_16260,N_10088);
nand U29328 (N_29328,N_19750,N_15172);
nand U29329 (N_29329,N_16599,N_11807);
nor U29330 (N_29330,N_17808,N_16256);
and U29331 (N_29331,N_16736,N_15735);
nand U29332 (N_29332,N_16172,N_15174);
or U29333 (N_29333,N_19112,N_17324);
or U29334 (N_29334,N_18573,N_12703);
and U29335 (N_29335,N_14104,N_19636);
or U29336 (N_29336,N_17073,N_14095);
or U29337 (N_29337,N_17880,N_12658);
xor U29338 (N_29338,N_18041,N_17395);
nand U29339 (N_29339,N_13313,N_19553);
nor U29340 (N_29340,N_16617,N_18086);
nand U29341 (N_29341,N_17530,N_17360);
and U29342 (N_29342,N_11113,N_11883);
nand U29343 (N_29343,N_17125,N_15939);
xor U29344 (N_29344,N_19049,N_13258);
and U29345 (N_29345,N_16965,N_19982);
or U29346 (N_29346,N_11798,N_19063);
and U29347 (N_29347,N_18553,N_11003);
xnor U29348 (N_29348,N_12279,N_13709);
nor U29349 (N_29349,N_13983,N_11809);
xor U29350 (N_29350,N_14622,N_17440);
xnor U29351 (N_29351,N_13791,N_17706);
and U29352 (N_29352,N_16456,N_15644);
nor U29353 (N_29353,N_11701,N_18947);
nor U29354 (N_29354,N_13849,N_17791);
nand U29355 (N_29355,N_17697,N_16503);
nor U29356 (N_29356,N_19449,N_15647);
and U29357 (N_29357,N_10128,N_19241);
nand U29358 (N_29358,N_16416,N_19402);
xnor U29359 (N_29359,N_14698,N_15751);
or U29360 (N_29360,N_19537,N_15221);
and U29361 (N_29361,N_10719,N_15888);
or U29362 (N_29362,N_14884,N_18415);
nand U29363 (N_29363,N_12088,N_15360);
or U29364 (N_29364,N_13868,N_12950);
nor U29365 (N_29365,N_19164,N_15088);
nand U29366 (N_29366,N_12912,N_15891);
and U29367 (N_29367,N_19420,N_17183);
or U29368 (N_29368,N_10373,N_16906);
and U29369 (N_29369,N_19323,N_16160);
xor U29370 (N_29370,N_17256,N_17230);
nand U29371 (N_29371,N_18222,N_13447);
xnor U29372 (N_29372,N_10389,N_19666);
xor U29373 (N_29373,N_17701,N_15410);
or U29374 (N_29374,N_18438,N_13624);
or U29375 (N_29375,N_19733,N_16786);
or U29376 (N_29376,N_19801,N_16407);
or U29377 (N_29377,N_16011,N_16922);
or U29378 (N_29378,N_10141,N_15774);
xnor U29379 (N_29379,N_13004,N_11892);
nand U29380 (N_29380,N_18223,N_15532);
and U29381 (N_29381,N_15363,N_11195);
or U29382 (N_29382,N_15403,N_11140);
or U29383 (N_29383,N_14676,N_17517);
nor U29384 (N_29384,N_11531,N_18280);
nand U29385 (N_29385,N_15513,N_14663);
and U29386 (N_29386,N_15325,N_12775);
or U29387 (N_29387,N_14248,N_19343);
or U29388 (N_29388,N_17922,N_13862);
or U29389 (N_29389,N_12643,N_12659);
nor U29390 (N_29390,N_14914,N_11415);
nor U29391 (N_29391,N_13061,N_12835);
nor U29392 (N_29392,N_11907,N_11469);
nor U29393 (N_29393,N_19815,N_16818);
xnor U29394 (N_29394,N_10407,N_16187);
nand U29395 (N_29395,N_13160,N_13923);
xor U29396 (N_29396,N_12659,N_11956);
nor U29397 (N_29397,N_16674,N_10826);
and U29398 (N_29398,N_17283,N_11229);
nor U29399 (N_29399,N_19706,N_15687);
xor U29400 (N_29400,N_17251,N_19866);
and U29401 (N_29401,N_12636,N_11235);
or U29402 (N_29402,N_16097,N_16997);
nor U29403 (N_29403,N_17815,N_10525);
and U29404 (N_29404,N_19595,N_10056);
or U29405 (N_29405,N_10919,N_13483);
xor U29406 (N_29406,N_14633,N_15938);
nand U29407 (N_29407,N_14053,N_13606);
nor U29408 (N_29408,N_16607,N_12502);
nor U29409 (N_29409,N_19576,N_13585);
nor U29410 (N_29410,N_18651,N_16072);
or U29411 (N_29411,N_11370,N_13839);
nand U29412 (N_29412,N_12296,N_18589);
xnor U29413 (N_29413,N_13188,N_13866);
and U29414 (N_29414,N_12454,N_15842);
xnor U29415 (N_29415,N_13818,N_17624);
and U29416 (N_29416,N_14035,N_17892);
or U29417 (N_29417,N_10702,N_15431);
or U29418 (N_29418,N_11353,N_11628);
xor U29419 (N_29419,N_13293,N_13343);
nand U29420 (N_29420,N_13316,N_15931);
xnor U29421 (N_29421,N_14133,N_16728);
xnor U29422 (N_29422,N_17070,N_17890);
nand U29423 (N_29423,N_13249,N_10315);
nand U29424 (N_29424,N_13107,N_18920);
nor U29425 (N_29425,N_16721,N_12273);
and U29426 (N_29426,N_10448,N_18381);
nand U29427 (N_29427,N_19839,N_11740);
nor U29428 (N_29428,N_10204,N_19495);
nand U29429 (N_29429,N_19123,N_13009);
xnor U29430 (N_29430,N_19403,N_13069);
or U29431 (N_29431,N_12248,N_18745);
and U29432 (N_29432,N_11899,N_15493);
nor U29433 (N_29433,N_10347,N_19491);
and U29434 (N_29434,N_18099,N_15921);
nand U29435 (N_29435,N_17483,N_12327);
and U29436 (N_29436,N_11506,N_15308);
nor U29437 (N_29437,N_14523,N_19706);
xnor U29438 (N_29438,N_13438,N_17391);
and U29439 (N_29439,N_11105,N_13421);
and U29440 (N_29440,N_16939,N_14317);
xor U29441 (N_29441,N_19804,N_15534);
xnor U29442 (N_29442,N_18120,N_12313);
or U29443 (N_29443,N_13990,N_13983);
nand U29444 (N_29444,N_13330,N_16143);
xor U29445 (N_29445,N_13049,N_11947);
or U29446 (N_29446,N_14842,N_13652);
and U29447 (N_29447,N_11359,N_15625);
and U29448 (N_29448,N_19877,N_13638);
and U29449 (N_29449,N_15294,N_18693);
and U29450 (N_29450,N_15555,N_18302);
or U29451 (N_29451,N_16822,N_15940);
and U29452 (N_29452,N_11592,N_16282);
nor U29453 (N_29453,N_11030,N_11974);
and U29454 (N_29454,N_13959,N_10196);
and U29455 (N_29455,N_15956,N_18435);
nand U29456 (N_29456,N_10455,N_10645);
nor U29457 (N_29457,N_14975,N_10061);
or U29458 (N_29458,N_14773,N_13184);
or U29459 (N_29459,N_19270,N_13101);
nor U29460 (N_29460,N_10703,N_13019);
or U29461 (N_29461,N_17092,N_19410);
and U29462 (N_29462,N_16641,N_12703);
xor U29463 (N_29463,N_19903,N_14822);
nor U29464 (N_29464,N_14199,N_15247);
or U29465 (N_29465,N_14872,N_16125);
and U29466 (N_29466,N_13347,N_13195);
xnor U29467 (N_29467,N_15987,N_19507);
or U29468 (N_29468,N_11963,N_18896);
nand U29469 (N_29469,N_10737,N_14064);
or U29470 (N_29470,N_15145,N_16218);
xnor U29471 (N_29471,N_16419,N_10957);
nand U29472 (N_29472,N_13651,N_12027);
nand U29473 (N_29473,N_12102,N_11378);
xnor U29474 (N_29474,N_18795,N_18335);
or U29475 (N_29475,N_12347,N_18357);
nand U29476 (N_29476,N_12436,N_16134);
xor U29477 (N_29477,N_11776,N_19132);
and U29478 (N_29478,N_15657,N_14744);
nor U29479 (N_29479,N_14289,N_18837);
nand U29480 (N_29480,N_12667,N_12718);
and U29481 (N_29481,N_16489,N_11530);
nor U29482 (N_29482,N_16356,N_18501);
or U29483 (N_29483,N_12136,N_14828);
nor U29484 (N_29484,N_15674,N_14813);
nor U29485 (N_29485,N_18280,N_11848);
nand U29486 (N_29486,N_18832,N_12732);
nand U29487 (N_29487,N_15130,N_16495);
xor U29488 (N_29488,N_13304,N_18995);
or U29489 (N_29489,N_12045,N_18486);
nand U29490 (N_29490,N_14001,N_12469);
nor U29491 (N_29491,N_15343,N_16441);
or U29492 (N_29492,N_11877,N_16958);
nand U29493 (N_29493,N_10032,N_17660);
nand U29494 (N_29494,N_13150,N_17063);
and U29495 (N_29495,N_14987,N_16623);
nor U29496 (N_29496,N_13281,N_19253);
or U29497 (N_29497,N_15101,N_14686);
or U29498 (N_29498,N_11222,N_11556);
xnor U29499 (N_29499,N_15980,N_16959);
nand U29500 (N_29500,N_10646,N_19167);
xor U29501 (N_29501,N_18772,N_13605);
xnor U29502 (N_29502,N_17422,N_16925);
nand U29503 (N_29503,N_15747,N_17725);
and U29504 (N_29504,N_14972,N_18536);
nand U29505 (N_29505,N_15358,N_11905);
and U29506 (N_29506,N_17640,N_11076);
nor U29507 (N_29507,N_14128,N_13589);
xor U29508 (N_29508,N_16335,N_14523);
and U29509 (N_29509,N_15940,N_10307);
or U29510 (N_29510,N_14332,N_15594);
xor U29511 (N_29511,N_17446,N_19438);
or U29512 (N_29512,N_11431,N_17030);
and U29513 (N_29513,N_13603,N_12782);
and U29514 (N_29514,N_11331,N_16114);
nor U29515 (N_29515,N_19370,N_10826);
and U29516 (N_29516,N_12649,N_15386);
nor U29517 (N_29517,N_17162,N_17765);
and U29518 (N_29518,N_16379,N_12099);
xor U29519 (N_29519,N_14789,N_16480);
nor U29520 (N_29520,N_17835,N_12970);
or U29521 (N_29521,N_19580,N_17918);
and U29522 (N_29522,N_13611,N_11184);
nor U29523 (N_29523,N_10539,N_11897);
and U29524 (N_29524,N_12701,N_12000);
nor U29525 (N_29525,N_14427,N_19183);
and U29526 (N_29526,N_17169,N_18988);
and U29527 (N_29527,N_18024,N_16430);
xnor U29528 (N_29528,N_14381,N_16780);
and U29529 (N_29529,N_13950,N_14798);
xor U29530 (N_29530,N_11782,N_12619);
nor U29531 (N_29531,N_14324,N_11027);
and U29532 (N_29532,N_15839,N_17165);
nand U29533 (N_29533,N_14010,N_17746);
and U29534 (N_29534,N_17830,N_14482);
xor U29535 (N_29535,N_16503,N_12757);
xor U29536 (N_29536,N_15272,N_16653);
xnor U29537 (N_29537,N_14119,N_19525);
and U29538 (N_29538,N_12822,N_16880);
nand U29539 (N_29539,N_15629,N_19269);
and U29540 (N_29540,N_17988,N_18459);
or U29541 (N_29541,N_17262,N_16153);
nor U29542 (N_29542,N_12757,N_15132);
or U29543 (N_29543,N_17078,N_12039);
nand U29544 (N_29544,N_16353,N_10180);
and U29545 (N_29545,N_11642,N_15243);
nor U29546 (N_29546,N_18557,N_11568);
and U29547 (N_29547,N_10319,N_18203);
or U29548 (N_29548,N_16489,N_12075);
or U29549 (N_29549,N_12650,N_18262);
and U29550 (N_29550,N_10047,N_15079);
or U29551 (N_29551,N_14450,N_17217);
xor U29552 (N_29552,N_16371,N_11420);
nand U29553 (N_29553,N_10578,N_10123);
and U29554 (N_29554,N_11003,N_13792);
nor U29555 (N_29555,N_16654,N_16206);
xnor U29556 (N_29556,N_16600,N_13867);
and U29557 (N_29557,N_11971,N_15963);
xnor U29558 (N_29558,N_13219,N_13585);
xor U29559 (N_29559,N_17557,N_15521);
nor U29560 (N_29560,N_12421,N_18523);
nor U29561 (N_29561,N_13873,N_11021);
or U29562 (N_29562,N_13226,N_12503);
or U29563 (N_29563,N_14861,N_12207);
and U29564 (N_29564,N_15755,N_18164);
and U29565 (N_29565,N_13589,N_11402);
or U29566 (N_29566,N_12091,N_18843);
nand U29567 (N_29567,N_14570,N_15516);
nor U29568 (N_29568,N_18896,N_11855);
and U29569 (N_29569,N_10733,N_16359);
and U29570 (N_29570,N_11724,N_10418);
nand U29571 (N_29571,N_16878,N_12321);
nor U29572 (N_29572,N_16030,N_14783);
nand U29573 (N_29573,N_11562,N_13350);
or U29574 (N_29574,N_18772,N_15538);
nand U29575 (N_29575,N_11183,N_11961);
or U29576 (N_29576,N_15012,N_13507);
nor U29577 (N_29577,N_16628,N_19933);
nor U29578 (N_29578,N_11147,N_12553);
nand U29579 (N_29579,N_18003,N_18257);
nand U29580 (N_29580,N_13194,N_14936);
nand U29581 (N_29581,N_14224,N_14340);
or U29582 (N_29582,N_19378,N_11549);
xnor U29583 (N_29583,N_14463,N_15618);
or U29584 (N_29584,N_17895,N_16037);
nand U29585 (N_29585,N_12572,N_11087);
nand U29586 (N_29586,N_12745,N_19525);
and U29587 (N_29587,N_18035,N_10732);
or U29588 (N_29588,N_18368,N_18076);
or U29589 (N_29589,N_10394,N_11198);
xnor U29590 (N_29590,N_10814,N_13614);
nand U29591 (N_29591,N_12888,N_12145);
and U29592 (N_29592,N_10015,N_19739);
or U29593 (N_29593,N_11983,N_12093);
or U29594 (N_29594,N_15021,N_11866);
nand U29595 (N_29595,N_10603,N_14340);
nand U29596 (N_29596,N_19949,N_19132);
or U29597 (N_29597,N_18850,N_17018);
nand U29598 (N_29598,N_19088,N_18213);
or U29599 (N_29599,N_18538,N_18070);
and U29600 (N_29600,N_17988,N_15069);
nand U29601 (N_29601,N_17462,N_18854);
and U29602 (N_29602,N_10213,N_17922);
xnor U29603 (N_29603,N_10388,N_15633);
or U29604 (N_29604,N_14735,N_18199);
nand U29605 (N_29605,N_13280,N_11935);
or U29606 (N_29606,N_12696,N_13558);
nand U29607 (N_29607,N_16854,N_18786);
and U29608 (N_29608,N_10415,N_15903);
and U29609 (N_29609,N_16412,N_18040);
or U29610 (N_29610,N_16422,N_15100);
nor U29611 (N_29611,N_17199,N_14791);
or U29612 (N_29612,N_18516,N_12965);
and U29613 (N_29613,N_13194,N_18296);
and U29614 (N_29614,N_11169,N_13164);
xor U29615 (N_29615,N_12746,N_15431);
nor U29616 (N_29616,N_14089,N_16919);
nand U29617 (N_29617,N_19880,N_13524);
xnor U29618 (N_29618,N_13687,N_16525);
and U29619 (N_29619,N_13496,N_10185);
nor U29620 (N_29620,N_19257,N_12367);
and U29621 (N_29621,N_18987,N_15437);
nand U29622 (N_29622,N_19159,N_17482);
or U29623 (N_29623,N_14058,N_19506);
and U29624 (N_29624,N_13165,N_11275);
and U29625 (N_29625,N_18783,N_12196);
and U29626 (N_29626,N_19699,N_19340);
nor U29627 (N_29627,N_11793,N_15257);
xnor U29628 (N_29628,N_12959,N_13726);
nor U29629 (N_29629,N_10010,N_15362);
or U29630 (N_29630,N_17106,N_15818);
and U29631 (N_29631,N_10563,N_19886);
or U29632 (N_29632,N_10128,N_15951);
or U29633 (N_29633,N_12256,N_13081);
or U29634 (N_29634,N_14654,N_10305);
nor U29635 (N_29635,N_10506,N_17623);
nor U29636 (N_29636,N_13567,N_16958);
nand U29637 (N_29637,N_17497,N_19393);
or U29638 (N_29638,N_14555,N_10361);
nand U29639 (N_29639,N_18926,N_10024);
or U29640 (N_29640,N_16094,N_14342);
nand U29641 (N_29641,N_14716,N_15064);
and U29642 (N_29642,N_11032,N_15278);
or U29643 (N_29643,N_10108,N_14351);
and U29644 (N_29644,N_12819,N_15828);
or U29645 (N_29645,N_18125,N_13467);
xor U29646 (N_29646,N_19310,N_10310);
xnor U29647 (N_29647,N_11448,N_11360);
nor U29648 (N_29648,N_12104,N_10227);
xnor U29649 (N_29649,N_19126,N_15683);
or U29650 (N_29650,N_18526,N_17700);
nor U29651 (N_29651,N_16504,N_10285);
and U29652 (N_29652,N_15200,N_12771);
nor U29653 (N_29653,N_10782,N_18036);
nand U29654 (N_29654,N_14534,N_13016);
and U29655 (N_29655,N_18261,N_12453);
xor U29656 (N_29656,N_15016,N_14048);
nor U29657 (N_29657,N_13441,N_10522);
or U29658 (N_29658,N_11386,N_10322);
or U29659 (N_29659,N_12818,N_12205);
xnor U29660 (N_29660,N_14062,N_16485);
xnor U29661 (N_29661,N_13300,N_14220);
and U29662 (N_29662,N_12824,N_11397);
xor U29663 (N_29663,N_16496,N_10593);
nand U29664 (N_29664,N_14721,N_15912);
nor U29665 (N_29665,N_17191,N_11950);
and U29666 (N_29666,N_18182,N_15565);
and U29667 (N_29667,N_16011,N_11560);
or U29668 (N_29668,N_16842,N_11393);
xnor U29669 (N_29669,N_18947,N_16164);
nand U29670 (N_29670,N_16026,N_12392);
or U29671 (N_29671,N_14667,N_19166);
and U29672 (N_29672,N_10411,N_17379);
and U29673 (N_29673,N_12057,N_16345);
and U29674 (N_29674,N_17642,N_16679);
xor U29675 (N_29675,N_14943,N_13016);
xor U29676 (N_29676,N_14742,N_11252);
or U29677 (N_29677,N_17034,N_19027);
and U29678 (N_29678,N_10723,N_11265);
nor U29679 (N_29679,N_18232,N_13050);
or U29680 (N_29680,N_13531,N_12700);
and U29681 (N_29681,N_17839,N_15593);
and U29682 (N_29682,N_17251,N_17760);
or U29683 (N_29683,N_10157,N_17104);
nand U29684 (N_29684,N_14083,N_17587);
nand U29685 (N_29685,N_11164,N_18410);
nor U29686 (N_29686,N_10092,N_10143);
nor U29687 (N_29687,N_14971,N_18942);
or U29688 (N_29688,N_17662,N_12704);
nand U29689 (N_29689,N_18928,N_15579);
or U29690 (N_29690,N_17887,N_10535);
xor U29691 (N_29691,N_11499,N_19831);
nor U29692 (N_29692,N_15485,N_12326);
xor U29693 (N_29693,N_18356,N_16170);
xnor U29694 (N_29694,N_13284,N_16112);
and U29695 (N_29695,N_11056,N_17740);
and U29696 (N_29696,N_16916,N_14605);
or U29697 (N_29697,N_19617,N_12032);
nor U29698 (N_29698,N_18550,N_17131);
nor U29699 (N_29699,N_18949,N_19120);
xor U29700 (N_29700,N_18563,N_16087);
nor U29701 (N_29701,N_10372,N_13617);
or U29702 (N_29702,N_19643,N_16509);
nand U29703 (N_29703,N_12756,N_19158);
or U29704 (N_29704,N_15427,N_13600);
nand U29705 (N_29705,N_19756,N_12551);
and U29706 (N_29706,N_12075,N_15358);
xnor U29707 (N_29707,N_19803,N_19319);
or U29708 (N_29708,N_17855,N_10687);
nor U29709 (N_29709,N_17463,N_11749);
xnor U29710 (N_29710,N_17950,N_16485);
and U29711 (N_29711,N_14787,N_15951);
and U29712 (N_29712,N_17143,N_16156);
nand U29713 (N_29713,N_13859,N_16931);
nor U29714 (N_29714,N_18910,N_17630);
nor U29715 (N_29715,N_18337,N_19270);
and U29716 (N_29716,N_19902,N_18569);
nor U29717 (N_29717,N_16626,N_16612);
xor U29718 (N_29718,N_18310,N_15850);
and U29719 (N_29719,N_14725,N_18796);
or U29720 (N_29720,N_11052,N_14456);
or U29721 (N_29721,N_10492,N_10744);
nand U29722 (N_29722,N_13506,N_10470);
and U29723 (N_29723,N_14637,N_17670);
xor U29724 (N_29724,N_17619,N_18467);
xnor U29725 (N_29725,N_15961,N_15279);
or U29726 (N_29726,N_13517,N_12481);
nand U29727 (N_29727,N_16973,N_10091);
xor U29728 (N_29728,N_10705,N_17788);
nor U29729 (N_29729,N_15328,N_11075);
nand U29730 (N_29730,N_12457,N_11058);
or U29731 (N_29731,N_11554,N_13615);
xor U29732 (N_29732,N_12163,N_14513);
nand U29733 (N_29733,N_13867,N_12238);
and U29734 (N_29734,N_19115,N_15441);
and U29735 (N_29735,N_11782,N_11538);
or U29736 (N_29736,N_11877,N_14889);
nor U29737 (N_29737,N_15588,N_11565);
nand U29738 (N_29738,N_19645,N_12416);
and U29739 (N_29739,N_17872,N_16041);
or U29740 (N_29740,N_17844,N_14425);
and U29741 (N_29741,N_16893,N_12134);
xnor U29742 (N_29742,N_16458,N_11453);
nor U29743 (N_29743,N_12621,N_16297);
nor U29744 (N_29744,N_18372,N_19254);
nor U29745 (N_29745,N_16181,N_11101);
xor U29746 (N_29746,N_12798,N_11491);
nor U29747 (N_29747,N_19780,N_19621);
and U29748 (N_29748,N_17508,N_16768);
xor U29749 (N_29749,N_18339,N_15168);
nor U29750 (N_29750,N_16462,N_14901);
nand U29751 (N_29751,N_11991,N_15373);
nor U29752 (N_29752,N_11105,N_17442);
and U29753 (N_29753,N_17551,N_14481);
and U29754 (N_29754,N_10246,N_16235);
nor U29755 (N_29755,N_14619,N_10263);
nor U29756 (N_29756,N_15058,N_16308);
xnor U29757 (N_29757,N_16969,N_14503);
or U29758 (N_29758,N_13458,N_13792);
xor U29759 (N_29759,N_16198,N_19656);
or U29760 (N_29760,N_14323,N_12242);
nand U29761 (N_29761,N_14351,N_16968);
nand U29762 (N_29762,N_14693,N_14144);
nor U29763 (N_29763,N_19568,N_17366);
or U29764 (N_29764,N_19942,N_19782);
nor U29765 (N_29765,N_19772,N_17045);
nand U29766 (N_29766,N_10632,N_19691);
or U29767 (N_29767,N_16765,N_14810);
nand U29768 (N_29768,N_14104,N_19989);
xor U29769 (N_29769,N_18656,N_13081);
nor U29770 (N_29770,N_14038,N_16879);
nor U29771 (N_29771,N_16744,N_10790);
or U29772 (N_29772,N_12518,N_18572);
nand U29773 (N_29773,N_14996,N_17870);
or U29774 (N_29774,N_19188,N_15148);
or U29775 (N_29775,N_18626,N_15273);
xnor U29776 (N_29776,N_10994,N_16409);
xor U29777 (N_29777,N_15190,N_18690);
xnor U29778 (N_29778,N_18397,N_18538);
xnor U29779 (N_29779,N_15277,N_17077);
nor U29780 (N_29780,N_13772,N_17315);
and U29781 (N_29781,N_18820,N_19792);
or U29782 (N_29782,N_10385,N_16802);
nand U29783 (N_29783,N_10101,N_11105);
nand U29784 (N_29784,N_14293,N_12986);
or U29785 (N_29785,N_12510,N_10649);
nand U29786 (N_29786,N_12644,N_12818);
nand U29787 (N_29787,N_12208,N_11463);
and U29788 (N_29788,N_10978,N_17279);
or U29789 (N_29789,N_14108,N_12030);
nor U29790 (N_29790,N_10195,N_17196);
and U29791 (N_29791,N_16333,N_12430);
xnor U29792 (N_29792,N_10767,N_13529);
and U29793 (N_29793,N_13629,N_12773);
nand U29794 (N_29794,N_18001,N_18422);
xor U29795 (N_29795,N_12295,N_13725);
nand U29796 (N_29796,N_11715,N_13408);
or U29797 (N_29797,N_15029,N_15753);
nand U29798 (N_29798,N_14283,N_16936);
xor U29799 (N_29799,N_19562,N_13762);
xnor U29800 (N_29800,N_14689,N_15182);
nor U29801 (N_29801,N_12661,N_14806);
and U29802 (N_29802,N_10080,N_15739);
or U29803 (N_29803,N_17472,N_18257);
xnor U29804 (N_29804,N_14724,N_12794);
xnor U29805 (N_29805,N_15445,N_12170);
xnor U29806 (N_29806,N_15605,N_10412);
xor U29807 (N_29807,N_19908,N_16646);
nor U29808 (N_29808,N_16069,N_13488);
nand U29809 (N_29809,N_12236,N_16529);
or U29810 (N_29810,N_12512,N_18152);
nor U29811 (N_29811,N_16303,N_12223);
or U29812 (N_29812,N_11744,N_14365);
nand U29813 (N_29813,N_13538,N_16488);
nor U29814 (N_29814,N_18615,N_15232);
nor U29815 (N_29815,N_17220,N_16458);
nand U29816 (N_29816,N_14538,N_10131);
and U29817 (N_29817,N_12408,N_18179);
nor U29818 (N_29818,N_19170,N_13567);
or U29819 (N_29819,N_18641,N_19535);
nor U29820 (N_29820,N_13681,N_18563);
and U29821 (N_29821,N_13844,N_10648);
xnor U29822 (N_29822,N_17847,N_19834);
xnor U29823 (N_29823,N_16718,N_15904);
nor U29824 (N_29824,N_16778,N_19221);
and U29825 (N_29825,N_19630,N_12653);
or U29826 (N_29826,N_10564,N_14633);
nor U29827 (N_29827,N_17378,N_16826);
xnor U29828 (N_29828,N_12267,N_16855);
or U29829 (N_29829,N_16140,N_15969);
and U29830 (N_29830,N_11032,N_19492);
or U29831 (N_29831,N_15754,N_12759);
and U29832 (N_29832,N_16886,N_11718);
xnor U29833 (N_29833,N_18201,N_15946);
or U29834 (N_29834,N_13788,N_19157);
nand U29835 (N_29835,N_13913,N_19918);
nand U29836 (N_29836,N_14148,N_15299);
nor U29837 (N_29837,N_11790,N_19334);
or U29838 (N_29838,N_13755,N_17236);
xor U29839 (N_29839,N_16630,N_14665);
or U29840 (N_29840,N_13117,N_11286);
nor U29841 (N_29841,N_18124,N_18396);
or U29842 (N_29842,N_15078,N_16924);
and U29843 (N_29843,N_16656,N_17756);
or U29844 (N_29844,N_17452,N_17331);
or U29845 (N_29845,N_16217,N_10880);
nor U29846 (N_29846,N_15786,N_13230);
nand U29847 (N_29847,N_14142,N_17100);
nand U29848 (N_29848,N_13843,N_13266);
nand U29849 (N_29849,N_10943,N_18785);
nand U29850 (N_29850,N_15816,N_13733);
nand U29851 (N_29851,N_19525,N_19769);
and U29852 (N_29852,N_11266,N_17211);
nor U29853 (N_29853,N_10766,N_18401);
nand U29854 (N_29854,N_12544,N_11126);
or U29855 (N_29855,N_10534,N_16266);
nor U29856 (N_29856,N_19450,N_10269);
and U29857 (N_29857,N_15622,N_10024);
or U29858 (N_29858,N_14405,N_12940);
xor U29859 (N_29859,N_16358,N_18024);
xnor U29860 (N_29860,N_17680,N_16757);
xor U29861 (N_29861,N_12121,N_19052);
and U29862 (N_29862,N_13406,N_17681);
or U29863 (N_29863,N_13167,N_15015);
and U29864 (N_29864,N_13905,N_10120);
xor U29865 (N_29865,N_11167,N_16225);
nor U29866 (N_29866,N_10850,N_16456);
nand U29867 (N_29867,N_10947,N_11081);
nor U29868 (N_29868,N_13500,N_14655);
xnor U29869 (N_29869,N_12267,N_19627);
and U29870 (N_29870,N_16994,N_17283);
xor U29871 (N_29871,N_14631,N_19566);
nand U29872 (N_29872,N_14244,N_17967);
nor U29873 (N_29873,N_19946,N_17685);
nand U29874 (N_29874,N_17915,N_14596);
nor U29875 (N_29875,N_11816,N_11341);
nor U29876 (N_29876,N_15970,N_11473);
xor U29877 (N_29877,N_15209,N_19701);
nand U29878 (N_29878,N_12344,N_17500);
xor U29879 (N_29879,N_18491,N_18591);
nor U29880 (N_29880,N_17976,N_12274);
nor U29881 (N_29881,N_12739,N_12309);
or U29882 (N_29882,N_11457,N_14908);
nor U29883 (N_29883,N_12143,N_13428);
xnor U29884 (N_29884,N_11664,N_18689);
or U29885 (N_29885,N_15988,N_12997);
or U29886 (N_29886,N_17802,N_14345);
nand U29887 (N_29887,N_14589,N_14990);
nor U29888 (N_29888,N_13659,N_17471);
xnor U29889 (N_29889,N_18731,N_10453);
xnor U29890 (N_29890,N_12468,N_14135);
xnor U29891 (N_29891,N_14058,N_19698);
nand U29892 (N_29892,N_17084,N_14059);
or U29893 (N_29893,N_12612,N_16141);
nand U29894 (N_29894,N_12888,N_18053);
xor U29895 (N_29895,N_12528,N_14557);
nand U29896 (N_29896,N_12049,N_13783);
or U29897 (N_29897,N_19707,N_16710);
or U29898 (N_29898,N_10184,N_17880);
nor U29899 (N_29899,N_16853,N_12368);
nand U29900 (N_29900,N_15902,N_12030);
or U29901 (N_29901,N_18491,N_15988);
nor U29902 (N_29902,N_12830,N_14593);
xor U29903 (N_29903,N_12052,N_18877);
and U29904 (N_29904,N_18947,N_19007);
nor U29905 (N_29905,N_16724,N_17651);
nor U29906 (N_29906,N_10815,N_17602);
or U29907 (N_29907,N_17369,N_17728);
and U29908 (N_29908,N_14158,N_12219);
nand U29909 (N_29909,N_13114,N_13572);
and U29910 (N_29910,N_15350,N_10393);
or U29911 (N_29911,N_11713,N_17099);
and U29912 (N_29912,N_18561,N_18177);
or U29913 (N_29913,N_17138,N_18589);
or U29914 (N_29914,N_16072,N_17997);
nor U29915 (N_29915,N_17905,N_19560);
or U29916 (N_29916,N_10486,N_13333);
and U29917 (N_29917,N_10916,N_13782);
and U29918 (N_29918,N_15075,N_11243);
nand U29919 (N_29919,N_10825,N_10201);
nand U29920 (N_29920,N_13188,N_18222);
xor U29921 (N_29921,N_10779,N_15216);
xor U29922 (N_29922,N_16501,N_15738);
nor U29923 (N_29923,N_13928,N_12107);
nor U29924 (N_29924,N_19713,N_13618);
nand U29925 (N_29925,N_18678,N_15829);
xnor U29926 (N_29926,N_15354,N_16437);
nand U29927 (N_29927,N_11783,N_13094);
or U29928 (N_29928,N_10001,N_17532);
and U29929 (N_29929,N_19587,N_12402);
nor U29930 (N_29930,N_12298,N_13663);
nand U29931 (N_29931,N_11335,N_15011);
xor U29932 (N_29932,N_19549,N_13967);
nand U29933 (N_29933,N_19689,N_15339);
xnor U29934 (N_29934,N_10873,N_19387);
or U29935 (N_29935,N_13965,N_19923);
xor U29936 (N_29936,N_13984,N_18405);
and U29937 (N_29937,N_10160,N_10807);
nor U29938 (N_29938,N_11413,N_18767);
nand U29939 (N_29939,N_12516,N_18771);
nand U29940 (N_29940,N_17399,N_15228);
or U29941 (N_29941,N_16563,N_16914);
and U29942 (N_29942,N_19767,N_10453);
xnor U29943 (N_29943,N_12319,N_15947);
or U29944 (N_29944,N_10869,N_12389);
and U29945 (N_29945,N_17440,N_19628);
or U29946 (N_29946,N_16332,N_17824);
xnor U29947 (N_29947,N_19643,N_11226);
nor U29948 (N_29948,N_19761,N_19287);
nor U29949 (N_29949,N_12328,N_12581);
xnor U29950 (N_29950,N_12381,N_11965);
and U29951 (N_29951,N_11166,N_18208);
xnor U29952 (N_29952,N_14328,N_16895);
nand U29953 (N_29953,N_18341,N_10665);
and U29954 (N_29954,N_12887,N_16780);
xor U29955 (N_29955,N_10688,N_11088);
or U29956 (N_29956,N_14079,N_10633);
nor U29957 (N_29957,N_14893,N_16213);
nor U29958 (N_29958,N_11572,N_19242);
nor U29959 (N_29959,N_12772,N_17230);
xor U29960 (N_29960,N_14578,N_17816);
xor U29961 (N_29961,N_17130,N_13139);
nor U29962 (N_29962,N_15972,N_12036);
or U29963 (N_29963,N_12656,N_18902);
and U29964 (N_29964,N_18631,N_10513);
nor U29965 (N_29965,N_17125,N_15136);
or U29966 (N_29966,N_14502,N_17438);
nand U29967 (N_29967,N_19261,N_19358);
nor U29968 (N_29968,N_10322,N_17078);
nor U29969 (N_29969,N_18789,N_10205);
nand U29970 (N_29970,N_12037,N_18082);
xnor U29971 (N_29971,N_17641,N_16113);
nor U29972 (N_29972,N_13630,N_11078);
and U29973 (N_29973,N_16609,N_17659);
xnor U29974 (N_29974,N_17762,N_11596);
xor U29975 (N_29975,N_11617,N_15984);
and U29976 (N_29976,N_14381,N_10424);
xor U29977 (N_29977,N_19991,N_12496);
or U29978 (N_29978,N_16050,N_18963);
nor U29979 (N_29979,N_10989,N_11399);
nor U29980 (N_29980,N_12267,N_13307);
nor U29981 (N_29981,N_17556,N_10364);
and U29982 (N_29982,N_18044,N_16460);
nand U29983 (N_29983,N_16461,N_10560);
nand U29984 (N_29984,N_19574,N_17319);
or U29985 (N_29985,N_12989,N_19437);
xnor U29986 (N_29986,N_16258,N_13896);
and U29987 (N_29987,N_17069,N_17352);
and U29988 (N_29988,N_16104,N_18302);
xor U29989 (N_29989,N_19034,N_11436);
and U29990 (N_29990,N_15063,N_12537);
xor U29991 (N_29991,N_16441,N_17552);
and U29992 (N_29992,N_11958,N_15543);
or U29993 (N_29993,N_14984,N_16633);
or U29994 (N_29994,N_13592,N_11979);
nor U29995 (N_29995,N_14053,N_19987);
nor U29996 (N_29996,N_12197,N_13489);
xor U29997 (N_29997,N_17680,N_18937);
xnor U29998 (N_29998,N_18994,N_13247);
xor U29999 (N_29999,N_12147,N_13908);
and UO_0 (O_0,N_29312,N_20225);
xnor UO_1 (O_1,N_23298,N_27885);
and UO_2 (O_2,N_28090,N_20129);
nand UO_3 (O_3,N_23486,N_25701);
or UO_4 (O_4,N_29581,N_22255);
and UO_5 (O_5,N_22416,N_28852);
and UO_6 (O_6,N_23022,N_22237);
and UO_7 (O_7,N_20700,N_20396);
xor UO_8 (O_8,N_26641,N_21068);
or UO_9 (O_9,N_27682,N_22883);
nor UO_10 (O_10,N_23907,N_22011);
xor UO_11 (O_11,N_28969,N_27952);
and UO_12 (O_12,N_27382,N_28935);
xnor UO_13 (O_13,N_27645,N_27573);
and UO_14 (O_14,N_22104,N_24061);
or UO_15 (O_15,N_22711,N_21005);
nor UO_16 (O_16,N_21976,N_25627);
and UO_17 (O_17,N_28584,N_26707);
nor UO_18 (O_18,N_23375,N_28717);
and UO_19 (O_19,N_25224,N_25575);
or UO_20 (O_20,N_23152,N_28418);
xnor UO_21 (O_21,N_21850,N_22658);
xor UO_22 (O_22,N_22777,N_23004);
or UO_23 (O_23,N_25038,N_28232);
nand UO_24 (O_24,N_21905,N_23985);
and UO_25 (O_25,N_26511,N_28641);
nor UO_26 (O_26,N_29493,N_29571);
and UO_27 (O_27,N_28086,N_25415);
or UO_28 (O_28,N_29250,N_22103);
or UO_29 (O_29,N_21172,N_25337);
nand UO_30 (O_30,N_28849,N_28588);
and UO_31 (O_31,N_28972,N_23822);
nor UO_32 (O_32,N_24533,N_20207);
and UO_33 (O_33,N_21477,N_23772);
nor UO_34 (O_34,N_28026,N_26014);
or UO_35 (O_35,N_22623,N_29427);
and UO_36 (O_36,N_20272,N_25120);
nand UO_37 (O_37,N_26938,N_20021);
xor UO_38 (O_38,N_22153,N_21938);
nand UO_39 (O_39,N_21699,N_23497);
nor UO_40 (O_40,N_28455,N_26686);
nand UO_41 (O_41,N_29221,N_20805);
or UO_42 (O_42,N_29759,N_22119);
nor UO_43 (O_43,N_27889,N_25113);
nor UO_44 (O_44,N_20955,N_27252);
nand UO_45 (O_45,N_22782,N_20151);
nor UO_46 (O_46,N_22144,N_24855);
nor UO_47 (O_47,N_25072,N_27405);
nand UO_48 (O_48,N_21369,N_20008);
nor UO_49 (O_49,N_23823,N_29095);
xnor UO_50 (O_50,N_20914,N_20310);
and UO_51 (O_51,N_24249,N_25323);
nor UO_52 (O_52,N_24543,N_20152);
or UO_53 (O_53,N_21420,N_27718);
xor UO_54 (O_54,N_20439,N_24148);
or UO_55 (O_55,N_24549,N_25200);
and UO_56 (O_56,N_28134,N_21982);
or UO_57 (O_57,N_20414,N_29796);
or UO_58 (O_58,N_23141,N_20244);
xor UO_59 (O_59,N_20067,N_21050);
nand UO_60 (O_60,N_24833,N_21849);
xor UO_61 (O_61,N_29174,N_25125);
nor UO_62 (O_62,N_24540,N_21985);
xnor UO_63 (O_63,N_26138,N_29382);
xnor UO_64 (O_64,N_27568,N_27759);
or UO_65 (O_65,N_27843,N_28457);
xor UO_66 (O_66,N_25062,N_21291);
and UO_67 (O_67,N_27555,N_21088);
or UO_68 (O_68,N_24985,N_20673);
xor UO_69 (O_69,N_24534,N_21160);
or UO_70 (O_70,N_26103,N_29670);
nor UO_71 (O_71,N_21688,N_25880);
nor UO_72 (O_72,N_27280,N_27501);
xnor UO_73 (O_73,N_28348,N_28580);
and UO_74 (O_74,N_25871,N_29959);
or UO_75 (O_75,N_20444,N_27419);
nand UO_76 (O_76,N_20234,N_22302);
and UO_77 (O_77,N_22474,N_21353);
nor UO_78 (O_78,N_24299,N_22213);
xnor UO_79 (O_79,N_28900,N_28998);
xor UO_80 (O_80,N_24021,N_28072);
xnor UO_81 (O_81,N_24486,N_20556);
xor UO_82 (O_82,N_26474,N_28763);
xnor UO_83 (O_83,N_21865,N_23150);
nand UO_84 (O_84,N_24680,N_26912);
or UO_85 (O_85,N_24296,N_26637);
or UO_86 (O_86,N_23793,N_28014);
nand UO_87 (O_87,N_29369,N_22385);
xnor UO_88 (O_88,N_28645,N_27196);
or UO_89 (O_89,N_20395,N_24467);
and UO_90 (O_90,N_24685,N_26328);
or UO_91 (O_91,N_29912,N_24491);
nand UO_92 (O_92,N_25819,N_20066);
xor UO_93 (O_93,N_25074,N_20848);
or UO_94 (O_94,N_28111,N_27527);
or UO_95 (O_95,N_25037,N_20488);
nand UO_96 (O_96,N_22996,N_25287);
nor UO_97 (O_97,N_29529,N_27213);
xnor UO_98 (O_98,N_20859,N_25303);
nor UO_99 (O_99,N_27586,N_23393);
or UO_100 (O_100,N_28652,N_28591);
and UO_101 (O_101,N_22028,N_25041);
nor UO_102 (O_102,N_29471,N_24251);
nor UO_103 (O_103,N_26362,N_23941);
xnor UO_104 (O_104,N_24140,N_22865);
and UO_105 (O_105,N_27074,N_27095);
nand UO_106 (O_106,N_23628,N_23271);
nand UO_107 (O_107,N_27687,N_22425);
xor UO_108 (O_108,N_20044,N_25246);
nor UO_109 (O_109,N_26858,N_27785);
and UO_110 (O_110,N_25802,N_25257);
and UO_111 (O_111,N_21701,N_27587);
nor UO_112 (O_112,N_28015,N_20979);
or UO_113 (O_113,N_20206,N_27865);
or UO_114 (O_114,N_24667,N_25829);
and UO_115 (O_115,N_25308,N_20241);
xor UO_116 (O_116,N_22525,N_24239);
and UO_117 (O_117,N_25558,N_24503);
or UO_118 (O_118,N_25610,N_20355);
or UO_119 (O_119,N_27651,N_28871);
nand UO_120 (O_120,N_23684,N_21304);
xnor UO_121 (O_121,N_21512,N_28131);
xor UO_122 (O_122,N_24247,N_26643);
nor UO_123 (O_123,N_25625,N_28210);
or UO_124 (O_124,N_23200,N_26546);
nand UO_125 (O_125,N_20335,N_24117);
and UO_126 (O_126,N_24943,N_23122);
nand UO_127 (O_127,N_28476,N_25548);
nand UO_128 (O_128,N_20452,N_25915);
xor UO_129 (O_129,N_27678,N_28405);
xor UO_130 (O_130,N_29035,N_29321);
nand UO_131 (O_131,N_22240,N_25359);
and UO_132 (O_132,N_22704,N_29367);
nor UO_133 (O_133,N_22598,N_23219);
and UO_134 (O_134,N_24529,N_23549);
nor UO_135 (O_135,N_21346,N_21713);
nand UO_136 (O_136,N_27558,N_20931);
or UO_137 (O_137,N_25352,N_22647);
or UO_138 (O_138,N_27858,N_21661);
nor UO_139 (O_139,N_27390,N_25143);
nor UO_140 (O_140,N_27663,N_26326);
xnor UO_141 (O_141,N_27788,N_20057);
nor UO_142 (O_142,N_29729,N_27649);
xor UO_143 (O_143,N_25397,N_21556);
or UO_144 (O_144,N_21354,N_28599);
xor UO_145 (O_145,N_28189,N_22204);
or UO_146 (O_146,N_25727,N_24179);
nand UO_147 (O_147,N_24232,N_22599);
xor UO_148 (O_148,N_21957,N_20503);
nor UO_149 (O_149,N_20600,N_26088);
or UO_150 (O_150,N_24926,N_24399);
xor UO_151 (O_151,N_24902,N_28762);
xor UO_152 (O_152,N_23079,N_20183);
nand UO_153 (O_153,N_25122,N_29913);
or UO_154 (O_154,N_23460,N_23093);
or UO_155 (O_155,N_29875,N_26124);
or UO_156 (O_156,N_25156,N_21253);
nand UO_157 (O_157,N_21906,N_26589);
xnor UO_158 (O_158,N_21712,N_21561);
or UO_159 (O_159,N_29014,N_27323);
nand UO_160 (O_160,N_24259,N_25853);
or UO_161 (O_161,N_21028,N_28235);
nand UO_162 (O_162,N_21004,N_22667);
and UO_163 (O_163,N_23094,N_20155);
and UO_164 (O_164,N_27079,N_22800);
nand UO_165 (O_165,N_26714,N_22306);
nand UO_166 (O_166,N_26015,N_23268);
and UO_167 (O_167,N_23256,N_26634);
or UO_168 (O_168,N_29425,N_29706);
and UO_169 (O_169,N_21680,N_28727);
nand UO_170 (O_170,N_28567,N_28667);
nor UO_171 (O_171,N_20907,N_20506);
xor UO_172 (O_172,N_22211,N_26115);
xnor UO_173 (O_173,N_20938,N_28637);
nor UO_174 (O_174,N_29326,N_26000);
or UO_175 (O_175,N_25071,N_21084);
nor UO_176 (O_176,N_23517,N_26481);
nand UO_177 (O_177,N_27255,N_24721);
nor UO_178 (O_178,N_22352,N_26904);
nand UO_179 (O_179,N_26120,N_24068);
nor UO_180 (O_180,N_24212,N_21241);
nand UO_181 (O_181,N_25263,N_20061);
xnor UO_182 (O_182,N_23888,N_29399);
nor UO_183 (O_183,N_20386,N_26770);
or UO_184 (O_184,N_21239,N_22417);
or UO_185 (O_185,N_28214,N_24306);
nand UO_186 (O_186,N_21468,N_24350);
xor UO_187 (O_187,N_23522,N_24941);
and UO_188 (O_188,N_26924,N_24102);
nand UO_189 (O_189,N_23365,N_27604);
nand UO_190 (O_190,N_27495,N_29205);
or UO_191 (O_191,N_26741,N_25053);
or UO_192 (O_192,N_27026,N_22860);
or UO_193 (O_193,N_27871,N_29076);
xnor UO_194 (O_194,N_23518,N_26220);
and UO_195 (O_195,N_22070,N_22069);
or UO_196 (O_196,N_21414,N_24581);
nand UO_197 (O_197,N_26162,N_29791);
or UO_198 (O_198,N_20409,N_28574);
or UO_199 (O_199,N_20991,N_26930);
xnor UO_200 (O_200,N_25520,N_29660);
or UO_201 (O_201,N_23090,N_21835);
nor UO_202 (O_202,N_23561,N_27088);
nand UO_203 (O_203,N_22679,N_23423);
nand UO_204 (O_204,N_27704,N_27376);
nand UO_205 (O_205,N_27679,N_29755);
or UO_206 (O_206,N_26418,N_22513);
or UO_207 (O_207,N_29903,N_22630);
xnor UO_208 (O_208,N_28556,N_28912);
xnor UO_209 (O_209,N_26501,N_25140);
nand UO_210 (O_210,N_27765,N_26218);
or UO_211 (O_211,N_26303,N_20588);
or UO_212 (O_212,N_25979,N_26885);
nor UO_213 (O_213,N_25652,N_29292);
xor UO_214 (O_214,N_27379,N_21806);
xor UO_215 (O_215,N_21179,N_28164);
and UO_216 (O_216,N_29091,N_23433);
and UO_217 (O_217,N_23547,N_24601);
and UO_218 (O_218,N_25613,N_21555);
nand UO_219 (O_219,N_23294,N_29685);
nand UO_220 (O_220,N_23956,N_22124);
or UO_221 (O_221,N_23237,N_27856);
and UO_222 (O_222,N_28788,N_24550);
or UO_223 (O_223,N_23444,N_23623);
and UO_224 (O_224,N_26297,N_23220);
nand UO_225 (O_225,N_27993,N_22972);
or UO_226 (O_226,N_29950,N_27263);
nand UO_227 (O_227,N_21319,N_22230);
and UO_228 (O_228,N_25087,N_24542);
nand UO_229 (O_229,N_29462,N_23028);
nor UO_230 (O_230,N_27018,N_21021);
or UO_231 (O_231,N_23916,N_25533);
and UO_232 (O_232,N_27365,N_23412);
or UO_233 (O_233,N_27948,N_23875);
xnor UO_234 (O_234,N_24272,N_28867);
nand UO_235 (O_235,N_23894,N_24107);
and UO_236 (O_236,N_25391,N_24050);
xnor UO_237 (O_237,N_29436,N_21023);
and UO_238 (O_238,N_23051,N_29662);
nand UO_239 (O_239,N_27894,N_23148);
nor UO_240 (O_240,N_28471,N_28790);
and UO_241 (O_241,N_23356,N_23750);
xnor UO_242 (O_242,N_28101,N_25779);
nor UO_243 (O_243,N_24580,N_25205);
xor UO_244 (O_244,N_21485,N_27647);
xnor UO_245 (O_245,N_26794,N_20944);
nor UO_246 (O_246,N_28597,N_21756);
and UO_247 (O_247,N_24127,N_24914);
and UO_248 (O_248,N_25602,N_28674);
and UO_249 (O_249,N_26573,N_29335);
or UO_250 (O_250,N_25767,N_27052);
nand UO_251 (O_251,N_28263,N_27083);
or UO_252 (O_252,N_26996,N_22173);
nand UO_253 (O_253,N_25192,N_29547);
nor UO_254 (O_254,N_26646,N_25799);
nand UO_255 (O_255,N_25286,N_24265);
nor UO_256 (O_256,N_28916,N_28927);
xnor UO_257 (O_257,N_23685,N_26555);
and UO_258 (O_258,N_20231,N_28562);
and UO_259 (O_259,N_20612,N_28376);
and UO_260 (O_260,N_22741,N_25810);
or UO_261 (O_261,N_24559,N_29297);
nand UO_262 (O_262,N_29290,N_28314);
and UO_263 (O_263,N_25183,N_21036);
nand UO_264 (O_264,N_27686,N_22043);
nor UO_265 (O_265,N_25050,N_22516);
nor UO_266 (O_266,N_28618,N_27508);
nand UO_267 (O_267,N_26074,N_26541);
and UO_268 (O_268,N_21355,N_24031);
xor UO_269 (O_269,N_20367,N_27186);
and UO_270 (O_270,N_26237,N_23490);
nor UO_271 (O_271,N_29837,N_26467);
or UO_272 (O_272,N_26593,N_20048);
nor UO_273 (O_273,N_25262,N_21518);
nand UO_274 (O_274,N_28384,N_29589);
and UO_275 (O_275,N_20752,N_23273);
nand UO_276 (O_276,N_27328,N_26049);
and UO_277 (O_277,N_29924,N_24091);
xnor UO_278 (O_278,N_26421,N_21930);
xnor UO_279 (O_279,N_24798,N_26915);
and UO_280 (O_280,N_28328,N_22214);
xnor UO_281 (O_281,N_29413,N_23025);
and UO_282 (O_282,N_22483,N_29942);
nor UO_283 (O_283,N_20982,N_25392);
or UO_284 (O_284,N_29974,N_22523);
nand UO_285 (O_285,N_24098,N_21515);
and UO_286 (O_286,N_26485,N_29743);
nor UO_287 (O_287,N_21394,N_27939);
nand UO_288 (O_288,N_24092,N_29977);
xnor UO_289 (O_289,N_29029,N_26213);
nor UO_290 (O_290,N_20166,N_25467);
nand UO_291 (O_291,N_29510,N_29626);
nor UO_292 (O_292,N_20123,N_26903);
xor UO_293 (O_293,N_26189,N_23275);
and UO_294 (O_294,N_29995,N_23502);
nor UO_295 (O_295,N_28308,N_27067);
nand UO_296 (O_296,N_24975,N_23933);
and UO_297 (O_297,N_25433,N_26656);
nor UO_298 (O_298,N_21206,N_28163);
xor UO_299 (O_299,N_21049,N_24434);
and UO_300 (O_300,N_28954,N_28712);
xnor UO_301 (O_301,N_29621,N_28932);
or UO_302 (O_302,N_25996,N_22465);
or UO_303 (O_303,N_29204,N_23942);
nor UO_304 (O_304,N_25428,N_20385);
or UO_305 (O_305,N_29537,N_25436);
xnor UO_306 (O_306,N_28527,N_22359);
nand UO_307 (O_307,N_29473,N_24401);
xor UO_308 (O_308,N_28811,N_29691);
and UO_309 (O_309,N_23981,N_28453);
or UO_310 (O_310,N_29444,N_26462);
nand UO_311 (O_311,N_27728,N_29516);
nor UO_312 (O_312,N_29343,N_28253);
xnor UO_313 (O_313,N_25978,N_26772);
nor UO_314 (O_314,N_21915,N_20286);
xnor UO_315 (O_315,N_21125,N_21509);
xor UO_316 (O_316,N_23687,N_22958);
and UO_317 (O_317,N_21466,N_28627);
nor UO_318 (O_318,N_29971,N_25547);
nand UO_319 (O_319,N_21597,N_22015);
and UO_320 (O_320,N_22581,N_20482);
xor UO_321 (O_321,N_22934,N_28904);
or UO_322 (O_322,N_24541,N_26999);
xor UO_323 (O_323,N_26702,N_28897);
nand UO_324 (O_324,N_20472,N_27172);
and UO_325 (O_325,N_22781,N_24166);
xnor UO_326 (O_326,N_20992,N_20086);
xnor UO_327 (O_327,N_28483,N_24508);
and UO_328 (O_328,N_23054,N_29676);
or UO_329 (O_329,N_22315,N_26260);
or UO_330 (O_330,N_25088,N_28672);
nand UO_331 (O_331,N_23248,N_28054);
nand UO_332 (O_332,N_29910,N_28862);
xnor UO_333 (O_333,N_24822,N_26872);
nand UO_334 (O_334,N_23466,N_28403);
nor UO_335 (O_335,N_25942,N_29570);
nor UO_336 (O_336,N_22221,N_27970);
nand UO_337 (O_337,N_26395,N_29252);
or UO_338 (O_338,N_24426,N_29655);
and UO_339 (O_339,N_28411,N_23543);
xnor UO_340 (O_340,N_22900,N_24560);
nor UO_341 (O_341,N_22452,N_26572);
and UO_342 (O_342,N_28989,N_22320);
or UO_343 (O_343,N_22205,N_22401);
or UO_344 (O_344,N_24199,N_22438);
or UO_345 (O_345,N_25776,N_21995);
nor UO_346 (O_346,N_20978,N_22999);
and UO_347 (O_347,N_23193,N_23195);
nor UO_348 (O_348,N_21243,N_22330);
nor UO_349 (O_349,N_21975,N_24838);
and UO_350 (O_350,N_22990,N_21795);
or UO_351 (O_351,N_21948,N_27378);
or UO_352 (O_352,N_20292,N_21735);
and UO_353 (O_353,N_21069,N_20913);
nor UO_354 (O_354,N_26809,N_23679);
xor UO_355 (O_355,N_26013,N_20954);
xnor UO_356 (O_356,N_23788,N_28292);
xor UO_357 (O_357,N_21374,N_20906);
nand UO_358 (O_358,N_20419,N_25118);
and UO_359 (O_359,N_28644,N_28070);
nor UO_360 (O_360,N_24643,N_21145);
nand UO_361 (O_361,N_27322,N_25031);
xnor UO_362 (O_362,N_26948,N_29144);
xor UO_363 (O_363,N_22715,N_21208);
and UO_364 (O_364,N_25939,N_21237);
nand UO_365 (O_365,N_22314,N_24123);
or UO_366 (O_366,N_26038,N_26113);
xor UO_367 (O_367,N_21506,N_24590);
or UO_368 (O_368,N_25235,N_22755);
xnor UO_369 (O_369,N_21811,N_20222);
and UO_370 (O_370,N_25043,N_24824);
and UO_371 (O_371,N_26361,N_28234);
or UO_372 (O_372,N_21583,N_21902);
nand UO_373 (O_373,N_23633,N_20772);
xnor UO_374 (O_374,N_26508,N_26958);
nor UO_375 (O_375,N_24255,N_25867);
xnor UO_376 (O_376,N_28450,N_24725);
and UO_377 (O_377,N_29781,N_29178);
and UO_378 (O_378,N_26438,N_22998);
nor UO_379 (O_379,N_26763,N_25046);
nand UO_380 (O_380,N_22568,N_29500);
nand UO_381 (O_381,N_21582,N_28829);
xnor UO_382 (O_382,N_23738,N_26587);
nor UO_383 (O_383,N_23850,N_23613);
nand UO_384 (O_384,N_26808,N_25596);
nand UO_385 (O_385,N_27893,N_25967);
and UO_386 (O_386,N_23331,N_24263);
or UO_387 (O_387,N_23076,N_29438);
and UO_388 (O_388,N_26684,N_23147);
nor UO_389 (O_389,N_24490,N_29806);
and UO_390 (O_390,N_21729,N_23109);
or UO_391 (O_391,N_27325,N_23014);
xor UO_392 (O_392,N_25682,N_24499);
or UO_393 (O_393,N_20273,N_29301);
or UO_394 (O_394,N_26201,N_28332);
nor UO_395 (O_395,N_25772,N_24528);
xor UO_396 (O_396,N_20512,N_26072);
or UO_397 (O_397,N_22253,N_29307);
xnor UO_398 (O_398,N_20749,N_23723);
and UO_399 (O_399,N_24891,N_28919);
and UO_400 (O_400,N_25376,N_21095);
or UO_401 (O_401,N_22447,N_29992);
or UO_402 (O_402,N_29891,N_22486);
or UO_403 (O_403,N_28045,N_24788);
nand UO_404 (O_404,N_27283,N_27915);
and UO_405 (O_405,N_26651,N_29164);
or UO_406 (O_406,N_27577,N_22379);
nand UO_407 (O_407,N_27846,N_20646);
and UO_408 (O_408,N_27812,N_22199);
or UO_409 (O_409,N_20710,N_26472);
nand UO_410 (O_410,N_21747,N_21122);
nand UO_411 (O_411,N_28512,N_27468);
xnor UO_412 (O_412,N_28447,N_26222);
or UO_413 (O_413,N_28639,N_23635);
or UO_414 (O_414,N_26112,N_26839);
nor UO_415 (O_415,N_20112,N_23711);
or UO_416 (O_416,N_22514,N_25442);
xnor UO_417 (O_417,N_20633,N_21492);
and UO_418 (O_418,N_23794,N_27119);
and UO_419 (O_419,N_23461,N_26860);
or UO_420 (O_420,N_23611,N_21154);
or UO_421 (O_421,N_25838,N_29238);
nand UO_422 (O_422,N_21242,N_20669);
and UO_423 (O_423,N_21071,N_24354);
and UO_424 (O_424,N_21008,N_24175);
nor UO_425 (O_425,N_27592,N_26217);
xnor UO_426 (O_426,N_24849,N_22080);
or UO_427 (O_427,N_26936,N_29771);
xor UO_428 (O_428,N_26020,N_22061);
and UO_429 (O_429,N_25028,N_27727);
and UO_430 (O_430,N_20376,N_20617);
or UO_431 (O_431,N_27125,N_24230);
nor UO_432 (O_432,N_24322,N_21904);
nor UO_433 (O_433,N_21896,N_20179);
xnor UO_434 (O_434,N_23784,N_21530);
nand UO_435 (O_435,N_26516,N_21333);
or UO_436 (O_436,N_24246,N_24723);
or UO_437 (O_437,N_21349,N_28694);
xor UO_438 (O_438,N_27016,N_23255);
nor UO_439 (O_439,N_27639,N_23763);
or UO_440 (O_440,N_26601,N_22653);
nand UO_441 (O_441,N_24922,N_22722);
or UO_442 (O_442,N_26874,N_20025);
or UO_443 (O_443,N_29863,N_28933);
nand UO_444 (O_444,N_20724,N_23389);
or UO_445 (O_445,N_27772,N_23917);
xor UO_446 (O_446,N_24205,N_20963);
and UO_447 (O_447,N_20664,N_28196);
and UO_448 (O_448,N_25066,N_28141);
or UO_449 (O_449,N_25760,N_28740);
and UO_450 (O_450,N_23265,N_29475);
or UO_451 (O_451,N_29116,N_23144);
and UO_452 (O_452,N_28282,N_24270);
nand UO_453 (O_453,N_20125,N_22424);
nand UO_454 (O_454,N_26529,N_23787);
or UO_455 (O_455,N_27518,N_29682);
xnor UO_456 (O_456,N_25385,N_23217);
nand UO_457 (O_457,N_29721,N_20528);
nor UO_458 (O_458,N_25751,N_24382);
or UO_459 (O_459,N_22166,N_22909);
or UO_460 (O_460,N_22319,N_22000);
or UO_461 (O_461,N_23886,N_27448);
xnor UO_462 (O_462,N_22249,N_24911);
nor UO_463 (O_463,N_22074,N_28963);
and UO_464 (O_464,N_23993,N_24796);
xor UO_465 (O_465,N_28857,N_22948);
nand UO_466 (O_466,N_29128,N_22884);
and UO_467 (O_467,N_29577,N_23621);
nand UO_468 (O_468,N_25109,N_28393);
nor UO_469 (O_469,N_23746,N_29047);
and UO_470 (O_470,N_22362,N_24720);
and UO_471 (O_471,N_28456,N_26613);
nor UO_472 (O_472,N_21168,N_27046);
and UO_473 (O_473,N_20330,N_24664);
xnor UO_474 (O_474,N_21900,N_23211);
nand UO_475 (O_475,N_22120,N_23602);
and UO_476 (O_476,N_27386,N_28333);
xor UO_477 (O_477,N_21647,N_27660);
nor UO_478 (O_478,N_26673,N_25569);
nor UO_479 (O_479,N_27807,N_22605);
or UO_480 (O_480,N_22446,N_25860);
xor UO_481 (O_481,N_29106,N_26003);
or UO_482 (O_482,N_22340,N_20535);
nor UO_483 (O_483,N_28479,N_20174);
and UO_484 (O_484,N_25124,N_27701);
and UO_485 (O_485,N_28749,N_25646);
nor UO_486 (O_486,N_25675,N_29293);
nor UO_487 (O_487,N_25980,N_25791);
and UO_488 (O_488,N_27972,N_21800);
nand UO_489 (O_489,N_21877,N_21110);
xor UO_490 (O_490,N_24652,N_22740);
nand UO_491 (O_491,N_28280,N_21379);
nor UO_492 (O_492,N_26047,N_28646);
and UO_493 (O_493,N_28175,N_26765);
and UO_494 (O_494,N_23057,N_20322);
nor UO_495 (O_495,N_20893,N_20426);
and UO_496 (O_496,N_28178,N_27147);
xnor UO_497 (O_497,N_22463,N_23596);
nand UO_498 (O_498,N_26611,N_21015);
xor UO_499 (O_499,N_21694,N_22664);
nand UO_500 (O_500,N_27169,N_27874);
and UO_501 (O_501,N_26704,N_27299);
nor UO_502 (O_502,N_28521,N_26185);
and UO_503 (O_503,N_25993,N_27839);
nand UO_504 (O_504,N_20391,N_24466);
nand UO_505 (O_505,N_22949,N_21097);
or UO_506 (O_506,N_20841,N_25892);
and UO_507 (O_507,N_21495,N_28844);
or UO_508 (O_508,N_20433,N_29485);
nand UO_509 (O_509,N_23173,N_25540);
and UO_510 (O_510,N_20235,N_21707);
nand UO_511 (O_511,N_20983,N_29658);
xnor UO_512 (O_512,N_28842,N_22660);
xnor UO_513 (O_513,N_26321,N_21790);
nor UO_514 (O_514,N_29772,N_20793);
xnor UO_515 (O_515,N_25111,N_27453);
xor UO_516 (O_516,N_27713,N_24473);
or UO_517 (O_517,N_27392,N_23732);
and UO_518 (O_518,N_22591,N_24141);
nand UO_519 (O_519,N_23092,N_25460);
nand UO_520 (O_520,N_28258,N_24913);
nand UO_521 (O_521,N_27474,N_20972);
and UO_522 (O_522,N_22720,N_20853);
xor UO_523 (O_523,N_26106,N_29253);
or UO_524 (O_524,N_28362,N_20595);
and UO_525 (O_525,N_29998,N_21058);
nand UO_526 (O_526,N_26797,N_22977);
xor UO_527 (O_527,N_20758,N_26137);
nand UO_528 (O_528,N_28546,N_23185);
and UO_529 (O_529,N_25474,N_25306);
nand UO_530 (O_530,N_26221,N_26785);
or UO_531 (O_531,N_23453,N_27093);
and UO_532 (O_532,N_28551,N_27339);
and UO_533 (O_533,N_22258,N_29575);
and UO_534 (O_534,N_20774,N_23330);
and UO_535 (O_535,N_28434,N_21940);
nor UO_536 (O_536,N_27277,N_21480);
nor UO_537 (O_537,N_25907,N_25989);
or UO_538 (O_538,N_25349,N_23398);
xnor UO_539 (O_539,N_27268,N_21928);
and UO_540 (O_540,N_27245,N_27087);
nand UO_541 (O_541,N_21803,N_26931);
and UO_542 (O_542,N_24330,N_25084);
and UO_543 (O_543,N_21157,N_29149);
xor UO_544 (O_544,N_28304,N_21309);
nand UO_545 (O_545,N_26151,N_28702);
nand UO_546 (O_546,N_23311,N_29230);
xnor UO_547 (O_547,N_28522,N_21683);
and UO_548 (O_548,N_23584,N_29853);
nand UO_549 (O_549,N_27835,N_26405);
and UO_550 (O_550,N_25094,N_26869);
and UO_551 (O_551,N_22648,N_23416);
xnor UO_552 (O_552,N_20594,N_23863);
nand UO_553 (O_553,N_27773,N_21884);
xor UO_554 (O_554,N_20280,N_29526);
xor UO_555 (O_555,N_29006,N_21898);
nand UO_556 (O_556,N_29848,N_28699);
nand UO_557 (O_557,N_24925,N_21637);
nor UO_558 (O_558,N_20263,N_25230);
and UO_559 (O_559,N_21225,N_21432);
or UO_560 (O_560,N_24520,N_20113);
xor UO_561 (O_561,N_22944,N_23228);
and UO_562 (O_562,N_25346,N_29988);
xor UO_563 (O_563,N_20420,N_26678);
xor UO_564 (O_564,N_22206,N_28690);
nand UO_565 (O_565,N_25137,N_26916);
nor UO_566 (O_566,N_25742,N_26128);
or UO_567 (O_567,N_20417,N_25403);
or UO_568 (O_568,N_29654,N_20817);
xnor UO_569 (O_569,N_20769,N_24688);
nand UO_570 (O_570,N_24498,N_26341);
nand UO_571 (O_571,N_23050,N_23554);
xor UO_572 (O_572,N_20831,N_23533);
and UO_573 (O_573,N_20331,N_29479);
or UO_574 (O_574,N_28432,N_26122);
and UO_575 (O_575,N_28010,N_29303);
nand UO_576 (O_576,N_28064,N_24128);
nand UO_577 (O_577,N_28953,N_23366);
and UO_578 (O_578,N_23493,N_26699);
and UO_579 (O_579,N_22835,N_22457);
xor UO_580 (O_580,N_22824,N_24794);
or UO_581 (O_581,N_20049,N_23164);
and UO_582 (O_582,N_20495,N_29689);
nor UO_583 (O_583,N_29879,N_25959);
nand UO_584 (O_584,N_24947,N_28062);
nand UO_585 (O_585,N_22443,N_20598);
nor UO_586 (O_586,N_22965,N_25065);
or UO_587 (O_587,N_20291,N_20271);
and UO_588 (O_588,N_22878,N_27753);
or UO_589 (O_589,N_29960,N_23158);
and UO_590 (O_590,N_27171,N_26676);
and UO_591 (O_591,N_20450,N_27776);
nand UO_592 (O_592,N_21429,N_29745);
and UO_593 (O_593,N_26698,N_29090);
nor UO_594 (O_594,N_29226,N_26258);
or UO_595 (O_595,N_20866,N_23995);
and UO_596 (O_596,N_24281,N_24965);
xnor UO_597 (O_597,N_24589,N_21431);
nand UO_598 (O_598,N_26866,N_25788);
and UO_599 (O_599,N_24754,N_21151);
and UO_600 (O_600,N_20971,N_21257);
or UO_601 (O_601,N_22499,N_23903);
and UO_602 (O_602,N_27711,N_27570);
and UO_603 (O_603,N_22923,N_28970);
xnor UO_604 (O_604,N_26093,N_22501);
or UO_605 (O_605,N_21964,N_20212);
and UO_606 (O_606,N_23341,N_21175);
nor UO_607 (O_607,N_22172,N_21240);
and UO_608 (O_608,N_27425,N_22311);
nor UO_609 (O_609,N_26401,N_21844);
nand UO_610 (O_610,N_23911,N_28083);
nand UO_611 (O_611,N_26720,N_27973);
nand UO_612 (O_612,N_23890,N_29207);
nor UO_613 (O_613,N_20483,N_21141);
nor UO_614 (O_614,N_23540,N_21655);
nand UO_615 (O_615,N_22461,N_29907);
xnor UO_616 (O_616,N_25394,N_28524);
or UO_617 (O_617,N_22476,N_25049);
xnor UO_618 (O_618,N_23108,N_20532);
or UO_619 (O_619,N_20712,N_27541);
nor UO_620 (O_620,N_26121,N_24022);
nor UO_621 (O_621,N_21025,N_22779);
or UO_622 (O_622,N_29211,N_25503);
and UO_623 (O_623,N_23666,N_27954);
or UO_624 (O_624,N_28255,N_20530);
xor UO_625 (O_625,N_29890,N_23053);
xnor UO_626 (O_626,N_23996,N_23722);
nand UO_627 (O_627,N_25007,N_25325);
xnor UO_628 (O_628,N_20953,N_26461);
or UO_629 (O_629,N_22164,N_21186);
nand UO_630 (O_630,N_24953,N_25382);
nor UO_631 (O_631,N_21463,N_23627);
nand UO_632 (O_632,N_29719,N_24004);
and UO_633 (O_633,N_28715,N_20959);
nor UO_634 (O_634,N_27606,N_22469);
xor UO_635 (O_635,N_20674,N_23809);
nor UO_636 (O_636,N_23680,N_23812);
nor UO_637 (O_637,N_25412,N_23162);
xnor UO_638 (O_638,N_29309,N_28595);
nand UO_639 (O_639,N_27533,N_24229);
or UO_640 (O_640,N_29448,N_25822);
xnor UO_641 (O_641,N_28858,N_24383);
nor UO_642 (O_642,N_28596,N_20510);
nand UO_643 (O_643,N_20270,N_28143);
nor UO_644 (O_644,N_24719,N_25777);
nor UO_645 (O_645,N_21426,N_28686);
xor UO_646 (O_646,N_26239,N_24262);
nand UO_647 (O_647,N_23819,N_21214);
and UO_648 (O_648,N_20949,N_22400);
nor UO_649 (O_649,N_29385,N_27118);
nand UO_650 (O_650,N_23487,N_27105);
and UO_651 (O_651,N_29333,N_29266);
xnor UO_652 (O_652,N_26272,N_26010);
xnor UO_653 (O_653,N_25817,N_20374);
or UO_654 (O_654,N_27675,N_25465);
nand UO_655 (O_655,N_22729,N_21303);
nor UO_656 (O_656,N_22115,N_22775);
nand UO_657 (O_657,N_28168,N_22145);
nor UO_658 (O_658,N_25454,N_27389);
xnor UO_659 (O_659,N_22506,N_26017);
xor UO_660 (O_660,N_29920,N_21192);
nand UO_661 (O_661,N_23636,N_27430);
or UO_662 (O_662,N_26308,N_24878);
and UO_663 (O_663,N_21599,N_20201);
nand UO_664 (O_664,N_22391,N_29043);
xor UO_665 (O_665,N_25773,N_20933);
and UO_666 (O_666,N_26367,N_25703);
nand UO_667 (O_667,N_20020,N_26653);
nor UO_668 (O_668,N_27363,N_26751);
nor UO_669 (O_669,N_28771,N_26782);
nand UO_670 (O_670,N_23660,N_26721);
or UO_671 (O_671,N_26956,N_23339);
and UO_672 (O_672,N_29443,N_29071);
and UO_673 (O_673,N_26034,N_24848);
and UO_674 (O_674,N_25592,N_25893);
xnor UO_675 (O_675,N_20052,N_29511);
and UO_676 (O_676,N_25237,N_24787);
nor UO_677 (O_677,N_20184,N_20540);
nand UO_678 (O_678,N_24186,N_22468);
or UO_679 (O_679,N_25146,N_22585);
nand UO_680 (O_680,N_26660,N_29060);
and UO_681 (O_681,N_23404,N_29683);
nor UO_682 (O_682,N_24961,N_24215);
and UO_683 (O_683,N_29376,N_27658);
nor UO_684 (O_684,N_29667,N_29722);
and UO_685 (O_685,N_20660,N_22783);
and UO_686 (O_686,N_29159,N_25298);
or UO_687 (O_687,N_29084,N_28793);
and UO_688 (O_688,N_26412,N_21665);
nand UO_689 (O_689,N_25933,N_25781);
and UO_690 (O_690,N_24018,N_27996);
and UO_691 (O_691,N_24211,N_27097);
nand UO_692 (O_692,N_23036,N_20371);
nor UO_693 (O_693,N_20628,N_24669);
and UO_694 (O_694,N_24220,N_29156);
xor UO_695 (O_695,N_26071,N_22108);
nor UO_696 (O_696,N_22666,N_28778);
and UO_697 (O_697,N_29501,N_27547);
xor UO_698 (O_698,N_25567,N_20312);
or UO_699 (O_699,N_20804,N_21892);
and UO_700 (O_700,N_21670,N_20050);
nand UO_701 (O_701,N_26193,N_26195);
and UO_702 (O_702,N_22535,N_22122);
xnor UO_703 (O_703,N_27029,N_25778);
nor UO_704 (O_704,N_22897,N_28903);
and UO_705 (O_705,N_27719,N_28295);
nor UO_706 (O_706,N_28950,N_23080);
nand UO_707 (O_707,N_20726,N_22682);
nor UO_708 (O_708,N_25139,N_20802);
xnor UO_709 (O_709,N_24058,N_24155);
or UO_710 (O_710,N_25476,N_23134);
xor UO_711 (O_711,N_20478,N_20464);
nor UO_712 (O_712,N_25138,N_28029);
and UO_713 (O_713,N_22684,N_27828);
or UO_714 (O_714,N_25399,N_26053);
or UO_715 (O_715,N_27123,N_27158);
and UO_716 (O_716,N_27232,N_28194);
or UO_717 (O_717,N_22578,N_28800);
or UO_718 (O_718,N_25416,N_26582);
and UO_719 (O_719,N_22512,N_24409);
or UO_720 (O_720,N_21528,N_25747);
and UO_721 (O_721,N_29009,N_22327);
or UO_722 (O_722,N_25056,N_23182);
and UO_723 (O_723,N_22559,N_22064);
and UO_724 (O_724,N_29637,N_28606);
or UO_725 (O_725,N_21105,N_23604);
xor UO_726 (O_726,N_29107,N_27608);
or UO_727 (O_727,N_20800,N_29460);
nand UO_728 (O_728,N_22959,N_27467);
and UO_729 (O_729,N_24915,N_28755);
and UO_730 (O_730,N_22739,N_29003);
or UO_731 (O_731,N_26557,N_29671);
nand UO_732 (O_732,N_26985,N_21029);
nand UO_733 (O_733,N_22395,N_23421);
or UO_734 (O_734,N_26562,N_27203);
nor UO_735 (O_735,N_22955,N_22298);
xor UO_736 (O_736,N_24962,N_29940);
nor UO_737 (O_737,N_29748,N_26114);
xnor UO_738 (O_738,N_25642,N_28018);
or UO_739 (O_739,N_22435,N_24457);
xor UO_740 (O_740,N_26450,N_29147);
xnor UO_741 (O_741,N_24315,N_24321);
nand UO_742 (O_742,N_26517,N_26639);
and UO_743 (O_743,N_28995,N_20032);
and UO_744 (O_744,N_25380,N_21484);
nor UO_745 (O_745,N_22552,N_20768);
nand UO_746 (O_746,N_27932,N_24582);
and UO_747 (O_747,N_22920,N_29400);
nand UO_748 (O_748,N_21682,N_23003);
or UO_749 (O_749,N_27182,N_21411);
nor UO_750 (O_750,N_25152,N_20780);
nand UO_751 (O_751,N_27375,N_25249);
xor UO_752 (O_752,N_24196,N_28046);
nor UO_753 (O_753,N_28737,N_28984);
nand UO_754 (O_754,N_21502,N_20544);
xnor UO_755 (O_755,N_20662,N_21378);
xnor UO_756 (O_756,N_21755,N_27936);
or UO_757 (O_757,N_28153,N_24496);
xor UO_758 (O_758,N_27153,N_28869);
nand UO_759 (O_759,N_25108,N_28767);
and UO_760 (O_760,N_22546,N_26142);
and UO_761 (O_761,N_28601,N_23020);
nand UO_762 (O_762,N_20122,N_21081);
and UO_763 (O_763,N_22932,N_23473);
or UO_764 (O_764,N_29218,N_25583);
or UO_765 (O_765,N_26825,N_25981);
and UO_766 (O_766,N_25713,N_20369);
nor UO_767 (O_767,N_26986,N_27111);
nand UO_768 (O_768,N_21859,N_29678);
or UO_769 (O_769,N_29932,N_28781);
nor UO_770 (O_770,N_29099,N_25841);
nor UO_771 (O_771,N_25620,N_29761);
nand UO_772 (O_772,N_24165,N_20224);
xor UO_773 (O_773,N_21924,N_28825);
nor UO_774 (O_774,N_25895,N_26416);
nor UO_775 (O_775,N_20722,N_29185);
or UO_776 (O_776,N_26090,N_26942);
nand UO_777 (O_777,N_25443,N_24075);
xnor UO_778 (O_778,N_24735,N_23323);
xor UO_779 (O_779,N_21608,N_28207);
xnor UO_780 (O_780,N_26062,N_23385);
nand UO_781 (O_781,N_21234,N_25350);
nand UO_782 (O_782,N_22375,N_25008);
nand UO_783 (O_783,N_22906,N_25764);
or UO_784 (O_784,N_27797,N_22594);
or UO_785 (O_785,N_22092,N_29864);
and UO_786 (O_786,N_26520,N_20950);
xnor UO_787 (O_787,N_26618,N_29124);
and UO_788 (O_788,N_21344,N_25889);
or UO_789 (O_789,N_25794,N_27671);
nor UO_790 (O_790,N_25265,N_22873);
nor UO_791 (O_791,N_29018,N_22290);
and UO_792 (O_792,N_24195,N_27837);
and UO_793 (O_793,N_28499,N_21138);
xnor UO_794 (O_794,N_29978,N_21451);
xnor UO_795 (O_795,N_27135,N_23467);
or UO_796 (O_796,N_20733,N_22964);
xor UO_797 (O_797,N_23800,N_28985);
xnor UO_798 (O_798,N_28581,N_27584);
or UO_799 (O_799,N_25271,N_29421);
nor UO_800 (O_800,N_28723,N_20164);
nor UO_801 (O_801,N_25577,N_28167);
nand UO_802 (O_802,N_28915,N_21345);
xor UO_803 (O_803,N_24260,N_27580);
or UO_804 (O_804,N_22307,N_27600);
and UO_805 (O_805,N_20014,N_28034);
and UO_806 (O_806,N_23957,N_20943);
xnor UO_807 (O_807,N_28538,N_26801);
xnor UO_808 (O_808,N_29630,N_27341);
xnor UO_809 (O_809,N_22636,N_26837);
xnor UO_810 (O_810,N_24924,N_28334);
and UO_811 (O_811,N_20822,N_26759);
or UO_812 (O_812,N_20999,N_23867);
xor UO_813 (O_813,N_28589,N_25505);
nand UO_814 (O_814,N_25324,N_27857);
xor UO_815 (O_815,N_28728,N_21576);
or UO_816 (O_816,N_25212,N_22810);
nand UO_817 (O_817,N_29862,N_28240);
nor UO_818 (O_818,N_20071,N_22176);
xor UO_819 (O_819,N_28392,N_24976);
nor UO_820 (O_820,N_25141,N_23439);
nand UO_821 (O_821,N_27145,N_29470);
nor UO_822 (O_822,N_27833,N_27820);
nand UO_823 (O_823,N_28766,N_29336);
and UO_824 (O_824,N_26532,N_29801);
xor UO_825 (O_825,N_28760,N_23432);
nor UO_826 (O_826,N_27132,N_21692);
nor UO_827 (O_827,N_29657,N_25696);
xor UO_828 (O_828,N_20111,N_23950);
nand UO_829 (O_829,N_25664,N_28149);
and UO_830 (O_830,N_25881,N_26749);
or UO_831 (O_831,N_29546,N_28910);
and UO_832 (O_832,N_27114,N_26586);
nand UO_833 (O_833,N_27454,N_29580);
nor UO_834 (O_834,N_23739,N_29272);
or UO_835 (O_835,N_24152,N_23320);
xor UO_836 (O_836,N_22245,N_29563);
and UO_837 (O_837,N_26104,N_27722);
xnor UO_838 (O_838,N_23649,N_22444);
or UO_839 (O_839,N_23400,N_27291);
or UO_840 (O_840,N_28338,N_24879);
and UO_841 (O_841,N_21705,N_21180);
and UO_842 (O_842,N_27116,N_29778);
nor UO_843 (O_843,N_21026,N_26991);
and UO_844 (O_844,N_23697,N_22046);
xnor UO_845 (O_845,N_27876,N_23362);
nor UO_846 (O_846,N_22197,N_21112);
nor UO_847 (O_847,N_21679,N_20867);
and UO_848 (O_848,N_24216,N_21788);
and UO_849 (O_849,N_24132,N_26380);
and UO_850 (O_850,N_23360,N_26052);
xor UO_851 (O_851,N_25218,N_28377);
nor UO_852 (O_852,N_22049,N_23716);
or UO_853 (O_853,N_25716,N_24681);
and UO_854 (O_854,N_25985,N_20746);
nor UO_855 (O_855,N_24865,N_22838);
or UO_856 (O_856,N_22278,N_20854);
nand UO_857 (O_857,N_22905,N_21471);
xor UO_858 (O_858,N_24460,N_23326);
or UO_859 (O_859,N_27381,N_28350);
nor UO_860 (O_860,N_27281,N_22803);
xnor UO_861 (O_861,N_22138,N_26323);
and UO_862 (O_862,N_20051,N_28429);
and UO_863 (O_863,N_22843,N_24945);
and UO_864 (O_864,N_27210,N_28417);
xnor UO_865 (O_865,N_29536,N_25916);
xor UO_866 (O_866,N_29102,N_26292);
and UO_867 (O_867,N_21275,N_28203);
nand UO_868 (O_868,N_27409,N_29059);
and UO_869 (O_869,N_23983,N_23381);
xor UO_870 (O_870,N_27529,N_23891);
xnor UO_871 (O_871,N_23292,N_25189);
and UO_872 (O_872,N_24623,N_24480);
nand UO_873 (O_873,N_25245,N_26692);
nor UO_874 (O_874,N_29857,N_20582);
or UO_875 (O_875,N_27944,N_24323);
xor UO_876 (O_876,N_24275,N_29941);
nor UO_877 (O_877,N_22832,N_20194);
and UO_878 (O_878,N_20154,N_20083);
or UO_879 (O_879,N_20634,N_25765);
nand UO_880 (O_880,N_28642,N_21818);
or UO_881 (O_881,N_20249,N_20159);
nand UO_882 (O_882,N_22619,N_27346);
or UO_883 (O_883,N_28040,N_24256);
xor UO_884 (O_884,N_29152,N_29954);
xnor UO_885 (O_885,N_23847,N_25126);
nor UO_886 (O_886,N_28495,N_20994);
and UO_887 (O_887,N_27034,N_27521);
and UO_888 (O_888,N_26132,N_21657);
xor UO_889 (O_889,N_27597,N_29555);
and UO_890 (O_890,N_27180,N_25831);
nor UO_891 (O_891,N_28057,N_25131);
nor UO_892 (O_892,N_28003,N_27302);
nor UO_893 (O_893,N_26475,N_24991);
xnor UO_894 (O_894,N_23671,N_20076);
nand UO_895 (O_895,N_28464,N_24125);
nor UO_896 (O_896,N_27082,N_20012);
or UO_897 (O_897,N_23695,N_26861);
or UO_898 (O_898,N_20789,N_26466);
nand UO_899 (O_899,N_24045,N_24101);
nand UO_900 (O_900,N_22938,N_26925);
and UO_901 (O_901,N_24425,N_28257);
or UO_902 (O_902,N_21640,N_22083);
or UO_903 (O_903,N_27064,N_29445);
or UO_904 (O_904,N_21946,N_27108);
xnor UO_905 (O_905,N_22159,N_29979);
xnor UO_906 (O_906,N_25733,N_21458);
nand UO_907 (O_907,N_24353,N_27729);
nor UO_908 (O_908,N_26432,N_29788);
or UO_909 (O_909,N_28682,N_20302);
xor UO_910 (O_910,N_21604,N_29236);
nor UO_911 (O_911,N_23103,N_23452);
nor UO_912 (O_912,N_28854,N_22409);
nor UO_913 (O_913,N_26795,N_26658);
or UO_914 (O_914,N_25196,N_20827);
and UO_915 (O_915,N_22480,N_26615);
or UO_916 (O_916,N_21761,N_27373);
xor UO_917 (O_917,N_20840,N_23455);
nor UO_918 (O_918,N_29562,N_23494);
and UO_919 (O_919,N_21276,N_29323);
nor UO_920 (O_920,N_25483,N_20881);
or UO_921 (O_921,N_26061,N_23954);
or UO_922 (O_922,N_27384,N_25462);
nand UO_923 (O_923,N_25082,N_29224);
and UO_924 (O_924,N_25932,N_27769);
nor UO_925 (O_925,N_23568,N_28502);
or UO_926 (O_926,N_27300,N_23588);
nand UO_927 (O_927,N_26975,N_27565);
nor UO_928 (O_928,N_28106,N_27628);
and UO_929 (O_929,N_27475,N_27219);
nor UO_930 (O_930,N_29967,N_23034);
nand UO_931 (O_931,N_25500,N_29062);
nand UO_932 (O_932,N_27199,N_26389);
xnor UO_933 (O_933,N_20686,N_24182);
xnor UO_934 (O_934,N_20730,N_24077);
nor UO_935 (O_935,N_25965,N_26600);
xnor UO_936 (O_936,N_20519,N_26584);
nand UO_937 (O_937,N_23121,N_28052);
nor UO_938 (O_938,N_28883,N_27275);
and UO_939 (O_939,N_23302,N_22641);
and UO_940 (O_940,N_29640,N_22616);
xor UO_941 (O_941,N_22241,N_21098);
nand UO_942 (O_942,N_25179,N_22600);
nor UO_943 (O_943,N_26834,N_24970);
nor UO_944 (O_944,N_22673,N_21926);
nand UO_945 (O_945,N_21171,N_27902);
xor UO_946 (O_946,N_20382,N_28299);
nor UO_947 (O_947,N_23456,N_24187);
and UO_948 (O_948,N_22728,N_20671);
xor UO_949 (O_949,N_29319,N_26492);
nor UO_950 (O_950,N_24521,N_29136);
nand UO_951 (O_951,N_28951,N_28394);
nor UO_952 (O_952,N_21501,N_26377);
and UO_953 (O_953,N_21155,N_20706);
nand UO_954 (O_954,N_22392,N_27292);
nand UO_955 (O_955,N_28577,N_25427);
nor UO_956 (O_956,N_25429,N_23128);
nand UO_957 (O_957,N_23437,N_21127);
and UO_958 (O_958,N_22057,N_24385);
xnor UO_959 (O_959,N_21216,N_27167);
nor UO_960 (O_960,N_29033,N_28422);
xor UO_961 (O_961,N_29277,N_21676);
nand UO_962 (O_962,N_26262,N_21944);
nand UO_963 (O_963,N_22045,N_22562);
nor UO_964 (O_964,N_20707,N_27151);
or UO_965 (O_965,N_20705,N_23579);
nand UO_966 (O_966,N_23177,N_26522);
and UO_967 (O_967,N_29410,N_26188);
and UO_968 (O_968,N_26539,N_29803);
nor UO_969 (O_969,N_24602,N_20653);
nor UO_970 (O_970,N_24191,N_20604);
xnor UO_971 (O_971,N_28939,N_21947);
and UO_972 (O_972,N_28821,N_26609);
nor UO_973 (O_973,N_29109,N_23449);
xor UO_974 (O_974,N_20845,N_20578);
xnor UO_975 (O_975,N_24314,N_27342);
and UO_976 (O_976,N_29263,N_20477);
or UO_977 (O_977,N_28138,N_25157);
nand UO_978 (O_978,N_27674,N_28848);
or UO_979 (O_979,N_28130,N_27733);
and UO_980 (O_980,N_26388,N_20250);
or UO_981 (O_981,N_24218,N_20082);
xnor UO_982 (O_982,N_27427,N_24403);
and UO_983 (O_983,N_28162,N_21751);
nand UO_984 (O_984,N_22202,N_24986);
xor UO_985 (O_985,N_21563,N_23428);
and UO_986 (O_986,N_21542,N_28120);
and UO_987 (O_987,N_24465,N_20922);
or UO_988 (O_988,N_20958,N_23946);
xnor UO_989 (O_989,N_22799,N_29012);
and UO_990 (O_990,N_28038,N_28269);
or UO_991 (O_991,N_25478,N_25095);
xnor UO_992 (O_992,N_29968,N_29364);
nor UO_993 (O_993,N_29219,N_20878);
and UO_994 (O_994,N_28529,N_28043);
xor UO_995 (O_995,N_28071,N_26465);
and UO_996 (O_996,N_20110,N_23895);
and UO_997 (O_997,N_21352,N_23840);
or UO_998 (O_998,N_28383,N_29300);
and UO_999 (O_999,N_22744,N_24411);
xor UO_1000 (O_1000,N_25954,N_26169);
xnor UO_1001 (O_1001,N_24968,N_23844);
and UO_1002 (O_1002,N_22526,N_25149);
or UO_1003 (O_1003,N_28687,N_27818);
or UO_1004 (O_1004,N_20139,N_26927);
xnor UO_1005 (O_1005,N_22262,N_22102);
xnor UO_1006 (O_1006,N_23184,N_22353);
or UO_1007 (O_1007,N_28863,N_26553);
xor UO_1008 (O_1008,N_26548,N_25338);
or UO_1009 (O_1009,N_21041,N_26006);
and UO_1010 (O_1010,N_27851,N_23753);
nor UO_1011 (O_1011,N_26080,N_23290);
nand UO_1012 (O_1012,N_25635,N_25461);
and UO_1013 (O_1013,N_23519,N_22317);
and UO_1014 (O_1014,N_21516,N_23654);
nor UO_1015 (O_1015,N_28491,N_21894);
and UO_1016 (O_1016,N_22784,N_28135);
nand UO_1017 (O_1017,N_20128,N_21016);
or UO_1018 (O_1018,N_27642,N_20172);
or UO_1019 (O_1019,N_28112,N_22582);
xor UO_1020 (O_1020,N_20351,N_22813);
nand UO_1021 (O_1021,N_22848,N_29909);
and UO_1022 (O_1022,N_21662,N_22357);
or UO_1023 (O_1023,N_22207,N_22343);
xnor UO_1024 (O_1024,N_27157,N_24842);
nor UO_1025 (O_1025,N_25530,N_24455);
xnor UO_1026 (O_1026,N_24717,N_20559);
xnor UO_1027 (O_1027,N_27138,N_22455);
nand UO_1028 (O_1028,N_24629,N_22294);
xnor UO_1029 (O_1029,N_21079,N_26024);
nand UO_1030 (O_1030,N_24271,N_23011);
or UO_1031 (O_1031,N_28233,N_22095);
xor UO_1032 (O_1032,N_26854,N_20170);
xor UO_1033 (O_1033,N_28136,N_21524);
xnor UO_1034 (O_1034,N_20909,N_22126);
and UO_1035 (O_1035,N_22449,N_25669);
nor UO_1036 (O_1036,N_26342,N_23169);
nor UO_1037 (O_1037,N_21052,N_25970);
and UO_1038 (O_1038,N_26073,N_28158);
nor UO_1039 (O_1039,N_25590,N_26846);
or UO_1040 (O_1040,N_29760,N_29552);
nand UO_1041 (O_1041,N_21807,N_24039);
and UO_1042 (O_1042,N_29270,N_29217);
xor UO_1043 (O_1043,N_23948,N_23470);
and UO_1044 (O_1044,N_27519,N_27796);
and UO_1045 (O_1045,N_22086,N_25698);
nor UO_1046 (O_1046,N_25379,N_28992);
or UO_1047 (O_1047,N_21140,N_20957);
and UO_1048 (O_1048,N_21538,N_21504);
nand UO_1049 (O_1049,N_28230,N_29198);
xor UO_1050 (O_1050,N_22324,N_25691);
and UO_1051 (O_1051,N_20466,N_25439);
or UO_1052 (O_1052,N_23647,N_29490);
xor UO_1053 (O_1053,N_23253,N_21269);
and UO_1054 (O_1054,N_28691,N_29787);
nand UO_1055 (O_1055,N_23107,N_27576);
nor UO_1056 (O_1056,N_20956,N_22649);
xnor UO_1057 (O_1057,N_29165,N_25290);
or UO_1058 (O_1058,N_28976,N_27534);
or UO_1059 (O_1059,N_27107,N_23629);
nor UO_1060 (O_1060,N_22725,N_28482);
nand UO_1061 (O_1061,N_22263,N_28943);
or UO_1062 (O_1062,N_28346,N_25309);
and UO_1063 (O_1063,N_29143,N_23411);
nand UO_1064 (O_1064,N_20577,N_21764);
nand UO_1065 (O_1065,N_22874,N_28381);
and UO_1066 (O_1066,N_23962,N_28400);
and UO_1067 (O_1067,N_23066,N_27262);
and UO_1068 (O_1068,N_28994,N_22058);
nand UO_1069 (O_1069,N_22244,N_26359);
xnor UO_1070 (O_1070,N_27170,N_20073);
nand UO_1071 (O_1071,N_21164,N_23833);
and UO_1072 (O_1072,N_21039,N_28891);
xor UO_1073 (O_1073,N_26899,N_26727);
nor UO_1074 (O_1074,N_28497,N_24516);
nand UO_1075 (O_1075,N_23321,N_29478);
and UO_1076 (O_1076,N_27193,N_22754);
or UO_1077 (O_1077,N_21300,N_27827);
nand UO_1078 (O_1078,N_25619,N_26815);
xor UO_1079 (O_1079,N_20157,N_27396);
or UO_1080 (O_1080,N_23013,N_25862);
and UO_1081 (O_1081,N_28554,N_22403);
nor UO_1082 (O_1082,N_26657,N_29800);
or UO_1083 (O_1083,N_20485,N_26301);
xor UO_1084 (O_1084,N_28541,N_27190);
or UO_1085 (O_1085,N_24859,N_28239);
xnor UO_1086 (O_1086,N_21289,N_26680);
and UO_1087 (O_1087,N_26616,N_21351);
or UO_1088 (O_1088,N_22356,N_23161);
nand UO_1089 (O_1089,N_25560,N_23642);
xor UO_1090 (O_1090,N_29093,N_27832);
nor UO_1091 (O_1091,N_24890,N_28022);
nand UO_1092 (O_1092,N_25537,N_23700);
or UO_1093 (O_1093,N_20299,N_25793);
and UO_1094 (O_1094,N_22321,N_24984);
xnor UO_1095 (O_1095,N_21749,N_21246);
nand UO_1096 (O_1096,N_29285,N_27633);
or UO_1097 (O_1097,N_21950,N_23930);
and UO_1098 (O_1098,N_28115,N_23619);
and UO_1099 (O_1099,N_27680,N_27226);
nand UO_1100 (O_1100,N_25655,N_20192);
xor UO_1101 (O_1101,N_29898,N_28000);
xor UO_1102 (O_1102,N_28327,N_20456);
or UO_1103 (O_1103,N_29945,N_27113);
and UO_1104 (O_1104,N_27331,N_22227);
nor UO_1105 (O_1105,N_24248,N_26558);
xor UO_1106 (O_1106,N_24277,N_24027);
or UO_1107 (O_1107,N_27156,N_21328);
xnor UO_1108 (O_1108,N_26853,N_29412);
nand UO_1109 (O_1109,N_21562,N_23534);
or UO_1110 (O_1110,N_28133,N_21793);
nand UO_1111 (O_1111,N_22622,N_23088);
and UO_1112 (O_1112,N_28721,N_20997);
nand UO_1113 (O_1113,N_27619,N_23001);
and UO_1114 (O_1114,N_23811,N_24059);
xnor UO_1115 (O_1115,N_28033,N_28768);
xnor UO_1116 (O_1116,N_25922,N_26706);
and UO_1117 (O_1117,N_24041,N_21706);
xnor UO_1118 (O_1118,N_26033,N_22631);
or UO_1119 (O_1119,N_27011,N_28256);
xor UO_1120 (O_1120,N_28537,N_21645);
and UO_1121 (O_1121,N_20372,N_23538);
xnor UO_1122 (O_1122,N_27359,N_28390);
nor UO_1123 (O_1123,N_24505,N_27531);
and UO_1124 (O_1124,N_25410,N_22178);
or UO_1125 (O_1125,N_24443,N_29673);
or UO_1126 (O_1126,N_28140,N_25377);
nor UO_1127 (O_1127,N_22946,N_28926);
xnor UO_1128 (O_1128,N_23282,N_21387);
xnor UO_1129 (O_1129,N_22545,N_21327);
nor UO_1130 (O_1130,N_23016,N_29715);
and UO_1131 (O_1131,N_28827,N_25238);
xnor UO_1132 (O_1132,N_29707,N_26364);
nor UO_1133 (O_1133,N_28890,N_29056);
nand UO_1134 (O_1134,N_23491,N_27841);
and UO_1135 (O_1135,N_24846,N_24948);
or UO_1136 (O_1136,N_28738,N_23289);
or UO_1137 (O_1137,N_24567,N_27408);
or UO_1138 (O_1138,N_21650,N_21614);
or UO_1139 (O_1139,N_21261,N_27545);
or UO_1140 (O_1140,N_26845,N_24087);
nand UO_1141 (O_1141,N_25564,N_27589);
nor UO_1142 (O_1142,N_24933,N_25814);
nor UO_1143 (O_1143,N_21366,N_27594);
xor UO_1144 (O_1144,N_24067,N_28208);
nor UO_1145 (O_1145,N_23551,N_23278);
nand UO_1146 (O_1146,N_24514,N_23600);
nand UO_1147 (O_1147,N_26944,N_26488);
and UO_1148 (O_1148,N_21991,N_20127);
xnor UO_1149 (O_1149,N_26740,N_29282);
nand UO_1150 (O_1150,N_23503,N_28357);
or UO_1151 (O_1151,N_29170,N_26796);
xnor UO_1152 (O_1152,N_20666,N_29997);
or UO_1153 (O_1153,N_25479,N_24603);
nor UO_1154 (O_1154,N_24279,N_23064);
nand UO_1155 (O_1155,N_26044,N_27629);
xor UO_1156 (O_1156,N_22547,N_24483);
and UO_1157 (O_1157,N_23361,N_28660);
and UO_1158 (O_1158,N_26979,N_23082);
xor UO_1159 (O_1159,N_20988,N_25676);
and UO_1160 (O_1160,N_23862,N_27924);
nor UO_1161 (O_1161,N_26981,N_25423);
and UO_1162 (O_1162,N_25809,N_28798);
nor UO_1163 (O_1163,N_26711,N_26900);
nand UO_1164 (O_1164,N_27767,N_27489);
nand UO_1165 (O_1165,N_28416,N_25523);
or UO_1166 (O_1166,N_29982,N_21921);
xor UO_1167 (O_1167,N_24939,N_22493);
xnor UO_1168 (O_1168,N_29877,N_24856);
or UO_1169 (O_1169,N_28669,N_21969);
and UO_1170 (O_1170,N_23741,N_22695);
and UO_1171 (O_1171,N_29249,N_28572);
nand UO_1172 (O_1172,N_23720,N_28708);
and UO_1173 (O_1173,N_27603,N_26506);
and UO_1174 (O_1174,N_29016,N_26780);
xnor UO_1175 (O_1175,N_28494,N_21281);
nand UO_1176 (O_1176,N_21447,N_28958);
nor UO_1177 (O_1177,N_27343,N_21571);
or UO_1178 (O_1178,N_29700,N_29730);
nor UO_1179 (O_1179,N_27732,N_25605);
xor UO_1180 (O_1180,N_29476,N_25992);
nand UO_1181 (O_1181,N_22758,N_23104);
or UO_1182 (O_1182,N_29716,N_27925);
nor UO_1183 (O_1183,N_24956,N_26768);
or UO_1184 (O_1184,N_20830,N_28570);
xor UO_1185 (O_1185,N_25674,N_21287);
nor UO_1186 (O_1186,N_24839,N_28150);
nand UO_1187 (O_1187,N_29747,N_25561);
xnor UO_1188 (O_1188,N_27266,N_20531);
xnor UO_1189 (O_1189,N_27224,N_23426);
or UO_1190 (O_1190,N_28406,N_22283);
or UO_1191 (O_1191,N_20037,N_20046);
or UO_1192 (O_1192,N_25135,N_26011);
nor UO_1193 (O_1193,N_28697,N_27310);
and UO_1194 (O_1194,N_24525,N_20236);
nand UO_1195 (O_1195,N_24469,N_22881);
or UO_1196 (O_1196,N_27051,N_24672);
nor UO_1197 (O_1197,N_28182,N_26385);
nor UO_1198 (O_1198,N_29371,N_22854);
or UO_1199 (O_1199,N_27959,N_20935);
or UO_1200 (O_1200,N_26198,N_25285);
nand UO_1201 (O_1201,N_27422,N_25498);
nand UO_1202 (O_1202,N_26149,N_22081);
xor UO_1203 (O_1203,N_23582,N_24326);
nand UO_1204 (O_1204,N_23075,N_29904);
nand UO_1205 (O_1205,N_29695,N_25441);
or UO_1206 (O_1206,N_27931,N_21605);
xor UO_1207 (O_1207,N_24208,N_20006);
xnor UO_1208 (O_1208,N_24290,N_29895);
nor UO_1209 (O_1209,N_24743,N_25722);
and UO_1210 (O_1210,N_26440,N_21715);
and UO_1211 (O_1211,N_25797,N_25531);
nand UO_1212 (O_1212,N_25197,N_26400);
xnor UO_1213 (O_1213,N_27763,N_25988);
xor UO_1214 (O_1214,N_20033,N_29193);
xor UO_1215 (O_1215,N_24821,N_22888);
nand UO_1216 (O_1216,N_20095,N_23448);
or UO_1217 (O_1217,N_29558,N_24526);
or UO_1218 (O_1218,N_27668,N_26139);
nor UO_1219 (O_1219,N_21931,N_24512);
or UO_1220 (O_1220,N_28545,N_27237);
and UO_1221 (O_1221,N_24221,N_23914);
nand UO_1222 (O_1222,N_27106,N_28165);
and UO_1223 (O_1223,N_28187,N_25475);
xor UO_1224 (O_1224,N_23322,N_25695);
or UO_1225 (O_1225,N_25174,N_23777);
and UO_1226 (O_1226,N_22114,N_26223);
and UO_1227 (O_1227,N_27329,N_23157);
or UO_1228 (O_1228,N_20316,N_23083);
or UO_1229 (O_1229,N_27877,N_25904);
nor UO_1230 (O_1230,N_21401,N_29420);
xor UO_1231 (O_1231,N_20850,N_21072);
and UO_1232 (O_1232,N_23427,N_26414);
nor UO_1233 (O_1233,N_22066,N_28459);
or UO_1234 (O_1234,N_25579,N_24728);
nor UO_1235 (O_1235,N_24817,N_20967);
nand UO_1236 (O_1236,N_26867,N_22220);
and UO_1237 (O_1237,N_29429,N_21494);
nor UO_1238 (O_1238,N_28902,N_28531);
xnor UO_1239 (O_1239,N_25668,N_20028);
or UO_1240 (O_1240,N_29672,N_27994);
and UO_1241 (O_1241,N_25966,N_20807);
and UO_1242 (O_1242,N_20703,N_29328);
and UO_1243 (O_1243,N_22277,N_27648);
nand UO_1244 (O_1244,N_22724,N_27549);
nand UO_1245 (O_1245,N_28656,N_27814);
nand UO_1246 (O_1246,N_29565,N_27987);
or UO_1247 (O_1247,N_21042,N_29970);
nand UO_1248 (O_1248,N_29015,N_25358);
and UO_1249 (O_1249,N_26629,N_28802);
nor UO_1250 (O_1250,N_25283,N_26598);
nand UO_1251 (O_1251,N_23913,N_24044);
or UO_1252 (O_1252,N_26171,N_29377);
xnor UO_1253 (O_1253,N_20884,N_27233);
or UO_1254 (O_1254,N_27802,N_26542);
and UO_1255 (O_1255,N_26348,N_29477);
and UO_1256 (O_1256,N_29764,N_27115);
xnor UO_1257 (O_1257,N_28806,N_23126);
nor UO_1258 (O_1258,N_24190,N_22389);
and UO_1259 (O_1259,N_23897,N_28266);
nor UO_1260 (O_1260,N_22183,N_21489);
and UO_1261 (O_1261,N_29491,N_29798);
xnor UO_1262 (O_1262,N_27747,N_21577);
xor UO_1263 (O_1263,N_25184,N_25735);
nand UO_1264 (O_1264,N_26295,N_29078);
nor UO_1265 (O_1265,N_26949,N_25859);
or UO_1266 (O_1266,N_29775,N_22030);
xor UO_1267 (O_1267,N_27340,N_23170);
nor UO_1268 (O_1268,N_21770,N_27257);
nor UO_1269 (O_1269,N_28948,N_29397);
nor UO_1270 (O_1270,N_24057,N_23506);
or UO_1271 (O_1271,N_25807,N_23492);
xor UO_1272 (O_1272,N_26355,N_23776);
nor UO_1273 (O_1273,N_22624,N_25846);
and UO_1274 (O_1274,N_21532,N_20332);
nand UO_1275 (O_1275,N_20150,N_26622);
or UO_1276 (O_1276,N_23468,N_25160);
nand UO_1277 (O_1277,N_21360,N_24958);
and UO_1278 (O_1278,N_23187,N_24060);
nand UO_1279 (O_1279,N_29714,N_23789);
and UO_1280 (O_1280,N_27344,N_25789);
and UO_1281 (O_1281,N_20934,N_25758);
xor UO_1282 (O_1282,N_27969,N_22773);
nor UO_1283 (O_1283,N_22769,N_24402);
or UO_1284 (O_1284,N_28364,N_28463);
xnor UO_1285 (O_1285,N_24355,N_26427);
nand UO_1286 (O_1286,N_27626,N_25440);
and UO_1287 (O_1287,N_21212,N_28251);
nor UO_1288 (O_1288,N_22574,N_22536);
or UO_1289 (O_1289,N_20672,N_29085);
and UO_1290 (O_1290,N_24919,N_23658);
or UO_1291 (O_1291,N_21224,N_27032);
and UO_1292 (O_1292,N_21481,N_29900);
nand UO_1293 (O_1293,N_23683,N_21887);
nand UO_1294 (O_1294,N_26804,N_29480);
xnor UO_1295 (O_1295,N_25573,N_27462);
nor UO_1296 (O_1296,N_24147,N_23760);
nand UO_1297 (O_1297,N_23583,N_22678);
nand UO_1298 (O_1298,N_25790,N_23929);
nor UO_1299 (O_1299,N_24789,N_29847);
nand UO_1300 (O_1300,N_28496,N_22688);
and UO_1301 (O_1301,N_23260,N_25608);
nor UO_1302 (O_1302,N_29965,N_29645);
nand UO_1303 (O_1303,N_22342,N_26043);
nor UO_1304 (O_1304,N_28706,N_22565);
xor UO_1305 (O_1305,N_25929,N_26470);
or UO_1306 (O_1306,N_29830,N_28306);
and UO_1307 (O_1307,N_21978,N_28688);
nor UO_1308 (O_1308,N_23295,N_28443);
or UO_1309 (O_1309,N_21158,N_21817);
nor UO_1310 (O_1310,N_26451,N_21794);
nand UO_1311 (O_1311,N_21251,N_24909);
xor UO_1312 (O_1312,N_26031,N_26533);
xor UO_1313 (O_1313,N_21306,N_20323);
nor UO_1314 (O_1314,N_28215,N_24840);
or UO_1315 (O_1315,N_28859,N_24145);
xor UO_1316 (O_1316,N_21066,N_23367);
or UO_1317 (O_1317,N_29450,N_24811);
and UO_1318 (O_1318,N_24407,N_22271);
and UO_1319 (O_1319,N_28509,N_28366);
xnor UO_1320 (O_1320,N_20297,N_25241);
xnor UO_1321 (O_1321,N_27571,N_26760);
or UO_1322 (O_1322,N_22039,N_23430);
and UO_1323 (O_1323,N_27023,N_29789);
or UO_1324 (O_1324,N_20300,N_27092);
or UO_1325 (O_1325,N_25869,N_26458);
or UO_1326 (O_1326,N_25958,N_22518);
nand UO_1327 (O_1327,N_28876,N_25653);
and UO_1328 (O_1328,N_22077,N_29598);
nor UO_1329 (O_1329,N_29762,N_24081);
nor UO_1330 (O_1330,N_24014,N_21264);
nor UO_1331 (O_1331,N_25327,N_27173);
nand UO_1332 (O_1332,N_23262,N_26569);
nor UO_1333 (O_1333,N_21629,N_29845);
xor UO_1334 (O_1334,N_23545,N_20890);
or UO_1335 (O_1335,N_27748,N_22184);
nand UO_1336 (O_1336,N_27094,N_23826);
nor UO_1337 (O_1337,N_21994,N_24519);
or UO_1338 (O_1338,N_20354,N_23820);
nand UO_1339 (O_1339,N_23017,N_20937);
nand UO_1340 (O_1340,N_21843,N_23609);
nor UO_1341 (O_1341,N_23481,N_21270);
or UO_1342 (O_1342,N_20360,N_29865);
and UO_1343 (O_1343,N_25496,N_24159);
xnor UO_1344 (O_1344,N_22428,N_23472);
xnor UO_1345 (O_1345,N_25148,N_23231);
and UO_1346 (O_1346,N_24318,N_24378);
nor UO_1347 (O_1347,N_21196,N_21672);
nor UO_1348 (O_1348,N_20424,N_22042);
and UO_1349 (O_1349,N_23884,N_26305);
nor UO_1350 (O_1350,N_20740,N_26307);
nand UO_1351 (O_1351,N_26306,N_28032);
nand UO_1352 (O_1352,N_28467,N_26619);
or UO_1353 (O_1353,N_20219,N_20581);
xnor UO_1354 (O_1354,N_20042,N_27909);
nor UO_1355 (O_1355,N_29196,N_26187);
nor UO_1356 (O_1356,N_25159,N_24959);
nor UO_1357 (O_1357,N_22979,N_26493);
nor UO_1358 (O_1358,N_29115,N_26847);
and UO_1359 (O_1359,N_21441,N_28632);
xnor UO_1360 (O_1360,N_26373,N_27248);
and UO_1361 (O_1361,N_20892,N_24084);
xor UO_1362 (O_1362,N_29131,N_23203);
xor UO_1363 (O_1363,N_26155,N_27005);
and UO_1364 (O_1364,N_27222,N_25331);
or UO_1365 (O_1365,N_23901,N_23727);
or UO_1366 (O_1366,N_29492,N_23477);
or UO_1367 (O_1367,N_20601,N_28378);
nor UO_1368 (O_1368,N_28568,N_21445);
nor UO_1369 (O_1369,N_23155,N_27951);
or UO_1370 (O_1370,N_28050,N_28272);
nand UO_1371 (O_1371,N_26032,N_22575);
xnor UO_1372 (O_1372,N_23855,N_21675);
nand UO_1373 (O_1373,N_24286,N_25221);
xor UO_1374 (O_1374,N_27774,N_28229);
xor UO_1375 (O_1375,N_24446,N_28808);
nand UO_1376 (O_1376,N_27040,N_25972);
nand UO_1377 (O_1377,N_25903,N_28161);
xnor UO_1378 (O_1378,N_25398,N_24524);
nand UO_1379 (O_1379,N_29057,N_29681);
xnor UO_1380 (O_1380,N_27333,N_22894);
or UO_1381 (O_1381,N_29045,N_27509);
xor UO_1382 (O_1382,N_27638,N_20555);
nor UO_1383 (O_1383,N_23556,N_27978);
or UO_1384 (O_1384,N_21188,N_20966);
or UO_1385 (O_1385,N_20239,N_20309);
or UO_1386 (O_1386,N_22022,N_27353);
nand UO_1387 (O_1387,N_20527,N_25010);
nor UO_1388 (O_1388,N_25801,N_20342);
nand UO_1389 (O_1389,N_24547,N_26921);
and UO_1390 (O_1390,N_23542,N_25150);
or UO_1391 (O_1391,N_20114,N_20676);
nor UO_1392 (O_1392,N_28635,N_20605);
nand UO_1393 (O_1393,N_27824,N_27205);
nand UO_1394 (O_1394,N_20748,N_28804);
xnor UO_1395 (O_1395,N_28810,N_21819);
nor UO_1396 (O_1396,N_24795,N_29030);
xor UO_1397 (O_1397,N_21255,N_22109);
and UO_1398 (O_1398,N_23175,N_23378);
nand UO_1399 (O_1399,N_24468,N_22859);
and UO_1400 (O_1400,N_21945,N_26638);
nand UO_1401 (O_1401,N_23065,N_27861);
and UO_1402 (O_1402,N_26252,N_29324);
nor UO_1403 (O_1403,N_28322,N_23831);
and UO_1404 (O_1404,N_27685,N_25182);
nand UO_1405 (O_1405,N_22460,N_21830);
nand UO_1406 (O_1406,N_29669,N_25951);
nor UO_1407 (O_1407,N_20215,N_29615);
and UO_1408 (O_1408,N_28227,N_23027);
and UO_1409 (O_1409,N_23852,N_20692);
or UO_1410 (O_1410,N_29495,N_23513);
and UO_1411 (O_1411,N_24554,N_22007);
or UO_1412 (O_1412,N_25009,N_21813);
and UO_1413 (O_1413,N_23436,N_24176);
nor UO_1414 (O_1414,N_28213,N_20379);
nor UO_1415 (O_1415,N_21006,N_25654);
nand UO_1416 (O_1416,N_20806,N_29737);
xor UO_1417 (O_1417,N_23756,N_28105);
and UO_1418 (O_1418,N_22749,N_25092);
nand UO_1419 (O_1419,N_24080,N_21143);
and UO_1420 (O_1420,N_27977,N_20515);
nand UO_1421 (O_1421,N_21132,N_29161);
nand UO_1422 (O_1422,N_23940,N_24507);
nor UO_1423 (O_1423,N_29966,N_28273);
or UO_1424 (O_1424,N_28166,N_27540);
nand UO_1425 (O_1425,N_23562,N_27862);
nor UO_1426 (O_1426,N_22217,N_27906);
or UO_1427 (O_1427,N_26691,N_26724);
or UO_1428 (O_1428,N_27456,N_22381);
and UO_1429 (O_1429,N_24750,N_26875);
nor UO_1430 (O_1430,N_20739,N_22502);
nor UO_1431 (O_1431,N_29933,N_29888);
nor UO_1432 (O_1432,N_28424,N_20925);
nor UO_1433 (O_1433,N_22024,N_29002);
and UO_1434 (O_1434,N_20384,N_25378);
xor UO_1435 (O_1435,N_24333,N_29783);
nand UO_1436 (O_1436,N_22196,N_24950);
nand UO_1437 (O_1437,N_27860,N_27585);
nand UO_1438 (O_1438,N_24412,N_28503);
xor UO_1439 (O_1439,N_24592,N_24921);
nor UO_1440 (O_1440,N_22033,N_25553);
nor UO_1441 (O_1441,N_29162,N_23631);
nor UO_1442 (O_1442,N_22875,N_24390);
or UO_1443 (O_1443,N_23097,N_22607);
or UO_1444 (O_1444,N_23188,N_29430);
xor UO_1445 (O_1445,N_26612,N_21802);
xnor UO_1446 (O_1446,N_28741,N_26662);
or UO_1447 (O_1447,N_24020,N_24801);
xnor UO_1448 (O_1448,N_20089,N_27221);
and UO_1449 (O_1449,N_23338,N_20407);
xor UO_1450 (O_1450,N_27721,N_29256);
nor UO_1451 (O_1451,N_27654,N_28945);
nand UO_1452 (O_1452,N_20160,N_26358);
xnor UO_1453 (O_1453,N_25522,N_23383);
nand UO_1454 (O_1454,N_28936,N_26001);
nand UO_1455 (O_1455,N_21176,N_28865);
nand UO_1456 (O_1456,N_28268,N_26585);
and UO_1457 (O_1457,N_28838,N_24977);
nand UO_1458 (O_1458,N_26254,N_26567);
and UO_1459 (O_1459,N_20346,N_21070);
or UO_1460 (O_1460,N_27631,N_23652);
nand UO_1461 (O_1461,N_25117,N_22182);
and UO_1462 (O_1462,N_21339,N_24790);
nand UO_1463 (O_1463,N_21646,N_24745);
nand UO_1464 (O_1464,N_28004,N_26821);
nand UO_1465 (O_1465,N_26345,N_21086);
nand UO_1466 (O_1466,N_21691,N_25300);
nand UO_1467 (O_1467,N_24535,N_29129);
xnor UO_1468 (O_1468,N_20762,N_27236);
and UO_1469 (O_1469,N_21546,N_21283);
nor UO_1470 (O_1470,N_22517,N_26025);
and UO_1471 (O_1471,N_24431,N_28344);
xor UO_1472 (O_1472,N_29732,N_23617);
or UO_1473 (O_1473,N_29070,N_20470);
and UO_1474 (O_1474,N_24444,N_22349);
and UO_1475 (O_1475,N_22252,N_24302);
xor UO_1476 (O_1476,N_29548,N_29389);
and UO_1477 (O_1477,N_22957,N_22031);
or UO_1478 (O_1478,N_25029,N_20070);
nor UO_1479 (O_1479,N_21020,N_29554);
or UO_1480 (O_1480,N_24808,N_27270);
or UO_1481 (O_1481,N_28583,N_22801);
or UO_1482 (O_1482,N_20140,N_26253);
xnor UO_1483 (O_1483,N_26182,N_23303);
xnor UO_1484 (O_1484,N_20826,N_22423);
nand UO_1485 (O_1485,N_21185,N_24857);
or UO_1486 (O_1486,N_25291,N_23563);
or UO_1487 (O_1487,N_25941,N_22558);
or UO_1488 (O_1488,N_23085,N_21060);
and UO_1489 (O_1489,N_27048,N_21108);
nand UO_1490 (O_1490,N_20735,N_25161);
and UO_1491 (O_1491,N_24386,N_25326);
and UO_1492 (O_1492,N_22650,N_25645);
xor UO_1493 (O_1493,N_26757,N_29613);
or UO_1494 (O_1494,N_21348,N_24722);
xor UO_1495 (O_1495,N_28615,N_25599);
nand UO_1496 (O_1496,N_29010,N_20132);
nor UO_1497 (O_1497,N_25493,N_24404);
and UO_1498 (O_1498,N_25585,N_22427);
or UO_1499 (O_1499,N_26159,N_22384);
and UO_1500 (O_1500,N_23704,N_21796);
nor UO_1501 (O_1501,N_22084,N_26271);
or UO_1502 (O_1502,N_26170,N_23961);
nor UO_1503 (O_1503,N_23239,N_21350);
and UO_1504 (O_1504,N_22504,N_22017);
xor UO_1505 (O_1505,N_24269,N_22076);
and UO_1506 (O_1506,N_21096,N_28285);
xor UO_1507 (O_1507,N_22169,N_22571);
xnor UO_1508 (O_1508,N_20624,N_21690);
or UO_1509 (O_1509,N_21322,N_20462);
and UO_1510 (O_1510,N_21123,N_28368);
nor UO_1511 (O_1511,N_27768,N_21167);
or UO_1512 (O_1512,N_24036,N_20345);
xor UO_1513 (O_1513,N_28514,N_24749);
or UO_1514 (O_1514,N_28398,N_20318);
or UO_1515 (O_1515,N_22928,N_22065);
nor UO_1516 (O_1516,N_24158,N_21092);
or UO_1517 (O_1517,N_28216,N_24691);
nand UO_1518 (O_1518,N_21169,N_28875);
and UO_1519 (O_1519,N_23077,N_29350);
and UO_1520 (O_1520,N_26023,N_29976);
and UO_1521 (O_1521,N_26879,N_26664);
or UO_1522 (O_1522,N_27488,N_24099);
nor UO_1523 (O_1523,N_29561,N_24052);
nor UO_1524 (O_1524,N_24005,N_22829);
nand UO_1525 (O_1525,N_25396,N_24481);
nand UO_1526 (O_1526,N_25417,N_23293);
xor UO_1527 (O_1527,N_25096,N_23770);
and UO_1528 (O_1528,N_20667,N_23151);
and UO_1529 (O_1529,N_28023,N_26997);
nor UO_1530 (O_1530,N_26144,N_27777);
or UO_1531 (O_1531,N_20121,N_27426);
nor UO_1532 (O_1532,N_21062,N_25449);
nor UO_1533 (O_1533,N_22148,N_26035);
or UO_1534 (O_1534,N_27880,N_22533);
nor UO_1535 (O_1535,N_23132,N_25317);
and UO_1536 (O_1536,N_20305,N_23235);
or UO_1537 (O_1537,N_26608,N_28549);
and UO_1538 (O_1538,N_28892,N_27267);
nor UO_1539 (O_1539,N_28648,N_20880);
nor UO_1540 (O_1540,N_24097,N_27072);
nand UO_1541 (O_1541,N_26962,N_28598);
nand UO_1542 (O_1542,N_23019,N_24478);
xor UO_1543 (O_1543,N_22014,N_28634);
or UO_1544 (O_1544,N_27578,N_21497);
and UO_1545 (O_1545,N_26856,N_22075);
nor UO_1546 (O_1546,N_25185,N_28152);
or UO_1547 (O_1547,N_25451,N_23377);
and UO_1548 (O_1548,N_25818,N_22162);
nand UO_1549 (O_1549,N_21590,N_23055);
and UO_1550 (O_1550,N_25100,N_25129);
and UO_1551 (O_1551,N_25516,N_22437);
and UO_1552 (O_1552,N_24604,N_23900);
xnor UO_1553 (O_1553,N_22748,N_25963);
nor UO_1554 (O_1554,N_24532,N_27830);
xnor UO_1555 (O_1555,N_22654,N_26829);
or UO_1556 (O_1556,N_23774,N_28613);
xor UO_1557 (O_1557,N_24700,N_25689);
xor UO_1558 (O_1558,N_27090,N_24222);
or UO_1559 (O_1559,N_28442,N_21100);
or UO_1560 (O_1560,N_22898,N_26826);
and UO_1561 (O_1561,N_20484,N_27988);
nor UO_1562 (O_1562,N_25058,N_22212);
or UO_1563 (O_1563,N_25313,N_25630);
or UO_1564 (O_1564,N_25555,N_23905);
and UO_1565 (O_1565,N_21223,N_27640);
xor UO_1566 (O_1566,N_23058,N_27957);
nor UO_1567 (O_1567,N_26604,N_20136);
and UO_1568 (O_1568,N_20255,N_23070);
xor UO_1569 (O_1569,N_29233,N_21170);
or UO_1570 (O_1570,N_28125,N_25373);
or UO_1571 (O_1571,N_22368,N_25408);
and UO_1572 (O_1572,N_27406,N_24733);
nor UO_1573 (O_1573,N_23286,N_23304);
xnor UO_1574 (O_1574,N_25369,N_29604);
and UO_1575 (O_1575,N_29079,N_26473);
and UO_1576 (O_1576,N_20810,N_26087);
and UO_1577 (O_1577,N_24137,N_28940);
or UO_1578 (O_1578,N_29560,N_27869);
xor UO_1579 (O_1579,N_26868,N_23768);
or UO_1580 (O_1580,N_24146,N_20678);
nand UO_1581 (O_1581,N_22292,N_25464);
and UO_1582 (O_1582,N_23692,N_28647);
nor UO_1583 (O_1583,N_24803,N_28031);
and UO_1584 (O_1584,N_24065,N_26181);
or UO_1585 (O_1585,N_25365,N_27798);
xor UO_1586 (O_1586,N_27212,N_20616);
nor UO_1587 (O_1587,N_27625,N_29167);
or UO_1588 (O_1588,N_28611,N_28157);
nor UO_1589 (O_1589,N_21952,N_28676);
xor UO_1590 (O_1590,N_28974,N_25536);
and UO_1591 (O_1591,N_24586,N_25214);
xor UO_1592 (O_1592,N_20870,N_21826);
xor UO_1593 (O_1593,N_28488,N_27126);
xnor UO_1594 (O_1594,N_27078,N_29774);
nor UO_1595 (O_1595,N_28298,N_25294);
or UO_1596 (O_1596,N_27542,N_21080);
xnor UO_1597 (O_1597,N_28534,N_27230);
nand UO_1598 (O_1598,N_28925,N_24951);
nor UO_1599 (O_1599,N_21320,N_21486);
xnor UO_1600 (O_1600,N_24339,N_26234);
nand UO_1601 (O_1601,N_20679,N_23714);
or UO_1602 (O_1602,N_28410,N_29628);
xnor UO_1603 (O_1603,N_28199,N_22421);
and UO_1604 (O_1604,N_20090,N_28027);
nand UO_1605 (O_1605,N_20343,N_22620);
xor UO_1606 (O_1606,N_28518,N_20455);
nand UO_1607 (O_1607,N_25715,N_27974);
nand UO_1608 (O_1608,N_25178,N_20534);
xnor UO_1609 (O_1609,N_24366,N_23922);
nor UO_1610 (O_1610,N_22997,N_28882);
xor UO_1611 (O_1611,N_29327,N_21598);
nor UO_1612 (O_1612,N_29958,N_22918);
nor UO_1613 (O_1613,N_24210,N_25497);
nand UO_1614 (O_1614,N_26709,N_22454);
nand UO_1615 (O_1615,N_27742,N_20328);
and UO_1616 (O_1616,N_27460,N_22131);
nand UO_1617 (O_1617,N_25665,N_23496);
xnor UO_1618 (O_1618,N_26219,N_27562);
nor UO_1619 (O_1619,N_23570,N_21109);
and UO_1620 (O_1620,N_26966,N_26713);
nor UO_1621 (O_1621,N_23571,N_26439);
nand UO_1622 (O_1622,N_23530,N_22714);
nand UO_1623 (O_1623,N_26396,N_24766);
or UO_1624 (O_1624,N_29831,N_22580);
nand UO_1625 (O_1625,N_28461,N_24635);
and UO_1626 (O_1626,N_25957,N_23703);
nor UO_1627 (O_1627,N_29622,N_27069);
nor UO_1628 (O_1628,N_29824,N_28458);
or UO_1629 (O_1629,N_25604,N_24679);
or UO_1630 (O_1630,N_26054,N_25746);
xnor UO_1631 (O_1631,N_20708,N_27314);
and UO_1632 (O_1632,N_23992,N_26310);
and UO_1633 (O_1633,N_28777,N_25986);
xor UO_1634 (O_1634,N_23575,N_29316);
nand UO_1635 (O_1635,N_22921,N_26460);
xor UO_1636 (O_1636,N_22549,N_23039);
nor UO_1637 (O_1637,N_20256,N_23327);
or UO_1638 (O_1638,N_29533,N_20043);
or UO_1639 (O_1639,N_26209,N_20901);
nand UO_1640 (O_1640,N_24095,N_25374);
and UO_1641 (O_1641,N_27478,N_29026);
or UO_1642 (O_1642,N_25612,N_27799);
xor UO_1643 (O_1643,N_27183,N_25670);
and UO_1644 (O_1644,N_28369,N_27500);
and UO_1645 (O_1645,N_27867,N_22002);
or UO_1646 (O_1646,N_24741,N_23299);
nor UO_1647 (O_1647,N_20053,N_21514);
nand UO_1648 (O_1648,N_22180,N_21832);
xor UO_1649 (O_1649,N_24659,N_23081);
and UO_1650 (O_1650,N_21228,N_23866);
and UO_1651 (O_1651,N_27466,N_23541);
nand UO_1652 (O_1652,N_24427,N_23221);
xor UO_1653 (O_1653,N_26242,N_24636);
nor UO_1654 (O_1654,N_28671,N_24495);
nor UO_1655 (O_1655,N_23612,N_23191);
xnor UO_1656 (O_1656,N_20282,N_24702);
and UO_1657 (O_1657,N_26179,N_22797);
nor UO_1658 (O_1658,N_29254,N_20566);
or UO_1659 (O_1659,N_22309,N_28665);
or UO_1660 (O_1660,N_27019,N_20650);
nand UO_1661 (O_1661,N_27366,N_23347);
and UO_1662 (O_1662,N_27014,N_25768);
and UO_1663 (O_1663,N_29269,N_20237);
or UO_1664 (O_1664,N_25684,N_21812);
nand UO_1665 (O_1665,N_21150,N_29048);
or UO_1666 (O_1666,N_21453,N_22335);
nor UO_1667 (O_1667,N_26579,N_26943);
nor UO_1668 (O_1668,N_20373,N_29861);
xor UO_1669 (O_1669,N_22200,N_21886);
and UO_1670 (O_1670,N_26081,N_27141);
and UO_1671 (O_1671,N_21338,N_29753);
nand UO_1672 (O_1672,N_23091,N_28659);
xnor UO_1673 (O_1673,N_21871,N_26742);
or UO_1674 (O_1674,N_22762,N_22032);
nand UO_1675 (O_1675,N_23878,N_23510);
nand UO_1676 (O_1676,N_20034,N_25231);
and UO_1677 (O_1677,N_21277,N_26620);
and UO_1678 (O_1678,N_29585,N_29893);
and UO_1679 (O_1679,N_23166,N_29183);
nand UO_1680 (O_1680,N_23591,N_22969);
and UO_1681 (O_1681,N_24372,N_20627);
xor UO_1682 (O_1682,N_27702,N_27804);
and UO_1683 (O_1683,N_25899,N_27960);
xor UO_1684 (O_1684,N_27104,N_21162);
nand UO_1685 (O_1685,N_21827,N_26266);
nor UO_1686 (O_1686,N_28901,N_24809);
or UO_1687 (O_1687,N_27434,N_22967);
and UO_1688 (O_1688,N_26807,N_21359);
xor UO_1689 (O_1689,N_28009,N_26753);
nor UO_1690 (O_1690,N_24841,N_27826);
nand UO_1691 (O_1691,N_21177,N_26498);
and UO_1692 (O_1692,N_24557,N_27782);
xor UO_1693 (O_1693,N_29432,N_29073);
xor UO_1694 (O_1694,N_29582,N_22345);
and UO_1695 (O_1695,N_25128,N_26244);
nand UO_1696 (O_1696,N_20614,N_29231);
or UO_1697 (O_1697,N_20087,N_29418);
or UO_1698 (O_1698,N_22656,N_22752);
and UO_1699 (O_1699,N_26382,N_29574);
nor UO_1700 (O_1700,N_25356,N_24169);
nand UO_1701 (O_1701,N_23488,N_23006);
and UO_1702 (O_1702,N_28566,N_25099);
and UO_1703 (O_1703,N_23440,N_29080);
nor UO_1704 (O_1704,N_22037,N_29633);
and UO_1705 (O_1705,N_28725,N_27483);
xnor UO_1706 (O_1706,N_26476,N_20576);
or UO_1707 (O_1707,N_24180,N_28340);
and UO_1708 (O_1708,N_27103,N_25948);
nor UO_1709 (O_1709,N_20265,N_29206);
xor UO_1710 (O_1710,N_22995,N_29127);
nand UO_1711 (O_1711,N_21890,N_24805);
nand UO_1712 (O_1712,N_27260,N_28830);
nand UO_1713 (O_1713,N_26479,N_29194);
and UO_1714 (O_1714,N_26918,N_24110);
nor UO_1715 (O_1715,N_24791,N_25047);
xnor UO_1716 (O_1716,N_21686,N_23489);
and UO_1717 (O_1717,N_29686,N_23978);
xor UO_1718 (O_1718,N_23872,N_26229);
or UO_1719 (O_1719,N_24701,N_20030);
nor UO_1720 (O_1720,N_20024,N_25947);
or UO_1721 (O_1721,N_26413,N_29184);
nand UO_1722 (O_1722,N_25044,N_27838);
and UO_1723 (O_1723,N_22060,N_20989);
xor UO_1724 (O_1724,N_29625,N_29650);
nand UO_1725 (O_1725,N_24800,N_26820);
or UO_1726 (O_1726,N_22665,N_20928);
nand UO_1727 (O_1727,N_20659,N_26431);
nor UO_1728 (O_1728,N_25975,N_29596);
nor UO_1729 (O_1729,N_25355,N_27122);
nor UO_1730 (O_1730,N_28238,N_25731);
xor UO_1731 (O_1731,N_20131,N_27933);
nor UO_1732 (O_1732,N_22572,N_27303);
nor UO_1733 (O_1733,N_22707,N_21055);
nand UO_1734 (O_1734,N_21519,N_22242);
or UO_1735 (O_1735,N_23113,N_27999);
nand UO_1736 (O_1736,N_29158,N_23087);
or UO_1737 (O_1737,N_27209,N_25473);
and UO_1738 (O_1738,N_27146,N_28920);
or UO_1739 (O_1739,N_25217,N_20745);
or UO_1740 (O_1740,N_22826,N_27228);
nand UO_1741 (O_1741,N_23691,N_22593);
or UO_1742 (O_1742,N_21475,N_29375);
xnor UO_1743 (O_1743,N_29664,N_22689);
nor UO_1744 (O_1744,N_25407,N_28784);
nand UO_1745 (O_1745,N_29338,N_24417);
nand UO_1746 (O_1746,N_28831,N_24641);
and UO_1747 (O_1747,N_21823,N_27795);
nor UO_1748 (O_1748,N_26828,N_29666);
xor UO_1749 (O_1749,N_24016,N_23415);
nor UO_1750 (O_1750,N_25017,N_27661);
nor UO_1751 (O_1751,N_24646,N_27395);
nor UO_1752 (O_1752,N_24396,N_26487);
or UO_1753 (O_1753,N_25167,N_25195);
or UO_1754 (O_1754,N_22177,N_24595);
xnor UO_1755 (O_1755,N_29225,N_25977);
nor UO_1756 (O_1756,N_21500,N_22940);
and UO_1757 (O_1757,N_28061,N_22870);
or UO_1758 (O_1758,N_20985,N_28593);
nor UO_1759 (O_1759,N_22857,N_21754);
or UO_1760 (O_1760,N_29549,N_20609);
nand UO_1761 (O_1761,N_25762,N_28446);
xnor UO_1762 (O_1762,N_28743,N_20795);
nor UO_1763 (O_1763,N_22041,N_28814);
or UO_1764 (O_1764,N_27160,N_27229);
or UO_1765 (O_1765,N_27444,N_27794);
nand UO_1766 (O_1766,N_20001,N_26041);
nand UO_1767 (O_1767,N_26800,N_26197);
or UO_1768 (O_1768,N_23702,N_26491);
or UO_1769 (O_1769,N_20682,N_25699);
and UO_1770 (O_1770,N_20920,N_29168);
and UO_1771 (O_1771,N_28552,N_21543);
or UO_1772 (O_1772,N_28121,N_24764);
xor UO_1773 (O_1773,N_22697,N_27737);
nand UO_1774 (O_1774,N_26521,N_25517);
nor UO_1775 (O_1775,N_29096,N_27681);
xnor UO_1776 (O_1776,N_20923,N_20303);
or UO_1777 (O_1777,N_29602,N_29736);
nand UO_1778 (O_1778,N_21731,N_25456);
nor UO_1779 (O_1779,N_25366,N_26933);
nand UO_1780 (O_1780,N_24266,N_23975);
nor UO_1781 (O_1781,N_21046,N_22268);
nor UO_1782 (O_1782,N_21958,N_29434);
or UO_1783 (O_1783,N_29601,N_25495);
or UO_1784 (O_1784,N_22047,N_28619);
or UO_1785 (O_1785,N_26045,N_21839);
xnor UO_1786 (O_1786,N_24761,N_28498);
xor UO_1787 (O_1787,N_23098,N_27472);
nor UO_1788 (O_1788,N_24301,N_28845);
nor UO_1789 (O_1789,N_24596,N_27726);
nor UO_1790 (O_1790,N_20522,N_21091);
or UO_1791 (O_1791,N_29118,N_20704);
or UO_1792 (O_1792,N_23501,N_24450);
nand UO_1793 (O_1793,N_22406,N_23040);
xor UO_1794 (O_1794,N_22751,N_22879);
or UO_1795 (O_1795,N_21778,N_23117);
and UO_1796 (O_1796,N_23816,N_26877);
and UO_1797 (O_1797,N_25589,N_24692);
nor UO_1798 (O_1798,N_24042,N_27201);
xnor UO_1799 (O_1799,N_20451,N_21704);
or UO_1800 (O_1800,N_28714,N_29464);
or UO_1801 (O_1801,N_24996,N_27875);
nor UO_1802 (O_1802,N_26500,N_27634);
or UO_1803 (O_1803,N_28036,N_20096);
nor UO_1804 (O_1804,N_26744,N_25032);
nor UO_1805 (O_1805,N_23931,N_21569);
nor UO_1806 (O_1806,N_20750,N_21341);
xnor UO_1807 (O_1807,N_25406,N_22334);
nor UO_1808 (O_1808,N_25821,N_20809);
and UO_1809 (O_1809,N_20266,N_27720);
xnor UO_1810 (O_1810,N_22366,N_29157);
nor UO_1811 (O_1811,N_27966,N_24342);
nand UO_1812 (O_1812,N_29372,N_22078);
xor UO_1813 (O_1813,N_25437,N_20507);
xnor UO_1814 (O_1814,N_28284,N_23197);
nor UO_1815 (O_1815,N_26914,N_29279);
or UO_1816 (O_1816,N_29494,N_23848);
and UO_1817 (O_1817,N_25681,N_21090);
or UO_1818 (O_1818,N_27525,N_27740);
xor UO_1819 (O_1819,N_23186,N_26588);
nor UO_1820 (O_1820,N_28913,N_24178);
and UO_1821 (O_1821,N_25526,N_24332);
or UO_1822 (O_1822,N_21282,N_20757);
and UO_1823 (O_1823,N_24373,N_25018);
or UO_1824 (O_1824,N_20796,N_28342);
and UO_1825 (O_1825,N_21364,N_21211);
xnor UO_1826 (O_1826,N_24823,N_29454);
xnor UO_1827 (O_1827,N_26407,N_20064);
and UO_1828 (O_1828,N_21462,N_21997);
nand UO_1829 (O_1829,N_23988,N_23564);
or UO_1830 (O_1830,N_22023,N_28590);
xor UO_1831 (O_1831,N_29623,N_20415);
nand UO_1832 (O_1832,N_22376,N_20138);
nand UO_1833 (O_1833,N_29069,N_21421);
and UO_1834 (O_1834,N_29639,N_23640);
nand UO_1835 (O_1835,N_21783,N_22611);
nor UO_1836 (O_1836,N_25729,N_24807);
nand UO_1837 (O_1837,N_25061,N_22788);
nor UO_1838 (O_1838,N_25426,N_28650);
nand UO_1839 (O_1839,N_25518,N_28809);
or UO_1840 (O_1840,N_28335,N_20756);
or UO_1841 (O_1841,N_20434,N_24008);
nand UO_1842 (O_1842,N_20261,N_23199);
or UO_1843 (O_1843,N_24089,N_25617);
xor UO_1844 (O_1844,N_28868,N_24969);
nand UO_1845 (O_1845,N_22844,N_28923);
or UO_1846 (O_1846,N_27256,N_21863);
and UO_1847 (O_1847,N_21434,N_20397);
or UO_1848 (O_1848,N_28908,N_20553);
and UO_1849 (O_1849,N_28779,N_21716);
nand UO_1850 (O_1850,N_22690,N_28176);
or UO_1851 (O_1851,N_22528,N_22510);
or UO_1852 (O_1852,N_24023,N_21286);
or UO_1853 (O_1853,N_22336,N_20911);
and UO_1854 (O_1854,N_22542,N_29134);
xnor UO_1855 (O_1855,N_23484,N_28986);
xnor UO_1856 (O_1856,N_27569,N_29624);
nand UO_1857 (O_1857,N_28425,N_21772);
nor UO_1858 (O_1858,N_22029,N_26190);
nand UO_1859 (O_1859,N_26518,N_21677);
or UO_1860 (O_1860,N_29661,N_28988);
and UO_1861 (O_1861,N_23101,N_24236);
xnor UO_1862 (O_1862,N_20193,N_20654);
xnor UO_1863 (O_1863,N_29889,N_25059);
or UO_1864 (O_1864,N_25866,N_20698);
nor UO_1865 (O_1865,N_29878,N_27130);
xnor UO_1866 (O_1866,N_21564,N_28894);
nor UO_1867 (O_1867,N_27321,N_22383);
nor UO_1868 (O_1868,N_27537,N_22862);
nor UO_1869 (O_1869,N_29243,N_25576);
nor UO_1870 (O_1870,N_27947,N_23778);
xnor UO_1871 (O_1871,N_27964,N_26143);
nand UO_1872 (O_1872,N_24882,N_21076);
nand UO_1873 (O_1873,N_23740,N_24291);
or UO_1874 (O_1874,N_24736,N_29318);
and UO_1875 (O_1875,N_20882,N_22911);
and UO_1876 (O_1876,N_29063,N_27962);
xor UO_1877 (O_1877,N_21198,N_25641);
nor UO_1878 (O_1878,N_21014,N_24364);
or UO_1879 (O_1879,N_25142,N_24112);
and UO_1880 (O_1880,N_23280,N_25289);
or UO_1881 (O_1881,N_23977,N_27076);
and UO_1882 (O_1882,N_22194,N_25704);
xnor UO_1883 (O_1883,N_20394,N_23815);
or UO_1884 (O_1884,N_28055,N_21403);
nand UO_1885 (O_1885,N_29885,N_20054);
xor UO_1886 (O_1886,N_29852,N_26437);
xnor UO_1887 (O_1887,N_23308,N_24718);
nor UO_1888 (O_1888,N_28899,N_24932);
or UO_1889 (O_1889,N_27673,N_28293);
and UO_1890 (O_1890,N_20513,N_23310);
nand UO_1891 (O_1891,N_20107,N_29311);
or UO_1892 (O_1892,N_29037,N_22912);
or UO_1893 (O_1893,N_21883,N_29054);
or UO_1894 (O_1894,N_29828,N_28420);
nor UO_1895 (O_1895,N_20195,N_24357);
and UO_1896 (O_1896,N_21917,N_26945);
xor UO_1897 (O_1897,N_23924,N_21664);
nand UO_1898 (O_1898,N_26723,N_28078);
nor UO_1899 (O_1899,N_23767,N_21258);
or UO_1900 (O_1900,N_24894,N_24244);
nand UO_1901 (O_1901,N_24307,N_28437);
nor UO_1902 (O_1902,N_29310,N_23577);
nand UO_1903 (O_1903,N_29869,N_25220);
or UO_1904 (O_1904,N_29481,N_22750);
and UO_1905 (O_1905,N_26478,N_22573);
nor UO_1906 (O_1906,N_25562,N_27895);
nand UO_1907 (O_1907,N_23359,N_20916);
xor UO_1908 (O_1908,N_28181,N_20430);
or UO_1909 (O_1909,N_20145,N_21163);
nor UO_1910 (O_1910,N_27775,N_21693);
and UO_1911 (O_1911,N_28278,N_23938);
xor UO_1912 (O_1912,N_25805,N_23465);
or UO_1913 (O_1913,N_25601,N_28300);
nor UO_1914 (O_1914,N_24131,N_27557);
and UO_1915 (O_1915,N_21929,N_22325);
and UO_1916 (O_1916,N_21417,N_24238);
nor UO_1917 (O_1917,N_22586,N_21797);
or UO_1918 (O_1918,N_26452,N_22817);
xor UO_1919 (O_1919,N_29592,N_20063);
and UO_1920 (O_1920,N_23712,N_24368);
and UO_1921 (O_1921,N_22553,N_26781);
and UO_1922 (O_1922,N_29827,N_21358);
nor UO_1923 (O_1923,N_28067,N_21545);
xnor UO_1924 (O_1924,N_27919,N_21037);
nand UO_1925 (O_1925,N_25528,N_20187);
nand UO_1926 (O_1926,N_26241,N_23297);
nor UO_1927 (O_1927,N_20557,N_29251);
nand UO_1928 (O_1928,N_25204,N_22373);
nand UO_1929 (O_1929,N_25130,N_20041);
xnor UO_1930 (O_1930,N_27211,N_23254);
or UO_1931 (O_1931,N_22915,N_21427);
nand UO_1932 (O_1932,N_24309,N_28709);
and UO_1933 (O_1933,N_23241,N_23480);
or UO_1934 (O_1934,N_21567,N_26324);
nor UO_1935 (O_1935,N_26898,N_20490);
nor UO_1936 (O_1936,N_27961,N_23073);
xnor UO_1937 (O_1937,N_25035,N_23478);
xor UO_1938 (O_1938,N_27613,N_21968);
xor UO_1939 (O_1939,N_25905,N_26383);
or UO_1940 (O_1940,N_29209,N_22346);
or UO_1941 (O_1941,N_27465,N_24257);
or UO_1942 (O_1942,N_28206,N_27596);
and UO_1943 (O_1943,N_23910,N_29867);
xor UO_1944 (O_1944,N_22927,N_26974);
nor UO_1945 (O_1945,N_20562,N_25885);
xnor UO_1946 (O_1946,N_27306,N_27646);
nand UO_1947 (O_1947,N_23669,N_27056);
xnor UO_1948 (O_1948,N_23603,N_20996);
and UO_1949 (O_1949,N_26129,N_29052);
or UO_1950 (O_1950,N_22175,N_28397);
nand UO_1951 (O_1951,N_21297,N_25808);
nand UO_1952 (O_1952,N_28301,N_23706);
and UO_1953 (O_1953,N_29553,N_25687);
and UO_1954 (O_1954,N_23532,N_21259);
nor UO_1955 (O_1955,N_28799,N_20040);
nor UO_1956 (O_1956,N_25012,N_28159);
nand UO_1957 (O_1957,N_24049,N_24896);
nand UO_1958 (O_1958,N_25102,N_29776);
or UO_1959 (O_1959,N_25770,N_28506);
nor UO_1960 (O_1960,N_24818,N_28107);
and UO_1961 (O_1961,N_20306,N_25223);
nand UO_1962 (O_1962,N_29278,N_27063);
nor UO_1963 (O_1963,N_26207,N_29795);
or UO_1964 (O_1964,N_28670,N_28211);
or UO_1965 (O_1965,N_29360,N_23724);
or UO_1966 (O_1966,N_22910,N_20579);
nand UO_1967 (O_1967,N_27402,N_20767);
nand UO_1968 (O_1968,N_20269,N_21618);
or UO_1969 (O_1969,N_26444,N_23837);
or UO_1970 (O_1970,N_23364,N_24070);
xor UO_1971 (O_1971,N_20832,N_28990);
or UO_1972 (O_1972,N_21148,N_26597);
nor UO_1973 (O_1973,N_22827,N_27458);
and UO_1974 (O_1974,N_22917,N_21615);
and UO_1975 (O_1975,N_27361,N_26331);
xor UO_1976 (O_1976,N_26116,N_28490);
and UO_1977 (O_1977,N_28307,N_21302);
nand UO_1978 (O_1978,N_27298,N_22492);
nand UO_1979 (O_1979,N_29583,N_20039);
xor UO_1980 (O_1980,N_28783,N_26293);
and UO_1981 (O_1981,N_24880,N_25550);
and UO_1982 (O_1982,N_23450,N_29201);
or UO_1983 (O_1983,N_29599,N_29606);
nand UO_1984 (O_1984,N_27693,N_23335);
and UO_1985 (O_1985,N_23630,N_24130);
xnor UO_1986 (O_1986,N_22136,N_24967);
nand UO_1987 (O_1987,N_21606,N_25489);
and UO_1988 (O_1988,N_25953,N_26685);
or UO_1989 (O_1989,N_24964,N_27149);
and UO_1990 (O_1990,N_23245,N_22522);
xor UO_1991 (O_1991,N_27572,N_23009);
or UO_1992 (O_1992,N_20626,N_20130);
nand UO_1993 (O_1993,N_22478,N_23721);
nor UO_1994 (O_1994,N_22789,N_26200);
nand UO_1995 (O_1995,N_20074,N_28358);
nand UO_1996 (O_1996,N_21722,N_29081);
xor UO_1997 (O_1997,N_22680,N_22541);
nor UO_1998 (O_1998,N_25752,N_21018);
nand UO_1999 (O_1999,N_24153,N_27567);
nor UO_2000 (O_2000,N_21048,N_21717);
nand UO_2001 (O_2001,N_24133,N_21013);
xnor UO_2002 (O_2002,N_24944,N_23925);
and UO_2003 (O_2003,N_23593,N_27657);
xnor UO_2004 (O_2004,N_21381,N_27288);
or UO_2005 (O_2005,N_24143,N_21415);
xor UO_2006 (O_2006,N_29229,N_23442);
or UO_2007 (O_2007,N_25463,N_24313);
or UO_2008 (O_2008,N_22524,N_22322);
nand UO_2009 (O_2009,N_20663,N_21746);
and UO_2010 (O_2010,N_25386,N_25351);
and UO_2011 (O_2011,N_24379,N_20514);
and UO_2012 (O_2012,N_21592,N_29105);
nor UO_2013 (O_2013,N_22886,N_21878);
or UO_2014 (O_2014,N_22143,N_24995);
xnor UO_2015 (O_2015,N_21159,N_25239);
or UO_2016 (O_2016,N_29089,N_21673);
and UO_2017 (O_2017,N_23346,N_25594);
xnor UO_2018 (O_2018,N_29994,N_25332);
or UO_2019 (O_2019,N_25563,N_27308);
nor UO_2020 (O_2020,N_20501,N_29794);
or UO_2021 (O_2021,N_29175,N_21998);
or UO_2022 (O_2022,N_22968,N_20347);
nor UO_2023 (O_2023,N_23751,N_24288);
nand UO_2024 (O_2024,N_26163,N_26512);
or UO_2025 (O_2025,N_25632,N_27803);
nand UO_2026 (O_2026,N_24697,N_23325);
nor UO_2027 (O_2027,N_22331,N_27786);
or UO_2028 (O_2028,N_20120,N_25187);
or UO_2029 (O_2029,N_22540,N_21450);
or UO_2030 (O_2030,N_26379,N_27897);
nor UO_2031 (O_2031,N_26178,N_20865);
nor UO_2032 (O_2032,N_28938,N_25554);
and UO_2033 (O_2033,N_26728,N_20862);
nor UO_2034 (O_2034,N_28924,N_26746);
or UO_2035 (O_2035,N_27326,N_24606);
or UO_2036 (O_2036,N_24154,N_28636);
xnor UO_2037 (O_2037,N_26352,N_21174);
nand UO_2038 (O_2038,N_26135,N_22885);
and UO_2039 (O_2039,N_29082,N_23665);
nand UO_2040 (O_2040,N_24079,N_25233);
xor UO_2041 (O_2041,N_20383,N_28993);
xnor UO_2042 (O_2042,N_27225,N_24258);
and UO_2043 (O_2043,N_22503,N_22216);
and UO_2044 (O_2044,N_22090,N_29566);
xnor UO_2045 (O_2045,N_29780,N_25370);
nand UO_2046 (O_2046,N_21780,N_29305);
and UO_2047 (O_2047,N_20568,N_27385);
xor UO_2048 (O_2048,N_22285,N_29690);
xnor UO_2049 (O_2049,N_20635,N_21335);
nor UO_2050 (O_2050,N_28409,N_21404);
nand UO_2051 (O_2051,N_29754,N_20919);
or UO_2052 (O_2052,N_22820,N_28095);
nand UO_2053 (O_2053,N_26806,N_29952);
nor UO_2054 (O_2054,N_29098,N_25597);
and UO_2055 (O_2055,N_27692,N_27955);
nor UO_2056 (O_2056,N_28118,N_25448);
nor UO_2057 (O_2057,N_22137,N_23012);
and UO_2058 (O_2058,N_22093,N_23214);
nand UO_2059 (O_2059,N_27080,N_21613);
nand UO_2060 (O_2060,N_26666,N_26803);
nand UO_2061 (O_2061,N_22890,N_20760);
nand UO_2062 (O_2062,N_21595,N_21368);
nor UO_2063 (O_2063,N_21834,N_25093);
xor UO_2064 (O_2064,N_20651,N_29584);
and UO_2065 (O_2065,N_26094,N_26968);
and UO_2066 (O_2066,N_29799,N_21869);
or UO_2067 (O_2067,N_21193,N_21332);
xnor UO_2068 (O_2068,N_20723,N_27017);
nand UO_2069 (O_2069,N_23853,N_22521);
nor UO_2070 (O_2070,N_29406,N_28419);
xor UO_2071 (O_2071,N_20448,N_28359);
and UO_2072 (O_2072,N_24365,N_25176);
or UO_2073 (O_2073,N_26317,N_27315);
nor UO_2074 (O_2074,N_20267,N_24886);
or UO_2075 (O_2075,N_28614,N_21278);
nor UO_2076 (O_2076,N_27652,N_24873);
and UO_2077 (O_2077,N_27605,N_28204);
and UO_2078 (O_2078,N_28663,N_28931);
or UO_2079 (O_2079,N_21649,N_21106);
nor UO_2080 (O_2080,N_28732,N_22849);
or UO_2081 (O_2081,N_25302,N_23980);
xor UO_2082 (O_2082,N_20571,N_26077);
or UO_2083 (O_2083,N_27901,N_25069);
xor UO_2084 (O_2084,N_24837,N_25281);
nor UO_2085 (O_2085,N_26818,N_29641);
or UO_2086 (O_2086,N_27162,N_24674);
nand UO_2087 (O_2087,N_29121,N_24908);
xnor UO_2088 (O_2088,N_25964,N_27000);
xnor UO_2089 (O_2089,N_23791,N_29482);
nand UO_2090 (O_2090,N_29647,N_29451);
and UO_2091 (O_2091,N_25472,N_20537);
or UO_2092 (O_2092,N_21412,N_28209);
nand UO_2093 (O_2093,N_27128,N_26670);
and UO_2094 (O_2094,N_29697,N_21184);
nand UO_2095 (O_2095,N_20775,N_20013);
nor UO_2096 (O_2096,N_21288,N_26176);
or UO_2097 (O_2097,N_23999,N_29023);
nor UO_2098 (O_2098,N_22185,N_20915);
nand UO_2099 (O_2099,N_23887,N_28139);
xor UO_2100 (O_2100,N_22807,N_21064);
nor UO_2101 (O_2101,N_24778,N_29313);
or UO_2102 (O_2102,N_29449,N_28523);
xor UO_2103 (O_2103,N_21925,N_29985);
nor UO_2104 (O_2104,N_29087,N_20406);
xor UO_2105 (O_2105,N_28319,N_29257);
and UO_2106 (O_2106,N_25864,N_21653);
nand UO_2107 (O_2107,N_20399,N_26880);
xnor UO_2108 (O_2108,N_28773,N_27503);
and UO_2109 (O_2109,N_25621,N_28657);
nor UO_2110 (O_2110,N_24579,N_27486);
nand UO_2111 (O_2111,N_28402,N_28349);
nor UO_2112 (O_2112,N_21660,N_21831);
or UO_2113 (O_2113,N_29212,N_29568);
nor UO_2114 (O_2114,N_21953,N_29634);
nor UO_2115 (O_2115,N_28578,N_22896);
xnor UO_2116 (O_2116,N_28129,N_22595);
and UO_2117 (O_2117,N_20592,N_26042);
xor UO_2118 (O_2118,N_24538,N_26290);
and UO_2119 (O_2119,N_22683,N_25795);
or UO_2120 (O_2120,N_29518,N_28528);
xnor UO_2121 (O_2121,N_24445,N_26951);
xor UO_2122 (O_2122,N_24156,N_24241);
nand UO_2123 (O_2123,N_25730,N_24544);
nor UO_2124 (O_2124,N_27816,N_26457);
nor UO_2125 (O_2125,N_28302,N_24047);
nor UO_2126 (O_2126,N_21651,N_28526);
nand UO_2127 (O_2127,N_23908,N_20652);
or UO_2128 (O_2128,N_27821,N_29820);
and UO_2129 (O_2129,N_28508,N_21144);
xnor UO_2130 (O_2130,N_20899,N_24100);
xnor UO_2131 (O_2131,N_21762,N_22603);
and UO_2132 (O_2132,N_20846,N_21875);
nor UO_2133 (O_2133,N_26881,N_20007);
or UO_2134 (O_2134,N_26595,N_26076);
and UO_2135 (O_2135,N_23142,N_21032);
and UO_2136 (O_2136,N_24983,N_23434);
and UO_2137 (O_2137,N_21768,N_28053);
or UO_2138 (O_2138,N_25445,N_25328);
or UO_2139 (O_2139,N_25166,N_27398);
and UO_2140 (O_2140,N_29353,N_27042);
nand UO_2141 (O_2141,N_29591,N_20561);
or UO_2142 (O_2142,N_28704,N_23031);
xnor UO_2143 (O_2143,N_23972,N_26363);
or UO_2144 (O_2144,N_24826,N_28751);
xor UO_2145 (O_2145,N_24771,N_27452);
xor UO_2146 (O_2146,N_23424,N_24782);
or UO_2147 (O_2147,N_25020,N_25168);
or UO_2148 (O_2148,N_28700,N_24035);
nand UO_2149 (O_2149,N_23578,N_22975);
or UO_2150 (O_2150,N_23883,N_24374);
nand UO_2151 (O_2151,N_21517,N_25136);
nand UO_2152 (O_2152,N_29411,N_22951);
xor UO_2153 (O_2153,N_21425,N_24304);
and UO_2154 (O_2154,N_27916,N_29860);
and UO_2155 (O_2155,N_25636,N_23386);
or UO_2156 (O_2156,N_28739,N_24420);
nor UO_2157 (O_2157,N_28439,N_20681);
nor UO_2158 (O_2158,N_23535,N_20190);
nand UO_2159 (O_2159,N_20572,N_25080);
or UO_2160 (O_2160,N_20741,N_20137);
xor UO_2161 (O_2161,N_20520,N_28477);
xor UO_2162 (O_2162,N_24562,N_25114);
nor UO_2163 (O_2163,N_26302,N_29609);
xnor UO_2164 (O_2164,N_25545,N_26805);
xor UO_2165 (O_2165,N_20442,N_22947);
nand UO_2166 (O_2166,N_26661,N_21643);
nand UO_2167 (O_2167,N_22834,N_24830);
nor UO_2168 (O_2168,N_26791,N_20295);
xnor UO_2169 (O_2169,N_21040,N_24607);
nor UO_2170 (O_2170,N_26934,N_20169);
nor UO_2171 (O_2171,N_24163,N_21558);
nor UO_2172 (O_2172,N_24419,N_27009);
nand UO_2173 (O_2173,N_28530,N_28928);
xor UO_2174 (O_2174,N_27526,N_24539);
nor UO_2175 (O_2175,N_28160,N_29359);
nor UO_2176 (O_2176,N_21521,N_29826);
xnor UO_2177 (O_2177,N_24727,N_21965);
nand UO_2178 (O_2178,N_28310,N_26056);
xnor UO_2179 (O_2179,N_25837,N_25697);
nand UO_2180 (O_2180,N_28543,N_28191);
or UO_2181 (O_2181,N_24730,N_26735);
nand UO_2182 (O_2182,N_27284,N_23668);
and UO_2183 (O_2183,N_22323,N_26538);
nand UO_2184 (O_2184,N_20498,N_29396);
nand UO_2185 (O_2185,N_25389,N_29191);
nand UO_2186 (O_2186,N_29176,N_26333);
or UO_2187 (O_2187,N_28973,N_29370);
or UO_2188 (O_2188,N_22388,N_22150);
nor UO_2189 (O_2189,N_29442,N_27926);
and UO_2190 (O_2190,N_20887,N_21290);
or UO_2191 (O_2191,N_27007,N_21559);
xor UO_2192 (O_2192,N_28084,N_24998);
xor UO_2193 (O_2193,N_26009,N_23227);
nor UO_2194 (O_2194,N_22646,N_20100);
nor UO_2195 (O_2195,N_23238,N_28399);
or UO_2196 (O_2196,N_25188,N_20590);
nor UO_2197 (O_2197,N_21149,N_29203);
and UO_2198 (O_2198,N_20364,N_24711);
nand UO_2199 (O_2199,N_20874,N_22105);
and UO_2200 (O_2200,N_24449,N_26429);
xnor UO_2201 (O_2201,N_20186,N_29504);
nand UO_2202 (O_2202,N_27287,N_28444);
and UO_2203 (O_2203,N_29125,N_24343);
and UO_2204 (O_2204,N_29733,N_23699);
nor UO_2205 (O_2205,N_21405,N_21529);
or UO_2206 (O_2206,N_28172,N_21073);
xnor UO_2207 (O_2207,N_22508,N_23114);
or UO_2208 (O_2208,N_27062,N_29946);
nor UO_2209 (O_2209,N_24292,N_29280);
xor UO_2210 (O_2210,N_26824,N_24392);
xnor UO_2211 (O_2211,N_23659,N_25277);
nand UO_2212 (O_2212,N_20964,N_21001);
or UO_2213 (O_2213,N_29605,N_28117);
and UO_2214 (O_2214,N_27414,N_20486);
nor UO_2215 (O_2215,N_21889,N_21419);
nand UO_2216 (O_2216,N_23458,N_24138);
and UO_2217 (O_2217,N_21888,N_22534);
or UO_2218 (O_2218,N_22814,N_29758);
xor UO_2219 (O_2219,N_25371,N_26617);
and UO_2220 (O_2220,N_27779,N_28898);
nor UO_2221 (O_2221,N_25215,N_27204);
and UO_2222 (O_2222,N_26206,N_29440);
nand UO_2223 (O_2223,N_22632,N_27667);
xnor UO_2224 (O_2224,N_23483,N_21846);
xor UO_2225 (O_2225,N_21295,N_26693);
xnor UO_2226 (O_2226,N_25586,N_27911);
nor UO_2227 (O_2227,N_22118,N_27940);
or UO_2228 (O_2228,N_29833,N_26852);
nand UO_2229 (O_2229,N_20445,N_28770);
nor UO_2230 (O_2230,N_26107,N_23677);
or UO_2231 (O_2231,N_23259,N_28879);
xor UO_2232 (O_2232,N_21316,N_27653);
and UO_2233 (O_2233,N_25785,N_20404);
nor UO_2234 (O_2234,N_23548,N_20742);
nand UO_2235 (O_2235,N_26748,N_26075);
xor UO_2236 (O_2236,N_26659,N_23288);
xor UO_2237 (O_2237,N_26863,N_29868);
nand UO_2238 (O_2238,N_20480,N_28851);
xor UO_2239 (O_2239,N_23589,N_20105);
and UO_2240 (O_2240,N_21932,N_22713);
and UO_2241 (O_2241,N_21436,N_24583);
nor UO_2242 (O_2242,N_23119,N_26499);
or UO_2243 (O_2243,N_23388,N_23376);
or UO_2244 (O_2244,N_27923,N_22877);
and UO_2245 (O_2245,N_27764,N_21356);
nand UO_2246 (O_2246,N_29244,N_25615);
nand UO_2247 (O_2247,N_26883,N_20658);
or UO_2248 (O_2248,N_28414,N_24493);
nand UO_2249 (O_2249,N_22129,N_25896);
nor UO_2250 (O_2250,N_24763,N_28681);
and UO_2251 (O_2251,N_20839,N_22919);
nor UO_2252 (O_2252,N_26277,N_23743);
xnor UO_2253 (O_2253,N_27469,N_23754);
xor UO_2254 (O_2254,N_26140,N_24689);
and UO_2255 (O_2255,N_22265,N_29424);
nor UO_2256 (O_2256,N_21272,N_28100);
nor UO_2257 (O_2257,N_25997,N_25413);
nor UO_2258 (O_2258,N_28316,N_22852);
and UO_2259 (O_2259,N_24671,N_27432);
xnor UO_2260 (O_2260,N_25040,N_27312);
xor UO_2261 (O_2261,N_24225,N_29334);
nand UO_2262 (O_2262,N_28873,N_22351);
nand UO_2263 (O_2263,N_28540,N_23586);
nand UO_2264 (O_2264,N_20240,N_22981);
and UO_2265 (O_2265,N_21774,N_20689);
nand UO_2266 (O_2266,N_20939,N_28474);
nand UO_2267 (O_2267,N_23715,N_26089);
nand UO_2268 (O_2268,N_24570,N_22284);
xor UO_2269 (O_2269,N_24895,N_27716);
xnor UO_2270 (O_2270,N_25004,N_22464);
and UO_2271 (O_2271,N_27582,N_27612);
nand UO_2272 (O_2272,N_22966,N_26430);
xor UO_2273 (O_2273,N_20075,N_28761);
nor UO_2274 (O_2274,N_23856,N_28184);
or UO_2275 (O_2275,N_26513,N_26982);
xnor UO_2276 (O_2276,N_24942,N_28720);
nor UO_2277 (O_2277,N_23943,N_28947);
and UO_2278 (O_2278,N_23606,N_23216);
nor UO_2279 (O_2279,N_27520,N_29519);
or UO_2280 (O_2280,N_24829,N_27643);
or UO_2281 (O_2281,N_23371,N_28007);
xnor UO_2282 (O_2282,N_27220,N_24618);
nor UO_2283 (O_2283,N_24957,N_29962);
and UO_2284 (O_2284,N_28081,N_26910);
nor UO_2285 (O_2285,N_22668,N_27998);
and UO_2286 (O_2286,N_20823,N_26368);
or UO_2287 (O_2287,N_24863,N_20777);
or UO_2288 (O_2288,N_23276,N_22692);
and UO_2289 (O_2289,N_20552,N_21702);
xnor UO_2290 (O_2290,N_29752,N_21200);
and UO_2291 (O_2291,N_20973,N_21732);
and UO_2292 (O_2292,N_29629,N_23932);
or UO_2293 (O_2293,N_20094,N_28525);
nand UO_2294 (O_2294,N_25341,N_29286);
nand UO_2295 (O_2295,N_28188,N_24320);
nand UO_2296 (O_2296,N_22839,N_25110);
nor UO_2297 (O_2297,N_28855,N_26590);
xnor UO_2298 (O_2298,N_21362,N_28247);
nor UO_2299 (O_2299,N_27517,N_26036);
xor UO_2300 (O_2300,N_20727,N_27731);
or UO_2301 (O_2301,N_22709,N_26950);
and UO_2302 (O_2302,N_26372,N_22986);
or UO_2303 (O_2303,N_28539,N_27574);
xor UO_2304 (O_2304,N_20388,N_23757);
xnor UO_2305 (O_2305,N_24693,N_21983);
nor UO_2306 (O_2306,N_26369,N_28171);
xnor UO_2307 (O_2307,N_27391,N_28828);
and UO_2308 (O_2308,N_26160,N_26689);
nand UO_2309 (O_2309,N_20465,N_24360);
nand UO_2310 (O_2310,N_29190,N_26471);
xor UO_2311 (O_2311,N_24716,N_27189);
xnor UO_2312 (O_2312,N_21659,N_24361);
and UO_2313 (O_2313,N_22367,N_20358);
and UO_2314 (O_2314,N_22491,N_24531);
nand UO_2315 (O_2315,N_29873,N_29503);
nand UO_2316 (O_2316,N_23838,N_22734);
nor UO_2317 (O_2317,N_24482,N_25707);
xnor UO_2318 (O_2318,N_28226,N_25890);
nor UO_2319 (O_2319,N_20200,N_21418);
nor UO_2320 (O_2320,N_27318,N_26667);
nand UO_2321 (O_2321,N_29725,N_25055);
and UO_2322 (O_2322,N_23676,N_24194);
nand UO_2323 (O_2323,N_24207,N_22926);
nand UO_2324 (O_2324,N_24438,N_21710);
or UO_2325 (O_2325,N_28629,N_20469);
xor UO_2326 (O_2326,N_28048,N_23431);
nand UO_2327 (O_2327,N_24768,N_29677);
xor UO_2328 (O_2328,N_21867,N_27045);
nand UO_2329 (O_2329,N_26526,N_21022);
and UO_2330 (O_2330,N_22850,N_21575);
nor UO_2331 (O_2331,N_29200,N_21759);
and UO_2332 (O_2332,N_28116,N_24433);
xor UO_2333 (O_2333,N_24907,N_26810);
or UO_2334 (O_2334,N_26282,N_21612);
nand UO_2335 (O_2335,N_20946,N_22805);
nor UO_2336 (O_2336,N_26920,N_28113);
xnor UO_2337 (O_2337,N_26786,N_28555);
nor UO_2338 (O_2338,N_20277,N_21078);
xor UO_2339 (O_2339,N_25067,N_24083);
nor UO_2340 (O_2340,N_25190,N_23555);
nand UO_2341 (O_2341,N_28137,N_21410);
and UO_2342 (O_2342,N_20276,N_25726);
or UO_2343 (O_2343,N_24007,N_24227);
xor UO_2344 (O_2344,N_27455,N_25618);
nor UO_2345 (O_2345,N_20092,N_28017);
or UO_2346 (O_2346,N_27878,N_27293);
or UO_2347 (O_2347,N_27393,N_26327);
nor UO_2348 (O_2348,N_20648,N_21388);
xor UO_2349 (O_2349,N_20970,N_24621);
nor UO_2350 (O_2350,N_28796,N_28812);
nand UO_2351 (O_2351,N_20429,N_24858);
xor UO_2352 (O_2352,N_24308,N_22787);
xnor UO_2353 (O_2353,N_25021,N_25486);
or UO_2354 (O_2354,N_28431,N_24213);
nor UO_2355 (O_2355,N_28096,N_29544);
xor UO_2356 (O_2356,N_25430,N_21534);
nand UO_2357 (O_2357,N_22399,N_23672);
nand UO_2358 (O_2358,N_24048,N_22796);
or UO_2359 (O_2359,N_29939,N_25297);
and UO_2360 (O_2360,N_28325,N_20208);
and UO_2361 (O_2361,N_21550,N_27370);
or UO_2362 (O_2362,N_26173,N_20851);
xnor UO_2363 (O_2363,N_25660,N_29972);
xor UO_2364 (O_2364,N_25353,N_22497);
nor UO_2365 (O_2365,N_26274,N_25552);
or UO_2366 (O_2366,N_29659,N_22621);
or UO_2367 (O_2367,N_21989,N_22952);
or UO_2368 (O_2368,N_22544,N_23915);
nand UO_2369 (O_2369,N_23207,N_20631);
or UO_2370 (O_2370,N_24695,N_26249);
nand UO_2371 (O_2371,N_25005,N_29597);
nand UO_2372 (O_2372,N_28605,N_27847);
or UO_2373 (O_2373,N_20649,N_24428);
nor UO_2374 (O_2374,N_28975,N_27992);
and UO_2375 (O_2375,N_25458,N_27024);
and UO_2376 (O_2376,N_28249,N_22687);
nor UO_2377 (O_2377,N_26687,N_27134);
nor UO_2378 (O_2378,N_21024,N_26816);
and UO_2379 (O_2379,N_23355,N_25388);
nor UO_2380 (O_2380,N_27388,N_24648);
nand UO_2381 (O_2381,N_22761,N_28520);
and UO_2382 (O_2382,N_24115,N_26848);
or UO_2383 (O_2383,N_23860,N_29299);
nor UO_2384 (O_2384,N_20402,N_20844);
or UO_2385 (O_2385,N_26147,N_28021);
and UO_2386 (O_2386,N_29608,N_22701);
xnor UO_2387 (O_2387,N_21523,N_27739);
nor UO_2388 (O_2388,N_26992,N_21848);
nor UO_2389 (O_2389,N_24056,N_22556);
nand UO_2390 (O_2390,N_25155,N_26649);
and UO_2391 (O_2391,N_27127,N_22130);
nor UO_2392 (O_2392,N_29245,N_25077);
nor UO_2393 (O_2393,N_20976,N_28661);
xor UO_2394 (O_2394,N_23342,N_23061);
xnor UO_2395 (O_2395,N_23264,N_23508);
nor UO_2396 (O_2396,N_22280,N_24121);
nand UO_2397 (O_2397,N_26624,N_25855);
or UO_2398 (O_2398,N_20349,N_29419);
nand UO_2399 (O_2399,N_23574,N_20427);
nand UO_2400 (O_2400,N_21895,N_22589);
nor UO_2401 (O_2401,N_28252,N_26998);
or UO_2402 (O_2402,N_20838,N_27941);
or UO_2403 (O_2403,N_27583,N_22930);
xnor UO_2404 (O_2404,N_25304,N_29112);
nor UO_2405 (O_2405,N_22584,N_21866);
xor UO_2406 (O_2406,N_24484,N_27622);
xnor UO_2407 (O_2407,N_21607,N_22539);
xor UO_2408 (O_2408,N_27852,N_23934);
and UO_2409 (O_2409,N_22063,N_26459);
xor UO_2410 (O_2410,N_25629,N_20858);
nor UO_2411 (O_2411,N_29458,N_27265);
xnor UO_2412 (O_2412,N_26917,N_20084);
and UO_2413 (O_2413,N_22617,N_27853);
and UO_2414 (O_2414,N_28731,N_26897);
nand UO_2415 (O_2415,N_20308,N_29384);
xor UO_2416 (O_2416,N_24192,N_20668);
xor UO_2417 (O_2417,N_24638,N_23616);
or UO_2418 (O_2418,N_20352,N_28241);
xor UO_2419 (O_2419,N_24759,N_29595);
nor UO_2420 (O_2420,N_22167,N_26851);
or UO_2421 (O_2421,N_22700,N_28780);
xnor UO_2422 (O_2422,N_28602,N_20056);
nor UO_2423 (O_2423,N_23747,N_29169);
or UO_2424 (O_2424,N_29539,N_21907);
nand UO_2425 (O_2425,N_23309,N_23737);
nand UO_2426 (O_2426,N_29521,N_22260);
or UO_2427 (O_2427,N_20474,N_28680);
xor UO_2428 (O_2428,N_29260,N_22414);
nor UO_2429 (O_2429,N_21611,N_23316);
xor UO_2430 (O_2430,N_29092,N_20238);
nand UO_2431 (O_2431,N_27320,N_25330);
or UO_2432 (O_2432,N_25269,N_22433);
xnor UO_2433 (O_2433,N_28412,N_22863);
xor UO_2434 (O_2434,N_29619,N_20078);
xnor UO_2435 (O_2435,N_20773,N_25721);
and UO_2436 (O_2436,N_27770,N_25201);
nor UO_2437 (O_2437,N_21626,N_22291);
or UO_2438 (O_2438,N_27863,N_21111);
and UO_2439 (O_2439,N_26688,N_29542);
or UO_2440 (O_2440,N_20620,N_27913);
or UO_2441 (O_2441,N_21089,N_24038);
xor UO_2442 (O_2442,N_21392,N_28024);
xor UO_2443 (O_2443,N_22008,N_20101);
or UO_2444 (O_2444,N_26817,N_25284);
nand UO_2445 (O_2445,N_25974,N_26776);
or UO_2446 (O_2446,N_26417,N_22555);
and UO_2447 (O_2447,N_25631,N_24436);
nand UO_2448 (O_2448,N_25256,N_29110);
nor UO_2449 (O_2449,N_23675,N_21266);
nand UO_2450 (O_2450,N_27809,N_24303);
nor UO_2451 (O_2451,N_25367,N_24502);
nor UO_2452 (O_2452,N_28415,N_26841);
or UO_2453 (O_2453,N_20779,N_27677);
and UO_2454 (O_2454,N_24476,N_21535);
or UO_2455 (O_2455,N_23904,N_22411);
and UO_2456 (O_2456,N_27403,N_27942);
xor UO_2457 (O_2457,N_26402,N_22500);
nor UO_2458 (O_2458,N_27494,N_27920);
nand UO_2459 (O_2459,N_25812,N_26614);
and UO_2460 (O_2460,N_28630,N_21197);
nor UO_2461 (O_2461,N_27588,N_22068);
xnor UO_2462 (O_2462,N_27383,N_20587);
nand UO_2463 (O_2463,N_25897,N_23441);
nand UO_2464 (O_2464,N_29964,N_21901);
nand UO_2465 (O_2465,N_22485,N_22188);
and UO_2466 (O_2466,N_26971,N_26336);
nand UO_2467 (O_2467,N_29522,N_29216);
xor UO_2468 (O_2468,N_28967,N_26409);
nor UO_2469 (O_2469,N_29223,N_24599);
nor UO_2470 (O_2470,N_20632,N_23224);
nor UO_2471 (O_2471,N_26315,N_26750);
nor UO_2472 (O_2472,N_20055,N_28668);
and UO_2473 (O_2473,N_26535,N_26865);
nor UO_2474 (O_2474,N_20436,N_21314);
or UO_2475 (O_2475,N_21730,N_25581);
xor UO_2476 (O_2476,N_21267,N_21949);
or UO_2477 (O_2477,N_27165,N_22407);
xor UO_2478 (O_2478,N_28695,N_21067);
nand UO_2479 (O_2479,N_29315,N_22685);
and UO_2480 (O_2480,N_24513,N_25348);
and UO_2481 (O_2481,N_28575,N_27022);
nand UO_2482 (O_2482,N_23438,N_24234);
xnor UO_2483 (O_2483,N_21115,N_29823);
and UO_2484 (O_2484,N_21019,N_25003);
nor UO_2485 (O_2485,N_24973,N_29378);
nor UO_2486 (O_2486,N_27480,N_25591);
and UO_2487 (O_2487,N_25680,N_29235);
nand UO_2488 (O_2488,N_23525,N_26350);
xor UO_2489 (O_2489,N_20242,N_20457);
nor UO_2490 (O_2490,N_25089,N_28059);
and UO_2491 (O_2491,N_21470,N_20847);
or UO_2492 (O_2492,N_23192,N_23240);
or UO_2493 (O_2493,N_24116,N_24954);
nand UO_2494 (O_2494,N_27010,N_20389);
or UO_2495 (O_2495,N_29390,N_29314);
or UO_2496 (O_2496,N_25042,N_26300);
xor UO_2497 (O_2497,N_29514,N_24358);
xor UO_2498 (O_2498,N_27556,N_24982);
nand UO_2499 (O_2499,N_26830,N_29489);
xnor UO_2500 (O_2500,N_25107,N_27039);
and UO_2501 (O_2501,N_27899,N_21974);
nor UO_2502 (O_2502,N_26243,N_26596);
nor UO_2503 (O_2503,N_25248,N_21139);
nor UO_2504 (O_2504,N_24946,N_21219);
and UO_2505 (O_2505,N_20603,N_29739);
nand UO_2506 (O_2506,N_24362,N_23536);
or UO_2507 (O_2507,N_26947,N_22628);
xor UO_2508 (O_2508,N_20945,N_25199);
and UO_2509 (O_2509,N_24935,N_21498);
and UO_2510 (O_2510,N_22097,N_29341);
nor UO_2511 (O_2511,N_29956,N_22370);
or UO_2512 (O_2512,N_21591,N_21853);
nor UO_2513 (O_2513,N_28144,N_29291);
and UO_2514 (O_2514,N_22627,N_28020);
nand UO_2515 (O_2515,N_27496,N_23870);
or UO_2516 (O_2516,N_23828,N_22819);
or UO_2517 (O_2517,N_25116,N_22299);
or UO_2518 (O_2518,N_21838,N_22732);
nor UO_2519 (O_2519,N_26665,N_27918);
nand UO_2520 (O_2520,N_22386,N_24463);
xor UO_2521 (O_2521,N_26118,N_25693);
nand UO_2522 (O_2522,N_21630,N_22718);
xnor UO_2523 (O_2523,N_24015,N_26838);
and UO_2524 (O_2524,N_28154,N_26212);
nand UO_2525 (O_2525,N_22155,N_26610);
nand UO_2526 (O_2526,N_22100,N_26700);
or UO_2527 (O_2527,N_24297,N_24588);
nand UO_2528 (O_2528,N_26606,N_20491);
nand UO_2529 (O_2529,N_29049,N_23708);
xor UO_2530 (O_2530,N_20428,N_25431);
and UO_2531 (O_2531,N_28978,N_27423);
xnor UO_2532 (O_2532,N_25935,N_24447);
and UO_2533 (O_2533,N_24901,N_22659);
and UO_2534 (O_2534,N_23959,N_27623);
xnor UO_2535 (O_2535,N_28719,N_28841);
xor UO_2536 (O_2536,N_28386,N_28087);
xnor UO_2537 (O_2537,N_26635,N_29532);
and UO_2538 (O_2538,N_25123,N_22963);
xnor UO_2539 (O_2539,N_27033,N_29894);
or UO_2540 (O_2540,N_28037,N_27036);
or UO_2541 (O_2541,N_28696,N_22275);
nor UO_2542 (O_2542,N_22670,N_23892);
nand UO_2543 (O_2543,N_21293,N_29287);
xnor UO_2544 (O_2544,N_28533,N_26836);
nor UO_2545 (O_2545,N_29040,N_21728);
xnor UO_2546 (O_2546,N_20803,N_27185);
or UO_2547 (O_2547,N_28485,N_20301);
and UO_2548 (O_2548,N_28759,N_25477);
nand UO_2549 (O_2549,N_23130,N_23313);
nand UO_2550 (O_2550,N_25222,N_24836);
nor UO_2551 (O_2551,N_29866,N_20554);
nand UO_2552 (O_2552,N_25234,N_27935);
nand UO_2553 (O_2553,N_20362,N_23419);
xnor UO_2554 (O_2554,N_26490,N_20644);
and UO_2555 (O_2555,N_28012,N_22842);
or UO_2556 (O_2556,N_28519,N_29986);
nand UO_2557 (O_2557,N_21552,N_24760);
nor UO_2558 (O_2558,N_27730,N_25481);
or UO_2559 (O_2559,N_27898,N_23710);
nand UO_2560 (O_2560,N_21054,N_25725);
nor UO_2561 (O_2561,N_20625,N_27043);
or UO_2562 (O_2562,N_25995,N_23179);
and UO_2563 (O_2563,N_21581,N_27194);
and UO_2564 (O_2564,N_23071,N_27632);
nand UO_2565 (O_2565,N_22882,N_28110);
nand UO_2566 (O_2566,N_23222,N_20782);
nor UO_2567 (O_2567,N_23780,N_26028);
nand UO_2568 (O_2568,N_22960,N_23145);
xor UO_2569 (O_2569,N_23174,N_28423);
nand UO_2570 (O_2570,N_27949,N_26769);
xor UO_2571 (O_2571,N_29874,N_29502);
and UO_2572 (O_2572,N_20792,N_21372);
or UO_2573 (O_2573,N_26831,N_20622);
xor UO_2574 (O_2574,N_25813,N_22772);
and UO_2575 (O_2575,N_29126,N_21624);
xnor UO_2576 (O_2576,N_20005,N_25551);
and UO_2577 (O_2577,N_25470,N_20560);
or UO_2578 (O_2578,N_23958,N_28734);
nor UO_2579 (O_2579,N_29053,N_25702);
and UO_2580 (O_2580,N_20877,N_21454);
nand UO_2581 (O_2581,N_29564,N_24555);
nor UO_2582 (O_2582,N_25851,N_29777);
nand UO_2583 (O_2583,N_25444,N_22365);
nand UO_2584 (O_2584,N_24073,N_24875);
and UO_2585 (O_2585,N_20759,N_21435);
and UO_2586 (O_2586,N_20563,N_22001);
nor UO_2587 (O_2587,N_26184,N_25119);
nor UO_2588 (O_2588,N_27980,N_27725);
nand UO_2589 (O_2589,N_22543,N_23344);
nand UO_2590 (O_2590,N_20929,N_23912);
nor UO_2591 (O_2591,N_26183,N_23655);
xor UO_2592 (O_2592,N_24454,N_23374);
or UO_2593 (O_2593,N_27538,N_24334);
xor UO_2594 (O_2594,N_27666,N_20017);
xor UO_2595 (O_2595,N_29989,N_21201);
nand UO_2596 (O_2596,N_20262,N_27177);
or UO_2597 (O_2597,N_29345,N_23340);
nand UO_2598 (O_2598,N_25280,N_22991);
xnor UO_2599 (O_2599,N_25559,N_28843);
or UO_2600 (O_2600,N_20173,N_27546);
nand UO_2601 (O_2601,N_25872,N_27487);
or UO_2602 (O_2602,N_25172,N_24834);
nor UO_2603 (O_2603,N_22861,N_23118);
xnor UO_2604 (O_2604,N_24992,N_22404);
or UO_2605 (O_2605,N_25344,N_25013);
and UO_2606 (O_2606,N_26410,N_26505);
xor UO_2607 (O_2607,N_25414,N_26039);
nand UO_2608 (O_2608,N_27510,N_23624);
xnor UO_2609 (O_2609,N_27710,N_27433);
nand UO_2610 (O_2610,N_29180,N_23749);
or UO_2611 (O_2611,N_27415,N_23008);
nor UO_2612 (O_2612,N_28030,N_24660);
or UO_2613 (O_2613,N_21296,N_20288);
nor UO_2614 (O_2614,N_23135,N_29273);
nor UO_2615 (O_2615,N_22098,N_27945);
nor UO_2616 (O_2616,N_24344,N_29114);
xnor UO_2617 (O_2617,N_21748,N_21113);
xnor UO_2618 (O_2618,N_26152,N_22269);
nor UO_2619 (O_2619,N_24094,N_20202);
and UO_2620 (O_2620,N_23212,N_20009);
and UO_2621 (O_2621,N_20597,N_22369);
xnor UO_2622 (O_2622,N_20463,N_29805);
and UO_2623 (O_2623,N_24487,N_24773);
nor UO_2624 (O_2624,N_29288,N_25830);
nor UO_2625 (O_2625,N_28448,N_26204);
nand UO_2626 (O_2626,N_28013,N_24337);
nand UO_2627 (O_2627,N_23926,N_23030);
or UO_2628 (O_2628,N_26977,N_26726);
nand UO_2629 (O_2629,N_24987,N_21511);
or UO_2630 (O_2630,N_21725,N_29459);
nand UO_2631 (O_2631,N_20047,N_24162);
xor UO_2632 (O_2632,N_24363,N_21681);
nand UO_2633 (O_2633,N_28201,N_29957);
nand UO_2634 (O_2634,N_25804,N_28791);
nor UO_2635 (O_2635,N_22071,N_24356);
xnor UO_2636 (O_2636,N_27879,N_22993);
or UO_2637 (O_2637,N_29177,N_21437);
nor UO_2638 (O_2638,N_28190,N_23558);
nand UO_2639 (O_2639,N_23632,N_25098);
nand UO_2640 (O_2640,N_23208,N_22982);
nand UO_2641 (O_2641,N_27285,N_20584);
nand UO_2642 (O_2642,N_24451,N_25755);
and UO_2643 (O_2643,N_27215,N_23251);
and UO_2644 (O_2644,N_25485,N_26633);
xnor UO_2645 (O_2645,N_27815,N_28451);
nand UO_2646 (O_2646,N_21584,N_25360);
nor UO_2647 (O_2647,N_25710,N_24076);
and UO_2648 (O_2648,N_28202,N_26560);
and UO_2649 (O_2649,N_29635,N_28833);
or UO_2650 (O_2650,N_29528,N_22382);
nand UO_2651 (O_2651,N_21027,N_26267);
xnor UO_2652 (O_2652,N_23250,N_26939);
nand UO_2653 (O_2653,N_21851,N_26482);
xor UO_2654 (O_2654,N_20607,N_25393);
nor UO_2655 (O_2655,N_27591,N_22451);
xnor UO_2656 (O_2656,N_20824,N_27380);
nand UO_2657 (O_2657,N_21446,N_23797);
and UO_2658 (O_2658,N_28564,N_29616);
nand UO_2659 (O_2659,N_27044,N_23384);
or UO_2660 (O_2660,N_21636,N_29031);
or UO_2661 (O_2661,N_22657,N_21568);
or UO_2662 (O_2662,N_28887,N_23454);
and UO_2663 (O_2663,N_27560,N_22347);
nand UO_2664 (O_2664,N_24295,N_26695);
nand UO_2665 (O_2665,N_26455,N_25868);
xnor UO_2666 (O_2666,N_24726,N_25952);
nor UO_2667 (O_2667,N_23560,N_27259);
or UO_2668 (O_2668,N_28846,N_20492);
or UO_2669 (O_2669,N_22604,N_23973);
and UO_2670 (O_2670,N_28753,N_22733);
or UO_2671 (O_2671,N_23007,N_28640);
nor UO_2672 (O_2672,N_21195,N_23305);
and UO_2673 (O_2673,N_29996,N_27842);
nand UO_2674 (O_2674,N_25544,N_23111);
nand UO_2675 (O_2675,N_23565,N_26291);
nor UO_2676 (O_2676,N_26509,N_26681);
nand UO_2677 (O_2677,N_25816,N_27927);
or UO_2678 (O_2678,N_28834,N_21993);
nor UO_2679 (O_2679,N_27447,N_23139);
or UO_2680 (O_2680,N_24654,N_26625);
and UO_2681 (O_2681,N_27502,N_25640);
xor UO_2682 (O_2682,N_23726,N_25347);
and UO_2683 (O_2683,N_26524,N_27700);
nand UO_2684 (O_2684,N_22731,N_24938);
and UO_2685 (O_2685,N_26166,N_23667);
nor UO_2686 (O_2686,N_20541,N_20468);
nor UO_2687 (O_2687,N_29620,N_29366);
xor UO_2688 (O_2688,N_27003,N_22596);
xnor UO_2689 (O_2689,N_26141,N_21099);
xor UO_2690 (O_2690,N_29744,N_22936);
nand UO_2691 (O_2691,N_28698,N_23514);
or UO_2692 (O_2692,N_26279,N_29969);
nor UO_2693 (O_2693,N_22168,N_28297);
nand UO_2694 (O_2694,N_23537,N_20353);
xnor UO_2695 (O_2695,N_26248,N_26932);
and UO_2696 (O_2696,N_27429,N_21433);
or UO_2697 (O_2697,N_20808,N_23744);
nand UO_2698 (O_2698,N_24999,N_24475);
nand UO_2699 (O_2699,N_24656,N_29135);
or UO_2700 (O_2700,N_23670,N_28733);
nand UO_2701 (O_2701,N_28330,N_23363);
and UO_2702 (O_2702,N_28991,N_27745);
or UO_2703 (O_2703,N_29712,N_29387);
nor UO_2704 (O_2704,N_27049,N_25538);
nand UO_2705 (O_2705,N_26370,N_23218);
or UO_2706 (O_2706,N_26913,N_29038);
nand UO_2707 (O_2707,N_23937,N_23861);
nor UO_2708 (O_2708,N_26570,N_27703);
nor UO_2709 (O_2709,N_20656,N_20104);
or UO_2710 (O_2710,N_29851,N_20158);
or UO_2711 (O_2711,N_24319,N_22085);
nand UO_2712 (O_2712,N_28242,N_23798);
nand UO_2713 (O_2713,N_25949,N_23951);
nor UO_2714 (O_2714,N_22851,N_22745);
or UO_2715 (O_2715,N_26109,N_23512);
nor UO_2716 (O_2716,N_24546,N_24576);
and UO_2717 (O_2717,N_25898,N_23357);
and UO_2718 (O_2718,N_25334,N_25039);
xnor UO_2719 (O_2719,N_22901,N_25877);
nor UO_2720 (O_2720,N_20778,N_22146);
nand UO_2721 (O_2721,N_22219,N_22295);
nand UO_2722 (O_2722,N_20852,N_29465);
nor UO_2723 (O_2723,N_25833,N_25924);
xor UO_2724 (O_2724,N_26636,N_29679);
nand UO_2725 (O_2725,N_28965,N_25508);
nand UO_2726 (O_2726,N_22790,N_29497);
or UO_2727 (O_2727,N_21438,N_29199);
nand UO_2728 (O_2728,N_22735,N_28835);
and UO_2729 (O_2729,N_26086,N_24658);
and UO_2730 (O_2730,N_20253,N_26420);
xnor UO_2731 (O_2731,N_25917,N_27910);
nor UO_2732 (O_2732,N_24452,N_28960);
nor UO_2733 (O_2733,N_27110,N_28840);
nor UO_2734 (O_2734,N_26066,N_29983);
nor UO_2735 (O_2735,N_24336,N_22560);
xor UO_2736 (O_2736,N_27272,N_28966);
or UO_2737 (O_2737,N_24712,N_24391);
xor UO_2738 (O_2738,N_20837,N_23893);
nand UO_2739 (O_2739,N_24769,N_24715);
xor UO_2740 (O_2740,N_25732,N_24530);
or UO_2741 (O_2741,N_26690,N_22402);
nand UO_2742 (O_2742,N_22378,N_26281);
nand UO_2743 (O_2743,N_27930,N_29467);
or UO_2744 (O_2744,N_24545,N_22712);
xor UO_2745 (O_2745,N_23397,N_26743);
and UO_2746 (O_2746,N_20611,N_23287);
xor UO_2747 (O_2747,N_20109,N_25990);
and UO_2748 (O_2748,N_20545,N_20825);
xnor UO_2749 (O_2749,N_29455,N_23418);
and UO_2750 (O_2750,N_27836,N_23626);
xor UO_2751 (O_2751,N_26096,N_21043);
or UO_2752 (O_2752,N_21503,N_26871);
xor UO_2753 (O_2753,N_27637,N_27015);
and UO_2754 (O_2754,N_28291,N_24109);
or UO_2755 (O_2755,N_22035,N_25242);
nand UO_2756 (O_2756,N_28173,N_24198);
xnor UO_2757 (O_2757,N_29930,N_24776);
and UO_2758 (O_2758,N_20324,N_22372);
nor UO_2759 (O_2759,N_20199,N_29011);
nand UO_2760 (O_2760,N_23829,N_28156);
nor UO_2761 (O_2761,N_24587,N_26480);
and UO_2762 (O_2762,N_29505,N_20960);
xnor UO_2763 (O_2763,N_29610,N_20794);
or UO_2764 (O_2764,N_21684,N_24019);
nor UO_2765 (O_2765,N_27140,N_28949);
and UO_2766 (O_2766,N_24644,N_25225);
nand UO_2767 (O_2767,N_21954,N_21263);
nor UO_2768 (O_2768,N_26273,N_26864);
nor UO_2769 (O_2769,N_26161,N_24813);
nand UO_2770 (O_2770,N_27071,N_22246);
or UO_2771 (O_2771,N_25647,N_22123);
or UO_2772 (O_2772,N_29702,N_22634);
nor UO_2773 (O_2773,N_24501,N_20259);
and UO_2774 (O_2774,N_21217,N_28094);
nor UO_2775 (O_2775,N_20900,N_25452);
or UO_2776 (O_2776,N_23010,N_28748);
and UO_2777 (O_2777,N_26669,N_22566);
xor UO_2778 (O_2778,N_23818,N_28934);
nor UO_2779 (O_2779,N_28756,N_28801);
nand UO_2780 (O_2780,N_24013,N_29766);
nor UO_2781 (O_2781,N_24569,N_23133);
xor UO_2782 (O_2782,N_28296,N_27332);
nand UO_2783 (O_2783,N_25048,N_29166);
nand UO_2784 (O_2784,N_28701,N_25459);
xor UO_2785 (O_2785,N_22753,N_28389);
xor UO_2786 (O_2786,N_21622,N_29704);
nand UO_2787 (O_2787,N_20279,N_20320);
nand UO_2788 (O_2788,N_20283,N_29832);
nor UO_2789 (O_2789,N_20508,N_27760);
or UO_2790 (O_2790,N_26216,N_24663);
and UO_2791 (O_2791,N_21881,N_27850);
xnor UO_2792 (O_2792,N_25714,N_27946);
nor UO_2793 (O_2793,N_29769,N_22462);
nor UO_2794 (O_2794,N_26764,N_23529);
nor UO_2795 (O_2795,N_24762,N_25466);
nor UO_2796 (O_2796,N_26092,N_21617);
nor UO_2797 (O_2797,N_27055,N_26642);
xnor UO_2798 (O_2798,N_20080,N_22259);
and UO_2799 (O_2799,N_29807,N_21544);
or UO_2800 (O_2800,N_22313,N_29947);
xor UO_2801 (O_2801,N_27364,N_27461);
nand UO_2802 (O_2802,N_23277,N_28271);
or UO_2803 (O_2803,N_26873,N_26347);
nor UO_2804 (O_2804,N_25420,N_28726);
xor UO_2805 (O_2805,N_21370,N_27050);
or UO_2806 (O_2806,N_21666,N_23896);
or UO_2807 (O_2807,N_25267,N_29145);
nor UO_2808 (O_2808,N_21318,N_27187);
nand UO_2809 (O_2809,N_25847,N_27174);
nand UO_2810 (O_2810,N_20829,N_28782);
nor UO_2811 (O_2811,N_24144,N_21862);
nand UO_2812 (O_2812,N_26967,N_23836);
and UO_2813 (O_2813,N_22279,N_27575);
nor UO_2814 (O_2814,N_21030,N_28427);
nand UO_2815 (O_2815,N_27394,N_29663);
or UO_2816 (O_2816,N_23349,N_26180);
nand UO_2817 (O_2817,N_20476,N_25175);
or UO_2818 (O_2818,N_23226,N_22795);
or UO_2819 (O_2819,N_21547,N_21104);
and UO_2820 (O_2820,N_24713,N_23877);
and UO_2821 (O_2821,N_25666,N_26928);
or UO_2822 (O_2822,N_21593,N_27368);
or UO_2823 (O_2823,N_25244,N_27471);
nor UO_2824 (O_2824,N_27504,N_20229);
nand UO_2825 (O_2825,N_20115,N_29347);
xnor UO_2826 (O_2826,N_22106,N_22286);
and UO_2827 (O_2827,N_29578,N_20116);
nor UO_2828 (O_2828,N_25900,N_29160);
and UO_2829 (O_2829,N_27917,N_23678);
nor UO_2830 (O_2830,N_24634,N_24001);
xor UO_2831 (O_2831,N_23969,N_22867);
xnor UO_2832 (O_2832,N_20165,N_20185);
or UO_2833 (O_2833,N_22053,N_25852);
and UO_2834 (O_2834,N_25912,N_25796);
nand UO_2835 (O_2835,N_22719,N_28222);
nand UO_2836 (O_2836,N_28060,N_29600);
xnor UO_2837 (O_2837,N_24395,N_22396);
xnor UO_2838 (O_2838,N_22333,N_22243);
xor UO_2839 (O_2839,N_20511,N_27792);
nand UO_2840 (O_2840,N_28039,N_28803);
or UO_2841 (O_2841,N_29051,N_28470);
or UO_2842 (O_2842,N_23656,N_29767);
nand UO_2843 (O_2843,N_21390,N_23387);
nand UO_2844 (O_2844,N_20248,N_28028);
nand UO_2845 (O_2845,N_26225,N_21738);
nor UO_2846 (O_2846,N_24832,N_27766);
xor UO_2847 (O_2847,N_28608,N_25339);
xor UO_2848 (O_2848,N_25584,N_29646);
xnor UO_2849 (O_2849,N_28747,N_26545);
nand UO_2850 (O_2850,N_28261,N_21882);
nand UO_2851 (O_2851,N_22924,N_28705);
and UO_2852 (O_2852,N_27872,N_20296);
or UO_2853 (O_2853,N_29973,N_26628);
and UO_2854 (O_2854,N_28283,N_28710);
nand UO_2855 (O_2855,N_24168,N_20539);
nand UO_2856 (O_2856,N_26312,N_22012);
or UO_2857 (O_2857,N_22674,N_23056);
nand UO_2858 (O_2858,N_28735,N_21357);
nand UO_2859 (O_2859,N_26255,N_20812);
or UO_2860 (O_2860,N_27133,N_26030);
xor UO_2861 (O_2861,N_28169,N_24071);
or UO_2862 (O_2862,N_20814,N_24876);
nand UO_2863 (O_2863,N_29074,N_22626);
and UO_2864 (O_2864,N_22746,N_21505);
nand UO_2865 (O_2865,N_29797,N_21897);
nor UO_2866 (O_2866,N_25836,N_29763);
xor UO_2867 (O_2867,N_21384,N_20701);
nor UO_2868 (O_2868,N_29742,N_25194);
nand UO_2869 (O_2869,N_23369,N_23851);
nor UO_2870 (O_2870,N_20995,N_28684);
or UO_2871 (O_2871,N_20411,N_21934);
nor UO_2872 (O_2872,N_21247,N_27086);
nor UO_2873 (O_2873,N_23043,N_20981);
or UO_2874 (O_2874,N_23229,N_25961);
nand UO_2875 (O_2875,N_29466,N_27250);
or UO_2876 (O_2876,N_29834,N_29357);
and UO_2877 (O_2877,N_27438,N_21422);
xor UO_2878 (O_2878,N_29007,N_25075);
nand UO_2879 (O_2879,N_29593,N_22488);
nor UO_2880 (O_2880,N_21860,N_25090);
nand UO_2881 (O_2881,N_23718,N_27984);
and UO_2882 (O_2882,N_25678,N_23648);
or UO_2883 (O_2883,N_21034,N_23358);
nor UO_2884 (O_2884,N_28679,N_23827);
and UO_2885 (O_2885,N_20475,N_21757);
xor UO_2886 (O_2886,N_23765,N_28638);
nand UO_2887 (O_2887,N_22671,N_21510);
xor UO_2888 (O_2888,N_29858,N_25623);
or UO_2889 (O_2889,N_22694,N_26814);
nor UO_2890 (O_2890,N_24792,N_25856);
nor UO_2891 (O_2891,N_22651,N_22398);
nand UO_2892 (O_2892,N_23345,N_24474);
or UO_2893 (O_2893,N_20843,N_29840);
and UO_2894 (O_2894,N_26603,N_26987);
xnor UO_2895 (O_2895,N_28180,N_25073);
xor UO_2896 (O_2896,N_23759,N_20720);
nand UO_2897 (O_2897,N_26005,N_23499);
nor UO_2898 (O_2898,N_26980,N_20630);
and UO_2899 (O_2899,N_25556,N_23399);
xor UO_2900 (O_2900,N_21540,N_20737);
nor UO_2901 (O_2901,N_28452,N_21669);
xor UO_2902 (O_2902,N_25570,N_23315);
or UO_2903 (O_2903,N_21760,N_24415);
nor UO_2904 (O_2904,N_21922,N_25316);
xor UO_2905 (O_2905,N_24847,N_22629);
and UO_2906 (O_2906,N_26671,N_25908);
nor UO_2907 (O_2907,N_22606,N_26097);
and UO_2908 (O_2908,N_24929,N_20638);
and UO_2909 (O_2909,N_26268,N_23244);
nor UO_2910 (O_2910,N_26390,N_26133);
xor UO_2911 (O_2911,N_24224,N_27749);
or UO_2912 (O_2912,N_27659,N_20060);
nand UO_2913 (O_2913,N_21536,N_20834);
nand UO_2914 (O_2914,N_26442,N_21580);
nand UO_2915 (O_2915,N_24785,N_22236);
nand UO_2916 (O_2916,N_22569,N_21325);
xor UO_2917 (O_2917,N_26812,N_26069);
xnor UO_2918 (O_2918,N_29222,N_29349);
nor UO_2919 (O_2919,N_21972,N_20542);
nand UO_2920 (O_2920,N_22390,N_26978);
nand UO_2921 (O_2921,N_26250,N_20467);
or UO_2922 (O_2922,N_24082,N_23944);
and UO_2923 (O_2923,N_23154,N_29066);
or UO_2924 (O_2924,N_22792,N_27937);
nor UO_2925 (O_2925,N_26503,N_22405);
and UO_2926 (O_2926,N_23165,N_26164);
and UO_2927 (O_2927,N_28837,N_22163);
nor UO_2928 (O_2928,N_25153,N_24665);
and UO_2929 (O_2929,N_27247,N_24453);
xnor UO_2930 (O_2930,N_29240,N_29428);
xnor UO_2931 (O_2931,N_29103,N_26156);
nand UO_2932 (O_2932,N_27991,N_29358);
and UO_2933 (O_2933,N_27351,N_20753);
nor UO_2934 (O_2934,N_29496,N_29835);
nand UO_2935 (O_2935,N_27243,N_26645);
and UO_2936 (O_2936,N_25424,N_29296);
and UO_2937 (O_2937,N_21589,N_26960);
nor UO_2938 (O_2938,N_24043,N_21658);
or UO_2939 (O_2939,N_29298,N_21308);
nor UO_2940 (O_2940,N_22256,N_25910);
nor UO_2941 (O_2941,N_22434,N_29750);
xor UO_2942 (O_2942,N_25014,N_29220);
nand UO_2943 (O_2943,N_23102,N_25926);
nor UO_2944 (O_2944,N_27012,N_21483);
nand UO_2945 (O_2945,N_23062,N_22643);
nor UO_2946 (O_2946,N_25800,N_23881);
nand UO_2947 (O_2947,N_20228,N_29405);
nor UO_2948 (O_2948,N_20647,N_29698);
nor UO_2949 (O_2949,N_25946,N_25078);
xnor UO_2950 (O_2950,N_25945,N_26084);
xor UO_2951 (O_2951,N_27979,N_24699);
and UO_2952 (O_2952,N_27664,N_29838);
and UO_2953 (O_2953,N_26175,N_28807);
nand UO_2954 (O_2954,N_21129,N_20876);
and UO_2955 (O_2955,N_23037,N_21315);
nand UO_2956 (O_2956,N_23350,N_21402);
and UO_2957 (O_2957,N_27278,N_28044);
xor UO_2958 (O_2958,N_29680,N_21736);
nor UO_2959 (O_2959,N_21133,N_23803);
nand UO_2960 (O_2960,N_20377,N_23546);
xnor UO_2961 (O_2961,N_29373,N_21229);
nand UO_2962 (O_2962,N_27624,N_28102);
and UO_2963 (O_2963,N_23761,N_21709);
nor UO_2964 (O_2964,N_23762,N_29086);
nor UO_2965 (O_2965,N_24418,N_23935);
nor UO_2966 (O_2966,N_20883,N_29703);
xor UO_2967 (O_2967,N_28373,N_28075);
or UO_2968 (O_2968,N_26261,N_27181);
nor UO_2969 (O_2969,N_23796,N_24639);
nand UO_2970 (O_2970,N_22902,N_25022);
and UO_2971 (O_2971,N_26738,N_21313);
nor UO_2972 (O_2972,N_20216,N_27511);
nand UO_2973 (O_2973,N_24862,N_26445);
or UO_2974 (O_2974,N_21842,N_29872);
or UO_2975 (O_2975,N_21116,N_21959);
xor UO_2976 (O_2976,N_27563,N_20905);
and UO_2977 (O_2977,N_24677,N_28391);
nand UO_2978 (O_2978,N_24705,N_22082);
nand UO_2979 (O_2979,N_21271,N_25759);
and UO_2980 (O_2980,N_23701,N_22495);
nand UO_2981 (O_2981,N_29768,N_20987);
and UO_2982 (O_2982,N_22044,N_21711);
or UO_2983 (O_2983,N_29404,N_27362);
and UO_2984 (O_2984,N_27697,N_27207);
xnor UO_2985 (O_2985,N_20314,N_26284);
and UO_2986 (O_2986,N_29403,N_24920);
nand UO_2987 (O_2987,N_20836,N_28744);
nor UO_2988 (O_2988,N_26891,N_27008);
and UO_2989 (O_2989,N_20567,N_28303);
and UO_2990 (O_2990,N_20260,N_21809);
or UO_2991 (O_2991,N_22931,N_28757);
nand UO_2992 (O_2992,N_29264,N_20819);
nor UO_2993 (O_2993,N_26599,N_28889);
and UO_2994 (O_2994,N_25260,N_24134);
and UO_2995 (O_2995,N_23372,N_27066);
nor UO_2996 (O_2996,N_28693,N_25016);
nand UO_2997 (O_2997,N_22026,N_26766);
or UO_2998 (O_2998,N_28874,N_25679);
nor UO_2999 (O_2999,N_29811,N_23443);
nand UO_3000 (O_3000,N_28132,N_28056);
and UO_3001 (O_3001,N_26701,N_20828);
nand UO_3002 (O_3002,N_24979,N_23198);
nand UO_3003 (O_3003,N_21700,N_25882);
or UO_3004 (O_3004,N_24867,N_21444);
nor UO_3005 (O_3005,N_25858,N_21988);
xor UO_3006 (O_3006,N_28088,N_24597);
nand UO_3007 (O_3007,N_25683,N_22608);
nand UO_3008 (O_3008,N_23681,N_22615);
xor UO_3009 (O_3009,N_23553,N_23644);
nor UO_3010 (O_3010,N_24228,N_25994);
and UO_3011 (O_3011,N_27073,N_29901);
and UO_3012 (O_3012,N_21861,N_29588);
and UO_3013 (O_3013,N_25891,N_21199);
nand UO_3014 (O_3014,N_28956,N_21393);
nor UO_3015 (O_3015,N_20717,N_20962);
and UO_3016 (O_3016,N_21586,N_21385);
and UO_3017 (O_3017,N_22316,N_24183);
and UO_3018 (O_3018,N_21220,N_22866);
or UO_3019 (O_3019,N_29612,N_28224);
nand UO_3020 (O_3020,N_23334,N_25000);
nand UO_3021 (O_3021,N_28436,N_20693);
xor UO_3022 (O_3022,N_23317,N_23858);
nor UO_3023 (O_3023,N_27943,N_28911);
or UO_3024 (O_3024,N_21909,N_22837);
nand UO_3025 (O_3025,N_26232,N_20965);
and UO_3026 (O_3026,N_20820,N_26902);
or UO_3027 (O_3027,N_26007,N_26226);
nor UO_3028 (O_3028,N_29693,N_22858);
or UO_3029 (O_3029,N_29822,N_26436);
xor UO_3030 (O_3030,N_29756,N_24517);
nand UO_3031 (O_3031,N_26594,N_24753);
nand UO_3032 (O_3032,N_22913,N_20421);
xor UO_3033 (O_3033,N_27304,N_21398);
xnor UO_3034 (O_3034,N_20334,N_26674);
xnor UO_3035 (O_3035,N_22229,N_22479);
and UO_3036 (O_3036,N_22094,N_22675);
or UO_3037 (O_3037,N_24598,N_27514);
nand UO_3038 (O_3038,N_28347,N_28375);
and UO_3039 (O_3039,N_23673,N_24276);
and UO_3040 (O_3040,N_24285,N_25250);
and UO_3041 (O_3041,N_21815,N_29573);
nor UO_3042 (O_3042,N_29696,N_21808);
and UO_3043 (O_3043,N_20274,N_28626);
or UO_3044 (O_3044,N_29239,N_20517);
or UO_3045 (O_3045,N_28997,N_21416);
nor UO_3046 (O_3046,N_20784,N_23945);
or UO_3047 (O_3047,N_28560,N_25236);
or UO_3048 (O_3048,N_28561,N_21868);
and UO_3049 (O_3049,N_21038,N_20400);
or UO_3050 (O_3050,N_21063,N_27178);
xnor UO_3051 (O_3051,N_28909,N_24197);
nand UO_3052 (O_3052,N_22767,N_29825);
xor UO_3053 (O_3053,N_29829,N_22348);
or UO_3054 (O_3054,N_20106,N_24111);
or UO_3055 (O_3055,N_27683,N_23213);
or UO_3056 (O_3056,N_29352,N_21962);
nand UO_3057 (O_3057,N_27470,N_20894);
xor UO_3058 (O_3058,N_22992,N_20232);
or UO_3059 (O_3059,N_21428,N_23989);
nand UO_3060 (O_3060,N_23968,N_21061);
nand UO_3061 (O_3061,N_26710,N_21573);
xnor UO_3062 (O_3062,N_21971,N_21566);
nor UO_3063 (O_3063,N_28367,N_21719);
nand UO_3064 (O_3064,N_28051,N_27607);
or UO_3065 (O_3065,N_27528,N_29119);
nor UO_3066 (O_3066,N_28408,N_26819);
xor UO_3067 (O_3067,N_26194,N_24278);
xor UO_3068 (O_3068,N_28893,N_20461);
nand UO_3069 (O_3069,N_24827,N_29731);
nor UO_3070 (O_3070,N_27269,N_29786);
and UO_3071 (O_3071,N_21638,N_21880);
xor UO_3072 (O_3072,N_25783,N_29028);
xnor UO_3073 (O_3073,N_21923,N_26082);
xnor UO_3074 (O_3074,N_25158,N_22520);
xnor UO_3075 (O_3075,N_21474,N_25976);
nor UO_3076 (O_3076,N_28600,N_20801);
or UO_3077 (O_3077,N_26857,N_20337);
or UO_3078 (O_3078,N_28819,N_20418);
and UO_3079 (O_3079,N_25151,N_27006);
or UO_3080 (O_3080,N_23032,N_26543);
nor UO_3081 (O_3081,N_25171,N_25270);
nor UO_3082 (O_3082,N_28492,N_21745);
and UO_3083 (O_3083,N_28462,N_24770);
nand UO_3084 (O_3084,N_28042,N_22125);
xor UO_3085 (O_3085,N_20755,N_28016);
or UO_3086 (O_3086,N_22939,N_22471);
nand UO_3087 (O_3087,N_27335,N_22054);
and UO_3088 (O_3088,N_23707,N_25342);
nor UO_3089 (O_3089,N_24405,N_27031);
xnor UO_3090 (O_3090,N_27601,N_23717);
or UO_3091 (O_3091,N_27831,N_21621);
and UO_3092 (O_3092,N_27752,N_23435);
or UO_3093 (O_3093,N_20811,N_22210);
and UO_3094 (O_3094,N_29627,N_24777);
nand UO_3095 (O_3095,N_25769,N_27387);
and UO_3096 (O_3096,N_27539,N_20313);
nor UO_3097 (O_3097,N_22034,N_23595);
and UO_3098 (O_3098,N_23573,N_27890);
and UO_3099 (O_3099,N_22305,N_21279);
or UO_3100 (O_3100,N_26108,N_26725);
nor UO_3101 (O_3101,N_21828,N_21334);
xor UO_3102 (O_3102,N_23590,N_25626);
or UO_3103 (O_3103,N_26813,N_21668);
xnor UO_3104 (O_3104,N_28126,N_22364);
and UO_3105 (O_3105,N_22669,N_28866);
nand UO_3106 (O_3106,N_26647,N_20888);
nand UO_3107 (O_3107,N_28510,N_28816);
xor UO_3108 (O_3108,N_26955,N_27553);
xor UO_3109 (O_3109,N_21473,N_20871);
xnor UO_3110 (O_3110,N_25825,N_24731);
nand UO_3111 (O_3111,N_28245,N_20350);
or UO_3112 (O_3112,N_23523,N_25886);
nor UO_3113 (O_3113,N_24593,N_24852);
and UO_3114 (O_3114,N_22174,N_27559);
xnor UO_3115 (O_3115,N_28343,N_22892);
and UO_3116 (O_3116,N_27581,N_25921);
xor UO_3117 (O_3117,N_23599,N_26177);
xnor UO_3118 (O_3118,N_28080,N_28441);
nor UO_3119 (O_3119,N_25651,N_24000);
nor UO_3120 (O_3120,N_27859,N_27421);
nor UO_3121 (O_3121,N_25255,N_28789);
or UO_3122 (O_3122,N_20940,N_25782);
nor UO_3123 (O_3123,N_20268,N_23234);
xor UO_3124 (O_3124,N_22475,N_26722);
and UO_3125 (O_3125,N_28225,N_23024);
or UO_3126 (O_3126,N_20585,N_26203);
and UO_3127 (O_3127,N_25659,N_28649);
and UO_3128 (O_3128,N_24126,N_26046);
and UO_3129 (O_3129,N_29108,N_22764);
nand UO_3130 (O_3130,N_25906,N_21323);
nand UO_3131 (O_3131,N_21181,N_20687);
xor UO_3132 (O_3132,N_26447,N_20380);
nand UO_3133 (O_3133,N_24804,N_29651);
nor UO_3134 (O_3134,N_20290,N_20864);
nand UO_3135 (O_3135,N_20986,N_21233);
and UO_3136 (O_3136,N_21603,N_28435);
nor UO_3137 (O_3137,N_24422,N_25718);
nor UO_3138 (O_3138,N_24600,N_27449);
and UO_3139 (O_3139,N_29892,N_25402);
nand UO_3140 (O_3140,N_25409,N_29426);
or UO_3141 (O_3141,N_24851,N_21814);
nor UO_3142 (O_3142,N_27124,N_23752);
and UO_3143 (O_3143,N_29607,N_24627);
nor UO_3144 (O_3144,N_26286,N_24214);
and UO_3145 (O_3145,N_28870,N_20438);
nand UO_3146 (O_3146,N_29171,N_22160);
nand UO_3147 (O_3147,N_26117,N_22721);
xor UO_3148 (O_3148,N_23598,N_26311);
xnor UO_3149 (O_3149,N_27200,N_21087);
and UO_3150 (O_3150,N_28193,N_27357);
or UO_3151 (O_3151,N_29713,N_25571);
nor UO_3152 (O_3152,N_28341,N_28946);
nand UO_3153 (O_3153,N_26415,N_26434);
and UO_3154 (O_3154,N_23713,N_23143);
nor UO_3155 (O_3155,N_21986,N_21967);
xnor UO_3156 (O_3156,N_20252,N_21262);
nand UO_3157 (O_3157,N_27498,N_29975);
nor UO_3158 (O_3158,N_26134,N_27566);
nor UO_3159 (O_3159,N_27112,N_29262);
nor UO_3160 (O_3160,N_21423,N_20618);
and UO_3161 (O_3161,N_24287,N_20167);
and UO_3162 (O_3162,N_29948,N_20254);
xnor UO_3163 (O_3163,N_28792,N_29186);
xor UO_3164 (O_3164,N_23936,N_24565);
nand UO_3165 (O_3165,N_29228,N_27136);
xnor UO_3166 (O_3166,N_27708,N_27347);
xnor UO_3167 (O_3167,N_24905,N_25132);
xnor UO_3168 (O_3168,N_21202,N_24088);
nor UO_3169 (O_3169,N_21467,N_22344);
and UO_3170 (O_3170,N_26259,N_22113);
nor UO_3171 (O_3171,N_29391,N_25723);
or UO_3172 (O_3172,N_20344,N_26581);
nor UO_3173 (O_3173,N_24489,N_28516);
or UO_3174 (O_3174,N_20220,N_22149);
or UO_3175 (O_3175,N_21891,N_24167);
nor UO_3176 (O_3176,N_27416,N_22893);
nand UO_3177 (O_3177,N_26580,N_24655);
xor UO_3178 (O_3178,N_22550,N_28794);
nor UO_3179 (O_3179,N_28955,N_25878);
xnor UO_3180 (O_3180,N_24744,N_24614);
xnor UO_3181 (O_3181,N_27735,N_24548);
and UO_3182 (O_3182,N_26371,N_27217);
or UO_3183 (O_3183,N_22079,N_29401);
nand UO_3184 (O_3184,N_29258,N_27561);
xnor UO_3185 (O_3185,N_26965,N_23786);
nand UO_3186 (O_3186,N_26199,N_28585);
nor UO_3187 (O_3187,N_20583,N_28454);
or UO_3188 (O_3188,N_23140,N_22816);
and UO_3189 (O_3189,N_22296,N_25844);
xnor UO_3190 (O_3190,N_23409,N_25775);
and UO_3191 (O_3191,N_25705,N_24642);
nand UO_3192 (O_3192,N_20764,N_24819);
nor UO_3193 (O_3193,N_22361,N_24471);
or UO_3194 (O_3194,N_24710,N_21376);
or UO_3195 (O_3195,N_21183,N_22945);
nand UO_3196 (O_3196,N_29351,N_25279);
nand UO_3197 (O_3197,N_28565,N_21674);
nand UO_3198 (O_3198,N_29487,N_27037);
nand UO_3199 (O_3199,N_22812,N_29808);
and UO_3200 (O_3200,N_26843,N_22429);
nand UO_3201 (O_3201,N_24696,N_23834);
or UO_3202 (O_3202,N_25272,N_28336);
xor UO_3203 (O_3203,N_20203,N_26111);
or UO_3204 (O_3204,N_24884,N_21284);
nor UO_3205 (O_3205,N_26334,N_24955);
nor UO_3206 (O_3206,N_25806,N_23210);
xnor UO_3207 (O_3207,N_22809,N_29388);
nand UO_3208 (O_3208,N_20785,N_27845);
nand UO_3209 (O_3209,N_28824,N_24470);
and UO_3210 (O_3210,N_25756,N_24927);
xor UO_3211 (O_3211,N_27231,N_23842);
or UO_3212 (O_3212,N_21408,N_20072);
and UO_3213 (O_3213,N_25333,N_27305);
nor UO_3214 (O_3214,N_24960,N_26890);
xor UO_3215 (O_3215,N_20917,N_22984);
and UO_3216 (O_3216,N_20319,N_25085);
or UO_3217 (O_3217,N_21153,N_21248);
xnor UO_3218 (O_3218,N_25312,N_23038);
nor UO_3219 (O_3219,N_26246,N_21847);
or UO_3220 (O_3220,N_26386,N_27669);
or UO_3221 (O_3221,N_24510,N_29987);
or UO_3222 (O_3222,N_23403,N_23696);
xor UO_3223 (O_3223,N_22133,N_24877);
or UO_3224 (O_3224,N_23576,N_21231);
xor UO_3225 (O_3225,N_20412,N_29393);
nor UO_3226 (O_3226,N_20058,N_26145);
nand UO_3227 (O_3227,N_20257,N_29281);
or UO_3228 (O_3228,N_20543,N_27928);
nor UO_3229 (O_3229,N_28317,N_24209);
or UO_3230 (O_3230,N_29215,N_20771);
xnor UO_3231 (O_3231,N_27736,N_21908);
nand UO_3232 (O_3232,N_20533,N_27914);
and UO_3233 (O_3233,N_29474,N_29883);
or UO_3234 (O_3234,N_27021,N_23232);
xor UO_3235 (O_3235,N_25750,N_29208);
and UO_3236 (O_3236,N_25361,N_29793);
nor UO_3237 (O_3237,N_25019,N_27041);
nand UO_3238 (O_3238,N_24729,N_20375);
nor UO_3239 (O_3239,N_24799,N_20621);
nand UO_3240 (O_3240,N_28128,N_21574);
or UO_3241 (O_3241,N_29617,N_21235);
nor UO_3242 (O_3242,N_20293,N_21260);
nor UO_3243 (O_3243,N_27896,N_26325);
xnor UO_3244 (O_3244,N_27714,N_26630);
nor UO_3245 (O_3245,N_29275,N_20849);
xnor UO_3246 (O_3246,N_25170,N_22453);
xnor UO_3247 (O_3247,N_23205,N_26275);
nand UO_3248 (O_3248,N_28754,N_20178);
and UO_3249 (O_3249,N_22198,N_26048);
or UO_3250 (O_3250,N_28603,N_25521);
nor UO_3251 (O_3251,N_27620,N_24881);
xor UO_3252 (O_3252,N_21635,N_29734);
nand UO_3253 (O_3253,N_23921,N_23597);
xor UO_3254 (O_3254,N_23230,N_20146);
and UO_3255 (O_3255,N_27771,N_24202);
nor UO_3256 (O_3256,N_25840,N_27670);
and UO_3257 (O_3257,N_21189,N_26167);
or UO_3258 (O_3258,N_24237,N_28275);
and UO_3259 (O_3259,N_28179,N_22786);
and UO_3260 (O_3260,N_24515,N_29453);
nor UO_3261 (O_3261,N_21903,N_22602);
and UO_3262 (O_3262,N_27355,N_23067);
and UO_3263 (O_3263,N_27512,N_22644);
and UO_3264 (O_3264,N_26761,N_23457);
nor UO_3265 (O_3265,N_29123,N_27109);
nor UO_3266 (O_3266,N_26870,N_21781);
nor UO_3267 (O_3267,N_25512,N_22765);
and UO_3268 (O_3268,N_25343,N_24786);
and UO_3269 (O_3269,N_29024,N_27246);
and UO_3270 (O_3270,N_26605,N_21744);
and UO_3271 (O_3271,N_24461,N_27781);
nand UO_3272 (O_3272,N_29000,N_27864);
xor UO_3273 (O_3273,N_23089,N_26153);
xnor UO_3274 (O_3274,N_22171,N_29984);
nor UO_3275 (O_3275,N_22189,N_22903);
nor UO_3276 (O_3276,N_26131,N_29340);
nor UO_3277 (O_3277,N_26719,N_29146);
xnor UO_3278 (O_3278,N_27060,N_22872);
xor UO_3279 (O_3279,N_21012,N_20570);
xnor UO_3280 (O_3280,N_20162,N_24523);
or UO_3281 (O_3281,N_26063,N_27120);
nand UO_3282 (O_3282,N_21703,N_28504);
xnor UO_3283 (O_3283,N_22766,N_23410);
nand UO_3284 (O_3284,N_23902,N_25784);
nand UO_3285 (O_3285,N_21777,N_23773);
or UO_3286 (O_3286,N_26391,N_24797);
nor UO_3287 (O_3287,N_20281,N_25030);
nand UO_3288 (O_3288,N_23764,N_26734);
nand UO_3289 (O_3289,N_24910,N_23002);
nor UO_3290 (O_3290,N_27507,N_24709);
and UO_3291 (O_3291,N_29810,N_27413);
and UO_3292 (O_3292,N_23817,N_26736);
or UO_3293 (O_3293,N_24571,N_26882);
and UO_3294 (O_3294,N_25274,N_26784);
xor UO_3295 (O_3295,N_28091,N_20298);
or UO_3296 (O_3296,N_26788,N_29506);
or UO_3297 (O_3297,N_22747,N_24608);
and UO_3298 (O_3298,N_20670,N_29849);
and UO_3299 (O_3299,N_20143,N_28895);
and UO_3300 (O_3300,N_24472,N_24619);
nor UO_3301 (O_3301,N_23801,N_23526);
and UO_3302 (O_3302,N_26100,N_29844);
or UO_3303 (O_3303,N_23086,N_20069);
nand UO_3304 (O_3304,N_24774,N_24226);
xor UO_3305 (O_3305,N_26210,N_24828);
xor UO_3306 (O_3306,N_27599,N_29856);
or UO_3307 (O_3307,N_27463,N_27985);
or UO_3308 (O_3308,N_29790,N_21822);
xor UO_3309 (O_3309,N_21737,N_25603);
and UO_3310 (O_3310,N_26990,N_20855);
nor UO_3311 (O_3311,N_23029,N_29362);
and UO_3312 (O_3312,N_26504,N_20580);
or UO_3313 (O_3313,N_29508,N_22743);
nand UO_3314 (O_3314,N_29938,N_26894);
nand UO_3315 (O_3315,N_26304,N_26191);
xnor UO_3316 (O_3316,N_26697,N_20227);
nor UO_3317 (O_3317,N_29727,N_24898);
or UO_3318 (O_3318,N_27579,N_24063);
or UO_3319 (O_3319,N_20910,N_29317);
xnor UO_3320 (O_3320,N_27882,N_29041);
xnor UO_3321 (O_3321,N_27035,N_21740);
nor UO_3322 (O_3322,N_27986,N_29469);
or UO_3323 (O_3323,N_24605,N_27254);
nand UO_3324 (O_3324,N_27307,N_28982);
nand UO_3325 (O_3325,N_22855,N_28507);
or UO_3326 (O_3326,N_26463,N_24698);
xnor UO_3327 (O_3327,N_20102,N_24860);
or UO_3328 (O_3328,N_28355,N_24485);
nand UO_3329 (O_3329,N_29757,N_25744);
nor UO_3330 (O_3330,N_24072,N_28421);
nor UO_3331 (O_3331,N_28438,N_23063);
nor UO_3332 (O_3332,N_25960,N_23909);
or UO_3333 (O_3333,N_26425,N_21553);
or UO_3334 (O_3334,N_26394,N_24940);
nor UO_3335 (O_3335,N_27218,N_24885);
nor UO_3336 (O_3336,N_21161,N_21178);
nor UO_3337 (O_3337,N_25611,N_27650);
or UO_3338 (O_3338,N_22111,N_27431);
nor UO_3339 (O_3339,N_26733,N_29163);
or UO_3340 (O_3340,N_25823,N_28722);
nand UO_3341 (O_3341,N_27621,N_26119);
nand UO_3342 (O_3342,N_29077,N_28093);
and UO_3343 (O_3343,N_29138,N_20359);
nand UO_3344 (O_3344,N_21671,N_26215);
nand UO_3345 (O_3345,N_21250,N_26257);
xor UO_3346 (O_3346,N_21317,N_27934);
nor UO_3347 (O_3347,N_21324,N_26349);
and UO_3348 (O_3348,N_25288,N_26085);
nand UO_3349 (O_3349,N_28878,N_25253);
and UO_3350 (O_3350,N_22140,N_27800);
xor UO_3351 (O_3351,N_20766,N_27741);
and UO_3352 (O_3352,N_29843,N_28276);
and UO_3353 (O_3353,N_25015,N_22577);
nor UO_3354 (O_3354,N_26537,N_20502);
xor UO_3355 (O_3355,N_24683,N_28468);
or UO_3356 (O_3356,N_25259,N_21126);
nand UO_3357 (O_3357,N_20370,N_29394);
nand UO_3358 (O_3358,N_24572,N_29439);
nor UO_3359 (O_3359,N_22672,N_24136);
nor UO_3360 (O_3360,N_26351,N_21741);
or UO_3361 (O_3361,N_25296,N_20357);
or UO_3362 (O_3362,N_25724,N_25515);
xnor UO_3363 (O_3363,N_29457,N_20018);
and UO_3364 (O_3364,N_25293,N_27627);
and UO_3365 (O_3365,N_21596,N_27672);
xor UO_3366 (O_3366,N_22639,N_29836);
nor UO_3367 (O_3367,N_25103,N_24869);
nand UO_3368 (O_3368,N_28267,N_28123);
and UO_3369 (O_3369,N_20842,N_25876);
and UO_3370 (O_3370,N_26583,N_25320);
and UO_3371 (O_3371,N_22354,N_20496);
or UO_3372 (O_3372,N_23300,N_22768);
and UO_3373 (O_3373,N_20657,N_28265);
nand UO_3374 (O_3374,N_22267,N_21628);
nor UO_3375 (O_3375,N_27535,N_27706);
xnor UO_3376 (O_3376,N_26269,N_28320);
and UO_3377 (O_3377,N_22891,N_23927);
nand UO_3378 (O_3378,N_26576,N_28999);
or UO_3379 (O_3379,N_21855,N_26230);
nor UO_3380 (O_3380,N_20435,N_22592);
nor UO_3381 (O_3381,N_25468,N_22408);
and UO_3382 (O_3382,N_23180,N_21265);
or UO_3383 (O_3383,N_21631,N_21963);
nand UO_3384 (O_3384,N_29636,N_21377);
xnor UO_3385 (O_3385,N_24479,N_23183);
xnor UO_3386 (O_3386,N_23585,N_27484);
xnor UO_3387 (O_3387,N_21340,N_27499);
nand UO_3388 (O_3388,N_25034,N_24993);
and UO_3389 (O_3389,N_23153,N_24174);
nand UO_3390 (O_3390,N_27806,N_22141);
nor UO_3391 (O_3391,N_21750,N_25999);
nor UO_3392 (O_3392,N_23928,N_28445);
xor UO_3393 (O_3393,N_27057,N_25700);
or UO_3394 (O_3394,N_28324,N_20278);
nand UO_3395 (O_3395,N_24703,N_25363);
nor UO_3396 (O_3396,N_24537,N_26592);
nand UO_3397 (O_3397,N_28805,N_24273);
nor UO_3398 (O_3398,N_20550,N_24340);
or UO_3399 (O_3399,N_27975,N_24988);
nand UO_3400 (O_3400,N_21292,N_22601);
xnor UO_3401 (O_3401,N_29955,N_20926);
and UO_3402 (O_3402,N_24294,N_21478);
nor UO_3403 (O_3403,N_27903,N_21752);
nor UO_3404 (O_3404,N_20509,N_20361);
nor UO_3405 (O_3405,N_26058,N_21007);
xor UO_3406 (O_3406,N_29188,N_22511);
nor UO_3407 (O_3407,N_27091,N_20564);
or UO_3408 (O_3408,N_21311,N_20547);
xor UO_3409 (O_3409,N_24414,N_21513);
nor UO_3410 (O_3410,N_23509,N_20356);
xor UO_3411 (O_3411,N_20275,N_22529);
or UO_3412 (O_3412,N_24170,N_25663);
nor UO_3413 (O_3413,N_29302,N_27443);
or UO_3414 (O_3414,N_27464,N_20327);
nor UO_3415 (O_3415,N_25206,N_21791);
nand UO_3416 (O_3416,N_24617,N_21695);
nor UO_3417 (O_3417,N_29896,N_25315);
nand UO_3418 (O_3418,N_27440,N_23719);
and UO_3419 (O_3419,N_20889,N_23520);
and UO_3420 (O_3420,N_29943,N_24923);
xnor UO_3421 (O_3421,N_20636,N_22040);
xor UO_3422 (O_3422,N_24690,N_28587);
nor UO_3423 (O_3423,N_25419,N_22432);
nor UO_3424 (O_3424,N_25450,N_23233);
and UO_3425 (O_3425,N_28379,N_28836);
nand UO_3426 (O_3426,N_20348,N_28197);
nand UO_3427 (O_3427,N_25728,N_25252);
or UO_3428 (O_3428,N_24456,N_28076);
or UO_3429 (O_3429,N_26983,N_25432);
xnor UO_3430 (O_3430,N_27264,N_23955);
and UO_3431 (O_3431,N_26051,N_22846);
and UO_3432 (O_3432,N_26961,N_21156);
nor UO_3433 (O_3433,N_21047,N_29202);
nor UO_3434 (O_3434,N_29355,N_23967);
and UO_3435 (O_3435,N_27691,N_20497);
nand UO_3436 (O_3436,N_26536,N_20770);
or UO_3437 (O_3437,N_24714,N_24028);
and UO_3438 (O_3438,N_20709,N_25741);
and UO_3439 (O_3439,N_20835,N_27905);
nor UO_3440 (O_3440,N_20947,N_25828);
nor UO_3441 (O_3441,N_22971,N_20718);
and UO_3442 (O_3442,N_29294,N_27338);
xor UO_3443 (O_3443,N_28356,N_20119);
nor UO_3444 (O_3444,N_26745,N_23406);
xor UO_3445 (O_3445,N_27295,N_21307);
xor UO_3446 (O_3446,N_23266,N_26648);
and UO_3447 (O_3447,N_28607,N_23115);
and UO_3448 (O_3448,N_28200,N_24380);
or UO_3449 (O_3449,N_24477,N_23408);
nor UO_3450 (O_3450,N_27350,N_20924);
xnor UO_3451 (O_3451,N_29576,N_24883);
nand UO_3452 (O_3452,N_25147,N_21984);
or UO_3453 (O_3453,N_25919,N_21456);
or UO_3454 (O_3454,N_26329,N_28573);
xnor UO_3455 (O_3455,N_25595,N_27907);
or UO_3456 (O_3456,N_26247,N_22808);
and UO_3457 (O_3457,N_24772,N_29993);
and UO_3458 (O_3458,N_20927,N_21218);
and UO_3459 (O_3459,N_24149,N_22151);
nor UO_3460 (O_3460,N_21121,N_24825);
nor UO_3461 (O_3461,N_23868,N_26065);
or UO_3462 (O_3462,N_26322,N_28655);
and UO_3463 (O_3463,N_20500,N_26779);
xnor UO_3464 (O_3464,N_26022,N_23401);
xnor UO_3465 (O_3465,N_29674,N_27989);
and UO_3466 (O_3466,N_20857,N_25076);
nand UO_3467 (O_3467,N_29773,N_20117);
and UO_3468 (O_3468,N_22869,N_28918);
nor UO_3469 (O_3469,N_29337,N_25827);
and UO_3470 (O_3470,N_22663,N_21602);
nand UO_3471 (O_3471,N_29483,N_20696);
nor UO_3472 (O_3472,N_22597,N_26811);
and UO_3473 (O_3473,N_27754,N_23615);
xnor UO_3474 (O_3474,N_20038,N_28277);
or UO_3475 (O_3475,N_23429,N_23035);
or UO_3476 (O_3476,N_24408,N_23352);
and UO_3477 (O_3477,N_21977,N_25364);
xnor UO_3478 (O_3478,N_20886,N_25671);
and UO_3479 (O_3479,N_20437,N_21135);
xnor UO_3480 (O_3480,N_26946,N_22736);
xnor UO_3481 (O_3481,N_27593,N_27476);
nor UO_3482 (O_3482,N_29545,N_27372);
or UO_3483 (O_3483,N_24631,N_20813);
nor UO_3484 (O_3484,N_21858,N_27883);
nor UO_3485 (O_3485,N_24781,N_22038);
nor UO_3486 (O_3486,N_25511,N_25991);
or UO_3487 (O_3487,N_23646,N_24328);
or UO_3488 (O_3488,N_29513,N_23614);
nand UO_3489 (O_3489,N_21609,N_29094);
xnor UO_3490 (O_3490,N_20026,N_21966);
or UO_3491 (O_3491,N_26423,N_21256);
or UO_3492 (O_3492,N_25863,N_21836);
or UO_3493 (O_3493,N_24410,N_25937);
nand UO_3494 (O_3494,N_24871,N_23391);
xnor UO_3495 (O_3495,N_24536,N_24740);
or UO_3496 (O_3496,N_25934,N_22726);
nand UO_3497 (O_3497,N_22440,N_25658);
nand UO_3498 (O_3498,N_28885,N_28517);
xor UO_3499 (O_3499,N_21343,N_22301);
endmodule