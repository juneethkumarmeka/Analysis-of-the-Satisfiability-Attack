module basic_3000_30000_3500_6_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_2357,In_2051);
or U1 (N_1,In_1438,In_962);
or U2 (N_2,In_2031,In_1035);
xor U3 (N_3,In_632,In_292);
nand U4 (N_4,In_2272,In_2907);
nor U5 (N_5,In_839,In_1126);
or U6 (N_6,In_2347,In_2615);
and U7 (N_7,In_2525,In_2395);
nor U8 (N_8,In_730,In_1159);
and U9 (N_9,In_2631,In_1474);
xor U10 (N_10,In_600,In_1161);
or U11 (N_11,In_174,In_1489);
and U12 (N_12,In_2024,In_1901);
or U13 (N_13,In_43,In_2796);
or U14 (N_14,In_112,In_1208);
nand U15 (N_15,In_2021,In_888);
xnor U16 (N_16,In_2586,In_252);
or U17 (N_17,In_489,In_1639);
and U18 (N_18,In_2405,In_2354);
or U19 (N_19,In_2559,In_1278);
xnor U20 (N_20,In_2949,In_986);
nor U21 (N_21,In_2565,In_1670);
or U22 (N_22,In_2532,In_2128);
nand U23 (N_23,In_2613,In_224);
and U24 (N_24,In_760,In_2281);
or U25 (N_25,In_2713,In_1733);
or U26 (N_26,In_2132,In_2098);
nor U27 (N_27,In_1596,In_1120);
xnor U28 (N_28,In_540,In_2492);
xnor U29 (N_29,In_1478,In_1884);
and U30 (N_30,In_889,In_2429);
nand U31 (N_31,In_1349,In_1079);
nand U32 (N_32,In_2014,In_1512);
xnor U33 (N_33,In_687,In_793);
xnor U34 (N_34,In_1954,In_1076);
nor U35 (N_35,In_2044,In_812);
xnor U36 (N_36,In_729,In_2574);
xor U37 (N_37,In_827,In_755);
or U38 (N_38,In_1694,In_204);
and U39 (N_39,In_2498,In_543);
nand U40 (N_40,In_138,In_2570);
xor U41 (N_41,In_2939,In_1855);
and U42 (N_42,In_906,In_2287);
nand U43 (N_43,In_2725,In_518);
nor U44 (N_44,In_1889,In_1946);
xor U45 (N_45,In_2428,In_1168);
xor U46 (N_46,In_738,In_2798);
or U47 (N_47,In_2439,In_660);
or U48 (N_48,In_1647,In_1460);
nand U49 (N_49,In_2776,In_2487);
nand U50 (N_50,In_2847,In_1949);
xor U51 (N_51,In_1007,In_2566);
or U52 (N_52,In_716,In_2434);
nor U53 (N_53,In_1722,In_2511);
xnor U54 (N_54,In_1535,In_1108);
nor U55 (N_55,In_1741,In_461);
and U56 (N_56,In_573,In_2900);
nor U57 (N_57,In_2137,In_1262);
xnor U58 (N_58,In_1899,In_2087);
and U59 (N_59,In_864,In_711);
and U60 (N_60,In_1685,In_2226);
nor U61 (N_61,In_1854,In_918);
nand U62 (N_62,In_858,In_1246);
nor U63 (N_63,In_39,In_2368);
or U64 (N_64,In_1545,In_1338);
nor U65 (N_65,In_2076,In_1216);
nand U66 (N_66,In_780,In_2469);
nand U67 (N_67,In_1784,In_1215);
and U68 (N_68,In_1140,In_1156);
nand U69 (N_69,In_1307,In_1731);
or U70 (N_70,In_395,In_968);
nor U71 (N_71,In_1498,In_18);
and U72 (N_72,In_8,In_1888);
nor U73 (N_73,In_1905,In_2546);
and U74 (N_74,In_616,In_647);
or U75 (N_75,In_2743,In_2874);
nand U76 (N_76,In_1525,In_2540);
xnor U77 (N_77,In_26,In_25);
and U78 (N_78,In_1196,In_2111);
and U79 (N_79,In_2928,In_1265);
or U80 (N_80,In_1983,In_1031);
and U81 (N_81,In_1255,In_1241);
nor U82 (N_82,In_1470,In_2916);
and U83 (N_83,In_820,In_2812);
or U84 (N_84,In_2034,In_2188);
and U85 (N_85,In_2698,In_879);
xnor U86 (N_86,In_1613,In_2504);
xnor U87 (N_87,In_2501,In_1048);
nand U88 (N_88,In_41,In_2079);
xor U89 (N_89,In_2551,In_46);
or U90 (N_90,In_603,In_1394);
nand U91 (N_91,In_1198,In_577);
nand U92 (N_92,In_2058,In_12);
or U93 (N_93,In_185,In_1938);
and U94 (N_94,In_13,In_923);
and U95 (N_95,In_1017,In_1866);
xnor U96 (N_96,In_2769,In_2976);
xor U97 (N_97,In_2389,In_1443);
and U98 (N_98,In_662,In_1038);
nor U99 (N_99,In_1147,In_2040);
and U100 (N_100,In_939,In_1520);
and U101 (N_101,In_1092,In_506);
nand U102 (N_102,In_98,In_741);
and U103 (N_103,In_291,In_2249);
nand U104 (N_104,In_1734,In_1605);
xor U105 (N_105,In_439,In_2482);
nor U106 (N_106,In_2609,In_2314);
nor U107 (N_107,In_1936,In_2445);
xor U108 (N_108,In_173,In_1100);
or U109 (N_109,In_2390,In_708);
nor U110 (N_110,In_2107,In_2260);
xor U111 (N_111,In_2625,In_1451);
nor U112 (N_112,In_285,In_628);
nand U113 (N_113,In_424,In_2601);
or U114 (N_114,In_757,In_2484);
nand U115 (N_115,In_1423,In_2538);
nand U116 (N_116,In_2215,In_239);
or U117 (N_117,In_2035,In_1067);
or U118 (N_118,In_2396,In_2801);
or U119 (N_119,In_1886,In_1664);
or U120 (N_120,In_1740,In_750);
nand U121 (N_121,In_474,In_2708);
nor U122 (N_122,In_1912,In_2295);
nor U123 (N_123,In_1948,In_672);
nor U124 (N_124,In_902,In_2481);
xnor U125 (N_125,In_1125,In_592);
nor U126 (N_126,In_2223,In_1167);
nor U127 (N_127,In_1226,In_823);
nand U128 (N_128,In_2321,In_2459);
or U129 (N_129,In_1051,In_2290);
nor U130 (N_130,In_323,In_1206);
nand U131 (N_131,In_1422,In_1466);
or U132 (N_132,In_153,In_2756);
xnor U133 (N_133,In_1687,In_2746);
nand U134 (N_134,In_2921,In_2029);
nor U135 (N_135,In_2239,In_1069);
nand U136 (N_136,In_1700,In_289);
or U137 (N_137,In_1229,In_2787);
nand U138 (N_138,In_1153,In_1080);
xnor U139 (N_139,In_2810,In_122);
or U140 (N_140,In_2773,In_2213);
and U141 (N_141,In_2261,In_1698);
nor U142 (N_142,In_1404,In_2224);
or U143 (N_143,In_1078,In_142);
nand U144 (N_144,In_693,In_208);
nand U145 (N_145,In_2041,In_2608);
xor U146 (N_146,In_818,In_1292);
xnor U147 (N_147,In_2760,In_2083);
nor U148 (N_148,In_453,In_372);
nor U149 (N_149,In_2156,In_1251);
nor U150 (N_150,In_278,In_2997);
nand U151 (N_151,In_264,In_2503);
nand U152 (N_152,In_1524,In_1207);
and U153 (N_153,In_960,In_131);
nand U154 (N_154,In_1186,In_193);
and U155 (N_155,In_211,In_219);
nand U156 (N_156,In_1406,In_1461);
nand U157 (N_157,In_2174,In_2596);
xnor U158 (N_158,In_1675,In_1143);
xnor U159 (N_159,In_1641,In_852);
nor U160 (N_160,In_51,In_2234);
and U161 (N_161,In_1157,In_557);
nor U162 (N_162,In_2788,In_2605);
xnor U163 (N_163,In_2641,In_4);
nor U164 (N_164,In_2387,In_1094);
xor U165 (N_165,In_854,In_1961);
nand U166 (N_166,In_1789,In_2919);
xnor U167 (N_167,In_1809,In_949);
nor U168 (N_168,In_56,In_761);
and U169 (N_169,In_250,In_240);
or U170 (N_170,In_2818,In_2175);
xor U171 (N_171,In_1297,In_2946);
nand U172 (N_172,In_1832,In_1608);
nor U173 (N_173,In_1926,In_578);
nor U174 (N_174,In_1367,In_1539);
nand U175 (N_175,In_764,In_574);
and U176 (N_176,In_1804,In_58);
xnor U177 (N_177,In_1458,In_1577);
or U178 (N_178,In_2729,In_2531);
nand U179 (N_179,In_2150,In_629);
and U180 (N_180,In_587,In_2467);
nand U181 (N_181,In_2251,In_2894);
or U182 (N_182,In_245,In_1454);
and U183 (N_183,In_2100,In_649);
nor U184 (N_184,In_200,In_2284);
nand U185 (N_185,In_2977,In_350);
nand U186 (N_186,In_1324,In_1202);
and U187 (N_187,In_1074,In_899);
xor U188 (N_188,In_2248,In_329);
or U189 (N_189,In_1752,In_642);
and U190 (N_190,In_1591,In_352);
nand U191 (N_191,In_973,In_984);
and U192 (N_192,In_859,In_2816);
and U193 (N_193,In_2211,In_1021);
nor U194 (N_194,In_2673,In_105);
xor U195 (N_195,In_1183,In_1558);
or U196 (N_196,In_2136,In_2587);
nand U197 (N_197,In_2312,In_1385);
nor U198 (N_198,In_2005,In_1584);
xor U199 (N_199,In_2981,In_2697);
nor U200 (N_200,In_2583,In_2862);
nor U201 (N_201,In_874,In_732);
or U202 (N_202,In_465,In_281);
nand U203 (N_203,In_405,In_494);
or U204 (N_204,In_1293,In_2356);
nor U205 (N_205,In_2351,In_2856);
nand U206 (N_206,In_1341,In_581);
nand U207 (N_207,In_2264,In_2783);
nand U208 (N_208,In_1298,In_1362);
xnor U209 (N_209,In_1791,In_928);
xnor U210 (N_210,In_1402,In_917);
nor U211 (N_211,In_810,In_2651);
nor U212 (N_212,In_1321,In_1010);
and U213 (N_213,In_1838,In_322);
nor U214 (N_214,In_109,In_1672);
nand U215 (N_215,In_511,In_802);
nand U216 (N_216,In_2344,In_325);
and U217 (N_217,In_2747,In_2336);
and U218 (N_218,In_976,In_1531);
and U219 (N_219,In_608,In_2162);
and U220 (N_220,In_719,In_32);
or U221 (N_221,In_2302,In_2600);
xnor U222 (N_222,In_381,In_2706);
and U223 (N_223,In_2008,In_2696);
nor U224 (N_224,In_157,In_95);
or U225 (N_225,In_2055,In_754);
and U226 (N_226,In_2388,In_2549);
nor U227 (N_227,In_2966,In_2122);
or U228 (N_228,In_2176,In_113);
or U229 (N_229,In_624,In_2508);
xor U230 (N_230,In_510,In_2967);
or U231 (N_231,In_735,In_167);
and U232 (N_232,In_1066,In_1743);
and U233 (N_233,In_1086,In_2075);
nand U234 (N_234,In_2377,In_2449);
xnor U235 (N_235,In_1121,In_1070);
nor U236 (N_236,In_1767,In_903);
nand U237 (N_237,In_2789,In_2210);
or U238 (N_238,In_1413,In_2320);
or U239 (N_239,In_900,In_1450);
and U240 (N_240,In_2443,In_2927);
nand U241 (N_241,In_2384,In_952);
xnor U242 (N_242,In_2984,In_568);
or U243 (N_243,In_2635,In_1697);
xnor U244 (N_244,In_368,In_295);
or U245 (N_245,In_1075,In_2971);
nor U246 (N_246,In_396,In_1118);
and U247 (N_247,In_569,In_29);
xor U248 (N_248,In_2640,In_2474);
nand U249 (N_249,In_2216,In_2456);
xor U250 (N_250,In_2716,In_1371);
or U251 (N_251,In_2313,In_2164);
xor U252 (N_252,In_2143,In_1538);
or U253 (N_253,In_297,In_438);
nand U254 (N_254,In_2319,In_2165);
nor U255 (N_255,In_1097,In_1704);
nor U256 (N_256,In_2127,In_123);
xnor U257 (N_257,In_1530,In_2373);
nor U258 (N_258,In_1440,In_1477);
or U259 (N_259,In_82,In_2010);
or U260 (N_260,In_2832,In_1570);
nor U261 (N_261,In_1653,In_429);
or U262 (N_262,In_658,In_2218);
and U263 (N_263,In_144,In_31);
nand U264 (N_264,In_2096,In_62);
and U265 (N_265,In_1314,In_1669);
xor U266 (N_266,In_894,In_2734);
or U267 (N_267,In_1415,In_821);
nor U268 (N_268,In_2723,In_831);
xor U269 (N_269,In_759,In_1148);
xor U270 (N_270,In_320,In_1057);
or U271 (N_271,In_2733,In_2870);
nor U272 (N_272,In_998,In_1785);
nor U273 (N_273,In_773,In_857);
and U274 (N_274,In_117,In_304);
and U275 (N_275,In_695,In_1792);
nor U276 (N_276,In_644,In_2001);
nor U277 (N_277,In_988,In_2674);
xor U278 (N_278,In_2857,In_572);
nand U279 (N_279,In_1011,In_1453);
or U280 (N_280,In_290,In_1873);
nor U281 (N_281,In_1906,In_1171);
xnor U282 (N_282,In_2996,In_523);
nor U283 (N_283,In_2705,In_2990);
xor U284 (N_284,In_1276,In_740);
nor U285 (N_285,In_2271,In_1553);
nor U286 (N_286,In_1283,In_1318);
and U287 (N_287,In_1841,In_1860);
or U288 (N_288,In_799,In_959);
nor U289 (N_289,In_1930,In_1029);
nor U290 (N_290,In_2629,In_1346);
and U291 (N_291,In_1678,In_2911);
and U292 (N_292,In_739,In_2661);
nor U293 (N_293,In_584,In_337);
and U294 (N_294,In_2408,In_1334);
or U295 (N_295,In_2550,In_1991);
or U296 (N_296,In_922,In_2555);
or U297 (N_297,In_688,In_2500);
and U298 (N_298,In_38,In_1237);
and U299 (N_299,In_1214,In_2027);
xnor U300 (N_300,In_2229,In_2973);
xnor U301 (N_301,In_1045,In_798);
nor U302 (N_302,In_1452,In_1746);
nand U303 (N_303,In_582,In_196);
or U304 (N_304,In_27,In_606);
nor U305 (N_305,In_2898,In_1662);
nor U306 (N_306,In_2123,In_1054);
and U307 (N_307,In_2867,In_1187);
nand U308 (N_308,In_1637,In_1636);
or U309 (N_309,In_2473,In_701);
nand U310 (N_310,In_1210,In_2642);
or U311 (N_311,In_1617,In_1264);
xnor U312 (N_312,In_528,In_2400);
xnor U313 (N_313,In_875,In_2230);
or U314 (N_314,In_2824,In_1027);
nand U315 (N_315,In_2761,In_14);
or U316 (N_316,In_2161,In_346);
or U317 (N_317,In_2440,In_10);
xor U318 (N_318,In_1881,In_490);
nand U319 (N_319,In_2114,In_751);
and U320 (N_320,In_576,In_1851);
nand U321 (N_321,In_1061,In_473);
xor U322 (N_322,In_656,In_2854);
nor U323 (N_323,In_966,In_1620);
nor U324 (N_324,In_421,In_867);
xor U325 (N_325,In_2536,In_950);
and U326 (N_326,In_1435,In_2422);
and U327 (N_327,In_2666,In_947);
and U328 (N_328,In_2004,In_872);
and U329 (N_329,In_1490,In_2653);
nor U330 (N_330,In_2339,In_2823);
or U331 (N_331,In_1732,In_727);
and U332 (N_332,In_2023,In_293);
or U333 (N_333,In_907,In_1124);
or U334 (N_334,In_630,In_2019);
or U335 (N_335,In_2375,In_2070);
xor U336 (N_336,In_463,In_948);
or U337 (N_337,In_2278,In_1115);
nand U338 (N_338,In_107,In_2941);
nor U339 (N_339,In_2078,In_534);
nor U340 (N_340,In_2257,In_1656);
nor U341 (N_341,In_814,In_1962);
nand U342 (N_342,In_868,In_2677);
xor U343 (N_343,In_2518,In_1372);
nand U344 (N_344,In_2703,In_1002);
nor U345 (N_345,In_2480,In_883);
or U346 (N_346,In_330,In_614);
and U347 (N_347,In_1885,In_1514);
xnor U348 (N_348,In_1555,In_2675);
and U349 (N_349,In_700,In_2332);
nor U350 (N_350,In_1446,In_734);
nand U351 (N_351,In_354,In_2770);
and U352 (N_352,In_2764,In_180);
or U353 (N_353,In_2866,In_1222);
nor U354 (N_354,In_1437,In_1374);
or U355 (N_355,In_251,In_406);
nand U356 (N_356,In_2245,In_1651);
nor U357 (N_357,In_2684,In_591);
or U358 (N_358,In_2554,In_2850);
and U359 (N_359,In_133,In_86);
and U360 (N_360,In_884,In_1279);
nor U361 (N_361,In_397,In_2607);
nand U362 (N_362,In_1462,In_2446);
nand U363 (N_363,In_2291,In_2419);
or U364 (N_364,In_1282,In_2833);
xor U365 (N_365,In_2630,In_1497);
or U366 (N_366,In_2193,In_2145);
or U367 (N_367,In_2370,In_2512);
nor U368 (N_368,In_865,In_669);
and U369 (N_369,In_1060,In_2961);
nor U370 (N_370,In_399,In_1642);
or U371 (N_371,In_2792,In_2335);
xor U372 (N_372,In_526,In_1114);
or U373 (N_373,In_2736,In_605);
nor U374 (N_374,In_2528,In_559);
or U375 (N_375,In_1152,In_1883);
xnor U376 (N_376,In_911,In_2802);
xnor U377 (N_377,In_2730,In_829);
nand U378 (N_378,In_985,In_331);
xnor U379 (N_379,In_2042,In_17);
and U380 (N_380,In_76,In_996);
xor U381 (N_381,In_1026,In_1797);
and U382 (N_382,In_1256,In_897);
nor U383 (N_383,In_736,In_1526);
nand U384 (N_384,In_2177,In_747);
or U385 (N_385,In_766,In_183);
or U386 (N_386,In_537,In_1622);
nand U387 (N_387,In_992,In_77);
nand U388 (N_388,In_1676,In_42);
nand U389 (N_389,In_125,In_1914);
xor U390 (N_390,In_989,In_2670);
nor U391 (N_391,In_2721,In_413);
nor U392 (N_392,In_1922,In_1981);
nor U393 (N_393,In_909,In_2380);
xor U394 (N_394,In_1880,In_593);
and U395 (N_395,In_535,In_1723);
nor U396 (N_396,In_2880,In_2829);
xnor U397 (N_397,In_307,In_1794);
nor U398 (N_398,In_1122,In_2516);
nand U399 (N_399,In_2054,In_493);
xnor U400 (N_400,In_2081,In_247);
and U401 (N_401,In_2057,In_314);
xor U402 (N_402,In_207,In_1049);
xor U403 (N_403,In_1380,In_2187);
xnor U404 (N_404,In_509,In_2073);
and U405 (N_405,In_963,In_861);
xor U406 (N_406,In_2648,In_1829);
and U407 (N_407,In_2196,In_550);
nor U408 (N_408,In_936,In_2950);
nand U409 (N_409,In_2731,In_746);
xnor U410 (N_410,In_2378,In_1467);
or U411 (N_411,In_446,In_2841);
nand U412 (N_412,In_1095,In_1379);
nand U413 (N_413,In_2914,In_2852);
nand U414 (N_414,In_981,In_2933);
xor U415 (N_415,In_2877,In_1893);
xor U416 (N_416,In_2863,In_83);
or U417 (N_417,In_1598,In_1518);
nor U418 (N_418,In_1875,In_1252);
nor U419 (N_419,In_1041,In_2737);
xnor U420 (N_420,In_308,In_2381);
and U421 (N_421,In_1505,In_1878);
or U422 (N_422,In_1516,In_1610);
nand U423 (N_423,In_525,In_1691);
xnor U424 (N_424,In_2668,In_1769);
nand U425 (N_425,In_1344,In_1311);
nand U426 (N_426,In_1817,In_2748);
nor U427 (N_427,In_1588,In_503);
and U428 (N_428,In_2153,In_666);
xnor U429 (N_429,In_1308,In_1907);
nand U430 (N_430,In_458,In_707);
xnor U431 (N_431,In_932,In_1287);
nor U432 (N_432,In_2955,In_995);
xnor U433 (N_433,In_1679,In_1790);
nand U434 (N_434,In_2785,In_154);
xor U435 (N_435,In_938,In_206);
or U436 (N_436,In_1129,In_1472);
nand U437 (N_437,In_2246,In_2735);
and U438 (N_438,In_2575,In_787);
or U439 (N_439,In_2752,In_2093);
nand U440 (N_440,In_1179,In_1064);
or U441 (N_441,In_1503,In_1680);
nand U442 (N_442,In_887,In_1688);
and U443 (N_443,In_621,In_143);
nand U444 (N_444,In_280,In_440);
or U445 (N_445,In_2690,In_671);
nand U446 (N_446,In_2269,In_1668);
nor U447 (N_447,In_703,In_2560);
or U448 (N_448,In_2464,In_2235);
nor U449 (N_449,In_1915,In_1169);
xnor U450 (N_450,In_811,In_2252);
nor U451 (N_451,In_1939,In_2688);
or U452 (N_452,In_1270,In_384);
xnor U453 (N_453,In_698,In_558);
nor U454 (N_454,In_796,In_1177);
and U455 (N_455,In_1508,In_2308);
nor U456 (N_456,In_638,In_2781);
nand U457 (N_457,In_676,In_2454);
nand U458 (N_458,In_679,In_404);
and U459 (N_459,In_385,In_1395);
and U460 (N_460,In_1382,In_2931);
nand U461 (N_461,In_2542,In_1576);
nand U462 (N_462,In_1828,In_2279);
nor U463 (N_463,In_2227,In_2367);
xor U464 (N_464,In_1399,In_565);
nor U465 (N_465,In_2940,In_2918);
or U466 (N_466,In_826,In_588);
nand U467 (N_467,In_910,In_2751);
and U468 (N_468,In_1476,In_1378);
and U469 (N_469,In_394,In_2831);
nand U470 (N_470,In_2263,In_541);
nand U471 (N_471,In_324,In_1568);
nor U472 (N_472,In_1299,In_1228);
xor U473 (N_473,In_2695,In_2039);
nand U474 (N_474,In_2365,In_1980);
and U475 (N_475,In_101,In_860);
or U476 (N_476,In_2000,In_1223);
or U477 (N_477,In_191,In_2935);
xnor U478 (N_478,In_2478,In_1944);
xor U479 (N_479,In_2169,In_374);
xnor U480 (N_480,In_1155,In_1376);
nor U481 (N_481,In_742,In_1635);
nand U482 (N_482,In_1655,In_226);
nand U483 (N_483,In_2876,In_1448);
xor U484 (N_484,In_1117,In_1400);
and U485 (N_485,In_2745,In_1985);
nor U486 (N_486,In_1389,In_552);
nand U487 (N_487,In_90,In_1105);
xnor U488 (N_488,In_2978,In_1941);
or U489 (N_489,In_2899,In_1260);
or U490 (N_490,In_1205,In_502);
xor U491 (N_491,In_492,In_2502);
nor U492 (N_492,In_2206,In_74);
or U493 (N_493,In_1877,In_1397);
and U494 (N_494,In_410,In_79);
nor U495 (N_495,In_305,In_1109);
nand U496 (N_496,In_594,In_483);
xnor U497 (N_497,In_2089,In_481);
nor U498 (N_498,In_2208,In_1840);
xnor U499 (N_499,In_1869,In_2598);
or U500 (N_500,In_517,In_646);
and U501 (N_501,In_2168,In_2527);
and U502 (N_502,In_1336,In_1759);
nand U503 (N_503,In_1291,In_89);
nand U504 (N_504,In_2717,In_2844);
and U505 (N_505,In_1003,In_667);
xor U506 (N_506,In_2348,In_2424);
and U507 (N_507,In_271,In_345);
nand U508 (N_508,In_1456,In_1504);
and U509 (N_509,In_1702,In_2633);
and U510 (N_510,In_1193,In_300);
nand U511 (N_511,In_794,In_1625);
and U512 (N_512,In_1527,In_1744);
nor U513 (N_513,In_1442,In_328);
and U514 (N_514,In_319,In_166);
nand U515 (N_515,In_570,In_1275);
or U516 (N_516,In_2962,In_246);
nor U517 (N_517,In_2460,In_256);
or U518 (N_518,In_838,In_2772);
or U519 (N_519,In_2762,In_1500);
xnor U520 (N_520,In_2709,In_2082);
xor U521 (N_521,In_1931,In_2425);
and U522 (N_522,In_44,In_361);
nand U523 (N_523,In_382,In_548);
nand U524 (N_524,In_163,In_1312);
nand U525 (N_525,In_155,In_392);
nor U526 (N_526,In_2683,In_1111);
xor U527 (N_527,In_156,In_1047);
xor U528 (N_528,In_1737,In_2391);
nand U529 (N_529,In_1071,In_2763);
and U530 (N_530,In_332,In_2826);
xnor U531 (N_531,In_919,In_2179);
nor U532 (N_532,In_994,In_2139);
nand U533 (N_533,In_341,In_2964);
nor U534 (N_534,In_1649,In_1974);
or U535 (N_535,In_1173,In_1493);
xor U536 (N_536,In_2623,In_2774);
nor U537 (N_537,In_1266,In_485);
nand U538 (N_538,In_1550,In_387);
xor U539 (N_539,In_2152,In_100);
nand U540 (N_540,In_15,In_249);
or U541 (N_541,In_2534,In_1028);
xor U542 (N_542,In_1195,In_2056);
nand U543 (N_543,In_2821,In_1765);
nand U544 (N_544,In_1567,In_1587);
or U545 (N_545,In_54,In_1507);
and U546 (N_546,In_1033,In_2101);
nor U547 (N_547,In_2341,In_2515);
nand U548 (N_548,In_1218,In_1416);
or U549 (N_549,In_199,In_2888);
and U550 (N_550,In_2659,In_70);
and U551 (N_551,In_377,In_836);
and U552 (N_552,In_2529,In_1693);
and U553 (N_553,In_961,In_1468);
nor U554 (N_554,In_1043,In_2447);
xnor U555 (N_555,In_1736,In_477);
or U556 (N_556,In_1856,In_1544);
xor U557 (N_557,In_198,In_1573);
and U558 (N_558,In_265,In_1181);
nor U559 (N_559,In_2750,In_2619);
nand U560 (N_560,In_1863,In_2217);
nand U561 (N_561,In_1082,In_64);
nor U562 (N_562,In_1348,In_2544);
nand U563 (N_563,In_1805,In_2450);
nand U564 (N_564,In_2883,In_1267);
nand U565 (N_565,In_2092,In_2297);
xnor U566 (N_566,In_2893,In_1248);
nand U567 (N_567,In_1023,In_333);
and U568 (N_568,In_2280,In_882);
and U569 (N_569,In_33,In_2414);
nand U570 (N_570,In_21,In_2277);
xor U571 (N_571,In_342,In_2458);
nand U572 (N_572,In_1300,In_486);
nor U573 (N_573,In_2360,In_2599);
and U574 (N_574,In_2214,In_2496);
xor U575 (N_575,In_1850,In_1657);
and U576 (N_576,In_2170,In_1638);
nand U577 (N_577,In_1919,In_2185);
xor U578 (N_578,In_615,In_2724);
xnor U579 (N_579,In_2691,In_969);
nor U580 (N_580,In_30,In_876);
nor U581 (N_581,In_132,In_2944);
nor U582 (N_582,In_1660,In_93);
nor U583 (N_583,In_2121,In_1830);
nor U584 (N_584,In_619,In_2233);
or U585 (N_585,In_1903,In_335);
and U586 (N_586,In_2738,In_57);
xnor U587 (N_587,In_1197,In_2477);
and U588 (N_588,In_1107,In_449);
nand U589 (N_589,In_445,In_231);
and U590 (N_590,In_2800,In_598);
xor U591 (N_591,In_1773,In_1747);
xor U592 (N_592,In_2806,In_1836);
nand U593 (N_593,In_141,In_1738);
nand U594 (N_594,In_205,In_152);
xor U595 (N_595,In_491,In_343);
nand U596 (N_596,In_505,In_715);
and U597 (N_597,In_1436,In_2436);
nand U598 (N_598,In_1822,In_1532);
and U599 (N_599,In_456,In_1988);
or U600 (N_600,In_1132,In_363);
xnor U601 (N_601,In_1062,In_562);
nand U602 (N_602,In_2435,In_129);
xnor U603 (N_603,In_2475,In_1599);
nor U604 (N_604,In_88,In_2805);
nand U605 (N_605,In_0,In_1630);
xnor U606 (N_606,In_987,In_60);
and U607 (N_607,In_2610,In_2399);
and U608 (N_608,In_114,In_937);
nor U609 (N_609,In_2744,In_2882);
and U610 (N_610,In_2557,In_181);
and U611 (N_611,In_1993,In_1585);
xnor U612 (N_612,In_1970,In_942);
nor U613 (N_613,In_2974,In_1257);
nor U614 (N_614,In_1053,In_407);
xnor U615 (N_615,In_1781,In_1842);
nor U616 (N_616,In_1018,In_2767);
or U617 (N_617,In_546,In_2652);
or U618 (N_618,In_312,In_1357);
xor U619 (N_619,In_2956,In_2397);
and U620 (N_620,In_355,In_1084);
nor U621 (N_621,In_1113,In_1063);
or U622 (N_622,In_1564,In_1479);
or U623 (N_623,In_804,In_2485);
and U624 (N_624,In_1646,In_2304);
xor U625 (N_625,In_2009,In_480);
and U626 (N_626,In_1288,In_412);
nor U627 (N_627,In_2672,In_934);
nand U628 (N_628,In_817,In_1964);
or U629 (N_629,In_563,In_139);
nand U630 (N_630,In_87,In_1245);
or U631 (N_631,In_441,In_1444);
nand U632 (N_632,In_2407,In_287);
or U633 (N_633,In_459,In_1760);
nor U634 (N_634,In_2535,In_1541);
xnor U635 (N_635,In_2398,In_659);
nand U636 (N_636,In_599,In_2349);
nor U637 (N_637,In_1849,In_2331);
nand U638 (N_638,In_1058,In_1480);
or U639 (N_639,In_2318,In_1659);
nor U640 (N_640,In_1174,In_2593);
or U641 (N_641,In_1331,In_978);
nor U642 (N_642,In_1284,In_2330);
xor U643 (N_643,In_2561,In_234);
and U644 (N_644,In_1990,In_2497);
xor U645 (N_645,In_696,In_134);
and U646 (N_646,In_1894,In_807);
or U647 (N_647,In_37,In_704);
xnor U648 (N_648,In_2975,In_1238);
xnor U649 (N_649,In_921,In_2418);
nor U650 (N_650,In_2881,In_2120);
nand U651 (N_651,In_2432,In_2637);
or U652 (N_652,In_2147,In_990);
nand U653 (N_653,In_428,In_2180);
nand U654 (N_654,In_426,In_2757);
nor U655 (N_655,In_499,In_391);
and U656 (N_656,In_2392,In_1145);
xnor U657 (N_657,In_2189,In_2563);
or U658 (N_658,In_2074,In_2340);
or U659 (N_659,In_2285,In_1286);
and U660 (N_660,In_2155,In_2342);
nand U661 (N_661,In_49,In_1019);
nor U662 (N_662,In_2393,In_1714);
or U663 (N_663,In_2926,In_210);
nor U664 (N_664,In_2207,In_2571);
xnor U665 (N_665,In_1650,In_2947);
and U666 (N_666,In_957,In_2552);
nand U667 (N_667,In_1088,In_2472);
nor U668 (N_668,In_913,In_1951);
xor U669 (N_669,In_625,In_2203);
nor U670 (N_670,In_159,In_179);
and U671 (N_671,In_681,In_1821);
and U672 (N_672,In_1303,In_1629);
xor U673 (N_673,In_2184,In_195);
xor U674 (N_674,In_965,In_1373);
xor U675 (N_675,In_835,In_35);
xnor U676 (N_676,In_2275,In_1592);
and U677 (N_677,In_2090,In_498);
nor U678 (N_678,In_1098,In_776);
nor U679 (N_679,In_1824,In_873);
nand U680 (N_680,In_652,In_2255);
and U681 (N_681,In_1151,In_2545);
nand U682 (N_682,In_1509,In_1754);
xor U683 (N_683,In_613,In_2992);
xnor U684 (N_684,In_1200,In_1431);
or U685 (N_685,In_1352,In_2817);
xnor U686 (N_686,In_1495,In_1582);
nand U687 (N_687,In_99,In_1005);
nand U688 (N_688,In_409,In_1523);
and U689 (N_689,In_521,In_2116);
xor U690 (N_690,In_2627,In_2020);
xor U691 (N_691,In_1831,In_1227);
or U692 (N_692,In_1745,In_2665);
nor U693 (N_693,In_1219,In_1295);
nand U694 (N_694,In_1093,In_1426);
or U695 (N_695,In_1496,In_1160);
and U696 (N_696,In_169,In_635);
and U697 (N_697,In_411,In_94);
xnor U698 (N_698,In_1194,In_452);
xor U699 (N_699,In_983,In_2682);
and U700 (N_700,In_816,In_2013);
and U701 (N_701,In_1556,In_2309);
nor U702 (N_702,In_168,In_856);
nor U703 (N_703,In_1614,In_1242);
nand U704 (N_704,In_2864,In_612);
nand U705 (N_705,In_431,In_1729);
xor U706 (N_706,In_2982,In_650);
and U707 (N_707,In_2886,In_1189);
and U708 (N_708,In_1777,In_2199);
or U709 (N_709,In_1277,In_2848);
or U710 (N_710,In_1910,In_2576);
nand U711 (N_711,In_1424,In_401);
xnor U712 (N_712,In_484,In_348);
nor U713 (N_713,In_1803,In_609);
nand U714 (N_714,In_2517,In_2507);
nor U715 (N_715,In_1801,In_1956);
or U716 (N_716,In_116,In_1482);
xnor U717 (N_717,In_2692,In_2465);
and U718 (N_718,In_1337,In_2306);
nor U719 (N_719,In_837,In_1923);
or U720 (N_720,In_2647,In_1325);
or U721 (N_721,In_437,In_28);
and U722 (N_722,In_1134,In_497);
nand U723 (N_723,In_2803,In_1945);
nand U724 (N_724,In_149,In_1192);
xor U725 (N_725,In_2603,In_217);
or U726 (N_726,In_1104,In_1771);
nand U727 (N_727,In_182,In_1645);
xor U728 (N_728,In_1806,In_1681);
nor U729 (N_729,In_529,In_487);
and U730 (N_730,In_877,In_2644);
nand U731 (N_731,In_2969,In_259);
and U732 (N_732,In_20,In_1742);
xnor U733 (N_733,In_1965,In_1459);
and U734 (N_734,In_2346,In_1847);
and U735 (N_735,In_1870,In_782);
xor U736 (N_736,In_2929,In_334);
or U737 (N_737,In_640,In_2327);
xnor U738 (N_738,In_1099,In_1327);
xor U739 (N_739,In_1992,In_895);
or U740 (N_740,In_2292,In_1231);
and U741 (N_741,In_1862,In_870);
xnor U742 (N_742,In_1667,In_1220);
or U743 (N_743,In_1865,In_991);
nor U744 (N_744,In_2906,In_2448);
nor U745 (N_745,In_1640,In_1652);
nor U746 (N_746,In_1952,In_2758);
or U747 (N_747,In_849,In_327);
xnor U748 (N_748,In_2835,In_862);
nor U749 (N_749,In_1934,In_2028);
nor U750 (N_750,In_1543,In_1859);
and U751 (N_751,In_119,In_846);
and U752 (N_752,In_944,In_2957);
and U753 (N_753,In_227,In_2842);
and U754 (N_754,In_1786,In_637);
nand U755 (N_755,In_2254,In_964);
nor U756 (N_756,In_2316,In_2755);
nor U757 (N_757,In_2628,In_2329);
xnor U758 (N_758,In_2305,In_2875);
nor U759 (N_759,In_1643,In_723);
nor U760 (N_760,In_2222,In_1712);
nor U761 (N_761,In_2951,In_2151);
nand U762 (N_762,In_2068,In_752);
and U763 (N_763,In_286,In_1250);
nor U764 (N_764,In_690,In_1274);
nor U765 (N_765,In_1320,In_2958);
xnor U766 (N_766,In_233,In_2288);
and U767 (N_767,In_257,In_2680);
or U768 (N_768,In_538,In_2896);
nand U769 (N_769,In_1916,In_2726);
or U770 (N_770,In_9,In_97);
nand U771 (N_771,In_532,In_1633);
nand U772 (N_772,In_1818,In_1563);
nand U773 (N_773,In_1929,In_110);
or U774 (N_774,In_1464,In_1201);
nand U775 (N_775,In_1616,In_73);
nor U776 (N_776,In_1823,In_2061);
xor U777 (N_777,In_1020,In_2112);
nand U778 (N_778,In_1932,In_1506);
nand U779 (N_779,In_1433,In_2220);
and U780 (N_780,In_1056,In_55);
nor U781 (N_781,In_2578,In_1799);
nand U782 (N_782,In_197,In_769);
or U783 (N_783,In_72,In_420);
and U784 (N_784,In_338,In_1024);
nor U785 (N_785,In_260,In_2259);
or U786 (N_786,In_1795,In_722);
nor U787 (N_787,In_2741,In_1239);
xor U788 (N_788,In_2676,In_161);
or U789 (N_789,In_2416,In_1612);
nand U790 (N_790,In_2361,In_560);
or U791 (N_791,In_2015,In_2790);
nor U792 (N_792,In_2582,In_845);
nor U793 (N_793,In_686,In_1235);
nand U794 (N_794,In_2366,In_519);
nor U795 (N_795,In_2699,In_261);
nand U796 (N_796,In_1977,In_1233);
nor U797 (N_797,In_726,In_1142);
or U798 (N_798,In_824,In_1994);
nor U799 (N_799,In_571,In_2577);
nand U800 (N_800,In_2138,In_1203);
xor U801 (N_801,In_745,In_1959);
nand U802 (N_802,In_1853,In_2558);
nand U803 (N_803,In_1175,In_2667);
nor U804 (N_804,In_2413,In_318);
or U805 (N_805,In_1383,In_1749);
xor U806 (N_806,In_1561,In_2242);
nand U807 (N_807,In_2433,In_1360);
or U808 (N_808,In_2225,In_1796);
xnor U809 (N_809,In_215,In_767);
and U810 (N_810,In_148,In_1684);
nand U811 (N_811,In_784,In_1340);
nor U812 (N_812,In_710,In_1928);
nor U813 (N_813,In_1013,In_2658);
xor U814 (N_814,In_2038,In_2195);
and U815 (N_815,In_2533,In_1557);
nand U816 (N_816,In_880,In_2200);
nand U817 (N_817,In_2626,In_941);
nand U818 (N_818,In_1874,In_2374);
nand U819 (N_819,In_16,In_2543);
nand U820 (N_820,In_176,In_2860);
nor U821 (N_821,In_1149,In_758);
xor U822 (N_822,In_296,In_209);
nor U823 (N_823,In_1368,In_2258);
and U824 (N_824,In_45,In_201);
or U825 (N_825,In_2172,In_2853);
and U826 (N_826,In_1254,In_2228);
and U827 (N_827,In_1943,In_2402);
or U828 (N_828,In_365,In_1690);
or U829 (N_829,In_2960,In_788);
nand U830 (N_830,In_2564,In_262);
and U831 (N_831,In_2845,In_1654);
xnor U832 (N_832,In_136,In_2085);
nor U833 (N_833,In_651,In_1486);
nor U834 (N_834,In_400,In_2791);
nand U835 (N_835,In_7,In_871);
nor U836 (N_836,In_2980,In_1359);
nand U837 (N_837,In_364,In_1313);
xor U838 (N_838,In_1717,In_2572);
or U839 (N_839,In_311,In_2506);
xnor U840 (N_840,In_1172,In_241);
nor U841 (N_841,In_1316,In_1182);
xor U842 (N_842,In_2106,In_2700);
nand U843 (N_843,In_1819,In_1188);
and U844 (N_844,In_2430,In_2495);
or U845 (N_845,In_2837,In_2358);
xor U846 (N_846,In_1756,In_2379);
nand U847 (N_847,In_2025,In_1405);
nand U848 (N_848,In_2237,In_2865);
nand U849 (N_849,In_1301,In_2509);
nor U850 (N_850,In_863,In_1987);
nand U851 (N_851,In_1534,In_466);
and U852 (N_852,In_1996,In_1162);
and U853 (N_853,In_1902,In_2103);
xor U854 (N_854,In_1782,In_2897);
and U855 (N_855,In_1665,In_633);
or U856 (N_856,In_699,In_1713);
and U857 (N_857,In_2711,In_1780);
and U858 (N_858,In_1920,In_1355);
nand U859 (N_859,In_639,In_482);
xor U860 (N_860,In_718,In_2912);
nand U861 (N_861,In_2753,In_302);
nor U862 (N_862,In_436,In_2310);
nand U863 (N_863,In_1391,In_1116);
and U864 (N_864,In_908,In_2129);
and U865 (N_865,In_1848,In_1716);
nand U866 (N_866,In_1548,In_2007);
or U867 (N_867,In_488,In_2846);
or U868 (N_868,In_2827,In_1364);
and U869 (N_869,In_2426,In_1857);
nand U870 (N_870,In_2890,In_1663);
and U871 (N_871,In_2303,In_507);
or U872 (N_872,In_1978,In_539);
xor U873 (N_873,In_2913,In_1006);
and U874 (N_874,In_433,In_269);
or U875 (N_875,In_2328,In_120);
or U876 (N_876,In_1421,In_1273);
xnor U877 (N_877,In_2144,In_1631);
nand U878 (N_878,In_1083,In_531);
and U879 (N_879,In_980,In_1718);
and U880 (N_880,In_1103,In_610);
and U881 (N_881,In_1473,In_2728);
xor U882 (N_882,In_725,In_772);
xnor U883 (N_883,In_2942,In_2855);
xor U884 (N_884,In_2836,In_2471);
and U885 (N_885,In_1549,In_2694);
nor U886 (N_886,In_1887,In_1261);
or U887 (N_887,In_1554,In_367);
and U888 (N_888,In_2868,In_2003);
xor U889 (N_889,In_781,In_69);
xnor U890 (N_890,In_187,In_1290);
and U891 (N_891,In_1249,In_1138);
xnor U892 (N_892,In_2825,In_2970);
nor U893 (N_893,In_2719,In_1022);
or U894 (N_894,In_108,In_705);
or U895 (N_895,In_2830,In_253);
nand U896 (N_896,In_1758,In_830);
nand U897 (N_897,In_2133,In_2183);
or U898 (N_898,In_2352,In_1695);
or U899 (N_899,In_2712,In_50);
nor U900 (N_900,In_2638,In_1342);
xnor U901 (N_901,In_135,In_1579);
nand U902 (N_902,In_213,In_645);
nor U903 (N_903,In_1706,In_1601);
xor U904 (N_904,In_1211,In_379);
nor U905 (N_905,In_709,In_2945);
nor U906 (N_906,In_770,In_1513);
nor U907 (N_907,In_2097,In_2602);
or U908 (N_908,In_1882,In_2326);
xnor U909 (N_909,In_2232,In_366);
nand U910 (N_910,In_2067,In_283);
nor U911 (N_911,In_2643,In_496);
and U912 (N_912,In_544,In_1547);
or U913 (N_913,In_2624,In_1603);
nand U914 (N_914,In_2547,In_2322);
nand U915 (N_915,In_927,In_1529);
and U916 (N_916,In_2113,In_1710);
xor U917 (N_917,In_347,In_2819);
nand U918 (N_918,In_1772,In_2851);
nor U919 (N_919,In_294,In_904);
nor U920 (N_920,In_165,In_1393);
or U921 (N_921,In_2212,In_2404);
or U922 (N_922,In_228,In_1940);
xnor U923 (N_923,In_1133,In_2994);
and U924 (N_924,In_306,In_126);
nor U925 (N_925,In_2995,In_2983);
and U926 (N_926,In_1937,In_1345);
nor U927 (N_927,In_1751,In_221);
nor U928 (N_928,In_2294,In_756);
nor U929 (N_929,In_1546,In_2793);
nor U930 (N_930,In_242,In_22);
nor U931 (N_931,In_1091,In_2462);
nor U932 (N_932,In_2181,In_2839);
xnor U933 (N_933,In_737,In_1158);
or U934 (N_934,In_2298,In_775);
nor U935 (N_935,In_2191,In_585);
or U936 (N_936,In_801,In_2240);
xor U937 (N_937,In_1960,In_692);
and U938 (N_938,In_1230,In_223);
nand U939 (N_939,In_2030,In_1455);
nor U940 (N_940,In_657,In_1326);
nand U941 (N_941,In_151,In_1037);
and U942 (N_942,In_2119,In_848);
xnor U943 (N_943,In_866,In_930);
nor U944 (N_944,In_2569,In_806);
and U945 (N_945,In_1030,In_2584);
nor U946 (N_946,In_714,In_1825);
nand U947 (N_947,In_1609,In_1199);
and U948 (N_948,In_415,In_243);
nor U949 (N_949,In_713,In_665);
and U950 (N_950,In_24,In_85);
nor U951 (N_951,In_235,In_2799);
or U952 (N_952,In_2173,In_2063);
and U953 (N_953,In_2963,In_514);
nor U954 (N_954,In_2808,In_2892);
xor U955 (N_955,In_326,In_890);
xnor U956 (N_956,In_1793,In_586);
or U957 (N_957,In_768,In_2125);
and U958 (N_958,In_1750,In_892);
nand U959 (N_959,In_1365,In_104);
and U960 (N_960,In_1709,In_258);
or U961 (N_961,In_2094,In_2959);
or U962 (N_962,In_2539,In_842);
xor U963 (N_963,In_2505,In_2952);
nand U964 (N_964,In_2779,In_1154);
nor U965 (N_965,In_1000,In_2409);
nand U966 (N_966,In_840,In_1329);
xor U967 (N_967,In_267,In_1044);
and U968 (N_968,In_1096,In_408);
or U969 (N_969,In_1967,In_931);
and U970 (N_970,In_2807,In_524);
or U971 (N_971,In_1762,In_2099);
and U972 (N_972,In_1166,In_146);
nor U973 (N_973,In_1521,In_1615);
or U974 (N_974,In_2022,In_2345);
xor U975 (N_975,In_706,In_2989);
or U976 (N_976,In_2902,In_1190);
or U977 (N_977,In_2221,In_797);
xnor U978 (N_978,In_1788,In_1414);
nand U979 (N_979,In_362,In_943);
and U980 (N_980,In_2333,In_1271);
or U981 (N_981,In_648,In_2059);
nand U982 (N_982,In_2871,In_238);
and U983 (N_983,In_789,In_2141);
nor U984 (N_984,In_214,In_1814);
and U985 (N_985,In_1644,In_59);
nand U986 (N_986,In_1487,In_2820);
xor U987 (N_987,In_5,In_2343);
or U988 (N_988,In_2567,In_1586);
nor U989 (N_989,In_1141,In_673);
nand U990 (N_990,In_2149,In_795);
or U991 (N_991,In_2993,In_771);
and U992 (N_992,In_1330,In_2493);
and U993 (N_993,In_1955,In_1289);
nor U994 (N_994,In_351,In_2080);
or U995 (N_995,In_1933,In_712);
and U996 (N_996,In_2307,In_2489);
nor U997 (N_997,In_2461,In_809);
and U998 (N_998,In_1347,In_2718);
xnor U999 (N_999,In_982,In_34);
nor U1000 (N_1000,In_1969,In_230);
xor U1001 (N_1001,In_2205,In_2104);
xnor U1002 (N_1002,In_1607,In_822);
nor U1003 (N_1003,In_373,In_516);
nand U1004 (N_1004,In_1217,In_791);
xnor U1005 (N_1005,In_457,In_1724);
xor U1006 (N_1006,In_2915,In_1807);
and U1007 (N_1007,In_375,In_1895);
nor U1008 (N_1008,In_1176,In_2274);
or U1009 (N_1009,In_850,In_2991);
or U1010 (N_1010,In_1658,In_721);
and U1011 (N_1011,In_844,In_2036);
xnor U1012 (N_1012,In_177,In_684);
nand U1013 (N_1013,In_1975,In_1628);
nor U1014 (N_1014,In_786,In_779);
nor U1015 (N_1015,In_2268,In_1090);
or U1016 (N_1016,In_1908,In_1410);
nand U1017 (N_1017,In_1533,In_2786);
nand U1018 (N_1018,In_356,In_1185);
nand U1019 (N_1019,In_891,In_2130);
or U1020 (N_1020,In_744,In_1073);
nand U1021 (N_1021,In_2253,In_2286);
and U1022 (N_1022,In_2262,In_2362);
nor U1023 (N_1023,In_896,In_2182);
or U1024 (N_1024,In_2714,In_1971);
nor U1025 (N_1025,In_2766,In_1123);
nand U1026 (N_1026,In_841,In_878);
or U1027 (N_1027,In_1562,In_1280);
nand U1028 (N_1028,In_2537,In_1463);
or U1029 (N_1029,In_2427,In_1178);
xor U1030 (N_1030,In_2580,In_912);
nand U1031 (N_1031,In_434,In_1081);
xnor U1032 (N_1032,In_1701,In_2814);
or U1033 (N_1033,In_1542,In_1835);
nor U1034 (N_1034,In_1682,In_1606);
and U1035 (N_1035,In_743,In_1351);
or U1036 (N_1036,In_3,In_303);
and U1037 (N_1037,In_1999,In_1689);
xor U1038 (N_1038,In_2687,In_1032);
or U1039 (N_1039,In_1966,In_313);
xor U1040 (N_1040,In_2702,In_2524);
nor U1041 (N_1041,In_2923,In_158);
xor U1042 (N_1042,In_935,In_1039);
nor U1043 (N_1043,In_1522,In_1578);
xnor U1044 (N_1044,In_1441,In_23);
and U1045 (N_1045,In_1973,In_1619);
nand U1046 (N_1046,In_1401,In_2660);
or U1047 (N_1047,In_2715,In_170);
or U1048 (N_1048,In_288,In_2026);
xnor U1049 (N_1049,In_1559,In_1725);
xnor U1050 (N_1050,In_1247,In_530);
nor U1051 (N_1051,In_2573,In_2858);
nand U1052 (N_1052,In_2062,In_1131);
xor U1053 (N_1053,In_2466,In_469);
xnor U1054 (N_1054,In_277,In_2813);
nor U1055 (N_1055,In_386,In_254);
and U1056 (N_1056,In_977,In_2047);
nor U1057 (N_1057,In_1517,In_2903);
xor U1058 (N_1058,In_617,In_2732);
and U1059 (N_1059,In_2884,In_435);
nor U1060 (N_1060,In_2148,In_1016);
nor U1061 (N_1061,In_1594,In_2618);
xor U1062 (N_1062,In_2463,In_1761);
nand U1063 (N_1063,In_2108,In_1502);
nand U1064 (N_1064,In_1913,In_1811);
nand U1065 (N_1065,In_1001,In_1306);
or U1066 (N_1066,In_2315,In_80);
nand U1067 (N_1067,In_1484,In_279);
nand U1068 (N_1068,In_924,In_47);
nor U1069 (N_1069,In_597,In_2372);
nand U1070 (N_1070,In_1381,In_1429);
nor U1071 (N_1071,In_430,In_728);
nand U1072 (N_1072,In_1827,In_1510);
or U1073 (N_1073,In_162,In_1634);
xnor U1074 (N_1074,In_229,In_2514);
nand U1075 (N_1075,In_636,In_2091);
and U1076 (N_1076,In_2936,In_1110);
or U1077 (N_1077,In_137,In_1666);
nor U1078 (N_1078,In_2476,In_1816);
and U1079 (N_1079,In_847,In_1236);
nand U1080 (N_1080,In_495,In_1388);
nor U1081 (N_1081,In_2046,In_1304);
nor U1082 (N_1082,In_1677,In_1012);
nand U1083 (N_1083,In_2878,In_2157);
or U1084 (N_1084,In_2300,In_527);
nor U1085 (N_1085,In_2523,In_1315);
nand U1086 (N_1086,In_2159,In_1891);
nor U1087 (N_1087,In_6,In_1204);
nand U1088 (N_1088,In_2590,In_749);
xor U1089 (N_1089,In_2371,In_2194);
and U1090 (N_1090,In_512,In_2722);
nor U1091 (N_1091,In_675,In_1112);
xor U1092 (N_1092,In_2166,In_1748);
and U1093 (N_1093,In_2979,In_2012);
nor U1094 (N_1094,In_1540,In_1135);
and U1095 (N_1095,In_1864,In_2050);
nand U1096 (N_1096,In_2158,In_299);
xnor U1097 (N_1097,In_2654,In_1305);
nand U1098 (N_1098,In_186,In_2186);
nor U1099 (N_1099,In_478,In_2556);
and U1100 (N_1100,In_2873,In_1826);
and U1101 (N_1101,In_471,In_956);
or U1102 (N_1102,In_2192,In_683);
nand U1103 (N_1103,In_972,In_1673);
xnor U1104 (N_1104,In_733,In_282);
nand U1105 (N_1105,In_1009,In_273);
and U1106 (N_1106,In_2649,In_65);
or U1107 (N_1107,In_520,In_556);
xor U1108 (N_1108,In_1963,In_2689);
nand U1109 (N_1109,In_2910,In_1119);
nand U1110 (N_1110,In_1707,In_1232);
nor U1111 (N_1111,In_115,In_2124);
nand U1112 (N_1112,In_1552,In_1571);
xor U1113 (N_1113,In_1595,In_694);
nand U1114 (N_1114,In_317,In_225);
xor U1115 (N_1115,In_1918,In_2244);
xor U1116 (N_1116,In_1212,In_2219);
or U1117 (N_1117,In_792,In_2922);
nor U1118 (N_1118,In_1686,In_915);
nand U1119 (N_1119,In_504,In_2470);
nor U1120 (N_1120,In_220,In_2140);
and U1121 (N_1121,In_389,In_111);
and U1122 (N_1122,In_1720,In_2681);
nand U1123 (N_1123,In_1224,In_2606);
nor U1124 (N_1124,In_2250,In_1386);
nand U1125 (N_1125,In_2704,In_1501);
nand U1126 (N_1126,In_2154,In_522);
or U1127 (N_1127,In_1674,In_2403);
xor U1128 (N_1128,In_1358,In_237);
nor U1129 (N_1129,In_1209,In_2646);
or U1130 (N_1130,In_178,In_1976);
or U1131 (N_1131,In_2581,In_1407);
and U1132 (N_1132,In_2838,In_1408);
nand U1133 (N_1133,In_2198,In_448);
nor U1134 (N_1134,In_777,In_1623);
xor U1135 (N_1135,In_2197,In_975);
and U1136 (N_1136,In_103,In_376);
or U1137 (N_1137,In_765,In_1412);
nor U1138 (N_1138,In_160,In_2334);
nor U1139 (N_1139,In_175,In_1491);
nand U1140 (N_1140,In_1942,In_1621);
nand U1141 (N_1141,In_2775,In_790);
nor U1142 (N_1142,In_2095,In_2011);
nor U1143 (N_1143,In_803,In_2656);
or U1144 (N_1144,In_805,In_808);
xor U1145 (N_1145,In_881,In_2323);
xnor U1146 (N_1146,In_1957,In_2889);
nor U1147 (N_1147,In_1240,In_378);
nand U1148 (N_1148,In_933,In_470);
nor U1149 (N_1149,In_1353,In_349);
and U1150 (N_1150,In_1927,In_425);
xnor U1151 (N_1151,In_1244,In_1566);
xor U1152 (N_1152,In_1699,In_2568);
xnor U1153 (N_1153,In_1755,In_1481);
xnor U1154 (N_1154,In_1872,In_2479);
nand U1155 (N_1155,In_2895,In_2548);
or U1156 (N_1156,In_1323,In_2664);
and U1157 (N_1157,In_2406,In_1485);
nand U1158 (N_1158,In_2887,In_358);
or U1159 (N_1159,In_369,In_1137);
xnor U1160 (N_1160,In_1837,In_2861);
and U1161 (N_1161,In_2686,In_583);
and U1162 (N_1162,In_2053,In_1876);
and U1163 (N_1163,In_1369,In_753);
nor U1164 (N_1164,In_680,In_1350);
nor U1165 (N_1165,In_2859,In_1572);
and U1166 (N_1166,In_2749,In_1072);
nor U1167 (N_1167,In_2066,In_1511);
or U1168 (N_1168,In_1735,In_1040);
and U1169 (N_1169,In_1377,In_244);
and U1170 (N_1170,In_940,In_1551);
nor U1171 (N_1171,In_946,In_1581);
or U1172 (N_1172,In_1144,In_2794);
or U1173 (N_1173,In_1234,In_472);
or U1174 (N_1174,In_1339,In_2759);
or U1175 (N_1175,In_689,In_885);
xor U1176 (N_1176,In_1310,In_66);
and U1177 (N_1177,In_2382,In_1268);
and U1178 (N_1178,In_2904,In_2146);
xnor U1179 (N_1179,In_2238,In_1356);
xor U1180 (N_1180,In_2740,In_2266);
and U1181 (N_1181,In_1366,In_2163);
xnor U1182 (N_1182,In_542,In_1569);
and U1183 (N_1183,In_2,In_1492);
and U1184 (N_1184,In_2679,In_464);
nor U1185 (N_1185,In_414,In_2109);
nand U1186 (N_1186,In_604,In_1420);
and U1187 (N_1187,In_353,In_2885);
xor U1188 (N_1188,In_2201,In_344);
or U1189 (N_1189,In_825,In_2650);
xor U1190 (N_1190,In_999,In_1624);
xnor U1191 (N_1191,In_974,In_1800);
nor U1192 (N_1192,In_979,In_359);
or U1193 (N_1193,In_1600,In_1890);
nand U1194 (N_1194,In_416,In_869);
nor U1195 (N_1195,In_1106,In_2386);
xor U1196 (N_1196,In_1285,In_2135);
and U1197 (N_1197,In_422,In_2604);
nand U1198 (N_1198,In_1213,In_834);
nor U1199 (N_1199,In_2273,In_2363);
nor U1200 (N_1200,In_2270,In_274);
nand U1201 (N_1201,In_641,In_2937);
nand U1202 (N_1202,In_618,In_1127);
nand U1203 (N_1203,In_1618,In_2693);
and U1204 (N_1204,In_1427,In_685);
or U1205 (N_1205,In_171,In_390);
and U1206 (N_1206,In_2457,In_2431);
or U1207 (N_1207,In_1165,In_1515);
and U1208 (N_1208,In_1180,In_1294);
nand U1209 (N_1209,In_1852,In_145);
and U1210 (N_1210,In_663,In_1778);
and U1211 (N_1211,In_2754,In_2353);
nand U1212 (N_1212,In_575,In_1243);
nor U1213 (N_1213,In_1726,In_2612);
nand U1214 (N_1214,In_1014,In_554);
and U1215 (N_1215,In_1008,In_1574);
xnor U1216 (N_1216,In_1627,In_1272);
or U1217 (N_1217,In_2037,In_1363);
and U1218 (N_1218,In_1387,In_1392);
and U1219 (N_1219,In_2663,In_1626);
and U1220 (N_1220,In_953,In_2972);
nand U1221 (N_1221,In_2276,In_2588);
or U1222 (N_1222,In_1602,In_901);
nand U1223 (N_1223,In_2869,In_1087);
nor U1224 (N_1224,In_1499,In_916);
or U1225 (N_1225,In_2369,In_75);
and U1226 (N_1226,In_2739,In_2795);
nor U1227 (N_1227,In_1537,In_1375);
or U1228 (N_1228,In_677,In_2488);
xnor U1229 (N_1229,In_564,In_2925);
nand U1230 (N_1230,In_40,In_1953);
or U1231 (N_1231,In_1768,In_2204);
or U1232 (N_1232,In_602,In_545);
nand U1233 (N_1233,In_2267,In_2727);
xnor U1234 (N_1234,In_398,In_1921);
or U1235 (N_1235,In_748,In_1833);
nand U1236 (N_1236,In_549,In_301);
xnor U1237 (N_1237,In_1332,In_2359);
nand U1238 (N_1238,In_360,In_2771);
or U1239 (N_1239,In_2241,In_2678);
nor U1240 (N_1240,In_1900,In_553);
or U1241 (N_1241,In_1984,In_2809);
or U1242 (N_1242,In_102,In_2171);
xnor U1243 (N_1243,In_172,In_68);
and U1244 (N_1244,In_595,In_655);
and U1245 (N_1245,In_2986,In_2917);
nand U1246 (N_1246,In_1361,In_1580);
and U1247 (N_1247,In_815,In_785);
xor U1248 (N_1248,In_140,In_1845);
or U1249 (N_1249,In_951,In_2620);
nor U1250 (N_1250,In_513,In_1077);
or U1251 (N_1251,In_1705,In_2417);
nor U1252 (N_1252,In_1770,In_1575);
nor U1253 (N_1253,In_2519,In_828);
and U1254 (N_1254,In_1004,In_1604);
nand U1255 (N_1255,In_533,In_547);
xor U1256 (N_1256,In_52,In_2236);
xor U1257 (N_1257,In_2293,In_551);
xor U1258 (N_1258,In_515,In_566);
xnor U1259 (N_1259,In_1457,In_1998);
nand U1260 (N_1260,In_248,In_2084);
nand U1261 (N_1261,In_2901,In_2811);
or U1262 (N_1262,In_536,In_2355);
or U1263 (N_1263,In_1411,In_383);
xnor U1264 (N_1264,In_2987,In_1834);
nand U1265 (N_1265,In_2768,In_1025);
or U1266 (N_1266,In_623,In_236);
nand U1267 (N_1267,In_467,In_1281);
nor U1268 (N_1268,In_298,In_427);
nand U1269 (N_1269,In_1434,In_1296);
and U1270 (N_1270,In_2639,In_2879);
nand U1271 (N_1271,In_631,In_455);
xor U1272 (N_1272,In_2595,In_222);
nand U1273 (N_1273,In_580,In_1101);
or U1274 (N_1274,In_2622,In_203);
nor U1275 (N_1275,In_2891,In_1892);
or U1276 (N_1276,In_763,In_118);
xor U1277 (N_1277,In_1812,In_1065);
and U1278 (N_1278,In_2110,In_607);
or U1279 (N_1279,In_2510,In_2685);
nor U1280 (N_1280,In_1986,In_1432);
xnor U1281 (N_1281,In_276,In_476);
nand U1282 (N_1282,In_2126,In_1958);
and U1283 (N_1283,In_202,In_1259);
xor U1284 (N_1284,In_2909,In_2102);
or U1285 (N_1285,In_2645,In_2077);
or U1286 (N_1286,In_1776,In_2780);
nand U1287 (N_1287,In_2513,In_1950);
xor U1288 (N_1288,In_1597,In_1050);
nand U1289 (N_1289,In_1925,In_2828);
nand U1290 (N_1290,In_1774,In_1924);
nand U1291 (N_1291,In_2072,In_920);
and U1292 (N_1292,In_2442,In_340);
and U1293 (N_1293,In_970,In_2585);
nor U1294 (N_1294,In_508,In_2985);
and U1295 (N_1295,In_2778,In_2045);
and U1296 (N_1296,In_106,In_2784);
and U1297 (N_1297,In_654,In_1972);
nor U1298 (N_1298,In_1764,In_682);
nand U1299 (N_1299,In_2562,In_929);
nor U1300 (N_1300,In_78,In_2385);
or U1301 (N_1301,In_2924,In_955);
or U1302 (N_1302,In_501,In_479);
and U1303 (N_1303,In_218,In_1163);
nand U1304 (N_1304,In_2438,In_2486);
nor U1305 (N_1305,In_2499,In_1398);
or U1306 (N_1306,In_1593,In_1719);
nor U1307 (N_1307,In_2655,In_1034);
or U1308 (N_1308,In_150,In_454);
xnor U1309 (N_1309,In_67,In_1783);
and U1310 (N_1310,In_2118,In_2765);
nor U1311 (N_1311,In_893,In_2671);
and U1312 (N_1312,In_2589,In_1146);
nor U1313 (N_1313,In_2616,In_1839);
and U1314 (N_1314,In_2411,In_1089);
and U1315 (N_1315,In_1428,In_2954);
and U1316 (N_1316,In_1565,In_1396);
xnor U1317 (N_1317,In_147,In_263);
nor U1318 (N_1318,In_275,In_1947);
xnor U1319 (N_1319,In_1317,In_1447);
or U1320 (N_1320,In_1184,In_1917);
nand U1321 (N_1321,In_321,In_121);
nand U1322 (N_1322,In_2289,In_2350);
or U1323 (N_1323,In_691,In_1979);
nor U1324 (N_1324,In_1419,In_2178);
xnor U1325 (N_1325,In_1753,In_664);
xnor U1326 (N_1326,In_460,In_2002);
nor U1327 (N_1327,In_2190,In_1583);
xor U1328 (N_1328,In_1384,In_2452);
nand U1329 (N_1329,In_1465,In_2777);
nor U1330 (N_1330,In_2301,In_2134);
xnor U1331 (N_1331,In_2282,In_2142);
nand U1332 (N_1332,In_702,In_53);
nor U1333 (N_1333,In_48,In_450);
xnor U1334 (N_1334,In_601,In_1055);
or U1335 (N_1335,In_189,In_1590);
and U1336 (N_1336,In_1322,In_316);
nand U1337 (N_1337,In_2324,In_403);
xor U1338 (N_1338,In_418,In_2908);
and U1339 (N_1339,In_2131,In_1798);
or U1340 (N_1340,In_1779,In_1648);
nand U1341 (N_1341,In_914,In_1868);
or U1342 (N_1342,In_2017,In_2032);
nand U1343 (N_1343,In_2376,In_216);
or U1344 (N_1344,In_1909,In_2494);
nand U1345 (N_1345,In_627,In_2490);
nand U1346 (N_1346,In_1335,In_2105);
nor U1347 (N_1347,In_2932,In_2483);
or U1348 (N_1348,In_1164,In_1982);
nor U1349 (N_1349,In_92,In_63);
xnor U1350 (N_1350,In_1528,In_1475);
or U1351 (N_1351,In_270,In_255);
or U1352 (N_1352,In_2522,In_36);
or U1353 (N_1353,In_1471,In_832);
nand U1354 (N_1354,In_774,In_127);
xor U1355 (N_1355,In_1989,In_164);
nand U1356 (N_1356,In_2115,In_2088);
nor U1357 (N_1357,In_2468,In_2338);
nand U1358 (N_1358,In_2591,In_2657);
xor U1359 (N_1359,In_2437,In_2621);
and U1360 (N_1360,In_1766,In_1102);
or U1361 (N_1361,In_91,In_444);
and U1362 (N_1362,In_2611,In_194);
nand U1363 (N_1363,In_1739,In_1068);
xnor U1364 (N_1364,In_2840,In_2707);
nor U1365 (N_1365,In_2710,In_2410);
nor U1366 (N_1366,In_2998,In_819);
nand U1367 (N_1367,In_1191,In_2720);
xnor U1368 (N_1368,In_1968,In_2018);
nor U1369 (N_1369,In_1052,In_762);
nand U1370 (N_1370,In_954,In_2420);
nand U1371 (N_1371,In_813,In_284);
xnor U1372 (N_1372,In_2934,In_1715);
nor U1373 (N_1373,In_1935,In_1810);
xnor U1374 (N_1374,In_1085,In_1692);
or U1375 (N_1375,In_1430,In_2742);
nand U1376 (N_1376,In_2938,In_2117);
or U1377 (N_1377,In_2265,In_2311);
nand U1378 (N_1378,In_589,In_731);
nor U1379 (N_1379,In_1844,In_2541);
and U1380 (N_1380,In_96,In_926);
and U1381 (N_1381,In_833,In_643);
and U1382 (N_1382,In_2815,In_310);
nand U1383 (N_1383,In_1843,In_61);
and U1384 (N_1384,In_958,In_451);
or U1385 (N_1385,In_1488,In_1253);
xor U1386 (N_1386,In_2920,In_2337);
or U1387 (N_1387,In_2283,In_1775);
or U1388 (N_1388,In_1519,In_2943);
nand U1389 (N_1389,In_84,In_855);
xor U1390 (N_1390,In_905,In_561);
or U1391 (N_1391,In_336,In_475);
and U1392 (N_1392,In_853,In_2043);
nand U1393 (N_1393,In_1409,In_380);
and U1394 (N_1394,In_1757,In_1059);
or U1395 (N_1395,In_611,In_925);
and U1396 (N_1396,In_2905,In_315);
nor U1397 (N_1397,In_393,In_423);
and U1398 (N_1398,In_661,In_2401);
and U1399 (N_1399,In_2930,In_2999);
nor U1400 (N_1400,In_2834,In_192);
or U1401 (N_1401,In_1536,In_2520);
nor U1402 (N_1402,In_2296,In_993);
nor U1403 (N_1403,In_2415,In_626);
nor U1404 (N_1404,In_843,In_653);
nor U1405 (N_1405,In_2167,In_1);
nand U1406 (N_1406,In_2383,In_2965);
nand U1407 (N_1407,In_1418,In_1802);
or U1408 (N_1408,In_898,In_188);
nor U1409 (N_1409,In_1871,In_668);
xor U1410 (N_1410,In_2016,In_1858);
or U1411 (N_1411,In_1469,In_2822);
nand U1412 (N_1412,In_419,In_886);
nand U1413 (N_1413,In_2412,In_212);
nand U1414 (N_1414,In_1861,In_468);
nand U1415 (N_1415,In_2782,In_1170);
nor U1416 (N_1416,In_1671,In_2988);
or U1417 (N_1417,In_2421,In_130);
or U1418 (N_1418,In_1225,In_971);
nor U1419 (N_1419,In_71,In_2701);
nand U1420 (N_1420,In_1302,In_2948);
nand U1421 (N_1421,In_2669,In_2160);
and U1422 (N_1422,In_2521,In_2592);
xor U1423 (N_1423,In_2872,In_2444);
xor U1424 (N_1424,In_1879,In_2953);
nor U1425 (N_1425,In_1136,In_579);
or U1426 (N_1426,In_967,In_2325);
or U1427 (N_1427,In_1696,In_1589);
or U1428 (N_1428,In_2614,In_2530);
or U1429 (N_1429,In_2033,In_2052);
nor U1430 (N_1430,In_555,In_1439);
xor U1431 (N_1431,In_1328,In_634);
nor U1432 (N_1432,In_1221,In_1721);
nor U1433 (N_1433,In_778,In_2843);
and U1434 (N_1434,In_2209,In_1258);
or U1435 (N_1435,In_2453,In_2065);
xor U1436 (N_1436,In_1128,In_2455);
or U1437 (N_1437,In_945,In_184);
xor U1438 (N_1438,In_2247,In_2243);
nand U1439 (N_1439,In_417,In_997);
and U1440 (N_1440,In_443,In_500);
nand U1441 (N_1441,In_2804,In_2069);
nor U1442 (N_1442,In_309,In_402);
or U1443 (N_1443,In_1449,In_124);
and U1444 (N_1444,In_1898,In_1494);
xor U1445 (N_1445,In_1808,In_622);
nor U1446 (N_1446,In_567,In_1997);
or U1447 (N_1447,In_800,In_1130);
nor U1448 (N_1448,In_2597,In_1611);
or U1449 (N_1449,In_1483,In_2071);
xor U1450 (N_1450,In_232,In_1150);
and U1451 (N_1451,In_2491,In_1661);
xnor U1452 (N_1452,In_1815,In_1263);
and U1453 (N_1453,In_2617,In_1904);
or U1454 (N_1454,In_1015,In_2423);
xor U1455 (N_1455,In_2231,In_2634);
nor U1456 (N_1456,In_2060,In_1417);
xor U1457 (N_1457,In_1813,In_81);
xnor U1458 (N_1458,In_1390,In_1343);
nand U1459 (N_1459,In_1846,In_670);
or U1460 (N_1460,In_266,In_2317);
or U1461 (N_1461,In_1708,In_1867);
nor U1462 (N_1462,In_2049,In_2364);
and U1463 (N_1463,In_128,In_1763);
xnor U1464 (N_1464,In_2299,In_11);
or U1465 (N_1465,In_2553,In_1319);
xnor U1466 (N_1466,In_1728,In_2451);
xor U1467 (N_1467,In_1425,In_1445);
xor U1468 (N_1468,In_1787,In_596);
nor U1469 (N_1469,In_2579,In_1820);
or U1470 (N_1470,In_1995,In_2441);
nor U1471 (N_1471,In_724,In_2662);
and U1472 (N_1472,In_1730,In_339);
nand U1473 (N_1473,In_2064,In_1333);
nor U1474 (N_1474,In_388,In_1632);
or U1475 (N_1475,In_620,In_697);
or U1476 (N_1476,In_442,In_268);
nand U1477 (N_1477,In_272,In_2256);
or U1478 (N_1478,In_370,In_1683);
or U1479 (N_1479,In_2594,In_357);
and U1480 (N_1480,In_2797,In_678);
nand U1481 (N_1481,In_783,In_2849);
or U1482 (N_1482,In_1370,In_2006);
xor U1483 (N_1483,In_2632,In_1711);
and U1484 (N_1484,In_447,In_1309);
nor U1485 (N_1485,In_1911,In_371);
and U1486 (N_1486,In_674,In_1139);
or U1487 (N_1487,In_1560,In_851);
and U1488 (N_1488,In_2526,In_1354);
and U1489 (N_1489,In_1046,In_590);
or U1490 (N_1490,In_2636,In_1703);
nor U1491 (N_1491,In_190,In_19);
nand U1492 (N_1492,In_2394,In_2048);
nand U1493 (N_1493,In_1727,In_2202);
xor U1494 (N_1494,In_1042,In_2968);
or U1495 (N_1495,In_462,In_1403);
or U1496 (N_1496,In_1036,In_1269);
or U1497 (N_1497,In_2086,In_720);
nor U1498 (N_1498,In_432,In_1896);
nand U1499 (N_1499,In_1897,In_717);
and U1500 (N_1500,In_1297,In_2538);
or U1501 (N_1501,In_2831,In_336);
xnor U1502 (N_1502,In_1268,In_1861);
and U1503 (N_1503,In_552,In_99);
xor U1504 (N_1504,In_1261,In_996);
and U1505 (N_1505,In_2041,In_317);
xor U1506 (N_1506,In_2413,In_2608);
nand U1507 (N_1507,In_2964,In_1769);
nor U1508 (N_1508,In_1594,In_184);
xnor U1509 (N_1509,In_1728,In_1363);
nand U1510 (N_1510,In_1741,In_1064);
and U1511 (N_1511,In_558,In_517);
nor U1512 (N_1512,In_2145,In_924);
xor U1513 (N_1513,In_2500,In_643);
xor U1514 (N_1514,In_1295,In_358);
nand U1515 (N_1515,In_999,In_75);
or U1516 (N_1516,In_1036,In_1433);
and U1517 (N_1517,In_1021,In_121);
or U1518 (N_1518,In_2986,In_493);
nand U1519 (N_1519,In_2292,In_2358);
and U1520 (N_1520,In_2990,In_2306);
or U1521 (N_1521,In_1966,In_1336);
nor U1522 (N_1522,In_1896,In_2758);
or U1523 (N_1523,In_765,In_823);
and U1524 (N_1524,In_503,In_2376);
and U1525 (N_1525,In_1111,In_1899);
xor U1526 (N_1526,In_1920,In_1502);
and U1527 (N_1527,In_2440,In_2512);
or U1528 (N_1528,In_1921,In_1942);
xor U1529 (N_1529,In_552,In_1122);
or U1530 (N_1530,In_2482,In_393);
or U1531 (N_1531,In_1929,In_2055);
nor U1532 (N_1532,In_2105,In_931);
and U1533 (N_1533,In_2399,In_1105);
or U1534 (N_1534,In_1875,In_2278);
xor U1535 (N_1535,In_1115,In_2371);
or U1536 (N_1536,In_1362,In_2703);
xor U1537 (N_1537,In_1,In_1926);
or U1538 (N_1538,In_2590,In_585);
and U1539 (N_1539,In_134,In_2855);
nand U1540 (N_1540,In_2012,In_1966);
xor U1541 (N_1541,In_2069,In_1903);
and U1542 (N_1542,In_2688,In_185);
nand U1543 (N_1543,In_2558,In_1683);
nor U1544 (N_1544,In_212,In_1816);
xnor U1545 (N_1545,In_2341,In_2029);
nand U1546 (N_1546,In_2132,In_2765);
xnor U1547 (N_1547,In_2751,In_2541);
or U1548 (N_1548,In_1107,In_2770);
nor U1549 (N_1549,In_487,In_1495);
nand U1550 (N_1550,In_1852,In_1066);
or U1551 (N_1551,In_2895,In_578);
nor U1552 (N_1552,In_2692,In_1517);
and U1553 (N_1553,In_275,In_1534);
nor U1554 (N_1554,In_2454,In_2090);
and U1555 (N_1555,In_1015,In_2144);
nand U1556 (N_1556,In_2380,In_2658);
or U1557 (N_1557,In_2302,In_1044);
nand U1558 (N_1558,In_2613,In_696);
and U1559 (N_1559,In_2170,In_341);
and U1560 (N_1560,In_1192,In_1586);
nor U1561 (N_1561,In_495,In_1171);
xnor U1562 (N_1562,In_240,In_219);
nor U1563 (N_1563,In_698,In_1184);
or U1564 (N_1564,In_615,In_1135);
or U1565 (N_1565,In_1189,In_918);
nand U1566 (N_1566,In_1711,In_1103);
nand U1567 (N_1567,In_864,In_1581);
nor U1568 (N_1568,In_662,In_1407);
xnor U1569 (N_1569,In_1221,In_2987);
or U1570 (N_1570,In_1306,In_1357);
nand U1571 (N_1571,In_2825,In_2743);
xnor U1572 (N_1572,In_1195,In_668);
nor U1573 (N_1573,In_933,In_1691);
xnor U1574 (N_1574,In_855,In_2693);
or U1575 (N_1575,In_164,In_2132);
nand U1576 (N_1576,In_1703,In_1125);
or U1577 (N_1577,In_2165,In_1369);
xnor U1578 (N_1578,In_375,In_2970);
xnor U1579 (N_1579,In_2596,In_1251);
and U1580 (N_1580,In_566,In_2775);
or U1581 (N_1581,In_254,In_971);
nand U1582 (N_1582,In_1515,In_1989);
nand U1583 (N_1583,In_1947,In_1396);
nor U1584 (N_1584,In_533,In_1354);
and U1585 (N_1585,In_2297,In_2982);
and U1586 (N_1586,In_1306,In_48);
and U1587 (N_1587,In_2650,In_747);
or U1588 (N_1588,In_56,In_1574);
or U1589 (N_1589,In_2559,In_1339);
xor U1590 (N_1590,In_1975,In_540);
xor U1591 (N_1591,In_545,In_566);
nand U1592 (N_1592,In_1823,In_2491);
nor U1593 (N_1593,In_2239,In_541);
nand U1594 (N_1594,In_2409,In_2301);
nor U1595 (N_1595,In_659,In_1361);
and U1596 (N_1596,In_475,In_111);
and U1597 (N_1597,In_151,In_1370);
xnor U1598 (N_1598,In_1059,In_1895);
xnor U1599 (N_1599,In_1065,In_1799);
xor U1600 (N_1600,In_910,In_1553);
nor U1601 (N_1601,In_2400,In_1079);
and U1602 (N_1602,In_378,In_1346);
nand U1603 (N_1603,In_2932,In_649);
nand U1604 (N_1604,In_2566,In_1323);
xor U1605 (N_1605,In_1666,In_133);
and U1606 (N_1606,In_201,In_1287);
nor U1607 (N_1607,In_2401,In_2975);
nand U1608 (N_1608,In_831,In_445);
nand U1609 (N_1609,In_2975,In_814);
or U1610 (N_1610,In_768,In_1133);
xor U1611 (N_1611,In_722,In_1826);
xor U1612 (N_1612,In_2058,In_2793);
xor U1613 (N_1613,In_259,In_2358);
and U1614 (N_1614,In_233,In_1314);
and U1615 (N_1615,In_2252,In_611);
xor U1616 (N_1616,In_660,In_2818);
nand U1617 (N_1617,In_2254,In_1376);
nand U1618 (N_1618,In_2183,In_1144);
or U1619 (N_1619,In_1989,In_1995);
or U1620 (N_1620,In_1700,In_1672);
and U1621 (N_1621,In_2102,In_2402);
nand U1622 (N_1622,In_73,In_1598);
xnor U1623 (N_1623,In_470,In_537);
nor U1624 (N_1624,In_2877,In_1033);
xor U1625 (N_1625,In_824,In_2399);
and U1626 (N_1626,In_1016,In_2155);
xnor U1627 (N_1627,In_808,In_1770);
nor U1628 (N_1628,In_1256,In_1280);
nor U1629 (N_1629,In_2631,In_1606);
xor U1630 (N_1630,In_2963,In_614);
or U1631 (N_1631,In_2921,In_421);
nor U1632 (N_1632,In_2381,In_604);
nand U1633 (N_1633,In_373,In_1454);
nor U1634 (N_1634,In_532,In_1505);
nand U1635 (N_1635,In_2549,In_884);
and U1636 (N_1636,In_1690,In_1163);
or U1637 (N_1637,In_1821,In_2867);
and U1638 (N_1638,In_1768,In_112);
xnor U1639 (N_1639,In_2641,In_1852);
nand U1640 (N_1640,In_2561,In_1886);
or U1641 (N_1641,In_1680,In_2711);
and U1642 (N_1642,In_1669,In_2072);
xor U1643 (N_1643,In_2140,In_56);
or U1644 (N_1644,In_1424,In_2896);
xnor U1645 (N_1645,In_1330,In_993);
nand U1646 (N_1646,In_2218,In_2422);
and U1647 (N_1647,In_1435,In_445);
nor U1648 (N_1648,In_2178,In_2027);
or U1649 (N_1649,In_1235,In_1364);
nand U1650 (N_1650,In_322,In_2991);
or U1651 (N_1651,In_629,In_1046);
or U1652 (N_1652,In_547,In_1474);
or U1653 (N_1653,In_1953,In_1893);
nor U1654 (N_1654,In_2710,In_925);
xnor U1655 (N_1655,In_587,In_1726);
and U1656 (N_1656,In_138,In_1336);
nand U1657 (N_1657,In_657,In_2421);
and U1658 (N_1658,In_61,In_142);
and U1659 (N_1659,In_176,In_413);
or U1660 (N_1660,In_2851,In_2679);
nand U1661 (N_1661,In_48,In_2923);
nand U1662 (N_1662,In_1873,In_672);
xnor U1663 (N_1663,In_1833,In_1215);
nand U1664 (N_1664,In_2810,In_1817);
and U1665 (N_1665,In_2653,In_289);
nand U1666 (N_1666,In_2405,In_329);
nor U1667 (N_1667,In_1788,In_1270);
nand U1668 (N_1668,In_2066,In_1712);
xor U1669 (N_1669,In_1933,In_1544);
or U1670 (N_1670,In_1728,In_1526);
nand U1671 (N_1671,In_2615,In_665);
nor U1672 (N_1672,In_830,In_1878);
nand U1673 (N_1673,In_1585,In_700);
nand U1674 (N_1674,In_1741,In_1568);
xor U1675 (N_1675,In_1492,In_701);
and U1676 (N_1676,In_2077,In_1162);
xnor U1677 (N_1677,In_504,In_1590);
xnor U1678 (N_1678,In_1163,In_1784);
xnor U1679 (N_1679,In_696,In_2395);
xor U1680 (N_1680,In_452,In_324);
nor U1681 (N_1681,In_2511,In_411);
or U1682 (N_1682,In_1362,In_1824);
and U1683 (N_1683,In_280,In_1101);
nor U1684 (N_1684,In_2638,In_2125);
xor U1685 (N_1685,In_2556,In_1603);
and U1686 (N_1686,In_925,In_2795);
and U1687 (N_1687,In_1052,In_1992);
nand U1688 (N_1688,In_641,In_20);
and U1689 (N_1689,In_275,In_996);
nand U1690 (N_1690,In_930,In_1590);
and U1691 (N_1691,In_2545,In_1771);
or U1692 (N_1692,In_1809,In_1671);
nand U1693 (N_1693,In_2025,In_928);
and U1694 (N_1694,In_2050,In_2089);
and U1695 (N_1695,In_1377,In_405);
and U1696 (N_1696,In_2729,In_303);
nand U1697 (N_1697,In_2804,In_1343);
or U1698 (N_1698,In_1157,In_1467);
and U1699 (N_1699,In_2352,In_1552);
xnor U1700 (N_1700,In_2778,In_1469);
or U1701 (N_1701,In_2330,In_1916);
xnor U1702 (N_1702,In_2355,In_1732);
xnor U1703 (N_1703,In_814,In_877);
or U1704 (N_1704,In_1832,In_2961);
and U1705 (N_1705,In_576,In_520);
xor U1706 (N_1706,In_632,In_2229);
or U1707 (N_1707,In_726,In_2282);
nand U1708 (N_1708,In_1692,In_1983);
and U1709 (N_1709,In_2793,In_2155);
or U1710 (N_1710,In_1552,In_1810);
xor U1711 (N_1711,In_1289,In_1957);
and U1712 (N_1712,In_397,In_2466);
nor U1713 (N_1713,In_1033,In_1127);
xnor U1714 (N_1714,In_2895,In_2883);
nor U1715 (N_1715,In_286,In_1328);
nor U1716 (N_1716,In_786,In_2836);
or U1717 (N_1717,In_809,In_2851);
or U1718 (N_1718,In_2892,In_346);
or U1719 (N_1719,In_1420,In_2728);
and U1720 (N_1720,In_2993,In_143);
and U1721 (N_1721,In_586,In_1219);
xnor U1722 (N_1722,In_367,In_258);
xnor U1723 (N_1723,In_462,In_2683);
nor U1724 (N_1724,In_2243,In_1679);
xor U1725 (N_1725,In_2859,In_295);
nor U1726 (N_1726,In_2971,In_877);
nand U1727 (N_1727,In_1308,In_1543);
and U1728 (N_1728,In_1893,In_2922);
or U1729 (N_1729,In_383,In_2321);
nor U1730 (N_1730,In_2454,In_1133);
xnor U1731 (N_1731,In_902,In_1937);
nor U1732 (N_1732,In_1572,In_349);
nor U1733 (N_1733,In_66,In_2606);
nand U1734 (N_1734,In_996,In_1219);
nand U1735 (N_1735,In_642,In_97);
xnor U1736 (N_1736,In_1455,In_1759);
and U1737 (N_1737,In_2791,In_376);
xnor U1738 (N_1738,In_40,In_2409);
nor U1739 (N_1739,In_2463,In_1872);
or U1740 (N_1740,In_1592,In_2080);
and U1741 (N_1741,In_1828,In_546);
nor U1742 (N_1742,In_2884,In_1253);
and U1743 (N_1743,In_1345,In_1711);
and U1744 (N_1744,In_1684,In_363);
and U1745 (N_1745,In_2661,In_2086);
nor U1746 (N_1746,In_1550,In_1755);
xor U1747 (N_1747,In_1146,In_2505);
or U1748 (N_1748,In_443,In_2441);
or U1749 (N_1749,In_901,In_1017);
or U1750 (N_1750,In_2664,In_2992);
and U1751 (N_1751,In_1862,In_2025);
or U1752 (N_1752,In_2494,In_2119);
nor U1753 (N_1753,In_1876,In_2192);
xor U1754 (N_1754,In_561,In_50);
nand U1755 (N_1755,In_2860,In_1006);
and U1756 (N_1756,In_590,In_249);
and U1757 (N_1757,In_1362,In_2515);
and U1758 (N_1758,In_1610,In_2099);
nor U1759 (N_1759,In_2318,In_356);
nand U1760 (N_1760,In_2678,In_2681);
and U1761 (N_1761,In_354,In_1145);
nand U1762 (N_1762,In_437,In_2176);
xor U1763 (N_1763,In_2852,In_472);
and U1764 (N_1764,In_2832,In_2888);
nor U1765 (N_1765,In_791,In_2079);
nand U1766 (N_1766,In_1011,In_2016);
nor U1767 (N_1767,In_1486,In_1954);
nor U1768 (N_1768,In_150,In_2836);
nand U1769 (N_1769,In_2683,In_528);
nand U1770 (N_1770,In_636,In_329);
and U1771 (N_1771,In_1731,In_1615);
nand U1772 (N_1772,In_2057,In_1652);
xor U1773 (N_1773,In_346,In_1198);
nor U1774 (N_1774,In_2401,In_1552);
nand U1775 (N_1775,In_2688,In_351);
nor U1776 (N_1776,In_791,In_1268);
nor U1777 (N_1777,In_1710,In_666);
xor U1778 (N_1778,In_2154,In_2827);
and U1779 (N_1779,In_960,In_2503);
and U1780 (N_1780,In_1541,In_1034);
nor U1781 (N_1781,In_2246,In_1546);
nand U1782 (N_1782,In_1198,In_974);
nor U1783 (N_1783,In_309,In_2516);
nand U1784 (N_1784,In_1347,In_1846);
xnor U1785 (N_1785,In_1483,In_2919);
and U1786 (N_1786,In_369,In_2724);
nand U1787 (N_1787,In_1261,In_1991);
or U1788 (N_1788,In_259,In_1868);
nand U1789 (N_1789,In_1407,In_1309);
nand U1790 (N_1790,In_4,In_556);
xnor U1791 (N_1791,In_1030,In_1763);
or U1792 (N_1792,In_2049,In_1199);
xor U1793 (N_1793,In_1822,In_484);
xor U1794 (N_1794,In_1036,In_142);
and U1795 (N_1795,In_1718,In_1399);
nand U1796 (N_1796,In_808,In_2749);
nand U1797 (N_1797,In_2355,In_521);
or U1798 (N_1798,In_621,In_2943);
nor U1799 (N_1799,In_1969,In_1045);
or U1800 (N_1800,In_1481,In_2524);
nor U1801 (N_1801,In_1599,In_25);
or U1802 (N_1802,In_2201,In_1976);
xnor U1803 (N_1803,In_1416,In_2670);
or U1804 (N_1804,In_588,In_2104);
xnor U1805 (N_1805,In_2821,In_2492);
nand U1806 (N_1806,In_1252,In_2776);
nor U1807 (N_1807,In_2134,In_890);
or U1808 (N_1808,In_22,In_409);
nand U1809 (N_1809,In_2049,In_1229);
xnor U1810 (N_1810,In_2979,In_42);
nand U1811 (N_1811,In_539,In_2159);
nand U1812 (N_1812,In_1572,In_2771);
and U1813 (N_1813,In_2560,In_145);
xnor U1814 (N_1814,In_2005,In_2514);
xor U1815 (N_1815,In_1148,In_2648);
and U1816 (N_1816,In_130,In_1899);
nor U1817 (N_1817,In_1092,In_959);
xor U1818 (N_1818,In_1864,In_1747);
nand U1819 (N_1819,In_2476,In_1921);
nor U1820 (N_1820,In_1756,In_1833);
or U1821 (N_1821,In_2183,In_1050);
or U1822 (N_1822,In_640,In_2244);
or U1823 (N_1823,In_1074,In_2446);
and U1824 (N_1824,In_178,In_2498);
nor U1825 (N_1825,In_1357,In_2815);
or U1826 (N_1826,In_2422,In_2720);
xnor U1827 (N_1827,In_1341,In_2683);
and U1828 (N_1828,In_2400,In_444);
or U1829 (N_1829,In_512,In_71);
nor U1830 (N_1830,In_1494,In_1725);
or U1831 (N_1831,In_2950,In_1321);
xor U1832 (N_1832,In_483,In_280);
or U1833 (N_1833,In_1724,In_1637);
nor U1834 (N_1834,In_40,In_968);
and U1835 (N_1835,In_69,In_1355);
nor U1836 (N_1836,In_1700,In_2292);
or U1837 (N_1837,In_1485,In_2619);
and U1838 (N_1838,In_2962,In_1701);
nand U1839 (N_1839,In_414,In_1494);
nand U1840 (N_1840,In_607,In_2958);
or U1841 (N_1841,In_1509,In_2476);
nor U1842 (N_1842,In_1619,In_1165);
nor U1843 (N_1843,In_82,In_2285);
nor U1844 (N_1844,In_2523,In_703);
xor U1845 (N_1845,In_2918,In_1122);
or U1846 (N_1846,In_2210,In_2174);
and U1847 (N_1847,In_436,In_1455);
xor U1848 (N_1848,In_2694,In_112);
or U1849 (N_1849,In_767,In_1982);
nand U1850 (N_1850,In_1777,In_2686);
and U1851 (N_1851,In_2297,In_1106);
xor U1852 (N_1852,In_319,In_1777);
nand U1853 (N_1853,In_174,In_2613);
or U1854 (N_1854,In_710,In_907);
xnor U1855 (N_1855,In_144,In_1805);
nor U1856 (N_1856,In_778,In_1379);
nand U1857 (N_1857,In_142,In_2518);
xor U1858 (N_1858,In_714,In_2259);
and U1859 (N_1859,In_1808,In_1226);
and U1860 (N_1860,In_627,In_2835);
or U1861 (N_1861,In_997,In_2813);
xnor U1862 (N_1862,In_1584,In_1054);
and U1863 (N_1863,In_2450,In_846);
and U1864 (N_1864,In_2307,In_2095);
and U1865 (N_1865,In_412,In_252);
xnor U1866 (N_1866,In_732,In_2593);
nor U1867 (N_1867,In_1170,In_1121);
nand U1868 (N_1868,In_1349,In_1148);
nand U1869 (N_1869,In_2582,In_2858);
nand U1870 (N_1870,In_122,In_260);
and U1871 (N_1871,In_2697,In_2499);
or U1872 (N_1872,In_4,In_2867);
or U1873 (N_1873,In_2310,In_1561);
or U1874 (N_1874,In_2219,In_424);
nand U1875 (N_1875,In_1867,In_1014);
nor U1876 (N_1876,In_2851,In_745);
nor U1877 (N_1877,In_2819,In_957);
xnor U1878 (N_1878,In_2290,In_2145);
xor U1879 (N_1879,In_171,In_2812);
nand U1880 (N_1880,In_2450,In_2324);
nand U1881 (N_1881,In_94,In_222);
xor U1882 (N_1882,In_286,In_1341);
nand U1883 (N_1883,In_2646,In_303);
and U1884 (N_1884,In_1058,In_1074);
nand U1885 (N_1885,In_2970,In_608);
xnor U1886 (N_1886,In_2872,In_703);
xnor U1887 (N_1887,In_1533,In_2685);
nor U1888 (N_1888,In_2461,In_1316);
and U1889 (N_1889,In_1699,In_1412);
and U1890 (N_1890,In_1595,In_456);
and U1891 (N_1891,In_346,In_2625);
and U1892 (N_1892,In_27,In_1169);
xor U1893 (N_1893,In_1083,In_2394);
nand U1894 (N_1894,In_1439,In_2622);
nand U1895 (N_1895,In_436,In_2347);
or U1896 (N_1896,In_1030,In_316);
or U1897 (N_1897,In_245,In_2125);
or U1898 (N_1898,In_2365,In_1098);
and U1899 (N_1899,In_2759,In_2270);
nand U1900 (N_1900,In_1569,In_2123);
and U1901 (N_1901,In_2843,In_2292);
nor U1902 (N_1902,In_1559,In_1236);
xnor U1903 (N_1903,In_2436,In_56);
xnor U1904 (N_1904,In_338,In_1702);
xnor U1905 (N_1905,In_2201,In_2068);
nand U1906 (N_1906,In_2392,In_1443);
nor U1907 (N_1907,In_831,In_2885);
xnor U1908 (N_1908,In_1991,In_2117);
or U1909 (N_1909,In_534,In_277);
and U1910 (N_1910,In_381,In_2585);
and U1911 (N_1911,In_2,In_2121);
and U1912 (N_1912,In_1418,In_240);
nand U1913 (N_1913,In_968,In_826);
xnor U1914 (N_1914,In_2890,In_2515);
or U1915 (N_1915,In_334,In_158);
xnor U1916 (N_1916,In_277,In_505);
nor U1917 (N_1917,In_1758,In_2032);
nor U1918 (N_1918,In_766,In_1956);
and U1919 (N_1919,In_5,In_2988);
or U1920 (N_1920,In_1582,In_2278);
xnor U1921 (N_1921,In_2987,In_1672);
or U1922 (N_1922,In_1453,In_480);
nor U1923 (N_1923,In_2757,In_1892);
nor U1924 (N_1924,In_2124,In_2706);
xnor U1925 (N_1925,In_1644,In_1324);
nor U1926 (N_1926,In_1279,In_1059);
nand U1927 (N_1927,In_2644,In_1075);
nor U1928 (N_1928,In_2054,In_1336);
or U1929 (N_1929,In_2931,In_326);
and U1930 (N_1930,In_689,In_927);
nor U1931 (N_1931,In_831,In_2279);
xor U1932 (N_1932,In_1390,In_2424);
and U1933 (N_1933,In_2998,In_1871);
xnor U1934 (N_1934,In_2104,In_741);
and U1935 (N_1935,In_2482,In_1798);
and U1936 (N_1936,In_1519,In_261);
xor U1937 (N_1937,In_1560,In_2075);
and U1938 (N_1938,In_1303,In_759);
and U1939 (N_1939,In_1810,In_1677);
xnor U1940 (N_1940,In_1610,In_1110);
and U1941 (N_1941,In_2623,In_632);
nand U1942 (N_1942,In_2286,In_1608);
and U1943 (N_1943,In_2029,In_2139);
and U1944 (N_1944,In_2913,In_834);
or U1945 (N_1945,In_598,In_388);
or U1946 (N_1946,In_2690,In_720);
or U1947 (N_1947,In_2141,In_1673);
xor U1948 (N_1948,In_2517,In_226);
and U1949 (N_1949,In_1240,In_2512);
and U1950 (N_1950,In_1599,In_2247);
nand U1951 (N_1951,In_2330,In_291);
or U1952 (N_1952,In_265,In_2989);
or U1953 (N_1953,In_2960,In_564);
nor U1954 (N_1954,In_1937,In_2288);
or U1955 (N_1955,In_2066,In_2866);
nor U1956 (N_1956,In_1620,In_1463);
or U1957 (N_1957,In_2204,In_475);
nor U1958 (N_1958,In_2370,In_530);
nor U1959 (N_1959,In_538,In_807);
and U1960 (N_1960,In_984,In_1438);
xnor U1961 (N_1961,In_967,In_1372);
nand U1962 (N_1962,In_1943,In_2478);
xnor U1963 (N_1963,In_675,In_1745);
nor U1964 (N_1964,In_1559,In_2196);
xnor U1965 (N_1965,In_2783,In_141);
and U1966 (N_1966,In_436,In_2277);
xor U1967 (N_1967,In_510,In_1432);
xnor U1968 (N_1968,In_2140,In_546);
or U1969 (N_1969,In_2214,In_1615);
or U1970 (N_1970,In_95,In_1509);
nor U1971 (N_1971,In_2130,In_731);
nor U1972 (N_1972,In_744,In_1892);
or U1973 (N_1973,In_2880,In_1576);
and U1974 (N_1974,In_280,In_2279);
xnor U1975 (N_1975,In_1089,In_1115);
and U1976 (N_1976,In_817,In_2635);
or U1977 (N_1977,In_1873,In_338);
or U1978 (N_1978,In_835,In_2572);
xor U1979 (N_1979,In_1521,In_1080);
or U1980 (N_1980,In_873,In_2317);
nand U1981 (N_1981,In_1529,In_1797);
nand U1982 (N_1982,In_850,In_763);
nor U1983 (N_1983,In_2522,In_1102);
xnor U1984 (N_1984,In_1867,In_249);
nand U1985 (N_1985,In_2530,In_1351);
and U1986 (N_1986,In_1649,In_1981);
and U1987 (N_1987,In_708,In_135);
or U1988 (N_1988,In_1725,In_1105);
nor U1989 (N_1989,In_1142,In_1463);
and U1990 (N_1990,In_1713,In_2189);
or U1991 (N_1991,In_1078,In_1330);
nor U1992 (N_1992,In_1962,In_1893);
and U1993 (N_1993,In_2058,In_2790);
nand U1994 (N_1994,In_976,In_2150);
nor U1995 (N_1995,In_2802,In_433);
nand U1996 (N_1996,In_317,In_2543);
xor U1997 (N_1997,In_2418,In_2405);
nand U1998 (N_1998,In_268,In_676);
nor U1999 (N_1999,In_2742,In_2486);
and U2000 (N_2000,In_185,In_173);
or U2001 (N_2001,In_733,In_89);
nor U2002 (N_2002,In_1575,In_908);
xnor U2003 (N_2003,In_119,In_693);
or U2004 (N_2004,In_1985,In_92);
nand U2005 (N_2005,In_2320,In_26);
nor U2006 (N_2006,In_2966,In_880);
xor U2007 (N_2007,In_7,In_8);
nand U2008 (N_2008,In_582,In_254);
xnor U2009 (N_2009,In_1330,In_2357);
nand U2010 (N_2010,In_1336,In_749);
and U2011 (N_2011,In_765,In_1621);
or U2012 (N_2012,In_2480,In_480);
nor U2013 (N_2013,In_1378,In_2900);
nor U2014 (N_2014,In_2234,In_1980);
and U2015 (N_2015,In_2798,In_681);
or U2016 (N_2016,In_499,In_1916);
and U2017 (N_2017,In_1203,In_283);
and U2018 (N_2018,In_1777,In_2577);
or U2019 (N_2019,In_706,In_2623);
xor U2020 (N_2020,In_481,In_1916);
or U2021 (N_2021,In_1603,In_2827);
and U2022 (N_2022,In_2221,In_2898);
xor U2023 (N_2023,In_2648,In_2553);
nand U2024 (N_2024,In_1507,In_2380);
or U2025 (N_2025,In_2662,In_1813);
and U2026 (N_2026,In_576,In_2385);
nor U2027 (N_2027,In_281,In_1742);
nor U2028 (N_2028,In_2636,In_276);
nor U2029 (N_2029,In_1784,In_558);
or U2030 (N_2030,In_926,In_1058);
nor U2031 (N_2031,In_451,In_1060);
nand U2032 (N_2032,In_2046,In_1436);
nor U2033 (N_2033,In_2657,In_2626);
nand U2034 (N_2034,In_240,In_124);
nand U2035 (N_2035,In_299,In_1897);
nand U2036 (N_2036,In_131,In_1268);
or U2037 (N_2037,In_1126,In_1531);
nand U2038 (N_2038,In_499,In_2533);
nor U2039 (N_2039,In_1091,In_2468);
or U2040 (N_2040,In_1247,In_713);
and U2041 (N_2041,In_1236,In_1670);
nor U2042 (N_2042,In_1971,In_2545);
and U2043 (N_2043,In_308,In_1563);
and U2044 (N_2044,In_1257,In_2914);
nor U2045 (N_2045,In_955,In_2564);
and U2046 (N_2046,In_697,In_2041);
nor U2047 (N_2047,In_2983,In_960);
nand U2048 (N_2048,In_859,In_1134);
xnor U2049 (N_2049,In_701,In_91);
or U2050 (N_2050,In_1303,In_544);
nor U2051 (N_2051,In_661,In_1977);
nor U2052 (N_2052,In_1238,In_2164);
nor U2053 (N_2053,In_2814,In_1957);
or U2054 (N_2054,In_320,In_2564);
xor U2055 (N_2055,In_1991,In_1050);
or U2056 (N_2056,In_275,In_453);
nor U2057 (N_2057,In_2936,In_2154);
nor U2058 (N_2058,In_1928,In_1237);
nor U2059 (N_2059,In_1110,In_1426);
xnor U2060 (N_2060,In_539,In_1121);
nand U2061 (N_2061,In_505,In_1668);
nor U2062 (N_2062,In_2946,In_1607);
nor U2063 (N_2063,In_2266,In_458);
and U2064 (N_2064,In_283,In_2375);
or U2065 (N_2065,In_491,In_1962);
xor U2066 (N_2066,In_354,In_2014);
nor U2067 (N_2067,In_1714,In_2662);
nor U2068 (N_2068,In_1247,In_686);
xor U2069 (N_2069,In_1067,In_1280);
and U2070 (N_2070,In_317,In_720);
nand U2071 (N_2071,In_173,In_870);
and U2072 (N_2072,In_1161,In_2495);
xor U2073 (N_2073,In_2952,In_699);
or U2074 (N_2074,In_867,In_2018);
nand U2075 (N_2075,In_2518,In_2952);
nand U2076 (N_2076,In_2251,In_2303);
and U2077 (N_2077,In_781,In_1033);
nor U2078 (N_2078,In_1678,In_842);
nand U2079 (N_2079,In_1932,In_886);
or U2080 (N_2080,In_1764,In_124);
nand U2081 (N_2081,In_860,In_1485);
nand U2082 (N_2082,In_1899,In_1279);
or U2083 (N_2083,In_2202,In_690);
nor U2084 (N_2084,In_2070,In_608);
and U2085 (N_2085,In_1662,In_1727);
nand U2086 (N_2086,In_362,In_1969);
xnor U2087 (N_2087,In_1719,In_1210);
nand U2088 (N_2088,In_285,In_2850);
xnor U2089 (N_2089,In_2015,In_1180);
xor U2090 (N_2090,In_2043,In_1825);
xor U2091 (N_2091,In_2077,In_370);
and U2092 (N_2092,In_460,In_2281);
nand U2093 (N_2093,In_699,In_2136);
or U2094 (N_2094,In_1650,In_389);
nand U2095 (N_2095,In_2843,In_2918);
and U2096 (N_2096,In_881,In_1709);
xor U2097 (N_2097,In_1016,In_44);
nand U2098 (N_2098,In_1598,In_265);
nor U2099 (N_2099,In_795,In_1233);
nor U2100 (N_2100,In_2115,In_2433);
or U2101 (N_2101,In_1035,In_68);
xor U2102 (N_2102,In_981,In_1664);
nand U2103 (N_2103,In_937,In_2352);
nand U2104 (N_2104,In_1392,In_1725);
nand U2105 (N_2105,In_1624,In_2303);
nand U2106 (N_2106,In_2067,In_1809);
nand U2107 (N_2107,In_2347,In_493);
and U2108 (N_2108,In_531,In_902);
nor U2109 (N_2109,In_50,In_2649);
and U2110 (N_2110,In_749,In_1953);
or U2111 (N_2111,In_1727,In_1491);
and U2112 (N_2112,In_2275,In_2716);
nor U2113 (N_2113,In_135,In_2435);
and U2114 (N_2114,In_2273,In_579);
xor U2115 (N_2115,In_2179,In_2775);
or U2116 (N_2116,In_283,In_2176);
or U2117 (N_2117,In_2081,In_2781);
nand U2118 (N_2118,In_356,In_2886);
and U2119 (N_2119,In_809,In_294);
nand U2120 (N_2120,In_2986,In_411);
nand U2121 (N_2121,In_1237,In_2369);
xnor U2122 (N_2122,In_2458,In_1397);
nand U2123 (N_2123,In_1837,In_2975);
nand U2124 (N_2124,In_2614,In_1026);
nand U2125 (N_2125,In_2565,In_2471);
nand U2126 (N_2126,In_1556,In_461);
and U2127 (N_2127,In_2771,In_601);
xor U2128 (N_2128,In_1177,In_1982);
nand U2129 (N_2129,In_1363,In_42);
xor U2130 (N_2130,In_64,In_571);
and U2131 (N_2131,In_1847,In_1088);
nor U2132 (N_2132,In_581,In_523);
and U2133 (N_2133,In_376,In_900);
xor U2134 (N_2134,In_2348,In_1230);
nor U2135 (N_2135,In_1587,In_2864);
and U2136 (N_2136,In_1753,In_1180);
or U2137 (N_2137,In_571,In_450);
or U2138 (N_2138,In_2859,In_2874);
or U2139 (N_2139,In_2397,In_2606);
nand U2140 (N_2140,In_1152,In_1715);
or U2141 (N_2141,In_2377,In_2084);
or U2142 (N_2142,In_2256,In_77);
nand U2143 (N_2143,In_1740,In_2207);
or U2144 (N_2144,In_2918,In_2711);
nand U2145 (N_2145,In_1949,In_2456);
xor U2146 (N_2146,In_2326,In_244);
and U2147 (N_2147,In_674,In_223);
xnor U2148 (N_2148,In_2675,In_832);
or U2149 (N_2149,In_647,In_2614);
nand U2150 (N_2150,In_1007,In_631);
and U2151 (N_2151,In_1583,In_2603);
or U2152 (N_2152,In_1689,In_1471);
nor U2153 (N_2153,In_2599,In_1272);
nand U2154 (N_2154,In_254,In_2777);
and U2155 (N_2155,In_774,In_1980);
xor U2156 (N_2156,In_838,In_12);
nand U2157 (N_2157,In_2657,In_25);
nand U2158 (N_2158,In_1365,In_308);
nand U2159 (N_2159,In_835,In_1368);
nand U2160 (N_2160,In_2818,In_257);
or U2161 (N_2161,In_1366,In_2445);
or U2162 (N_2162,In_389,In_1786);
xnor U2163 (N_2163,In_847,In_2752);
or U2164 (N_2164,In_2056,In_1860);
and U2165 (N_2165,In_2512,In_535);
and U2166 (N_2166,In_2237,In_2443);
and U2167 (N_2167,In_1532,In_2848);
and U2168 (N_2168,In_1835,In_1891);
nand U2169 (N_2169,In_65,In_447);
nand U2170 (N_2170,In_1242,In_129);
or U2171 (N_2171,In_1330,In_86);
nand U2172 (N_2172,In_410,In_2220);
nor U2173 (N_2173,In_1990,In_1918);
or U2174 (N_2174,In_2417,In_2848);
and U2175 (N_2175,In_1443,In_242);
and U2176 (N_2176,In_2535,In_1516);
or U2177 (N_2177,In_636,In_957);
and U2178 (N_2178,In_65,In_1729);
xor U2179 (N_2179,In_838,In_2476);
nand U2180 (N_2180,In_1868,In_2005);
nor U2181 (N_2181,In_2575,In_924);
or U2182 (N_2182,In_1262,In_573);
or U2183 (N_2183,In_1547,In_1384);
or U2184 (N_2184,In_1473,In_1546);
nand U2185 (N_2185,In_2247,In_457);
nor U2186 (N_2186,In_2614,In_271);
or U2187 (N_2187,In_1415,In_76);
nor U2188 (N_2188,In_1953,In_68);
xor U2189 (N_2189,In_157,In_1466);
nor U2190 (N_2190,In_1578,In_688);
or U2191 (N_2191,In_544,In_134);
nand U2192 (N_2192,In_2099,In_1254);
nand U2193 (N_2193,In_2044,In_1310);
xor U2194 (N_2194,In_2747,In_51);
nand U2195 (N_2195,In_1714,In_1580);
nand U2196 (N_2196,In_1659,In_1924);
and U2197 (N_2197,In_1485,In_2174);
nand U2198 (N_2198,In_1681,In_230);
or U2199 (N_2199,In_1801,In_872);
xnor U2200 (N_2200,In_2102,In_540);
or U2201 (N_2201,In_644,In_1978);
and U2202 (N_2202,In_1812,In_2351);
xor U2203 (N_2203,In_1591,In_1317);
and U2204 (N_2204,In_482,In_2606);
nor U2205 (N_2205,In_2858,In_138);
or U2206 (N_2206,In_498,In_1387);
and U2207 (N_2207,In_1409,In_1323);
nand U2208 (N_2208,In_2678,In_1368);
nand U2209 (N_2209,In_690,In_2999);
and U2210 (N_2210,In_214,In_814);
and U2211 (N_2211,In_231,In_2328);
and U2212 (N_2212,In_1862,In_2356);
xor U2213 (N_2213,In_1069,In_2243);
nand U2214 (N_2214,In_464,In_1421);
or U2215 (N_2215,In_1331,In_389);
and U2216 (N_2216,In_2638,In_1075);
or U2217 (N_2217,In_1616,In_1819);
nand U2218 (N_2218,In_2949,In_1589);
or U2219 (N_2219,In_1653,In_2154);
or U2220 (N_2220,In_1452,In_2503);
nor U2221 (N_2221,In_1021,In_1224);
xnor U2222 (N_2222,In_1003,In_199);
xnor U2223 (N_2223,In_71,In_2652);
nor U2224 (N_2224,In_2842,In_1284);
and U2225 (N_2225,In_1666,In_2511);
nor U2226 (N_2226,In_1837,In_2290);
nand U2227 (N_2227,In_2979,In_329);
or U2228 (N_2228,In_2458,In_235);
and U2229 (N_2229,In_2438,In_989);
or U2230 (N_2230,In_1780,In_953);
nand U2231 (N_2231,In_2719,In_765);
nand U2232 (N_2232,In_822,In_2521);
nor U2233 (N_2233,In_1780,In_87);
xor U2234 (N_2234,In_2432,In_782);
nand U2235 (N_2235,In_1479,In_2255);
or U2236 (N_2236,In_1555,In_2521);
xor U2237 (N_2237,In_1664,In_2852);
nor U2238 (N_2238,In_664,In_839);
or U2239 (N_2239,In_1983,In_806);
nand U2240 (N_2240,In_1738,In_1586);
or U2241 (N_2241,In_379,In_2555);
or U2242 (N_2242,In_1710,In_2815);
xnor U2243 (N_2243,In_993,In_152);
nand U2244 (N_2244,In_609,In_1759);
nor U2245 (N_2245,In_876,In_1119);
xor U2246 (N_2246,In_643,In_2088);
or U2247 (N_2247,In_67,In_2877);
and U2248 (N_2248,In_605,In_2944);
or U2249 (N_2249,In_2687,In_730);
nand U2250 (N_2250,In_1212,In_2035);
nor U2251 (N_2251,In_2540,In_661);
nand U2252 (N_2252,In_1206,In_2309);
nor U2253 (N_2253,In_2018,In_718);
xor U2254 (N_2254,In_1728,In_2946);
nand U2255 (N_2255,In_1599,In_324);
and U2256 (N_2256,In_1877,In_1779);
and U2257 (N_2257,In_1434,In_685);
xnor U2258 (N_2258,In_1020,In_193);
xor U2259 (N_2259,In_1946,In_2065);
xnor U2260 (N_2260,In_1287,In_463);
and U2261 (N_2261,In_1791,In_1034);
xor U2262 (N_2262,In_186,In_1473);
nand U2263 (N_2263,In_2223,In_2286);
nand U2264 (N_2264,In_1685,In_314);
and U2265 (N_2265,In_2177,In_1578);
nor U2266 (N_2266,In_869,In_2268);
and U2267 (N_2267,In_2710,In_2585);
xor U2268 (N_2268,In_1304,In_1695);
nor U2269 (N_2269,In_2977,In_306);
xor U2270 (N_2270,In_1491,In_1846);
and U2271 (N_2271,In_2112,In_2968);
xnor U2272 (N_2272,In_1268,In_2878);
and U2273 (N_2273,In_1,In_2485);
and U2274 (N_2274,In_2793,In_1556);
and U2275 (N_2275,In_1287,In_2488);
nor U2276 (N_2276,In_2553,In_443);
and U2277 (N_2277,In_2034,In_546);
and U2278 (N_2278,In_1204,In_2898);
xor U2279 (N_2279,In_721,In_1438);
nor U2280 (N_2280,In_1645,In_1278);
and U2281 (N_2281,In_372,In_192);
nor U2282 (N_2282,In_197,In_413);
or U2283 (N_2283,In_2262,In_187);
nand U2284 (N_2284,In_1020,In_2306);
or U2285 (N_2285,In_2965,In_2166);
xnor U2286 (N_2286,In_511,In_1676);
or U2287 (N_2287,In_2553,In_2996);
or U2288 (N_2288,In_188,In_2151);
nor U2289 (N_2289,In_2641,In_657);
nor U2290 (N_2290,In_1078,In_2379);
and U2291 (N_2291,In_831,In_2573);
or U2292 (N_2292,In_2854,In_34);
xor U2293 (N_2293,In_1065,In_804);
and U2294 (N_2294,In_1136,In_2938);
xor U2295 (N_2295,In_1686,In_1527);
and U2296 (N_2296,In_1529,In_2191);
xor U2297 (N_2297,In_1474,In_2683);
and U2298 (N_2298,In_2112,In_2150);
nor U2299 (N_2299,In_1959,In_2688);
xnor U2300 (N_2300,In_533,In_1164);
or U2301 (N_2301,In_335,In_3);
and U2302 (N_2302,In_2719,In_518);
or U2303 (N_2303,In_1860,In_2205);
or U2304 (N_2304,In_2101,In_1677);
and U2305 (N_2305,In_1662,In_955);
nand U2306 (N_2306,In_1512,In_2094);
xor U2307 (N_2307,In_178,In_1647);
xnor U2308 (N_2308,In_946,In_53);
nor U2309 (N_2309,In_2258,In_1283);
nand U2310 (N_2310,In_1337,In_2128);
or U2311 (N_2311,In_2289,In_451);
nor U2312 (N_2312,In_1634,In_1959);
and U2313 (N_2313,In_511,In_1909);
or U2314 (N_2314,In_2608,In_2571);
xnor U2315 (N_2315,In_344,In_2010);
nor U2316 (N_2316,In_1357,In_544);
or U2317 (N_2317,In_2738,In_1211);
xnor U2318 (N_2318,In_469,In_2311);
and U2319 (N_2319,In_2114,In_2758);
and U2320 (N_2320,In_2763,In_2445);
nor U2321 (N_2321,In_1381,In_1628);
nor U2322 (N_2322,In_2112,In_1681);
and U2323 (N_2323,In_1705,In_112);
nand U2324 (N_2324,In_1855,In_1189);
xnor U2325 (N_2325,In_2008,In_327);
xnor U2326 (N_2326,In_442,In_601);
nor U2327 (N_2327,In_2709,In_1561);
xnor U2328 (N_2328,In_533,In_644);
xnor U2329 (N_2329,In_2715,In_1780);
nor U2330 (N_2330,In_1931,In_1384);
nor U2331 (N_2331,In_1050,In_532);
nand U2332 (N_2332,In_681,In_2803);
nor U2333 (N_2333,In_426,In_1040);
xnor U2334 (N_2334,In_2498,In_653);
nand U2335 (N_2335,In_307,In_1256);
and U2336 (N_2336,In_1477,In_238);
nor U2337 (N_2337,In_2501,In_2295);
nand U2338 (N_2338,In_1492,In_255);
or U2339 (N_2339,In_309,In_2845);
xor U2340 (N_2340,In_1089,In_2677);
and U2341 (N_2341,In_2546,In_2686);
nor U2342 (N_2342,In_500,In_492);
xnor U2343 (N_2343,In_2384,In_2324);
nor U2344 (N_2344,In_429,In_1313);
nand U2345 (N_2345,In_1283,In_2187);
nand U2346 (N_2346,In_1587,In_2695);
xor U2347 (N_2347,In_287,In_2629);
and U2348 (N_2348,In_525,In_2849);
nand U2349 (N_2349,In_1578,In_1360);
and U2350 (N_2350,In_2214,In_1029);
xor U2351 (N_2351,In_1185,In_224);
nor U2352 (N_2352,In_888,In_74);
and U2353 (N_2353,In_188,In_1372);
nand U2354 (N_2354,In_842,In_61);
or U2355 (N_2355,In_2390,In_2779);
and U2356 (N_2356,In_2332,In_2064);
nand U2357 (N_2357,In_1754,In_1555);
and U2358 (N_2358,In_2729,In_485);
nand U2359 (N_2359,In_507,In_2546);
and U2360 (N_2360,In_2642,In_1844);
and U2361 (N_2361,In_1046,In_2215);
or U2362 (N_2362,In_850,In_1039);
xor U2363 (N_2363,In_753,In_2009);
and U2364 (N_2364,In_2925,In_2542);
nor U2365 (N_2365,In_1865,In_2662);
nand U2366 (N_2366,In_2764,In_2495);
xnor U2367 (N_2367,In_35,In_897);
nor U2368 (N_2368,In_2254,In_2555);
or U2369 (N_2369,In_683,In_1486);
and U2370 (N_2370,In_398,In_2094);
nor U2371 (N_2371,In_2185,In_2379);
nor U2372 (N_2372,In_2670,In_1785);
and U2373 (N_2373,In_2859,In_1438);
xnor U2374 (N_2374,In_1421,In_1785);
nand U2375 (N_2375,In_2431,In_1299);
or U2376 (N_2376,In_1772,In_372);
nand U2377 (N_2377,In_1208,In_2041);
nand U2378 (N_2378,In_2049,In_719);
or U2379 (N_2379,In_538,In_1804);
and U2380 (N_2380,In_221,In_715);
nor U2381 (N_2381,In_1333,In_1151);
and U2382 (N_2382,In_1959,In_118);
and U2383 (N_2383,In_1159,In_544);
nand U2384 (N_2384,In_515,In_1923);
or U2385 (N_2385,In_1505,In_1691);
xor U2386 (N_2386,In_424,In_1839);
and U2387 (N_2387,In_97,In_2721);
nor U2388 (N_2388,In_2944,In_1190);
nor U2389 (N_2389,In_917,In_466);
and U2390 (N_2390,In_1712,In_2216);
nand U2391 (N_2391,In_1286,In_1048);
or U2392 (N_2392,In_1222,In_2647);
and U2393 (N_2393,In_2568,In_1026);
xor U2394 (N_2394,In_2050,In_1725);
or U2395 (N_2395,In_2246,In_1871);
xor U2396 (N_2396,In_2880,In_802);
nor U2397 (N_2397,In_2140,In_1891);
xnor U2398 (N_2398,In_406,In_492);
nand U2399 (N_2399,In_152,In_40);
xor U2400 (N_2400,In_2236,In_1946);
nand U2401 (N_2401,In_358,In_1229);
or U2402 (N_2402,In_2819,In_1299);
nand U2403 (N_2403,In_2650,In_2042);
or U2404 (N_2404,In_48,In_836);
and U2405 (N_2405,In_2460,In_610);
or U2406 (N_2406,In_2785,In_2744);
nand U2407 (N_2407,In_1159,In_2701);
nand U2408 (N_2408,In_1290,In_1046);
or U2409 (N_2409,In_1172,In_2160);
nand U2410 (N_2410,In_1645,In_1117);
or U2411 (N_2411,In_2102,In_217);
nor U2412 (N_2412,In_474,In_1814);
and U2413 (N_2413,In_2104,In_2793);
and U2414 (N_2414,In_1967,In_1436);
or U2415 (N_2415,In_366,In_2990);
or U2416 (N_2416,In_1362,In_2801);
xor U2417 (N_2417,In_44,In_1717);
nand U2418 (N_2418,In_697,In_2915);
or U2419 (N_2419,In_762,In_1009);
and U2420 (N_2420,In_1400,In_248);
and U2421 (N_2421,In_2063,In_921);
xnor U2422 (N_2422,In_407,In_2675);
or U2423 (N_2423,In_789,In_1690);
nor U2424 (N_2424,In_565,In_478);
xnor U2425 (N_2425,In_724,In_1185);
nand U2426 (N_2426,In_1926,In_2056);
xor U2427 (N_2427,In_404,In_967);
or U2428 (N_2428,In_2967,In_1132);
xnor U2429 (N_2429,In_2087,In_1796);
and U2430 (N_2430,In_1746,In_1731);
xor U2431 (N_2431,In_2259,In_2410);
or U2432 (N_2432,In_2790,In_320);
nand U2433 (N_2433,In_1369,In_2220);
nor U2434 (N_2434,In_1311,In_2157);
nor U2435 (N_2435,In_1458,In_840);
nand U2436 (N_2436,In_260,In_1982);
and U2437 (N_2437,In_367,In_2951);
or U2438 (N_2438,In_2574,In_1917);
nor U2439 (N_2439,In_973,In_1291);
nand U2440 (N_2440,In_2441,In_1261);
nand U2441 (N_2441,In_1952,In_710);
or U2442 (N_2442,In_1155,In_2724);
xor U2443 (N_2443,In_1907,In_2661);
and U2444 (N_2444,In_1003,In_1131);
and U2445 (N_2445,In_360,In_335);
nor U2446 (N_2446,In_2382,In_2567);
nand U2447 (N_2447,In_1974,In_584);
or U2448 (N_2448,In_2107,In_2793);
nor U2449 (N_2449,In_1376,In_830);
and U2450 (N_2450,In_644,In_2193);
nor U2451 (N_2451,In_1880,In_1171);
xnor U2452 (N_2452,In_1350,In_1372);
and U2453 (N_2453,In_1631,In_2429);
xor U2454 (N_2454,In_2614,In_1870);
nor U2455 (N_2455,In_13,In_233);
or U2456 (N_2456,In_2559,In_2783);
xnor U2457 (N_2457,In_113,In_1348);
or U2458 (N_2458,In_1118,In_2363);
or U2459 (N_2459,In_972,In_2584);
and U2460 (N_2460,In_2570,In_2143);
nand U2461 (N_2461,In_879,In_1364);
xnor U2462 (N_2462,In_381,In_1332);
xor U2463 (N_2463,In_1087,In_1138);
or U2464 (N_2464,In_352,In_462);
nor U2465 (N_2465,In_1772,In_772);
or U2466 (N_2466,In_2805,In_1133);
nand U2467 (N_2467,In_628,In_1618);
nor U2468 (N_2468,In_1026,In_913);
nand U2469 (N_2469,In_1402,In_767);
nand U2470 (N_2470,In_1407,In_2566);
xor U2471 (N_2471,In_172,In_1496);
xor U2472 (N_2472,In_2682,In_317);
xor U2473 (N_2473,In_1844,In_2438);
nand U2474 (N_2474,In_1236,In_561);
and U2475 (N_2475,In_69,In_2315);
xor U2476 (N_2476,In_1656,In_391);
or U2477 (N_2477,In_729,In_961);
and U2478 (N_2478,In_637,In_684);
or U2479 (N_2479,In_2727,In_1681);
or U2480 (N_2480,In_1672,In_1349);
or U2481 (N_2481,In_2726,In_2653);
or U2482 (N_2482,In_1219,In_1400);
and U2483 (N_2483,In_555,In_1883);
and U2484 (N_2484,In_1300,In_1975);
nor U2485 (N_2485,In_197,In_2933);
nand U2486 (N_2486,In_515,In_2625);
nor U2487 (N_2487,In_881,In_1295);
or U2488 (N_2488,In_676,In_1497);
nand U2489 (N_2489,In_1388,In_2713);
and U2490 (N_2490,In_805,In_1095);
xor U2491 (N_2491,In_2240,In_1825);
xor U2492 (N_2492,In_1890,In_333);
xnor U2493 (N_2493,In_2023,In_1652);
xnor U2494 (N_2494,In_1561,In_1031);
or U2495 (N_2495,In_1727,In_517);
or U2496 (N_2496,In_1224,In_2131);
nand U2497 (N_2497,In_1533,In_2007);
nand U2498 (N_2498,In_1632,In_2933);
xnor U2499 (N_2499,In_2579,In_2226);
nor U2500 (N_2500,In_741,In_1784);
xnor U2501 (N_2501,In_995,In_2733);
nand U2502 (N_2502,In_2924,In_1241);
and U2503 (N_2503,In_2328,In_270);
and U2504 (N_2504,In_1362,In_1198);
and U2505 (N_2505,In_503,In_992);
or U2506 (N_2506,In_614,In_45);
or U2507 (N_2507,In_2615,In_438);
nor U2508 (N_2508,In_1598,In_1463);
nor U2509 (N_2509,In_1339,In_1087);
nor U2510 (N_2510,In_276,In_518);
nand U2511 (N_2511,In_1183,In_1769);
nor U2512 (N_2512,In_1515,In_507);
nand U2513 (N_2513,In_1609,In_110);
nor U2514 (N_2514,In_2146,In_2969);
nor U2515 (N_2515,In_2846,In_2919);
xor U2516 (N_2516,In_1727,In_1308);
xnor U2517 (N_2517,In_2518,In_2687);
xnor U2518 (N_2518,In_1079,In_2943);
and U2519 (N_2519,In_23,In_505);
and U2520 (N_2520,In_845,In_799);
nor U2521 (N_2521,In_2949,In_1323);
or U2522 (N_2522,In_677,In_2113);
nor U2523 (N_2523,In_1224,In_2546);
nor U2524 (N_2524,In_347,In_172);
nor U2525 (N_2525,In_1604,In_2457);
xor U2526 (N_2526,In_1107,In_2541);
and U2527 (N_2527,In_446,In_1739);
xor U2528 (N_2528,In_1622,In_462);
or U2529 (N_2529,In_358,In_656);
or U2530 (N_2530,In_2536,In_2903);
xor U2531 (N_2531,In_2758,In_1364);
xnor U2532 (N_2532,In_2910,In_1703);
or U2533 (N_2533,In_2570,In_284);
or U2534 (N_2534,In_807,In_208);
or U2535 (N_2535,In_1048,In_1141);
xnor U2536 (N_2536,In_2858,In_1101);
or U2537 (N_2537,In_272,In_2098);
or U2538 (N_2538,In_537,In_2798);
nor U2539 (N_2539,In_1035,In_364);
nor U2540 (N_2540,In_852,In_1820);
xnor U2541 (N_2541,In_763,In_1986);
xnor U2542 (N_2542,In_1495,In_1885);
nor U2543 (N_2543,In_2739,In_191);
nand U2544 (N_2544,In_1909,In_899);
nand U2545 (N_2545,In_909,In_2258);
nand U2546 (N_2546,In_2635,In_2989);
or U2547 (N_2547,In_2941,In_2709);
nor U2548 (N_2548,In_2352,In_2576);
xnor U2549 (N_2549,In_2360,In_2026);
or U2550 (N_2550,In_1651,In_1594);
nand U2551 (N_2551,In_2819,In_1605);
nor U2552 (N_2552,In_2773,In_2135);
and U2553 (N_2553,In_1272,In_2769);
nor U2554 (N_2554,In_1630,In_1193);
nor U2555 (N_2555,In_1839,In_413);
xor U2556 (N_2556,In_1056,In_2654);
or U2557 (N_2557,In_295,In_2035);
nor U2558 (N_2558,In_1265,In_1338);
nor U2559 (N_2559,In_75,In_2738);
nand U2560 (N_2560,In_1897,In_2203);
and U2561 (N_2561,In_172,In_1730);
nand U2562 (N_2562,In_2605,In_2362);
or U2563 (N_2563,In_2143,In_325);
nor U2564 (N_2564,In_1373,In_2891);
nand U2565 (N_2565,In_352,In_841);
and U2566 (N_2566,In_1230,In_991);
nand U2567 (N_2567,In_2341,In_850);
or U2568 (N_2568,In_1431,In_54);
or U2569 (N_2569,In_1642,In_1404);
or U2570 (N_2570,In_2190,In_207);
and U2571 (N_2571,In_1197,In_1854);
and U2572 (N_2572,In_2881,In_2568);
and U2573 (N_2573,In_2637,In_452);
or U2574 (N_2574,In_828,In_124);
and U2575 (N_2575,In_1790,In_1594);
and U2576 (N_2576,In_1619,In_2009);
nand U2577 (N_2577,In_2769,In_2099);
nand U2578 (N_2578,In_500,In_2451);
and U2579 (N_2579,In_1842,In_2132);
nand U2580 (N_2580,In_1541,In_687);
nand U2581 (N_2581,In_2941,In_2438);
nor U2582 (N_2582,In_2148,In_2991);
and U2583 (N_2583,In_2338,In_8);
or U2584 (N_2584,In_1736,In_2371);
nand U2585 (N_2585,In_717,In_1376);
nand U2586 (N_2586,In_2749,In_1315);
nor U2587 (N_2587,In_1412,In_870);
nor U2588 (N_2588,In_446,In_1654);
xnor U2589 (N_2589,In_1655,In_2122);
or U2590 (N_2590,In_2838,In_811);
nor U2591 (N_2591,In_1172,In_2279);
and U2592 (N_2592,In_2185,In_485);
nand U2593 (N_2593,In_2405,In_479);
or U2594 (N_2594,In_2406,In_5);
xnor U2595 (N_2595,In_2599,In_1279);
and U2596 (N_2596,In_623,In_390);
nand U2597 (N_2597,In_2457,In_2574);
or U2598 (N_2598,In_1362,In_2530);
or U2599 (N_2599,In_768,In_703);
nor U2600 (N_2600,In_2032,In_2835);
xnor U2601 (N_2601,In_1538,In_1567);
nand U2602 (N_2602,In_286,In_784);
or U2603 (N_2603,In_2999,In_2434);
nand U2604 (N_2604,In_2330,In_2659);
nand U2605 (N_2605,In_1954,In_212);
or U2606 (N_2606,In_2166,In_990);
nand U2607 (N_2607,In_358,In_1282);
or U2608 (N_2608,In_474,In_2992);
or U2609 (N_2609,In_2676,In_778);
or U2610 (N_2610,In_827,In_2599);
or U2611 (N_2611,In_8,In_1894);
nand U2612 (N_2612,In_2551,In_112);
nor U2613 (N_2613,In_186,In_1894);
or U2614 (N_2614,In_2036,In_2315);
and U2615 (N_2615,In_1964,In_1283);
and U2616 (N_2616,In_35,In_2045);
and U2617 (N_2617,In_1650,In_1689);
xor U2618 (N_2618,In_1292,In_2174);
nand U2619 (N_2619,In_1429,In_2953);
and U2620 (N_2620,In_781,In_435);
and U2621 (N_2621,In_2091,In_304);
nand U2622 (N_2622,In_1135,In_450);
or U2623 (N_2623,In_679,In_667);
xnor U2624 (N_2624,In_1809,In_16);
or U2625 (N_2625,In_1783,In_257);
xor U2626 (N_2626,In_2403,In_2561);
or U2627 (N_2627,In_1933,In_2609);
xor U2628 (N_2628,In_374,In_85);
xor U2629 (N_2629,In_72,In_2318);
nor U2630 (N_2630,In_868,In_1677);
nor U2631 (N_2631,In_2868,In_2127);
xor U2632 (N_2632,In_1701,In_1116);
nor U2633 (N_2633,In_474,In_2139);
xor U2634 (N_2634,In_1791,In_2228);
or U2635 (N_2635,In_1557,In_1721);
nand U2636 (N_2636,In_95,In_795);
and U2637 (N_2637,In_1674,In_97);
and U2638 (N_2638,In_1752,In_1665);
or U2639 (N_2639,In_2535,In_1125);
or U2640 (N_2640,In_237,In_309);
xnor U2641 (N_2641,In_2289,In_2623);
xnor U2642 (N_2642,In_1221,In_1934);
nand U2643 (N_2643,In_1538,In_2420);
nand U2644 (N_2644,In_985,In_53);
xor U2645 (N_2645,In_330,In_2479);
nand U2646 (N_2646,In_2054,In_1780);
xnor U2647 (N_2647,In_1140,In_207);
and U2648 (N_2648,In_1138,In_1931);
or U2649 (N_2649,In_1193,In_1501);
and U2650 (N_2650,In_372,In_1827);
xor U2651 (N_2651,In_1105,In_2818);
or U2652 (N_2652,In_1287,In_1019);
nand U2653 (N_2653,In_2464,In_200);
or U2654 (N_2654,In_1941,In_69);
and U2655 (N_2655,In_1169,In_1969);
nor U2656 (N_2656,In_1662,In_63);
and U2657 (N_2657,In_1600,In_2947);
or U2658 (N_2658,In_521,In_1607);
nand U2659 (N_2659,In_530,In_1892);
and U2660 (N_2660,In_1564,In_1638);
or U2661 (N_2661,In_2608,In_1242);
or U2662 (N_2662,In_178,In_2374);
and U2663 (N_2663,In_476,In_2452);
xor U2664 (N_2664,In_2685,In_2956);
xnor U2665 (N_2665,In_473,In_232);
and U2666 (N_2666,In_2281,In_1581);
xor U2667 (N_2667,In_458,In_682);
or U2668 (N_2668,In_1617,In_2763);
and U2669 (N_2669,In_77,In_1803);
or U2670 (N_2670,In_111,In_2843);
xor U2671 (N_2671,In_1620,In_455);
or U2672 (N_2672,In_2960,In_1458);
xnor U2673 (N_2673,In_1218,In_864);
nand U2674 (N_2674,In_2814,In_2259);
nor U2675 (N_2675,In_1911,In_2756);
xnor U2676 (N_2676,In_2596,In_1345);
nand U2677 (N_2677,In_2373,In_1051);
and U2678 (N_2678,In_2652,In_1397);
xnor U2679 (N_2679,In_747,In_2808);
xnor U2680 (N_2680,In_135,In_2908);
or U2681 (N_2681,In_2153,In_917);
and U2682 (N_2682,In_166,In_326);
xnor U2683 (N_2683,In_2095,In_1321);
and U2684 (N_2684,In_2473,In_234);
and U2685 (N_2685,In_2818,In_648);
nand U2686 (N_2686,In_747,In_895);
nor U2687 (N_2687,In_2803,In_1210);
xor U2688 (N_2688,In_854,In_758);
and U2689 (N_2689,In_467,In_2390);
xnor U2690 (N_2690,In_1295,In_865);
xnor U2691 (N_2691,In_1763,In_1109);
or U2692 (N_2692,In_1633,In_2284);
or U2693 (N_2693,In_1838,In_538);
nand U2694 (N_2694,In_387,In_893);
xnor U2695 (N_2695,In_1056,In_205);
xor U2696 (N_2696,In_1566,In_1549);
or U2697 (N_2697,In_719,In_1283);
nor U2698 (N_2698,In_1984,In_1622);
and U2699 (N_2699,In_2122,In_1760);
or U2700 (N_2700,In_477,In_841);
xnor U2701 (N_2701,In_175,In_400);
and U2702 (N_2702,In_719,In_1174);
and U2703 (N_2703,In_27,In_1292);
or U2704 (N_2704,In_2008,In_479);
nor U2705 (N_2705,In_596,In_1422);
nor U2706 (N_2706,In_2779,In_575);
nand U2707 (N_2707,In_2867,In_1075);
and U2708 (N_2708,In_1407,In_1952);
xnor U2709 (N_2709,In_1108,In_972);
and U2710 (N_2710,In_2500,In_1535);
nand U2711 (N_2711,In_2162,In_52);
xor U2712 (N_2712,In_2777,In_2672);
and U2713 (N_2713,In_1202,In_1177);
nor U2714 (N_2714,In_2311,In_2476);
or U2715 (N_2715,In_1194,In_2666);
nor U2716 (N_2716,In_2109,In_2516);
xnor U2717 (N_2717,In_1421,In_321);
nand U2718 (N_2718,In_2732,In_2224);
or U2719 (N_2719,In_439,In_972);
and U2720 (N_2720,In_2979,In_2232);
nand U2721 (N_2721,In_366,In_2067);
xor U2722 (N_2722,In_2254,In_1028);
and U2723 (N_2723,In_1490,In_1234);
xor U2724 (N_2724,In_2599,In_93);
or U2725 (N_2725,In_2581,In_268);
and U2726 (N_2726,In_704,In_2618);
nand U2727 (N_2727,In_63,In_2896);
nand U2728 (N_2728,In_1305,In_2243);
xor U2729 (N_2729,In_319,In_2099);
or U2730 (N_2730,In_1589,In_2979);
nor U2731 (N_2731,In_1450,In_450);
and U2732 (N_2732,In_1932,In_630);
xor U2733 (N_2733,In_58,In_1456);
nand U2734 (N_2734,In_2142,In_817);
nor U2735 (N_2735,In_1240,In_41);
nor U2736 (N_2736,In_1213,In_1020);
and U2737 (N_2737,In_1254,In_603);
or U2738 (N_2738,In_1726,In_2464);
xor U2739 (N_2739,In_839,In_1650);
xor U2740 (N_2740,In_1453,In_1268);
xnor U2741 (N_2741,In_2590,In_1234);
xnor U2742 (N_2742,In_1011,In_2662);
nand U2743 (N_2743,In_1335,In_1393);
and U2744 (N_2744,In_1664,In_2105);
xor U2745 (N_2745,In_545,In_895);
nor U2746 (N_2746,In_1414,In_2800);
and U2747 (N_2747,In_2117,In_1381);
or U2748 (N_2748,In_1886,In_1473);
nor U2749 (N_2749,In_545,In_548);
nor U2750 (N_2750,In_82,In_261);
xnor U2751 (N_2751,In_2101,In_1032);
nor U2752 (N_2752,In_2960,In_865);
nand U2753 (N_2753,In_446,In_2561);
and U2754 (N_2754,In_1644,In_537);
nand U2755 (N_2755,In_2709,In_1972);
nand U2756 (N_2756,In_935,In_224);
and U2757 (N_2757,In_517,In_1775);
nor U2758 (N_2758,In_1849,In_1596);
xnor U2759 (N_2759,In_1448,In_330);
xor U2760 (N_2760,In_76,In_997);
xnor U2761 (N_2761,In_2654,In_353);
nor U2762 (N_2762,In_2172,In_1154);
and U2763 (N_2763,In_696,In_1135);
or U2764 (N_2764,In_1695,In_2760);
xor U2765 (N_2765,In_1042,In_471);
nand U2766 (N_2766,In_405,In_126);
and U2767 (N_2767,In_99,In_2027);
nor U2768 (N_2768,In_1705,In_192);
and U2769 (N_2769,In_2967,In_1908);
xor U2770 (N_2770,In_318,In_1875);
nand U2771 (N_2771,In_139,In_1751);
nand U2772 (N_2772,In_1254,In_2757);
and U2773 (N_2773,In_1802,In_532);
nand U2774 (N_2774,In_590,In_2509);
and U2775 (N_2775,In_22,In_1525);
and U2776 (N_2776,In_2031,In_2365);
nand U2777 (N_2777,In_135,In_935);
or U2778 (N_2778,In_2654,In_2982);
xor U2779 (N_2779,In_1847,In_2043);
and U2780 (N_2780,In_1957,In_548);
nand U2781 (N_2781,In_687,In_2937);
and U2782 (N_2782,In_1054,In_2103);
or U2783 (N_2783,In_2069,In_475);
nor U2784 (N_2784,In_1742,In_359);
or U2785 (N_2785,In_1275,In_1728);
or U2786 (N_2786,In_1171,In_401);
nor U2787 (N_2787,In_438,In_1744);
xnor U2788 (N_2788,In_799,In_2769);
nand U2789 (N_2789,In_491,In_1354);
xor U2790 (N_2790,In_2853,In_1797);
xor U2791 (N_2791,In_2003,In_1286);
or U2792 (N_2792,In_2426,In_1177);
nor U2793 (N_2793,In_2483,In_2650);
xor U2794 (N_2794,In_1600,In_733);
or U2795 (N_2795,In_2720,In_2881);
nand U2796 (N_2796,In_2565,In_1431);
or U2797 (N_2797,In_301,In_589);
or U2798 (N_2798,In_312,In_2208);
and U2799 (N_2799,In_629,In_511);
nand U2800 (N_2800,In_2887,In_1191);
nor U2801 (N_2801,In_1719,In_1731);
nand U2802 (N_2802,In_927,In_2488);
nor U2803 (N_2803,In_692,In_1);
or U2804 (N_2804,In_1294,In_1520);
or U2805 (N_2805,In_734,In_831);
nand U2806 (N_2806,In_837,In_2748);
or U2807 (N_2807,In_1886,In_1257);
and U2808 (N_2808,In_564,In_32);
or U2809 (N_2809,In_2989,In_234);
or U2810 (N_2810,In_1023,In_418);
and U2811 (N_2811,In_2347,In_1103);
xnor U2812 (N_2812,In_589,In_1560);
xnor U2813 (N_2813,In_2064,In_2121);
xor U2814 (N_2814,In_2464,In_1925);
nand U2815 (N_2815,In_2264,In_2598);
or U2816 (N_2816,In_83,In_348);
nor U2817 (N_2817,In_2445,In_829);
nor U2818 (N_2818,In_459,In_2071);
nand U2819 (N_2819,In_279,In_519);
nor U2820 (N_2820,In_340,In_571);
xor U2821 (N_2821,In_592,In_2141);
nand U2822 (N_2822,In_1433,In_2905);
nor U2823 (N_2823,In_1424,In_92);
xnor U2824 (N_2824,In_1371,In_2016);
and U2825 (N_2825,In_831,In_181);
nand U2826 (N_2826,In_694,In_420);
and U2827 (N_2827,In_1376,In_410);
or U2828 (N_2828,In_412,In_969);
or U2829 (N_2829,In_1595,In_2824);
and U2830 (N_2830,In_871,In_112);
xnor U2831 (N_2831,In_2047,In_1807);
xnor U2832 (N_2832,In_72,In_515);
nor U2833 (N_2833,In_120,In_97);
or U2834 (N_2834,In_2309,In_984);
and U2835 (N_2835,In_2249,In_1425);
and U2836 (N_2836,In_2752,In_2947);
xor U2837 (N_2837,In_2896,In_359);
nor U2838 (N_2838,In_2658,In_2704);
nor U2839 (N_2839,In_624,In_1290);
nand U2840 (N_2840,In_1249,In_68);
nor U2841 (N_2841,In_2778,In_2810);
and U2842 (N_2842,In_1720,In_1916);
xnor U2843 (N_2843,In_1072,In_2011);
xor U2844 (N_2844,In_159,In_616);
or U2845 (N_2845,In_2335,In_2264);
or U2846 (N_2846,In_808,In_1671);
nor U2847 (N_2847,In_293,In_2781);
nor U2848 (N_2848,In_1785,In_2539);
and U2849 (N_2849,In_2917,In_2476);
or U2850 (N_2850,In_647,In_1288);
or U2851 (N_2851,In_2013,In_963);
nor U2852 (N_2852,In_1880,In_1764);
nand U2853 (N_2853,In_2826,In_216);
nand U2854 (N_2854,In_540,In_2769);
or U2855 (N_2855,In_1381,In_2857);
nor U2856 (N_2856,In_2119,In_2299);
nor U2857 (N_2857,In_354,In_487);
xor U2858 (N_2858,In_2232,In_2827);
nand U2859 (N_2859,In_2117,In_1767);
or U2860 (N_2860,In_1684,In_1300);
nor U2861 (N_2861,In_1063,In_2587);
xor U2862 (N_2862,In_2367,In_303);
or U2863 (N_2863,In_309,In_827);
nor U2864 (N_2864,In_1492,In_139);
or U2865 (N_2865,In_562,In_105);
nand U2866 (N_2866,In_523,In_712);
or U2867 (N_2867,In_35,In_2419);
nor U2868 (N_2868,In_2447,In_1119);
or U2869 (N_2869,In_1459,In_2081);
nand U2870 (N_2870,In_137,In_2642);
nor U2871 (N_2871,In_1283,In_2329);
xnor U2872 (N_2872,In_829,In_2468);
or U2873 (N_2873,In_1983,In_1697);
nand U2874 (N_2874,In_2522,In_2501);
nand U2875 (N_2875,In_1825,In_2727);
and U2876 (N_2876,In_258,In_999);
xor U2877 (N_2877,In_2539,In_216);
or U2878 (N_2878,In_599,In_1877);
xnor U2879 (N_2879,In_1037,In_1726);
and U2880 (N_2880,In_960,In_1946);
xor U2881 (N_2881,In_2091,In_463);
or U2882 (N_2882,In_554,In_349);
and U2883 (N_2883,In_1349,In_2764);
xnor U2884 (N_2884,In_1393,In_1668);
nand U2885 (N_2885,In_50,In_2244);
xor U2886 (N_2886,In_562,In_47);
or U2887 (N_2887,In_179,In_623);
or U2888 (N_2888,In_2604,In_232);
or U2889 (N_2889,In_558,In_1291);
or U2890 (N_2890,In_518,In_1970);
or U2891 (N_2891,In_1666,In_2304);
nor U2892 (N_2892,In_2836,In_2734);
and U2893 (N_2893,In_1234,In_892);
and U2894 (N_2894,In_1243,In_1746);
xnor U2895 (N_2895,In_888,In_1966);
xnor U2896 (N_2896,In_2478,In_726);
nor U2897 (N_2897,In_91,In_2641);
nor U2898 (N_2898,In_1502,In_1390);
xor U2899 (N_2899,In_2886,In_951);
or U2900 (N_2900,In_2802,In_1781);
or U2901 (N_2901,In_837,In_2000);
xnor U2902 (N_2902,In_785,In_283);
nand U2903 (N_2903,In_1342,In_310);
nand U2904 (N_2904,In_1384,In_1446);
or U2905 (N_2905,In_513,In_1354);
xor U2906 (N_2906,In_2938,In_1188);
nand U2907 (N_2907,In_2865,In_522);
and U2908 (N_2908,In_1490,In_2704);
and U2909 (N_2909,In_1170,In_647);
or U2910 (N_2910,In_2345,In_1488);
or U2911 (N_2911,In_2240,In_2933);
nand U2912 (N_2912,In_591,In_1477);
and U2913 (N_2913,In_1413,In_1441);
nand U2914 (N_2914,In_1941,In_1942);
nor U2915 (N_2915,In_1880,In_2751);
xnor U2916 (N_2916,In_1596,In_264);
xor U2917 (N_2917,In_1641,In_966);
nand U2918 (N_2918,In_701,In_2142);
xnor U2919 (N_2919,In_259,In_2487);
and U2920 (N_2920,In_1039,In_292);
and U2921 (N_2921,In_1672,In_375);
and U2922 (N_2922,In_2335,In_107);
nor U2923 (N_2923,In_2161,In_639);
xor U2924 (N_2924,In_1809,In_678);
or U2925 (N_2925,In_361,In_2100);
nand U2926 (N_2926,In_2832,In_2889);
and U2927 (N_2927,In_1282,In_2967);
nor U2928 (N_2928,In_2026,In_421);
nor U2929 (N_2929,In_1553,In_195);
nor U2930 (N_2930,In_947,In_2159);
nand U2931 (N_2931,In_2231,In_982);
or U2932 (N_2932,In_1675,In_843);
xnor U2933 (N_2933,In_1533,In_986);
or U2934 (N_2934,In_1164,In_1463);
xor U2935 (N_2935,In_388,In_1846);
or U2936 (N_2936,In_2814,In_2746);
and U2937 (N_2937,In_1064,In_1025);
or U2938 (N_2938,In_1196,In_22);
nand U2939 (N_2939,In_1880,In_909);
nand U2940 (N_2940,In_618,In_2979);
and U2941 (N_2941,In_633,In_1980);
and U2942 (N_2942,In_2418,In_809);
and U2943 (N_2943,In_2818,In_1284);
xnor U2944 (N_2944,In_838,In_617);
nand U2945 (N_2945,In_906,In_1972);
or U2946 (N_2946,In_1853,In_2690);
and U2947 (N_2947,In_1087,In_2871);
xnor U2948 (N_2948,In_2642,In_298);
xnor U2949 (N_2949,In_1359,In_204);
or U2950 (N_2950,In_1391,In_2130);
or U2951 (N_2951,In_2088,In_54);
and U2952 (N_2952,In_1614,In_1340);
xnor U2953 (N_2953,In_773,In_379);
nand U2954 (N_2954,In_2287,In_707);
xor U2955 (N_2955,In_2270,In_1652);
and U2956 (N_2956,In_2606,In_1852);
and U2957 (N_2957,In_298,In_24);
or U2958 (N_2958,In_2212,In_133);
nand U2959 (N_2959,In_819,In_1256);
or U2960 (N_2960,In_656,In_2295);
or U2961 (N_2961,In_213,In_1031);
xnor U2962 (N_2962,In_2486,In_2355);
nor U2963 (N_2963,In_790,In_1104);
and U2964 (N_2964,In_806,In_15);
or U2965 (N_2965,In_2365,In_2285);
nor U2966 (N_2966,In_894,In_1791);
nor U2967 (N_2967,In_2659,In_277);
xnor U2968 (N_2968,In_47,In_749);
and U2969 (N_2969,In_2483,In_2800);
nor U2970 (N_2970,In_524,In_2647);
xor U2971 (N_2971,In_2563,In_2775);
or U2972 (N_2972,In_52,In_2302);
xnor U2973 (N_2973,In_2873,In_1911);
nor U2974 (N_2974,In_1426,In_2677);
and U2975 (N_2975,In_1711,In_2833);
nor U2976 (N_2976,In_2376,In_2077);
xnor U2977 (N_2977,In_1087,In_2930);
nor U2978 (N_2978,In_746,In_1539);
or U2979 (N_2979,In_950,In_1478);
or U2980 (N_2980,In_2086,In_854);
nand U2981 (N_2981,In_1460,In_1222);
nand U2982 (N_2982,In_1782,In_1475);
and U2983 (N_2983,In_677,In_47);
and U2984 (N_2984,In_2494,In_2042);
or U2985 (N_2985,In_2512,In_381);
nand U2986 (N_2986,In_1988,In_2961);
and U2987 (N_2987,In_1525,In_882);
or U2988 (N_2988,In_2641,In_381);
nor U2989 (N_2989,In_2590,In_2179);
or U2990 (N_2990,In_7,In_2892);
and U2991 (N_2991,In_1456,In_634);
and U2992 (N_2992,In_2411,In_34);
xnor U2993 (N_2993,In_473,In_2790);
or U2994 (N_2994,In_1074,In_628);
xnor U2995 (N_2995,In_1036,In_866);
or U2996 (N_2996,In_1007,In_223);
or U2997 (N_2997,In_104,In_889);
nand U2998 (N_2998,In_591,In_1390);
nand U2999 (N_2999,In_681,In_1167);
nor U3000 (N_3000,In_470,In_2601);
and U3001 (N_3001,In_960,In_421);
nor U3002 (N_3002,In_1234,In_2247);
xnor U3003 (N_3003,In_1122,In_1329);
and U3004 (N_3004,In_708,In_744);
xnor U3005 (N_3005,In_1772,In_1565);
nand U3006 (N_3006,In_790,In_1966);
and U3007 (N_3007,In_2231,In_1263);
or U3008 (N_3008,In_1788,In_1634);
and U3009 (N_3009,In_581,In_2536);
and U3010 (N_3010,In_2662,In_2352);
and U3011 (N_3011,In_2837,In_1765);
nand U3012 (N_3012,In_1736,In_2558);
xor U3013 (N_3013,In_543,In_1689);
and U3014 (N_3014,In_471,In_1027);
and U3015 (N_3015,In_2377,In_1480);
and U3016 (N_3016,In_2503,In_923);
or U3017 (N_3017,In_1143,In_2373);
and U3018 (N_3018,In_2523,In_1477);
and U3019 (N_3019,In_140,In_1620);
and U3020 (N_3020,In_2155,In_2049);
and U3021 (N_3021,In_468,In_428);
nand U3022 (N_3022,In_1086,In_2771);
xor U3023 (N_3023,In_2544,In_2003);
nand U3024 (N_3024,In_1928,In_1126);
nand U3025 (N_3025,In_1555,In_2047);
xor U3026 (N_3026,In_914,In_329);
xnor U3027 (N_3027,In_681,In_1693);
nand U3028 (N_3028,In_544,In_1205);
xnor U3029 (N_3029,In_1562,In_83);
xor U3030 (N_3030,In_376,In_2681);
or U3031 (N_3031,In_251,In_2563);
nor U3032 (N_3032,In_908,In_1033);
xor U3033 (N_3033,In_1351,In_2613);
or U3034 (N_3034,In_2760,In_888);
xor U3035 (N_3035,In_2564,In_2447);
xor U3036 (N_3036,In_1898,In_1753);
xor U3037 (N_3037,In_2541,In_1745);
or U3038 (N_3038,In_955,In_450);
and U3039 (N_3039,In_487,In_901);
nor U3040 (N_3040,In_2794,In_498);
nand U3041 (N_3041,In_59,In_2563);
nand U3042 (N_3042,In_1226,In_179);
or U3043 (N_3043,In_888,In_2320);
nor U3044 (N_3044,In_913,In_988);
xor U3045 (N_3045,In_1921,In_205);
xnor U3046 (N_3046,In_179,In_2829);
nor U3047 (N_3047,In_1387,In_371);
and U3048 (N_3048,In_693,In_2606);
nand U3049 (N_3049,In_1295,In_2176);
nand U3050 (N_3050,In_2051,In_667);
or U3051 (N_3051,In_2662,In_760);
and U3052 (N_3052,In_467,In_2178);
or U3053 (N_3053,In_642,In_2581);
or U3054 (N_3054,In_653,In_756);
nor U3055 (N_3055,In_1694,In_2414);
nor U3056 (N_3056,In_396,In_501);
and U3057 (N_3057,In_1011,In_2307);
xor U3058 (N_3058,In_1797,In_485);
or U3059 (N_3059,In_999,In_1802);
nand U3060 (N_3060,In_1739,In_867);
or U3061 (N_3061,In_2468,In_2851);
xnor U3062 (N_3062,In_1749,In_668);
nand U3063 (N_3063,In_1195,In_99);
nand U3064 (N_3064,In_143,In_272);
xnor U3065 (N_3065,In_1772,In_2071);
and U3066 (N_3066,In_1990,In_553);
or U3067 (N_3067,In_1293,In_1268);
or U3068 (N_3068,In_575,In_2203);
xor U3069 (N_3069,In_2705,In_2726);
nor U3070 (N_3070,In_1066,In_1591);
or U3071 (N_3071,In_2987,In_1324);
xor U3072 (N_3072,In_495,In_1674);
or U3073 (N_3073,In_1080,In_1874);
nand U3074 (N_3074,In_1315,In_2291);
xor U3075 (N_3075,In_2116,In_2133);
nor U3076 (N_3076,In_1863,In_2253);
xnor U3077 (N_3077,In_2136,In_1208);
and U3078 (N_3078,In_2698,In_2462);
nand U3079 (N_3079,In_1848,In_1084);
and U3080 (N_3080,In_582,In_2962);
nor U3081 (N_3081,In_1396,In_2474);
or U3082 (N_3082,In_2700,In_626);
xor U3083 (N_3083,In_1495,In_1841);
xnor U3084 (N_3084,In_1910,In_2991);
nand U3085 (N_3085,In_218,In_1274);
or U3086 (N_3086,In_541,In_1627);
and U3087 (N_3087,In_289,In_963);
xor U3088 (N_3088,In_2141,In_1572);
nand U3089 (N_3089,In_2386,In_2020);
nor U3090 (N_3090,In_1119,In_1548);
nor U3091 (N_3091,In_1189,In_2943);
nor U3092 (N_3092,In_1587,In_684);
nor U3093 (N_3093,In_876,In_2204);
nor U3094 (N_3094,In_1287,In_886);
nand U3095 (N_3095,In_2459,In_1328);
nand U3096 (N_3096,In_447,In_649);
and U3097 (N_3097,In_2054,In_2124);
xor U3098 (N_3098,In_673,In_1236);
nand U3099 (N_3099,In_902,In_1079);
nor U3100 (N_3100,In_1955,In_1730);
or U3101 (N_3101,In_426,In_1599);
xor U3102 (N_3102,In_1636,In_2599);
xor U3103 (N_3103,In_1707,In_2581);
and U3104 (N_3104,In_922,In_809);
nor U3105 (N_3105,In_2001,In_2583);
nor U3106 (N_3106,In_1145,In_633);
nand U3107 (N_3107,In_92,In_882);
nand U3108 (N_3108,In_885,In_777);
nand U3109 (N_3109,In_363,In_1367);
or U3110 (N_3110,In_651,In_2395);
or U3111 (N_3111,In_2583,In_2849);
xor U3112 (N_3112,In_785,In_2214);
nand U3113 (N_3113,In_1740,In_455);
and U3114 (N_3114,In_102,In_621);
nor U3115 (N_3115,In_2217,In_1064);
nand U3116 (N_3116,In_2788,In_1471);
and U3117 (N_3117,In_736,In_559);
and U3118 (N_3118,In_1512,In_2410);
or U3119 (N_3119,In_416,In_2464);
xor U3120 (N_3120,In_373,In_1458);
xnor U3121 (N_3121,In_663,In_1989);
and U3122 (N_3122,In_64,In_1975);
or U3123 (N_3123,In_1654,In_1289);
or U3124 (N_3124,In_480,In_947);
and U3125 (N_3125,In_954,In_1886);
or U3126 (N_3126,In_2718,In_28);
and U3127 (N_3127,In_2564,In_2381);
nand U3128 (N_3128,In_1659,In_1512);
xor U3129 (N_3129,In_1130,In_228);
or U3130 (N_3130,In_666,In_303);
and U3131 (N_3131,In_2583,In_1585);
nor U3132 (N_3132,In_979,In_1820);
nand U3133 (N_3133,In_2582,In_1536);
nand U3134 (N_3134,In_187,In_1538);
xor U3135 (N_3135,In_2451,In_1475);
and U3136 (N_3136,In_893,In_1434);
nand U3137 (N_3137,In_577,In_1591);
xnor U3138 (N_3138,In_1456,In_1778);
xnor U3139 (N_3139,In_2791,In_912);
and U3140 (N_3140,In_1340,In_2593);
and U3141 (N_3141,In_1597,In_1200);
xnor U3142 (N_3142,In_1108,In_689);
nand U3143 (N_3143,In_2065,In_2323);
nor U3144 (N_3144,In_248,In_2148);
or U3145 (N_3145,In_1845,In_2860);
nor U3146 (N_3146,In_512,In_2195);
nor U3147 (N_3147,In_2044,In_1860);
nand U3148 (N_3148,In_1944,In_2276);
or U3149 (N_3149,In_2495,In_2482);
and U3150 (N_3150,In_1156,In_1712);
nor U3151 (N_3151,In_1825,In_786);
xor U3152 (N_3152,In_904,In_1167);
and U3153 (N_3153,In_1410,In_246);
and U3154 (N_3154,In_26,In_2581);
and U3155 (N_3155,In_90,In_12);
or U3156 (N_3156,In_831,In_1458);
xor U3157 (N_3157,In_2900,In_2680);
or U3158 (N_3158,In_1436,In_1716);
nand U3159 (N_3159,In_668,In_2337);
nand U3160 (N_3160,In_2162,In_1620);
nor U3161 (N_3161,In_1640,In_1088);
and U3162 (N_3162,In_1786,In_1606);
nor U3163 (N_3163,In_2805,In_1783);
nor U3164 (N_3164,In_727,In_2056);
or U3165 (N_3165,In_827,In_2838);
and U3166 (N_3166,In_910,In_954);
and U3167 (N_3167,In_157,In_1288);
nor U3168 (N_3168,In_1486,In_328);
or U3169 (N_3169,In_355,In_1471);
nand U3170 (N_3170,In_156,In_602);
and U3171 (N_3171,In_2554,In_1894);
nand U3172 (N_3172,In_1666,In_683);
xnor U3173 (N_3173,In_1843,In_2375);
nor U3174 (N_3174,In_2507,In_694);
nor U3175 (N_3175,In_2137,In_1545);
nand U3176 (N_3176,In_95,In_1003);
and U3177 (N_3177,In_2679,In_2255);
nor U3178 (N_3178,In_2524,In_1462);
xnor U3179 (N_3179,In_1,In_1598);
nor U3180 (N_3180,In_1631,In_2804);
and U3181 (N_3181,In_2306,In_2546);
nand U3182 (N_3182,In_2667,In_1383);
and U3183 (N_3183,In_1461,In_1599);
nand U3184 (N_3184,In_372,In_1176);
nor U3185 (N_3185,In_709,In_204);
xor U3186 (N_3186,In_1138,In_1157);
or U3187 (N_3187,In_1156,In_981);
nand U3188 (N_3188,In_2321,In_2310);
nand U3189 (N_3189,In_322,In_2260);
and U3190 (N_3190,In_1993,In_1470);
xnor U3191 (N_3191,In_941,In_812);
and U3192 (N_3192,In_2827,In_500);
nand U3193 (N_3193,In_2659,In_837);
and U3194 (N_3194,In_2682,In_1432);
or U3195 (N_3195,In_2590,In_360);
xnor U3196 (N_3196,In_888,In_2597);
nand U3197 (N_3197,In_299,In_1962);
xor U3198 (N_3198,In_1655,In_1672);
or U3199 (N_3199,In_467,In_1160);
nor U3200 (N_3200,In_764,In_1468);
nand U3201 (N_3201,In_622,In_1491);
and U3202 (N_3202,In_401,In_2400);
nand U3203 (N_3203,In_2221,In_624);
xnor U3204 (N_3204,In_2145,In_2088);
xor U3205 (N_3205,In_2305,In_933);
nor U3206 (N_3206,In_2434,In_1829);
and U3207 (N_3207,In_1950,In_2209);
or U3208 (N_3208,In_1290,In_1242);
and U3209 (N_3209,In_386,In_1415);
nand U3210 (N_3210,In_895,In_2071);
and U3211 (N_3211,In_1533,In_1915);
and U3212 (N_3212,In_2316,In_2068);
nor U3213 (N_3213,In_2950,In_2737);
xnor U3214 (N_3214,In_1372,In_1012);
nand U3215 (N_3215,In_2969,In_512);
or U3216 (N_3216,In_691,In_422);
or U3217 (N_3217,In_685,In_2811);
xor U3218 (N_3218,In_2060,In_123);
nand U3219 (N_3219,In_2780,In_2824);
nand U3220 (N_3220,In_12,In_1367);
and U3221 (N_3221,In_2733,In_328);
nand U3222 (N_3222,In_2843,In_691);
xnor U3223 (N_3223,In_1772,In_2090);
and U3224 (N_3224,In_1121,In_808);
xnor U3225 (N_3225,In_26,In_1542);
nor U3226 (N_3226,In_1234,In_1604);
nor U3227 (N_3227,In_2809,In_1140);
and U3228 (N_3228,In_323,In_2895);
or U3229 (N_3229,In_381,In_1667);
xor U3230 (N_3230,In_601,In_924);
xnor U3231 (N_3231,In_2057,In_2135);
nor U3232 (N_3232,In_1914,In_961);
and U3233 (N_3233,In_2820,In_1428);
or U3234 (N_3234,In_1599,In_1983);
xor U3235 (N_3235,In_100,In_710);
nand U3236 (N_3236,In_2344,In_2427);
nand U3237 (N_3237,In_1906,In_1030);
nor U3238 (N_3238,In_2560,In_2800);
nand U3239 (N_3239,In_22,In_2934);
or U3240 (N_3240,In_1034,In_1213);
nor U3241 (N_3241,In_2350,In_2143);
and U3242 (N_3242,In_1464,In_2285);
or U3243 (N_3243,In_1422,In_2561);
xor U3244 (N_3244,In_1685,In_1018);
and U3245 (N_3245,In_2529,In_21);
nor U3246 (N_3246,In_7,In_1806);
or U3247 (N_3247,In_967,In_1469);
nand U3248 (N_3248,In_726,In_1761);
or U3249 (N_3249,In_986,In_1896);
xnor U3250 (N_3250,In_945,In_1200);
or U3251 (N_3251,In_801,In_2454);
nand U3252 (N_3252,In_1804,In_1680);
or U3253 (N_3253,In_2763,In_2329);
nand U3254 (N_3254,In_2876,In_2488);
or U3255 (N_3255,In_399,In_2805);
nand U3256 (N_3256,In_2133,In_1033);
nand U3257 (N_3257,In_2739,In_1429);
or U3258 (N_3258,In_1658,In_560);
xor U3259 (N_3259,In_1089,In_2008);
nand U3260 (N_3260,In_2775,In_2366);
nor U3261 (N_3261,In_1901,In_24);
and U3262 (N_3262,In_1769,In_704);
and U3263 (N_3263,In_2864,In_1619);
nor U3264 (N_3264,In_2417,In_2351);
nor U3265 (N_3265,In_496,In_1144);
or U3266 (N_3266,In_753,In_208);
or U3267 (N_3267,In_801,In_1166);
xnor U3268 (N_3268,In_1555,In_134);
nand U3269 (N_3269,In_2956,In_1242);
nand U3270 (N_3270,In_69,In_1019);
nand U3271 (N_3271,In_2189,In_2309);
nor U3272 (N_3272,In_1612,In_2597);
xnor U3273 (N_3273,In_1068,In_1868);
nor U3274 (N_3274,In_475,In_134);
or U3275 (N_3275,In_147,In_711);
and U3276 (N_3276,In_2796,In_1357);
and U3277 (N_3277,In_791,In_1124);
and U3278 (N_3278,In_1473,In_1402);
or U3279 (N_3279,In_2208,In_1144);
or U3280 (N_3280,In_1988,In_8);
nor U3281 (N_3281,In_2594,In_2968);
xor U3282 (N_3282,In_1227,In_1911);
xnor U3283 (N_3283,In_2802,In_397);
nor U3284 (N_3284,In_1654,In_673);
nor U3285 (N_3285,In_2125,In_2655);
xnor U3286 (N_3286,In_305,In_143);
nand U3287 (N_3287,In_1292,In_945);
xor U3288 (N_3288,In_159,In_7);
and U3289 (N_3289,In_2251,In_2395);
nand U3290 (N_3290,In_2415,In_1619);
xnor U3291 (N_3291,In_2329,In_72);
xor U3292 (N_3292,In_576,In_1902);
xor U3293 (N_3293,In_2195,In_394);
xnor U3294 (N_3294,In_833,In_1772);
or U3295 (N_3295,In_2444,In_2652);
or U3296 (N_3296,In_866,In_987);
or U3297 (N_3297,In_1630,In_2367);
or U3298 (N_3298,In_1463,In_2990);
nor U3299 (N_3299,In_1391,In_517);
and U3300 (N_3300,In_2474,In_1543);
nand U3301 (N_3301,In_1458,In_1968);
xnor U3302 (N_3302,In_309,In_1626);
and U3303 (N_3303,In_1022,In_1946);
nand U3304 (N_3304,In_2323,In_834);
or U3305 (N_3305,In_2589,In_2159);
and U3306 (N_3306,In_2504,In_1058);
nand U3307 (N_3307,In_2929,In_420);
xnor U3308 (N_3308,In_697,In_364);
nand U3309 (N_3309,In_2068,In_391);
nand U3310 (N_3310,In_1285,In_621);
or U3311 (N_3311,In_81,In_2688);
xor U3312 (N_3312,In_1693,In_1746);
nor U3313 (N_3313,In_723,In_661);
xnor U3314 (N_3314,In_2119,In_1660);
nor U3315 (N_3315,In_349,In_50);
nor U3316 (N_3316,In_2742,In_2138);
and U3317 (N_3317,In_1644,In_550);
xor U3318 (N_3318,In_709,In_2100);
and U3319 (N_3319,In_299,In_2267);
nor U3320 (N_3320,In_2198,In_962);
or U3321 (N_3321,In_2499,In_1890);
nand U3322 (N_3322,In_2177,In_995);
nor U3323 (N_3323,In_188,In_1460);
nor U3324 (N_3324,In_468,In_24);
nor U3325 (N_3325,In_1390,In_2134);
nand U3326 (N_3326,In_2642,In_2129);
or U3327 (N_3327,In_2398,In_2917);
or U3328 (N_3328,In_2401,In_1095);
nand U3329 (N_3329,In_532,In_2179);
nor U3330 (N_3330,In_2360,In_2420);
or U3331 (N_3331,In_930,In_1616);
nand U3332 (N_3332,In_1056,In_1430);
nand U3333 (N_3333,In_1525,In_1688);
nand U3334 (N_3334,In_1089,In_2964);
or U3335 (N_3335,In_1659,In_1048);
nand U3336 (N_3336,In_1577,In_2907);
and U3337 (N_3337,In_1439,In_1121);
nor U3338 (N_3338,In_2492,In_1624);
nand U3339 (N_3339,In_1667,In_2025);
and U3340 (N_3340,In_2514,In_624);
or U3341 (N_3341,In_584,In_2418);
nand U3342 (N_3342,In_1333,In_1978);
nor U3343 (N_3343,In_237,In_1291);
nor U3344 (N_3344,In_2324,In_663);
nand U3345 (N_3345,In_987,In_67);
and U3346 (N_3346,In_1854,In_420);
nand U3347 (N_3347,In_378,In_45);
xnor U3348 (N_3348,In_1799,In_2878);
nand U3349 (N_3349,In_2871,In_2138);
or U3350 (N_3350,In_495,In_1791);
nor U3351 (N_3351,In_2677,In_2592);
xnor U3352 (N_3352,In_2488,In_2617);
or U3353 (N_3353,In_547,In_999);
and U3354 (N_3354,In_2813,In_2784);
nand U3355 (N_3355,In_853,In_342);
xnor U3356 (N_3356,In_1587,In_1382);
xnor U3357 (N_3357,In_1177,In_2704);
nand U3358 (N_3358,In_2537,In_1904);
xor U3359 (N_3359,In_283,In_2169);
nor U3360 (N_3360,In_2555,In_2381);
nand U3361 (N_3361,In_1757,In_29);
and U3362 (N_3362,In_507,In_1181);
nor U3363 (N_3363,In_1461,In_2337);
or U3364 (N_3364,In_302,In_2319);
and U3365 (N_3365,In_1507,In_1038);
or U3366 (N_3366,In_2863,In_634);
nor U3367 (N_3367,In_1656,In_1102);
or U3368 (N_3368,In_1790,In_228);
nor U3369 (N_3369,In_645,In_2608);
xnor U3370 (N_3370,In_1448,In_251);
and U3371 (N_3371,In_2987,In_1773);
or U3372 (N_3372,In_1040,In_2944);
and U3373 (N_3373,In_1910,In_2586);
xnor U3374 (N_3374,In_1048,In_1359);
xnor U3375 (N_3375,In_418,In_2319);
and U3376 (N_3376,In_467,In_2774);
nand U3377 (N_3377,In_1971,In_1923);
or U3378 (N_3378,In_767,In_2901);
nand U3379 (N_3379,In_2267,In_1102);
nand U3380 (N_3380,In_2364,In_1012);
or U3381 (N_3381,In_40,In_851);
nor U3382 (N_3382,In_2583,In_804);
xnor U3383 (N_3383,In_1761,In_2541);
xor U3384 (N_3384,In_994,In_573);
xnor U3385 (N_3385,In_12,In_1800);
nand U3386 (N_3386,In_1158,In_1099);
and U3387 (N_3387,In_2764,In_1681);
nor U3388 (N_3388,In_1736,In_2902);
nor U3389 (N_3389,In_2518,In_2401);
or U3390 (N_3390,In_1477,In_1699);
xnor U3391 (N_3391,In_1247,In_1293);
xor U3392 (N_3392,In_735,In_961);
xnor U3393 (N_3393,In_1784,In_1005);
and U3394 (N_3394,In_1213,In_1961);
xnor U3395 (N_3395,In_2095,In_504);
and U3396 (N_3396,In_1677,In_691);
nand U3397 (N_3397,In_554,In_1732);
or U3398 (N_3398,In_281,In_2160);
and U3399 (N_3399,In_1255,In_983);
and U3400 (N_3400,In_1195,In_253);
and U3401 (N_3401,In_1537,In_2869);
or U3402 (N_3402,In_151,In_796);
nor U3403 (N_3403,In_604,In_2715);
nor U3404 (N_3404,In_124,In_2142);
nand U3405 (N_3405,In_258,In_1644);
nor U3406 (N_3406,In_628,In_1020);
and U3407 (N_3407,In_671,In_1463);
nand U3408 (N_3408,In_764,In_1358);
nor U3409 (N_3409,In_1016,In_2910);
nand U3410 (N_3410,In_2074,In_1970);
and U3411 (N_3411,In_2064,In_122);
nand U3412 (N_3412,In_2482,In_2915);
nand U3413 (N_3413,In_2843,In_1530);
or U3414 (N_3414,In_444,In_2310);
nor U3415 (N_3415,In_2194,In_1329);
and U3416 (N_3416,In_654,In_1997);
or U3417 (N_3417,In_2159,In_2440);
xor U3418 (N_3418,In_2515,In_1341);
nand U3419 (N_3419,In_108,In_2360);
nor U3420 (N_3420,In_930,In_1790);
nor U3421 (N_3421,In_2321,In_1107);
nor U3422 (N_3422,In_609,In_91);
nor U3423 (N_3423,In_1766,In_1036);
and U3424 (N_3424,In_2364,In_814);
xor U3425 (N_3425,In_1108,In_279);
xnor U3426 (N_3426,In_2731,In_10);
nor U3427 (N_3427,In_968,In_2079);
xor U3428 (N_3428,In_945,In_590);
nor U3429 (N_3429,In_1662,In_2989);
nand U3430 (N_3430,In_650,In_1937);
and U3431 (N_3431,In_102,In_2227);
xor U3432 (N_3432,In_2024,In_2267);
xnor U3433 (N_3433,In_2369,In_2003);
xnor U3434 (N_3434,In_1546,In_2933);
xor U3435 (N_3435,In_2054,In_2160);
and U3436 (N_3436,In_2202,In_1621);
and U3437 (N_3437,In_780,In_2542);
or U3438 (N_3438,In_1568,In_1550);
xor U3439 (N_3439,In_1643,In_1648);
xor U3440 (N_3440,In_2563,In_2891);
and U3441 (N_3441,In_1154,In_1141);
xor U3442 (N_3442,In_2162,In_694);
or U3443 (N_3443,In_846,In_2164);
and U3444 (N_3444,In_102,In_2746);
or U3445 (N_3445,In_978,In_997);
nand U3446 (N_3446,In_95,In_2648);
and U3447 (N_3447,In_1303,In_2920);
nor U3448 (N_3448,In_1801,In_782);
nor U3449 (N_3449,In_1101,In_1820);
nor U3450 (N_3450,In_2853,In_1709);
and U3451 (N_3451,In_119,In_776);
and U3452 (N_3452,In_477,In_511);
and U3453 (N_3453,In_2812,In_1574);
xor U3454 (N_3454,In_935,In_2371);
nor U3455 (N_3455,In_49,In_20);
or U3456 (N_3456,In_1071,In_931);
and U3457 (N_3457,In_432,In_482);
nand U3458 (N_3458,In_1794,In_973);
nor U3459 (N_3459,In_324,In_1252);
and U3460 (N_3460,In_2979,In_1007);
or U3461 (N_3461,In_2915,In_1746);
nand U3462 (N_3462,In_2980,In_609);
nand U3463 (N_3463,In_1489,In_143);
nor U3464 (N_3464,In_92,In_2153);
xnor U3465 (N_3465,In_2377,In_2341);
nand U3466 (N_3466,In_2381,In_1185);
xnor U3467 (N_3467,In_1871,In_2720);
and U3468 (N_3468,In_357,In_2324);
nand U3469 (N_3469,In_1788,In_546);
xor U3470 (N_3470,In_1444,In_2629);
nor U3471 (N_3471,In_2926,In_1015);
or U3472 (N_3472,In_542,In_1883);
or U3473 (N_3473,In_2140,In_1518);
or U3474 (N_3474,In_1516,In_2264);
nand U3475 (N_3475,In_1943,In_1078);
nand U3476 (N_3476,In_918,In_1425);
xnor U3477 (N_3477,In_894,In_2311);
or U3478 (N_3478,In_1938,In_1739);
xnor U3479 (N_3479,In_1903,In_1699);
nand U3480 (N_3480,In_1748,In_310);
xor U3481 (N_3481,In_1109,In_1875);
or U3482 (N_3482,In_1794,In_1007);
and U3483 (N_3483,In_724,In_593);
or U3484 (N_3484,In_2583,In_863);
nor U3485 (N_3485,In_1899,In_1025);
nand U3486 (N_3486,In_2370,In_2779);
and U3487 (N_3487,In_208,In_1297);
nand U3488 (N_3488,In_38,In_1044);
and U3489 (N_3489,In_411,In_863);
xor U3490 (N_3490,In_1384,In_1463);
xor U3491 (N_3491,In_2022,In_1887);
and U3492 (N_3492,In_1353,In_1038);
and U3493 (N_3493,In_717,In_1612);
or U3494 (N_3494,In_1474,In_1561);
or U3495 (N_3495,In_1026,In_367);
nand U3496 (N_3496,In_228,In_838);
nand U3497 (N_3497,In_2959,In_2379);
nor U3498 (N_3498,In_480,In_2966);
xnor U3499 (N_3499,In_732,In_330);
nor U3500 (N_3500,In_293,In_402);
xnor U3501 (N_3501,In_1399,In_1148);
nand U3502 (N_3502,In_2175,In_1051);
nor U3503 (N_3503,In_574,In_2333);
nor U3504 (N_3504,In_288,In_1902);
xor U3505 (N_3505,In_2926,In_434);
nand U3506 (N_3506,In_2430,In_2499);
nand U3507 (N_3507,In_909,In_714);
nor U3508 (N_3508,In_1135,In_620);
xor U3509 (N_3509,In_2296,In_2864);
and U3510 (N_3510,In_2105,In_758);
xor U3511 (N_3511,In_2003,In_1101);
or U3512 (N_3512,In_2493,In_2026);
or U3513 (N_3513,In_2903,In_104);
nand U3514 (N_3514,In_1624,In_2338);
nand U3515 (N_3515,In_988,In_911);
or U3516 (N_3516,In_2269,In_2069);
or U3517 (N_3517,In_2650,In_1311);
nand U3518 (N_3518,In_1962,In_202);
and U3519 (N_3519,In_1117,In_974);
or U3520 (N_3520,In_1329,In_2507);
xor U3521 (N_3521,In_675,In_2763);
xor U3522 (N_3522,In_2232,In_2482);
or U3523 (N_3523,In_1743,In_397);
and U3524 (N_3524,In_93,In_2311);
and U3525 (N_3525,In_1944,In_932);
nor U3526 (N_3526,In_2303,In_1609);
xnor U3527 (N_3527,In_93,In_1353);
nor U3528 (N_3528,In_1854,In_237);
nor U3529 (N_3529,In_70,In_1848);
and U3530 (N_3530,In_1098,In_1894);
or U3531 (N_3531,In_1027,In_597);
nand U3532 (N_3532,In_1605,In_558);
nand U3533 (N_3533,In_463,In_2346);
nor U3534 (N_3534,In_1245,In_2935);
nor U3535 (N_3535,In_1906,In_2195);
or U3536 (N_3536,In_739,In_471);
nor U3537 (N_3537,In_1181,In_1448);
and U3538 (N_3538,In_2646,In_1293);
nor U3539 (N_3539,In_440,In_2856);
and U3540 (N_3540,In_573,In_1782);
xor U3541 (N_3541,In_773,In_1130);
or U3542 (N_3542,In_370,In_683);
nor U3543 (N_3543,In_1831,In_2938);
nor U3544 (N_3544,In_2610,In_1815);
nand U3545 (N_3545,In_2536,In_2339);
nand U3546 (N_3546,In_2851,In_2398);
or U3547 (N_3547,In_1768,In_1493);
nand U3548 (N_3548,In_466,In_2529);
and U3549 (N_3549,In_1952,In_715);
or U3550 (N_3550,In_2056,In_1374);
nor U3551 (N_3551,In_2956,In_1346);
nand U3552 (N_3552,In_2643,In_1817);
xor U3553 (N_3553,In_2534,In_672);
xor U3554 (N_3554,In_1361,In_2192);
nor U3555 (N_3555,In_1310,In_2818);
nand U3556 (N_3556,In_2417,In_2485);
and U3557 (N_3557,In_1933,In_601);
nand U3558 (N_3558,In_542,In_1276);
or U3559 (N_3559,In_649,In_388);
or U3560 (N_3560,In_810,In_2684);
or U3561 (N_3561,In_1808,In_1259);
nor U3562 (N_3562,In_1544,In_80);
and U3563 (N_3563,In_2305,In_854);
nor U3564 (N_3564,In_1420,In_663);
and U3565 (N_3565,In_505,In_1873);
nor U3566 (N_3566,In_629,In_1267);
nor U3567 (N_3567,In_2136,In_673);
nand U3568 (N_3568,In_579,In_1704);
xnor U3569 (N_3569,In_2232,In_1259);
nand U3570 (N_3570,In_1446,In_2050);
or U3571 (N_3571,In_2402,In_2994);
nor U3572 (N_3572,In_424,In_1980);
nand U3573 (N_3573,In_1847,In_2397);
or U3574 (N_3574,In_14,In_1946);
xnor U3575 (N_3575,In_2550,In_1059);
nand U3576 (N_3576,In_2456,In_2276);
xor U3577 (N_3577,In_1613,In_1703);
xnor U3578 (N_3578,In_2061,In_1043);
nand U3579 (N_3579,In_2864,In_2320);
nand U3580 (N_3580,In_2272,In_2639);
xnor U3581 (N_3581,In_785,In_10);
nand U3582 (N_3582,In_1522,In_1947);
nand U3583 (N_3583,In_1228,In_266);
or U3584 (N_3584,In_1885,In_1893);
nor U3585 (N_3585,In_405,In_1606);
or U3586 (N_3586,In_2803,In_574);
nand U3587 (N_3587,In_1399,In_2157);
and U3588 (N_3588,In_2503,In_629);
and U3589 (N_3589,In_1772,In_1133);
nand U3590 (N_3590,In_476,In_1753);
nor U3591 (N_3591,In_791,In_1089);
xor U3592 (N_3592,In_2584,In_2305);
xnor U3593 (N_3593,In_384,In_2344);
and U3594 (N_3594,In_891,In_1138);
nand U3595 (N_3595,In_2099,In_1034);
nor U3596 (N_3596,In_2621,In_1201);
or U3597 (N_3597,In_2263,In_740);
and U3598 (N_3598,In_2648,In_1553);
nand U3599 (N_3599,In_1878,In_1124);
xnor U3600 (N_3600,In_324,In_2570);
xnor U3601 (N_3601,In_1080,In_2407);
or U3602 (N_3602,In_2799,In_354);
or U3603 (N_3603,In_1440,In_2740);
nand U3604 (N_3604,In_2553,In_860);
xor U3605 (N_3605,In_1845,In_2448);
xor U3606 (N_3606,In_2285,In_425);
or U3607 (N_3607,In_949,In_369);
nand U3608 (N_3608,In_794,In_2401);
nand U3609 (N_3609,In_741,In_565);
and U3610 (N_3610,In_2877,In_2980);
nand U3611 (N_3611,In_596,In_1858);
nor U3612 (N_3612,In_1234,In_2026);
xor U3613 (N_3613,In_1850,In_1076);
nand U3614 (N_3614,In_1724,In_2028);
xor U3615 (N_3615,In_752,In_1218);
or U3616 (N_3616,In_60,In_1683);
and U3617 (N_3617,In_2958,In_2387);
and U3618 (N_3618,In_1223,In_1816);
or U3619 (N_3619,In_1672,In_293);
and U3620 (N_3620,In_497,In_1832);
nor U3621 (N_3621,In_1561,In_2085);
nand U3622 (N_3622,In_2617,In_2590);
nand U3623 (N_3623,In_2979,In_2683);
nand U3624 (N_3624,In_1926,In_127);
nand U3625 (N_3625,In_424,In_1217);
and U3626 (N_3626,In_2457,In_1015);
nand U3627 (N_3627,In_149,In_9);
nand U3628 (N_3628,In_802,In_1574);
xor U3629 (N_3629,In_519,In_588);
nand U3630 (N_3630,In_665,In_1713);
or U3631 (N_3631,In_1374,In_68);
and U3632 (N_3632,In_1924,In_1929);
nand U3633 (N_3633,In_1070,In_952);
nor U3634 (N_3634,In_1263,In_1515);
and U3635 (N_3635,In_1580,In_654);
and U3636 (N_3636,In_639,In_2287);
nor U3637 (N_3637,In_589,In_1216);
or U3638 (N_3638,In_919,In_531);
or U3639 (N_3639,In_2113,In_2519);
and U3640 (N_3640,In_1060,In_262);
nor U3641 (N_3641,In_2390,In_1891);
nand U3642 (N_3642,In_523,In_1287);
nand U3643 (N_3643,In_642,In_869);
nand U3644 (N_3644,In_2266,In_1072);
nor U3645 (N_3645,In_1307,In_31);
xor U3646 (N_3646,In_2459,In_1423);
and U3647 (N_3647,In_2960,In_568);
and U3648 (N_3648,In_2537,In_2224);
or U3649 (N_3649,In_2121,In_2780);
nand U3650 (N_3650,In_1678,In_1575);
xor U3651 (N_3651,In_1652,In_1660);
or U3652 (N_3652,In_207,In_2168);
and U3653 (N_3653,In_1436,In_2566);
or U3654 (N_3654,In_1468,In_855);
or U3655 (N_3655,In_1966,In_1497);
xnor U3656 (N_3656,In_1100,In_1587);
nor U3657 (N_3657,In_844,In_2096);
nor U3658 (N_3658,In_1136,In_1721);
xnor U3659 (N_3659,In_1674,In_520);
nor U3660 (N_3660,In_2720,In_2409);
or U3661 (N_3661,In_2641,In_2478);
and U3662 (N_3662,In_1016,In_455);
nor U3663 (N_3663,In_1836,In_458);
or U3664 (N_3664,In_1999,In_78);
xor U3665 (N_3665,In_2973,In_1664);
xnor U3666 (N_3666,In_1066,In_1058);
or U3667 (N_3667,In_577,In_171);
xor U3668 (N_3668,In_1918,In_2143);
nand U3669 (N_3669,In_2381,In_2123);
and U3670 (N_3670,In_1931,In_236);
and U3671 (N_3671,In_60,In_265);
xor U3672 (N_3672,In_1548,In_1452);
or U3673 (N_3673,In_1326,In_859);
xor U3674 (N_3674,In_550,In_2839);
nand U3675 (N_3675,In_141,In_575);
and U3676 (N_3676,In_1444,In_685);
xor U3677 (N_3677,In_1371,In_631);
and U3678 (N_3678,In_316,In_2951);
and U3679 (N_3679,In_2502,In_2965);
or U3680 (N_3680,In_1520,In_750);
nand U3681 (N_3681,In_340,In_2348);
xor U3682 (N_3682,In_357,In_2416);
or U3683 (N_3683,In_733,In_1233);
nand U3684 (N_3684,In_1917,In_2493);
nor U3685 (N_3685,In_1559,In_550);
nand U3686 (N_3686,In_1046,In_1510);
xnor U3687 (N_3687,In_2423,In_2460);
nand U3688 (N_3688,In_1186,In_979);
or U3689 (N_3689,In_2999,In_2449);
and U3690 (N_3690,In_1595,In_2211);
nor U3691 (N_3691,In_2985,In_1098);
xnor U3692 (N_3692,In_1665,In_1405);
nand U3693 (N_3693,In_2938,In_2203);
or U3694 (N_3694,In_1790,In_1488);
or U3695 (N_3695,In_820,In_2343);
nand U3696 (N_3696,In_2875,In_822);
nor U3697 (N_3697,In_68,In_1659);
nand U3698 (N_3698,In_2641,In_735);
or U3699 (N_3699,In_2098,In_2061);
nand U3700 (N_3700,In_2993,In_2929);
xnor U3701 (N_3701,In_869,In_1944);
nand U3702 (N_3702,In_575,In_737);
xnor U3703 (N_3703,In_257,In_1192);
nand U3704 (N_3704,In_2506,In_875);
nor U3705 (N_3705,In_1099,In_2537);
nor U3706 (N_3706,In_461,In_1500);
nand U3707 (N_3707,In_2582,In_2012);
nor U3708 (N_3708,In_2394,In_1351);
nand U3709 (N_3709,In_2412,In_946);
xor U3710 (N_3710,In_2036,In_234);
or U3711 (N_3711,In_898,In_1116);
or U3712 (N_3712,In_1465,In_2689);
xor U3713 (N_3713,In_970,In_450);
xnor U3714 (N_3714,In_2589,In_1946);
and U3715 (N_3715,In_2782,In_2691);
and U3716 (N_3716,In_2498,In_1257);
xor U3717 (N_3717,In_1834,In_106);
nor U3718 (N_3718,In_1980,In_219);
xnor U3719 (N_3719,In_1217,In_1525);
xnor U3720 (N_3720,In_1588,In_1953);
or U3721 (N_3721,In_2767,In_153);
nand U3722 (N_3722,In_1646,In_2662);
nor U3723 (N_3723,In_1503,In_2074);
xnor U3724 (N_3724,In_900,In_1212);
and U3725 (N_3725,In_1544,In_2378);
nor U3726 (N_3726,In_1653,In_1441);
and U3727 (N_3727,In_2421,In_1504);
xor U3728 (N_3728,In_635,In_2475);
nand U3729 (N_3729,In_1958,In_478);
xnor U3730 (N_3730,In_1135,In_1036);
nor U3731 (N_3731,In_343,In_1486);
or U3732 (N_3732,In_2919,In_2803);
xor U3733 (N_3733,In_94,In_1408);
nor U3734 (N_3734,In_1714,In_1241);
and U3735 (N_3735,In_2712,In_2357);
nand U3736 (N_3736,In_21,In_1465);
or U3737 (N_3737,In_554,In_1659);
nor U3738 (N_3738,In_1904,In_812);
xor U3739 (N_3739,In_751,In_2295);
and U3740 (N_3740,In_2499,In_2535);
xnor U3741 (N_3741,In_2669,In_2067);
and U3742 (N_3742,In_2947,In_1007);
or U3743 (N_3743,In_1122,In_2410);
and U3744 (N_3744,In_256,In_1266);
or U3745 (N_3745,In_2333,In_1918);
nor U3746 (N_3746,In_2013,In_47);
nand U3747 (N_3747,In_143,In_519);
nand U3748 (N_3748,In_2416,In_1984);
xor U3749 (N_3749,In_2247,In_2503);
nand U3750 (N_3750,In_769,In_913);
and U3751 (N_3751,In_2354,In_1394);
and U3752 (N_3752,In_66,In_2536);
nor U3753 (N_3753,In_2711,In_2093);
or U3754 (N_3754,In_2178,In_1219);
nor U3755 (N_3755,In_1663,In_752);
or U3756 (N_3756,In_2879,In_2609);
or U3757 (N_3757,In_594,In_1221);
nor U3758 (N_3758,In_1943,In_1624);
nand U3759 (N_3759,In_1189,In_550);
nand U3760 (N_3760,In_1840,In_982);
nor U3761 (N_3761,In_1953,In_156);
nand U3762 (N_3762,In_403,In_2648);
or U3763 (N_3763,In_2458,In_2929);
nand U3764 (N_3764,In_1787,In_222);
xnor U3765 (N_3765,In_1963,In_1882);
nor U3766 (N_3766,In_193,In_2949);
or U3767 (N_3767,In_2652,In_2161);
and U3768 (N_3768,In_473,In_1460);
xnor U3769 (N_3769,In_1715,In_117);
or U3770 (N_3770,In_281,In_1355);
nor U3771 (N_3771,In_534,In_2676);
nor U3772 (N_3772,In_204,In_417);
and U3773 (N_3773,In_1734,In_2278);
and U3774 (N_3774,In_1806,In_266);
nor U3775 (N_3775,In_467,In_2895);
or U3776 (N_3776,In_2461,In_274);
or U3777 (N_3777,In_1316,In_2933);
nor U3778 (N_3778,In_2755,In_100);
or U3779 (N_3779,In_1234,In_1515);
and U3780 (N_3780,In_922,In_1424);
nor U3781 (N_3781,In_231,In_1098);
nand U3782 (N_3782,In_2109,In_1856);
or U3783 (N_3783,In_1811,In_2313);
and U3784 (N_3784,In_862,In_2808);
or U3785 (N_3785,In_2906,In_2501);
and U3786 (N_3786,In_486,In_1074);
nand U3787 (N_3787,In_1011,In_2955);
and U3788 (N_3788,In_1086,In_2114);
nor U3789 (N_3789,In_332,In_1203);
or U3790 (N_3790,In_1319,In_376);
and U3791 (N_3791,In_2976,In_1270);
or U3792 (N_3792,In_31,In_175);
and U3793 (N_3793,In_1473,In_2585);
nand U3794 (N_3794,In_1454,In_2768);
nor U3795 (N_3795,In_2278,In_1557);
or U3796 (N_3796,In_286,In_1787);
nand U3797 (N_3797,In_133,In_2333);
or U3798 (N_3798,In_296,In_1004);
xnor U3799 (N_3799,In_1801,In_2230);
nand U3800 (N_3800,In_2694,In_2025);
nand U3801 (N_3801,In_650,In_125);
xnor U3802 (N_3802,In_2010,In_449);
nand U3803 (N_3803,In_1870,In_1568);
nor U3804 (N_3804,In_2956,In_2350);
xor U3805 (N_3805,In_2651,In_2163);
xnor U3806 (N_3806,In_2800,In_315);
and U3807 (N_3807,In_21,In_1117);
nand U3808 (N_3808,In_2416,In_778);
and U3809 (N_3809,In_2961,In_516);
or U3810 (N_3810,In_1031,In_2320);
xnor U3811 (N_3811,In_1981,In_1756);
xor U3812 (N_3812,In_327,In_2782);
xnor U3813 (N_3813,In_969,In_799);
xor U3814 (N_3814,In_2173,In_2958);
nor U3815 (N_3815,In_458,In_754);
nor U3816 (N_3816,In_2237,In_921);
nor U3817 (N_3817,In_405,In_1013);
nand U3818 (N_3818,In_282,In_2897);
or U3819 (N_3819,In_338,In_1016);
nand U3820 (N_3820,In_2643,In_717);
and U3821 (N_3821,In_336,In_1630);
nor U3822 (N_3822,In_2821,In_272);
xnor U3823 (N_3823,In_965,In_313);
xor U3824 (N_3824,In_2481,In_2565);
xnor U3825 (N_3825,In_1504,In_1884);
or U3826 (N_3826,In_1954,In_405);
or U3827 (N_3827,In_2058,In_914);
and U3828 (N_3828,In_447,In_2608);
and U3829 (N_3829,In_455,In_2736);
and U3830 (N_3830,In_1805,In_670);
and U3831 (N_3831,In_1724,In_1686);
and U3832 (N_3832,In_2638,In_86);
and U3833 (N_3833,In_1923,In_2741);
or U3834 (N_3834,In_382,In_727);
and U3835 (N_3835,In_1567,In_1253);
or U3836 (N_3836,In_2055,In_2197);
nand U3837 (N_3837,In_1279,In_1658);
and U3838 (N_3838,In_715,In_1385);
xor U3839 (N_3839,In_537,In_957);
and U3840 (N_3840,In_2928,In_1423);
nor U3841 (N_3841,In_2900,In_835);
and U3842 (N_3842,In_1806,In_1203);
nor U3843 (N_3843,In_1504,In_511);
or U3844 (N_3844,In_2685,In_1089);
xor U3845 (N_3845,In_2816,In_1663);
and U3846 (N_3846,In_1959,In_1987);
and U3847 (N_3847,In_119,In_2737);
xnor U3848 (N_3848,In_550,In_2800);
or U3849 (N_3849,In_2486,In_2124);
nand U3850 (N_3850,In_2668,In_2286);
nor U3851 (N_3851,In_1327,In_625);
nand U3852 (N_3852,In_1696,In_1565);
or U3853 (N_3853,In_2541,In_1923);
or U3854 (N_3854,In_139,In_526);
nand U3855 (N_3855,In_991,In_502);
or U3856 (N_3856,In_2569,In_211);
nor U3857 (N_3857,In_759,In_1982);
nor U3858 (N_3858,In_2617,In_1736);
nor U3859 (N_3859,In_2758,In_1155);
xnor U3860 (N_3860,In_1090,In_1436);
xnor U3861 (N_3861,In_564,In_71);
nand U3862 (N_3862,In_1667,In_2297);
nand U3863 (N_3863,In_808,In_1892);
and U3864 (N_3864,In_1042,In_1649);
or U3865 (N_3865,In_2706,In_462);
xnor U3866 (N_3866,In_1685,In_2327);
or U3867 (N_3867,In_642,In_485);
nand U3868 (N_3868,In_860,In_1744);
and U3869 (N_3869,In_214,In_2016);
and U3870 (N_3870,In_885,In_1042);
xnor U3871 (N_3871,In_1909,In_1107);
or U3872 (N_3872,In_1722,In_1786);
xnor U3873 (N_3873,In_152,In_1278);
nor U3874 (N_3874,In_1995,In_2145);
nor U3875 (N_3875,In_2583,In_324);
and U3876 (N_3876,In_2865,In_2109);
nor U3877 (N_3877,In_2407,In_1331);
or U3878 (N_3878,In_916,In_2975);
or U3879 (N_3879,In_2860,In_2368);
and U3880 (N_3880,In_2730,In_5);
nand U3881 (N_3881,In_223,In_490);
or U3882 (N_3882,In_1163,In_1917);
xor U3883 (N_3883,In_1475,In_1180);
and U3884 (N_3884,In_272,In_1937);
nor U3885 (N_3885,In_662,In_837);
nand U3886 (N_3886,In_2808,In_2559);
nand U3887 (N_3887,In_2137,In_1574);
or U3888 (N_3888,In_157,In_1304);
nand U3889 (N_3889,In_1686,In_596);
or U3890 (N_3890,In_1372,In_2181);
and U3891 (N_3891,In_1981,In_506);
nand U3892 (N_3892,In_39,In_2950);
or U3893 (N_3893,In_494,In_2296);
nor U3894 (N_3894,In_2170,In_1101);
or U3895 (N_3895,In_1136,In_587);
or U3896 (N_3896,In_559,In_1704);
and U3897 (N_3897,In_1334,In_911);
nand U3898 (N_3898,In_1409,In_148);
xor U3899 (N_3899,In_2149,In_2802);
xnor U3900 (N_3900,In_2028,In_725);
or U3901 (N_3901,In_1380,In_90);
or U3902 (N_3902,In_2106,In_665);
and U3903 (N_3903,In_2334,In_1854);
and U3904 (N_3904,In_2166,In_754);
nand U3905 (N_3905,In_1042,In_2043);
and U3906 (N_3906,In_283,In_671);
and U3907 (N_3907,In_2337,In_1017);
nand U3908 (N_3908,In_405,In_1887);
and U3909 (N_3909,In_2901,In_1498);
xnor U3910 (N_3910,In_885,In_541);
nand U3911 (N_3911,In_2628,In_507);
or U3912 (N_3912,In_1750,In_120);
nor U3913 (N_3913,In_2059,In_395);
or U3914 (N_3914,In_812,In_2653);
or U3915 (N_3915,In_1200,In_2985);
and U3916 (N_3916,In_1519,In_1624);
nor U3917 (N_3917,In_1472,In_1414);
nor U3918 (N_3918,In_1337,In_1879);
nand U3919 (N_3919,In_2655,In_958);
nor U3920 (N_3920,In_706,In_75);
or U3921 (N_3921,In_819,In_521);
xnor U3922 (N_3922,In_941,In_1763);
or U3923 (N_3923,In_2433,In_920);
xor U3924 (N_3924,In_492,In_374);
nand U3925 (N_3925,In_2222,In_563);
or U3926 (N_3926,In_1668,In_2123);
or U3927 (N_3927,In_455,In_2026);
xor U3928 (N_3928,In_2519,In_1746);
or U3929 (N_3929,In_1839,In_2403);
nor U3930 (N_3930,In_1215,In_2738);
xnor U3931 (N_3931,In_376,In_658);
nor U3932 (N_3932,In_1043,In_2177);
xor U3933 (N_3933,In_1370,In_1132);
xor U3934 (N_3934,In_2389,In_1037);
or U3935 (N_3935,In_889,In_1983);
nand U3936 (N_3936,In_161,In_2571);
nand U3937 (N_3937,In_2664,In_2498);
and U3938 (N_3938,In_2689,In_1566);
nand U3939 (N_3939,In_174,In_1105);
xor U3940 (N_3940,In_2289,In_2124);
nand U3941 (N_3941,In_360,In_1777);
or U3942 (N_3942,In_466,In_330);
nand U3943 (N_3943,In_1572,In_1762);
nand U3944 (N_3944,In_535,In_1852);
and U3945 (N_3945,In_1154,In_655);
xor U3946 (N_3946,In_473,In_98);
and U3947 (N_3947,In_2136,In_8);
or U3948 (N_3948,In_2352,In_2107);
nor U3949 (N_3949,In_2418,In_1243);
nand U3950 (N_3950,In_542,In_1460);
nand U3951 (N_3951,In_286,In_762);
xnor U3952 (N_3952,In_900,In_2408);
nor U3953 (N_3953,In_2484,In_2420);
nand U3954 (N_3954,In_2931,In_2589);
xnor U3955 (N_3955,In_2727,In_270);
nor U3956 (N_3956,In_607,In_2182);
and U3957 (N_3957,In_896,In_599);
or U3958 (N_3958,In_1264,In_2987);
and U3959 (N_3959,In_818,In_2573);
xor U3960 (N_3960,In_344,In_733);
xnor U3961 (N_3961,In_2051,In_2362);
nand U3962 (N_3962,In_1742,In_2092);
nor U3963 (N_3963,In_2552,In_1132);
and U3964 (N_3964,In_2599,In_293);
xor U3965 (N_3965,In_2262,In_311);
nand U3966 (N_3966,In_1128,In_1329);
or U3967 (N_3967,In_709,In_2154);
nor U3968 (N_3968,In_2368,In_276);
nor U3969 (N_3969,In_27,In_1477);
and U3970 (N_3970,In_2751,In_1140);
or U3971 (N_3971,In_1874,In_1749);
or U3972 (N_3972,In_476,In_233);
or U3973 (N_3973,In_1600,In_681);
nand U3974 (N_3974,In_313,In_895);
nor U3975 (N_3975,In_1359,In_417);
xor U3976 (N_3976,In_937,In_2207);
or U3977 (N_3977,In_1650,In_1046);
nor U3978 (N_3978,In_990,In_1655);
xnor U3979 (N_3979,In_2001,In_2277);
nand U3980 (N_3980,In_2835,In_1653);
or U3981 (N_3981,In_1139,In_1514);
and U3982 (N_3982,In_1062,In_2843);
xnor U3983 (N_3983,In_3,In_1315);
or U3984 (N_3984,In_2767,In_2530);
and U3985 (N_3985,In_1245,In_819);
and U3986 (N_3986,In_2670,In_1435);
and U3987 (N_3987,In_2374,In_1188);
nor U3988 (N_3988,In_515,In_261);
nor U3989 (N_3989,In_998,In_1313);
or U3990 (N_3990,In_32,In_484);
and U3991 (N_3991,In_2186,In_2443);
nor U3992 (N_3992,In_1219,In_820);
nand U3993 (N_3993,In_2385,In_172);
nor U3994 (N_3994,In_1921,In_991);
and U3995 (N_3995,In_893,In_269);
nor U3996 (N_3996,In_1999,In_2825);
xor U3997 (N_3997,In_189,In_251);
xnor U3998 (N_3998,In_269,In_2062);
nand U3999 (N_3999,In_2081,In_2548);
nand U4000 (N_4000,In_1386,In_708);
or U4001 (N_4001,In_2717,In_1602);
xor U4002 (N_4002,In_316,In_1895);
nor U4003 (N_4003,In_1604,In_1448);
and U4004 (N_4004,In_2348,In_223);
or U4005 (N_4005,In_774,In_1655);
or U4006 (N_4006,In_1376,In_2856);
or U4007 (N_4007,In_1753,In_1708);
and U4008 (N_4008,In_2597,In_2585);
and U4009 (N_4009,In_1292,In_206);
xnor U4010 (N_4010,In_2623,In_953);
nor U4011 (N_4011,In_627,In_2234);
nor U4012 (N_4012,In_2534,In_2086);
xor U4013 (N_4013,In_1585,In_2197);
or U4014 (N_4014,In_1831,In_1584);
and U4015 (N_4015,In_802,In_1282);
or U4016 (N_4016,In_2415,In_2981);
nor U4017 (N_4017,In_1424,In_356);
or U4018 (N_4018,In_1805,In_85);
nand U4019 (N_4019,In_2512,In_2963);
or U4020 (N_4020,In_1261,In_1432);
nand U4021 (N_4021,In_2308,In_942);
nor U4022 (N_4022,In_688,In_964);
and U4023 (N_4023,In_249,In_2171);
nand U4024 (N_4024,In_2454,In_585);
nor U4025 (N_4025,In_1047,In_2623);
nand U4026 (N_4026,In_2476,In_1927);
nand U4027 (N_4027,In_1325,In_2502);
and U4028 (N_4028,In_947,In_267);
xnor U4029 (N_4029,In_2937,In_2812);
nor U4030 (N_4030,In_1852,In_2821);
nand U4031 (N_4031,In_2873,In_2255);
and U4032 (N_4032,In_1913,In_989);
nand U4033 (N_4033,In_1856,In_1182);
and U4034 (N_4034,In_332,In_70);
or U4035 (N_4035,In_1603,In_363);
or U4036 (N_4036,In_449,In_1371);
xnor U4037 (N_4037,In_416,In_1159);
and U4038 (N_4038,In_1632,In_2670);
nor U4039 (N_4039,In_431,In_2985);
nor U4040 (N_4040,In_984,In_885);
nand U4041 (N_4041,In_33,In_1915);
xnor U4042 (N_4042,In_1877,In_2257);
and U4043 (N_4043,In_1484,In_63);
xor U4044 (N_4044,In_528,In_1368);
and U4045 (N_4045,In_1432,In_713);
xnor U4046 (N_4046,In_2071,In_1786);
nor U4047 (N_4047,In_2646,In_2347);
xor U4048 (N_4048,In_1162,In_1160);
nor U4049 (N_4049,In_1566,In_2948);
nand U4050 (N_4050,In_447,In_665);
and U4051 (N_4051,In_1409,In_1578);
nor U4052 (N_4052,In_289,In_1611);
nor U4053 (N_4053,In_637,In_2763);
or U4054 (N_4054,In_1337,In_1726);
xor U4055 (N_4055,In_2361,In_1205);
xnor U4056 (N_4056,In_1492,In_1060);
and U4057 (N_4057,In_1469,In_2364);
and U4058 (N_4058,In_573,In_2008);
xor U4059 (N_4059,In_1025,In_1069);
or U4060 (N_4060,In_1451,In_1232);
or U4061 (N_4061,In_755,In_1586);
xor U4062 (N_4062,In_419,In_2348);
and U4063 (N_4063,In_2331,In_923);
or U4064 (N_4064,In_524,In_496);
nor U4065 (N_4065,In_959,In_2757);
or U4066 (N_4066,In_1803,In_1720);
nor U4067 (N_4067,In_325,In_960);
xor U4068 (N_4068,In_2403,In_2770);
xnor U4069 (N_4069,In_734,In_2918);
xnor U4070 (N_4070,In_704,In_2497);
nand U4071 (N_4071,In_863,In_2214);
and U4072 (N_4072,In_2529,In_774);
nor U4073 (N_4073,In_627,In_1237);
and U4074 (N_4074,In_1235,In_220);
nor U4075 (N_4075,In_1975,In_1117);
nand U4076 (N_4076,In_628,In_1782);
xnor U4077 (N_4077,In_2549,In_2566);
xor U4078 (N_4078,In_1864,In_2995);
nor U4079 (N_4079,In_2041,In_1397);
nand U4080 (N_4080,In_1590,In_484);
nand U4081 (N_4081,In_2396,In_540);
nand U4082 (N_4082,In_2844,In_408);
xnor U4083 (N_4083,In_1038,In_1180);
nand U4084 (N_4084,In_175,In_1197);
xnor U4085 (N_4085,In_1559,In_2470);
and U4086 (N_4086,In_2253,In_2783);
or U4087 (N_4087,In_2602,In_2596);
nor U4088 (N_4088,In_2118,In_1322);
nand U4089 (N_4089,In_187,In_1453);
or U4090 (N_4090,In_1608,In_1550);
xor U4091 (N_4091,In_941,In_2721);
or U4092 (N_4092,In_2169,In_1904);
and U4093 (N_4093,In_1240,In_1951);
nor U4094 (N_4094,In_788,In_706);
xnor U4095 (N_4095,In_606,In_2631);
nand U4096 (N_4096,In_2059,In_2027);
nand U4097 (N_4097,In_525,In_1765);
nor U4098 (N_4098,In_1165,In_1847);
xnor U4099 (N_4099,In_937,In_2768);
xor U4100 (N_4100,In_1722,In_2245);
or U4101 (N_4101,In_2337,In_569);
and U4102 (N_4102,In_1142,In_1383);
xor U4103 (N_4103,In_2224,In_2931);
nand U4104 (N_4104,In_1932,In_1256);
or U4105 (N_4105,In_1302,In_2979);
xnor U4106 (N_4106,In_1363,In_2619);
nand U4107 (N_4107,In_2589,In_459);
or U4108 (N_4108,In_2999,In_420);
and U4109 (N_4109,In_1708,In_605);
nand U4110 (N_4110,In_68,In_1920);
and U4111 (N_4111,In_1960,In_1443);
xor U4112 (N_4112,In_1393,In_637);
nor U4113 (N_4113,In_2636,In_2069);
nand U4114 (N_4114,In_2175,In_1461);
xor U4115 (N_4115,In_2133,In_1649);
and U4116 (N_4116,In_1969,In_780);
nand U4117 (N_4117,In_2477,In_2641);
and U4118 (N_4118,In_1867,In_1024);
or U4119 (N_4119,In_2242,In_1997);
xnor U4120 (N_4120,In_2047,In_2599);
and U4121 (N_4121,In_627,In_122);
and U4122 (N_4122,In_360,In_212);
nand U4123 (N_4123,In_1627,In_3);
xor U4124 (N_4124,In_2825,In_2231);
nand U4125 (N_4125,In_2165,In_77);
nor U4126 (N_4126,In_2283,In_510);
nor U4127 (N_4127,In_323,In_181);
nand U4128 (N_4128,In_1946,In_2620);
and U4129 (N_4129,In_2906,In_1158);
nor U4130 (N_4130,In_1173,In_1230);
or U4131 (N_4131,In_2231,In_347);
or U4132 (N_4132,In_695,In_2564);
nor U4133 (N_4133,In_1691,In_2352);
and U4134 (N_4134,In_1599,In_1166);
nor U4135 (N_4135,In_2915,In_731);
xor U4136 (N_4136,In_1223,In_1712);
or U4137 (N_4137,In_444,In_2015);
nand U4138 (N_4138,In_2986,In_806);
nor U4139 (N_4139,In_2811,In_2798);
or U4140 (N_4140,In_1045,In_2540);
and U4141 (N_4141,In_2831,In_1178);
and U4142 (N_4142,In_2273,In_446);
and U4143 (N_4143,In_1516,In_979);
nor U4144 (N_4144,In_1491,In_750);
nor U4145 (N_4145,In_2670,In_713);
and U4146 (N_4146,In_120,In_2192);
nand U4147 (N_4147,In_2414,In_2967);
nand U4148 (N_4148,In_931,In_2452);
xnor U4149 (N_4149,In_2341,In_1730);
xnor U4150 (N_4150,In_1877,In_952);
nor U4151 (N_4151,In_1890,In_484);
or U4152 (N_4152,In_66,In_1777);
xor U4153 (N_4153,In_321,In_1455);
xnor U4154 (N_4154,In_1390,In_2777);
nor U4155 (N_4155,In_700,In_2654);
nor U4156 (N_4156,In_1145,In_1237);
or U4157 (N_4157,In_2833,In_2503);
and U4158 (N_4158,In_248,In_2596);
nand U4159 (N_4159,In_1265,In_630);
or U4160 (N_4160,In_1243,In_2204);
or U4161 (N_4161,In_518,In_2647);
nor U4162 (N_4162,In_2660,In_2346);
and U4163 (N_4163,In_615,In_1417);
xor U4164 (N_4164,In_2864,In_750);
nand U4165 (N_4165,In_2843,In_2111);
nor U4166 (N_4166,In_2287,In_2580);
nor U4167 (N_4167,In_2288,In_1405);
or U4168 (N_4168,In_1038,In_986);
nand U4169 (N_4169,In_2368,In_947);
nand U4170 (N_4170,In_2312,In_1731);
and U4171 (N_4171,In_217,In_1131);
or U4172 (N_4172,In_1952,In_1273);
nand U4173 (N_4173,In_2572,In_1472);
xor U4174 (N_4174,In_1029,In_1794);
nand U4175 (N_4175,In_1905,In_1891);
or U4176 (N_4176,In_463,In_595);
nand U4177 (N_4177,In_494,In_2095);
nand U4178 (N_4178,In_2647,In_1201);
nor U4179 (N_4179,In_2412,In_191);
and U4180 (N_4180,In_36,In_2237);
or U4181 (N_4181,In_2196,In_1220);
xor U4182 (N_4182,In_1234,In_797);
nor U4183 (N_4183,In_1153,In_2775);
and U4184 (N_4184,In_989,In_1130);
and U4185 (N_4185,In_2969,In_1436);
nor U4186 (N_4186,In_2189,In_142);
nand U4187 (N_4187,In_1204,In_2223);
xor U4188 (N_4188,In_1211,In_2546);
nor U4189 (N_4189,In_150,In_1008);
nand U4190 (N_4190,In_311,In_437);
and U4191 (N_4191,In_1733,In_2534);
nand U4192 (N_4192,In_775,In_1404);
or U4193 (N_4193,In_1570,In_2203);
nand U4194 (N_4194,In_1628,In_1480);
nand U4195 (N_4195,In_1246,In_885);
nand U4196 (N_4196,In_158,In_1677);
and U4197 (N_4197,In_809,In_2235);
and U4198 (N_4198,In_2781,In_737);
and U4199 (N_4199,In_1633,In_2013);
nor U4200 (N_4200,In_594,In_2659);
nor U4201 (N_4201,In_2730,In_2700);
or U4202 (N_4202,In_1917,In_1418);
and U4203 (N_4203,In_1247,In_454);
nor U4204 (N_4204,In_1920,In_2904);
and U4205 (N_4205,In_1997,In_901);
xor U4206 (N_4206,In_2342,In_2366);
xnor U4207 (N_4207,In_1889,In_49);
nand U4208 (N_4208,In_149,In_675);
xor U4209 (N_4209,In_2905,In_1440);
and U4210 (N_4210,In_1193,In_1865);
nor U4211 (N_4211,In_1129,In_1623);
and U4212 (N_4212,In_536,In_2832);
or U4213 (N_4213,In_720,In_11);
and U4214 (N_4214,In_1364,In_1242);
and U4215 (N_4215,In_2635,In_1016);
and U4216 (N_4216,In_1485,In_2611);
nor U4217 (N_4217,In_2378,In_1010);
or U4218 (N_4218,In_2276,In_990);
and U4219 (N_4219,In_520,In_2624);
and U4220 (N_4220,In_2981,In_2762);
and U4221 (N_4221,In_2924,In_2512);
or U4222 (N_4222,In_826,In_883);
nand U4223 (N_4223,In_2939,In_1891);
xnor U4224 (N_4224,In_2978,In_1426);
nor U4225 (N_4225,In_537,In_1183);
and U4226 (N_4226,In_184,In_100);
nand U4227 (N_4227,In_1350,In_1279);
nand U4228 (N_4228,In_2124,In_1287);
or U4229 (N_4229,In_735,In_1907);
or U4230 (N_4230,In_465,In_2500);
or U4231 (N_4231,In_2050,In_2537);
or U4232 (N_4232,In_1170,In_537);
or U4233 (N_4233,In_1830,In_1913);
and U4234 (N_4234,In_68,In_1304);
and U4235 (N_4235,In_2634,In_2147);
xnor U4236 (N_4236,In_2161,In_804);
or U4237 (N_4237,In_2599,In_471);
and U4238 (N_4238,In_759,In_2542);
nand U4239 (N_4239,In_2906,In_2381);
and U4240 (N_4240,In_2345,In_144);
nor U4241 (N_4241,In_2450,In_451);
and U4242 (N_4242,In_2737,In_1353);
or U4243 (N_4243,In_829,In_833);
xor U4244 (N_4244,In_191,In_2309);
nor U4245 (N_4245,In_2690,In_2724);
nor U4246 (N_4246,In_293,In_2726);
nor U4247 (N_4247,In_1859,In_2904);
and U4248 (N_4248,In_1583,In_1137);
xor U4249 (N_4249,In_1900,In_1964);
nand U4250 (N_4250,In_1871,In_2855);
xnor U4251 (N_4251,In_944,In_22);
xnor U4252 (N_4252,In_158,In_109);
or U4253 (N_4253,In_1366,In_34);
nand U4254 (N_4254,In_2504,In_2825);
or U4255 (N_4255,In_1223,In_772);
nand U4256 (N_4256,In_2782,In_299);
xor U4257 (N_4257,In_1010,In_107);
xnor U4258 (N_4258,In_1548,In_2341);
nor U4259 (N_4259,In_459,In_1260);
nor U4260 (N_4260,In_2408,In_1634);
nor U4261 (N_4261,In_2086,In_2694);
nand U4262 (N_4262,In_2623,In_2435);
and U4263 (N_4263,In_2471,In_1859);
xnor U4264 (N_4264,In_1430,In_970);
xor U4265 (N_4265,In_2047,In_2424);
or U4266 (N_4266,In_235,In_2119);
nor U4267 (N_4267,In_817,In_1881);
nor U4268 (N_4268,In_446,In_2643);
nand U4269 (N_4269,In_1658,In_945);
nand U4270 (N_4270,In_2834,In_1031);
nor U4271 (N_4271,In_1556,In_2315);
or U4272 (N_4272,In_1971,In_564);
or U4273 (N_4273,In_2872,In_2434);
or U4274 (N_4274,In_2848,In_1156);
nand U4275 (N_4275,In_999,In_1567);
nand U4276 (N_4276,In_918,In_205);
xor U4277 (N_4277,In_2094,In_2512);
nor U4278 (N_4278,In_1907,In_981);
nand U4279 (N_4279,In_1683,In_903);
nand U4280 (N_4280,In_2007,In_699);
and U4281 (N_4281,In_716,In_611);
nand U4282 (N_4282,In_1102,In_616);
and U4283 (N_4283,In_1188,In_2234);
xnor U4284 (N_4284,In_1984,In_1111);
or U4285 (N_4285,In_854,In_149);
and U4286 (N_4286,In_27,In_2755);
xnor U4287 (N_4287,In_1032,In_2819);
and U4288 (N_4288,In_2815,In_2859);
or U4289 (N_4289,In_1282,In_763);
xor U4290 (N_4290,In_10,In_1961);
nand U4291 (N_4291,In_1346,In_2659);
nand U4292 (N_4292,In_327,In_48);
or U4293 (N_4293,In_1183,In_1790);
nor U4294 (N_4294,In_1052,In_2984);
and U4295 (N_4295,In_1293,In_222);
and U4296 (N_4296,In_1416,In_48);
nor U4297 (N_4297,In_1579,In_1488);
or U4298 (N_4298,In_733,In_2123);
and U4299 (N_4299,In_1356,In_371);
and U4300 (N_4300,In_2687,In_1584);
nor U4301 (N_4301,In_1033,In_1784);
nor U4302 (N_4302,In_964,In_2247);
xnor U4303 (N_4303,In_71,In_213);
xor U4304 (N_4304,In_811,In_2644);
or U4305 (N_4305,In_273,In_964);
nand U4306 (N_4306,In_415,In_973);
and U4307 (N_4307,In_1643,In_20);
xnor U4308 (N_4308,In_2932,In_1498);
nand U4309 (N_4309,In_2609,In_892);
nand U4310 (N_4310,In_1473,In_1941);
nor U4311 (N_4311,In_2720,In_973);
xor U4312 (N_4312,In_938,In_2593);
xnor U4313 (N_4313,In_1900,In_1189);
nor U4314 (N_4314,In_1858,In_938);
nor U4315 (N_4315,In_254,In_271);
or U4316 (N_4316,In_165,In_97);
xor U4317 (N_4317,In_2402,In_2129);
or U4318 (N_4318,In_311,In_1667);
xnor U4319 (N_4319,In_1426,In_300);
nor U4320 (N_4320,In_766,In_2137);
or U4321 (N_4321,In_1524,In_2113);
nand U4322 (N_4322,In_2047,In_1791);
xnor U4323 (N_4323,In_391,In_1357);
nor U4324 (N_4324,In_2256,In_203);
nand U4325 (N_4325,In_1098,In_852);
nand U4326 (N_4326,In_2999,In_224);
nand U4327 (N_4327,In_884,In_1890);
xor U4328 (N_4328,In_226,In_1250);
or U4329 (N_4329,In_2851,In_1965);
or U4330 (N_4330,In_2322,In_193);
nand U4331 (N_4331,In_2416,In_584);
or U4332 (N_4332,In_184,In_2509);
or U4333 (N_4333,In_782,In_2706);
nor U4334 (N_4334,In_1572,In_1746);
xor U4335 (N_4335,In_1250,In_240);
nor U4336 (N_4336,In_1357,In_693);
or U4337 (N_4337,In_2060,In_1396);
and U4338 (N_4338,In_1167,In_982);
nor U4339 (N_4339,In_1272,In_1379);
and U4340 (N_4340,In_1245,In_2936);
and U4341 (N_4341,In_22,In_893);
or U4342 (N_4342,In_500,In_581);
nor U4343 (N_4343,In_106,In_1798);
and U4344 (N_4344,In_1231,In_2942);
or U4345 (N_4345,In_183,In_1420);
xor U4346 (N_4346,In_664,In_2516);
or U4347 (N_4347,In_1471,In_2413);
or U4348 (N_4348,In_1165,In_1684);
xnor U4349 (N_4349,In_743,In_2844);
nor U4350 (N_4350,In_2088,In_2089);
xor U4351 (N_4351,In_2665,In_1584);
or U4352 (N_4352,In_1511,In_1803);
nor U4353 (N_4353,In_537,In_2574);
and U4354 (N_4354,In_936,In_1845);
nor U4355 (N_4355,In_2002,In_1639);
nor U4356 (N_4356,In_2782,In_2768);
nand U4357 (N_4357,In_1756,In_2522);
nand U4358 (N_4358,In_2329,In_1868);
or U4359 (N_4359,In_1849,In_1033);
and U4360 (N_4360,In_2301,In_2155);
or U4361 (N_4361,In_2737,In_138);
and U4362 (N_4362,In_1880,In_342);
or U4363 (N_4363,In_2120,In_977);
nor U4364 (N_4364,In_924,In_2728);
and U4365 (N_4365,In_590,In_1881);
nand U4366 (N_4366,In_1027,In_1547);
or U4367 (N_4367,In_1863,In_1096);
or U4368 (N_4368,In_738,In_1011);
xor U4369 (N_4369,In_2585,In_980);
nand U4370 (N_4370,In_691,In_2207);
nor U4371 (N_4371,In_554,In_177);
or U4372 (N_4372,In_2526,In_2);
nand U4373 (N_4373,In_1486,In_512);
or U4374 (N_4374,In_2362,In_2027);
xor U4375 (N_4375,In_76,In_2075);
nand U4376 (N_4376,In_2129,In_2811);
and U4377 (N_4377,In_1036,In_1917);
nand U4378 (N_4378,In_1150,In_181);
and U4379 (N_4379,In_215,In_2302);
and U4380 (N_4380,In_1740,In_1561);
nand U4381 (N_4381,In_300,In_1143);
nor U4382 (N_4382,In_821,In_1329);
xor U4383 (N_4383,In_2994,In_1014);
nor U4384 (N_4384,In_1936,In_2207);
xor U4385 (N_4385,In_414,In_1631);
or U4386 (N_4386,In_906,In_189);
or U4387 (N_4387,In_2591,In_694);
xor U4388 (N_4388,In_2176,In_2186);
and U4389 (N_4389,In_1571,In_2699);
xor U4390 (N_4390,In_1211,In_2647);
nor U4391 (N_4391,In_2959,In_759);
nor U4392 (N_4392,In_1981,In_2754);
xnor U4393 (N_4393,In_1617,In_1818);
nand U4394 (N_4394,In_2694,In_274);
nor U4395 (N_4395,In_1896,In_2501);
xor U4396 (N_4396,In_2191,In_2791);
nor U4397 (N_4397,In_2051,In_1058);
and U4398 (N_4398,In_1660,In_2680);
nand U4399 (N_4399,In_2065,In_1945);
or U4400 (N_4400,In_1346,In_547);
xor U4401 (N_4401,In_1003,In_530);
nor U4402 (N_4402,In_1370,In_1207);
nand U4403 (N_4403,In_2211,In_1218);
and U4404 (N_4404,In_14,In_2718);
and U4405 (N_4405,In_1342,In_1102);
nand U4406 (N_4406,In_891,In_1898);
xor U4407 (N_4407,In_2916,In_1408);
or U4408 (N_4408,In_1913,In_2830);
nand U4409 (N_4409,In_2009,In_2799);
or U4410 (N_4410,In_1670,In_2125);
and U4411 (N_4411,In_274,In_2477);
xor U4412 (N_4412,In_1699,In_2149);
xnor U4413 (N_4413,In_456,In_2559);
and U4414 (N_4414,In_2097,In_2242);
xor U4415 (N_4415,In_2779,In_132);
and U4416 (N_4416,In_733,In_2991);
nor U4417 (N_4417,In_1405,In_1635);
xor U4418 (N_4418,In_57,In_1587);
xor U4419 (N_4419,In_2300,In_1318);
nand U4420 (N_4420,In_1534,In_38);
and U4421 (N_4421,In_951,In_2492);
xnor U4422 (N_4422,In_2035,In_1743);
or U4423 (N_4423,In_620,In_2884);
nor U4424 (N_4424,In_2155,In_1046);
nor U4425 (N_4425,In_1221,In_197);
nand U4426 (N_4426,In_1256,In_2004);
xnor U4427 (N_4427,In_495,In_686);
nor U4428 (N_4428,In_106,In_2825);
and U4429 (N_4429,In_1680,In_2998);
or U4430 (N_4430,In_2795,In_448);
nand U4431 (N_4431,In_54,In_2322);
nand U4432 (N_4432,In_2553,In_2423);
or U4433 (N_4433,In_2941,In_1694);
xnor U4434 (N_4434,In_1750,In_148);
nand U4435 (N_4435,In_493,In_618);
or U4436 (N_4436,In_167,In_2995);
nand U4437 (N_4437,In_461,In_496);
xnor U4438 (N_4438,In_249,In_703);
or U4439 (N_4439,In_469,In_1471);
and U4440 (N_4440,In_2455,In_186);
or U4441 (N_4441,In_1868,In_1471);
xnor U4442 (N_4442,In_1247,In_935);
and U4443 (N_4443,In_2132,In_1866);
and U4444 (N_4444,In_1452,In_2265);
xnor U4445 (N_4445,In_2769,In_1781);
nor U4446 (N_4446,In_2341,In_805);
and U4447 (N_4447,In_998,In_2657);
or U4448 (N_4448,In_2054,In_2930);
or U4449 (N_4449,In_796,In_2230);
and U4450 (N_4450,In_1678,In_2489);
or U4451 (N_4451,In_956,In_1859);
xor U4452 (N_4452,In_187,In_176);
nand U4453 (N_4453,In_1931,In_1661);
xor U4454 (N_4454,In_818,In_414);
nor U4455 (N_4455,In_2950,In_241);
nor U4456 (N_4456,In_2312,In_1031);
or U4457 (N_4457,In_2101,In_224);
nor U4458 (N_4458,In_2857,In_527);
nor U4459 (N_4459,In_1652,In_1997);
nor U4460 (N_4460,In_1605,In_807);
nor U4461 (N_4461,In_2030,In_2850);
nand U4462 (N_4462,In_2745,In_1876);
xor U4463 (N_4463,In_1982,In_873);
nand U4464 (N_4464,In_2804,In_2661);
and U4465 (N_4465,In_1613,In_1202);
xnor U4466 (N_4466,In_1313,In_988);
and U4467 (N_4467,In_2252,In_1452);
nand U4468 (N_4468,In_2854,In_2529);
or U4469 (N_4469,In_1986,In_1003);
nor U4470 (N_4470,In_2424,In_220);
xnor U4471 (N_4471,In_1082,In_2614);
xor U4472 (N_4472,In_2157,In_1678);
nand U4473 (N_4473,In_207,In_554);
or U4474 (N_4474,In_629,In_2303);
xnor U4475 (N_4475,In_475,In_1103);
nor U4476 (N_4476,In_2382,In_842);
nand U4477 (N_4477,In_32,In_1777);
or U4478 (N_4478,In_2644,In_1780);
nand U4479 (N_4479,In_1084,In_2987);
nor U4480 (N_4480,In_1624,In_1328);
and U4481 (N_4481,In_2730,In_1502);
xor U4482 (N_4482,In_179,In_2251);
or U4483 (N_4483,In_1028,In_1545);
nor U4484 (N_4484,In_2955,In_2727);
or U4485 (N_4485,In_2642,In_1391);
or U4486 (N_4486,In_607,In_2934);
and U4487 (N_4487,In_2161,In_2970);
or U4488 (N_4488,In_512,In_2284);
nand U4489 (N_4489,In_297,In_1719);
nor U4490 (N_4490,In_1639,In_1715);
nand U4491 (N_4491,In_2537,In_302);
nor U4492 (N_4492,In_1371,In_1698);
nand U4493 (N_4493,In_1399,In_984);
and U4494 (N_4494,In_1114,In_2547);
or U4495 (N_4495,In_2733,In_758);
and U4496 (N_4496,In_712,In_2624);
nor U4497 (N_4497,In_2203,In_981);
nand U4498 (N_4498,In_1007,In_2442);
nand U4499 (N_4499,In_1163,In_2994);
nor U4500 (N_4500,In_2924,In_2238);
nor U4501 (N_4501,In_2076,In_1506);
or U4502 (N_4502,In_2340,In_1379);
xor U4503 (N_4503,In_2770,In_339);
nand U4504 (N_4504,In_133,In_2115);
or U4505 (N_4505,In_1023,In_2333);
and U4506 (N_4506,In_2776,In_1928);
or U4507 (N_4507,In_2699,In_743);
and U4508 (N_4508,In_309,In_57);
nand U4509 (N_4509,In_2816,In_2874);
xor U4510 (N_4510,In_295,In_1388);
nor U4511 (N_4511,In_1809,In_1317);
nor U4512 (N_4512,In_1273,In_1591);
nand U4513 (N_4513,In_1595,In_132);
xor U4514 (N_4514,In_1286,In_457);
and U4515 (N_4515,In_1528,In_1399);
xnor U4516 (N_4516,In_403,In_942);
nor U4517 (N_4517,In_1886,In_596);
or U4518 (N_4518,In_1310,In_851);
xor U4519 (N_4519,In_885,In_1187);
nor U4520 (N_4520,In_305,In_1170);
xnor U4521 (N_4521,In_576,In_1566);
and U4522 (N_4522,In_2149,In_957);
and U4523 (N_4523,In_1277,In_1466);
and U4524 (N_4524,In_1191,In_1590);
nand U4525 (N_4525,In_1244,In_2722);
and U4526 (N_4526,In_308,In_691);
nand U4527 (N_4527,In_1516,In_1788);
and U4528 (N_4528,In_1734,In_2201);
nand U4529 (N_4529,In_1939,In_428);
nand U4530 (N_4530,In_1266,In_1772);
nor U4531 (N_4531,In_2807,In_1373);
and U4532 (N_4532,In_2166,In_1718);
or U4533 (N_4533,In_137,In_1416);
xnor U4534 (N_4534,In_801,In_2812);
and U4535 (N_4535,In_2037,In_2812);
nand U4536 (N_4536,In_1157,In_1409);
nor U4537 (N_4537,In_2494,In_2184);
and U4538 (N_4538,In_996,In_2599);
or U4539 (N_4539,In_1292,In_474);
nand U4540 (N_4540,In_1313,In_2791);
nand U4541 (N_4541,In_535,In_530);
nand U4542 (N_4542,In_1308,In_202);
nor U4543 (N_4543,In_1524,In_2101);
or U4544 (N_4544,In_2413,In_2127);
xnor U4545 (N_4545,In_1728,In_154);
or U4546 (N_4546,In_1826,In_2660);
nor U4547 (N_4547,In_1479,In_2484);
and U4548 (N_4548,In_2942,In_926);
xor U4549 (N_4549,In_217,In_837);
nand U4550 (N_4550,In_882,In_1037);
and U4551 (N_4551,In_862,In_644);
or U4552 (N_4552,In_1758,In_1844);
or U4553 (N_4553,In_2775,In_1930);
or U4554 (N_4554,In_1389,In_190);
xnor U4555 (N_4555,In_622,In_860);
nand U4556 (N_4556,In_1138,In_1679);
or U4557 (N_4557,In_1035,In_2600);
and U4558 (N_4558,In_965,In_2177);
nor U4559 (N_4559,In_525,In_70);
nor U4560 (N_4560,In_1147,In_1252);
xnor U4561 (N_4561,In_2506,In_827);
xnor U4562 (N_4562,In_612,In_1088);
xnor U4563 (N_4563,In_1142,In_2121);
nand U4564 (N_4564,In_1961,In_1553);
or U4565 (N_4565,In_37,In_675);
or U4566 (N_4566,In_1282,In_1046);
xnor U4567 (N_4567,In_2007,In_2765);
nor U4568 (N_4568,In_246,In_1440);
and U4569 (N_4569,In_2645,In_2759);
xnor U4570 (N_4570,In_1050,In_2258);
nor U4571 (N_4571,In_2663,In_1117);
nor U4572 (N_4572,In_676,In_1355);
or U4573 (N_4573,In_2454,In_1705);
or U4574 (N_4574,In_990,In_1367);
nand U4575 (N_4575,In_1903,In_2350);
and U4576 (N_4576,In_944,In_371);
nor U4577 (N_4577,In_1175,In_2172);
or U4578 (N_4578,In_297,In_1736);
nor U4579 (N_4579,In_787,In_2771);
or U4580 (N_4580,In_209,In_2678);
xor U4581 (N_4581,In_756,In_2408);
and U4582 (N_4582,In_411,In_1350);
nand U4583 (N_4583,In_1789,In_1804);
nand U4584 (N_4584,In_400,In_1888);
nor U4585 (N_4585,In_683,In_2385);
nor U4586 (N_4586,In_175,In_1939);
or U4587 (N_4587,In_302,In_284);
or U4588 (N_4588,In_2432,In_781);
nor U4589 (N_4589,In_1802,In_743);
nand U4590 (N_4590,In_551,In_1989);
or U4591 (N_4591,In_2900,In_2193);
and U4592 (N_4592,In_2179,In_2321);
xnor U4593 (N_4593,In_530,In_851);
xor U4594 (N_4594,In_840,In_2755);
nor U4595 (N_4595,In_649,In_1784);
and U4596 (N_4596,In_1165,In_1647);
nand U4597 (N_4597,In_2702,In_193);
or U4598 (N_4598,In_1329,In_919);
nand U4599 (N_4599,In_2973,In_632);
and U4600 (N_4600,In_2374,In_1819);
nor U4601 (N_4601,In_2723,In_483);
nor U4602 (N_4602,In_2863,In_547);
and U4603 (N_4603,In_398,In_966);
nor U4604 (N_4604,In_1629,In_1943);
and U4605 (N_4605,In_2585,In_2887);
nand U4606 (N_4606,In_1420,In_2649);
and U4607 (N_4607,In_2473,In_420);
nand U4608 (N_4608,In_227,In_632);
nor U4609 (N_4609,In_1594,In_1810);
and U4610 (N_4610,In_491,In_972);
and U4611 (N_4611,In_1835,In_1487);
xnor U4612 (N_4612,In_206,In_1464);
nor U4613 (N_4613,In_1434,In_1764);
xor U4614 (N_4614,In_900,In_2964);
nand U4615 (N_4615,In_2146,In_2763);
and U4616 (N_4616,In_1791,In_782);
xnor U4617 (N_4617,In_757,In_1563);
xnor U4618 (N_4618,In_2611,In_1907);
xor U4619 (N_4619,In_718,In_2061);
nor U4620 (N_4620,In_1555,In_1341);
or U4621 (N_4621,In_1816,In_734);
xor U4622 (N_4622,In_346,In_2347);
xnor U4623 (N_4623,In_1442,In_800);
or U4624 (N_4624,In_123,In_494);
nand U4625 (N_4625,In_2594,In_836);
and U4626 (N_4626,In_850,In_979);
nand U4627 (N_4627,In_1322,In_2305);
or U4628 (N_4628,In_2096,In_2296);
nand U4629 (N_4629,In_2566,In_1226);
nor U4630 (N_4630,In_679,In_122);
xor U4631 (N_4631,In_1453,In_154);
xor U4632 (N_4632,In_1833,In_2182);
nor U4633 (N_4633,In_2688,In_2066);
nor U4634 (N_4634,In_430,In_332);
nor U4635 (N_4635,In_194,In_2550);
nor U4636 (N_4636,In_752,In_1780);
xnor U4637 (N_4637,In_2171,In_848);
nand U4638 (N_4638,In_1742,In_2473);
xnor U4639 (N_4639,In_2876,In_1948);
or U4640 (N_4640,In_1734,In_412);
xnor U4641 (N_4641,In_1506,In_438);
nor U4642 (N_4642,In_1489,In_2929);
nor U4643 (N_4643,In_1044,In_478);
nor U4644 (N_4644,In_1696,In_1300);
and U4645 (N_4645,In_1155,In_730);
nor U4646 (N_4646,In_2243,In_2892);
nand U4647 (N_4647,In_851,In_1337);
and U4648 (N_4648,In_741,In_1979);
xor U4649 (N_4649,In_2382,In_479);
or U4650 (N_4650,In_922,In_305);
nor U4651 (N_4651,In_168,In_2624);
xnor U4652 (N_4652,In_1356,In_1251);
or U4653 (N_4653,In_2198,In_1528);
nor U4654 (N_4654,In_245,In_1735);
nand U4655 (N_4655,In_1016,In_180);
and U4656 (N_4656,In_831,In_1340);
nand U4657 (N_4657,In_2352,In_2841);
nor U4658 (N_4658,In_133,In_2095);
xnor U4659 (N_4659,In_110,In_1964);
and U4660 (N_4660,In_1389,In_1047);
nor U4661 (N_4661,In_978,In_2842);
nor U4662 (N_4662,In_2814,In_1301);
or U4663 (N_4663,In_953,In_2271);
nor U4664 (N_4664,In_2836,In_203);
nand U4665 (N_4665,In_46,In_284);
nand U4666 (N_4666,In_1216,In_2509);
or U4667 (N_4667,In_2147,In_1997);
xor U4668 (N_4668,In_2304,In_986);
xnor U4669 (N_4669,In_2424,In_1613);
or U4670 (N_4670,In_1775,In_668);
nand U4671 (N_4671,In_2316,In_2124);
and U4672 (N_4672,In_2288,In_84);
xnor U4673 (N_4673,In_534,In_936);
nor U4674 (N_4674,In_1633,In_2082);
xor U4675 (N_4675,In_1941,In_2934);
or U4676 (N_4676,In_482,In_998);
xnor U4677 (N_4677,In_1732,In_89);
and U4678 (N_4678,In_2665,In_303);
and U4679 (N_4679,In_594,In_1284);
or U4680 (N_4680,In_2134,In_2979);
or U4681 (N_4681,In_2316,In_2143);
nor U4682 (N_4682,In_2965,In_1001);
nand U4683 (N_4683,In_2507,In_2675);
xnor U4684 (N_4684,In_1665,In_1411);
nand U4685 (N_4685,In_321,In_2280);
and U4686 (N_4686,In_2574,In_212);
nor U4687 (N_4687,In_1210,In_114);
or U4688 (N_4688,In_536,In_1548);
or U4689 (N_4689,In_2532,In_1540);
xor U4690 (N_4690,In_1850,In_2114);
or U4691 (N_4691,In_1772,In_394);
xor U4692 (N_4692,In_2274,In_2029);
nor U4693 (N_4693,In_1766,In_2215);
or U4694 (N_4694,In_1451,In_652);
xnor U4695 (N_4695,In_1307,In_433);
xnor U4696 (N_4696,In_975,In_2358);
or U4697 (N_4697,In_848,In_560);
nor U4698 (N_4698,In_1631,In_816);
xor U4699 (N_4699,In_223,In_1492);
xor U4700 (N_4700,In_713,In_61);
or U4701 (N_4701,In_2089,In_1818);
xor U4702 (N_4702,In_2377,In_2506);
nor U4703 (N_4703,In_1596,In_283);
and U4704 (N_4704,In_263,In_1720);
or U4705 (N_4705,In_1210,In_2245);
xnor U4706 (N_4706,In_1394,In_1413);
and U4707 (N_4707,In_1792,In_2271);
or U4708 (N_4708,In_2364,In_2105);
or U4709 (N_4709,In_2295,In_829);
and U4710 (N_4710,In_2441,In_92);
and U4711 (N_4711,In_1140,In_1532);
nor U4712 (N_4712,In_2066,In_1786);
nor U4713 (N_4713,In_1895,In_2153);
or U4714 (N_4714,In_341,In_1818);
xor U4715 (N_4715,In_2738,In_1256);
nor U4716 (N_4716,In_1578,In_698);
or U4717 (N_4717,In_680,In_804);
xor U4718 (N_4718,In_431,In_2781);
or U4719 (N_4719,In_2711,In_2994);
xor U4720 (N_4720,In_343,In_2443);
xor U4721 (N_4721,In_1787,In_1066);
xor U4722 (N_4722,In_674,In_1357);
and U4723 (N_4723,In_2206,In_1712);
nand U4724 (N_4724,In_467,In_607);
and U4725 (N_4725,In_231,In_2447);
and U4726 (N_4726,In_1362,In_449);
or U4727 (N_4727,In_2636,In_1240);
and U4728 (N_4728,In_2637,In_2651);
nand U4729 (N_4729,In_1676,In_1563);
nand U4730 (N_4730,In_281,In_835);
and U4731 (N_4731,In_265,In_2784);
xnor U4732 (N_4732,In_659,In_1561);
nor U4733 (N_4733,In_194,In_548);
xor U4734 (N_4734,In_2134,In_284);
xnor U4735 (N_4735,In_2143,In_2665);
nand U4736 (N_4736,In_1804,In_1753);
and U4737 (N_4737,In_1341,In_1950);
and U4738 (N_4738,In_177,In_2767);
or U4739 (N_4739,In_1666,In_275);
nor U4740 (N_4740,In_2179,In_949);
or U4741 (N_4741,In_1315,In_39);
and U4742 (N_4742,In_2789,In_1321);
nor U4743 (N_4743,In_1477,In_2524);
nor U4744 (N_4744,In_1831,In_2790);
and U4745 (N_4745,In_2304,In_2347);
xor U4746 (N_4746,In_2970,In_2243);
and U4747 (N_4747,In_2607,In_840);
nor U4748 (N_4748,In_396,In_912);
nand U4749 (N_4749,In_2044,In_445);
and U4750 (N_4750,In_548,In_2312);
nand U4751 (N_4751,In_2278,In_597);
xnor U4752 (N_4752,In_2693,In_849);
nor U4753 (N_4753,In_284,In_589);
nor U4754 (N_4754,In_699,In_2998);
nor U4755 (N_4755,In_2083,In_1746);
nand U4756 (N_4756,In_2407,In_2107);
xor U4757 (N_4757,In_346,In_1387);
nand U4758 (N_4758,In_152,In_1870);
nand U4759 (N_4759,In_1564,In_2613);
xor U4760 (N_4760,In_491,In_258);
and U4761 (N_4761,In_242,In_592);
xnor U4762 (N_4762,In_2340,In_1543);
nor U4763 (N_4763,In_2517,In_1582);
nor U4764 (N_4764,In_226,In_417);
xor U4765 (N_4765,In_1284,In_2820);
xor U4766 (N_4766,In_1944,In_276);
nand U4767 (N_4767,In_490,In_1755);
xor U4768 (N_4768,In_2388,In_2356);
nor U4769 (N_4769,In_1400,In_118);
nor U4770 (N_4770,In_1870,In_1455);
or U4771 (N_4771,In_2750,In_2652);
or U4772 (N_4772,In_586,In_2658);
or U4773 (N_4773,In_2106,In_728);
nand U4774 (N_4774,In_1580,In_999);
or U4775 (N_4775,In_242,In_949);
or U4776 (N_4776,In_1624,In_179);
xor U4777 (N_4777,In_580,In_1801);
nand U4778 (N_4778,In_2872,In_2809);
xor U4779 (N_4779,In_2835,In_1578);
and U4780 (N_4780,In_2176,In_752);
and U4781 (N_4781,In_2224,In_1980);
xnor U4782 (N_4782,In_1072,In_1163);
or U4783 (N_4783,In_1023,In_1938);
or U4784 (N_4784,In_2011,In_2498);
or U4785 (N_4785,In_782,In_2196);
xnor U4786 (N_4786,In_1222,In_1390);
and U4787 (N_4787,In_451,In_2643);
xnor U4788 (N_4788,In_570,In_2126);
nor U4789 (N_4789,In_2400,In_955);
xor U4790 (N_4790,In_1552,In_1095);
nor U4791 (N_4791,In_1752,In_2761);
and U4792 (N_4792,In_2834,In_424);
nor U4793 (N_4793,In_1847,In_1334);
and U4794 (N_4794,In_2084,In_1111);
xor U4795 (N_4795,In_804,In_2326);
or U4796 (N_4796,In_2704,In_1882);
or U4797 (N_4797,In_2089,In_865);
nor U4798 (N_4798,In_2007,In_906);
and U4799 (N_4799,In_1271,In_2239);
nand U4800 (N_4800,In_975,In_2866);
nor U4801 (N_4801,In_2237,In_638);
nand U4802 (N_4802,In_695,In_1227);
and U4803 (N_4803,In_791,In_2034);
nor U4804 (N_4804,In_2026,In_1199);
xnor U4805 (N_4805,In_136,In_1280);
nor U4806 (N_4806,In_2013,In_944);
xor U4807 (N_4807,In_798,In_368);
or U4808 (N_4808,In_1075,In_1736);
xor U4809 (N_4809,In_2747,In_2433);
nand U4810 (N_4810,In_893,In_366);
or U4811 (N_4811,In_577,In_2823);
nor U4812 (N_4812,In_1080,In_644);
and U4813 (N_4813,In_1465,In_2850);
nor U4814 (N_4814,In_978,In_145);
nor U4815 (N_4815,In_1909,In_2469);
and U4816 (N_4816,In_827,In_1260);
nand U4817 (N_4817,In_2274,In_2980);
nor U4818 (N_4818,In_1788,In_2843);
xor U4819 (N_4819,In_265,In_2707);
or U4820 (N_4820,In_331,In_2248);
nor U4821 (N_4821,In_1811,In_1065);
nand U4822 (N_4822,In_2018,In_440);
nor U4823 (N_4823,In_51,In_2385);
xor U4824 (N_4824,In_2004,In_1565);
or U4825 (N_4825,In_2837,In_2428);
and U4826 (N_4826,In_337,In_2096);
and U4827 (N_4827,In_2012,In_2043);
and U4828 (N_4828,In_67,In_2715);
xor U4829 (N_4829,In_2125,In_2737);
nand U4830 (N_4830,In_1302,In_245);
nand U4831 (N_4831,In_2840,In_1284);
nand U4832 (N_4832,In_269,In_2988);
or U4833 (N_4833,In_1202,In_213);
nand U4834 (N_4834,In_2223,In_1424);
xnor U4835 (N_4835,In_269,In_1738);
or U4836 (N_4836,In_2099,In_1584);
and U4837 (N_4837,In_2202,In_2950);
and U4838 (N_4838,In_853,In_631);
nand U4839 (N_4839,In_86,In_2943);
and U4840 (N_4840,In_962,In_649);
and U4841 (N_4841,In_260,In_716);
and U4842 (N_4842,In_1551,In_2060);
nor U4843 (N_4843,In_2071,In_2760);
or U4844 (N_4844,In_2427,In_2307);
and U4845 (N_4845,In_1581,In_2295);
xnor U4846 (N_4846,In_2796,In_2328);
and U4847 (N_4847,In_170,In_546);
nor U4848 (N_4848,In_2007,In_752);
xor U4849 (N_4849,In_771,In_1003);
and U4850 (N_4850,In_129,In_217);
xor U4851 (N_4851,In_2950,In_1280);
and U4852 (N_4852,In_2407,In_792);
or U4853 (N_4853,In_1998,In_1947);
nand U4854 (N_4854,In_230,In_2092);
or U4855 (N_4855,In_463,In_2750);
xnor U4856 (N_4856,In_1716,In_1926);
and U4857 (N_4857,In_1617,In_1793);
and U4858 (N_4858,In_1169,In_959);
and U4859 (N_4859,In_2705,In_2793);
nand U4860 (N_4860,In_235,In_1191);
nor U4861 (N_4861,In_231,In_2756);
xnor U4862 (N_4862,In_2003,In_1594);
or U4863 (N_4863,In_590,In_428);
and U4864 (N_4864,In_596,In_1971);
nand U4865 (N_4865,In_1279,In_605);
nand U4866 (N_4866,In_1867,In_364);
or U4867 (N_4867,In_65,In_1756);
and U4868 (N_4868,In_1020,In_2384);
or U4869 (N_4869,In_135,In_1126);
nor U4870 (N_4870,In_695,In_1812);
or U4871 (N_4871,In_449,In_2011);
nor U4872 (N_4872,In_2901,In_194);
or U4873 (N_4873,In_1523,In_1435);
nand U4874 (N_4874,In_2967,In_2216);
and U4875 (N_4875,In_1888,In_1512);
nor U4876 (N_4876,In_938,In_2888);
or U4877 (N_4877,In_1568,In_2928);
and U4878 (N_4878,In_2698,In_1808);
and U4879 (N_4879,In_1829,In_739);
or U4880 (N_4880,In_1378,In_2553);
and U4881 (N_4881,In_2414,In_2651);
or U4882 (N_4882,In_627,In_1745);
or U4883 (N_4883,In_300,In_2766);
nor U4884 (N_4884,In_1796,In_997);
nand U4885 (N_4885,In_1316,In_1573);
or U4886 (N_4886,In_2616,In_2411);
xor U4887 (N_4887,In_1194,In_1264);
nand U4888 (N_4888,In_296,In_1386);
or U4889 (N_4889,In_2799,In_697);
nand U4890 (N_4890,In_146,In_2262);
xor U4891 (N_4891,In_1585,In_618);
and U4892 (N_4892,In_930,In_158);
xnor U4893 (N_4893,In_2753,In_2215);
xor U4894 (N_4894,In_536,In_1152);
xnor U4895 (N_4895,In_1907,In_630);
or U4896 (N_4896,In_1195,In_1855);
nand U4897 (N_4897,In_2590,In_1382);
or U4898 (N_4898,In_2155,In_2679);
nand U4899 (N_4899,In_1085,In_2776);
or U4900 (N_4900,In_165,In_145);
nand U4901 (N_4901,In_2630,In_1178);
or U4902 (N_4902,In_368,In_2795);
nand U4903 (N_4903,In_2954,In_1237);
nand U4904 (N_4904,In_1597,In_2418);
and U4905 (N_4905,In_132,In_2648);
nand U4906 (N_4906,In_730,In_2263);
nor U4907 (N_4907,In_860,In_73);
or U4908 (N_4908,In_2047,In_127);
or U4909 (N_4909,In_2637,In_1332);
and U4910 (N_4910,In_91,In_2291);
or U4911 (N_4911,In_1224,In_2159);
or U4912 (N_4912,In_2043,In_1515);
nand U4913 (N_4913,In_2604,In_1320);
nand U4914 (N_4914,In_940,In_1588);
or U4915 (N_4915,In_2895,In_163);
xnor U4916 (N_4916,In_1633,In_1238);
and U4917 (N_4917,In_2149,In_290);
xnor U4918 (N_4918,In_221,In_19);
nor U4919 (N_4919,In_1600,In_2078);
nand U4920 (N_4920,In_1949,In_856);
nor U4921 (N_4921,In_817,In_756);
xor U4922 (N_4922,In_2835,In_2667);
and U4923 (N_4923,In_2547,In_2197);
xor U4924 (N_4924,In_2864,In_1634);
or U4925 (N_4925,In_539,In_894);
or U4926 (N_4926,In_731,In_799);
nor U4927 (N_4927,In_1211,In_1375);
nor U4928 (N_4928,In_1709,In_2786);
nand U4929 (N_4929,In_2473,In_2779);
and U4930 (N_4930,In_1389,In_1946);
nor U4931 (N_4931,In_1930,In_113);
nor U4932 (N_4932,In_657,In_726);
nor U4933 (N_4933,In_1035,In_134);
nand U4934 (N_4934,In_2430,In_1039);
xor U4935 (N_4935,In_1523,In_284);
nand U4936 (N_4936,In_1381,In_2906);
and U4937 (N_4937,In_1026,In_1295);
and U4938 (N_4938,In_1639,In_2397);
nand U4939 (N_4939,In_223,In_1224);
xnor U4940 (N_4940,In_1824,In_2939);
or U4941 (N_4941,In_2957,In_2178);
nand U4942 (N_4942,In_351,In_593);
nor U4943 (N_4943,In_2247,In_740);
xnor U4944 (N_4944,In_2636,In_868);
nor U4945 (N_4945,In_2696,In_728);
nor U4946 (N_4946,In_1223,In_336);
xor U4947 (N_4947,In_1908,In_1126);
and U4948 (N_4948,In_2106,In_2344);
xnor U4949 (N_4949,In_1325,In_44);
nand U4950 (N_4950,In_1332,In_1937);
xor U4951 (N_4951,In_2010,In_267);
and U4952 (N_4952,In_439,In_601);
xor U4953 (N_4953,In_593,In_860);
xnor U4954 (N_4954,In_1313,In_873);
nand U4955 (N_4955,In_2297,In_1986);
and U4956 (N_4956,In_541,In_1924);
xnor U4957 (N_4957,In_1495,In_2042);
nor U4958 (N_4958,In_1279,In_1078);
nand U4959 (N_4959,In_1133,In_45);
and U4960 (N_4960,In_1006,In_748);
nand U4961 (N_4961,In_1045,In_1724);
nor U4962 (N_4962,In_1121,In_567);
nor U4963 (N_4963,In_919,In_2880);
nand U4964 (N_4964,In_769,In_2491);
nor U4965 (N_4965,In_2758,In_2524);
xor U4966 (N_4966,In_1295,In_1333);
nor U4967 (N_4967,In_347,In_534);
and U4968 (N_4968,In_882,In_323);
or U4969 (N_4969,In_539,In_1433);
nand U4970 (N_4970,In_987,In_2910);
nor U4971 (N_4971,In_885,In_1427);
or U4972 (N_4972,In_2763,In_2579);
and U4973 (N_4973,In_889,In_1658);
xor U4974 (N_4974,In_1497,In_1801);
xor U4975 (N_4975,In_1610,In_281);
nand U4976 (N_4976,In_2189,In_784);
nand U4977 (N_4977,In_185,In_2233);
nand U4978 (N_4978,In_2657,In_2534);
xnor U4979 (N_4979,In_702,In_398);
xor U4980 (N_4980,In_770,In_2337);
nor U4981 (N_4981,In_1422,In_676);
or U4982 (N_4982,In_2267,In_1098);
nor U4983 (N_4983,In_1456,In_2552);
and U4984 (N_4984,In_2214,In_1900);
xnor U4985 (N_4985,In_1869,In_1614);
or U4986 (N_4986,In_1209,In_333);
nand U4987 (N_4987,In_66,In_2995);
and U4988 (N_4988,In_518,In_1081);
nor U4989 (N_4989,In_2368,In_1736);
nor U4990 (N_4990,In_700,In_1447);
nor U4991 (N_4991,In_1482,In_561);
or U4992 (N_4992,In_1974,In_2598);
or U4993 (N_4993,In_62,In_698);
and U4994 (N_4994,In_2097,In_2968);
and U4995 (N_4995,In_572,In_777);
and U4996 (N_4996,In_1442,In_1770);
or U4997 (N_4997,In_724,In_2083);
nand U4998 (N_4998,In_1009,In_809);
nand U4999 (N_4999,In_974,In_348);
nand U5000 (N_5000,N_581,N_4844);
nand U5001 (N_5001,N_1087,N_2268);
nor U5002 (N_5002,N_3975,N_928);
or U5003 (N_5003,N_3521,N_490);
xnor U5004 (N_5004,N_2702,N_1300);
nor U5005 (N_5005,N_4416,N_1549);
xnor U5006 (N_5006,N_712,N_113);
or U5007 (N_5007,N_4345,N_2709);
xor U5008 (N_5008,N_4239,N_1535);
nand U5009 (N_5009,N_2732,N_4802);
xnor U5010 (N_5010,N_3827,N_2599);
nor U5011 (N_5011,N_375,N_4380);
nor U5012 (N_5012,N_105,N_887);
xor U5013 (N_5013,N_4728,N_4328);
xor U5014 (N_5014,N_2627,N_547);
nor U5015 (N_5015,N_3548,N_1272);
nor U5016 (N_5016,N_4562,N_2923);
nand U5017 (N_5017,N_2551,N_3971);
xor U5018 (N_5018,N_1738,N_4329);
and U5019 (N_5019,N_1135,N_2340);
and U5020 (N_5020,N_1279,N_2484);
xnor U5021 (N_5021,N_4398,N_3883);
or U5022 (N_5022,N_3390,N_4367);
and U5023 (N_5023,N_2930,N_4491);
nor U5024 (N_5024,N_3957,N_4619);
nand U5025 (N_5025,N_3638,N_4637);
and U5026 (N_5026,N_3698,N_1862);
xor U5027 (N_5027,N_497,N_2854);
and U5028 (N_5028,N_1129,N_1899);
xor U5029 (N_5029,N_4001,N_926);
nand U5030 (N_5030,N_445,N_4130);
xnor U5031 (N_5031,N_2160,N_1451);
xnor U5032 (N_5032,N_1554,N_227);
or U5033 (N_5033,N_291,N_754);
or U5034 (N_5034,N_3876,N_1785);
and U5035 (N_5035,N_2515,N_319);
and U5036 (N_5036,N_4667,N_3872);
nand U5037 (N_5037,N_808,N_1583);
nand U5038 (N_5038,N_4630,N_3882);
nand U5039 (N_5039,N_3018,N_431);
or U5040 (N_5040,N_3157,N_1650);
and U5041 (N_5041,N_2757,N_4670);
nor U5042 (N_5042,N_4264,N_4395);
nand U5043 (N_5043,N_1842,N_4701);
nand U5044 (N_5044,N_4094,N_31);
nand U5045 (N_5045,N_2448,N_1482);
nor U5046 (N_5046,N_2740,N_4864);
or U5047 (N_5047,N_1128,N_278);
nand U5048 (N_5048,N_312,N_1218);
and U5049 (N_5049,N_4714,N_4982);
xnor U5050 (N_5050,N_1231,N_3649);
nor U5051 (N_5051,N_4096,N_4731);
nand U5052 (N_5052,N_4471,N_2253);
and U5053 (N_5053,N_2048,N_2027);
nand U5054 (N_5054,N_3010,N_1860);
xor U5055 (N_5055,N_4474,N_1876);
xnor U5056 (N_5056,N_3910,N_407);
nand U5057 (N_5057,N_2910,N_132);
or U5058 (N_5058,N_4241,N_1080);
nand U5059 (N_5059,N_3080,N_2250);
or U5060 (N_5060,N_1735,N_4648);
xor U5061 (N_5061,N_3011,N_1301);
and U5062 (N_5062,N_1179,N_797);
xor U5063 (N_5063,N_2783,N_2667);
or U5064 (N_5064,N_4773,N_3084);
and U5065 (N_5065,N_4876,N_4254);
xor U5066 (N_5066,N_332,N_1149);
nand U5067 (N_5067,N_3111,N_1161);
nand U5068 (N_5068,N_2018,N_4422);
xor U5069 (N_5069,N_1696,N_4616);
nor U5070 (N_5070,N_4358,N_3878);
or U5071 (N_5071,N_662,N_3246);
nor U5072 (N_5072,N_2470,N_2557);
and U5073 (N_5073,N_3518,N_3982);
xnor U5074 (N_5074,N_4321,N_416);
nor U5075 (N_5075,N_145,N_115);
xor U5076 (N_5076,N_1756,N_2016);
and U5077 (N_5077,N_3278,N_42);
nand U5078 (N_5078,N_3424,N_1572);
nor U5079 (N_5079,N_3286,N_3729);
nand U5080 (N_5080,N_3269,N_4739);
and U5081 (N_5081,N_1020,N_4850);
or U5082 (N_5082,N_2257,N_4308);
xnor U5083 (N_5083,N_3807,N_3926);
xor U5084 (N_5084,N_1284,N_2525);
nand U5085 (N_5085,N_914,N_2315);
nor U5086 (N_5086,N_583,N_430);
nand U5087 (N_5087,N_463,N_1626);
and U5088 (N_5088,N_221,N_1186);
or U5089 (N_5089,N_4512,N_83);
xnor U5090 (N_5090,N_1745,N_4995);
nand U5091 (N_5091,N_4436,N_3567);
nor U5092 (N_5092,N_972,N_2066);
or U5093 (N_5093,N_2648,N_2722);
nand U5094 (N_5094,N_386,N_1809);
and U5095 (N_5095,N_3853,N_4266);
nand U5096 (N_5096,N_88,N_1564);
or U5097 (N_5097,N_772,N_213);
xor U5098 (N_5098,N_1000,N_1901);
and U5099 (N_5099,N_2073,N_411);
nor U5100 (N_5100,N_4755,N_1023);
xor U5101 (N_5101,N_654,N_2208);
nor U5102 (N_5102,N_3583,N_3506);
nand U5103 (N_5103,N_399,N_3757);
xnor U5104 (N_5104,N_2405,N_1251);
nand U5105 (N_5105,N_2365,N_2180);
or U5106 (N_5106,N_4617,N_4100);
and U5107 (N_5107,N_4245,N_2922);
xor U5108 (N_5108,N_2869,N_3469);
nor U5109 (N_5109,N_396,N_442);
nor U5110 (N_5110,N_571,N_247);
nand U5111 (N_5111,N_4277,N_2453);
xor U5112 (N_5112,N_483,N_2200);
nor U5113 (N_5113,N_3481,N_4414);
nand U5114 (N_5114,N_2621,N_3662);
xnor U5115 (N_5115,N_3375,N_2611);
xor U5116 (N_5116,N_3299,N_4407);
or U5117 (N_5117,N_822,N_1406);
or U5118 (N_5118,N_4257,N_1173);
and U5119 (N_5119,N_2356,N_477);
nand U5120 (N_5120,N_4752,N_2789);
and U5121 (N_5121,N_3162,N_2086);
nand U5122 (N_5122,N_3262,N_3947);
nor U5123 (N_5123,N_448,N_3444);
or U5124 (N_5124,N_2805,N_4806);
nor U5125 (N_5125,N_1728,N_2796);
and U5126 (N_5126,N_3879,N_1539);
nand U5127 (N_5127,N_4510,N_693);
or U5128 (N_5128,N_865,N_1877);
nor U5129 (N_5129,N_546,N_3364);
xor U5130 (N_5130,N_4333,N_3171);
nor U5131 (N_5131,N_2670,N_905);
nand U5132 (N_5132,N_2110,N_2215);
xnor U5133 (N_5133,N_1935,N_3956);
and U5134 (N_5134,N_3029,N_1648);
nor U5135 (N_5135,N_2028,N_1146);
xor U5136 (N_5136,N_1663,N_4354);
nor U5137 (N_5137,N_4720,N_1096);
xnor U5138 (N_5138,N_3692,N_557);
nor U5139 (N_5139,N_2010,N_1387);
nand U5140 (N_5140,N_2764,N_2843);
nor U5141 (N_5141,N_2972,N_1404);
xnor U5142 (N_5142,N_4852,N_1844);
or U5143 (N_5143,N_1355,N_530);
nand U5144 (N_5144,N_2755,N_952);
nor U5145 (N_5145,N_3789,N_362);
and U5146 (N_5146,N_1617,N_2947);
and U5147 (N_5147,N_2068,N_2905);
and U5148 (N_5148,N_2337,N_1959);
nand U5149 (N_5149,N_4206,N_1085);
or U5150 (N_5150,N_4223,N_1979);
xor U5151 (N_5151,N_858,N_3577);
nor U5152 (N_5152,N_2339,N_3932);
xor U5153 (N_5153,N_4332,N_2478);
nor U5154 (N_5154,N_1646,N_1873);
and U5155 (N_5155,N_3991,N_1900);
xor U5156 (N_5156,N_2111,N_487);
nand U5157 (N_5157,N_2247,N_2326);
xnor U5158 (N_5158,N_3183,N_982);
or U5159 (N_5159,N_158,N_4887);
xnor U5160 (N_5160,N_3132,N_3476);
and U5161 (N_5161,N_3857,N_4676);
nand U5162 (N_5162,N_3595,N_4950);
xnor U5163 (N_5163,N_3530,N_1577);
and U5164 (N_5164,N_2071,N_651);
or U5165 (N_5165,N_3273,N_727);
nor U5166 (N_5166,N_3027,N_2975);
xnor U5167 (N_5167,N_3345,N_1551);
or U5168 (N_5168,N_3682,N_1513);
and U5169 (N_5169,N_1758,N_3373);
xnor U5170 (N_5170,N_714,N_4727);
nand U5171 (N_5171,N_2043,N_717);
nand U5172 (N_5172,N_3621,N_3124);
xor U5173 (N_5173,N_832,N_4338);
and U5174 (N_5174,N_1721,N_2521);
nand U5175 (N_5175,N_3720,N_2304);
xnor U5176 (N_5176,N_3768,N_4009);
xor U5177 (N_5177,N_370,N_2629);
nand U5178 (N_5178,N_4372,N_601);
nand U5179 (N_5179,N_1148,N_4208);
and U5180 (N_5180,N_4896,N_3533);
and U5181 (N_5181,N_4229,N_3938);
or U5182 (N_5182,N_3202,N_3684);
nand U5183 (N_5183,N_4658,N_1528);
nand U5184 (N_5184,N_1007,N_2449);
nor U5185 (N_5185,N_3116,N_3282);
xnor U5186 (N_5186,N_3811,N_3405);
xnor U5187 (N_5187,N_572,N_241);
or U5188 (N_5188,N_218,N_1292);
or U5189 (N_5189,N_3922,N_4168);
nand U5190 (N_5190,N_2392,N_2848);
nand U5191 (N_5191,N_1285,N_3306);
or U5192 (N_5192,N_338,N_921);
or U5193 (N_5193,N_3635,N_1523);
xnor U5194 (N_5194,N_618,N_1731);
or U5195 (N_5195,N_4353,N_1589);
nor U5196 (N_5196,N_3865,N_2772);
nor U5197 (N_5197,N_2004,N_1070);
nand U5198 (N_5198,N_149,N_2784);
nor U5199 (N_5199,N_3646,N_1910);
and U5200 (N_5200,N_1599,N_2876);
nor U5201 (N_5201,N_1636,N_3687);
or U5202 (N_5202,N_682,N_4342);
and U5203 (N_5203,N_1444,N_2756);
nand U5204 (N_5204,N_181,N_1048);
nand U5205 (N_5205,N_4006,N_4113);
nor U5206 (N_5206,N_4230,N_117);
nor U5207 (N_5207,N_2959,N_2329);
xnor U5208 (N_5208,N_3175,N_78);
and U5209 (N_5209,N_3316,N_4035);
or U5210 (N_5210,N_1770,N_1530);
xnor U5211 (N_5211,N_4234,N_3560);
and U5212 (N_5212,N_3397,N_1401);
nor U5213 (N_5213,N_398,N_3025);
xnor U5214 (N_5214,N_2428,N_4810);
nand U5215 (N_5215,N_3417,N_1982);
nor U5216 (N_5216,N_93,N_3398);
or U5217 (N_5217,N_3674,N_1260);
nand U5218 (N_5218,N_3877,N_919);
and U5219 (N_5219,N_2852,N_76);
nand U5220 (N_5220,N_1452,N_831);
nor U5221 (N_5221,N_3748,N_4629);
and U5222 (N_5222,N_1180,N_4819);
nand U5223 (N_5223,N_2371,N_2167);
xnor U5224 (N_5224,N_846,N_4460);
and U5225 (N_5225,N_1291,N_4984);
xor U5226 (N_5226,N_470,N_53);
nand U5227 (N_5227,N_2683,N_2292);
and U5228 (N_5228,N_4051,N_4833);
xor U5229 (N_5229,N_390,N_453);
nor U5230 (N_5230,N_3115,N_4893);
xor U5231 (N_5231,N_2572,N_3203);
xnor U5232 (N_5232,N_273,N_2079);
nand U5233 (N_5233,N_2656,N_4697);
nand U5234 (N_5234,N_2067,N_509);
or U5235 (N_5235,N_2929,N_4722);
and U5236 (N_5236,N_3970,N_4786);
nand U5237 (N_5237,N_1158,N_1392);
nor U5238 (N_5238,N_3055,N_3458);
xnor U5239 (N_5239,N_368,N_4974);
and U5240 (N_5240,N_2089,N_3494);
or U5241 (N_5241,N_1229,N_45);
or U5242 (N_5242,N_1062,N_734);
nor U5243 (N_5243,N_3448,N_4285);
or U5244 (N_5244,N_3146,N_1916);
nor U5245 (N_5245,N_1361,N_261);
nand U5246 (N_5246,N_140,N_4016);
xnor U5247 (N_5247,N_2862,N_3313);
nand U5248 (N_5248,N_2858,N_755);
nand U5249 (N_5249,N_2005,N_3047);
xor U5250 (N_5250,N_1372,N_1647);
or U5251 (N_5251,N_2890,N_1664);
nor U5252 (N_5252,N_1089,N_2322);
and U5253 (N_5253,N_2896,N_1418);
nand U5254 (N_5254,N_3048,N_3507);
or U5255 (N_5255,N_2276,N_4290);
xnor U5256 (N_5256,N_4817,N_315);
xor U5257 (N_5257,N_4917,N_896);
xnor U5258 (N_5258,N_1851,N_1483);
xnor U5259 (N_5259,N_16,N_1861);
nor U5260 (N_5260,N_237,N_4440);
nand U5261 (N_5261,N_787,N_3322);
or U5262 (N_5262,N_343,N_2694);
nand U5263 (N_5263,N_1220,N_4596);
xor U5264 (N_5264,N_4749,N_1475);
nand U5265 (N_5265,N_3172,N_769);
xnor U5266 (N_5266,N_244,N_3230);
nor U5267 (N_5267,N_3579,N_1937);
nand U5268 (N_5268,N_192,N_1618);
and U5269 (N_5269,N_2230,N_3988);
and U5270 (N_5270,N_258,N_993);
and U5271 (N_5271,N_3454,N_923);
nand U5272 (N_5272,N_957,N_3867);
xor U5273 (N_5273,N_984,N_4700);
nor U5274 (N_5274,N_2127,N_3484);
and U5275 (N_5275,N_3263,N_424);
and U5276 (N_5276,N_562,N_4260);
or U5277 (N_5277,N_2968,N_4082);
and U5278 (N_5278,N_1039,N_58);
or U5279 (N_5279,N_4915,N_4712);
xor U5280 (N_5280,N_1038,N_4832);
xor U5281 (N_5281,N_1722,N_2939);
and U5282 (N_5282,N_650,N_2260);
nor U5283 (N_5283,N_1083,N_99);
xor U5284 (N_5284,N_3223,N_1332);
xor U5285 (N_5285,N_3228,N_2049);
nand U5286 (N_5286,N_4964,N_635);
and U5287 (N_5287,N_2446,N_2888);
nand U5288 (N_5288,N_4603,N_1115);
or U5289 (N_5289,N_4278,N_1026);
nand U5290 (N_5290,N_4800,N_32);
nor U5291 (N_5291,N_413,N_4078);
and U5292 (N_5292,N_2914,N_4678);
and U5293 (N_5293,N_3056,N_563);
nand U5294 (N_5294,N_2948,N_2314);
or U5295 (N_5295,N_2361,N_959);
xnor U5296 (N_5296,N_2794,N_1184);
and U5297 (N_5297,N_4976,N_1967);
and U5298 (N_5298,N_3350,N_821);
or U5299 (N_5299,N_2823,N_657);
and U5300 (N_5300,N_4164,N_2149);
nor U5301 (N_5301,N_3792,N_3571);
or U5302 (N_5302,N_1710,N_2941);
or U5303 (N_5303,N_3088,N_1030);
xnor U5304 (N_5304,N_2800,N_2150);
nor U5305 (N_5305,N_3090,N_2135);
nand U5306 (N_5306,N_2891,N_4726);
or U5307 (N_5307,N_2139,N_2133);
nor U5308 (N_5308,N_3917,N_1690);
and U5309 (N_5309,N_1852,N_41);
or U5310 (N_5310,N_2989,N_2826);
and U5311 (N_5311,N_46,N_2567);
and U5312 (N_5312,N_328,N_3414);
or U5313 (N_5313,N_4531,N_3944);
or U5314 (N_5314,N_2785,N_507);
nor U5315 (N_5315,N_534,N_403);
and U5316 (N_5316,N_1928,N_541);
nor U5317 (N_5317,N_2509,N_4565);
or U5318 (N_5318,N_3788,N_1364);
nand U5319 (N_5319,N_3667,N_3436);
nor U5320 (N_5320,N_354,N_4303);
and U5321 (N_5321,N_2185,N_1088);
or U5322 (N_5322,N_2672,N_2353);
or U5323 (N_5323,N_4317,N_4190);
and U5324 (N_5324,N_359,N_933);
or U5325 (N_5325,N_3831,N_1866);
nand U5326 (N_5326,N_607,N_2717);
nand U5327 (N_5327,N_2926,N_410);
xor U5328 (N_5328,N_3064,N_3532);
or U5329 (N_5329,N_1338,N_2597);
nand U5330 (N_5330,N_3960,N_1059);
nand U5331 (N_5331,N_2205,N_3180);
nand U5332 (N_5332,N_1494,N_848);
and U5333 (N_5333,N_765,N_2729);
and U5334 (N_5334,N_190,N_1981);
nor U5335 (N_5335,N_2918,N_2343);
and U5336 (N_5336,N_3200,N_3834);
and U5337 (N_5337,N_4275,N_231);
nand U5338 (N_5338,N_1133,N_324);
and U5339 (N_5339,N_974,N_1134);
nand U5340 (N_5340,N_1490,N_3509);
nor U5341 (N_5341,N_2737,N_3429);
and U5342 (N_5342,N_1189,N_1267);
nand U5343 (N_5343,N_2346,N_2380);
and U5344 (N_5344,N_1357,N_2282);
and U5345 (N_5345,N_1233,N_4926);
xor U5346 (N_5346,N_14,N_367);
and U5347 (N_5347,N_1014,N_1055);
or U5348 (N_5348,N_1420,N_2194);
and U5349 (N_5349,N_3733,N_1704);
nor U5350 (N_5350,N_4425,N_326);
or U5351 (N_5351,N_3707,N_773);
and U5352 (N_5352,N_2791,N_4665);
nand U5353 (N_5353,N_2708,N_3978);
or U5354 (N_5354,N_2466,N_4989);
nor U5355 (N_5355,N_1840,N_4117);
nand U5356 (N_5356,N_404,N_4729);
nor U5357 (N_5357,N_4319,N_852);
xnor U5358 (N_5358,N_4000,N_1765);
xor U5359 (N_5359,N_2903,N_3589);
xor U5360 (N_5360,N_1829,N_302);
or U5361 (N_5361,N_4450,N_3997);
nand U5362 (N_5362,N_4088,N_4520);
or U5363 (N_5363,N_2798,N_4962);
xor U5364 (N_5364,N_1805,N_591);
nand U5365 (N_5365,N_4788,N_2938);
or U5366 (N_5366,N_2184,N_1340);
nor U5367 (N_5367,N_1819,N_1571);
nand U5368 (N_5368,N_1653,N_2088);
or U5369 (N_5369,N_3137,N_4948);
and U5370 (N_5370,N_671,N_3093);
nor U5371 (N_5371,N_1709,N_309);
and U5372 (N_5372,N_4740,N_1703);
nand U5373 (N_5373,N_2999,N_1330);
nor U5374 (N_5374,N_2494,N_1421);
or U5375 (N_5375,N_1563,N_570);
xnor U5376 (N_5376,N_1061,N_4977);
nand U5377 (N_5377,N_3452,N_389);
or U5378 (N_5378,N_2703,N_3451);
xnor U5379 (N_5379,N_2302,N_316);
xor U5380 (N_5380,N_967,N_3858);
nor U5381 (N_5381,N_4718,N_2991);
nor U5382 (N_5382,N_21,N_1514);
xor U5383 (N_5383,N_4542,N_4042);
or U5384 (N_5384,N_2677,N_2698);
nand U5385 (N_5385,N_893,N_3310);
xnor U5386 (N_5386,N_439,N_835);
nor U5387 (N_5387,N_874,N_4886);
xnor U5388 (N_5388,N_3184,N_1397);
nor U5389 (N_5389,N_1001,N_2472);
and U5390 (N_5390,N_3937,N_2916);
and U5391 (N_5391,N_2024,N_2602);
nor U5392 (N_5392,N_593,N_3095);
nor U5393 (N_5393,N_1101,N_692);
or U5394 (N_5394,N_4438,N_3948);
or U5395 (N_5395,N_489,N_3089);
nand U5396 (N_5396,N_2265,N_3083);
nor U5397 (N_5397,N_3652,N_1655);
xor U5398 (N_5398,N_783,N_899);
nand U5399 (N_5399,N_2015,N_2394);
nor U5400 (N_5400,N_2499,N_3987);
nand U5401 (N_5401,N_353,N_2639);
nor U5402 (N_5402,N_1907,N_3079);
xnor U5403 (N_5403,N_2270,N_3076);
xor U5404 (N_5404,N_556,N_2822);
or U5405 (N_5405,N_4043,N_438);
xnor U5406 (N_5406,N_299,N_1657);
or U5407 (N_5407,N_4897,N_4177);
nand U5408 (N_5408,N_4040,N_2299);
or U5409 (N_5409,N_397,N_11);
xnor U5410 (N_5410,N_4368,N_3040);
xnor U5411 (N_5411,N_1651,N_3468);
nand U5412 (N_5412,N_4821,N_4487);
nor U5413 (N_5413,N_2885,N_1224);
or U5414 (N_5414,N_1593,N_2512);
xnor U5415 (N_5415,N_123,N_111);
and U5416 (N_5416,N_4517,N_499);
nor U5417 (N_5417,N_1058,N_3252);
nand U5418 (N_5418,N_4889,N_548);
xnor U5419 (N_5419,N_4932,N_1402);
xor U5420 (N_5420,N_1309,N_2650);
xor U5421 (N_5421,N_4627,N_2174);
and U5422 (N_5422,N_2691,N_738);
and U5423 (N_5423,N_4966,N_3379);
or U5424 (N_5424,N_4608,N_1348);
and U5425 (N_5425,N_1543,N_3820);
and U5426 (N_5426,N_839,N_2955);
xnor U5427 (N_5427,N_861,N_3120);
xor U5428 (N_5428,N_1455,N_3873);
or U5429 (N_5429,N_3958,N_4990);
and U5430 (N_5430,N_1195,N_1323);
xnor U5431 (N_5431,N_851,N_4635);
xnor U5432 (N_5432,N_3845,N_3372);
and U5433 (N_5433,N_3486,N_529);
nor U5434 (N_5434,N_2091,N_3527);
xnor U5435 (N_5435,N_4150,N_2839);
and U5436 (N_5436,N_339,N_2342);
nor U5437 (N_5437,N_1449,N_3890);
or U5438 (N_5438,N_3655,N_3283);
and U5439 (N_5439,N_643,N_1202);
and U5440 (N_5440,N_4157,N_3367);
or U5441 (N_5441,N_4281,N_2931);
nand U5442 (N_5442,N_2207,N_3994);
nor U5443 (N_5443,N_2338,N_2859);
xor U5444 (N_5444,N_1671,N_3799);
nor U5445 (N_5445,N_1958,N_4271);
nand U5446 (N_5446,N_3437,N_3403);
xnor U5447 (N_5447,N_68,N_1586);
nand U5448 (N_5448,N_4331,N_1744);
nand U5449 (N_5449,N_4205,N_4767);
xor U5450 (N_5450,N_736,N_102);
nor U5451 (N_5451,N_1373,N_1911);
nor U5452 (N_5452,N_3099,N_1970);
xor U5453 (N_5453,N_201,N_515);
and U5454 (N_5454,N_4099,N_2186);
xor U5455 (N_5455,N_681,N_4508);
nor U5456 (N_5456,N_2684,N_3690);
xor U5457 (N_5457,N_1383,N_677);
xor U5458 (N_5458,N_1232,N_3888);
or U5459 (N_5459,N_4680,N_1286);
or U5460 (N_5460,N_3256,N_2956);
or U5461 (N_5461,N_3150,N_2598);
xor U5462 (N_5462,N_2324,N_2395);
and U5463 (N_5463,N_3411,N_3965);
and U5464 (N_5464,N_2408,N_3568);
nand U5465 (N_5465,N_3701,N_243);
nor U5466 (N_5466,N_1424,N_1500);
nand U5467 (N_5467,N_1906,N_108);
and U5468 (N_5468,N_385,N_4550);
or U5469 (N_5469,N_1912,N_1416);
or U5470 (N_5470,N_311,N_2192);
xor U5471 (N_5471,N_325,N_2435);
nand U5472 (N_5472,N_970,N_1649);
nor U5473 (N_5473,N_2424,N_2155);
or U5474 (N_5474,N_2264,N_2196);
nor U5475 (N_5475,N_3547,N_642);
or U5476 (N_5476,N_1591,N_2105);
and U5477 (N_5477,N_3607,N_4660);
nand U5478 (N_5478,N_1028,N_4685);
or U5479 (N_5479,N_1707,N_285);
xnor U5480 (N_5480,N_3393,N_4656);
nand U5481 (N_5481,N_2765,N_2415);
nand U5482 (N_5482,N_4859,N_2370);
nand U5483 (N_5483,N_3192,N_3308);
or U5484 (N_5484,N_2498,N_4169);
nand U5485 (N_5485,N_2526,N_1848);
nor U5486 (N_5486,N_3526,N_3522);
nand U5487 (N_5487,N_1227,N_2420);
nand U5488 (N_5488,N_3995,N_1266);
xnor U5489 (N_5489,N_4796,N_4944);
or U5490 (N_5490,N_909,N_1201);
xnor U5491 (N_5491,N_2770,N_2510);
nor U5492 (N_5492,N_3678,N_2003);
and U5493 (N_5493,N_2144,N_4534);
and U5494 (N_5494,N_3087,N_2502);
and U5495 (N_5495,N_3474,N_4336);
nor U5496 (N_5496,N_491,N_2833);
nand U5497 (N_5497,N_2595,N_945);
or U5498 (N_5498,N_2219,N_3033);
xnor U5499 (N_5499,N_4444,N_2871);
xnor U5500 (N_5500,N_203,N_4909);
and U5501 (N_5501,N_4936,N_3128);
nand U5502 (N_5502,N_2347,N_1798);
nor U5503 (N_5503,N_162,N_3512);
or U5504 (N_5504,N_3374,N_1033);
or U5505 (N_5505,N_2036,N_61);
and U5506 (N_5506,N_4794,N_4465);
nor U5507 (N_5507,N_876,N_2078);
nand U5508 (N_5508,N_62,N_3817);
and U5509 (N_5509,N_1385,N_2577);
nor U5510 (N_5510,N_4705,N_436);
xnor U5511 (N_5511,N_4121,N_1010);
nand U5512 (N_5512,N_3779,N_992);
nand U5513 (N_5513,N_695,N_3231);
nand U5514 (N_5514,N_3921,N_3710);
and U5515 (N_5515,N_4539,N_2372);
or U5516 (N_5516,N_163,N_2305);
nand U5517 (N_5517,N_3351,N_1717);
and U5518 (N_5518,N_892,N_1193);
and U5519 (N_5519,N_3304,N_3147);
xnor U5520 (N_5520,N_1943,N_4227);
nor U5521 (N_5521,N_742,N_4757);
and U5522 (N_5522,N_4702,N_2383);
and U5523 (N_5523,N_3179,N_4552);
or U5524 (N_5524,N_4938,N_4013);
or U5525 (N_5525,N_1190,N_1157);
or U5526 (N_5526,N_3542,N_3100);
and U5527 (N_5527,N_165,N_2283);
nor U5528 (N_5528,N_460,N_59);
and U5529 (N_5529,N_481,N_3220);
nor U5530 (N_5530,N_2272,N_39);
and U5531 (N_5531,N_1510,N_2720);
nor U5532 (N_5532,N_1737,N_4584);
xor U5533 (N_5533,N_2280,N_4771);
nand U5534 (N_5534,N_1817,N_561);
nand U5535 (N_5535,N_3572,N_2065);
or U5536 (N_5536,N_4511,N_3062);
or U5537 (N_5537,N_4840,N_2355);
nor U5538 (N_5538,N_2454,N_3097);
xnor U5539 (N_5539,N_33,N_1199);
nand U5540 (N_5540,N_1429,N_1097);
or U5541 (N_5541,N_3242,N_1130);
nor U5542 (N_5542,N_3327,N_224);
xor U5543 (N_5543,N_629,N_79);
or U5544 (N_5544,N_4265,N_4614);
and U5545 (N_5545,N_153,N_4502);
and U5546 (N_5546,N_260,N_1630);
nand U5547 (N_5547,N_3569,N_2625);
nor U5548 (N_5548,N_915,N_4778);
nand U5549 (N_5549,N_466,N_3537);
nand U5550 (N_5550,N_3801,N_2777);
or U5551 (N_5551,N_1432,N_4588);
and U5552 (N_5552,N_2183,N_845);
and U5553 (N_5553,N_2399,N_711);
nor U5554 (N_5554,N_1965,N_3848);
nand U5555 (N_5555,N_372,N_4361);
or U5556 (N_5556,N_2148,N_564);
and U5557 (N_5557,N_2021,N_3787);
or U5558 (N_5558,N_400,N_1386);
xnor U5559 (N_5559,N_4543,N_701);
nor U5560 (N_5560,N_3764,N_810);
xnor U5561 (N_5561,N_1019,N_4894);
nor U5562 (N_5562,N_4405,N_2902);
nand U5563 (N_5563,N_3410,N_4315);
and U5564 (N_5564,N_4625,N_253);
nor U5565 (N_5565,N_2094,N_2511);
nand U5566 (N_5566,N_833,N_532);
nor U5567 (N_5567,N_2386,N_1932);
or U5568 (N_5568,N_4377,N_3950);
or U5569 (N_5569,N_3604,N_3859);
xnor U5570 (N_5570,N_495,N_3830);
nand U5571 (N_5571,N_3868,N_2427);
or U5572 (N_5572,N_2838,N_3248);
or U5573 (N_5573,N_199,N_3836);
or U5574 (N_5574,N_3319,N_2492);
nand U5575 (N_5575,N_1110,N_4054);
or U5576 (N_5576,N_3239,N_1896);
xnor U5577 (N_5577,N_725,N_440);
and U5578 (N_5578,N_3665,N_284);
xor U5579 (N_5579,N_3616,N_2334);
or U5580 (N_5580,N_1567,N_4455);
nand U5581 (N_5581,N_3255,N_2224);
or U5582 (N_5582,N_1431,N_4949);
nor U5583 (N_5583,N_3348,N_114);
xor U5584 (N_5584,N_753,N_2190);
nand U5585 (N_5585,N_1947,N_2875);
and U5586 (N_5586,N_8,N_2735);
xnor U5587 (N_5587,N_96,N_3092);
and U5588 (N_5588,N_817,N_2084);
nor U5589 (N_5589,N_2830,N_2);
xnor U5590 (N_5590,N_2895,N_587);
and U5591 (N_5591,N_3786,N_4784);
nor U5592 (N_5592,N_3973,N_1076);
xnor U5593 (N_5593,N_1217,N_4129);
nand U5594 (N_5594,N_4716,N_2993);
xor U5595 (N_5595,N_3466,N_2828);
or U5596 (N_5596,N_590,N_2977);
nand U5597 (N_5597,N_880,N_433);
and U5598 (N_5598,N_216,N_4369);
xor U5599 (N_5599,N_3185,N_4313);
or U5600 (N_5600,N_1403,N_4055);
nand U5601 (N_5601,N_1290,N_4537);
xor U5602 (N_5602,N_369,N_3415);
nor U5603 (N_5603,N_2032,N_1075);
or U5604 (N_5604,N_2357,N_2063);
xnor U5605 (N_5605,N_1336,N_864);
xor U5606 (N_5606,N_4519,N_4953);
and U5607 (N_5607,N_2460,N_2744);
nor U5608 (N_5608,N_847,N_1141);
nor U5609 (N_5609,N_2285,N_1305);
nor U5610 (N_5610,N_318,N_3218);
or U5611 (N_5611,N_4418,N_414);
xor U5612 (N_5612,N_971,N_998);
nor U5613 (N_5613,N_1760,N_2465);
nand U5614 (N_5614,N_2560,N_4356);
xor U5615 (N_5615,N_1468,N_250);
xnor U5616 (N_5616,N_4002,N_2564);
nand U5617 (N_5617,N_3736,N_2842);
or U5618 (N_5618,N_49,N_2145);
or U5619 (N_5619,N_2437,N_718);
xor U5620 (N_5620,N_4152,N_4963);
nor U5621 (N_5621,N_4586,N_1700);
nand U5622 (N_5622,N_2335,N_4244);
nand U5623 (N_5623,N_3703,N_4737);
or U5624 (N_5624,N_595,N_1306);
and U5625 (N_5625,N_4692,N_4498);
nor U5626 (N_5626,N_2739,N_2104);
xor U5627 (N_5627,N_263,N_4935);
xor U5628 (N_5628,N_3505,N_4214);
or U5629 (N_5629,N_3144,N_4185);
or U5630 (N_5630,N_803,N_4004);
or U5631 (N_5631,N_1716,N_10);
and U5632 (N_5632,N_1063,N_4836);
and U5633 (N_5633,N_2962,N_960);
nand U5634 (N_5634,N_4388,N_4943);
and U5635 (N_5635,N_4175,N_4744);
and U5636 (N_5636,N_1016,N_1230);
nor U5637 (N_5637,N_3261,N_1448);
or U5638 (N_5638,N_4791,N_329);
and U5639 (N_5639,N_4914,N_1534);
xor U5640 (N_5640,N_4397,N_694);
nor U5641 (N_5641,N_469,N_1188);
nand U5642 (N_5642,N_87,N_43);
nand U5643 (N_5643,N_1398,N_1031);
xor U5644 (N_5644,N_2029,N_3480);
nand U5645 (N_5645,N_2932,N_3809);
nor U5646 (N_5646,N_2976,N_2000);
and U5647 (N_5647,N_2491,N_310);
or U5648 (N_5648,N_3266,N_679);
or U5649 (N_5649,N_3344,N_3758);
nor U5650 (N_5650,N_1548,N_879);
xnor U5651 (N_5651,N_3204,N_1497);
xnor U5652 (N_5652,N_2607,N_4435);
nor U5653 (N_5653,N_1846,N_3026);
xnor U5654 (N_5654,N_3385,N_322);
xnor U5655 (N_5655,N_321,N_1547);
nand U5656 (N_5656,N_1839,N_1837);
or U5657 (N_5657,N_3818,N_1678);
or U5658 (N_5658,N_2908,N_4869);
xor U5659 (N_5659,N_906,N_3737);
xnor U5660 (N_5660,N_2248,N_3609);
or U5661 (N_5661,N_2969,N_1964);
nand U5662 (N_5662,N_809,N_18);
nor U5663 (N_5663,N_4364,N_2191);
or U5664 (N_5664,N_2459,N_4954);
or U5665 (N_5665,N_2780,N_4933);
xnor U5666 (N_5666,N_1025,N_4882);
xor U5667 (N_5667,N_3394,N_1108);
nor U5668 (N_5668,N_1624,N_4795);
and U5669 (N_5669,N_3719,N_4288);
and U5670 (N_5670,N_2669,N_4919);
and U5671 (N_5671,N_743,N_819);
and U5672 (N_5672,N_3931,N_3177);
or U5673 (N_5673,N_456,N_2378);
nand U5674 (N_5674,N_2136,N_1371);
and U5675 (N_5675,N_1612,N_2644);
xnor U5676 (N_5676,N_1827,N_2390);
nand U5677 (N_5677,N_2434,N_4107);
xor U5678 (N_5678,N_4693,N_1865);
and U5679 (N_5679,N_2037,N_1637);
xnor U5680 (N_5680,N_3307,N_4741);
or U5681 (N_5681,N_2189,N_4626);
xnor U5682 (N_5682,N_3581,N_4939);
and U5683 (N_5683,N_867,N_1461);
nand U5684 (N_5684,N_2927,N_1814);
xor U5685 (N_5685,N_178,N_3490);
and U5686 (N_5686,N_3866,N_4807);
or U5687 (N_5687,N_3176,N_4469);
nand U5688 (N_5688,N_1498,N_1095);
nand U5689 (N_5689,N_297,N_2025);
and U5690 (N_5690,N_3819,N_678);
xnor U5691 (N_5691,N_3594,N_2223);
or U5692 (N_5692,N_4114,N_2209);
nor U5693 (N_5693,N_4681,N_2581);
xor U5694 (N_5694,N_3449,N_334);
xor U5695 (N_5695,N_2401,N_4337);
and U5696 (N_5696,N_2810,N_4960);
nor U5697 (N_5697,N_1147,N_930);
nand U5698 (N_5698,N_3031,N_3110);
or U5699 (N_5699,N_1393,N_1441);
nor U5700 (N_5700,N_4868,N_409);
or U5701 (N_5701,N_3250,N_2748);
xor U5702 (N_5702,N_1047,N_920);
xnor U5703 (N_5703,N_2109,N_2767);
nor U5704 (N_5704,N_3510,N_3245);
or U5705 (N_5705,N_2658,N_3311);
nand U5706 (N_5706,N_3284,N_1712);
nand U5707 (N_5707,N_2475,N_1480);
nand U5708 (N_5708,N_4570,N_2591);
or U5709 (N_5709,N_4022,N_4870);
or U5710 (N_5710,N_4297,N_524);
xor U5711 (N_5711,N_4865,N_2821);
xor U5712 (N_5712,N_3035,N_944);
or U5713 (N_5713,N_973,N_585);
nor U5714 (N_5714,N_1064,N_1343);
and U5715 (N_5715,N_1767,N_1245);
nand U5716 (N_5716,N_358,N_2412);
or U5717 (N_5717,N_4147,N_995);
nand U5718 (N_5718,N_3689,N_980);
nor U5719 (N_5719,N_3501,N_356);
xnor U5720 (N_5720,N_2009,N_3317);
xnor U5721 (N_5721,N_886,N_1820);
and U5722 (N_5722,N_378,N_2236);
nor U5723 (N_5723,N_3550,N_2178);
or U5724 (N_5724,N_4684,N_4477);
nand U5725 (N_5725,N_3191,N_3182);
nor U5726 (N_5726,N_475,N_214);
nor U5727 (N_5727,N_207,N_4219);
nand U5728 (N_5728,N_669,N_3435);
or U5729 (N_5729,N_3821,N_184);
and U5730 (N_5730,N_2500,N_3695);
or U5731 (N_5731,N_2655,N_2713);
and U5732 (N_5732,N_1749,N_2741);
or U5733 (N_5733,N_1349,N_3636);
nand U5734 (N_5734,N_922,N_2206);
nand U5735 (N_5735,N_3717,N_1427);
or U5736 (N_5736,N_579,N_3752);
nand U5737 (N_5737,N_4276,N_4753);
and U5738 (N_5738,N_983,N_1694);
xnor U5739 (N_5739,N_4124,N_4581);
and U5740 (N_5740,N_3874,N_4632);
and U5741 (N_5741,N_2336,N_1702);
nor U5742 (N_5742,N_3380,N_3240);
nand U5743 (N_5743,N_4518,N_2853);
or U5744 (N_5744,N_3722,N_2034);
xnor U5745 (N_5745,N_3457,N_994);
xor U5746 (N_5746,N_1008,N_2497);
nand U5747 (N_5747,N_1859,N_1106);
and U5748 (N_5748,N_3826,N_60);
nor U5749 (N_5749,N_638,N_2216);
xor U5750 (N_5750,N_2600,N_1454);
nor U5751 (N_5751,N_4898,N_188);
nand U5752 (N_5752,N_4076,N_1116);
nor U5753 (N_5753,N_2188,N_2107);
or U5754 (N_5754,N_4590,N_4351);
nand U5755 (N_5755,N_2953,N_4582);
nand U5756 (N_5756,N_1856,N_4605);
or U5757 (N_5757,N_1665,N_280);
or U5758 (N_5758,N_4561,N_3487);
xnor U5759 (N_5759,N_1903,N_3065);
nor U5760 (N_5760,N_3163,N_4267);
or U5761 (N_5761,N_1369,N_2878);
or U5762 (N_5762,N_2064,N_2716);
or U5763 (N_5763,N_4657,N_2837);
xor U5764 (N_5764,N_9,N_781);
nor U5765 (N_5765,N_3658,N_4480);
nor U5766 (N_5766,N_2804,N_4556);
nor U5767 (N_5767,N_1711,N_3331);
nand U5768 (N_5768,N_4623,N_4327);
nand U5769 (N_5769,N_3908,N_1044);
and U5770 (N_5770,N_2163,N_953);
nand U5771 (N_5771,N_1685,N_454);
nand U5772 (N_5772,N_1909,N_2603);
nor U5773 (N_5773,N_2398,N_597);
nand U5774 (N_5774,N_4125,N_1512);
nand U5775 (N_5775,N_4452,N_4867);
xor U5776 (N_5776,N_2530,N_4863);
and U5777 (N_5777,N_1321,N_568);
nor U5778 (N_5778,N_3381,N_4299);
or U5779 (N_5779,N_200,N_1382);
or U5780 (N_5780,N_4613,N_1643);
xnor U5781 (N_5781,N_4703,N_3940);
nand U5782 (N_5782,N_4952,N_746);
nand U5783 (N_5783,N_116,N_2364);
nor U5784 (N_5784,N_1897,N_1682);
xnor U5785 (N_5785,N_4507,N_3072);
nand U5786 (N_5786,N_4120,N_4375);
nor U5787 (N_5787,N_4008,N_3949);
nand U5788 (N_5788,N_580,N_3660);
nand U5789 (N_5789,N_3164,N_3840);
xnor U5790 (N_5790,N_705,N_3020);
nand U5791 (N_5791,N_1131,N_962);
or U5792 (N_5792,N_179,N_4430);
or U5793 (N_5793,N_4643,N_330);
xnor U5794 (N_5794,N_2633,N_2588);
nor U5795 (N_5795,N_4902,N_4034);
nor U5796 (N_5796,N_4210,N_3959);
or U5797 (N_5797,N_4083,N_4818);
xnor U5798 (N_5798,N_1930,N_4620);
nor U5799 (N_5799,N_418,N_615);
or U5800 (N_5800,N_4109,N_4569);
xnor U5801 (N_5801,N_520,N_4826);
or U5802 (N_5802,N_594,N_4506);
nor U5803 (N_5803,N_3942,N_4843);
or U5804 (N_5804,N_1705,N_3901);
or U5805 (N_5805,N_1376,N_4017);
and U5806 (N_5806,N_2766,N_1797);
nand U5807 (N_5807,N_3712,N_3069);
and U5808 (N_5808,N_2080,N_2213);
nor U5809 (N_5809,N_1610,N_3053);
and U5810 (N_5810,N_347,N_4032);
and U5811 (N_5811,N_2323,N_4816);
nand U5812 (N_5812,N_1875,N_432);
nor U5813 (N_5813,N_428,N_1521);
and U5814 (N_5814,N_522,N_1243);
xor U5815 (N_5815,N_1695,N_242);
and U5816 (N_5816,N_3524,N_537);
and U5817 (N_5817,N_3142,N_3427);
or U5818 (N_5818,N_4812,N_697);
and U5819 (N_5819,N_661,N_189);
xor U5820 (N_5820,N_3113,N_1121);
nand U5821 (N_5821,N_1561,N_4568);
and U5822 (N_5822,N_2646,N_1172);
xnor U5823 (N_5823,N_3155,N_4668);
and U5824 (N_5824,N_194,N_3843);
nor U5825 (N_5825,N_2426,N_3446);
xor U5826 (N_5826,N_2966,N_560);
or U5827 (N_5827,N_1049,N_2464);
nand U5828 (N_5828,N_1052,N_4694);
or U5829 (N_5829,N_3564,N_890);
nor U5830 (N_5830,N_3885,N_239);
nand U5831 (N_5831,N_1312,N_3669);
and U5832 (N_5832,N_1159,N_1962);
xnor U5833 (N_5833,N_940,N_3747);
nor U5834 (N_5834,N_4597,N_4306);
nor U5835 (N_5835,N_3915,N_1219);
nand U5836 (N_5836,N_86,N_2996);
and U5837 (N_5837,N_3861,N_1098);
nor U5838 (N_5838,N_1550,N_3213);
xor U5839 (N_5839,N_505,N_4289);
nand U5840 (N_5840,N_3413,N_3694);
xor U5841 (N_5841,N_2044,N_4479);
nand U5842 (N_5842,N_806,N_437);
nand U5843 (N_5843,N_778,N_665);
and U5844 (N_5844,N_3140,N_1337);
or U5845 (N_5845,N_2311,N_4609);
and U5846 (N_5846,N_230,N_4780);
and U5847 (N_5847,N_3377,N_3361);
or U5848 (N_5848,N_3421,N_966);
or U5849 (N_5849,N_37,N_535);
or U5850 (N_5850,N_2085,N_2604);
and U5851 (N_5851,N_2758,N_4366);
or U5852 (N_5852,N_3969,N_1204);
nand U5853 (N_5853,N_210,N_963);
xnor U5854 (N_5854,N_2724,N_3101);
or U5855 (N_5855,N_1919,N_4766);
and U5856 (N_5856,N_1985,N_1289);
xor U5857 (N_5857,N_1200,N_1363);
xnor U5858 (N_5858,N_4745,N_2457);
nand U5859 (N_5859,N_2535,N_807);
nand U5860 (N_5860,N_388,N_2911);
nand U5861 (N_5861,N_3528,N_3201);
or U5862 (N_5862,N_3061,N_1339);
and U5863 (N_5863,N_2433,N_2074);
or U5864 (N_5864,N_4046,N_2541);
and U5865 (N_5865,N_602,N_4018);
or U5866 (N_5866,N_3005,N_2070);
and U5867 (N_5867,N_3766,N_4996);
or U5868 (N_5868,N_1249,N_1518);
xnor U5869 (N_5869,N_2529,N_1997);
nor U5870 (N_5870,N_652,N_4246);
xnor U5871 (N_5871,N_2522,N_4615);
or U5872 (N_5872,N_4193,N_3916);
and U5873 (N_5873,N_327,N_3152);
or U5874 (N_5874,N_2933,N_647);
nand U5875 (N_5875,N_220,N_999);
nand U5876 (N_5876,N_2847,N_4072);
nor U5877 (N_5877,N_308,N_2618);
xnor U5878 (N_5878,N_4411,N_1238);
xnor U5879 (N_5879,N_3354,N_2552);
xor U5880 (N_5880,N_3045,N_3586);
xnor U5881 (N_5881,N_3891,N_3541);
nor U5882 (N_5882,N_4387,N_2204);
or U5883 (N_5883,N_3105,N_4412);
nand U5884 (N_5884,N_4975,N_510);
and U5885 (N_5885,N_796,N_24);
or U5886 (N_5886,N_2369,N_2083);
nand U5887 (N_5887,N_1592,N_4160);
xor U5888 (N_5888,N_1488,N_4010);
or U5889 (N_5889,N_1092,N_1746);
or U5890 (N_5890,N_1961,N_592);
xnor U5891 (N_5891,N_3741,N_1216);
or U5892 (N_5892,N_610,N_760);
nor U5893 (N_5893,N_3841,N_889);
nor U5894 (N_5894,N_4815,N_3000);
nand U5895 (N_5895,N_1462,N_419);
xor U5896 (N_5896,N_3760,N_4071);
xor U5897 (N_5897,N_2375,N_3920);
or U5898 (N_5898,N_4785,N_908);
or U5899 (N_5899,N_3135,N_2946);
and U5900 (N_5900,N_2747,N_2616);
nand U5901 (N_5901,N_3077,N_625);
nor U5902 (N_5902,N_176,N_1807);
and U5903 (N_5903,N_4750,N_4980);
and U5904 (N_5904,N_3992,N_3013);
and U5905 (N_5905,N_3219,N_4196);
xnor U5906 (N_5906,N_1107,N_3578);
and U5907 (N_5907,N_3464,N_3422);
xnor U5908 (N_5908,N_3556,N_3396);
xnor U5909 (N_5909,N_596,N_4913);
nor U5910 (N_5910,N_3909,N_3529);
nor U5911 (N_5911,N_166,N_3517);
nor U5912 (N_5912,N_1915,N_799);
and U5913 (N_5913,N_2803,N_1793);
and U5914 (N_5914,N_2402,N_2587);
or U5915 (N_5915,N_1174,N_2154);
xor U5916 (N_5916,N_1374,N_2418);
or U5917 (N_5917,N_3085,N_4155);
xor U5918 (N_5918,N_624,N_3661);
xnor U5919 (N_5919,N_3423,N_3460);
nand U5920 (N_5920,N_2259,N_2840);
or U5921 (N_5921,N_1400,N_3704);
nand U5922 (N_5922,N_1720,N_4041);
or U5923 (N_5923,N_617,N_3050);
xor U5924 (N_5924,N_1764,N_1788);
or U5925 (N_5925,N_1841,N_4451);
nor U5926 (N_5926,N_3479,N_3293);
nand U5927 (N_5927,N_1697,N_4910);
nand U5928 (N_5928,N_2759,N_4804);
nand U5929 (N_5929,N_903,N_4486);
nor U5930 (N_5930,N_3023,N_4912);
xor U5931 (N_5931,N_3209,N_2951);
and U5932 (N_5932,N_4968,N_2056);
nand U5933 (N_5933,N_1872,N_4272);
or U5934 (N_5934,N_2179,N_1660);
or U5935 (N_5935,N_2241,N_1352);
and U5936 (N_5936,N_3406,N_3215);
nor U5937 (N_5937,N_2092,N_1754);
or U5938 (N_5938,N_645,N_2548);
xnor U5939 (N_5939,N_2146,N_1914);
or U5940 (N_5940,N_249,N_1670);
and U5941 (N_5941,N_2647,N_688);
or U5942 (N_5942,N_2856,N_2325);
xnor U5943 (N_5943,N_3270,N_492);
nor U5944 (N_5944,N_3106,N_2786);
or U5945 (N_5945,N_2490,N_4853);
nor U5946 (N_5946,N_4176,N_251);
and U5947 (N_5947,N_1177,N_4972);
or U5948 (N_5948,N_3603,N_3519);
nand U5949 (N_5949,N_2330,N_2640);
xnor U5950 (N_5950,N_2119,N_2973);
or U5951 (N_5951,N_1661,N_1304);
xnor U5952 (N_5952,N_3318,N_1153);
nor U5953 (N_5953,N_2681,N_2501);
nor U5954 (N_5954,N_4250,N_48);
or U5955 (N_5955,N_3057,N_3601);
nor U5956 (N_5956,N_1952,N_1730);
nor U5957 (N_5957,N_989,N_1652);
nor U5958 (N_5958,N_4019,N_716);
nand U5959 (N_5959,N_3315,N_1790);
nand U5960 (N_5960,N_763,N_840);
and U5961 (N_5961,N_1307,N_2517);
or U5962 (N_5962,N_4633,N_4698);
nor U5963 (N_5963,N_2934,N_708);
and U5964 (N_5964,N_605,N_2396);
and U5965 (N_5965,N_1600,N_1614);
and U5966 (N_5966,N_3573,N_4834);
nand U5967 (N_5967,N_4399,N_3059);
nor U5968 (N_5968,N_267,N_4873);
xor U5969 (N_5969,N_794,N_4618);
xnor U5970 (N_5970,N_55,N_2665);
nand U5971 (N_5971,N_1621,N_907);
nand U5972 (N_5972,N_689,N_1698);
or U5973 (N_5973,N_4501,N_2637);
nand U5974 (N_5974,N_3420,N_3833);
or U5975 (N_5975,N_2596,N_3713);
nand U5976 (N_5976,N_3976,N_1160);
and U5977 (N_5977,N_3906,N_1766);
or U5978 (N_5978,N_1850,N_4005);
and U5979 (N_5979,N_1437,N_883);
and U5980 (N_5980,N_2297,N_395);
xor U5981 (N_5981,N_3998,N_225);
or U5982 (N_5982,N_3333,N_1275);
or U5983 (N_5983,N_3851,N_2108);
and U5984 (N_5984,N_382,N_3754);
or U5985 (N_5985,N_4611,N_3074);
and U5986 (N_5986,N_2897,N_197);
or U5987 (N_5987,N_2385,N_2711);
and U5988 (N_5988,N_4671,N_565);
nor U5989 (N_5989,N_3352,N_1360);
and U5990 (N_5990,N_1081,N_3784);
xnor U5991 (N_5991,N_3060,N_1105);
nand U5992 (N_5992,N_4128,N_1316);
nand U5993 (N_5993,N_640,N_3314);
nor U5994 (N_5994,N_2430,N_1762);
xnor U5995 (N_5995,N_3904,N_3022);
or U5996 (N_5996,N_4760,N_156);
nand U5997 (N_5997,N_1503,N_4106);
nand U5998 (N_5998,N_855,N_528);
nand U5999 (N_5999,N_3691,N_3771);
and U6000 (N_6000,N_72,N_3249);
xor U6001 (N_6001,N_751,N_731);
and U6002 (N_6002,N_2559,N_667);
nand U6003 (N_6003,N_1318,N_784);
xor U6004 (N_6004,N_3570,N_1929);
nor U6005 (N_6005,N_3742,N_506);
xnor U6006 (N_6006,N_1320,N_4776);
xor U6007 (N_6007,N_3939,N_2750);
xnor U6008 (N_6008,N_4062,N_2227);
nor U6009 (N_6009,N_1507,N_4965);
and U6010 (N_6010,N_4592,N_1687);
or U6011 (N_6011,N_4173,N_4296);
nand U6012 (N_6012,N_1975,N_1662);
and U6013 (N_6013,N_3181,N_2990);
or U6014 (N_6014,N_3151,N_1144);
nor U6015 (N_6015,N_4166,N_4490);
xnor U6016 (N_6016,N_2052,N_2860);
nor U6017 (N_6017,N_3404,N_1582);
and U6018 (N_6018,N_3504,N_3118);
or U6019 (N_6019,N_4580,N_3822);
nor U6020 (N_6020,N_2534,N_4045);
or U6021 (N_6021,N_4242,N_4247);
xnor U6022 (N_6022,N_4473,N_3905);
nand U6023 (N_6023,N_3794,N_2801);
nor U6024 (N_6024,N_658,N_4270);
nand U6025 (N_6025,N_3706,N_259);
and U6026 (N_6026,N_2790,N_272);
nand U6027 (N_6027,N_4488,N_2693);
or U6028 (N_6028,N_3587,N_3574);
xnor U6029 (N_6029,N_2407,N_3966);
nor U6030 (N_6030,N_2689,N_1783);
or U6031 (N_6031,N_1596,N_1533);
and U6032 (N_6032,N_73,N_1395);
or U6033 (N_6033,N_586,N_1732);
nor U6034 (N_6034,N_1013,N_3326);
nand U6035 (N_6035,N_1060,N_3455);
and U6036 (N_6036,N_1422,N_1654);
or U6037 (N_6037,N_2493,N_573);
nor U6038 (N_6038,N_1620,N_1);
and U6039 (N_6039,N_3426,N_198);
and U6040 (N_6040,N_1252,N_805);
xnor U6041 (N_6041,N_3357,N_1341);
xor U6042 (N_6042,N_2825,N_3514);
nor U6043 (N_6043,N_3,N_4790);
or U6044 (N_6044,N_1328,N_3407);
or U6045 (N_6045,N_3205,N_1433);
or U6046 (N_6046,N_2222,N_3382);
nor U6047 (N_6047,N_2834,N_1895);
nor U6048 (N_6048,N_4736,N_4075);
xor U6049 (N_6049,N_4401,N_3338);
or U6050 (N_6050,N_623,N_3775);
or U6051 (N_6051,N_4456,N_2289);
nand U6052 (N_6052,N_2952,N_296);
and U6053 (N_6053,N_2518,N_508);
or U6054 (N_6054,N_2760,N_1194);
or U6055 (N_6055,N_3623,N_744);
nor U6056 (N_6056,N_4348,N_2022);
xor U6057 (N_6057,N_2169,N_2061);
or U6058 (N_6058,N_670,N_3098);
xor U6059 (N_6059,N_1777,N_183);
xnor U6060 (N_6060,N_566,N_4651);
nor U6061 (N_6061,N_1439,N_1011);
and U6062 (N_6062,N_2967,N_1242);
or U6063 (N_6063,N_1925,N_1024);
nor U6064 (N_6064,N_206,N_925);
or U6065 (N_6065,N_2682,N_1100);
nand U6066 (N_6066,N_56,N_4857);
nor U6067 (N_6067,N_286,N_1603);
xor U6068 (N_6068,N_3332,N_4316);
xnor U6069 (N_6069,N_1389,N_2819);
xnor U6070 (N_6070,N_373,N_2731);
nor U6071 (N_6071,N_1890,N_4595);
xnor U6072 (N_6072,N_3894,N_1122);
or U6073 (N_6073,N_1384,N_4907);
or U6074 (N_6074,N_884,N_2059);
xnor U6075 (N_6075,N_4182,N_4012);
and U6076 (N_6076,N_2879,N_2623);
or U6077 (N_6077,N_2393,N_355);
or U6078 (N_6078,N_64,N_3459);
nor U6079 (N_6079,N_2686,N_4878);
nor U6080 (N_6080,N_3006,N_4655);
and U6081 (N_6081,N_4931,N_0);
and U6082 (N_6082,N_3443,N_2419);
nand U6083 (N_6083,N_300,N_2546);
nand U6084 (N_6084,N_1425,N_3941);
nor U6085 (N_6085,N_4961,N_1308);
nand U6086 (N_6086,N_1635,N_2978);
nor U6087 (N_6087,N_2495,N_1417);
nor U6088 (N_6088,N_3637,N_4400);
or U6089 (N_6089,N_1086,N_1996);
nand U6090 (N_6090,N_4847,N_4349);
or U6091 (N_6091,N_2143,N_2358);
nor U6092 (N_6092,N_2101,N_2387);
nand U6093 (N_6093,N_4772,N_134);
nor U6094 (N_6094,N_3968,N_4127);
nand U6095 (N_6095,N_4073,N_2714);
or U6096 (N_6096,N_4937,N_1465);
and U6097 (N_6097,N_4064,N_4942);
or U6098 (N_6098,N_4946,N_3897);
or U6099 (N_6099,N_3862,N_3478);
nand U6100 (N_6100,N_3685,N_1459);
and U6101 (N_6101,N_212,N_2985);
or U6102 (N_6102,N_2367,N_3360);
and U6103 (N_6103,N_1515,N_1940);
nand U6104 (N_6104,N_2652,N_3565);
nor U6105 (N_6105,N_935,N_23);
xnor U6106 (N_6106,N_182,N_1287);
and U6107 (N_6107,N_4225,N_3129);
and U6108 (N_6108,N_1326,N_3497);
or U6109 (N_6109,N_3359,N_1206);
or U6110 (N_6110,N_1041,N_533);
nor U6111 (N_6111,N_1271,N_4191);
xnor U6112 (N_6112,N_4325,N_3702);
or U6113 (N_6113,N_913,N_2444);
and U6114 (N_6114,N_3109,N_4758);
nor U6115 (N_6115,N_4081,N_3392);
nor U6116 (N_6116,N_1280,N_4304);
nor U6117 (N_6117,N_3445,N_2307);
nand U6118 (N_6118,N_826,N_4945);
nand U6119 (N_6119,N_941,N_916);
nand U6120 (N_6120,N_2877,N_2795);
nand U6121 (N_6121,N_1187,N_2773);
nor U6122 (N_6122,N_4918,N_4831);
nor U6123 (N_6123,N_3582,N_4689);
and U6124 (N_6124,N_4970,N_3254);
xor U6125 (N_6125,N_2039,N_2177);
nor U6126 (N_6126,N_3647,N_897);
nor U6127 (N_6127,N_898,N_4814);
xor U6128 (N_6128,N_1054,N_4606);
and U6129 (N_6129,N_1419,N_3038);
nor U6130 (N_6130,N_844,N_30);
nor U6131 (N_6131,N_3590,N_4640);
nor U6132 (N_6132,N_2974,N_2544);
or U6133 (N_6133,N_4200,N_3743);
xnor U6134 (N_6134,N_3039,N_3058);
xnor U6135 (N_6135,N_3275,N_3295);
nand U6136 (N_6136,N_384,N_3804);
or U6137 (N_6137,N_3563,N_4554);
nor U6138 (N_6138,N_4156,N_4470);
and U6139 (N_6139,N_3123,N_2727);
nand U6140 (N_6140,N_2583,N_888);
xnor U6141 (N_6141,N_2349,N_3371);
or U6142 (N_6142,N_1297,N_3993);
and U6143 (N_6143,N_2505,N_1706);
nand U6144 (N_6144,N_1053,N_3699);
or U6145 (N_6145,N_4199,N_2166);
and U6146 (N_6146,N_3265,N_616);
nand U6147 (N_6147,N_4343,N_2287);
and U6148 (N_6148,N_4851,N_1792);
nand U6149 (N_6149,N_4408,N_4298);
xor U6150 (N_6150,N_3936,N_1960);
nor U6151 (N_6151,N_1163,N_4461);
nand U6152 (N_6152,N_2982,N_589);
or U6153 (N_6153,N_122,N_1442);
nand U6154 (N_6154,N_788,N_3918);
xnor U6155 (N_6155,N_2463,N_3207);
and U6156 (N_6156,N_4835,N_1763);
xor U6157 (N_6157,N_964,N_3483);
nand U6158 (N_6158,N_2820,N_4376);
and U6159 (N_6159,N_4464,N_3963);
or U6160 (N_6160,N_3068,N_3425);
and U6161 (N_6161,N_4663,N_1396);
nand U6162 (N_6162,N_3141,N_1347);
nor U6163 (N_6163,N_4365,N_885);
nor U6164 (N_6164,N_863,N_2861);
nor U6165 (N_6165,N_276,N_3257);
or U6166 (N_6166,N_3400,N_3933);
and U6167 (N_6167,N_2806,N_2303);
nand U6168 (N_6168,N_2176,N_3610);
or U6169 (N_6169,N_3847,N_4458);
or U6170 (N_6170,N_4704,N_1113);
xnor U6171 (N_6171,N_3014,N_3067);
and U6172 (N_6172,N_3378,N_3697);
nor U6173 (N_6173,N_2841,N_1638);
nand U6174 (N_6174,N_1640,N_1093);
nor U6175 (N_6175,N_818,N_558);
nor U6176 (N_6176,N_3337,N_929);
or U6177 (N_6177,N_4717,N_4310);
nor U6178 (N_6178,N_4359,N_1082);
xnor U6179 (N_6179,N_3274,N_3502);
xor U6180 (N_6180,N_801,N_236);
nand U6181 (N_6181,N_80,N_447);
and U6182 (N_6182,N_1281,N_1921);
nor U6183 (N_6183,N_3138,N_155);
xnor U6184 (N_6184,N_2549,N_902);
nor U6185 (N_6185,N_81,N_482);
and U6186 (N_6186,N_2865,N_341);
xor U6187 (N_6187,N_2696,N_737);
xor U6188 (N_6188,N_2298,N_1629);
xor U6189 (N_6189,N_2613,N_4255);
and U6190 (N_6190,N_1414,N_4485);
nand U6191 (N_6191,N_4768,N_205);
nand U6192 (N_6192,N_2771,N_2368);
and U6193 (N_6193,N_2450,N_2182);
or U6194 (N_6194,N_4792,N_2479);
nand U6195 (N_6195,N_1607,N_3122);
or U6196 (N_6196,N_1017,N_4030);
xor U6197 (N_6197,N_4098,N_25);
or U6198 (N_6198,N_1800,N_2060);
nor U6199 (N_6199,N_3063,N_1789);
and U6200 (N_6200,N_4593,N_4738);
or U6201 (N_6201,N_3166,N_381);
and U6202 (N_6202,N_4188,N_2115);
nand U6203 (N_6203,N_968,N_517);
nand U6204 (N_6204,N_472,N_3953);
nor U6205 (N_6205,N_4362,N_3139);
and U6206 (N_6206,N_168,N_824);
nor U6207 (N_6207,N_3614,N_4228);
xor U6208 (N_6208,N_17,N_4350);
and U6209 (N_6209,N_1274,N_245);
and U6210 (N_6210,N_1878,N_4969);
and U6211 (N_6211,N_4232,N_3929);
or U6212 (N_6212,N_457,N_4775);
nand U6213 (N_6213,N_2328,N_4639);
or U6214 (N_6214,N_2138,N_4647);
xor U6215 (N_6215,N_3021,N_3499);
or U6216 (N_6216,N_1034,N_3981);
and U6217 (N_6217,N_2893,N_4427);
nor U6218 (N_6218,N_4457,N_4453);
nand U6219 (N_6219,N_4516,N_248);
or U6220 (N_6220,N_2707,N_3815);
and U6221 (N_6221,N_1811,N_4141);
nor U6222 (N_6222,N_673,N_3212);
and U6223 (N_6223,N_1602,N_4602);
or U6224 (N_6224,N_4428,N_4137);
nor U6225 (N_6225,N_1986,N_800);
xor U6226 (N_6226,N_4881,N_4690);
nand U6227 (N_6227,N_3143,N_292);
and U6228 (N_6228,N_2131,N_4986);
or U6229 (N_6229,N_1505,N_4594);
nor U6230 (N_6230,N_1140,N_161);
or U6231 (N_6231,N_3346,N_3778);
xnor U6232 (N_6232,N_3753,N_1370);
or U6233 (N_6233,N_704,N_2606);
and U6234 (N_6234,N_1379,N_3688);
and U6235 (N_6235,N_4057,N_4828);
nand U6236 (N_6236,N_3017,N_4922);
xnor U6237 (N_6237,N_1112,N_757);
nand U6238 (N_6238,N_233,N_1508);
xnor U6239 (N_6239,N_2436,N_1496);
or U6240 (N_6240,N_4759,N_2140);
and U6241 (N_6241,N_2439,N_2429);
xor U6242 (N_6242,N_3462,N_1684);
or U6243 (N_6243,N_2654,N_4536);
nand U6244 (N_6244,N_307,N_4546);
and U6245 (N_6245,N_1228,N_4797);
xor U6246 (N_6246,N_3402,N_735);
xor U6247 (N_6247,N_4515,N_3276);
nand U6248 (N_6248,N_2624,N_1989);
and U6249 (N_6249,N_4163,N_2246);
and U6250 (N_6250,N_1726,N_2928);
and U6251 (N_6251,N_2007,N_434);
and U6252 (N_6252,N_335,N_3498);
nand U6253 (N_6253,N_3898,N_1954);
nand U6254 (N_6254,N_148,N_723);
nand U6255 (N_6255,N_4056,N_4389);
or U6256 (N_6256,N_4165,N_4973);
and U6257 (N_6257,N_802,N_1595);
and U6258 (N_6258,N_1430,N_304);
nor U6259 (N_6259,N_323,N_4069);
and U6260 (N_6260,N_1210,N_435);
nand U6261 (N_6261,N_1880,N_4997);
and U6262 (N_6262,N_1927,N_138);
and U6263 (N_6263,N_2198,N_4326);
nand U6264 (N_6264,N_2477,N_1864);
and U6265 (N_6265,N_4762,N_1257);
or U6266 (N_6266,N_69,N_766);
nand U6267 (N_6267,N_4021,N_4132);
nor U6268 (N_6268,N_2520,N_187);
nand U6269 (N_6269,N_1545,N_2763);
or U6270 (N_6270,N_544,N_2400);
or U6271 (N_6271,N_3681,N_1248);
nor U6272 (N_6272,N_3666,N_3728);
xor U6273 (N_6273,N_4575,N_3472);
or U6274 (N_6274,N_3336,N_1329);
nand U6275 (N_6275,N_2045,N_1889);
and U6276 (N_6276,N_2617,N_1335);
or U6277 (N_6277,N_1886,N_2533);
xnor U6278 (N_6278,N_620,N_3186);
nand U6279 (N_6279,N_2631,N_2845);
xnor U6280 (N_6280,N_1672,N_4101);
nor U6281 (N_6281,N_2442,N_950);
nor U6282 (N_6282,N_1559,N_1562);
nand U6283 (N_6283,N_2296,N_4879);
and U6284 (N_6284,N_4145,N_4533);
nand U6285 (N_6285,N_4787,N_4645);
nand U6286 (N_6286,N_2835,N_777);
nor U6287 (N_6287,N_146,N_2256);
xnor U6288 (N_6288,N_4053,N_150);
xor U6289 (N_6289,N_3133,N_4659);
nand U6290 (N_6290,N_4621,N_500);
or U6291 (N_6291,N_488,N_1795);
or U6292 (N_6292,N_3418,N_4087);
or U6293 (N_6293,N_3173,N_4092);
or U6294 (N_6294,N_1255,N_4341);
xor U6295 (N_6295,N_4063,N_955);
and U6296 (N_6296,N_2423,N_208);
or U6297 (N_6297,N_3608,N_4146);
and U6298 (N_6298,N_1208,N_2831);
and U6299 (N_6299,N_112,N_4871);
xor U6300 (N_6300,N_4194,N_3724);
or U6301 (N_6301,N_614,N_2971);
xor U6302 (N_6302,N_2769,N_2844);
nor U6303 (N_6303,N_3746,N_131);
nor U6304 (N_6304,N_4628,N_180);
and U6305 (N_6305,N_4286,N_3399);
nor U6306 (N_6306,N_3349,N_1615);
or U6307 (N_6307,N_3576,N_1342);
nor U6308 (N_6308,N_1506,N_2381);
nor U6309 (N_6309,N_2874,N_2254);
and U6310 (N_6310,N_849,N_632);
nor U6311 (N_6311,N_4483,N_3277);
nand U6312 (N_6312,N_2867,N_4068);
nor U6313 (N_6313,N_1771,N_4764);
nand U6314 (N_6314,N_4111,N_3285);
xor U6315 (N_6315,N_3552,N_3756);
nand U6316 (N_6316,N_1676,N_4253);
or U6317 (N_6317,N_4066,N_1057);
or U6318 (N_6318,N_4434,N_4683);
xor U6319 (N_6319,N_2894,N_2345);
nand U6320 (N_6320,N_3534,N_3597);
xnor U6321 (N_6321,N_1126,N_2745);
nand U6322 (N_6322,N_1004,N_1679);
or U6323 (N_6323,N_2561,N_4799);
xnor U6324 (N_6324,N_446,N_4300);
or U6325 (N_6325,N_4820,N_1632);
or U6326 (N_6326,N_1074,N_2872);
nor U6327 (N_6327,N_2121,N_3980);
and U6328 (N_6328,N_550,N_1825);
xnor U6329 (N_6329,N_2023,N_137);
xor U6330 (N_6330,N_1036,N_553);
and U6331 (N_6331,N_3051,N_2576);
nor U6332 (N_6332,N_4149,N_2642);
xnor U6333 (N_6333,N_4866,N_2351);
and U6334 (N_6334,N_1117,N_2619);
and U6335 (N_6335,N_3566,N_3696);
nor U6336 (N_6336,N_228,N_2680);
xnor U6337 (N_6337,N_2913,N_1835);
or U6338 (N_6338,N_383,N_232);
xnor U6339 (N_6339,N_3683,N_2471);
nor U6340 (N_6340,N_204,N_4424);
and U6341 (N_6341,N_503,N_3785);
xor U6342 (N_6342,N_2397,N_1743);
nand U6343 (N_6343,N_2126,N_2041);
xnor U6344 (N_6344,N_3871,N_2235);
nor U6345 (N_6345,N_1078,N_1077);
nand U6346 (N_6346,N_1578,N_4691);
and U6347 (N_6347,N_1334,N_934);
and U6348 (N_6348,N_776,N_768);
nor U6349 (N_6349,N_408,N_160);
xnor U6350 (N_6350,N_4577,N_1575);
nor U6351 (N_6351,N_1934,N_3493);
nand U6352 (N_6352,N_3362,N_3363);
nand U6353 (N_6353,N_1296,N_3773);
and U6354 (N_6354,N_1585,N_2197);
or U6355 (N_6355,N_1317,N_379);
nand U6356 (N_6356,N_793,N_293);
or U6357 (N_6357,N_377,N_3679);
and U6358 (N_6358,N_4719,N_4906);
or U6359 (N_6359,N_3770,N_3864);
and U6360 (N_6360,N_4079,N_1489);
xnor U6361 (N_6361,N_2082,N_4687);
xnor U6362 (N_6362,N_2924,N_4269);
and U6363 (N_6363,N_536,N_4497);
or U6364 (N_6364,N_979,N_3369);
xnor U6365 (N_6365,N_856,N_4139);
nand U6366 (N_6366,N_1573,N_4579);
nor U6367 (N_6367,N_4783,N_4779);
nor U6368 (N_6368,N_40,N_1239);
nor U6369 (N_6369,N_2556,N_1922);
nand U6370 (N_6370,N_3071,N_402);
and U6371 (N_6371,N_1293,N_1311);
and U6372 (N_6372,N_1570,N_2318);
xnor U6373 (N_6373,N_1150,N_4908);
and U6374 (N_6374,N_2129,N_3233);
and U6375 (N_6375,N_3442,N_1941);
nand U6376 (N_6376,N_4553,N_871);
xnor U6377 (N_6377,N_1541,N_57);
and U6378 (N_6378,N_1212,N_676);
or U6379 (N_6379,N_4442,N_1871);
nand U6380 (N_6380,N_741,N_2761);
nor U6381 (N_6381,N_785,N_2811);
xor U6382 (N_6382,N_4504,N_4500);
nand U6383 (N_6383,N_4159,N_2354);
nor U6384 (N_6384,N_621,N_1164);
or U6385 (N_6385,N_211,N_19);
and U6386 (N_6386,N_3227,N_365);
or U6387 (N_6387,N_2278,N_1012);
xnor U6388 (N_6388,N_1458,N_4743);
or U6389 (N_6389,N_1138,N_739);
nand U6390 (N_6390,N_2097,N_3886);
or U6391 (N_6391,N_790,N_47);
and U6392 (N_6392,N_4526,N_2570);
nor U6393 (N_6393,N_1542,N_1322);
or U6394 (N_6394,N_1584,N_1127);
or U6395 (N_6395,N_1009,N_4927);
xor U6396 (N_6396,N_582,N_3913);
or U6397 (N_6397,N_2168,N_2132);
or U6398 (N_6398,N_2547,N_4020);
and U6399 (N_6399,N_2295,N_2935);
nor U6400 (N_6400,N_2134,N_1742);
nand U6401 (N_6401,N_1540,N_4947);
nand U6402 (N_6402,N_820,N_1118);
xnor U6403 (N_6403,N_1198,N_1782);
or U6404 (N_6404,N_219,N_4544);
and U6405 (N_6405,N_4545,N_4203);
and U6406 (N_6406,N_3525,N_1812);
or U6407 (N_6407,N_191,N_4116);
and U6408 (N_6408,N_1485,N_975);
nand U6409 (N_6409,N_2238,N_1276);
nor U6410 (N_6410,N_3453,N_2792);
and U6411 (N_6411,N_2940,N_3244);
nand U6412 (N_6412,N_265,N_2942);
xnor U6413 (N_6413,N_2310,N_2580);
nand U6414 (N_6414,N_480,N_1155);
nand U6415 (N_6415,N_630,N_1445);
xnor U6416 (N_6416,N_1810,N_2455);
nand U6417 (N_6417,N_3052,N_724);
or U6418 (N_6418,N_107,N_2925);
nand U6419 (N_6419,N_4382,N_4211);
xor U6420 (N_6420,N_627,N_2313);
or U6421 (N_6421,N_792,N_3721);
or U6422 (N_6422,N_3723,N_4709);
xnor U6423 (N_6423,N_3912,N_1359);
nor U6424 (N_6424,N_4748,N_4198);
or U6425 (N_6425,N_2917,N_1464);
xor U6426 (N_6426,N_2692,N_2245);
nor U6427 (N_6427,N_3232,N_1469);
and U6428 (N_6428,N_521,N_170);
xnor U6429 (N_6429,N_987,N_350);
nand U6430 (N_6430,N_3767,N_1688);
or U6431 (N_6431,N_4151,N_2240);
nor U6432 (N_6432,N_2151,N_3985);
nand U6433 (N_6433,N_1434,N_4838);
and U6434 (N_6434,N_2366,N_240);
nand U6435 (N_6435,N_4378,N_301);
nand U6436 (N_6436,N_2909,N_3340);
nand U6437 (N_6437,N_1109,N_1084);
nor U6438 (N_6438,N_4037,N_167);
xnor U6439 (N_6439,N_4723,N_1223);
xor U6440 (N_6440,N_196,N_2147);
xnor U6441 (N_6441,N_2697,N_3911);
nand U6442 (N_6442,N_1714,N_4134);
or U6443 (N_6443,N_4573,N_4824);
nor U6444 (N_6444,N_1949,N_26);
or U6445 (N_6445,N_1972,N_2483);
and U6446 (N_6446,N_1350,N_1277);
nand U6447 (N_6447,N_4751,N_3653);
nor U6448 (N_6448,N_2102,N_4967);
and U6449 (N_6449,N_1898,N_3644);
nand U6450 (N_6450,N_2742,N_3341);
or U6451 (N_6451,N_4675,N_415);
nor U6452 (N_6452,N_4243,N_4153);
and U6453 (N_6453,N_1944,N_954);
and U6454 (N_6454,N_3611,N_256);
or U6455 (N_6455,N_3823,N_4216);
nor U6456 (N_6456,N_4122,N_3288);
xnor U6457 (N_6457,N_2413,N_3292);
and U6458 (N_6458,N_1689,N_1258);
or U6459 (N_6459,N_685,N_3160);
or U6460 (N_6460,N_3555,N_1175);
and U6461 (N_6461,N_2915,N_2162);
nor U6462 (N_6462,N_539,N_3972);
and U6463 (N_6463,N_3673,N_2632);
nor U6464 (N_6464,N_3645,N_1574);
nand U6465 (N_6465,N_1412,N_2164);
xnor U6466 (N_6466,N_1806,N_2797);
nand U6467 (N_6467,N_3744,N_2630);
xor U6468 (N_6468,N_3648,N_4179);
or U6469 (N_6469,N_451,N_2331);
and U6470 (N_6470,N_1799,N_1211);
nor U6471 (N_6471,N_752,N_2193);
nor U6472 (N_6472,N_730,N_3615);
xor U6473 (N_6473,N_3538,N_3440);
or U6474 (N_6474,N_684,N_209);
nand U6475 (N_6475,N_2813,N_3546);
xnor U6476 (N_6476,N_2212,N_3241);
nand U6477 (N_6477,N_4431,N_4197);
and U6478 (N_6478,N_1623,N_1378);
and U6479 (N_6479,N_2267,N_2341);
or U6480 (N_6480,N_1641,N_2661);
xnor U6481 (N_6481,N_1222,N_1536);
nor U6482 (N_6482,N_1590,N_3165);
nand U6483 (N_6483,N_151,N_3875);
and U6484 (N_6484,N_2220,N_4324);
and U6485 (N_6485,N_1673,N_2317);
xnor U6486 (N_6486,N_1197,N_2726);
xnor U6487 (N_6487,N_1857,N_1858);
xnor U6488 (N_6488,N_3485,N_1822);
or U6489 (N_6489,N_4911,N_3347);
or U6490 (N_6490,N_3531,N_1755);
or U6491 (N_6491,N_4774,N_3495);
or U6492 (N_6492,N_2626,N_1099);
nand U6493 (N_6493,N_4058,N_3054);
or U6494 (N_6494,N_4548,N_3290);
nor U6495 (N_6495,N_4528,N_2738);
or U6496 (N_6496,N_1525,N_3066);
and U6497 (N_6497,N_20,N_728);
or U6498 (N_6498,N_1998,N_3633);
nand U6499 (N_6499,N_2425,N_3740);
or U6500 (N_6500,N_3334,N_812);
nand U6501 (N_6501,N_366,N_2660);
or U6502 (N_6502,N_3551,N_599);
or U6503 (N_6503,N_4468,N_2565);
nand U6504 (N_6504,N_4601,N_1478);
xor U6505 (N_6505,N_798,N_3170);
nand U6506 (N_6506,N_3007,N_2262);
and U6507 (N_6507,N_3037,N_7);
xnor U6508 (N_6508,N_4688,N_4441);
or U6509 (N_6509,N_2814,N_2753);
nand U6510 (N_6510,N_3439,N_552);
and U6511 (N_6511,N_762,N_791);
or U6512 (N_6512,N_4916,N_1463);
and U6513 (N_6513,N_3750,N_4721);
nor U6514 (N_6514,N_1891,N_4360);
xnor U6515 (N_6515,N_4007,N_3725);
or U6516 (N_6516,N_2746,N_1440);
nand U6517 (N_6517,N_1225,N_2221);
and U6518 (N_6518,N_1955,N_4599);
nand U6519 (N_6519,N_3430,N_2988);
xor U6520 (N_6520,N_1005,N_4564);
nor U6521 (N_6521,N_3946,N_948);
nand U6522 (N_6522,N_3243,N_1479);
or U6523 (N_6523,N_1353,N_450);
or U6524 (N_6524,N_938,N_1032);
nand U6525 (N_6525,N_4186,N_1674);
nor U6526 (N_6526,N_4065,N_660);
nor U6527 (N_6527,N_2775,N_2725);
nor U6528 (N_6528,N_2050,N_3131);
nand U6529 (N_6529,N_268,N_3718);
and U6530 (N_6530,N_4138,N_3383);
nand U6531 (N_6531,N_3114,N_1750);
xor U6532 (N_6532,N_2836,N_2904);
and U6533 (N_6533,N_3777,N_4604);
xor U6534 (N_6534,N_364,N_3893);
nand U6535 (N_6535,N_1594,N_2944);
and U6536 (N_6536,N_1214,N_719);
and U6537 (N_6537,N_3432,N_2685);
nand U6538 (N_6538,N_50,N_4419);
nand U6539 (N_6539,N_4634,N_2723);
and U6540 (N_6540,N_2569,N_2550);
or U6541 (N_6541,N_27,N_169);
xnor U6542 (N_6542,N_641,N_193);
nand U6543 (N_6543,N_4981,N_2170);
and U6544 (N_6544,N_901,N_1111);
or U6545 (N_6545,N_700,N_4417);
nand U6546 (N_6546,N_1686,N_3134);
and U6547 (N_6547,N_4314,N_317);
nor U6548 (N_6548,N_1278,N_4884);
and U6549 (N_6549,N_4679,N_3693);
nand U6550 (N_6550,N_1942,N_4855);
or U6551 (N_6551,N_3670,N_1040);
nand U6552 (N_6552,N_4513,N_2327);
and U6553 (N_6553,N_1207,N_36);
xor U6554 (N_6554,N_1978,N_2384);
and U6555 (N_6555,N_2284,N_4379);
or U6556 (N_6556,N_633,N_3012);
nand U6557 (N_6557,N_3631,N_3952);
nand U6558 (N_6558,N_262,N_3208);
or U6559 (N_6559,N_655,N_4383);
nor U6560 (N_6560,N_4538,N_2096);
nor U6561 (N_6561,N_609,N_1905);
and U6562 (N_6562,N_4220,N_703);
or U6563 (N_6563,N_4105,N_3221);
xor U6564 (N_6564,N_3989,N_1209);
xor U6565 (N_6565,N_3046,N_4202);
nor U6566 (N_6566,N_3387,N_828);
nand U6567 (N_6567,N_1499,N_804);
xnor U6568 (N_6568,N_3456,N_3210);
and U6569 (N_6569,N_2979,N_2886);
xnor U6570 (N_6570,N_829,N_1604);
xnor U6571 (N_6571,N_551,N_2046);
xnor U6572 (N_6572,N_1351,N_3545);
or U6573 (N_6573,N_2992,N_3824);
nand U6574 (N_6574,N_271,N_2432);
or U6575 (N_6575,N_3032,N_2300);
and U6576 (N_6576,N_4119,N_427);
nor U6577 (N_6577,N_644,N_3465);
or U6578 (N_6578,N_549,N_4115);
nor U6579 (N_6579,N_4172,N_363);
nand U6580 (N_6580,N_1493,N_3714);
or U6581 (N_6581,N_1566,N_3329);
nor U6582 (N_6582,N_2705,N_1473);
xnor U6583 (N_6583,N_2945,N_1191);
xor U6584 (N_6584,N_2128,N_496);
nor U6585 (N_6585,N_342,N_2829);
and U6586 (N_6586,N_1446,N_2035);
nor U6587 (N_6587,N_4649,N_3731);
nand U6588 (N_6588,N_779,N_1826);
nand U6589 (N_6589,N_3335,N_3289);
nand U6590 (N_6590,N_4209,N_1408);
and U6591 (N_6591,N_2539,N_4956);
nand U6592 (N_6592,N_3003,N_2095);
xor U6593 (N_6593,N_4854,N_120);
nor U6594 (N_6594,N_29,N_2832);
or U6595 (N_6595,N_4014,N_3447);
and U6596 (N_6596,N_1504,N_2421);
and U6597 (N_6597,N_3880,N_4529);
nand U6598 (N_6598,N_2507,N_3238);
nand U6599 (N_6599,N_4650,N_4217);
and U6600 (N_6600,N_2634,N_628);
xor U6601 (N_6601,N_2020,N_28);
and U6602 (N_6602,N_3974,N_1936);
xor U6603 (N_6603,N_4330,N_4085);
or U6604 (N_6604,N_2269,N_758);
and U6605 (N_6605,N_2620,N_4396);
or U6606 (N_6606,N_2573,N_3798);
nor U6607 (N_6607,N_3795,N_4301);
and U6608 (N_6608,N_479,N_3294);
xor U6609 (N_6609,N_870,N_721);
or U6610 (N_6610,N_2320,N_4540);
nor U6611 (N_6611,N_2496,N_1995);
or U6612 (N_6612,N_1608,N_3802);
nor U6613 (N_6613,N_3889,N_4340);
nor U6614 (N_6614,N_2943,N_266);
nor U6615 (N_6615,N_2251,N_843);
nor U6616 (N_6616,N_1855,N_2058);
nand U6617 (N_6617,N_2214,N_3887);
or U6618 (N_6618,N_1867,N_3924);
and U6619 (N_6619,N_2447,N_1902);
and U6620 (N_6620,N_2519,N_1046);
or U6621 (N_6621,N_1923,N_1957);
or U6622 (N_6622,N_4446,N_144);
xor U6623 (N_6623,N_1298,N_531);
or U6624 (N_6624,N_1237,N_357);
nor U6625 (N_6625,N_3339,N_2414);
and U6626 (N_6626,N_3828,N_1102);
or U6627 (N_6627,N_1259,N_4523);
nand U6628 (N_6628,N_202,N_65);
and U6629 (N_6629,N_4710,N_4672);
xnor U6630 (N_6630,N_853,N_4025);
nor U6631 (N_6631,N_142,N_900);
nor U6632 (N_6632,N_1977,N_976);
or U6633 (N_6633,N_709,N_3419);
and U6634 (N_6634,N_4872,N_349);
or U6635 (N_6635,N_3624,N_4462);
nor U6636 (N_6636,N_2984,N_147);
nor U6637 (N_6637,N_3605,N_2555);
and U6638 (N_6638,N_1375,N_3808);
and U6639 (N_6639,N_815,N_2963);
xnor U6640 (N_6640,N_965,N_1747);
nor U6641 (N_6641,N_3388,N_2666);
nand U6642 (N_6642,N_331,N_3606);
nand U6643 (N_6643,N_3042,N_3044);
xnor U6644 (N_6644,N_186,N_991);
xor U6645 (N_6645,N_3902,N_866);
or U6646 (N_6646,N_2452,N_3281);
or U6647 (N_6647,N_3919,N_1094);
nand U6648 (N_6648,N_825,N_4433);
or U6649 (N_6649,N_1868,N_1310);
nor U6650 (N_6650,N_2229,N_4309);
nand U6651 (N_6651,N_3628,N_1869);
xor U6652 (N_6652,N_504,N_1529);
xor U6653 (N_6653,N_2271,N_2950);
nand U6654 (N_6654,N_3409,N_4077);
or U6655 (N_6655,N_2881,N_1367);
and U6656 (N_6656,N_3287,N_4763);
xnor U6657 (N_6657,N_4052,N_2752);
xnor U6658 (N_6658,N_4384,N_912);
or U6659 (N_6659,N_1456,N_1244);
nor U6660 (N_6660,N_4409,N_713);
or U6661 (N_6661,N_2857,N_3561);
or U6662 (N_6662,N_4475,N_3513);
nand U6663 (N_6663,N_3622,N_904);
and U6664 (N_6664,N_4142,N_1885);
nor U6665 (N_6665,N_171,N_2001);
xnor U6666 (N_6666,N_1729,N_2218);
nand U6667 (N_6667,N_464,N_3639);
or U6668 (N_6668,N_401,N_4454);
nor U6669 (N_6669,N_4334,N_1675);
nand U6670 (N_6670,N_2937,N_4027);
or U6671 (N_6671,N_875,N_2645);
nor U6672 (N_6672,N_478,N_3626);
and U6673 (N_6673,N_1470,N_118);
xor U6674 (N_6674,N_1775,N_3178);
nand U6675 (N_6675,N_1569,N_94);
nor U6676 (N_6676,N_1345,N_2592);
nand U6677 (N_6677,N_862,N_3838);
xnor U6678 (N_6678,N_100,N_3190);
xnor U6679 (N_6679,N_1598,N_3091);
or U6680 (N_6680,N_1145,N_598);
and U6681 (N_6681,N_2695,N_857);
or U6682 (N_6682,N_4036,N_1152);
xor U6683 (N_6683,N_1294,N_3540);
and U6684 (N_6684,N_2075,N_3161);
xnor U6685 (N_6685,N_4644,N_4777);
nand U6686 (N_6686,N_1741,N_990);
or U6687 (N_6687,N_2983,N_172);
and U6688 (N_6688,N_4080,N_4284);
nor U6689 (N_6689,N_3814,N_110);
and U6690 (N_6690,N_443,N_444);
or U6691 (N_6691,N_143,N_4638);
nand U6692 (N_6692,N_656,N_1557);
or U6693 (N_6693,N_4158,N_2406);
and U6694 (N_6694,N_1968,N_1522);
nand U6695 (N_6695,N_1537,N_3816);
or U6696 (N_6696,N_1466,N_2920);
nand U6697 (N_6697,N_95,N_2536);
nand U6698 (N_6698,N_2799,N_3986);
and U6699 (N_6699,N_1863,N_542);
nand U6700 (N_6700,N_626,N_4983);
nand U6701 (N_6701,N_4572,N_3395);
nand U6702 (N_6702,N_2776,N_3301);
and U6703 (N_6703,N_391,N_1832);
xnor U6704 (N_6704,N_2344,N_1719);
nand U6705 (N_6705,N_1501,N_3562);
and U6706 (N_6706,N_4305,N_279);
and U6707 (N_6707,N_2558,N_3535);
or U6708 (N_6708,N_2244,N_2817);
nand U6709 (N_6709,N_141,N_1913);
and U6710 (N_6710,N_4754,N_2883);
xnor U6711 (N_6711,N_121,N_1683);
and U6712 (N_6712,N_3954,N_3928);
nand U6713 (N_6713,N_458,N_175);
nand U6714 (N_6714,N_1365,N_67);
xnor U6715 (N_6715,N_4885,N_4443);
and U6716 (N_6716,N_3272,N_1778);
nor U6717 (N_6717,N_4494,N_1631);
xor U6718 (N_6718,N_2958,N_2422);
nand U6719 (N_6719,N_3211,N_136);
or U6720 (N_6720,N_4535,N_425);
and U6721 (N_6721,N_4781,N_1622);
or U6722 (N_6722,N_3145,N_3716);
or U6723 (N_6723,N_4123,N_3553);
nand U6724 (N_6724,N_3234,N_2461);
and U6725 (N_6725,N_1780,N_4195);
xor U6726 (N_6726,N_4686,N_698);
nand U6727 (N_6727,N_3544,N_2062);
and U6728 (N_6728,N_3829,N_3194);
and U6729 (N_6729,N_2503,N_3214);
nor U6730 (N_6730,N_1988,N_1587);
or U6731 (N_6731,N_4823,N_3668);
nand U6732 (N_6732,N_4047,N_3389);
and U6733 (N_6733,N_2098,N_2659);
or U6734 (N_6734,N_2995,N_4725);
and U6735 (N_6735,N_748,N_2489);
and U6736 (N_6736,N_4292,N_2643);
xnor U6737 (N_6737,N_4463,N_2026);
or U6738 (N_6738,N_1409,N_2441);
and U6739 (N_6739,N_2362,N_3641);
or U6740 (N_6740,N_878,N_2568);
nand U6741 (N_6741,N_577,N_3996);
nor U6742 (N_6742,N_2202,N_2506);
nand U6743 (N_6743,N_2263,N_4235);
nand U6744 (N_6744,N_3738,N_502);
nand U6745 (N_6745,N_2090,N_683);
nor U6746 (N_6746,N_4503,N_1565);
and U6747 (N_6747,N_2586,N_1544);
or U6748 (N_6748,N_3096,N_2870);
and U6749 (N_6749,N_3297,N_3496);
xor U6750 (N_6750,N_3855,N_360);
and U6751 (N_6751,N_946,N_2699);
nor U6752 (N_6752,N_1071,N_1659);
nand U6753 (N_6753,N_3598,N_4747);
nand U6754 (N_6754,N_426,N_1405);
and U6755 (N_6755,N_3759,N_4641);
nand U6756 (N_6756,N_3125,N_2712);
and U6757 (N_6757,N_405,N_459);
nand U6758 (N_6758,N_3745,N_270);
xnor U6759 (N_6759,N_4374,N_4204);
or U6760 (N_6760,N_2360,N_4524);
or U6761 (N_6761,N_956,N_4);
xnor U6762 (N_6762,N_4991,N_1634);
and U6763 (N_6763,N_4249,N_2277);
nor U6764 (N_6764,N_881,N_3863);
nand U6765 (N_6765,N_106,N_1381);
nor U6766 (N_6766,N_1182,N_1894);
nand U6767 (N_6767,N_2584,N_2516);
nand U6768 (N_6768,N_3198,N_1270);
nand U6769 (N_6769,N_2087,N_3617);
xor U6770 (N_6770,N_4631,N_2006);
xor U6771 (N_6771,N_1616,N_3762);
and U6772 (N_6772,N_2537,N_3353);
nor U6773 (N_6773,N_3260,N_2532);
nand U6774 (N_6774,N_4559,N_2099);
xnor U6775 (N_6775,N_1834,N_2578);
nand U6776 (N_6776,N_2864,N_3019);
and U6777 (N_6777,N_2017,N_2377);
nor U6778 (N_6778,N_3832,N_4782);
nor U6779 (N_6779,N_3618,N_3416);
or U6780 (N_6780,N_707,N_4212);
xnor U6781 (N_6781,N_2980,N_3640);
and U6782 (N_6782,N_3119,N_2038);
or U6783 (N_6783,N_1773,N_1132);
nand U6784 (N_6784,N_3755,N_3835);
xor U6785 (N_6785,N_2657,N_2701);
nor U6786 (N_6786,N_35,N_3302);
xor U6787 (N_6787,N_2389,N_4849);
nand U6788 (N_6788,N_2077,N_1302);
nand U6789 (N_6789,N_3328,N_3772);
nand U6790 (N_6790,N_514,N_3515);
nand U6791 (N_6791,N_1477,N_4733);
or U6792 (N_6792,N_2538,N_691);
or U6793 (N_6793,N_1824,N_1715);
nand U6794 (N_6794,N_4283,N_4895);
and U6795 (N_6795,N_1774,N_4842);
xnor U6796 (N_6796,N_303,N_1236);
xor U6797 (N_6797,N_931,N_3188);
xor U6798 (N_6798,N_3837,N_3408);
nor U6799 (N_6799,N_2818,N_1066);
nor U6800 (N_6800,N_4711,N_1881);
nand U6801 (N_6801,N_639,N_2301);
xnor U6802 (N_6802,N_3159,N_345);
nor U6803 (N_6803,N_4558,N_4880);
nand U6804 (N_6804,N_525,N_4390);
or U6805 (N_6805,N_2849,N_3199);
xnor U6806 (N_6806,N_4699,N_555);
nor U6807 (N_6807,N_4015,N_4600);
nor U6808 (N_6808,N_1691,N_119);
and U6809 (N_6809,N_3251,N_4557);
or U6810 (N_6810,N_732,N_139);
and U6811 (N_6811,N_1918,N_2474);
or U6812 (N_6812,N_603,N_1748);
xor U6813 (N_6813,N_1487,N_2456);
and U6814 (N_6814,N_3559,N_981);
or U6815 (N_6815,N_3732,N_2566);
nor U6816 (N_6816,N_1692,N_2275);
nor U6817 (N_6817,N_3094,N_4335);
and U6818 (N_6818,N_4730,N_2308);
nand U6819 (N_6819,N_3126,N_3967);
or U6820 (N_6820,N_1642,N_4403);
nand U6821 (N_6821,N_2782,N_38);
nor U6822 (N_6822,N_2106,N_1931);
nand U6823 (N_6823,N_4756,N_4845);
nor U6824 (N_6824,N_2961,N_1882);
or U6825 (N_6825,N_15,N_3149);
or U6826 (N_6826,N_4801,N_3491);
and U6827 (N_6827,N_634,N_1029);
nor U6828 (N_6828,N_320,N_1410);
and U6829 (N_6829,N_234,N_4809);
xor U6830 (N_6830,N_4103,N_1658);
nand U6831 (N_6831,N_1169,N_2486);
xnor U6832 (N_6832,N_4555,N_4449);
xnor U6833 (N_6833,N_1853,N_2438);
nand U6834 (N_6834,N_3810,N_3391);
nand U6835 (N_6835,N_70,N_4706);
xnor U6836 (N_6836,N_2636,N_4144);
and U6837 (N_6837,N_275,N_3979);
and U6838 (N_6838,N_3117,N_133);
and U6839 (N_6839,N_1699,N_2609);
and U6840 (N_6840,N_4636,N_2293);
and U6841 (N_6841,N_814,N_3769);
or U6842 (N_6842,N_2734,N_2635);
nor U6843 (N_6843,N_3539,N_4837);
and U6844 (N_6844,N_4074,N_2382);
and U6845 (N_6845,N_4761,N_4061);
or U6846 (N_6846,N_3999,N_2373);
nor U6847 (N_6847,N_1816,N_2255);
and U6848 (N_6848,N_782,N_3896);
or U6849 (N_6849,N_340,N_1976);
nand U6850 (N_6850,N_2112,N_1669);
and U6851 (N_6851,N_2476,N_3520);
or U6852 (N_6852,N_3780,N_2076);
and U6853 (N_6853,N_4713,N_2882);
xor U6854 (N_6854,N_687,N_1619);
xor U6855 (N_6855,N_1984,N_3711);
and U6856 (N_6856,N_3806,N_2998);
or U6857 (N_6857,N_305,N_1196);
and U6858 (N_6858,N_3895,N_130);
or U6859 (N_6859,N_4481,N_1426);
xor U6860 (N_6860,N_4371,N_2579);
or U6861 (N_6861,N_1966,N_4610);
or U6862 (N_6862,N_2042,N_3384);
nor U6863 (N_6863,N_1613,N_924);
xor U6864 (N_6864,N_767,N_1579);
nand U6865 (N_6865,N_298,N_2391);
or U6866 (N_6866,N_1325,N_1971);
and U6867 (N_6867,N_2562,N_4654);
nand U6868 (N_6868,N_1394,N_3028);
or U6869 (N_6869,N_4273,N_951);
or U6870 (N_6870,N_2431,N_3825);
or U6871 (N_6871,N_1644,N_1933);
nor U6872 (N_6872,N_1609,N_387);
and U6873 (N_6873,N_4268,N_3593);
or U6874 (N_6874,N_608,N_1261);
nor U6875 (N_6875,N_2778,N_1183);
and U6876 (N_6876,N_4394,N_1156);
or U6877 (N_6877,N_3793,N_947);
nor U6878 (N_6878,N_764,N_2887);
and U6879 (N_6879,N_3206,N_4233);
or U6880 (N_6880,N_1234,N_4307);
xnor U6881 (N_6881,N_4143,N_4829);
nand U6882 (N_6882,N_2721,N_3803);
nor U6883 (N_6883,N_2388,N_4499);
xnor U6884 (N_6884,N_412,N_747);
and U6885 (N_6885,N_1154,N_961);
xnor U6886 (N_6886,N_1192,N_3216);
nor U6887 (N_6887,N_3739,N_1471);
nor U6888 (N_6888,N_1625,N_1950);
or U6889 (N_6889,N_44,N_2664);
and U6890 (N_6890,N_937,N_346);
and U6891 (N_6891,N_894,N_4930);
nand U6892 (N_6892,N_4848,N_932);
and U6893 (N_6893,N_3955,N_4505);
and U6894 (N_6894,N_1042,N_1879);
and U6895 (N_6895,N_3575,N_2122);
and U6896 (N_6896,N_4118,N_4070);
and U6897 (N_6897,N_1502,N_2850);
xor U6898 (N_6898,N_1205,N_2203);
and U6899 (N_6899,N_2614,N_600);
xor U6900 (N_6900,N_1999,N_4029);
and U6901 (N_6901,N_473,N_1546);
or U6902 (N_6902,N_1079,N_4905);
nand U6903 (N_6903,N_2554,N_1068);
or U6904 (N_6904,N_3136,N_4875);
nor U6905 (N_6905,N_4131,N_4421);
or U6906 (N_6906,N_4213,N_3783);
nor U6907 (N_6907,N_4033,N_2411);
nand U6908 (N_6908,N_977,N_3008);
nand U6909 (N_6909,N_1486,N_2051);
or U6910 (N_6910,N_2057,N_545);
nor U6911 (N_6911,N_4263,N_3749);
xnor U6912 (N_6912,N_1520,N_2641);
or U6913 (N_6913,N_2172,N_1796);
xnor U6914 (N_6914,N_3235,N_4059);
nor U6915 (N_6915,N_3934,N_4574);
nor U6916 (N_6916,N_939,N_1597);
xnor U6917 (N_6917,N_1956,N_1065);
nor U6918 (N_6918,N_2628,N_4923);
or U6919 (N_6919,N_811,N_3903);
nor U6920 (N_6920,N_1693,N_2473);
or U6921 (N_6921,N_4770,N_2898);
xor U6922 (N_6922,N_1945,N_2802);
nor U6923 (N_6923,N_690,N_4765);
nor U6924 (N_6924,N_1581,N_4664);
nor U6925 (N_6925,N_1354,N_3471);
or U6926 (N_6926,N_1904,N_125);
and U6927 (N_6927,N_3627,N_1815);
or U6928 (N_6928,N_4920,N_3557);
nand U6929 (N_6929,N_1170,N_2575);
or U6930 (N_6930,N_376,N_2266);
or U6931 (N_6931,N_4482,N_128);
and U6932 (N_6932,N_997,N_978);
or U6933 (N_6933,N_4184,N_1476);
xnor U6934 (N_6934,N_756,N_3300);
nor U6935 (N_6935,N_1282,N_720);
and U6936 (N_6936,N_1295,N_3073);
nand U6937 (N_6937,N_1472,N_2788);
or U6938 (N_6938,N_4661,N_3511);
or U6939 (N_6939,N_1724,N_4410);
nand U6940 (N_6940,N_4957,N_313);
and U6941 (N_6941,N_4682,N_4136);
nor U6942 (N_6942,N_1983,N_1556);
or U6943 (N_6943,N_3676,N_4437);
and U6944 (N_6944,N_2540,N_4381);
and U6945 (N_6945,N_3102,N_4402);
or U6946 (N_6946,N_2481,N_3167);
nor U6947 (N_6947,N_3296,N_873);
and U6948 (N_6948,N_674,N_393);
nor U6949 (N_6949,N_294,N_1002);
nor U6950 (N_6950,N_2638,N_1327);
nor U6951 (N_6951,N_3543,N_1380);
and U6952 (N_6952,N_2002,N_1784);
nand U6953 (N_6953,N_1761,N_3664);
nor U6954 (N_6954,N_4925,N_4484);
nor U6955 (N_6955,N_1666,N_4357);
nor U6956 (N_6956,N_3613,N_2751);
xor U6957 (N_6957,N_2563,N_4901);
and U6958 (N_6958,N_4090,N_4432);
nor U6959 (N_6959,N_4746,N_1708);
and U6960 (N_6960,N_3358,N_1484);
nand U6961 (N_6961,N_2332,N_215);
xnor U6962 (N_6962,N_4339,N_1481);
and U6963 (N_6963,N_3549,N_2986);
nand U6964 (N_6964,N_4940,N_4662);
and U6965 (N_6965,N_4201,N_4903);
and U6966 (N_6966,N_4951,N_4551);
nor U6967 (N_6967,N_2743,N_1531);
xnor U6968 (N_6968,N_4841,N_3271);
xnor U6969 (N_6969,N_2513,N_2054);
nor U6970 (N_6970,N_1283,N_4459);
xor U6971 (N_6971,N_4566,N_1993);
nand U6972 (N_6972,N_3237,N_461);
and U6973 (N_6973,N_4696,N_4038);
or U6974 (N_6974,N_4587,N_287);
or U6975 (N_6975,N_3907,N_3983);
nand U6976 (N_6976,N_4110,N_423);
nand U6977 (N_6977,N_4549,N_653);
xor U6978 (N_6978,N_2809,N_4447);
nor U6979 (N_6979,N_3500,N_2445);
nand U6980 (N_6980,N_2543,N_1727);
and U6981 (N_6981,N_3475,N_2730);
nor U6982 (N_6982,N_2312,N_4238);
and U6983 (N_6983,N_127,N_859);
xnor U6984 (N_6984,N_2201,N_3259);
and U6985 (N_6985,N_2288,N_3643);
and U6986 (N_6986,N_2290,N_2921);
nand U6987 (N_6987,N_4385,N_2458);
and U6988 (N_6988,N_869,N_2228);
nor U6989 (N_6989,N_1269,N_4715);
nand U6990 (N_6990,N_352,N_2706);
nand U6991 (N_6991,N_2153,N_4466);
nand U6992 (N_6992,N_2124,N_2704);
and U6993 (N_6993,N_154,N_4322);
nand U6994 (N_6994,N_66,N_837);
nor U6995 (N_6995,N_4941,N_3236);
nand U6996 (N_6996,N_1273,N_4846);
nor U6997 (N_6997,N_1250,N_3620);
xnor U6998 (N_6998,N_82,N_1973);
nand U6999 (N_6999,N_269,N_3016);
nand U7000 (N_7000,N_2873,N_3153);
and U7001 (N_7001,N_2528,N_1677);
nand U7002 (N_7002,N_584,N_648);
xnor U7003 (N_7003,N_2901,N_554);
or U7004 (N_7004,N_2273,N_4839);
nand U7005 (N_7005,N_1215,N_4530);
nand U7006 (N_7006,N_4514,N_3189);
nor U7007 (N_7007,N_1558,N_1450);
xor U7008 (N_7008,N_4222,N_4011);
xor U7009 (N_7009,N_4171,N_1980);
nor U7010 (N_7010,N_4067,N_91);
or U7011 (N_7011,N_3376,N_4492);
nor U7012 (N_7012,N_1969,N_1804);
xor U7013 (N_7013,N_830,N_3325);
and U7014 (N_7014,N_686,N_789);
or U7015 (N_7015,N_3049,N_4256);
nand U7016 (N_7016,N_1104,N_4934);
and U7017 (N_7017,N_3482,N_4262);
or U7018 (N_7018,N_1628,N_543);
and U7019 (N_7019,N_1027,N_4393);
xor U7020 (N_7020,N_2281,N_1120);
xnor U7021 (N_7021,N_578,N_3663);
nor U7022 (N_7022,N_1833,N_3401);
nor U7023 (N_7023,N_2306,N_588);
nor U7024 (N_7024,N_2679,N_4978);
xor U7025 (N_7025,N_1779,N_1056);
xor U7026 (N_7026,N_949,N_775);
xor U7027 (N_7027,N_152,N_540);
nand U7028 (N_7028,N_1125,N_516);
or U7029 (N_7029,N_4666,N_89);
or U7030 (N_7030,N_4346,N_1254);
nand U7031 (N_7031,N_157,N_1830);
xor U7032 (N_7032,N_2553,N_1018);
or U7033 (N_7033,N_2855,N_1801);
xor U7034 (N_7034,N_985,N_4031);
nand U7035 (N_7035,N_1399,N_3700);
nand U7036 (N_7036,N_740,N_1143);
or U7037 (N_7037,N_1114,N_257);
or U7038 (N_7038,N_1185,N_2593);
xnor U7039 (N_7039,N_1854,N_3488);
or U7040 (N_7040,N_195,N_2688);
or U7041 (N_7041,N_4874,N_4735);
and U7042 (N_7042,N_2589,N_4856);
nor U7043 (N_7043,N_1725,N_4476);
nor U7044 (N_7044,N_2379,N_1526);
nor U7045 (N_7045,N_3247,N_2233);
nand U7046 (N_7046,N_3727,N_4827);
or U7047 (N_7047,N_3812,N_1701);
or U7048 (N_7048,N_4320,N_1992);
nor U7049 (N_7049,N_92,N_3320);
xnor U7050 (N_7050,N_1368,N_1802);
nor U7051 (N_7051,N_2410,N_4048);
nor U7052 (N_7052,N_2316,N_2488);
nor U7053 (N_7053,N_2508,N_2987);
nand U7054 (N_7054,N_3961,N_1605);
nor U7055 (N_7055,N_3751,N_417);
or U7056 (N_7056,N_2907,N_3813);
and U7057 (N_7057,N_1003,N_2319);
xor U7058 (N_7058,N_1781,N_1423);
nor U7059 (N_7059,N_34,N_1253);
and U7060 (N_7060,N_1022,N_3805);
xor U7061 (N_7061,N_4813,N_911);
nor U7062 (N_7062,N_4154,N_2469);
nor U7063 (N_7063,N_1362,N_51);
or U7064 (N_7064,N_246,N_895);
and U7065 (N_7065,N_786,N_3463);
or U7066 (N_7066,N_3174,N_668);
xnor U7067 (N_7067,N_2649,N_1067);
nand U7068 (N_7068,N_3656,N_1407);
and U7069 (N_7069,N_523,N_3112);
xor U7070 (N_7070,N_4093,N_4091);
nand U7071 (N_7071,N_2359,N_2181);
xnor U7072 (N_7072,N_4724,N_1568);
xnor U7073 (N_7073,N_281,N_1974);
xnor U7074 (N_7074,N_3657,N_4567);
nor U7075 (N_7075,N_1588,N_1849);
xnor U7076 (N_7076,N_2173,N_637);
nor U7077 (N_7077,N_4677,N_4576);
or U7078 (N_7078,N_2787,N_3680);
xnor U7079 (N_7079,N_3428,N_1926);
and U7080 (N_7080,N_1411,N_1176);
or U7081 (N_7081,N_3438,N_726);
and U7082 (N_7082,N_2243,N_2053);
and U7083 (N_7083,N_1718,N_4312);
xor U7084 (N_7084,N_1893,N_3782);
and U7085 (N_7085,N_1453,N_1241);
nor U7086 (N_7086,N_4240,N_4998);
and U7087 (N_7087,N_4888,N_3869);
xnor U7088 (N_7088,N_3303,N_4291);
xor U7089 (N_7089,N_1263,N_3654);
nor U7090 (N_7090,N_3943,N_2175);
nor U7091 (N_7091,N_816,N_838);
nor U7092 (N_7092,N_1288,N_2662);
and U7093 (N_7093,N_3930,N_3070);
nor U7094 (N_7094,N_4891,N_1171);
nor U7095 (N_7095,N_3675,N_2116);
nand U7096 (N_7096,N_1203,N_4992);
xor U7097 (N_7097,N_2663,N_4803);
nand U7098 (N_7098,N_1167,N_710);
xor U7099 (N_7099,N_2013,N_722);
xnor U7100 (N_7100,N_1265,N_1734);
xnor U7101 (N_7101,N_1460,N_4521);
nand U7102 (N_7102,N_4489,N_3305);
nand U7103 (N_7103,N_3850,N_2258);
or U7104 (N_7104,N_1527,N_2524);
nand U7105 (N_7105,N_4496,N_1924);
and U7106 (N_7106,N_860,N_910);
nand U7107 (N_7107,N_1560,N_3554);
xnor U7108 (N_7108,N_1315,N_2137);
nand U7109 (N_7109,N_3900,N_3686);
xnor U7110 (N_7110,N_4192,N_4024);
nor U7111 (N_7111,N_4415,N_4344);
and U7112 (N_7112,N_3473,N_4883);
and U7113 (N_7113,N_2141,N_1823);
xor U7114 (N_7114,N_2582,N_4135);
xor U7115 (N_7115,N_1831,N_336);
xnor U7116 (N_7116,N_1668,N_1015);
or U7117 (N_7117,N_2239,N_2936);
xnor U7118 (N_7118,N_2252,N_3107);
and U7119 (N_7119,N_1821,N_2159);
and U7120 (N_7120,N_4674,N_3602);
nand U7121 (N_7121,N_3103,N_4825);
xor U7122 (N_7122,N_3312,N_4822);
nor U7123 (N_7123,N_3370,N_2404);
xnor U7124 (N_7124,N_4493,N_2291);
and U7125 (N_7125,N_2585,N_3187);
and U7126 (N_7126,N_3253,N_217);
or U7127 (N_7127,N_3433,N_4026);
and U7128 (N_7128,N_3634,N_371);
nand U7129 (N_7129,N_1736,N_2868);
or U7130 (N_7130,N_2574,N_612);
nor U7131 (N_7131,N_3632,N_1091);
nand U7132 (N_7132,N_3477,N_468);
and U7133 (N_7133,N_3168,N_2994);
and U7134 (N_7134,N_2462,N_1467);
nor U7135 (N_7135,N_2467,N_4607);
nand U7136 (N_7136,N_4311,N_4178);
and U7137 (N_7137,N_1874,N_4251);
nor U7138 (N_7138,N_3503,N_2350);
nor U7139 (N_7139,N_455,N_2480);
xor U7140 (N_7140,N_1324,N_4028);
nor U7141 (N_7141,N_3734,N_780);
or U7142 (N_7142,N_4180,N_771);
nor U7143 (N_7143,N_467,N_1181);
nor U7144 (N_7144,N_4583,N_3434);
nand U7145 (N_7145,N_3412,N_1436);
and U7146 (N_7146,N_1226,N_1103);
and U7147 (N_7147,N_173,N_4003);
or U7148 (N_7148,N_2416,N_4252);
or U7149 (N_7149,N_4259,N_2590);
or U7150 (N_7150,N_4472,N_2964);
nor U7151 (N_7151,N_2309,N_1555);
nor U7152 (N_7152,N_4318,N_3291);
nand U7153 (N_7153,N_4958,N_3508);
or U7154 (N_7154,N_4591,N_3366);
or U7155 (N_7155,N_4170,N_2610);
xnor U7156 (N_7156,N_3197,N_4039);
nand U7157 (N_7157,N_986,N_3884);
nand U7158 (N_7158,N_3267,N_4302);
nor U7159 (N_7159,N_3268,N_2485);
or U7160 (N_7160,N_429,N_1667);
nand U7161 (N_7161,N_1346,N_2033);
or U7162 (N_7162,N_2892,N_2409);
or U7163 (N_7163,N_4095,N_129);
and U7164 (N_7164,N_1240,N_3797);
or U7165 (N_7165,N_2012,N_4108);
nor U7166 (N_7166,N_1990,N_1836);
nand U7167 (N_7167,N_2863,N_3977);
nor U7168 (N_7168,N_2440,N_519);
nand U7169 (N_7169,N_3671,N_2055);
nand U7170 (N_7170,N_2118,N_2195);
nor U7171 (N_7171,N_675,N_761);
or U7172 (N_7172,N_1987,N_2957);
and U7173 (N_7173,N_4900,N_1213);
and U7174 (N_7174,N_841,N_4929);
nand U7175 (N_7175,N_3324,N_1532);
nor U7176 (N_7176,N_3229,N_646);
nor U7177 (N_7177,N_494,N_1495);
or U7178 (N_7178,N_3441,N_2333);
and U7179 (N_7179,N_2906,N_1627);
xor U7180 (N_7180,N_4525,N_649);
xor U7181 (N_7181,N_85,N_3196);
and U7182 (N_7182,N_2676,N_422);
nand U7183 (N_7183,N_4467,N_3536);
nor U7184 (N_7184,N_696,N_942);
xor U7185 (N_7185,N_1221,N_474);
nand U7186 (N_7186,N_351,N_1388);
nor U7187 (N_7187,N_2912,N_4928);
xnor U7188 (N_7188,N_1768,N_3763);
and U7189 (N_7189,N_2687,N_344);
xnor U7190 (N_7190,N_2919,N_3386);
xor U7191 (N_7191,N_4044,N_559);
xor U7192 (N_7192,N_1517,N_264);
xnor U7193 (N_7193,N_3130,N_3914);
and U7194 (N_7194,N_1139,N_868);
or U7195 (N_7195,N_619,N_774);
xnor U7196 (N_7196,N_4258,N_4890);
xor U7197 (N_7197,N_3600,N_518);
and U7198 (N_7198,N_420,N_2531);
and U7199 (N_7199,N_2030,N_4495);
or U7200 (N_7200,N_1035,N_3846);
and U7201 (N_7201,N_526,N_3791);
nand U7202 (N_7202,N_4181,N_745);
nand U7203 (N_7203,N_2571,N_1344);
nand U7204 (N_7204,N_3730,N_295);
and U7205 (N_7205,N_452,N_4830);
nand U7206 (N_7206,N_1492,N_1072);
nor U7207 (N_7207,N_3899,N_4860);
nor U7208 (N_7208,N_1474,N_1828);
nor U7209 (N_7209,N_333,N_4423);
xor U7210 (N_7210,N_235,N_2123);
or U7211 (N_7211,N_3467,N_3321);
and U7212 (N_7212,N_2880,N_1519);
nor U7213 (N_7213,N_289,N_4236);
and U7214 (N_7214,N_4104,N_1247);
or U7215 (N_7215,N_2970,N_2605);
or U7216 (N_7216,N_4622,N_3041);
nor U7217 (N_7217,N_4652,N_1892);
and U7218 (N_7218,N_3935,N_1888);
xnor U7219 (N_7219,N_2815,N_1438);
nor U7220 (N_7220,N_4858,N_1948);
nand U7221 (N_7221,N_3368,N_13);
nor U7222 (N_7222,N_3009,N_3781);
xnor U7223 (N_7223,N_3158,N_836);
and U7224 (N_7224,N_2884,N_943);
nand U7225 (N_7225,N_1162,N_4162);
or U7226 (N_7226,N_4653,N_3258);
or U7227 (N_7227,N_3154,N_1772);
or U7228 (N_7228,N_2816,N_74);
and U7229 (N_7229,N_2542,N_1681);
xnor U7230 (N_7230,N_4261,N_4060);
and U7231 (N_7231,N_2807,N_6);
or U7232 (N_7232,N_3224,N_1428);
nor U7233 (N_7233,N_1069,N_4439);
nor U7234 (N_7234,N_3086,N_666);
xnor U7235 (N_7235,N_3854,N_98);
nor U7236 (N_7236,N_3298,N_3516);
or U7237 (N_7237,N_2718,N_4391);
or U7238 (N_7238,N_2668,N_3677);
and U7239 (N_7239,N_277,N_2225);
or U7240 (N_7240,N_4445,N_486);
nor U7241 (N_7241,N_103,N_3659);
and U7242 (N_7242,N_4734,N_4167);
and U7243 (N_7243,N_126,N_663);
nand U7244 (N_7244,N_2403,N_2468);
or U7245 (N_7245,N_2103,N_1751);
and U7246 (N_7246,N_1166,N_4237);
xor U7247 (N_7247,N_3156,N_3193);
or U7248 (N_7248,N_2226,N_3226);
or U7249 (N_7249,N_834,N_2286);
or U7250 (N_7250,N_2019,N_2031);
and U7251 (N_7251,N_4148,N_2171);
nand U7252 (N_7252,N_4221,N_4707);
xor U7253 (N_7253,N_2781,N_222);
xnor U7254 (N_7254,N_813,N_1813);
or U7255 (N_7255,N_135,N_3765);
and U7256 (N_7256,N_4089,N_4955);
or U7257 (N_7257,N_4742,N_2232);
and U7258 (N_7258,N_3726,N_2851);
nor U7259 (N_7259,N_1413,N_1757);
and U7260 (N_7260,N_2674,N_4563);
xnor U7261 (N_7261,N_2199,N_449);
or U7262 (N_7262,N_3356,N_4086);
or U7263 (N_7263,N_1516,N_164);
and U7264 (N_7264,N_680,N_1331);
nor U7265 (N_7265,N_238,N_4732);
and U7266 (N_7266,N_3596,N_2728);
or U7267 (N_7267,N_1787,N_3030);
and U7268 (N_7268,N_1511,N_4218);
and U7269 (N_7269,N_4224,N_569);
or U7270 (N_7270,N_2242,N_2047);
nor U7271 (N_7271,N_2622,N_631);
nor U7272 (N_7272,N_2363,N_1580);
and U7273 (N_7273,N_3927,N_1680);
nor U7274 (N_7274,N_1552,N_2014);
nand U7275 (N_7275,N_1119,N_4363);
or U7276 (N_7276,N_2451,N_4140);
nand U7277 (N_7277,N_1794,N_4174);
nor U7278 (N_7278,N_4248,N_3355);
or U7279 (N_7279,N_3776,N_4959);
xor U7280 (N_7280,N_1246,N_2866);
xor U7281 (N_7281,N_485,N_2653);
nor U7282 (N_7282,N_2008,N_1314);
or U7283 (N_7283,N_3629,N_4578);
nor U7284 (N_7284,N_177,N_1786);
or U7285 (N_7285,N_2678,N_2011);
or U7286 (N_7286,N_3081,N_4420);
and U7287 (N_7287,N_1633,N_4994);
xor U7288 (N_7288,N_4547,N_4049);
nor U7289 (N_7289,N_52,N_174);
or U7290 (N_7290,N_101,N_574);
xnor U7291 (N_7291,N_254,N_1151);
nor U7292 (N_7292,N_850,N_4102);
and U7293 (N_7293,N_159,N_2673);
or U7294 (N_7294,N_4112,N_1752);
and U7295 (N_7295,N_1739,N_1791);
nor U7296 (N_7296,N_3461,N_71);
nor U7297 (N_7297,N_1262,N_4899);
and U7298 (N_7298,N_759,N_2615);
nand U7299 (N_7299,N_3588,N_1142);
nor U7300 (N_7300,N_124,N_1090);
and U7301 (N_7301,N_84,N_97);
and U7302 (N_7302,N_2374,N_1443);
and U7303 (N_7303,N_512,N_1006);
xnor U7304 (N_7304,N_1447,N_749);
nor U7305 (N_7305,N_1043,N_4352);
and U7306 (N_7306,N_2545,N_2594);
nor U7307 (N_7307,N_3849,N_575);
or U7308 (N_7308,N_3489,N_306);
and U7309 (N_7309,N_1818,N_1808);
xnor U7310 (N_7310,N_2733,N_1137);
and U7311 (N_7311,N_2113,N_1073);
nor U7312 (N_7312,N_1050,N_2231);
xor U7313 (N_7313,N_2487,N_2156);
and U7314 (N_7314,N_750,N_1051);
and U7315 (N_7315,N_374,N_2949);
xnor U7316 (N_7316,N_2981,N_1178);
nand U7317 (N_7317,N_2808,N_538);
and U7318 (N_7318,N_2321,N_1319);
xnor U7319 (N_7319,N_4695,N_2130);
xnor U7320 (N_7320,N_2997,N_441);
nand U7321 (N_7321,N_12,N_4478);
nand U7322 (N_7322,N_3450,N_3127);
xor U7323 (N_7323,N_2120,N_462);
nand U7324 (N_7324,N_1601,N_2114);
or U7325 (N_7325,N_854,N_3001);
nand U7326 (N_7326,N_918,N_226);
xor U7327 (N_7327,N_3651,N_3523);
or U7328 (N_7328,N_2812,N_3945);
and U7329 (N_7329,N_2274,N_4183);
nand U7330 (N_7330,N_2736,N_501);
nor U7331 (N_7331,N_4231,N_2187);
or U7332 (N_7332,N_2527,N_1845);
or U7333 (N_7333,N_3217,N_1994);
nor U7334 (N_7334,N_4541,N_2443);
and U7335 (N_7335,N_1538,N_2954);
xnor U7336 (N_7336,N_1606,N_1908);
nand U7337 (N_7337,N_274,N_4805);
xnor U7338 (N_7338,N_3761,N_4347);
or U7339 (N_7339,N_2237,N_2081);
nor U7340 (N_7340,N_4789,N_3619);
nand U7341 (N_7341,N_3709,N_1509);
nand U7342 (N_7342,N_606,N_2827);
xnor U7343 (N_7343,N_4522,N_3280);
and U7344 (N_7344,N_877,N_4226);
xnor U7345 (N_7345,N_1991,N_2234);
nand U7346 (N_7346,N_4811,N_4985);
or U7347 (N_7347,N_2608,N_4392);
nor U7348 (N_7348,N_282,N_4988);
nand U7349 (N_7349,N_3591,N_1256);
nor U7350 (N_7350,N_3264,N_2749);
or U7351 (N_7351,N_4133,N_2482);
or U7352 (N_7352,N_1264,N_75);
xor U7353 (N_7353,N_2504,N_63);
nor U7354 (N_7354,N_2754,N_988);
or U7355 (N_7355,N_348,N_3856);
nand U7356 (N_7356,N_3585,N_827);
or U7357 (N_7357,N_3842,N_4373);
nand U7358 (N_7358,N_4294,N_3672);
and U7359 (N_7359,N_4161,N_5);
nand U7360 (N_7360,N_1938,N_3148);
nor U7361 (N_7361,N_3892,N_3342);
nand U7362 (N_7362,N_2899,N_1333);
nor U7363 (N_7363,N_2142,N_3082);
nand U7364 (N_7364,N_2779,N_4769);
or U7365 (N_7365,N_3323,N_3104);
xor U7366 (N_7366,N_1124,N_4413);
nand U7367 (N_7367,N_4050,N_3279);
xnor U7368 (N_7368,N_3121,N_2612);
or U7369 (N_7369,N_3612,N_3169);
nand U7370 (N_7370,N_3839,N_4386);
and U7371 (N_7371,N_936,N_3043);
and U7372 (N_7372,N_4189,N_1639);
xor U7373 (N_7373,N_1740,N_4426);
nand U7374 (N_7374,N_2675,N_613);
nand U7375 (N_7375,N_664,N_672);
and U7376 (N_7376,N_421,N_3225);
nand U7377 (N_7377,N_2261,N_636);
xor U7378 (N_7378,N_3984,N_4993);
and U7379 (N_7379,N_1951,N_1776);
nand U7380 (N_7380,N_1457,N_3625);
and U7381 (N_7381,N_1713,N_1491);
and U7382 (N_7382,N_2710,N_3034);
and U7383 (N_7383,N_4295,N_337);
nor U7384 (N_7384,N_2211,N_3584);
and U7385 (N_7385,N_3951,N_229);
xnor U7386 (N_7386,N_4673,N_4023);
xnor U7387 (N_7387,N_1377,N_1366);
and U7388 (N_7388,N_513,N_4084);
or U7389 (N_7389,N_2217,N_917);
and U7390 (N_7390,N_1939,N_4532);
nand U7391 (N_7391,N_4979,N_3343);
nor U7392 (N_7392,N_4448,N_476);
or U7393 (N_7393,N_3599,N_1235);
or U7394 (N_7394,N_1769,N_3800);
xor U7395 (N_7395,N_77,N_4589);
xnor U7396 (N_7396,N_1953,N_4323);
and U7397 (N_7397,N_1946,N_471);
xnor U7398 (N_7398,N_2279,N_4355);
xor U7399 (N_7399,N_527,N_4798);
nand U7400 (N_7400,N_2158,N_283);
xnor U7401 (N_7401,N_611,N_2774);
and U7402 (N_7402,N_2117,N_4892);
nor U7403 (N_7403,N_2651,N_4862);
nand U7404 (N_7404,N_2690,N_4861);
xnor U7405 (N_7405,N_3708,N_465);
and U7406 (N_7406,N_4282,N_4279);
nor U7407 (N_7407,N_4404,N_1553);
and U7408 (N_7408,N_4971,N_842);
nand U7409 (N_7409,N_2793,N_1358);
nor U7410 (N_7410,N_3492,N_2960);
or U7411 (N_7411,N_3004,N_4987);
xor U7412 (N_7412,N_4097,N_1576);
nand U7413 (N_7413,N_2040,N_252);
xor U7414 (N_7414,N_104,N_3715);
xnor U7415 (N_7415,N_1611,N_1136);
or U7416 (N_7416,N_3630,N_493);
xnor U7417 (N_7417,N_54,N_392);
nor U7418 (N_7418,N_1759,N_1415);
nand U7419 (N_7419,N_2161,N_3852);
nand U7420 (N_7420,N_3024,N_1963);
or U7421 (N_7421,N_3015,N_4624);
and U7422 (N_7422,N_891,N_380);
xor U7423 (N_7423,N_4793,N_3075);
nand U7424 (N_7424,N_2965,N_1037);
or U7425 (N_7425,N_2210,N_2719);
xor U7426 (N_7426,N_3580,N_622);
nor U7427 (N_7427,N_3108,N_2072);
nand U7428 (N_7428,N_484,N_1313);
and U7429 (N_7429,N_659,N_1645);
or U7430 (N_7430,N_1883,N_3705);
nor U7431 (N_7431,N_729,N_2249);
nand U7432 (N_7432,N_1021,N_1656);
nand U7433 (N_7433,N_3870,N_361);
or U7434 (N_7434,N_567,N_4287);
or U7435 (N_7435,N_4921,N_4708);
nand U7436 (N_7436,N_3195,N_3735);
nand U7437 (N_7437,N_3990,N_1390);
xnor U7438 (N_7438,N_4527,N_1123);
nand U7439 (N_7439,N_4370,N_1723);
xor U7440 (N_7440,N_2523,N_3964);
or U7441 (N_7441,N_1268,N_3962);
nand U7442 (N_7442,N_4646,N_3923);
xor U7443 (N_7443,N_770,N_498);
xor U7444 (N_7444,N_1887,N_2165);
xnor U7445 (N_7445,N_4612,N_109);
xnor U7446 (N_7446,N_1884,N_3860);
or U7447 (N_7447,N_4598,N_4904);
nor U7448 (N_7448,N_3558,N_255);
or U7449 (N_7449,N_4571,N_1733);
nand U7450 (N_7450,N_969,N_2846);
xnor U7451 (N_7451,N_733,N_1299);
and U7452 (N_7452,N_1165,N_1870);
nand U7453 (N_7453,N_185,N_4585);
and U7454 (N_7454,N_604,N_3844);
or U7455 (N_7455,N_576,N_2125);
xor U7456 (N_7456,N_2900,N_223);
and U7457 (N_7457,N_1435,N_958);
nand U7458 (N_7458,N_2100,N_882);
xor U7459 (N_7459,N_2762,N_3365);
and U7460 (N_7460,N_406,N_3774);
or U7461 (N_7461,N_3036,N_3078);
and U7462 (N_7462,N_4187,N_4126);
or U7463 (N_7463,N_2157,N_2601);
nand U7464 (N_7464,N_795,N_2294);
xor U7465 (N_7465,N_823,N_3222);
or U7466 (N_7466,N_3796,N_3431);
nor U7467 (N_7467,N_2417,N_1168);
nor U7468 (N_7468,N_4293,N_1847);
nand U7469 (N_7469,N_1391,N_4429);
or U7470 (N_7470,N_4877,N_22);
nor U7471 (N_7471,N_715,N_3642);
nand U7472 (N_7472,N_2352,N_4215);
xor U7473 (N_7473,N_2152,N_3881);
nor U7474 (N_7474,N_1753,N_3470);
nand U7475 (N_7475,N_1045,N_1524);
xnor U7476 (N_7476,N_3592,N_3790);
and U7477 (N_7477,N_90,N_2671);
or U7478 (N_7478,N_706,N_3650);
nor U7479 (N_7479,N_4642,N_4669);
nand U7480 (N_7480,N_2768,N_2069);
and U7481 (N_7481,N_4274,N_1920);
nand U7482 (N_7482,N_4406,N_4280);
or U7483 (N_7483,N_3330,N_702);
nand U7484 (N_7484,N_4207,N_511);
nand U7485 (N_7485,N_2824,N_872);
or U7486 (N_7486,N_4808,N_2700);
or U7487 (N_7487,N_288,N_2348);
nor U7488 (N_7488,N_1917,N_4924);
nor U7489 (N_7489,N_314,N_290);
nand U7490 (N_7490,N_2514,N_4560);
and U7491 (N_7491,N_699,N_4999);
xor U7492 (N_7492,N_2889,N_1356);
or U7493 (N_7493,N_1803,N_996);
nor U7494 (N_7494,N_2376,N_2715);
and U7495 (N_7495,N_3002,N_3925);
and U7496 (N_7496,N_394,N_1838);
and U7497 (N_7497,N_4509,N_3309);
nand U7498 (N_7498,N_927,N_2093);
or U7499 (N_7499,N_1843,N_1303);
or U7500 (N_7500,N_1662,N_2262);
xor U7501 (N_7501,N_2811,N_1189);
xnor U7502 (N_7502,N_4407,N_4856);
nand U7503 (N_7503,N_2897,N_835);
and U7504 (N_7504,N_701,N_3022);
xnor U7505 (N_7505,N_3742,N_4353);
nand U7506 (N_7506,N_1316,N_367);
and U7507 (N_7507,N_4054,N_2679);
nor U7508 (N_7508,N_3211,N_2697);
nor U7509 (N_7509,N_735,N_737);
xnor U7510 (N_7510,N_2322,N_1283);
or U7511 (N_7511,N_1471,N_3824);
xnor U7512 (N_7512,N_396,N_3860);
and U7513 (N_7513,N_348,N_1941);
or U7514 (N_7514,N_1804,N_3590);
or U7515 (N_7515,N_1273,N_3534);
nor U7516 (N_7516,N_2623,N_4288);
xnor U7517 (N_7517,N_1303,N_2877);
and U7518 (N_7518,N_166,N_4202);
or U7519 (N_7519,N_4648,N_1012);
and U7520 (N_7520,N_3548,N_2294);
xnor U7521 (N_7521,N_607,N_4558);
nand U7522 (N_7522,N_3979,N_2434);
nor U7523 (N_7523,N_710,N_427);
or U7524 (N_7524,N_39,N_1287);
xnor U7525 (N_7525,N_3526,N_3555);
nor U7526 (N_7526,N_3334,N_2913);
or U7527 (N_7527,N_4895,N_1274);
or U7528 (N_7528,N_4660,N_1327);
xor U7529 (N_7529,N_665,N_2345);
nand U7530 (N_7530,N_2160,N_1275);
or U7531 (N_7531,N_3875,N_3568);
xor U7532 (N_7532,N_671,N_2109);
xnor U7533 (N_7533,N_3425,N_2288);
and U7534 (N_7534,N_4780,N_1202);
xor U7535 (N_7535,N_958,N_3552);
and U7536 (N_7536,N_4380,N_704);
nor U7537 (N_7537,N_4103,N_1968);
xnor U7538 (N_7538,N_331,N_3184);
xnor U7539 (N_7539,N_130,N_2164);
xor U7540 (N_7540,N_52,N_3314);
nor U7541 (N_7541,N_2044,N_2369);
nor U7542 (N_7542,N_3279,N_4853);
nor U7543 (N_7543,N_3758,N_1874);
or U7544 (N_7544,N_817,N_4526);
nor U7545 (N_7545,N_4728,N_910);
nand U7546 (N_7546,N_3517,N_1906);
nor U7547 (N_7547,N_2495,N_2236);
or U7548 (N_7548,N_904,N_970);
nor U7549 (N_7549,N_2894,N_1498);
and U7550 (N_7550,N_4010,N_3428);
nand U7551 (N_7551,N_3598,N_1734);
xnor U7552 (N_7552,N_2380,N_2211);
nand U7553 (N_7553,N_2082,N_1952);
xor U7554 (N_7554,N_3806,N_4288);
xnor U7555 (N_7555,N_249,N_238);
or U7556 (N_7556,N_823,N_2699);
and U7557 (N_7557,N_1821,N_2765);
nand U7558 (N_7558,N_4792,N_3737);
nand U7559 (N_7559,N_1531,N_2720);
nand U7560 (N_7560,N_2170,N_4544);
nor U7561 (N_7561,N_4742,N_1280);
nand U7562 (N_7562,N_2282,N_2205);
or U7563 (N_7563,N_3104,N_407);
nand U7564 (N_7564,N_1782,N_1923);
nor U7565 (N_7565,N_4639,N_4859);
xnor U7566 (N_7566,N_617,N_3240);
nor U7567 (N_7567,N_4549,N_3299);
xnor U7568 (N_7568,N_515,N_2965);
nand U7569 (N_7569,N_2803,N_3731);
or U7570 (N_7570,N_448,N_1895);
and U7571 (N_7571,N_2108,N_1085);
nor U7572 (N_7572,N_4318,N_3864);
nor U7573 (N_7573,N_1848,N_3236);
and U7574 (N_7574,N_1164,N_2143);
nor U7575 (N_7575,N_2997,N_3354);
and U7576 (N_7576,N_4442,N_4887);
xor U7577 (N_7577,N_4598,N_1229);
nor U7578 (N_7578,N_2807,N_2622);
xor U7579 (N_7579,N_824,N_1728);
nor U7580 (N_7580,N_3907,N_2161);
and U7581 (N_7581,N_1234,N_152);
xor U7582 (N_7582,N_2747,N_2389);
or U7583 (N_7583,N_3729,N_1774);
xnor U7584 (N_7584,N_3931,N_3133);
or U7585 (N_7585,N_4657,N_581);
xnor U7586 (N_7586,N_508,N_3107);
nand U7587 (N_7587,N_3869,N_3626);
or U7588 (N_7588,N_853,N_2372);
nand U7589 (N_7589,N_3500,N_2693);
or U7590 (N_7590,N_1985,N_4445);
nor U7591 (N_7591,N_2011,N_3735);
nand U7592 (N_7592,N_4112,N_2062);
xnor U7593 (N_7593,N_2277,N_1414);
nor U7594 (N_7594,N_2435,N_3960);
or U7595 (N_7595,N_2006,N_1316);
nor U7596 (N_7596,N_631,N_2764);
nor U7597 (N_7597,N_4726,N_1043);
nor U7598 (N_7598,N_4459,N_2308);
nand U7599 (N_7599,N_1001,N_3050);
nand U7600 (N_7600,N_2250,N_2369);
or U7601 (N_7601,N_3813,N_152);
nand U7602 (N_7602,N_3406,N_2068);
nor U7603 (N_7603,N_966,N_2970);
xor U7604 (N_7604,N_3916,N_682);
nand U7605 (N_7605,N_732,N_4181);
and U7606 (N_7606,N_972,N_4225);
nand U7607 (N_7607,N_4886,N_1406);
nand U7608 (N_7608,N_3814,N_2611);
nand U7609 (N_7609,N_4554,N_3756);
nand U7610 (N_7610,N_2639,N_588);
nor U7611 (N_7611,N_464,N_4518);
nand U7612 (N_7612,N_140,N_2640);
and U7613 (N_7613,N_3105,N_258);
and U7614 (N_7614,N_4832,N_1003);
xnor U7615 (N_7615,N_4943,N_2063);
and U7616 (N_7616,N_734,N_1271);
or U7617 (N_7617,N_2034,N_368);
and U7618 (N_7618,N_2386,N_3353);
and U7619 (N_7619,N_2034,N_3849);
or U7620 (N_7620,N_1899,N_4711);
nand U7621 (N_7621,N_3780,N_1529);
and U7622 (N_7622,N_2753,N_880);
xnor U7623 (N_7623,N_1495,N_1546);
nor U7624 (N_7624,N_113,N_1216);
nand U7625 (N_7625,N_4795,N_3196);
nor U7626 (N_7626,N_1427,N_2915);
nand U7627 (N_7627,N_3997,N_4877);
nand U7628 (N_7628,N_3958,N_3331);
xor U7629 (N_7629,N_4211,N_591);
nand U7630 (N_7630,N_3047,N_1611);
nor U7631 (N_7631,N_1194,N_2510);
and U7632 (N_7632,N_1695,N_2417);
nor U7633 (N_7633,N_1091,N_478);
xnor U7634 (N_7634,N_1291,N_1469);
xor U7635 (N_7635,N_1879,N_3078);
nand U7636 (N_7636,N_2652,N_4031);
nor U7637 (N_7637,N_4550,N_70);
xor U7638 (N_7638,N_2003,N_1777);
and U7639 (N_7639,N_644,N_2373);
nor U7640 (N_7640,N_2918,N_4655);
xnor U7641 (N_7641,N_125,N_3675);
nand U7642 (N_7642,N_4388,N_1097);
nand U7643 (N_7643,N_4007,N_4412);
nor U7644 (N_7644,N_122,N_4126);
or U7645 (N_7645,N_2142,N_618);
xor U7646 (N_7646,N_3137,N_3002);
or U7647 (N_7647,N_2814,N_2090);
xor U7648 (N_7648,N_603,N_4045);
xor U7649 (N_7649,N_3354,N_2789);
nor U7650 (N_7650,N_4136,N_1191);
and U7651 (N_7651,N_3770,N_2218);
or U7652 (N_7652,N_2954,N_3229);
or U7653 (N_7653,N_761,N_566);
nor U7654 (N_7654,N_3299,N_4731);
and U7655 (N_7655,N_2057,N_1111);
nand U7656 (N_7656,N_1787,N_4417);
xnor U7657 (N_7657,N_2346,N_4614);
nor U7658 (N_7658,N_2759,N_1884);
or U7659 (N_7659,N_4155,N_4688);
nor U7660 (N_7660,N_613,N_305);
nor U7661 (N_7661,N_168,N_2361);
xnor U7662 (N_7662,N_2726,N_4742);
or U7663 (N_7663,N_4301,N_108);
and U7664 (N_7664,N_2076,N_2879);
and U7665 (N_7665,N_2675,N_466);
and U7666 (N_7666,N_1801,N_4594);
or U7667 (N_7667,N_4382,N_1057);
xnor U7668 (N_7668,N_3870,N_2649);
nand U7669 (N_7669,N_2245,N_4656);
xor U7670 (N_7670,N_4175,N_2664);
nor U7671 (N_7671,N_1360,N_767);
and U7672 (N_7672,N_4812,N_3619);
or U7673 (N_7673,N_4325,N_4996);
xor U7674 (N_7674,N_2750,N_3745);
nor U7675 (N_7675,N_1155,N_375);
xnor U7676 (N_7676,N_108,N_1478);
nand U7677 (N_7677,N_2155,N_972);
nor U7678 (N_7678,N_2516,N_1389);
and U7679 (N_7679,N_1712,N_1665);
nand U7680 (N_7680,N_4674,N_3156);
or U7681 (N_7681,N_3449,N_4715);
xnor U7682 (N_7682,N_2324,N_855);
nand U7683 (N_7683,N_2962,N_3236);
and U7684 (N_7684,N_4795,N_3661);
nor U7685 (N_7685,N_4713,N_32);
or U7686 (N_7686,N_2359,N_4962);
nand U7687 (N_7687,N_3880,N_3230);
nand U7688 (N_7688,N_2599,N_878);
nor U7689 (N_7689,N_50,N_2147);
and U7690 (N_7690,N_4183,N_1984);
nor U7691 (N_7691,N_2416,N_1506);
or U7692 (N_7692,N_615,N_2953);
and U7693 (N_7693,N_4153,N_2105);
or U7694 (N_7694,N_1696,N_701);
xor U7695 (N_7695,N_2323,N_1372);
and U7696 (N_7696,N_2248,N_507);
nor U7697 (N_7697,N_4178,N_1552);
nand U7698 (N_7698,N_3918,N_528);
nand U7699 (N_7699,N_462,N_4839);
and U7700 (N_7700,N_2637,N_4772);
nor U7701 (N_7701,N_2040,N_2608);
nor U7702 (N_7702,N_4947,N_4015);
and U7703 (N_7703,N_3550,N_432);
nand U7704 (N_7704,N_2426,N_4155);
xnor U7705 (N_7705,N_1947,N_2563);
nor U7706 (N_7706,N_3847,N_4935);
nand U7707 (N_7707,N_852,N_4604);
nor U7708 (N_7708,N_2682,N_2153);
or U7709 (N_7709,N_1705,N_1883);
nand U7710 (N_7710,N_2691,N_410);
nand U7711 (N_7711,N_4234,N_4270);
or U7712 (N_7712,N_9,N_1292);
or U7713 (N_7713,N_4166,N_338);
or U7714 (N_7714,N_2827,N_3067);
nor U7715 (N_7715,N_538,N_2401);
nor U7716 (N_7716,N_4815,N_4882);
xor U7717 (N_7717,N_4406,N_4107);
and U7718 (N_7718,N_4081,N_2653);
nand U7719 (N_7719,N_3661,N_3197);
and U7720 (N_7720,N_2613,N_3050);
and U7721 (N_7721,N_1902,N_4813);
or U7722 (N_7722,N_2206,N_1208);
and U7723 (N_7723,N_3630,N_2522);
nand U7724 (N_7724,N_3006,N_1995);
and U7725 (N_7725,N_3367,N_1411);
xor U7726 (N_7726,N_1583,N_314);
xor U7727 (N_7727,N_2665,N_400);
xnor U7728 (N_7728,N_3574,N_4113);
xor U7729 (N_7729,N_1718,N_823);
xor U7730 (N_7730,N_1166,N_4335);
nand U7731 (N_7731,N_1844,N_1581);
nor U7732 (N_7732,N_2432,N_2683);
or U7733 (N_7733,N_2557,N_151);
or U7734 (N_7734,N_3504,N_641);
and U7735 (N_7735,N_2317,N_2925);
nor U7736 (N_7736,N_2923,N_4281);
nor U7737 (N_7737,N_1411,N_2624);
nand U7738 (N_7738,N_1320,N_1226);
nor U7739 (N_7739,N_4637,N_2869);
nand U7740 (N_7740,N_3143,N_3424);
and U7741 (N_7741,N_2084,N_290);
xnor U7742 (N_7742,N_3757,N_3579);
and U7743 (N_7743,N_3969,N_1949);
nand U7744 (N_7744,N_1172,N_2449);
nand U7745 (N_7745,N_3866,N_3571);
nor U7746 (N_7746,N_2048,N_2980);
and U7747 (N_7747,N_2520,N_622);
and U7748 (N_7748,N_2810,N_3789);
nor U7749 (N_7749,N_3128,N_3777);
nor U7750 (N_7750,N_952,N_2107);
nand U7751 (N_7751,N_1686,N_4575);
nor U7752 (N_7752,N_4389,N_2801);
xnor U7753 (N_7753,N_1058,N_1660);
nor U7754 (N_7754,N_4855,N_2857);
nor U7755 (N_7755,N_3246,N_1081);
or U7756 (N_7756,N_2102,N_51);
and U7757 (N_7757,N_3908,N_1124);
or U7758 (N_7758,N_1287,N_909);
nand U7759 (N_7759,N_706,N_1998);
and U7760 (N_7760,N_1317,N_1776);
and U7761 (N_7761,N_4847,N_4644);
xnor U7762 (N_7762,N_4500,N_2624);
xor U7763 (N_7763,N_969,N_54);
or U7764 (N_7764,N_2134,N_110);
or U7765 (N_7765,N_3303,N_946);
xor U7766 (N_7766,N_3473,N_1596);
nand U7767 (N_7767,N_1112,N_1792);
and U7768 (N_7768,N_3597,N_4261);
nand U7769 (N_7769,N_3944,N_1241);
nand U7770 (N_7770,N_3268,N_247);
or U7771 (N_7771,N_384,N_2288);
nor U7772 (N_7772,N_2675,N_615);
nand U7773 (N_7773,N_3949,N_1183);
nand U7774 (N_7774,N_1663,N_4169);
xnor U7775 (N_7775,N_1803,N_1145);
or U7776 (N_7776,N_2474,N_1000);
and U7777 (N_7777,N_2662,N_648);
or U7778 (N_7778,N_1012,N_2996);
xor U7779 (N_7779,N_4014,N_2047);
or U7780 (N_7780,N_4671,N_3979);
nor U7781 (N_7781,N_2168,N_447);
nand U7782 (N_7782,N_750,N_3405);
or U7783 (N_7783,N_1830,N_549);
or U7784 (N_7784,N_3109,N_4699);
nor U7785 (N_7785,N_3343,N_1027);
or U7786 (N_7786,N_3,N_1288);
nand U7787 (N_7787,N_781,N_4778);
nor U7788 (N_7788,N_4041,N_1864);
and U7789 (N_7789,N_2183,N_4707);
xnor U7790 (N_7790,N_3164,N_583);
or U7791 (N_7791,N_3101,N_2334);
or U7792 (N_7792,N_4710,N_924);
xnor U7793 (N_7793,N_569,N_4813);
nor U7794 (N_7794,N_2883,N_1167);
nor U7795 (N_7795,N_2931,N_4552);
xnor U7796 (N_7796,N_114,N_711);
nand U7797 (N_7797,N_2120,N_1546);
or U7798 (N_7798,N_3325,N_2448);
xnor U7799 (N_7799,N_727,N_2051);
or U7800 (N_7800,N_3434,N_3220);
nor U7801 (N_7801,N_2857,N_3308);
nor U7802 (N_7802,N_4401,N_65);
or U7803 (N_7803,N_105,N_3807);
or U7804 (N_7804,N_3937,N_1529);
nor U7805 (N_7805,N_2460,N_4385);
xor U7806 (N_7806,N_4601,N_3906);
nand U7807 (N_7807,N_1835,N_4486);
xor U7808 (N_7808,N_1556,N_4623);
and U7809 (N_7809,N_1516,N_2638);
nand U7810 (N_7810,N_1577,N_1898);
and U7811 (N_7811,N_1356,N_4813);
or U7812 (N_7812,N_1130,N_3166);
xor U7813 (N_7813,N_2233,N_4815);
xnor U7814 (N_7814,N_4150,N_3068);
and U7815 (N_7815,N_2887,N_4731);
or U7816 (N_7816,N_1452,N_4260);
nor U7817 (N_7817,N_4575,N_2893);
nand U7818 (N_7818,N_583,N_649);
or U7819 (N_7819,N_1469,N_2498);
nor U7820 (N_7820,N_4728,N_4296);
nor U7821 (N_7821,N_4426,N_4226);
xnor U7822 (N_7822,N_3565,N_3573);
xor U7823 (N_7823,N_1680,N_149);
or U7824 (N_7824,N_4889,N_11);
nor U7825 (N_7825,N_2837,N_850);
nand U7826 (N_7826,N_2024,N_67);
xnor U7827 (N_7827,N_2315,N_3);
nor U7828 (N_7828,N_3766,N_4901);
nor U7829 (N_7829,N_1786,N_4569);
nand U7830 (N_7830,N_2338,N_332);
or U7831 (N_7831,N_3415,N_2903);
or U7832 (N_7832,N_4804,N_969);
or U7833 (N_7833,N_2660,N_1127);
or U7834 (N_7834,N_2901,N_1290);
nand U7835 (N_7835,N_3441,N_1770);
nor U7836 (N_7836,N_3007,N_3050);
nand U7837 (N_7837,N_1652,N_3907);
nand U7838 (N_7838,N_816,N_2214);
or U7839 (N_7839,N_2725,N_2585);
or U7840 (N_7840,N_2287,N_358);
and U7841 (N_7841,N_2030,N_2371);
nand U7842 (N_7842,N_4186,N_1716);
xnor U7843 (N_7843,N_42,N_4229);
nor U7844 (N_7844,N_2001,N_2572);
and U7845 (N_7845,N_2930,N_2636);
and U7846 (N_7846,N_4265,N_4673);
or U7847 (N_7847,N_1403,N_1970);
nand U7848 (N_7848,N_4984,N_265);
xnor U7849 (N_7849,N_2754,N_1571);
xnor U7850 (N_7850,N_3665,N_3438);
nor U7851 (N_7851,N_3037,N_4509);
or U7852 (N_7852,N_3777,N_4334);
or U7853 (N_7853,N_11,N_2420);
xor U7854 (N_7854,N_2068,N_3150);
and U7855 (N_7855,N_2389,N_1633);
nand U7856 (N_7856,N_4066,N_4895);
nand U7857 (N_7857,N_1690,N_2925);
nor U7858 (N_7858,N_2265,N_139);
nor U7859 (N_7859,N_2495,N_1252);
nor U7860 (N_7860,N_4899,N_3384);
nor U7861 (N_7861,N_3032,N_3788);
nand U7862 (N_7862,N_988,N_493);
xnor U7863 (N_7863,N_1372,N_2611);
nor U7864 (N_7864,N_4739,N_4874);
xor U7865 (N_7865,N_2619,N_4942);
xnor U7866 (N_7866,N_988,N_3901);
xor U7867 (N_7867,N_4824,N_1088);
or U7868 (N_7868,N_1181,N_472);
nor U7869 (N_7869,N_4908,N_2374);
xor U7870 (N_7870,N_3866,N_3998);
or U7871 (N_7871,N_211,N_4430);
nor U7872 (N_7872,N_2051,N_4142);
and U7873 (N_7873,N_298,N_907);
nor U7874 (N_7874,N_806,N_3990);
or U7875 (N_7875,N_4954,N_4237);
nand U7876 (N_7876,N_795,N_4958);
and U7877 (N_7877,N_328,N_2275);
nor U7878 (N_7878,N_921,N_3075);
and U7879 (N_7879,N_4604,N_4001);
and U7880 (N_7880,N_1289,N_1481);
xor U7881 (N_7881,N_4226,N_4826);
nand U7882 (N_7882,N_874,N_4429);
nand U7883 (N_7883,N_4318,N_3328);
and U7884 (N_7884,N_2652,N_758);
nor U7885 (N_7885,N_3962,N_4807);
xor U7886 (N_7886,N_861,N_1081);
and U7887 (N_7887,N_4280,N_1748);
nor U7888 (N_7888,N_3407,N_3880);
nor U7889 (N_7889,N_4742,N_1888);
nor U7890 (N_7890,N_3166,N_1647);
and U7891 (N_7891,N_3965,N_1678);
or U7892 (N_7892,N_2842,N_74);
and U7893 (N_7893,N_3867,N_3771);
or U7894 (N_7894,N_2550,N_3407);
xor U7895 (N_7895,N_1370,N_3693);
and U7896 (N_7896,N_3911,N_3010);
and U7897 (N_7897,N_736,N_829);
and U7898 (N_7898,N_4278,N_2075);
nor U7899 (N_7899,N_2044,N_3005);
nand U7900 (N_7900,N_1149,N_58);
or U7901 (N_7901,N_2833,N_4681);
or U7902 (N_7902,N_1615,N_769);
or U7903 (N_7903,N_2863,N_4995);
or U7904 (N_7904,N_1980,N_2542);
nand U7905 (N_7905,N_2517,N_3516);
nand U7906 (N_7906,N_3015,N_1395);
nor U7907 (N_7907,N_1261,N_3517);
and U7908 (N_7908,N_138,N_3724);
and U7909 (N_7909,N_3261,N_3755);
nor U7910 (N_7910,N_2798,N_1222);
xnor U7911 (N_7911,N_121,N_1690);
nand U7912 (N_7912,N_827,N_27);
nor U7913 (N_7913,N_150,N_4449);
or U7914 (N_7914,N_578,N_1491);
and U7915 (N_7915,N_2381,N_4718);
or U7916 (N_7916,N_442,N_1022);
or U7917 (N_7917,N_4162,N_3761);
or U7918 (N_7918,N_1143,N_4988);
xnor U7919 (N_7919,N_1781,N_3112);
xnor U7920 (N_7920,N_2900,N_1836);
nor U7921 (N_7921,N_4964,N_800);
or U7922 (N_7922,N_3693,N_1453);
or U7923 (N_7923,N_3779,N_2547);
or U7924 (N_7924,N_2109,N_1100);
xnor U7925 (N_7925,N_1371,N_4705);
or U7926 (N_7926,N_1388,N_1290);
nor U7927 (N_7927,N_4883,N_489);
xnor U7928 (N_7928,N_4567,N_160);
nand U7929 (N_7929,N_1329,N_343);
nand U7930 (N_7930,N_4446,N_2584);
nand U7931 (N_7931,N_4756,N_539);
nor U7932 (N_7932,N_49,N_773);
xnor U7933 (N_7933,N_4000,N_4836);
nand U7934 (N_7934,N_2526,N_2069);
xnor U7935 (N_7935,N_3585,N_282);
nand U7936 (N_7936,N_4619,N_3623);
xor U7937 (N_7937,N_4294,N_558);
and U7938 (N_7938,N_954,N_4303);
nor U7939 (N_7939,N_195,N_2367);
xnor U7940 (N_7940,N_3545,N_3580);
xnor U7941 (N_7941,N_4205,N_2870);
xor U7942 (N_7942,N_2743,N_4331);
or U7943 (N_7943,N_4173,N_4106);
or U7944 (N_7944,N_2673,N_658);
and U7945 (N_7945,N_1124,N_260);
xor U7946 (N_7946,N_2358,N_297);
or U7947 (N_7947,N_2079,N_548);
nor U7948 (N_7948,N_4437,N_2118);
xor U7949 (N_7949,N_4912,N_4139);
nor U7950 (N_7950,N_2820,N_1590);
or U7951 (N_7951,N_2798,N_4545);
nor U7952 (N_7952,N_3999,N_2564);
and U7953 (N_7953,N_4475,N_319);
or U7954 (N_7954,N_4109,N_2983);
or U7955 (N_7955,N_3671,N_2642);
or U7956 (N_7956,N_1785,N_48);
xnor U7957 (N_7957,N_2853,N_3530);
nand U7958 (N_7958,N_3709,N_1331);
nor U7959 (N_7959,N_3900,N_1496);
or U7960 (N_7960,N_46,N_4066);
nand U7961 (N_7961,N_2754,N_4847);
nor U7962 (N_7962,N_617,N_329);
or U7963 (N_7963,N_211,N_1438);
xor U7964 (N_7964,N_1192,N_1701);
nor U7965 (N_7965,N_1922,N_3527);
xor U7966 (N_7966,N_725,N_4382);
nor U7967 (N_7967,N_1130,N_3401);
xnor U7968 (N_7968,N_3227,N_759);
xnor U7969 (N_7969,N_1029,N_3965);
nor U7970 (N_7970,N_624,N_3937);
nand U7971 (N_7971,N_2092,N_3902);
or U7972 (N_7972,N_251,N_1930);
xor U7973 (N_7973,N_1213,N_4966);
or U7974 (N_7974,N_4024,N_2696);
nand U7975 (N_7975,N_82,N_3385);
and U7976 (N_7976,N_1986,N_1803);
nor U7977 (N_7977,N_4379,N_960);
and U7978 (N_7978,N_4251,N_2830);
and U7979 (N_7979,N_1207,N_1290);
and U7980 (N_7980,N_588,N_4363);
nor U7981 (N_7981,N_814,N_22);
xnor U7982 (N_7982,N_596,N_3112);
nor U7983 (N_7983,N_899,N_723);
or U7984 (N_7984,N_4656,N_4143);
xor U7985 (N_7985,N_1580,N_4655);
nand U7986 (N_7986,N_1,N_440);
nand U7987 (N_7987,N_4672,N_4363);
nand U7988 (N_7988,N_2188,N_3162);
nand U7989 (N_7989,N_4004,N_4250);
xor U7990 (N_7990,N_3727,N_4376);
xor U7991 (N_7991,N_4541,N_2372);
and U7992 (N_7992,N_2754,N_2170);
or U7993 (N_7993,N_3713,N_123);
or U7994 (N_7994,N_904,N_934);
nor U7995 (N_7995,N_2766,N_1219);
nor U7996 (N_7996,N_4405,N_4273);
or U7997 (N_7997,N_4152,N_1963);
nand U7998 (N_7998,N_2147,N_4241);
nand U7999 (N_7999,N_895,N_1394);
or U8000 (N_8000,N_1389,N_1017);
xor U8001 (N_8001,N_1643,N_4240);
nand U8002 (N_8002,N_1311,N_512);
nand U8003 (N_8003,N_197,N_4310);
or U8004 (N_8004,N_1342,N_4545);
nor U8005 (N_8005,N_3498,N_4421);
xnor U8006 (N_8006,N_136,N_1589);
nand U8007 (N_8007,N_1853,N_3052);
and U8008 (N_8008,N_2665,N_3184);
xor U8009 (N_8009,N_726,N_1719);
nand U8010 (N_8010,N_1773,N_1893);
and U8011 (N_8011,N_4900,N_3311);
xnor U8012 (N_8012,N_2840,N_921);
nor U8013 (N_8013,N_2222,N_2525);
and U8014 (N_8014,N_969,N_4518);
or U8015 (N_8015,N_2994,N_1619);
or U8016 (N_8016,N_1508,N_597);
and U8017 (N_8017,N_4065,N_1178);
xor U8018 (N_8018,N_394,N_451);
or U8019 (N_8019,N_4518,N_654);
or U8020 (N_8020,N_1111,N_3352);
nand U8021 (N_8021,N_1934,N_3866);
or U8022 (N_8022,N_2573,N_4636);
nor U8023 (N_8023,N_814,N_2749);
and U8024 (N_8024,N_1561,N_2531);
and U8025 (N_8025,N_929,N_4223);
nor U8026 (N_8026,N_1232,N_4196);
nor U8027 (N_8027,N_2950,N_197);
or U8028 (N_8028,N_2324,N_2327);
or U8029 (N_8029,N_1104,N_1779);
and U8030 (N_8030,N_1422,N_2736);
xor U8031 (N_8031,N_1720,N_4774);
xor U8032 (N_8032,N_3888,N_3556);
xnor U8033 (N_8033,N_523,N_2450);
xor U8034 (N_8034,N_305,N_3060);
or U8035 (N_8035,N_2298,N_124);
xnor U8036 (N_8036,N_3710,N_4278);
nor U8037 (N_8037,N_4748,N_3122);
nor U8038 (N_8038,N_4490,N_4902);
xnor U8039 (N_8039,N_4380,N_3450);
nor U8040 (N_8040,N_959,N_2870);
or U8041 (N_8041,N_3538,N_4846);
nor U8042 (N_8042,N_1585,N_2152);
nand U8043 (N_8043,N_2473,N_3378);
nand U8044 (N_8044,N_4680,N_3946);
nand U8045 (N_8045,N_4061,N_2299);
xnor U8046 (N_8046,N_470,N_307);
nor U8047 (N_8047,N_3032,N_835);
or U8048 (N_8048,N_3388,N_2865);
xor U8049 (N_8049,N_4802,N_1990);
nor U8050 (N_8050,N_3479,N_4894);
and U8051 (N_8051,N_192,N_2332);
xnor U8052 (N_8052,N_1989,N_4883);
xor U8053 (N_8053,N_34,N_4015);
and U8054 (N_8054,N_1032,N_3222);
nand U8055 (N_8055,N_3438,N_1770);
xnor U8056 (N_8056,N_3816,N_4375);
and U8057 (N_8057,N_4970,N_4232);
and U8058 (N_8058,N_3706,N_4965);
or U8059 (N_8059,N_1648,N_2806);
and U8060 (N_8060,N_2807,N_2784);
xor U8061 (N_8061,N_722,N_2607);
xor U8062 (N_8062,N_2485,N_1131);
and U8063 (N_8063,N_4741,N_3731);
nor U8064 (N_8064,N_878,N_744);
and U8065 (N_8065,N_2170,N_2224);
xor U8066 (N_8066,N_4895,N_1317);
nor U8067 (N_8067,N_1650,N_3931);
or U8068 (N_8068,N_353,N_61);
nor U8069 (N_8069,N_1628,N_520);
xnor U8070 (N_8070,N_1769,N_1733);
xnor U8071 (N_8071,N_1848,N_3406);
xnor U8072 (N_8072,N_1234,N_2737);
nand U8073 (N_8073,N_4847,N_1607);
nor U8074 (N_8074,N_1594,N_3974);
nor U8075 (N_8075,N_2510,N_3720);
nand U8076 (N_8076,N_3776,N_838);
nand U8077 (N_8077,N_754,N_4570);
nor U8078 (N_8078,N_1571,N_4303);
xnor U8079 (N_8079,N_2814,N_4673);
or U8080 (N_8080,N_3700,N_4880);
nor U8081 (N_8081,N_4104,N_4480);
and U8082 (N_8082,N_2888,N_4417);
nor U8083 (N_8083,N_3954,N_1222);
nand U8084 (N_8084,N_1712,N_3404);
or U8085 (N_8085,N_1877,N_3558);
nor U8086 (N_8086,N_3845,N_1018);
nor U8087 (N_8087,N_2642,N_2592);
and U8088 (N_8088,N_3064,N_1295);
nand U8089 (N_8089,N_2562,N_1867);
nor U8090 (N_8090,N_2736,N_2405);
and U8091 (N_8091,N_4789,N_2321);
nand U8092 (N_8092,N_2595,N_2052);
and U8093 (N_8093,N_4250,N_1626);
or U8094 (N_8094,N_2891,N_4144);
nor U8095 (N_8095,N_1217,N_4103);
nand U8096 (N_8096,N_1766,N_905);
nand U8097 (N_8097,N_3900,N_1135);
nor U8098 (N_8098,N_777,N_4632);
xor U8099 (N_8099,N_2881,N_3244);
nand U8100 (N_8100,N_2872,N_3369);
nand U8101 (N_8101,N_4653,N_1891);
xor U8102 (N_8102,N_3027,N_4642);
nor U8103 (N_8103,N_4930,N_750);
nand U8104 (N_8104,N_2268,N_2562);
nand U8105 (N_8105,N_1953,N_3929);
nor U8106 (N_8106,N_587,N_2780);
or U8107 (N_8107,N_2172,N_2413);
xor U8108 (N_8108,N_2391,N_785);
nor U8109 (N_8109,N_4781,N_4339);
and U8110 (N_8110,N_3627,N_2017);
nor U8111 (N_8111,N_2456,N_3398);
and U8112 (N_8112,N_4242,N_1568);
and U8113 (N_8113,N_1686,N_2527);
xor U8114 (N_8114,N_1411,N_2637);
nor U8115 (N_8115,N_3380,N_531);
and U8116 (N_8116,N_1142,N_591);
xnor U8117 (N_8117,N_1432,N_3491);
or U8118 (N_8118,N_1452,N_2932);
xor U8119 (N_8119,N_1221,N_4537);
and U8120 (N_8120,N_814,N_2624);
and U8121 (N_8121,N_1551,N_2979);
nor U8122 (N_8122,N_2534,N_878);
or U8123 (N_8123,N_3995,N_3744);
nor U8124 (N_8124,N_735,N_3169);
or U8125 (N_8125,N_2777,N_2150);
and U8126 (N_8126,N_2286,N_2129);
and U8127 (N_8127,N_1095,N_3968);
nor U8128 (N_8128,N_2991,N_2957);
or U8129 (N_8129,N_1277,N_4473);
nor U8130 (N_8130,N_1727,N_1926);
nor U8131 (N_8131,N_3132,N_2212);
or U8132 (N_8132,N_2080,N_47);
nor U8133 (N_8133,N_2210,N_1884);
nor U8134 (N_8134,N_3397,N_629);
or U8135 (N_8135,N_4389,N_3375);
nor U8136 (N_8136,N_3386,N_1478);
or U8137 (N_8137,N_1336,N_4539);
or U8138 (N_8138,N_2396,N_2960);
nor U8139 (N_8139,N_128,N_996);
xor U8140 (N_8140,N_2387,N_2620);
or U8141 (N_8141,N_1323,N_1032);
nand U8142 (N_8142,N_1567,N_555);
nand U8143 (N_8143,N_4034,N_4463);
nor U8144 (N_8144,N_2168,N_250);
nor U8145 (N_8145,N_3427,N_2415);
nand U8146 (N_8146,N_3278,N_3191);
xor U8147 (N_8147,N_42,N_4649);
or U8148 (N_8148,N_417,N_2952);
and U8149 (N_8149,N_2310,N_4396);
or U8150 (N_8150,N_3436,N_1444);
xor U8151 (N_8151,N_4671,N_893);
nor U8152 (N_8152,N_2185,N_1514);
and U8153 (N_8153,N_3948,N_4005);
xor U8154 (N_8154,N_2095,N_4451);
nor U8155 (N_8155,N_4393,N_2048);
and U8156 (N_8156,N_4477,N_2963);
nand U8157 (N_8157,N_3004,N_1912);
or U8158 (N_8158,N_1276,N_2067);
and U8159 (N_8159,N_194,N_4043);
nor U8160 (N_8160,N_2537,N_2223);
nand U8161 (N_8161,N_1844,N_1972);
nand U8162 (N_8162,N_4407,N_983);
nor U8163 (N_8163,N_1133,N_3242);
or U8164 (N_8164,N_2320,N_4417);
nand U8165 (N_8165,N_1290,N_1939);
and U8166 (N_8166,N_910,N_249);
and U8167 (N_8167,N_4780,N_3335);
or U8168 (N_8168,N_416,N_3973);
and U8169 (N_8169,N_433,N_2376);
or U8170 (N_8170,N_2957,N_3551);
nor U8171 (N_8171,N_3279,N_925);
nand U8172 (N_8172,N_2245,N_3191);
nand U8173 (N_8173,N_3075,N_853);
xnor U8174 (N_8174,N_3000,N_827);
xnor U8175 (N_8175,N_3447,N_545);
and U8176 (N_8176,N_4576,N_2409);
nor U8177 (N_8177,N_3579,N_227);
and U8178 (N_8178,N_3851,N_4737);
xnor U8179 (N_8179,N_4343,N_4834);
nand U8180 (N_8180,N_4779,N_2508);
xor U8181 (N_8181,N_127,N_1172);
nor U8182 (N_8182,N_2143,N_1568);
nand U8183 (N_8183,N_3167,N_1262);
nor U8184 (N_8184,N_4092,N_2698);
xor U8185 (N_8185,N_4163,N_867);
and U8186 (N_8186,N_4465,N_1810);
xor U8187 (N_8187,N_3011,N_3318);
nor U8188 (N_8188,N_3675,N_1065);
or U8189 (N_8189,N_4981,N_1830);
and U8190 (N_8190,N_3035,N_4028);
nand U8191 (N_8191,N_372,N_3911);
nor U8192 (N_8192,N_984,N_4959);
or U8193 (N_8193,N_3867,N_3495);
nand U8194 (N_8194,N_3334,N_4734);
nor U8195 (N_8195,N_2206,N_656);
xor U8196 (N_8196,N_1562,N_492);
nand U8197 (N_8197,N_544,N_4416);
or U8198 (N_8198,N_4741,N_1734);
nand U8199 (N_8199,N_2406,N_1379);
or U8200 (N_8200,N_526,N_1419);
and U8201 (N_8201,N_1596,N_1561);
nand U8202 (N_8202,N_2298,N_4064);
or U8203 (N_8203,N_4189,N_3477);
xor U8204 (N_8204,N_1251,N_360);
nand U8205 (N_8205,N_3546,N_2673);
xnor U8206 (N_8206,N_1164,N_4341);
nand U8207 (N_8207,N_3689,N_2325);
nand U8208 (N_8208,N_2413,N_591);
and U8209 (N_8209,N_624,N_1133);
nand U8210 (N_8210,N_3970,N_2492);
and U8211 (N_8211,N_4432,N_2577);
or U8212 (N_8212,N_1391,N_437);
nor U8213 (N_8213,N_328,N_3326);
and U8214 (N_8214,N_802,N_3455);
nor U8215 (N_8215,N_4240,N_3461);
xnor U8216 (N_8216,N_3621,N_1655);
nand U8217 (N_8217,N_4899,N_1251);
nor U8218 (N_8218,N_2892,N_1974);
nor U8219 (N_8219,N_3768,N_1175);
nand U8220 (N_8220,N_1952,N_1406);
nor U8221 (N_8221,N_2155,N_1899);
or U8222 (N_8222,N_4658,N_3823);
and U8223 (N_8223,N_2937,N_2541);
or U8224 (N_8224,N_4928,N_4183);
nand U8225 (N_8225,N_2601,N_3039);
nor U8226 (N_8226,N_2661,N_91);
nor U8227 (N_8227,N_2686,N_1618);
nand U8228 (N_8228,N_405,N_464);
nor U8229 (N_8229,N_3685,N_2470);
or U8230 (N_8230,N_1856,N_2033);
or U8231 (N_8231,N_3973,N_3413);
xnor U8232 (N_8232,N_3238,N_315);
or U8233 (N_8233,N_1821,N_4210);
nor U8234 (N_8234,N_1490,N_4869);
xor U8235 (N_8235,N_1275,N_1702);
nor U8236 (N_8236,N_159,N_3959);
and U8237 (N_8237,N_3343,N_47);
or U8238 (N_8238,N_4094,N_323);
nand U8239 (N_8239,N_1563,N_3191);
and U8240 (N_8240,N_1303,N_3169);
and U8241 (N_8241,N_1744,N_3432);
xor U8242 (N_8242,N_864,N_3139);
xor U8243 (N_8243,N_3971,N_1802);
and U8244 (N_8244,N_231,N_3943);
and U8245 (N_8245,N_1698,N_4632);
or U8246 (N_8246,N_3730,N_4130);
xor U8247 (N_8247,N_3537,N_1935);
xor U8248 (N_8248,N_2667,N_866);
or U8249 (N_8249,N_4189,N_470);
or U8250 (N_8250,N_2711,N_4084);
nand U8251 (N_8251,N_4492,N_2283);
or U8252 (N_8252,N_3937,N_4355);
and U8253 (N_8253,N_4480,N_3058);
nand U8254 (N_8254,N_1308,N_517);
and U8255 (N_8255,N_2218,N_4065);
nor U8256 (N_8256,N_3411,N_1748);
and U8257 (N_8257,N_1422,N_4428);
and U8258 (N_8258,N_3024,N_634);
and U8259 (N_8259,N_146,N_1934);
nor U8260 (N_8260,N_525,N_1986);
and U8261 (N_8261,N_3756,N_1079);
or U8262 (N_8262,N_534,N_1379);
nand U8263 (N_8263,N_2176,N_4439);
or U8264 (N_8264,N_798,N_4722);
nor U8265 (N_8265,N_2509,N_1153);
nand U8266 (N_8266,N_225,N_1722);
or U8267 (N_8267,N_3617,N_4064);
and U8268 (N_8268,N_3807,N_864);
nand U8269 (N_8269,N_4077,N_4161);
nor U8270 (N_8270,N_4406,N_3136);
and U8271 (N_8271,N_2547,N_2882);
or U8272 (N_8272,N_878,N_4306);
or U8273 (N_8273,N_3467,N_1699);
nand U8274 (N_8274,N_1058,N_3178);
xor U8275 (N_8275,N_1485,N_3745);
xor U8276 (N_8276,N_2324,N_1733);
xnor U8277 (N_8277,N_4851,N_666);
xnor U8278 (N_8278,N_777,N_2157);
xnor U8279 (N_8279,N_2867,N_1794);
nand U8280 (N_8280,N_2166,N_3263);
and U8281 (N_8281,N_3495,N_1789);
nand U8282 (N_8282,N_2695,N_1298);
xor U8283 (N_8283,N_4719,N_642);
xor U8284 (N_8284,N_1076,N_1984);
nor U8285 (N_8285,N_985,N_2931);
nor U8286 (N_8286,N_466,N_4611);
xnor U8287 (N_8287,N_4251,N_381);
xnor U8288 (N_8288,N_1151,N_1108);
nor U8289 (N_8289,N_4683,N_3774);
or U8290 (N_8290,N_1677,N_3176);
xor U8291 (N_8291,N_438,N_3998);
nor U8292 (N_8292,N_4198,N_32);
xor U8293 (N_8293,N_3617,N_21);
xnor U8294 (N_8294,N_607,N_3929);
xor U8295 (N_8295,N_1154,N_198);
or U8296 (N_8296,N_2179,N_2957);
or U8297 (N_8297,N_2177,N_807);
nor U8298 (N_8298,N_3792,N_4048);
nand U8299 (N_8299,N_4561,N_97);
xnor U8300 (N_8300,N_1188,N_908);
nand U8301 (N_8301,N_2720,N_2901);
nand U8302 (N_8302,N_4959,N_2571);
nand U8303 (N_8303,N_2749,N_1964);
nor U8304 (N_8304,N_1191,N_1331);
nor U8305 (N_8305,N_4123,N_1167);
nand U8306 (N_8306,N_4252,N_2632);
nand U8307 (N_8307,N_919,N_3396);
nand U8308 (N_8308,N_2564,N_4736);
nand U8309 (N_8309,N_1161,N_4609);
or U8310 (N_8310,N_1474,N_71);
nand U8311 (N_8311,N_1201,N_1941);
nand U8312 (N_8312,N_1253,N_1092);
nor U8313 (N_8313,N_2458,N_2519);
and U8314 (N_8314,N_1792,N_3198);
xor U8315 (N_8315,N_740,N_588);
or U8316 (N_8316,N_344,N_668);
nand U8317 (N_8317,N_1509,N_908);
nor U8318 (N_8318,N_2474,N_622);
xor U8319 (N_8319,N_1929,N_4578);
or U8320 (N_8320,N_2951,N_4686);
and U8321 (N_8321,N_2302,N_807);
and U8322 (N_8322,N_1734,N_1080);
nor U8323 (N_8323,N_4647,N_1438);
or U8324 (N_8324,N_458,N_3755);
or U8325 (N_8325,N_3335,N_4535);
nor U8326 (N_8326,N_1863,N_4348);
xnor U8327 (N_8327,N_1894,N_1301);
nor U8328 (N_8328,N_2043,N_3114);
nor U8329 (N_8329,N_2901,N_3851);
and U8330 (N_8330,N_3756,N_1959);
or U8331 (N_8331,N_1320,N_1590);
nand U8332 (N_8332,N_3111,N_2958);
xor U8333 (N_8333,N_2940,N_798);
nand U8334 (N_8334,N_987,N_184);
nor U8335 (N_8335,N_4098,N_4506);
and U8336 (N_8336,N_4106,N_951);
and U8337 (N_8337,N_1324,N_953);
and U8338 (N_8338,N_179,N_4195);
and U8339 (N_8339,N_709,N_4406);
or U8340 (N_8340,N_3039,N_3637);
and U8341 (N_8341,N_4856,N_2805);
and U8342 (N_8342,N_1399,N_1889);
or U8343 (N_8343,N_3992,N_4950);
xnor U8344 (N_8344,N_1405,N_1976);
nand U8345 (N_8345,N_1357,N_1827);
and U8346 (N_8346,N_3364,N_4455);
and U8347 (N_8347,N_4590,N_4252);
nor U8348 (N_8348,N_4165,N_4386);
nor U8349 (N_8349,N_2894,N_1813);
xor U8350 (N_8350,N_2248,N_4841);
nand U8351 (N_8351,N_4703,N_3723);
nor U8352 (N_8352,N_4118,N_4503);
xnor U8353 (N_8353,N_131,N_2534);
and U8354 (N_8354,N_3556,N_1785);
or U8355 (N_8355,N_3120,N_73);
xnor U8356 (N_8356,N_314,N_3996);
xnor U8357 (N_8357,N_3467,N_1254);
nor U8358 (N_8358,N_1341,N_1344);
nand U8359 (N_8359,N_2411,N_1791);
xor U8360 (N_8360,N_4643,N_4178);
nor U8361 (N_8361,N_790,N_507);
nand U8362 (N_8362,N_3548,N_636);
nor U8363 (N_8363,N_2451,N_3492);
or U8364 (N_8364,N_296,N_4792);
nand U8365 (N_8365,N_347,N_1364);
and U8366 (N_8366,N_3353,N_2565);
nand U8367 (N_8367,N_609,N_120);
nor U8368 (N_8368,N_4726,N_2524);
nor U8369 (N_8369,N_4092,N_1720);
nor U8370 (N_8370,N_1862,N_3408);
or U8371 (N_8371,N_1290,N_3099);
xnor U8372 (N_8372,N_2506,N_2062);
or U8373 (N_8373,N_4015,N_2413);
xnor U8374 (N_8374,N_2716,N_4769);
nand U8375 (N_8375,N_3576,N_4501);
and U8376 (N_8376,N_1480,N_500);
xnor U8377 (N_8377,N_4437,N_3663);
and U8378 (N_8378,N_2381,N_2442);
and U8379 (N_8379,N_776,N_2034);
or U8380 (N_8380,N_2586,N_2977);
nor U8381 (N_8381,N_1588,N_1198);
and U8382 (N_8382,N_1204,N_1257);
and U8383 (N_8383,N_57,N_3671);
xor U8384 (N_8384,N_2823,N_4567);
and U8385 (N_8385,N_1669,N_4633);
nand U8386 (N_8386,N_3642,N_4138);
nand U8387 (N_8387,N_1526,N_1175);
nand U8388 (N_8388,N_1855,N_2022);
xnor U8389 (N_8389,N_2022,N_854);
nor U8390 (N_8390,N_2631,N_2508);
nand U8391 (N_8391,N_2345,N_3234);
nand U8392 (N_8392,N_2013,N_2656);
or U8393 (N_8393,N_1796,N_2106);
nand U8394 (N_8394,N_1639,N_983);
and U8395 (N_8395,N_4092,N_270);
nand U8396 (N_8396,N_3045,N_4891);
nand U8397 (N_8397,N_1588,N_1983);
nor U8398 (N_8398,N_1735,N_4069);
xor U8399 (N_8399,N_4703,N_4533);
and U8400 (N_8400,N_2186,N_3706);
or U8401 (N_8401,N_142,N_3607);
xnor U8402 (N_8402,N_495,N_4682);
nor U8403 (N_8403,N_579,N_1658);
xor U8404 (N_8404,N_4550,N_2535);
nand U8405 (N_8405,N_635,N_3366);
nor U8406 (N_8406,N_3651,N_2218);
xnor U8407 (N_8407,N_3512,N_1877);
nand U8408 (N_8408,N_3029,N_2305);
and U8409 (N_8409,N_1872,N_2405);
and U8410 (N_8410,N_3483,N_1217);
nand U8411 (N_8411,N_41,N_2586);
xnor U8412 (N_8412,N_1739,N_132);
nand U8413 (N_8413,N_3376,N_750);
or U8414 (N_8414,N_1332,N_3775);
and U8415 (N_8415,N_993,N_3083);
or U8416 (N_8416,N_3550,N_4262);
nand U8417 (N_8417,N_840,N_556);
nand U8418 (N_8418,N_3518,N_1237);
nand U8419 (N_8419,N_2101,N_2749);
and U8420 (N_8420,N_409,N_283);
nor U8421 (N_8421,N_2872,N_2441);
and U8422 (N_8422,N_1479,N_2828);
nor U8423 (N_8423,N_3875,N_3477);
nand U8424 (N_8424,N_4502,N_2099);
nor U8425 (N_8425,N_2627,N_2787);
and U8426 (N_8426,N_1237,N_714);
and U8427 (N_8427,N_2181,N_2959);
xor U8428 (N_8428,N_2152,N_4412);
nand U8429 (N_8429,N_3244,N_1830);
and U8430 (N_8430,N_4470,N_76);
and U8431 (N_8431,N_236,N_2829);
or U8432 (N_8432,N_3712,N_15);
or U8433 (N_8433,N_2291,N_4460);
nand U8434 (N_8434,N_803,N_1550);
xnor U8435 (N_8435,N_2403,N_581);
or U8436 (N_8436,N_3524,N_1660);
or U8437 (N_8437,N_118,N_4225);
nor U8438 (N_8438,N_4733,N_2150);
and U8439 (N_8439,N_4450,N_1017);
nand U8440 (N_8440,N_1093,N_1466);
nor U8441 (N_8441,N_823,N_2559);
or U8442 (N_8442,N_3552,N_1014);
or U8443 (N_8443,N_122,N_1312);
xor U8444 (N_8444,N_3305,N_2469);
and U8445 (N_8445,N_1177,N_1460);
and U8446 (N_8446,N_398,N_3083);
and U8447 (N_8447,N_1987,N_4135);
or U8448 (N_8448,N_3336,N_1708);
and U8449 (N_8449,N_233,N_2828);
xor U8450 (N_8450,N_3606,N_63);
nor U8451 (N_8451,N_1756,N_4170);
or U8452 (N_8452,N_4228,N_4657);
and U8453 (N_8453,N_2796,N_646);
nor U8454 (N_8454,N_3186,N_4919);
xnor U8455 (N_8455,N_1449,N_4186);
nor U8456 (N_8456,N_2089,N_4490);
or U8457 (N_8457,N_4754,N_4488);
or U8458 (N_8458,N_3421,N_37);
nand U8459 (N_8459,N_579,N_2026);
and U8460 (N_8460,N_865,N_4637);
nand U8461 (N_8461,N_289,N_1403);
and U8462 (N_8462,N_3650,N_901);
or U8463 (N_8463,N_3131,N_4625);
nand U8464 (N_8464,N_1157,N_3647);
xnor U8465 (N_8465,N_3136,N_2940);
xnor U8466 (N_8466,N_2665,N_1740);
or U8467 (N_8467,N_2271,N_4330);
or U8468 (N_8468,N_1976,N_4546);
xor U8469 (N_8469,N_2982,N_1637);
nor U8470 (N_8470,N_378,N_4364);
nand U8471 (N_8471,N_4858,N_3798);
or U8472 (N_8472,N_2765,N_388);
nand U8473 (N_8473,N_1772,N_4545);
xnor U8474 (N_8474,N_4712,N_4127);
xnor U8475 (N_8475,N_453,N_201);
and U8476 (N_8476,N_1636,N_4425);
nand U8477 (N_8477,N_2886,N_594);
nand U8478 (N_8478,N_695,N_1240);
nand U8479 (N_8479,N_105,N_240);
and U8480 (N_8480,N_857,N_3144);
nand U8481 (N_8481,N_4093,N_4985);
nand U8482 (N_8482,N_2461,N_1519);
or U8483 (N_8483,N_1996,N_4488);
xnor U8484 (N_8484,N_3013,N_2699);
nand U8485 (N_8485,N_3129,N_1790);
and U8486 (N_8486,N_1802,N_4762);
and U8487 (N_8487,N_2660,N_126);
nor U8488 (N_8488,N_4265,N_829);
and U8489 (N_8489,N_3067,N_4890);
xor U8490 (N_8490,N_2881,N_3825);
or U8491 (N_8491,N_3089,N_3905);
and U8492 (N_8492,N_171,N_4258);
xor U8493 (N_8493,N_1302,N_1754);
xnor U8494 (N_8494,N_2937,N_4680);
nor U8495 (N_8495,N_2949,N_3030);
and U8496 (N_8496,N_4242,N_4375);
nor U8497 (N_8497,N_1279,N_640);
nand U8498 (N_8498,N_2231,N_4592);
and U8499 (N_8499,N_1863,N_2242);
xor U8500 (N_8500,N_171,N_2423);
and U8501 (N_8501,N_3883,N_3351);
or U8502 (N_8502,N_2083,N_4724);
nand U8503 (N_8503,N_4333,N_2083);
nand U8504 (N_8504,N_1857,N_2217);
xor U8505 (N_8505,N_1710,N_739);
or U8506 (N_8506,N_4606,N_1286);
xor U8507 (N_8507,N_3861,N_1369);
nor U8508 (N_8508,N_3664,N_4918);
nand U8509 (N_8509,N_1771,N_2374);
or U8510 (N_8510,N_943,N_388);
or U8511 (N_8511,N_4880,N_2455);
and U8512 (N_8512,N_453,N_4782);
nand U8513 (N_8513,N_912,N_4351);
and U8514 (N_8514,N_4518,N_1464);
xor U8515 (N_8515,N_2856,N_3182);
and U8516 (N_8516,N_250,N_322);
xor U8517 (N_8517,N_971,N_3256);
xor U8518 (N_8518,N_1312,N_3721);
xor U8519 (N_8519,N_2962,N_4275);
xor U8520 (N_8520,N_4715,N_4069);
xnor U8521 (N_8521,N_2652,N_1897);
and U8522 (N_8522,N_1807,N_1078);
or U8523 (N_8523,N_2034,N_145);
nor U8524 (N_8524,N_4407,N_305);
xnor U8525 (N_8525,N_2869,N_4570);
nor U8526 (N_8526,N_423,N_2490);
xor U8527 (N_8527,N_1061,N_3661);
or U8528 (N_8528,N_824,N_861);
xor U8529 (N_8529,N_1512,N_2852);
or U8530 (N_8530,N_2402,N_4766);
nand U8531 (N_8531,N_4991,N_4228);
nand U8532 (N_8532,N_2979,N_3726);
xor U8533 (N_8533,N_1505,N_1631);
nand U8534 (N_8534,N_2784,N_4501);
or U8535 (N_8535,N_520,N_1932);
and U8536 (N_8536,N_3776,N_267);
and U8537 (N_8537,N_3068,N_2017);
nand U8538 (N_8538,N_1784,N_4628);
or U8539 (N_8539,N_3235,N_2198);
nor U8540 (N_8540,N_3549,N_3480);
or U8541 (N_8541,N_3648,N_2838);
and U8542 (N_8542,N_2897,N_4666);
nor U8543 (N_8543,N_4006,N_3392);
nand U8544 (N_8544,N_4737,N_4227);
xnor U8545 (N_8545,N_24,N_4438);
and U8546 (N_8546,N_3716,N_3317);
and U8547 (N_8547,N_2697,N_2245);
nor U8548 (N_8548,N_4825,N_2761);
or U8549 (N_8549,N_2346,N_214);
nand U8550 (N_8550,N_2962,N_660);
and U8551 (N_8551,N_4061,N_1647);
or U8552 (N_8552,N_3165,N_2665);
nor U8553 (N_8553,N_965,N_2906);
nand U8554 (N_8554,N_1192,N_2459);
or U8555 (N_8555,N_3402,N_4806);
xor U8556 (N_8556,N_667,N_4987);
and U8557 (N_8557,N_2752,N_2345);
nand U8558 (N_8558,N_2358,N_937);
nor U8559 (N_8559,N_4817,N_809);
and U8560 (N_8560,N_4407,N_4937);
or U8561 (N_8561,N_4098,N_4594);
nand U8562 (N_8562,N_515,N_1235);
or U8563 (N_8563,N_2367,N_791);
nor U8564 (N_8564,N_4806,N_1934);
nor U8565 (N_8565,N_4010,N_730);
nor U8566 (N_8566,N_18,N_1283);
or U8567 (N_8567,N_2347,N_2703);
xnor U8568 (N_8568,N_4716,N_221);
nand U8569 (N_8569,N_3624,N_2871);
or U8570 (N_8570,N_21,N_468);
xor U8571 (N_8571,N_2422,N_465);
or U8572 (N_8572,N_4682,N_4819);
nand U8573 (N_8573,N_3825,N_832);
and U8574 (N_8574,N_1287,N_4044);
and U8575 (N_8575,N_679,N_4774);
xor U8576 (N_8576,N_3213,N_3795);
xnor U8577 (N_8577,N_840,N_140);
nand U8578 (N_8578,N_2419,N_3066);
nand U8579 (N_8579,N_2445,N_2610);
nor U8580 (N_8580,N_734,N_206);
nand U8581 (N_8581,N_2256,N_2442);
nor U8582 (N_8582,N_249,N_2125);
and U8583 (N_8583,N_2916,N_4320);
or U8584 (N_8584,N_1282,N_3809);
nand U8585 (N_8585,N_2325,N_1942);
xor U8586 (N_8586,N_3261,N_3810);
or U8587 (N_8587,N_726,N_3623);
or U8588 (N_8588,N_4848,N_4015);
or U8589 (N_8589,N_1796,N_3428);
or U8590 (N_8590,N_368,N_1498);
nand U8591 (N_8591,N_1377,N_2986);
xor U8592 (N_8592,N_2591,N_4096);
and U8593 (N_8593,N_4972,N_901);
and U8594 (N_8594,N_3902,N_1098);
nor U8595 (N_8595,N_769,N_3299);
nand U8596 (N_8596,N_649,N_509);
xnor U8597 (N_8597,N_121,N_4932);
nor U8598 (N_8598,N_4024,N_3224);
or U8599 (N_8599,N_2100,N_3535);
and U8600 (N_8600,N_2647,N_3563);
and U8601 (N_8601,N_1390,N_3484);
nand U8602 (N_8602,N_441,N_1209);
xor U8603 (N_8603,N_888,N_1649);
or U8604 (N_8604,N_4467,N_2137);
xnor U8605 (N_8605,N_4334,N_2422);
or U8606 (N_8606,N_2715,N_1225);
nor U8607 (N_8607,N_2621,N_75);
nand U8608 (N_8608,N_3124,N_2653);
and U8609 (N_8609,N_4565,N_3336);
xnor U8610 (N_8610,N_676,N_4853);
and U8611 (N_8611,N_2852,N_198);
nand U8612 (N_8612,N_3116,N_1721);
and U8613 (N_8613,N_4828,N_128);
or U8614 (N_8614,N_1993,N_4355);
nor U8615 (N_8615,N_2132,N_3187);
or U8616 (N_8616,N_705,N_1481);
nand U8617 (N_8617,N_4384,N_2254);
nor U8618 (N_8618,N_4778,N_907);
nand U8619 (N_8619,N_4488,N_2847);
xnor U8620 (N_8620,N_2692,N_674);
nand U8621 (N_8621,N_3005,N_220);
nand U8622 (N_8622,N_4333,N_3257);
nand U8623 (N_8623,N_3740,N_1875);
and U8624 (N_8624,N_4598,N_1430);
nand U8625 (N_8625,N_655,N_169);
xnor U8626 (N_8626,N_3833,N_3098);
and U8627 (N_8627,N_582,N_4794);
nand U8628 (N_8628,N_4750,N_973);
nand U8629 (N_8629,N_3403,N_109);
and U8630 (N_8630,N_4560,N_3505);
nor U8631 (N_8631,N_1454,N_116);
or U8632 (N_8632,N_899,N_1271);
nand U8633 (N_8633,N_90,N_4386);
or U8634 (N_8634,N_4555,N_1907);
nor U8635 (N_8635,N_2524,N_2289);
and U8636 (N_8636,N_4706,N_2568);
nor U8637 (N_8637,N_989,N_945);
xnor U8638 (N_8638,N_882,N_1440);
and U8639 (N_8639,N_2968,N_851);
nor U8640 (N_8640,N_2740,N_2722);
xnor U8641 (N_8641,N_4990,N_3691);
nand U8642 (N_8642,N_1356,N_1648);
nor U8643 (N_8643,N_4044,N_336);
nor U8644 (N_8644,N_603,N_1383);
xnor U8645 (N_8645,N_335,N_329);
nor U8646 (N_8646,N_4737,N_2927);
and U8647 (N_8647,N_3263,N_1359);
nand U8648 (N_8648,N_1695,N_4582);
nand U8649 (N_8649,N_287,N_474);
xnor U8650 (N_8650,N_4834,N_941);
and U8651 (N_8651,N_2129,N_4481);
xor U8652 (N_8652,N_4646,N_1732);
and U8653 (N_8653,N_1139,N_1400);
and U8654 (N_8654,N_1255,N_3433);
nand U8655 (N_8655,N_869,N_4543);
or U8656 (N_8656,N_281,N_510);
nand U8657 (N_8657,N_2241,N_891);
nand U8658 (N_8658,N_3396,N_2328);
xor U8659 (N_8659,N_4453,N_970);
and U8660 (N_8660,N_1077,N_2414);
and U8661 (N_8661,N_3401,N_1061);
and U8662 (N_8662,N_2958,N_2537);
nor U8663 (N_8663,N_3603,N_1241);
xnor U8664 (N_8664,N_2884,N_2063);
nor U8665 (N_8665,N_4366,N_1776);
xnor U8666 (N_8666,N_430,N_718);
or U8667 (N_8667,N_4515,N_1696);
nor U8668 (N_8668,N_855,N_4084);
nor U8669 (N_8669,N_3748,N_3292);
nor U8670 (N_8670,N_1904,N_3102);
nand U8671 (N_8671,N_2205,N_4379);
nor U8672 (N_8672,N_611,N_2795);
nand U8673 (N_8673,N_672,N_40);
nand U8674 (N_8674,N_2688,N_4588);
and U8675 (N_8675,N_4523,N_3854);
xor U8676 (N_8676,N_2697,N_822);
or U8677 (N_8677,N_2061,N_2379);
xor U8678 (N_8678,N_3684,N_98);
and U8679 (N_8679,N_3747,N_4343);
xor U8680 (N_8680,N_1817,N_321);
nand U8681 (N_8681,N_2318,N_1113);
xnor U8682 (N_8682,N_719,N_356);
nor U8683 (N_8683,N_3162,N_3129);
or U8684 (N_8684,N_3364,N_2535);
and U8685 (N_8685,N_2387,N_4327);
nand U8686 (N_8686,N_2645,N_2808);
nor U8687 (N_8687,N_1062,N_4357);
nor U8688 (N_8688,N_4924,N_4939);
nand U8689 (N_8689,N_2720,N_2986);
or U8690 (N_8690,N_2401,N_3445);
xor U8691 (N_8691,N_1548,N_4055);
or U8692 (N_8692,N_59,N_2325);
nor U8693 (N_8693,N_3942,N_2221);
xnor U8694 (N_8694,N_718,N_3073);
xnor U8695 (N_8695,N_4038,N_953);
or U8696 (N_8696,N_2825,N_1211);
and U8697 (N_8697,N_271,N_626);
nand U8698 (N_8698,N_929,N_353);
or U8699 (N_8699,N_1580,N_1066);
or U8700 (N_8700,N_1971,N_4576);
or U8701 (N_8701,N_4209,N_535);
xnor U8702 (N_8702,N_3404,N_3914);
xnor U8703 (N_8703,N_4926,N_847);
or U8704 (N_8704,N_4308,N_592);
nor U8705 (N_8705,N_2435,N_873);
and U8706 (N_8706,N_2062,N_4361);
and U8707 (N_8707,N_1165,N_4235);
or U8708 (N_8708,N_3609,N_2494);
nand U8709 (N_8709,N_2530,N_802);
nand U8710 (N_8710,N_804,N_3385);
or U8711 (N_8711,N_1277,N_1850);
nor U8712 (N_8712,N_2403,N_3108);
nor U8713 (N_8713,N_3621,N_1289);
xor U8714 (N_8714,N_3700,N_1179);
or U8715 (N_8715,N_558,N_209);
nand U8716 (N_8716,N_392,N_965);
nor U8717 (N_8717,N_4587,N_4017);
or U8718 (N_8718,N_367,N_4804);
nor U8719 (N_8719,N_2015,N_3681);
xor U8720 (N_8720,N_4257,N_1191);
nand U8721 (N_8721,N_386,N_2459);
or U8722 (N_8722,N_2355,N_4702);
and U8723 (N_8723,N_3462,N_3503);
and U8724 (N_8724,N_4601,N_1964);
xnor U8725 (N_8725,N_3469,N_2118);
nor U8726 (N_8726,N_3303,N_1420);
nor U8727 (N_8727,N_3438,N_654);
and U8728 (N_8728,N_2041,N_1493);
nand U8729 (N_8729,N_3716,N_2669);
or U8730 (N_8730,N_3905,N_515);
xor U8731 (N_8731,N_836,N_3437);
or U8732 (N_8732,N_2312,N_4718);
xnor U8733 (N_8733,N_2027,N_4077);
nor U8734 (N_8734,N_277,N_2321);
nor U8735 (N_8735,N_4402,N_801);
or U8736 (N_8736,N_2918,N_224);
or U8737 (N_8737,N_792,N_570);
xor U8738 (N_8738,N_4717,N_2577);
or U8739 (N_8739,N_4280,N_1007);
or U8740 (N_8740,N_1616,N_2748);
and U8741 (N_8741,N_1947,N_1694);
xor U8742 (N_8742,N_1431,N_646);
nand U8743 (N_8743,N_2772,N_3778);
xor U8744 (N_8744,N_3604,N_2255);
nor U8745 (N_8745,N_3579,N_3735);
nand U8746 (N_8746,N_3931,N_2166);
nand U8747 (N_8747,N_4696,N_655);
or U8748 (N_8748,N_1397,N_2341);
nand U8749 (N_8749,N_4647,N_1928);
and U8750 (N_8750,N_96,N_3933);
xnor U8751 (N_8751,N_3170,N_42);
nand U8752 (N_8752,N_4378,N_3513);
nand U8753 (N_8753,N_1149,N_962);
nand U8754 (N_8754,N_1565,N_3898);
or U8755 (N_8755,N_1085,N_1013);
xnor U8756 (N_8756,N_4668,N_2429);
or U8757 (N_8757,N_1103,N_210);
xnor U8758 (N_8758,N_1380,N_229);
xnor U8759 (N_8759,N_4924,N_3489);
or U8760 (N_8760,N_4424,N_2783);
nor U8761 (N_8761,N_171,N_1096);
or U8762 (N_8762,N_3564,N_2552);
xnor U8763 (N_8763,N_2058,N_3528);
nand U8764 (N_8764,N_2128,N_3055);
xor U8765 (N_8765,N_151,N_977);
or U8766 (N_8766,N_2917,N_4936);
and U8767 (N_8767,N_1394,N_2122);
and U8768 (N_8768,N_4015,N_1060);
nand U8769 (N_8769,N_2049,N_3215);
nor U8770 (N_8770,N_2206,N_1527);
or U8771 (N_8771,N_1840,N_330);
xor U8772 (N_8772,N_2458,N_4665);
xnor U8773 (N_8773,N_4053,N_28);
or U8774 (N_8774,N_1133,N_2126);
nor U8775 (N_8775,N_2639,N_275);
or U8776 (N_8776,N_4328,N_4264);
or U8777 (N_8777,N_3678,N_4132);
or U8778 (N_8778,N_1850,N_3951);
and U8779 (N_8779,N_4608,N_994);
xor U8780 (N_8780,N_3611,N_4972);
xnor U8781 (N_8781,N_2437,N_299);
nor U8782 (N_8782,N_2208,N_3104);
nor U8783 (N_8783,N_4832,N_1168);
and U8784 (N_8784,N_2430,N_2190);
xnor U8785 (N_8785,N_2557,N_3719);
nor U8786 (N_8786,N_2292,N_745);
xnor U8787 (N_8787,N_4430,N_4558);
xor U8788 (N_8788,N_4043,N_3885);
and U8789 (N_8789,N_2458,N_3830);
nor U8790 (N_8790,N_2333,N_2974);
xor U8791 (N_8791,N_3266,N_1082);
nor U8792 (N_8792,N_1916,N_902);
nor U8793 (N_8793,N_3199,N_4005);
nor U8794 (N_8794,N_3362,N_3686);
nor U8795 (N_8795,N_2089,N_2321);
xnor U8796 (N_8796,N_4768,N_3229);
nand U8797 (N_8797,N_4503,N_2515);
nor U8798 (N_8798,N_3159,N_4059);
nand U8799 (N_8799,N_3466,N_3741);
nor U8800 (N_8800,N_643,N_1990);
xnor U8801 (N_8801,N_4520,N_4266);
nand U8802 (N_8802,N_613,N_3943);
or U8803 (N_8803,N_3204,N_2014);
nor U8804 (N_8804,N_866,N_50);
or U8805 (N_8805,N_4701,N_907);
nor U8806 (N_8806,N_2442,N_4185);
and U8807 (N_8807,N_2217,N_4669);
nor U8808 (N_8808,N_4821,N_1157);
or U8809 (N_8809,N_31,N_436);
nor U8810 (N_8810,N_3262,N_1257);
nand U8811 (N_8811,N_1244,N_1358);
or U8812 (N_8812,N_3976,N_192);
nand U8813 (N_8813,N_3055,N_751);
nor U8814 (N_8814,N_68,N_1938);
or U8815 (N_8815,N_2011,N_214);
nand U8816 (N_8816,N_799,N_592);
and U8817 (N_8817,N_2814,N_1558);
or U8818 (N_8818,N_4090,N_4144);
or U8819 (N_8819,N_869,N_2855);
nor U8820 (N_8820,N_918,N_760);
nand U8821 (N_8821,N_3593,N_4044);
xnor U8822 (N_8822,N_3133,N_327);
nand U8823 (N_8823,N_468,N_3106);
xor U8824 (N_8824,N_595,N_4427);
xnor U8825 (N_8825,N_282,N_500);
nor U8826 (N_8826,N_1428,N_857);
nor U8827 (N_8827,N_3362,N_1345);
and U8828 (N_8828,N_1976,N_2766);
nand U8829 (N_8829,N_4998,N_23);
xnor U8830 (N_8830,N_2941,N_1711);
or U8831 (N_8831,N_3542,N_1374);
nand U8832 (N_8832,N_1282,N_4404);
nand U8833 (N_8833,N_774,N_538);
nand U8834 (N_8834,N_4575,N_483);
xor U8835 (N_8835,N_2727,N_1526);
xnor U8836 (N_8836,N_408,N_4761);
and U8837 (N_8837,N_288,N_4830);
or U8838 (N_8838,N_2133,N_1049);
or U8839 (N_8839,N_2409,N_2905);
nor U8840 (N_8840,N_278,N_3599);
nor U8841 (N_8841,N_3206,N_1621);
nand U8842 (N_8842,N_2390,N_1446);
nand U8843 (N_8843,N_1287,N_2412);
nand U8844 (N_8844,N_2731,N_3194);
nor U8845 (N_8845,N_2265,N_3857);
or U8846 (N_8846,N_3312,N_1894);
and U8847 (N_8847,N_4924,N_938);
or U8848 (N_8848,N_1536,N_1569);
or U8849 (N_8849,N_3918,N_3318);
or U8850 (N_8850,N_766,N_4430);
xor U8851 (N_8851,N_3345,N_3659);
or U8852 (N_8852,N_4023,N_4737);
nand U8853 (N_8853,N_913,N_1306);
xnor U8854 (N_8854,N_2454,N_1373);
nand U8855 (N_8855,N_1414,N_3346);
nor U8856 (N_8856,N_2786,N_4927);
xnor U8857 (N_8857,N_962,N_4906);
or U8858 (N_8858,N_359,N_4969);
nand U8859 (N_8859,N_3298,N_2484);
xor U8860 (N_8860,N_3851,N_3245);
nand U8861 (N_8861,N_3236,N_154);
xor U8862 (N_8862,N_2361,N_2567);
nand U8863 (N_8863,N_2537,N_4426);
xor U8864 (N_8864,N_1000,N_4800);
nand U8865 (N_8865,N_3184,N_37);
nor U8866 (N_8866,N_3202,N_400);
or U8867 (N_8867,N_1758,N_1546);
or U8868 (N_8868,N_2798,N_1008);
xor U8869 (N_8869,N_1681,N_2937);
and U8870 (N_8870,N_3128,N_3985);
or U8871 (N_8871,N_2486,N_694);
xnor U8872 (N_8872,N_4483,N_1637);
or U8873 (N_8873,N_3878,N_627);
and U8874 (N_8874,N_3961,N_3860);
and U8875 (N_8875,N_1214,N_4640);
xnor U8876 (N_8876,N_4658,N_628);
nand U8877 (N_8877,N_1664,N_4394);
and U8878 (N_8878,N_1425,N_1022);
nand U8879 (N_8879,N_3892,N_1722);
xnor U8880 (N_8880,N_3617,N_1817);
nor U8881 (N_8881,N_1633,N_4648);
or U8882 (N_8882,N_4224,N_1206);
or U8883 (N_8883,N_2365,N_4233);
nor U8884 (N_8884,N_508,N_4484);
xnor U8885 (N_8885,N_3226,N_4819);
nor U8886 (N_8886,N_4390,N_1510);
xnor U8887 (N_8887,N_2970,N_432);
nand U8888 (N_8888,N_3503,N_3255);
and U8889 (N_8889,N_4382,N_2045);
nand U8890 (N_8890,N_2527,N_1335);
nand U8891 (N_8891,N_1555,N_3252);
or U8892 (N_8892,N_3135,N_729);
xnor U8893 (N_8893,N_218,N_310);
or U8894 (N_8894,N_4363,N_2737);
nand U8895 (N_8895,N_1034,N_2899);
xor U8896 (N_8896,N_2472,N_357);
or U8897 (N_8897,N_1538,N_2158);
and U8898 (N_8898,N_51,N_2626);
xor U8899 (N_8899,N_3472,N_1742);
nand U8900 (N_8900,N_4986,N_682);
nand U8901 (N_8901,N_3565,N_1494);
or U8902 (N_8902,N_3718,N_2869);
and U8903 (N_8903,N_2889,N_4251);
xor U8904 (N_8904,N_2680,N_1738);
nor U8905 (N_8905,N_1098,N_4622);
nand U8906 (N_8906,N_392,N_2850);
nand U8907 (N_8907,N_79,N_3858);
nor U8908 (N_8908,N_3947,N_3097);
or U8909 (N_8909,N_2496,N_1087);
or U8910 (N_8910,N_2009,N_263);
and U8911 (N_8911,N_4501,N_3932);
xnor U8912 (N_8912,N_123,N_2548);
or U8913 (N_8913,N_4400,N_2579);
nor U8914 (N_8914,N_4998,N_1296);
nor U8915 (N_8915,N_785,N_556);
or U8916 (N_8916,N_4941,N_1974);
or U8917 (N_8917,N_1526,N_3639);
nand U8918 (N_8918,N_1333,N_4418);
xnor U8919 (N_8919,N_3002,N_254);
nand U8920 (N_8920,N_4467,N_3635);
nand U8921 (N_8921,N_1713,N_3004);
nand U8922 (N_8922,N_2645,N_155);
nand U8923 (N_8923,N_4670,N_2818);
or U8924 (N_8924,N_1238,N_3325);
xnor U8925 (N_8925,N_2610,N_2245);
and U8926 (N_8926,N_2334,N_947);
and U8927 (N_8927,N_3419,N_3436);
and U8928 (N_8928,N_2115,N_1807);
nand U8929 (N_8929,N_3926,N_4745);
or U8930 (N_8930,N_3783,N_1836);
or U8931 (N_8931,N_2257,N_1375);
nand U8932 (N_8932,N_2110,N_4074);
nand U8933 (N_8933,N_1090,N_3091);
nor U8934 (N_8934,N_3424,N_1742);
and U8935 (N_8935,N_3277,N_3382);
nand U8936 (N_8936,N_1162,N_1651);
nand U8937 (N_8937,N_3904,N_1412);
and U8938 (N_8938,N_4413,N_3744);
or U8939 (N_8939,N_4204,N_4470);
nor U8940 (N_8940,N_4918,N_3036);
nand U8941 (N_8941,N_4972,N_795);
xor U8942 (N_8942,N_4819,N_2786);
xor U8943 (N_8943,N_1448,N_3659);
or U8944 (N_8944,N_3990,N_1307);
nand U8945 (N_8945,N_931,N_3941);
nor U8946 (N_8946,N_2676,N_604);
nor U8947 (N_8947,N_1755,N_2996);
and U8948 (N_8948,N_2391,N_1003);
nor U8949 (N_8949,N_497,N_4617);
nand U8950 (N_8950,N_1978,N_4304);
xnor U8951 (N_8951,N_2749,N_4630);
xor U8952 (N_8952,N_2168,N_3521);
nand U8953 (N_8953,N_4295,N_4137);
or U8954 (N_8954,N_2103,N_2618);
xnor U8955 (N_8955,N_2721,N_1455);
xor U8956 (N_8956,N_1864,N_1083);
xnor U8957 (N_8957,N_3314,N_387);
xnor U8958 (N_8958,N_3956,N_3453);
or U8959 (N_8959,N_3870,N_4008);
xnor U8960 (N_8960,N_3283,N_704);
and U8961 (N_8961,N_3024,N_1551);
and U8962 (N_8962,N_3084,N_4283);
and U8963 (N_8963,N_659,N_4716);
or U8964 (N_8964,N_2331,N_754);
or U8965 (N_8965,N_1911,N_1451);
xor U8966 (N_8966,N_1659,N_3712);
xnor U8967 (N_8967,N_618,N_4174);
xnor U8968 (N_8968,N_3057,N_733);
nor U8969 (N_8969,N_3104,N_2940);
nor U8970 (N_8970,N_2322,N_4752);
xor U8971 (N_8971,N_4836,N_1111);
and U8972 (N_8972,N_3890,N_2439);
and U8973 (N_8973,N_765,N_1937);
nand U8974 (N_8974,N_3378,N_3499);
and U8975 (N_8975,N_2501,N_3591);
or U8976 (N_8976,N_3102,N_1976);
or U8977 (N_8977,N_2094,N_3471);
nand U8978 (N_8978,N_1741,N_19);
or U8979 (N_8979,N_1236,N_4556);
nor U8980 (N_8980,N_618,N_4724);
xnor U8981 (N_8981,N_776,N_3090);
nand U8982 (N_8982,N_3553,N_2207);
xor U8983 (N_8983,N_1116,N_2314);
nor U8984 (N_8984,N_4672,N_811);
nand U8985 (N_8985,N_538,N_4090);
or U8986 (N_8986,N_3231,N_3344);
nor U8987 (N_8987,N_3739,N_3823);
and U8988 (N_8988,N_4866,N_1061);
and U8989 (N_8989,N_2648,N_2535);
xnor U8990 (N_8990,N_1694,N_1148);
xnor U8991 (N_8991,N_528,N_1500);
nand U8992 (N_8992,N_2456,N_1511);
nor U8993 (N_8993,N_2593,N_1763);
nand U8994 (N_8994,N_1384,N_2736);
nor U8995 (N_8995,N_513,N_4454);
nand U8996 (N_8996,N_233,N_3057);
nand U8997 (N_8997,N_1503,N_2473);
nand U8998 (N_8998,N_2989,N_4674);
or U8999 (N_8999,N_1179,N_4228);
and U9000 (N_9000,N_2468,N_3792);
xnor U9001 (N_9001,N_2374,N_344);
xor U9002 (N_9002,N_4736,N_3698);
or U9003 (N_9003,N_2130,N_2658);
xnor U9004 (N_9004,N_3818,N_2427);
nand U9005 (N_9005,N_4097,N_4319);
or U9006 (N_9006,N_1716,N_1724);
xor U9007 (N_9007,N_4281,N_3490);
and U9008 (N_9008,N_521,N_1032);
and U9009 (N_9009,N_1210,N_887);
and U9010 (N_9010,N_3702,N_864);
or U9011 (N_9011,N_1463,N_1182);
or U9012 (N_9012,N_510,N_1338);
nand U9013 (N_9013,N_570,N_501);
nor U9014 (N_9014,N_2715,N_3800);
xnor U9015 (N_9015,N_62,N_3982);
or U9016 (N_9016,N_853,N_544);
nand U9017 (N_9017,N_1848,N_2255);
xnor U9018 (N_9018,N_4401,N_1689);
nor U9019 (N_9019,N_4137,N_2096);
nor U9020 (N_9020,N_4361,N_121);
nand U9021 (N_9021,N_1566,N_1261);
xor U9022 (N_9022,N_629,N_3526);
xnor U9023 (N_9023,N_3582,N_3884);
nor U9024 (N_9024,N_1313,N_4277);
xor U9025 (N_9025,N_4537,N_2175);
nor U9026 (N_9026,N_1941,N_212);
nand U9027 (N_9027,N_4000,N_1041);
or U9028 (N_9028,N_48,N_2729);
or U9029 (N_9029,N_1185,N_1941);
or U9030 (N_9030,N_954,N_3872);
nor U9031 (N_9031,N_2027,N_1134);
and U9032 (N_9032,N_869,N_4367);
xor U9033 (N_9033,N_3302,N_4601);
xor U9034 (N_9034,N_2012,N_4342);
xnor U9035 (N_9035,N_944,N_4595);
xor U9036 (N_9036,N_4232,N_1702);
nor U9037 (N_9037,N_925,N_4930);
xor U9038 (N_9038,N_104,N_1519);
nand U9039 (N_9039,N_3142,N_1979);
xnor U9040 (N_9040,N_3278,N_4377);
or U9041 (N_9041,N_3722,N_3923);
nand U9042 (N_9042,N_1290,N_3825);
or U9043 (N_9043,N_3232,N_4722);
or U9044 (N_9044,N_2812,N_1176);
or U9045 (N_9045,N_2292,N_886);
and U9046 (N_9046,N_3403,N_4027);
or U9047 (N_9047,N_3674,N_4424);
nor U9048 (N_9048,N_4872,N_529);
nor U9049 (N_9049,N_4580,N_272);
nor U9050 (N_9050,N_172,N_3944);
nor U9051 (N_9051,N_3343,N_184);
nand U9052 (N_9052,N_1692,N_2146);
or U9053 (N_9053,N_1701,N_83);
and U9054 (N_9054,N_2514,N_2321);
and U9055 (N_9055,N_4079,N_4716);
or U9056 (N_9056,N_1479,N_3043);
xor U9057 (N_9057,N_4526,N_1659);
nor U9058 (N_9058,N_2875,N_3047);
and U9059 (N_9059,N_4383,N_658);
nand U9060 (N_9060,N_50,N_3528);
nand U9061 (N_9061,N_4860,N_4711);
nor U9062 (N_9062,N_1634,N_2429);
and U9063 (N_9063,N_4551,N_2735);
or U9064 (N_9064,N_2795,N_4104);
and U9065 (N_9065,N_3967,N_3478);
xnor U9066 (N_9066,N_420,N_691);
xnor U9067 (N_9067,N_1299,N_4558);
xor U9068 (N_9068,N_2009,N_1870);
xor U9069 (N_9069,N_3209,N_1479);
nor U9070 (N_9070,N_1706,N_2503);
xnor U9071 (N_9071,N_2394,N_564);
nand U9072 (N_9072,N_3536,N_4207);
nand U9073 (N_9073,N_4779,N_633);
nor U9074 (N_9074,N_106,N_471);
and U9075 (N_9075,N_4624,N_686);
xnor U9076 (N_9076,N_525,N_3838);
and U9077 (N_9077,N_3316,N_1421);
nand U9078 (N_9078,N_4624,N_4890);
xor U9079 (N_9079,N_1071,N_2287);
nand U9080 (N_9080,N_3946,N_1242);
xor U9081 (N_9081,N_2429,N_2615);
or U9082 (N_9082,N_2468,N_107);
nor U9083 (N_9083,N_4495,N_615);
xnor U9084 (N_9084,N_3506,N_2568);
or U9085 (N_9085,N_4344,N_2794);
nor U9086 (N_9086,N_4822,N_801);
and U9087 (N_9087,N_4525,N_125);
nor U9088 (N_9088,N_1544,N_4161);
nor U9089 (N_9089,N_1832,N_3944);
nand U9090 (N_9090,N_219,N_1098);
nand U9091 (N_9091,N_14,N_2962);
nand U9092 (N_9092,N_4555,N_2228);
or U9093 (N_9093,N_2841,N_2777);
or U9094 (N_9094,N_2547,N_104);
nor U9095 (N_9095,N_3960,N_1273);
and U9096 (N_9096,N_1838,N_2125);
or U9097 (N_9097,N_2650,N_806);
nor U9098 (N_9098,N_3833,N_171);
and U9099 (N_9099,N_3106,N_4773);
xnor U9100 (N_9100,N_217,N_2661);
and U9101 (N_9101,N_2549,N_4070);
and U9102 (N_9102,N_847,N_4221);
xor U9103 (N_9103,N_4229,N_3429);
nand U9104 (N_9104,N_3979,N_3464);
nor U9105 (N_9105,N_1792,N_4643);
and U9106 (N_9106,N_3734,N_4188);
nand U9107 (N_9107,N_2019,N_2945);
nor U9108 (N_9108,N_201,N_3252);
nor U9109 (N_9109,N_3500,N_1456);
or U9110 (N_9110,N_114,N_1196);
or U9111 (N_9111,N_843,N_1751);
and U9112 (N_9112,N_4071,N_2137);
nor U9113 (N_9113,N_2233,N_781);
and U9114 (N_9114,N_2630,N_4283);
or U9115 (N_9115,N_1728,N_777);
and U9116 (N_9116,N_1609,N_1138);
xor U9117 (N_9117,N_3369,N_2490);
or U9118 (N_9118,N_2439,N_3602);
xnor U9119 (N_9119,N_4896,N_3724);
nand U9120 (N_9120,N_4675,N_2091);
xnor U9121 (N_9121,N_4358,N_2340);
nor U9122 (N_9122,N_1268,N_1563);
nor U9123 (N_9123,N_1945,N_4478);
and U9124 (N_9124,N_3854,N_3845);
and U9125 (N_9125,N_3532,N_4387);
nor U9126 (N_9126,N_1357,N_4319);
nand U9127 (N_9127,N_424,N_1459);
and U9128 (N_9128,N_1785,N_417);
nor U9129 (N_9129,N_2585,N_1829);
and U9130 (N_9130,N_1786,N_1719);
xnor U9131 (N_9131,N_354,N_4635);
xor U9132 (N_9132,N_1703,N_1292);
nand U9133 (N_9133,N_209,N_2400);
xor U9134 (N_9134,N_1798,N_3126);
and U9135 (N_9135,N_2221,N_2747);
nand U9136 (N_9136,N_4713,N_4177);
and U9137 (N_9137,N_412,N_4310);
nand U9138 (N_9138,N_4013,N_1674);
nand U9139 (N_9139,N_4620,N_4948);
and U9140 (N_9140,N_2168,N_4337);
nand U9141 (N_9141,N_610,N_2678);
nor U9142 (N_9142,N_1284,N_4942);
or U9143 (N_9143,N_1059,N_3576);
nand U9144 (N_9144,N_626,N_88);
nand U9145 (N_9145,N_950,N_3439);
and U9146 (N_9146,N_4790,N_1567);
nor U9147 (N_9147,N_1894,N_907);
or U9148 (N_9148,N_4355,N_2904);
and U9149 (N_9149,N_445,N_3561);
and U9150 (N_9150,N_1041,N_1505);
nand U9151 (N_9151,N_1424,N_4678);
nor U9152 (N_9152,N_619,N_2953);
nor U9153 (N_9153,N_2423,N_2772);
and U9154 (N_9154,N_379,N_222);
xnor U9155 (N_9155,N_4324,N_136);
xnor U9156 (N_9156,N_801,N_2176);
nor U9157 (N_9157,N_4894,N_3298);
nor U9158 (N_9158,N_3711,N_837);
nand U9159 (N_9159,N_3157,N_4346);
or U9160 (N_9160,N_2372,N_3584);
nand U9161 (N_9161,N_2175,N_3187);
nor U9162 (N_9162,N_1775,N_3415);
xor U9163 (N_9163,N_831,N_3538);
nor U9164 (N_9164,N_1703,N_2337);
or U9165 (N_9165,N_1962,N_4882);
nor U9166 (N_9166,N_4893,N_2484);
or U9167 (N_9167,N_1586,N_2688);
nor U9168 (N_9168,N_3352,N_254);
xor U9169 (N_9169,N_4337,N_1392);
nor U9170 (N_9170,N_2973,N_1968);
and U9171 (N_9171,N_3787,N_1300);
xnor U9172 (N_9172,N_2392,N_4377);
nand U9173 (N_9173,N_1834,N_1749);
nand U9174 (N_9174,N_3664,N_3021);
nor U9175 (N_9175,N_723,N_789);
nor U9176 (N_9176,N_2975,N_1660);
xnor U9177 (N_9177,N_2223,N_169);
xnor U9178 (N_9178,N_3671,N_3282);
nand U9179 (N_9179,N_4384,N_1621);
nor U9180 (N_9180,N_2014,N_3989);
nand U9181 (N_9181,N_2779,N_2270);
nor U9182 (N_9182,N_3121,N_4700);
and U9183 (N_9183,N_3840,N_4979);
nor U9184 (N_9184,N_4182,N_534);
and U9185 (N_9185,N_4514,N_486);
and U9186 (N_9186,N_4451,N_1978);
nor U9187 (N_9187,N_3523,N_4901);
nand U9188 (N_9188,N_221,N_2343);
or U9189 (N_9189,N_1812,N_2156);
xnor U9190 (N_9190,N_520,N_4332);
nor U9191 (N_9191,N_678,N_4970);
xor U9192 (N_9192,N_770,N_1964);
or U9193 (N_9193,N_740,N_2301);
and U9194 (N_9194,N_781,N_283);
xnor U9195 (N_9195,N_4395,N_3223);
and U9196 (N_9196,N_2244,N_4060);
nand U9197 (N_9197,N_3220,N_3362);
and U9198 (N_9198,N_4465,N_1354);
or U9199 (N_9199,N_4271,N_2156);
or U9200 (N_9200,N_4410,N_4289);
and U9201 (N_9201,N_375,N_4940);
and U9202 (N_9202,N_1618,N_4134);
and U9203 (N_9203,N_2323,N_1169);
xnor U9204 (N_9204,N_948,N_1501);
or U9205 (N_9205,N_1939,N_2774);
and U9206 (N_9206,N_249,N_414);
xor U9207 (N_9207,N_4887,N_594);
nor U9208 (N_9208,N_743,N_689);
or U9209 (N_9209,N_1520,N_1327);
nor U9210 (N_9210,N_640,N_2397);
nand U9211 (N_9211,N_3044,N_1485);
or U9212 (N_9212,N_4439,N_2204);
or U9213 (N_9213,N_4650,N_237);
and U9214 (N_9214,N_2604,N_1350);
or U9215 (N_9215,N_1488,N_4990);
nor U9216 (N_9216,N_408,N_1890);
and U9217 (N_9217,N_2740,N_874);
nor U9218 (N_9218,N_1633,N_48);
and U9219 (N_9219,N_4020,N_2397);
nand U9220 (N_9220,N_4871,N_2196);
nand U9221 (N_9221,N_3450,N_2409);
and U9222 (N_9222,N_2856,N_339);
and U9223 (N_9223,N_2482,N_2516);
and U9224 (N_9224,N_407,N_848);
nand U9225 (N_9225,N_3708,N_1648);
xor U9226 (N_9226,N_3583,N_819);
nor U9227 (N_9227,N_474,N_2828);
and U9228 (N_9228,N_4085,N_2625);
nor U9229 (N_9229,N_325,N_2891);
nor U9230 (N_9230,N_2432,N_1041);
or U9231 (N_9231,N_714,N_4372);
xor U9232 (N_9232,N_1428,N_3457);
or U9233 (N_9233,N_4845,N_1743);
and U9234 (N_9234,N_4916,N_3878);
and U9235 (N_9235,N_215,N_3382);
and U9236 (N_9236,N_684,N_598);
nor U9237 (N_9237,N_3118,N_358);
or U9238 (N_9238,N_2608,N_2265);
nand U9239 (N_9239,N_891,N_1302);
nand U9240 (N_9240,N_2214,N_2793);
xor U9241 (N_9241,N_4271,N_1209);
nor U9242 (N_9242,N_1236,N_305);
nand U9243 (N_9243,N_1293,N_58);
and U9244 (N_9244,N_2296,N_1861);
nand U9245 (N_9245,N_3801,N_2009);
xor U9246 (N_9246,N_4623,N_2490);
and U9247 (N_9247,N_1190,N_2852);
nor U9248 (N_9248,N_1536,N_2938);
xnor U9249 (N_9249,N_852,N_1459);
nand U9250 (N_9250,N_237,N_615);
xnor U9251 (N_9251,N_2669,N_3577);
xnor U9252 (N_9252,N_704,N_106);
or U9253 (N_9253,N_451,N_398);
xor U9254 (N_9254,N_3996,N_1583);
and U9255 (N_9255,N_2615,N_3553);
or U9256 (N_9256,N_2950,N_2798);
xor U9257 (N_9257,N_3801,N_4546);
nor U9258 (N_9258,N_3981,N_1550);
xor U9259 (N_9259,N_494,N_2233);
xnor U9260 (N_9260,N_2444,N_4390);
nand U9261 (N_9261,N_1998,N_1798);
nand U9262 (N_9262,N_566,N_4936);
or U9263 (N_9263,N_1244,N_698);
and U9264 (N_9264,N_4743,N_4427);
nand U9265 (N_9265,N_1529,N_966);
nand U9266 (N_9266,N_1123,N_3748);
nand U9267 (N_9267,N_3317,N_1489);
and U9268 (N_9268,N_4248,N_4690);
nand U9269 (N_9269,N_949,N_3840);
xnor U9270 (N_9270,N_1646,N_1774);
nand U9271 (N_9271,N_1160,N_4465);
or U9272 (N_9272,N_2532,N_3772);
nand U9273 (N_9273,N_3871,N_1065);
xor U9274 (N_9274,N_1469,N_718);
xnor U9275 (N_9275,N_1304,N_4490);
nand U9276 (N_9276,N_2926,N_157);
xor U9277 (N_9277,N_3907,N_1078);
nand U9278 (N_9278,N_3855,N_4538);
xnor U9279 (N_9279,N_3847,N_244);
or U9280 (N_9280,N_2359,N_4547);
nor U9281 (N_9281,N_2741,N_3599);
nor U9282 (N_9282,N_2629,N_4847);
nor U9283 (N_9283,N_4461,N_2626);
xnor U9284 (N_9284,N_758,N_2683);
xor U9285 (N_9285,N_2972,N_2830);
xor U9286 (N_9286,N_698,N_2127);
or U9287 (N_9287,N_2817,N_1515);
xor U9288 (N_9288,N_2087,N_3517);
nor U9289 (N_9289,N_2816,N_4562);
or U9290 (N_9290,N_1057,N_2733);
nor U9291 (N_9291,N_1839,N_4424);
nand U9292 (N_9292,N_1142,N_905);
xnor U9293 (N_9293,N_3968,N_2197);
xnor U9294 (N_9294,N_4009,N_2726);
nor U9295 (N_9295,N_1387,N_206);
xnor U9296 (N_9296,N_3906,N_781);
xor U9297 (N_9297,N_3734,N_4634);
nand U9298 (N_9298,N_2919,N_3510);
or U9299 (N_9299,N_2882,N_1538);
and U9300 (N_9300,N_4248,N_4640);
nand U9301 (N_9301,N_1169,N_2389);
nand U9302 (N_9302,N_4548,N_3414);
xnor U9303 (N_9303,N_561,N_948);
or U9304 (N_9304,N_4102,N_3076);
nand U9305 (N_9305,N_1357,N_1313);
or U9306 (N_9306,N_143,N_2426);
nand U9307 (N_9307,N_2229,N_2017);
xnor U9308 (N_9308,N_4002,N_4775);
and U9309 (N_9309,N_2872,N_277);
nand U9310 (N_9310,N_1278,N_2412);
xor U9311 (N_9311,N_1540,N_3344);
or U9312 (N_9312,N_3713,N_2231);
nand U9313 (N_9313,N_1241,N_3539);
or U9314 (N_9314,N_4245,N_1847);
or U9315 (N_9315,N_4298,N_3770);
and U9316 (N_9316,N_4242,N_3116);
nand U9317 (N_9317,N_1888,N_4499);
nand U9318 (N_9318,N_4717,N_4783);
nand U9319 (N_9319,N_3610,N_1373);
and U9320 (N_9320,N_2310,N_4176);
and U9321 (N_9321,N_4349,N_2143);
xor U9322 (N_9322,N_3267,N_4586);
nand U9323 (N_9323,N_2464,N_4594);
or U9324 (N_9324,N_3714,N_108);
xor U9325 (N_9325,N_3229,N_3110);
or U9326 (N_9326,N_1941,N_391);
nor U9327 (N_9327,N_2226,N_4662);
nand U9328 (N_9328,N_1599,N_74);
nor U9329 (N_9329,N_1292,N_2022);
and U9330 (N_9330,N_3082,N_116);
nand U9331 (N_9331,N_2806,N_3766);
xor U9332 (N_9332,N_1174,N_2111);
or U9333 (N_9333,N_2455,N_4725);
nor U9334 (N_9334,N_408,N_3402);
nand U9335 (N_9335,N_2370,N_3252);
xor U9336 (N_9336,N_4278,N_1930);
nand U9337 (N_9337,N_1818,N_875);
and U9338 (N_9338,N_1593,N_3306);
nand U9339 (N_9339,N_3270,N_2054);
and U9340 (N_9340,N_39,N_4490);
and U9341 (N_9341,N_361,N_2650);
nand U9342 (N_9342,N_3458,N_4942);
or U9343 (N_9343,N_2568,N_2990);
xor U9344 (N_9344,N_715,N_4628);
nor U9345 (N_9345,N_3465,N_3612);
nor U9346 (N_9346,N_1523,N_4021);
and U9347 (N_9347,N_2455,N_2118);
and U9348 (N_9348,N_1507,N_2881);
nor U9349 (N_9349,N_4573,N_2097);
xor U9350 (N_9350,N_811,N_981);
nor U9351 (N_9351,N_164,N_4813);
nor U9352 (N_9352,N_364,N_3448);
nand U9353 (N_9353,N_253,N_36);
and U9354 (N_9354,N_481,N_1857);
xnor U9355 (N_9355,N_3833,N_3918);
nor U9356 (N_9356,N_4292,N_371);
nand U9357 (N_9357,N_4443,N_1682);
xor U9358 (N_9358,N_279,N_2456);
xor U9359 (N_9359,N_1746,N_791);
nand U9360 (N_9360,N_1657,N_2978);
or U9361 (N_9361,N_2216,N_1940);
or U9362 (N_9362,N_1356,N_2617);
or U9363 (N_9363,N_5,N_4575);
and U9364 (N_9364,N_2283,N_1402);
xor U9365 (N_9365,N_4957,N_172);
and U9366 (N_9366,N_2055,N_2586);
or U9367 (N_9367,N_582,N_2162);
nand U9368 (N_9368,N_2330,N_1339);
or U9369 (N_9369,N_3770,N_1371);
nand U9370 (N_9370,N_326,N_142);
or U9371 (N_9371,N_4690,N_4660);
xor U9372 (N_9372,N_3455,N_3559);
nor U9373 (N_9373,N_1050,N_114);
nor U9374 (N_9374,N_4937,N_3368);
xnor U9375 (N_9375,N_194,N_1721);
and U9376 (N_9376,N_2829,N_2970);
and U9377 (N_9377,N_1775,N_2950);
nand U9378 (N_9378,N_462,N_4835);
xor U9379 (N_9379,N_2135,N_2702);
nand U9380 (N_9380,N_886,N_876);
and U9381 (N_9381,N_786,N_3512);
or U9382 (N_9382,N_2499,N_391);
nor U9383 (N_9383,N_4127,N_2577);
nand U9384 (N_9384,N_2502,N_2746);
or U9385 (N_9385,N_1586,N_4543);
nand U9386 (N_9386,N_2005,N_3947);
nand U9387 (N_9387,N_4733,N_4247);
or U9388 (N_9388,N_2047,N_4501);
xor U9389 (N_9389,N_4286,N_3038);
xor U9390 (N_9390,N_2044,N_4753);
xor U9391 (N_9391,N_1759,N_1215);
nor U9392 (N_9392,N_875,N_1816);
and U9393 (N_9393,N_2240,N_2753);
xnor U9394 (N_9394,N_4096,N_4700);
xor U9395 (N_9395,N_1154,N_3192);
nor U9396 (N_9396,N_1230,N_2112);
or U9397 (N_9397,N_3638,N_2468);
nand U9398 (N_9398,N_2697,N_4531);
or U9399 (N_9399,N_1278,N_2438);
xnor U9400 (N_9400,N_1873,N_2698);
and U9401 (N_9401,N_425,N_4873);
xor U9402 (N_9402,N_2125,N_4948);
and U9403 (N_9403,N_2614,N_734);
nor U9404 (N_9404,N_4418,N_2241);
or U9405 (N_9405,N_1823,N_3521);
xor U9406 (N_9406,N_3969,N_4354);
xnor U9407 (N_9407,N_2310,N_2226);
and U9408 (N_9408,N_1192,N_3223);
and U9409 (N_9409,N_1630,N_3537);
nand U9410 (N_9410,N_3260,N_3880);
nand U9411 (N_9411,N_1857,N_4510);
or U9412 (N_9412,N_4282,N_4789);
and U9413 (N_9413,N_1489,N_4152);
and U9414 (N_9414,N_3054,N_3056);
nor U9415 (N_9415,N_1772,N_3145);
xor U9416 (N_9416,N_4623,N_677);
nor U9417 (N_9417,N_1175,N_3018);
nor U9418 (N_9418,N_3006,N_4378);
nand U9419 (N_9419,N_1480,N_2877);
nor U9420 (N_9420,N_481,N_2771);
and U9421 (N_9421,N_1949,N_3050);
nand U9422 (N_9422,N_3933,N_1110);
or U9423 (N_9423,N_2620,N_2297);
xnor U9424 (N_9424,N_4179,N_1483);
and U9425 (N_9425,N_3645,N_1149);
xnor U9426 (N_9426,N_65,N_2916);
or U9427 (N_9427,N_339,N_1721);
or U9428 (N_9428,N_4917,N_2506);
nor U9429 (N_9429,N_1112,N_2630);
and U9430 (N_9430,N_3997,N_3376);
nor U9431 (N_9431,N_4406,N_1029);
nand U9432 (N_9432,N_82,N_506);
nor U9433 (N_9433,N_2644,N_1086);
nand U9434 (N_9434,N_908,N_2565);
nand U9435 (N_9435,N_513,N_4584);
nand U9436 (N_9436,N_1308,N_1901);
nand U9437 (N_9437,N_450,N_1006);
and U9438 (N_9438,N_3272,N_748);
and U9439 (N_9439,N_1365,N_1537);
nand U9440 (N_9440,N_98,N_2661);
and U9441 (N_9441,N_3779,N_4392);
xor U9442 (N_9442,N_3587,N_1771);
and U9443 (N_9443,N_683,N_1089);
xor U9444 (N_9444,N_1583,N_2362);
nand U9445 (N_9445,N_3828,N_2851);
or U9446 (N_9446,N_237,N_4095);
xor U9447 (N_9447,N_2932,N_4198);
nor U9448 (N_9448,N_3856,N_2792);
nand U9449 (N_9449,N_2632,N_3798);
xnor U9450 (N_9450,N_911,N_2395);
and U9451 (N_9451,N_513,N_929);
xnor U9452 (N_9452,N_3701,N_4241);
nor U9453 (N_9453,N_4236,N_898);
xnor U9454 (N_9454,N_1344,N_1765);
xnor U9455 (N_9455,N_2300,N_4019);
and U9456 (N_9456,N_643,N_2881);
and U9457 (N_9457,N_2733,N_113);
xnor U9458 (N_9458,N_2435,N_2834);
or U9459 (N_9459,N_721,N_2101);
nor U9460 (N_9460,N_1686,N_454);
xor U9461 (N_9461,N_3410,N_3645);
or U9462 (N_9462,N_2052,N_3928);
nand U9463 (N_9463,N_3284,N_1679);
nand U9464 (N_9464,N_1407,N_3843);
nor U9465 (N_9465,N_3465,N_2317);
nand U9466 (N_9466,N_2172,N_2438);
xnor U9467 (N_9467,N_3022,N_2278);
nor U9468 (N_9468,N_4060,N_1644);
nand U9469 (N_9469,N_2001,N_62);
nand U9470 (N_9470,N_1468,N_3435);
nand U9471 (N_9471,N_754,N_4731);
nor U9472 (N_9472,N_706,N_452);
xnor U9473 (N_9473,N_2226,N_1996);
nor U9474 (N_9474,N_3789,N_2580);
nand U9475 (N_9475,N_1565,N_301);
nor U9476 (N_9476,N_3062,N_4752);
nand U9477 (N_9477,N_839,N_2664);
nand U9478 (N_9478,N_3927,N_3419);
xor U9479 (N_9479,N_959,N_2955);
nor U9480 (N_9480,N_4879,N_3987);
xnor U9481 (N_9481,N_2755,N_1160);
nor U9482 (N_9482,N_1536,N_2667);
xor U9483 (N_9483,N_4735,N_4770);
xnor U9484 (N_9484,N_3004,N_3719);
and U9485 (N_9485,N_3334,N_2620);
xor U9486 (N_9486,N_3688,N_2265);
nand U9487 (N_9487,N_4284,N_2640);
and U9488 (N_9488,N_4719,N_3233);
and U9489 (N_9489,N_1734,N_684);
nand U9490 (N_9490,N_3163,N_2989);
xor U9491 (N_9491,N_3552,N_1357);
nand U9492 (N_9492,N_1856,N_3090);
or U9493 (N_9493,N_1466,N_533);
nor U9494 (N_9494,N_3068,N_2653);
nor U9495 (N_9495,N_4099,N_3882);
nor U9496 (N_9496,N_1610,N_318);
nand U9497 (N_9497,N_4556,N_540);
nor U9498 (N_9498,N_4730,N_3767);
nand U9499 (N_9499,N_4758,N_3422);
nor U9500 (N_9500,N_1913,N_4602);
nand U9501 (N_9501,N_1771,N_3170);
nand U9502 (N_9502,N_1264,N_4612);
nand U9503 (N_9503,N_3384,N_3923);
nor U9504 (N_9504,N_2108,N_4333);
xnor U9505 (N_9505,N_1741,N_3921);
xor U9506 (N_9506,N_1195,N_2668);
xor U9507 (N_9507,N_3774,N_1946);
and U9508 (N_9508,N_1823,N_610);
xnor U9509 (N_9509,N_3821,N_2791);
nor U9510 (N_9510,N_4996,N_1177);
xnor U9511 (N_9511,N_341,N_3079);
nand U9512 (N_9512,N_3535,N_3463);
nand U9513 (N_9513,N_4518,N_4893);
xor U9514 (N_9514,N_509,N_1777);
or U9515 (N_9515,N_747,N_1445);
or U9516 (N_9516,N_3375,N_1977);
or U9517 (N_9517,N_3323,N_4691);
and U9518 (N_9518,N_4677,N_3331);
nand U9519 (N_9519,N_3294,N_3828);
nand U9520 (N_9520,N_1573,N_1480);
nand U9521 (N_9521,N_4946,N_1968);
nand U9522 (N_9522,N_2361,N_2301);
or U9523 (N_9523,N_4828,N_582);
or U9524 (N_9524,N_4699,N_2961);
and U9525 (N_9525,N_2858,N_2800);
or U9526 (N_9526,N_649,N_4897);
xor U9527 (N_9527,N_1293,N_2472);
xor U9528 (N_9528,N_2899,N_1285);
or U9529 (N_9529,N_506,N_4063);
nor U9530 (N_9530,N_4418,N_4976);
nor U9531 (N_9531,N_2055,N_1570);
or U9532 (N_9532,N_4165,N_3615);
xnor U9533 (N_9533,N_3295,N_1276);
nand U9534 (N_9534,N_1727,N_4771);
nand U9535 (N_9535,N_389,N_2436);
nand U9536 (N_9536,N_1726,N_4191);
nor U9537 (N_9537,N_4087,N_2252);
xor U9538 (N_9538,N_4942,N_4837);
and U9539 (N_9539,N_3497,N_542);
nor U9540 (N_9540,N_2333,N_3835);
nand U9541 (N_9541,N_1155,N_1483);
and U9542 (N_9542,N_2895,N_3375);
or U9543 (N_9543,N_3353,N_4603);
and U9544 (N_9544,N_1920,N_355);
nand U9545 (N_9545,N_72,N_3019);
nor U9546 (N_9546,N_3432,N_2812);
nand U9547 (N_9547,N_3568,N_3201);
xnor U9548 (N_9548,N_1002,N_4986);
nor U9549 (N_9549,N_4477,N_3150);
or U9550 (N_9550,N_3001,N_3574);
or U9551 (N_9551,N_345,N_1635);
or U9552 (N_9552,N_126,N_3371);
and U9553 (N_9553,N_4680,N_272);
nand U9554 (N_9554,N_3541,N_976);
nand U9555 (N_9555,N_3433,N_4816);
and U9556 (N_9556,N_3939,N_1550);
nand U9557 (N_9557,N_3427,N_1704);
nand U9558 (N_9558,N_4634,N_3389);
nor U9559 (N_9559,N_1334,N_3040);
and U9560 (N_9560,N_4930,N_2685);
nand U9561 (N_9561,N_1202,N_1137);
or U9562 (N_9562,N_1786,N_1754);
nor U9563 (N_9563,N_2533,N_720);
nand U9564 (N_9564,N_1806,N_2284);
nor U9565 (N_9565,N_4589,N_148);
and U9566 (N_9566,N_1160,N_4844);
nor U9567 (N_9567,N_1216,N_3992);
nand U9568 (N_9568,N_1982,N_2379);
nand U9569 (N_9569,N_4150,N_2437);
and U9570 (N_9570,N_4550,N_3460);
xor U9571 (N_9571,N_629,N_1285);
xnor U9572 (N_9572,N_2892,N_2255);
xnor U9573 (N_9573,N_1894,N_3296);
or U9574 (N_9574,N_3708,N_543);
or U9575 (N_9575,N_3678,N_4050);
xor U9576 (N_9576,N_34,N_2621);
xor U9577 (N_9577,N_2093,N_58);
nand U9578 (N_9578,N_2921,N_1686);
or U9579 (N_9579,N_4451,N_4318);
nor U9580 (N_9580,N_1271,N_4116);
nor U9581 (N_9581,N_2507,N_908);
nor U9582 (N_9582,N_826,N_1151);
or U9583 (N_9583,N_1024,N_1632);
nor U9584 (N_9584,N_1927,N_4444);
or U9585 (N_9585,N_3876,N_2738);
and U9586 (N_9586,N_3554,N_2021);
nor U9587 (N_9587,N_4384,N_1379);
xnor U9588 (N_9588,N_1350,N_179);
nand U9589 (N_9589,N_1107,N_4895);
nor U9590 (N_9590,N_1946,N_51);
xnor U9591 (N_9591,N_4030,N_3300);
and U9592 (N_9592,N_3226,N_1724);
xnor U9593 (N_9593,N_152,N_4249);
nand U9594 (N_9594,N_173,N_2417);
xnor U9595 (N_9595,N_2710,N_3696);
xnor U9596 (N_9596,N_158,N_4737);
or U9597 (N_9597,N_1692,N_4673);
xor U9598 (N_9598,N_535,N_3746);
xor U9599 (N_9599,N_551,N_4482);
xor U9600 (N_9600,N_4773,N_2880);
nand U9601 (N_9601,N_1065,N_3866);
nand U9602 (N_9602,N_3919,N_4156);
nor U9603 (N_9603,N_2520,N_95);
nand U9604 (N_9604,N_2422,N_4183);
or U9605 (N_9605,N_4556,N_173);
and U9606 (N_9606,N_1082,N_845);
nor U9607 (N_9607,N_4440,N_1712);
and U9608 (N_9608,N_2270,N_2720);
xor U9609 (N_9609,N_1991,N_2558);
nand U9610 (N_9610,N_3110,N_4909);
xnor U9611 (N_9611,N_4506,N_992);
and U9612 (N_9612,N_4454,N_3614);
xor U9613 (N_9613,N_613,N_3424);
and U9614 (N_9614,N_1420,N_389);
and U9615 (N_9615,N_4363,N_3594);
or U9616 (N_9616,N_950,N_3934);
nand U9617 (N_9617,N_171,N_2319);
or U9618 (N_9618,N_1227,N_2563);
xnor U9619 (N_9619,N_4054,N_1973);
nor U9620 (N_9620,N_1167,N_2574);
nor U9621 (N_9621,N_2181,N_442);
nand U9622 (N_9622,N_459,N_822);
nor U9623 (N_9623,N_3921,N_3077);
xor U9624 (N_9624,N_2147,N_459);
nand U9625 (N_9625,N_2490,N_3209);
and U9626 (N_9626,N_1211,N_615);
and U9627 (N_9627,N_673,N_123);
nor U9628 (N_9628,N_3408,N_572);
or U9629 (N_9629,N_1690,N_2078);
xnor U9630 (N_9630,N_4552,N_367);
xor U9631 (N_9631,N_4723,N_2158);
and U9632 (N_9632,N_4841,N_3904);
xnor U9633 (N_9633,N_2069,N_1946);
or U9634 (N_9634,N_2805,N_649);
nor U9635 (N_9635,N_2594,N_2300);
xnor U9636 (N_9636,N_1221,N_3884);
xnor U9637 (N_9637,N_4817,N_1193);
xor U9638 (N_9638,N_3180,N_2869);
and U9639 (N_9639,N_14,N_2606);
or U9640 (N_9640,N_2953,N_833);
nand U9641 (N_9641,N_4852,N_4108);
or U9642 (N_9642,N_658,N_1482);
nand U9643 (N_9643,N_307,N_3782);
and U9644 (N_9644,N_3447,N_457);
nand U9645 (N_9645,N_331,N_3713);
nand U9646 (N_9646,N_3701,N_2289);
xor U9647 (N_9647,N_1439,N_3957);
and U9648 (N_9648,N_896,N_3558);
nor U9649 (N_9649,N_4463,N_4686);
nor U9650 (N_9650,N_252,N_2056);
xor U9651 (N_9651,N_3597,N_3743);
nor U9652 (N_9652,N_779,N_1846);
nor U9653 (N_9653,N_4287,N_3223);
or U9654 (N_9654,N_2427,N_3267);
nor U9655 (N_9655,N_4049,N_2857);
and U9656 (N_9656,N_3768,N_187);
and U9657 (N_9657,N_3333,N_1027);
or U9658 (N_9658,N_4291,N_2881);
nor U9659 (N_9659,N_4910,N_3064);
xor U9660 (N_9660,N_4008,N_3627);
xnor U9661 (N_9661,N_4297,N_3602);
and U9662 (N_9662,N_1065,N_312);
and U9663 (N_9663,N_3921,N_3038);
xnor U9664 (N_9664,N_4579,N_1188);
or U9665 (N_9665,N_274,N_773);
nand U9666 (N_9666,N_3100,N_1118);
nor U9667 (N_9667,N_3916,N_778);
or U9668 (N_9668,N_592,N_456);
and U9669 (N_9669,N_1160,N_3971);
and U9670 (N_9670,N_1578,N_793);
or U9671 (N_9671,N_1078,N_2814);
nor U9672 (N_9672,N_377,N_3828);
xnor U9673 (N_9673,N_3445,N_278);
nor U9674 (N_9674,N_3354,N_1154);
or U9675 (N_9675,N_3290,N_1096);
and U9676 (N_9676,N_3818,N_3437);
nor U9677 (N_9677,N_1658,N_2219);
nor U9678 (N_9678,N_328,N_2416);
or U9679 (N_9679,N_976,N_1931);
xnor U9680 (N_9680,N_4642,N_1681);
or U9681 (N_9681,N_1456,N_193);
xnor U9682 (N_9682,N_3990,N_928);
xor U9683 (N_9683,N_3697,N_3376);
or U9684 (N_9684,N_3918,N_635);
xor U9685 (N_9685,N_2597,N_147);
xor U9686 (N_9686,N_1402,N_3749);
or U9687 (N_9687,N_3330,N_3082);
or U9688 (N_9688,N_1122,N_3639);
nor U9689 (N_9689,N_4541,N_637);
and U9690 (N_9690,N_408,N_65);
or U9691 (N_9691,N_4238,N_2861);
nand U9692 (N_9692,N_725,N_3849);
xor U9693 (N_9693,N_3151,N_669);
nor U9694 (N_9694,N_4037,N_3794);
nor U9695 (N_9695,N_2865,N_2601);
xnor U9696 (N_9696,N_4116,N_89);
or U9697 (N_9697,N_1252,N_4950);
and U9698 (N_9698,N_4054,N_1367);
xor U9699 (N_9699,N_4850,N_2956);
and U9700 (N_9700,N_3687,N_2357);
and U9701 (N_9701,N_1231,N_2187);
xnor U9702 (N_9702,N_3960,N_3838);
nor U9703 (N_9703,N_1668,N_933);
nor U9704 (N_9704,N_4705,N_377);
xnor U9705 (N_9705,N_1256,N_1534);
nand U9706 (N_9706,N_2217,N_4525);
nor U9707 (N_9707,N_2253,N_3611);
nand U9708 (N_9708,N_1687,N_4027);
xnor U9709 (N_9709,N_42,N_2480);
nor U9710 (N_9710,N_274,N_1938);
or U9711 (N_9711,N_1028,N_2552);
nand U9712 (N_9712,N_2590,N_2386);
nand U9713 (N_9713,N_2167,N_4186);
nand U9714 (N_9714,N_3596,N_1667);
nor U9715 (N_9715,N_2327,N_2554);
or U9716 (N_9716,N_2719,N_1705);
and U9717 (N_9717,N_825,N_2541);
nor U9718 (N_9718,N_864,N_465);
nor U9719 (N_9719,N_4257,N_3598);
nor U9720 (N_9720,N_3570,N_1396);
nor U9721 (N_9721,N_1916,N_2829);
nand U9722 (N_9722,N_985,N_1339);
nor U9723 (N_9723,N_4678,N_2700);
and U9724 (N_9724,N_3076,N_1103);
nor U9725 (N_9725,N_3374,N_285);
nor U9726 (N_9726,N_2851,N_3934);
xnor U9727 (N_9727,N_983,N_4401);
nand U9728 (N_9728,N_315,N_1486);
nor U9729 (N_9729,N_502,N_4031);
xor U9730 (N_9730,N_206,N_4454);
and U9731 (N_9731,N_1112,N_664);
xor U9732 (N_9732,N_459,N_2509);
nor U9733 (N_9733,N_4467,N_2698);
nand U9734 (N_9734,N_3692,N_4872);
xnor U9735 (N_9735,N_289,N_1050);
nand U9736 (N_9736,N_4230,N_1554);
and U9737 (N_9737,N_1133,N_3152);
nor U9738 (N_9738,N_4637,N_216);
and U9739 (N_9739,N_4053,N_4793);
and U9740 (N_9740,N_1951,N_15);
and U9741 (N_9741,N_2395,N_611);
xnor U9742 (N_9742,N_80,N_4716);
and U9743 (N_9743,N_3328,N_3073);
nand U9744 (N_9744,N_3811,N_3546);
and U9745 (N_9745,N_273,N_74);
xor U9746 (N_9746,N_4835,N_2947);
xor U9747 (N_9747,N_4520,N_181);
nand U9748 (N_9748,N_2801,N_4438);
nor U9749 (N_9749,N_3704,N_1547);
and U9750 (N_9750,N_3281,N_4463);
nand U9751 (N_9751,N_3747,N_3648);
or U9752 (N_9752,N_3072,N_2818);
or U9753 (N_9753,N_2220,N_97);
xor U9754 (N_9754,N_3503,N_854);
xor U9755 (N_9755,N_1648,N_552);
and U9756 (N_9756,N_2225,N_1587);
and U9757 (N_9757,N_1592,N_4746);
and U9758 (N_9758,N_872,N_2318);
and U9759 (N_9759,N_3852,N_925);
and U9760 (N_9760,N_4978,N_2363);
nand U9761 (N_9761,N_525,N_3006);
and U9762 (N_9762,N_529,N_4935);
and U9763 (N_9763,N_4667,N_3115);
or U9764 (N_9764,N_3706,N_1164);
or U9765 (N_9765,N_4987,N_1180);
nor U9766 (N_9766,N_3261,N_2925);
and U9767 (N_9767,N_3105,N_2837);
xor U9768 (N_9768,N_1094,N_3375);
and U9769 (N_9769,N_42,N_2923);
nor U9770 (N_9770,N_4242,N_4023);
nand U9771 (N_9771,N_3342,N_313);
and U9772 (N_9772,N_2833,N_3124);
or U9773 (N_9773,N_4859,N_1652);
nand U9774 (N_9774,N_3385,N_4235);
xor U9775 (N_9775,N_2740,N_1274);
or U9776 (N_9776,N_4517,N_4519);
xor U9777 (N_9777,N_1906,N_4224);
nor U9778 (N_9778,N_4772,N_3670);
nand U9779 (N_9779,N_354,N_1001);
xor U9780 (N_9780,N_1251,N_3218);
or U9781 (N_9781,N_1669,N_4080);
xor U9782 (N_9782,N_4984,N_270);
xor U9783 (N_9783,N_736,N_4327);
nand U9784 (N_9784,N_4612,N_2578);
or U9785 (N_9785,N_558,N_1332);
nor U9786 (N_9786,N_3130,N_4065);
or U9787 (N_9787,N_1782,N_2805);
and U9788 (N_9788,N_4860,N_4663);
or U9789 (N_9789,N_3588,N_339);
and U9790 (N_9790,N_2919,N_1871);
or U9791 (N_9791,N_1823,N_4092);
nand U9792 (N_9792,N_3221,N_916);
nand U9793 (N_9793,N_2488,N_1884);
nor U9794 (N_9794,N_2030,N_812);
nand U9795 (N_9795,N_4153,N_4618);
and U9796 (N_9796,N_4526,N_4132);
and U9797 (N_9797,N_498,N_708);
xnor U9798 (N_9798,N_1548,N_2112);
and U9799 (N_9799,N_1597,N_4023);
xor U9800 (N_9800,N_4110,N_491);
and U9801 (N_9801,N_3656,N_2265);
nand U9802 (N_9802,N_1268,N_2627);
nand U9803 (N_9803,N_863,N_2345);
nor U9804 (N_9804,N_616,N_2596);
and U9805 (N_9805,N_4722,N_2314);
and U9806 (N_9806,N_2230,N_3796);
xor U9807 (N_9807,N_863,N_4896);
nand U9808 (N_9808,N_4703,N_1476);
nand U9809 (N_9809,N_2267,N_3544);
and U9810 (N_9810,N_3101,N_1245);
nand U9811 (N_9811,N_1127,N_1785);
or U9812 (N_9812,N_2742,N_105);
xor U9813 (N_9813,N_296,N_626);
nand U9814 (N_9814,N_537,N_2302);
xor U9815 (N_9815,N_3454,N_2179);
nand U9816 (N_9816,N_93,N_287);
and U9817 (N_9817,N_2865,N_3748);
or U9818 (N_9818,N_1197,N_2572);
and U9819 (N_9819,N_669,N_3434);
xor U9820 (N_9820,N_2175,N_2712);
nand U9821 (N_9821,N_4661,N_3308);
and U9822 (N_9822,N_2124,N_359);
or U9823 (N_9823,N_173,N_2471);
xor U9824 (N_9824,N_2609,N_1610);
and U9825 (N_9825,N_1173,N_4374);
or U9826 (N_9826,N_3862,N_918);
or U9827 (N_9827,N_3554,N_1534);
and U9828 (N_9828,N_923,N_500);
and U9829 (N_9829,N_1349,N_445);
and U9830 (N_9830,N_2789,N_2828);
and U9831 (N_9831,N_3539,N_3180);
xor U9832 (N_9832,N_522,N_825);
xnor U9833 (N_9833,N_2522,N_618);
xnor U9834 (N_9834,N_20,N_364);
nand U9835 (N_9835,N_826,N_4197);
nand U9836 (N_9836,N_3061,N_4683);
xor U9837 (N_9837,N_3859,N_4117);
nor U9838 (N_9838,N_4183,N_2618);
xor U9839 (N_9839,N_2057,N_4921);
or U9840 (N_9840,N_4754,N_1167);
and U9841 (N_9841,N_4531,N_1268);
or U9842 (N_9842,N_1308,N_2182);
xor U9843 (N_9843,N_1790,N_2566);
nor U9844 (N_9844,N_1936,N_609);
or U9845 (N_9845,N_3669,N_3730);
xor U9846 (N_9846,N_4606,N_1019);
xnor U9847 (N_9847,N_3636,N_3390);
nand U9848 (N_9848,N_2864,N_2691);
xor U9849 (N_9849,N_3074,N_451);
nand U9850 (N_9850,N_3187,N_376);
xor U9851 (N_9851,N_619,N_1650);
and U9852 (N_9852,N_802,N_3986);
xor U9853 (N_9853,N_2317,N_4454);
and U9854 (N_9854,N_3289,N_243);
xor U9855 (N_9855,N_3809,N_406);
and U9856 (N_9856,N_1568,N_4502);
nor U9857 (N_9857,N_4407,N_2585);
or U9858 (N_9858,N_1433,N_1507);
or U9859 (N_9859,N_4653,N_3050);
nand U9860 (N_9860,N_3185,N_3205);
nor U9861 (N_9861,N_944,N_579);
xnor U9862 (N_9862,N_581,N_3316);
xnor U9863 (N_9863,N_4146,N_4261);
nand U9864 (N_9864,N_1780,N_1937);
nor U9865 (N_9865,N_608,N_1884);
and U9866 (N_9866,N_3000,N_1221);
nand U9867 (N_9867,N_3062,N_4723);
or U9868 (N_9868,N_1624,N_941);
nor U9869 (N_9869,N_274,N_1557);
and U9870 (N_9870,N_1645,N_1442);
or U9871 (N_9871,N_4897,N_4642);
or U9872 (N_9872,N_278,N_4174);
or U9873 (N_9873,N_4795,N_900);
nor U9874 (N_9874,N_3525,N_2693);
or U9875 (N_9875,N_1264,N_362);
nor U9876 (N_9876,N_3426,N_4263);
and U9877 (N_9877,N_2430,N_3075);
or U9878 (N_9878,N_157,N_4644);
xnor U9879 (N_9879,N_3260,N_1215);
nand U9880 (N_9880,N_496,N_3737);
and U9881 (N_9881,N_2085,N_2888);
nand U9882 (N_9882,N_741,N_174);
xor U9883 (N_9883,N_2667,N_3824);
xnor U9884 (N_9884,N_2473,N_2575);
and U9885 (N_9885,N_361,N_2439);
and U9886 (N_9886,N_3010,N_3538);
nor U9887 (N_9887,N_422,N_1451);
xor U9888 (N_9888,N_4146,N_3723);
nor U9889 (N_9889,N_4977,N_1428);
and U9890 (N_9890,N_3940,N_3623);
xor U9891 (N_9891,N_1184,N_3743);
xor U9892 (N_9892,N_3571,N_1006);
nor U9893 (N_9893,N_3938,N_4165);
nand U9894 (N_9894,N_4649,N_2733);
or U9895 (N_9895,N_4793,N_3977);
nor U9896 (N_9896,N_4107,N_3197);
xnor U9897 (N_9897,N_1885,N_4960);
nand U9898 (N_9898,N_236,N_4523);
xnor U9899 (N_9899,N_4449,N_124);
or U9900 (N_9900,N_2863,N_2491);
nor U9901 (N_9901,N_2384,N_2013);
nand U9902 (N_9902,N_443,N_3747);
or U9903 (N_9903,N_579,N_76);
xnor U9904 (N_9904,N_2471,N_3666);
or U9905 (N_9905,N_342,N_456);
xnor U9906 (N_9906,N_764,N_2284);
nor U9907 (N_9907,N_1449,N_4641);
xnor U9908 (N_9908,N_2255,N_327);
nor U9909 (N_9909,N_2313,N_3851);
or U9910 (N_9910,N_4715,N_1366);
and U9911 (N_9911,N_1917,N_1905);
nor U9912 (N_9912,N_242,N_322);
and U9913 (N_9913,N_3971,N_4546);
nand U9914 (N_9914,N_4527,N_1762);
nor U9915 (N_9915,N_4184,N_828);
nor U9916 (N_9916,N_1725,N_2681);
nand U9917 (N_9917,N_3438,N_1707);
xor U9918 (N_9918,N_2195,N_641);
or U9919 (N_9919,N_341,N_3005);
nand U9920 (N_9920,N_1470,N_651);
xnor U9921 (N_9921,N_909,N_1641);
or U9922 (N_9922,N_186,N_2583);
xor U9923 (N_9923,N_4256,N_153);
and U9924 (N_9924,N_107,N_458);
nand U9925 (N_9925,N_1816,N_4858);
xnor U9926 (N_9926,N_2467,N_96);
nor U9927 (N_9927,N_3129,N_260);
xor U9928 (N_9928,N_2813,N_2886);
and U9929 (N_9929,N_3233,N_4191);
nor U9930 (N_9930,N_1616,N_3914);
xnor U9931 (N_9931,N_175,N_1220);
nor U9932 (N_9932,N_3273,N_2092);
or U9933 (N_9933,N_330,N_2284);
or U9934 (N_9934,N_1828,N_1785);
xor U9935 (N_9935,N_3887,N_1493);
nand U9936 (N_9936,N_3969,N_3945);
and U9937 (N_9937,N_3026,N_1434);
or U9938 (N_9938,N_3146,N_1261);
nor U9939 (N_9939,N_4732,N_677);
or U9940 (N_9940,N_4334,N_421);
nor U9941 (N_9941,N_2894,N_1754);
and U9942 (N_9942,N_4255,N_2804);
or U9943 (N_9943,N_570,N_950);
nor U9944 (N_9944,N_2187,N_3894);
and U9945 (N_9945,N_1126,N_2103);
or U9946 (N_9946,N_2385,N_4502);
nand U9947 (N_9947,N_4240,N_2043);
and U9948 (N_9948,N_1921,N_3140);
nor U9949 (N_9949,N_4321,N_2701);
nand U9950 (N_9950,N_1373,N_1128);
or U9951 (N_9951,N_1584,N_4805);
nor U9952 (N_9952,N_917,N_2580);
nand U9953 (N_9953,N_4237,N_2179);
nor U9954 (N_9954,N_4314,N_4714);
xor U9955 (N_9955,N_2923,N_1946);
xor U9956 (N_9956,N_3404,N_4629);
and U9957 (N_9957,N_4725,N_1678);
nor U9958 (N_9958,N_2007,N_3712);
or U9959 (N_9959,N_3006,N_316);
or U9960 (N_9960,N_269,N_1120);
or U9961 (N_9961,N_3997,N_1159);
nor U9962 (N_9962,N_69,N_4367);
or U9963 (N_9963,N_3511,N_2024);
and U9964 (N_9964,N_1019,N_2713);
xor U9965 (N_9965,N_4141,N_3091);
or U9966 (N_9966,N_2328,N_975);
nand U9967 (N_9967,N_2845,N_1218);
and U9968 (N_9968,N_625,N_1096);
xor U9969 (N_9969,N_2837,N_1777);
nor U9970 (N_9970,N_1822,N_2504);
and U9971 (N_9971,N_3701,N_4929);
xor U9972 (N_9972,N_4050,N_212);
nor U9973 (N_9973,N_3215,N_4793);
and U9974 (N_9974,N_4073,N_1154);
or U9975 (N_9975,N_2913,N_3448);
nor U9976 (N_9976,N_3434,N_4410);
nand U9977 (N_9977,N_1978,N_426);
nor U9978 (N_9978,N_1270,N_4991);
xor U9979 (N_9979,N_849,N_4301);
or U9980 (N_9980,N_4159,N_4836);
or U9981 (N_9981,N_2102,N_4930);
nor U9982 (N_9982,N_2791,N_2182);
nor U9983 (N_9983,N_3508,N_4600);
and U9984 (N_9984,N_4326,N_467);
xor U9985 (N_9985,N_1215,N_2455);
nor U9986 (N_9986,N_2984,N_1433);
nand U9987 (N_9987,N_570,N_4347);
nor U9988 (N_9988,N_1662,N_1896);
nor U9989 (N_9989,N_506,N_3636);
or U9990 (N_9990,N_3658,N_284);
xor U9991 (N_9991,N_542,N_2430);
nand U9992 (N_9992,N_3548,N_1198);
or U9993 (N_9993,N_2823,N_4833);
nor U9994 (N_9994,N_2863,N_4577);
xor U9995 (N_9995,N_4368,N_4287);
nor U9996 (N_9996,N_4735,N_260);
xor U9997 (N_9997,N_1289,N_2923);
and U9998 (N_9998,N_287,N_309);
nand U9999 (N_9999,N_278,N_2894);
nor U10000 (N_10000,N_6368,N_7053);
or U10001 (N_10001,N_5944,N_8418);
or U10002 (N_10002,N_7369,N_8898);
nand U10003 (N_10003,N_9035,N_5893);
nor U10004 (N_10004,N_8951,N_5630);
xor U10005 (N_10005,N_5053,N_8431);
and U10006 (N_10006,N_6935,N_8481);
nand U10007 (N_10007,N_5478,N_8754);
nor U10008 (N_10008,N_6380,N_8844);
and U10009 (N_10009,N_8366,N_8330);
nand U10010 (N_10010,N_6026,N_8142);
and U10011 (N_10011,N_9261,N_7980);
and U10012 (N_10012,N_9347,N_7561);
nor U10013 (N_10013,N_7652,N_8342);
and U10014 (N_10014,N_5289,N_5751);
nor U10015 (N_10015,N_6811,N_7696);
nor U10016 (N_10016,N_5559,N_9431);
xnor U10017 (N_10017,N_8714,N_7386);
xnor U10018 (N_10018,N_5915,N_8201);
and U10019 (N_10019,N_8253,N_6256);
and U10020 (N_10020,N_9492,N_5250);
xnor U10021 (N_10021,N_6599,N_5083);
nor U10022 (N_10022,N_7345,N_6622);
nor U10023 (N_10023,N_5805,N_8640);
nand U10024 (N_10024,N_9168,N_9128);
xnor U10025 (N_10025,N_6769,N_5838);
or U10026 (N_10026,N_6985,N_9468);
and U10027 (N_10027,N_8089,N_5293);
or U10028 (N_10028,N_8775,N_8685);
xnor U10029 (N_10029,N_6150,N_5528);
and U10030 (N_10030,N_5829,N_7663);
nor U10031 (N_10031,N_6139,N_5457);
nor U10032 (N_10032,N_6080,N_7156);
nand U10033 (N_10033,N_8622,N_5632);
and U10034 (N_10034,N_7293,N_7276);
xnor U10035 (N_10035,N_7115,N_5583);
or U10036 (N_10036,N_6321,N_7752);
and U10037 (N_10037,N_9250,N_7299);
nor U10038 (N_10038,N_8061,N_7568);
and U10039 (N_10039,N_9724,N_7389);
and U10040 (N_10040,N_6420,N_7153);
xnor U10041 (N_10041,N_6748,N_5955);
and U10042 (N_10042,N_6651,N_7617);
or U10043 (N_10043,N_7729,N_9239);
nor U10044 (N_10044,N_9576,N_7608);
and U10045 (N_10045,N_8294,N_7998);
nand U10046 (N_10046,N_5309,N_7140);
xnor U10047 (N_10047,N_9318,N_7587);
and U10048 (N_10048,N_6400,N_9842);
xnor U10049 (N_10049,N_9582,N_8426);
or U10050 (N_10050,N_7230,N_6886);
or U10051 (N_10051,N_5948,N_5570);
nor U10052 (N_10052,N_8083,N_8214);
or U10053 (N_10053,N_8948,N_7219);
nor U10054 (N_10054,N_7987,N_8126);
and U10055 (N_10055,N_5049,N_8269);
nor U10056 (N_10056,N_7047,N_7307);
or U10057 (N_10057,N_7779,N_5160);
or U10058 (N_10058,N_8022,N_5611);
and U10059 (N_10059,N_9398,N_5364);
xnor U10060 (N_10060,N_8739,N_5777);
xnor U10061 (N_10061,N_7934,N_7968);
or U10062 (N_10062,N_7192,N_8581);
xor U10063 (N_10063,N_8930,N_5377);
nor U10064 (N_10064,N_7322,N_6175);
or U10065 (N_10065,N_6565,N_9254);
nand U10066 (N_10066,N_8892,N_9830);
and U10067 (N_10067,N_6242,N_6874);
xor U10068 (N_10068,N_8288,N_7812);
nor U10069 (N_10069,N_9943,N_7986);
or U10070 (N_10070,N_5897,N_8616);
xor U10071 (N_10071,N_6033,N_7187);
or U10072 (N_10072,N_8403,N_5140);
and U10073 (N_10073,N_9530,N_6958);
xor U10074 (N_10074,N_6771,N_6646);
xnor U10075 (N_10075,N_6952,N_8282);
nand U10076 (N_10076,N_6604,N_9288);
nand U10077 (N_10077,N_9799,N_8815);
nand U10078 (N_10078,N_6530,N_6743);
nand U10079 (N_10079,N_5175,N_9833);
and U10080 (N_10080,N_7073,N_7501);
nand U10081 (N_10081,N_8575,N_6361);
nand U10082 (N_10082,N_6853,N_8514);
or U10083 (N_10083,N_8504,N_5545);
and U10084 (N_10084,N_6701,N_7390);
and U10085 (N_10085,N_8752,N_9859);
and U10086 (N_10086,N_6427,N_8274);
or U10087 (N_10087,N_6404,N_5512);
nor U10088 (N_10088,N_9803,N_7081);
nand U10089 (N_10089,N_9666,N_5030);
or U10090 (N_10090,N_7712,N_8865);
and U10091 (N_10091,N_6645,N_5892);
nand U10092 (N_10092,N_7489,N_7315);
nor U10093 (N_10093,N_6971,N_5685);
nand U10094 (N_10094,N_6839,N_6178);
nand U10095 (N_10095,N_8726,N_6895);
or U10096 (N_10096,N_5676,N_7347);
nor U10097 (N_10097,N_6705,N_8814);
nor U10098 (N_10098,N_8800,N_7433);
nor U10099 (N_10099,N_6310,N_9969);
and U10100 (N_10100,N_7738,N_9702);
or U10101 (N_10101,N_6975,N_8797);
xor U10102 (N_10102,N_7923,N_5452);
or U10103 (N_10103,N_8636,N_7872);
nor U10104 (N_10104,N_8002,N_7973);
or U10105 (N_10105,N_7864,N_7842);
or U10106 (N_10106,N_6413,N_6672);
and U10107 (N_10107,N_5764,N_7348);
or U10108 (N_10108,N_8590,N_8679);
nor U10109 (N_10109,N_8630,N_9181);
nand U10110 (N_10110,N_6990,N_9466);
or U10111 (N_10111,N_9813,N_5850);
nand U10112 (N_10112,N_6838,N_8073);
or U10113 (N_10113,N_9759,N_5940);
nor U10114 (N_10114,N_7335,N_9024);
nand U10115 (N_10115,N_5108,N_5661);
nor U10116 (N_10116,N_8978,N_5907);
xor U10117 (N_10117,N_9015,N_7990);
or U10118 (N_10118,N_8146,N_9953);
and U10119 (N_10119,N_6348,N_6173);
xor U10120 (N_10120,N_6715,N_6077);
xnor U10121 (N_10121,N_6472,N_7191);
xnor U10122 (N_10122,N_8378,N_6916);
or U10123 (N_10123,N_5969,N_8984);
and U10124 (N_10124,N_5332,N_8200);
and U10125 (N_10125,N_9867,N_6823);
xnor U10126 (N_10126,N_8725,N_8990);
xor U10127 (N_10127,N_7952,N_7581);
nor U10128 (N_10128,N_5703,N_9452);
nor U10129 (N_10129,N_5608,N_6152);
and U10130 (N_10130,N_5280,N_5429);
xnor U10131 (N_10131,N_5151,N_5172);
and U10132 (N_10132,N_8343,N_8728);
xor U10133 (N_10133,N_6351,N_6213);
and U10134 (N_10134,N_7025,N_7228);
nor U10135 (N_10135,N_6738,N_6064);
and U10136 (N_10136,N_9743,N_8758);
xnor U10137 (N_10137,N_5016,N_5726);
nand U10138 (N_10138,N_7248,N_8000);
or U10139 (N_10139,N_5264,N_9723);
and U10140 (N_10140,N_8913,N_5261);
nor U10141 (N_10141,N_7136,N_8199);
and U10142 (N_10142,N_6439,N_8033);
nor U10143 (N_10143,N_8092,N_8664);
nand U10144 (N_10144,N_6263,N_6741);
or U10145 (N_10145,N_8009,N_6510);
nor U10146 (N_10146,N_6628,N_7280);
xor U10147 (N_10147,N_5900,N_9375);
nor U10148 (N_10148,N_7242,N_5563);
xnor U10149 (N_10149,N_8341,N_5345);
xnor U10150 (N_10150,N_9774,N_6953);
xnor U10151 (N_10151,N_9648,N_8662);
and U10152 (N_10152,N_7457,N_7849);
or U10153 (N_10153,N_9159,N_7567);
and U10154 (N_10154,N_8539,N_9081);
xor U10155 (N_10155,N_9342,N_7540);
xor U10156 (N_10156,N_9777,N_5371);
nor U10157 (N_10157,N_6896,N_6986);
xnor U10158 (N_10158,N_8748,N_8170);
nand U10159 (N_10159,N_5860,N_5472);
nand U10160 (N_10160,N_7971,N_5189);
nand U10161 (N_10161,N_7521,N_8076);
xnor U10162 (N_10162,N_7071,N_8138);
and U10163 (N_10163,N_7625,N_6485);
nor U10164 (N_10164,N_5741,N_6337);
or U10165 (N_10165,N_8498,N_8610);
nand U10166 (N_10166,N_5849,N_7977);
or U10167 (N_10167,N_9694,N_6180);
and U10168 (N_10168,N_6004,N_8899);
nand U10169 (N_10169,N_9495,N_5448);
nor U10170 (N_10170,N_5959,N_7377);
xor U10171 (N_10171,N_6970,N_9118);
nand U10172 (N_10172,N_8606,N_6829);
xnor U10173 (N_10173,N_8323,N_9682);
xor U10174 (N_10174,N_9605,N_9764);
nor U10175 (N_10175,N_9031,N_9243);
or U10176 (N_10176,N_7718,N_6461);
or U10177 (N_10177,N_6431,N_9965);
or U10178 (N_10178,N_5841,N_6317);
and U10179 (N_10179,N_8392,N_8968);
nand U10180 (N_10180,N_8793,N_8524);
or U10181 (N_10181,N_9802,N_9152);
nand U10182 (N_10182,N_9198,N_6383);
xnor U10183 (N_10183,N_6398,N_9073);
nand U10184 (N_10184,N_7095,N_5586);
and U10185 (N_10185,N_6155,N_7157);
xor U10186 (N_10186,N_6529,N_7430);
and U10187 (N_10187,N_9194,N_6775);
or U10188 (N_10188,N_6473,N_5567);
or U10189 (N_10189,N_7227,N_6136);
and U10190 (N_10190,N_6949,N_7897);
or U10191 (N_10191,N_9588,N_8600);
or U10192 (N_10192,N_6765,N_8154);
xnor U10193 (N_10193,N_8300,N_6883);
nor U10194 (N_10194,N_8568,N_6808);
xnor U10195 (N_10195,N_7520,N_6452);
and U10196 (N_10196,N_6225,N_9310);
nand U10197 (N_10197,N_6888,N_5961);
nand U10198 (N_10198,N_8667,N_5787);
and U10199 (N_10199,N_8565,N_8335);
xnor U10200 (N_10200,N_7126,N_9471);
xnor U10201 (N_10201,N_5395,N_8346);
or U10202 (N_10202,N_7488,N_7124);
nand U10203 (N_10203,N_8583,N_7671);
nand U10204 (N_10204,N_9522,N_5380);
nand U10205 (N_10205,N_8164,N_8046);
xor U10206 (N_10206,N_6846,N_6137);
and U10207 (N_10207,N_8897,N_9339);
and U10208 (N_10208,N_7077,N_6641);
nand U10209 (N_10209,N_5322,N_7648);
nor U10210 (N_10210,N_8976,N_5645);
xnor U10211 (N_10211,N_5483,N_9078);
nor U10212 (N_10212,N_5895,N_8571);
or U10213 (N_10213,N_6119,N_9560);
nor U10214 (N_10214,N_9658,N_5998);
nand U10215 (N_10215,N_8005,N_9422);
and U10216 (N_10216,N_5921,N_8143);
xor U10217 (N_10217,N_7471,N_9382);
or U10218 (N_10218,N_5052,N_7411);
and U10219 (N_10219,N_7757,N_9340);
and U10220 (N_10220,N_7667,N_7428);
or U10221 (N_10221,N_6484,N_8249);
xnor U10222 (N_10222,N_8988,N_5889);
xor U10223 (N_10223,N_7321,N_8543);
nand U10224 (N_10224,N_9356,N_7640);
nand U10225 (N_10225,N_8587,N_6603);
nor U10226 (N_10226,N_6643,N_9516);
or U10227 (N_10227,N_8557,N_6760);
nand U10228 (N_10228,N_6509,N_8133);
or U10229 (N_10229,N_9945,N_6303);
nand U10230 (N_10230,N_9806,N_7290);
xor U10231 (N_10231,N_7852,N_6982);
xor U10232 (N_10232,N_9855,N_9504);
xor U10233 (N_10233,N_7491,N_7658);
and U10234 (N_10234,N_5800,N_9814);
xor U10235 (N_10235,N_5300,N_6757);
nor U10236 (N_10236,N_5328,N_8961);
xnor U10237 (N_10237,N_9484,N_6746);
or U10238 (N_10238,N_6742,N_7068);
and U10239 (N_10239,N_7982,N_8649);
or U10240 (N_10240,N_9371,N_9532);
nand U10241 (N_10241,N_5865,N_5418);
nand U10242 (N_10242,N_7744,N_6496);
and U10243 (N_10243,N_5982,N_9866);
and U10244 (N_10244,N_6328,N_5144);
and U10245 (N_10245,N_5859,N_6695);
nand U10246 (N_10246,N_8210,N_9000);
xor U10247 (N_10247,N_9981,N_5212);
and U10248 (N_10248,N_7624,N_8205);
and U10249 (N_10249,N_9205,N_5562);
nand U10250 (N_10250,N_5158,N_6053);
or U10251 (N_10251,N_9987,N_9817);
xnor U10252 (N_10252,N_5027,N_6712);
or U10253 (N_10253,N_7423,N_8674);
xnor U10254 (N_10254,N_6716,N_8078);
nor U10255 (N_10255,N_6910,N_6056);
nor U10256 (N_10256,N_7586,N_9140);
nor U10257 (N_10257,N_7706,N_6983);
and U10258 (N_10258,N_7122,N_9584);
and U10259 (N_10259,N_8047,N_9919);
xor U10260 (N_10260,N_5600,N_7443);
or U10261 (N_10261,N_9272,N_8542);
nand U10262 (N_10262,N_9660,N_9569);
and U10263 (N_10263,N_8451,N_7856);
or U10264 (N_10264,N_5621,N_6795);
nor U10265 (N_10265,N_6831,N_9019);
and U10266 (N_10266,N_7459,N_6331);
or U10267 (N_10267,N_8429,N_9514);
xnor U10268 (N_10268,N_9600,N_5489);
and U10269 (N_10269,N_6890,N_6389);
xnor U10270 (N_10270,N_9596,N_5155);
and U10271 (N_10271,N_5626,N_7478);
nand U10272 (N_10272,N_9420,N_5691);
or U10273 (N_10273,N_6459,N_7629);
nand U10274 (N_10274,N_5042,N_5846);
or U10275 (N_10275,N_7109,N_9931);
xor U10276 (N_10276,N_7479,N_6306);
and U10277 (N_10277,N_8453,N_7070);
xnor U10278 (N_10278,N_6316,N_6777);
and U10279 (N_10279,N_6249,N_6430);
nand U10280 (N_10280,N_8842,N_9312);
and U10281 (N_10281,N_7450,N_7911);
xor U10282 (N_10282,N_7426,N_5762);
or U10283 (N_10283,N_8114,N_6934);
xnor U10284 (N_10284,N_5960,N_7253);
nor U10285 (N_10285,N_5941,N_5625);
or U10286 (N_10286,N_8601,N_8877);
nand U10287 (N_10287,N_6450,N_6796);
or U10288 (N_10288,N_7089,N_9552);
nor U10289 (N_10289,N_8982,N_7670);
xor U10290 (N_10290,N_5283,N_6907);
nand U10291 (N_10291,N_9918,N_5973);
or U10292 (N_10292,N_7027,N_6514);
and U10293 (N_10293,N_9556,N_8457);
nor U10294 (N_10294,N_5758,N_6592);
and U10295 (N_10295,N_7533,N_9069);
and U10296 (N_10296,N_5033,N_9824);
nand U10297 (N_10297,N_6616,N_8012);
xnor U10298 (N_10298,N_9700,N_8159);
nand U10299 (N_10299,N_5702,N_9841);
nand U10300 (N_10300,N_5252,N_7727);
or U10301 (N_10301,N_5084,N_7367);
nor U10302 (N_10302,N_5389,N_5336);
or U10303 (N_10303,N_8925,N_7167);
xnor U10304 (N_10304,N_6951,N_5825);
or U10305 (N_10305,N_8954,N_7364);
nand U10306 (N_10306,N_8141,N_7151);
xnor U10307 (N_10307,N_6267,N_8358);
xor U10308 (N_10308,N_6942,N_7094);
nand U10309 (N_10309,N_9735,N_9745);
or U10310 (N_10310,N_7113,N_5430);
nor U10311 (N_10311,N_8079,N_7205);
nor U10312 (N_10312,N_7879,N_8582);
and U10313 (N_10313,N_9022,N_5906);
and U10314 (N_10314,N_7957,N_5304);
xor U10315 (N_10315,N_9319,N_9904);
xnor U10316 (N_10316,N_8801,N_9107);
or U10317 (N_10317,N_5174,N_6878);
or U10318 (N_10318,N_6029,N_5811);
xor U10319 (N_10319,N_9646,N_7063);
xnor U10320 (N_10320,N_5864,N_6593);
or U10321 (N_10321,N_5058,N_7044);
nor U10322 (N_10322,N_6079,N_6656);
nor U10323 (N_10323,N_9898,N_6601);
nand U10324 (N_10324,N_8299,N_7370);
xor U10325 (N_10325,N_7300,N_5715);
nor U10326 (N_10326,N_7901,N_6370);
nor U10327 (N_10327,N_5254,N_5481);
xnor U10328 (N_10328,N_5997,N_8305);
nor U10329 (N_10329,N_7910,N_5890);
nand U10330 (N_10330,N_5383,N_6614);
and U10331 (N_10331,N_7424,N_6402);
and U10332 (N_10332,N_7352,N_6873);
nor U10333 (N_10333,N_5623,N_5116);
nand U10334 (N_10334,N_6073,N_9929);
and U10335 (N_10335,N_5749,N_9358);
or U10336 (N_10336,N_6806,N_6919);
or U10337 (N_10337,N_5885,N_6184);
xor U10338 (N_10338,N_9301,N_6470);
nand U10339 (N_10339,N_8672,N_8869);
nor U10340 (N_10340,N_6955,N_9470);
nand U10341 (N_10341,N_9831,N_9839);
and U10342 (N_10342,N_8713,N_7780);
nand U10343 (N_10343,N_7455,N_5072);
or U10344 (N_10344,N_9850,N_8338);
nand U10345 (N_10345,N_8522,N_6412);
xor U10346 (N_10346,N_9649,N_5592);
nand U10347 (N_10347,N_5015,N_6411);
and U10348 (N_10348,N_5008,N_5240);
nand U10349 (N_10349,N_9101,N_8056);
nand U10350 (N_10350,N_9882,N_5334);
or U10351 (N_10351,N_5359,N_7824);
xnor U10352 (N_10352,N_6954,N_7496);
and U10353 (N_10353,N_5017,N_5561);
xnor U10354 (N_10354,N_5228,N_6167);
and U10355 (N_10355,N_8123,N_5813);
nand U10356 (N_10356,N_9754,N_7395);
nand U10357 (N_10357,N_6763,N_8071);
nand U10358 (N_10358,N_9726,N_7504);
or U10359 (N_10359,N_6138,N_5496);
nor U10360 (N_10360,N_5077,N_6444);
and U10361 (N_10361,N_7653,N_6342);
nand U10362 (N_10362,N_7019,N_5205);
xnor U10363 (N_10363,N_7865,N_8651);
xor U10364 (N_10364,N_5752,N_9796);
and U10365 (N_10365,N_5678,N_9717);
nor U10366 (N_10366,N_6857,N_5223);
nand U10367 (N_10367,N_7638,N_8278);
and U10368 (N_10368,N_7907,N_9186);
xor U10369 (N_10369,N_6244,N_7030);
or U10370 (N_10370,N_7823,N_6751);
or U10371 (N_10371,N_9645,N_8715);
or U10372 (N_10372,N_5112,N_9713);
nand U10373 (N_10373,N_7554,N_5954);
or U10374 (N_10374,N_8761,N_8776);
and U10375 (N_10375,N_5115,N_8067);
nor U10376 (N_10376,N_9008,N_7464);
nand U10377 (N_10377,N_9822,N_5458);
nor U10378 (N_10378,N_5689,N_6471);
or U10379 (N_10379,N_7605,N_7143);
or U10380 (N_10380,N_9062,N_8952);
or U10381 (N_10381,N_6280,N_6639);
and U10382 (N_10382,N_6231,N_8433);
or U10383 (N_10383,N_9704,N_5615);
or U10384 (N_10384,N_8292,N_8983);
nor U10385 (N_10385,N_5089,N_7241);
or U10386 (N_10386,N_7273,N_8873);
or U10387 (N_10387,N_8093,N_6451);
nor U10388 (N_10388,N_8438,N_9265);
and U10389 (N_10389,N_7310,N_6581);
nor U10390 (N_10390,N_7735,N_6627);
xnor U10391 (N_10391,N_8189,N_8290);
and U10392 (N_10392,N_6237,N_5196);
xnor U10393 (N_10393,N_7378,N_8859);
and U10394 (N_10394,N_6127,N_5552);
xor U10395 (N_10395,N_9247,N_5476);
nor U10396 (N_10396,N_9651,N_7564);
and U10397 (N_10397,N_6475,N_8966);
and U10398 (N_10398,N_9574,N_7822);
nor U10399 (N_10399,N_8935,N_5603);
nand U10400 (N_10400,N_7085,N_5684);
or U10401 (N_10401,N_7356,N_6418);
nor U10402 (N_10402,N_8243,N_5657);
and U10403 (N_10403,N_8519,N_7788);
xor U10404 (N_10404,N_7532,N_5425);
or U10405 (N_10405,N_8777,N_7976);
xnor U10406 (N_10406,N_5248,N_8862);
nor U10407 (N_10407,N_5513,N_6074);
nor U10408 (N_10408,N_5078,N_8206);
nor U10409 (N_10409,N_9126,N_9013);
xnor U10410 (N_10410,N_9900,N_8687);
xnor U10411 (N_10411,N_7127,N_8548);
nand U10412 (N_10412,N_7412,N_9449);
or U10413 (N_10413,N_5556,N_7509);
nand U10414 (N_10414,N_8272,N_9609);
nand U10415 (N_10415,N_8906,N_7326);
nand U10416 (N_10416,N_9770,N_7200);
nor U10417 (N_10417,N_5307,N_6379);
or U10418 (N_10418,N_8363,N_5868);
nor U10419 (N_10419,N_7673,N_7777);
xnor U10420 (N_10420,N_6520,N_9188);
and U10421 (N_10421,N_6135,N_8497);
or U10422 (N_10422,N_9147,N_5402);
and U10423 (N_10423,N_9592,N_9630);
or U10424 (N_10424,N_7921,N_6677);
nor U10425 (N_10425,N_8441,N_6273);
nand U10426 (N_10426,N_6435,N_5674);
and U10427 (N_10427,N_7301,N_9045);
xnor U10428 (N_10428,N_7270,N_9323);
nor U10429 (N_10429,N_8150,N_8385);
and U10430 (N_10430,N_8684,N_6070);
and U10431 (N_10431,N_5319,N_5443);
xnor U10432 (N_10432,N_8436,N_9042);
or U10433 (N_10433,N_5866,N_7419);
xnor U10434 (N_10434,N_5574,N_7731);
or U10435 (N_10435,N_7139,N_9763);
nor U10436 (N_10436,N_8722,N_7551);
or U10437 (N_10437,N_8439,N_8698);
xor U10438 (N_10438,N_8821,N_6694);
or U10439 (N_10439,N_8317,N_7274);
and U10440 (N_10440,N_9037,N_6059);
xnor U10441 (N_10441,N_8069,N_8301);
and U10442 (N_10442,N_9878,N_5453);
or U10443 (N_10443,N_5344,N_8521);
or U10444 (N_10444,N_8847,N_5211);
xor U10445 (N_10445,N_8627,N_8449);
xor U10446 (N_10446,N_9054,N_8465);
nor U10447 (N_10447,N_9150,N_8202);
nor U10448 (N_10448,N_7938,N_8798);
or U10449 (N_10449,N_9417,N_6327);
nor U10450 (N_10450,N_6579,N_5742);
nor U10451 (N_10451,N_9948,N_9886);
and U10452 (N_10452,N_6010,N_8298);
or U10453 (N_10453,N_6114,N_5816);
xor U10454 (N_10454,N_7541,N_8320);
nand U10455 (N_10455,N_6159,N_7059);
or U10456 (N_10456,N_7913,N_5810);
xor U10457 (N_10457,N_9875,N_9368);
and U10458 (N_10458,N_8615,N_9184);
nand U10459 (N_10459,N_5981,N_5855);
xnor U10460 (N_10460,N_6595,N_8556);
and U10461 (N_10461,N_5209,N_7058);
or U10462 (N_10462,N_6493,N_5711);
and U10463 (N_10463,N_5492,N_6642);
xnor U10464 (N_10464,N_6735,N_9354);
and U10465 (N_10465,N_7407,N_5706);
nor U10466 (N_10466,N_6375,N_6414);
xor U10467 (N_10467,N_7915,N_5297);
or U10468 (N_10468,N_6703,N_9884);
or U10469 (N_10469,N_6403,N_5125);
nand U10470 (N_10470,N_9937,N_5584);
nand U10471 (N_10471,N_5793,N_5786);
and U10472 (N_10472,N_9388,N_6863);
xor U10473 (N_10473,N_6609,N_7552);
nand U10474 (N_10474,N_8607,N_7163);
xnor U10475 (N_10475,N_7708,N_7868);
xnor U10476 (N_10476,N_7018,N_8805);
and U10477 (N_10477,N_7700,N_6504);
and U10478 (N_10478,N_8510,N_6464);
nor U10479 (N_10479,N_7458,N_9742);
xor U10480 (N_10480,N_9396,N_9137);
and U10481 (N_10481,N_6502,N_8934);
or U10482 (N_10482,N_9027,N_9359);
nor U10483 (N_10483,N_6723,N_6453);
and U10484 (N_10484,N_8267,N_6872);
nand U10485 (N_10485,N_5235,N_9049);
nand U10486 (N_10486,N_5324,N_8738);
nand U10487 (N_10487,N_6876,N_5317);
or U10488 (N_10488,N_6683,N_8773);
nand U10489 (N_10489,N_8508,N_6113);
xnor U10490 (N_10490,N_7981,N_7674);
xor U10491 (N_10491,N_5641,N_7972);
xnor U10492 (N_10492,N_7715,N_5234);
nor U10493 (N_10493,N_5449,N_8941);
nor U10494 (N_10494,N_8487,N_8972);
or U10495 (N_10495,N_8186,N_8023);
nand U10496 (N_10496,N_5149,N_8746);
xor U10497 (N_10497,N_5409,N_9804);
nor U10498 (N_10498,N_9048,N_6497);
nor U10499 (N_10499,N_5862,N_8262);
and U10500 (N_10500,N_8377,N_9285);
xor U10501 (N_10501,N_5066,N_9047);
or U10502 (N_10502,N_8178,N_9860);
and U10503 (N_10503,N_8291,N_8768);
or U10504 (N_10504,N_8513,N_8007);
nor U10505 (N_10505,N_9920,N_6667);
nor U10506 (N_10506,N_9153,N_7515);
nand U10507 (N_10507,N_8165,N_9350);
and U10508 (N_10508,N_5514,N_9377);
and U10509 (N_10509,N_5358,N_8788);
or U10510 (N_10510,N_9084,N_8387);
or U10511 (N_10511,N_6662,N_7946);
nor U10512 (N_10512,N_8724,N_7877);
nor U10513 (N_10513,N_6882,N_6826);
xor U10514 (N_10514,N_8732,N_7832);
xor U10515 (N_10515,N_5074,N_8415);
or U10516 (N_10516,N_9345,N_9999);
nor U10517 (N_10517,N_8618,N_8389);
nor U10518 (N_10518,N_7284,N_6034);
or U10519 (N_10519,N_5485,N_5101);
nand U10520 (N_10520,N_6511,N_8979);
or U10521 (N_10521,N_5236,N_7396);
nor U10522 (N_10522,N_9427,N_8645);
or U10523 (N_10523,N_5904,N_5634);
nand U10524 (N_10524,N_7676,N_6663);
nor U10525 (N_10525,N_5748,N_8997);
nand U10526 (N_10526,N_8855,N_7125);
nand U10527 (N_10527,N_7792,N_8386);
nand U10528 (N_10528,N_9676,N_6240);
and U10529 (N_10529,N_7556,N_5423);
xnor U10530 (N_10530,N_7039,N_7258);
nor U10531 (N_10531,N_9281,N_6550);
and U10532 (N_10532,N_7578,N_9440);
nand U10533 (N_10533,N_8512,N_9141);
or U10534 (N_10534,N_7988,N_8489);
and U10535 (N_10535,N_7862,N_8675);
xor U10536 (N_10536,N_6512,N_8276);
or U10537 (N_10537,N_5836,N_9023);
xnor U10538 (N_10538,N_5853,N_8106);
and U10539 (N_10539,N_5949,N_8774);
nand U10540 (N_10540,N_6043,N_6937);
nand U10541 (N_10541,N_7265,N_9736);
and U10542 (N_10542,N_9650,N_9852);
or U10543 (N_10543,N_5043,N_5919);
or U10544 (N_10544,N_8336,N_6088);
nor U10545 (N_10545,N_9680,N_6416);
or U10546 (N_10546,N_8944,N_8766);
xnor U10547 (N_10547,N_9381,N_6582);
nand U10548 (N_10548,N_7557,N_8235);
nand U10549 (N_10549,N_8486,N_8177);
nand U10550 (N_10550,N_8090,N_7239);
or U10551 (N_10551,N_9551,N_7719);
nand U10552 (N_10552,N_8750,N_9565);
xor U10553 (N_10553,N_5660,N_5507);
xnor U10554 (N_10554,N_7753,N_8809);
xor U10555 (N_10555,N_6332,N_7002);
and U10556 (N_10556,N_8359,N_8779);
or U10557 (N_10557,N_8638,N_8911);
or U10558 (N_10558,N_9208,N_6397);
and U10559 (N_10559,N_7771,N_5502);
and U10560 (N_10560,N_8986,N_7184);
and U10561 (N_10561,N_8730,N_5061);
or U10562 (N_10562,N_8765,N_6668);
nor U10563 (N_10563,N_9762,N_6458);
nand U10564 (N_10564,N_7180,N_7524);
xor U10565 (N_10565,N_5311,N_5644);
and U10566 (N_10566,N_7894,N_8103);
nand U10567 (N_10567,N_8501,N_9076);
xor U10568 (N_10568,N_8500,N_5876);
and U10569 (N_10569,N_7790,N_5858);
and U10570 (N_10570,N_6078,N_8476);
and U10571 (N_10571,N_5387,N_8420);
nor U10572 (N_10572,N_8255,N_5617);
and U10573 (N_10573,N_6946,N_8880);
nor U10574 (N_10574,N_5398,N_5698);
nor U10575 (N_10575,N_5456,N_7092);
xor U10576 (N_10576,N_8810,N_5986);
and U10577 (N_10577,N_6259,N_7672);
or U10578 (N_10578,N_8101,N_9089);
xor U10579 (N_10579,N_6586,N_5601);
nor U10580 (N_10580,N_9325,N_5459);
and U10581 (N_10581,N_9262,N_9441);
or U10582 (N_10582,N_9095,N_5355);
and U10583 (N_10583,N_6232,N_9088);
xor U10584 (N_10584,N_8216,N_8566);
nand U10585 (N_10585,N_7511,N_6535);
or U10586 (N_10586,N_5822,N_7074);
nand U10587 (N_10587,N_8503,N_5754);
nand U10588 (N_10588,N_9276,N_5118);
or U10589 (N_10589,N_8435,N_9012);
xor U10590 (N_10590,N_9498,N_6038);
nand U10591 (N_10591,N_9056,N_8163);
nor U10592 (N_10592,N_6013,N_8643);
or U10593 (N_10593,N_5312,N_8130);
nand U10594 (N_10594,N_6417,N_5251);
and U10595 (N_10595,N_5046,N_7147);
nand U10596 (N_10596,N_5721,N_9219);
and U10597 (N_10597,N_8807,N_6922);
nor U10598 (N_10598,N_8271,N_9825);
nor U10599 (N_10599,N_6169,N_9138);
and U10600 (N_10600,N_9755,N_9765);
xnor U10601 (N_10601,N_7029,N_6532);
and U10602 (N_10602,N_8382,N_6679);
xor U10603 (N_10603,N_8703,N_7316);
nor U10604 (N_10604,N_6278,N_5385);
nor U10605 (N_10605,N_7732,N_7414);
xnor U10606 (N_10606,N_9952,N_7490);
nand U10607 (N_10607,N_5651,N_7108);
or U10608 (N_10608,N_8463,N_9300);
nor U10609 (N_10609,N_7784,N_8111);
nor U10610 (N_10610,N_8063,N_5832);
xnor U10611 (N_10611,N_7079,N_6562);
nor U10612 (N_10612,N_9989,N_7272);
and U10613 (N_10613,N_8794,N_9286);
xnor U10614 (N_10614,N_5226,N_7703);
xor U10615 (N_10615,N_9496,N_6596);
and U10616 (N_10616,N_7656,N_7655);
and U10617 (N_10617,N_9235,N_9572);
or U10618 (N_10618,N_9477,N_7801);
nand U10619 (N_10619,N_5446,N_5525);
nor U10620 (N_10620,N_7876,N_5145);
nor U10621 (N_10621,N_7161,N_7886);
xnor U10622 (N_10622,N_8390,N_6323);
xnor U10623 (N_10623,N_6966,N_8918);
and U10624 (N_10624,N_9714,N_9248);
nand U10625 (N_10625,N_9415,N_7435);
xnor U10626 (N_10626,N_5770,N_8927);
or U10627 (N_10627,N_9175,N_8525);
nor U10628 (N_10628,N_5794,N_6415);
or U10629 (N_10629,N_6577,N_5321);
and U10630 (N_10630,N_8350,N_7807);
nor U10631 (N_10631,N_6770,N_7434);
xor U10632 (N_10632,N_6217,N_7220);
and U10633 (N_10633,N_9647,N_6296);
nor U10634 (N_10634,N_6442,N_8888);
and U10635 (N_10635,N_6012,N_9407);
xnor U10636 (N_10636,N_7250,N_8057);
and U10637 (N_10637,N_7994,N_7380);
or U10638 (N_10638,N_7799,N_7006);
nor U10639 (N_10639,N_8180,N_9591);
and U10640 (N_10640,N_7863,N_6154);
xor U10641 (N_10641,N_9378,N_7831);
or U10642 (N_10642,N_5739,N_9299);
and U10643 (N_10643,N_7231,N_5680);
and U10644 (N_10644,N_6048,N_5025);
or U10645 (N_10645,N_9478,N_6871);
and U10646 (N_10646,N_6931,N_9633);
and U10647 (N_10647,N_9750,N_6906);
nor U10648 (N_10648,N_9136,N_8024);
nor U10649 (N_10649,N_9979,N_5511);
or U10650 (N_10650,N_7202,N_5606);
nand U10651 (N_10651,N_7916,N_5107);
xor U10652 (N_10652,N_6216,N_8612);
or U10653 (N_10653,N_5445,N_9856);
or U10654 (N_10654,N_8529,N_7213);
or U10655 (N_10655,N_7855,N_6684);
xor U10656 (N_10656,N_6141,N_6700);
nand U10657 (N_10657,N_7421,N_5256);
nor U10658 (N_10658,N_8652,N_5408);
and U10659 (N_10659,N_9476,N_8695);
or U10660 (N_10660,N_8995,N_8828);
nor U10661 (N_10661,N_7506,N_7043);
nor U10662 (N_10662,N_8098,N_9924);
xnor U10663 (N_10663,N_9039,N_6462);
or U10664 (N_10664,N_6793,N_6164);
nor U10665 (N_10665,N_7096,N_9121);
or U10666 (N_10666,N_8928,N_6024);
nand U10667 (N_10667,N_5067,N_6739);
and U10668 (N_10668,N_8875,N_6607);
and U10669 (N_10669,N_6850,N_9166);
xnor U10670 (N_10670,N_6784,N_8052);
nor U10671 (N_10671,N_9111,N_9734);
nor U10672 (N_10672,N_5214,N_5044);
and U10673 (N_10673,N_7492,N_9106);
xnor U10674 (N_10674,N_8589,N_5672);
nand U10675 (N_10675,N_8295,N_9784);
nor U10676 (N_10676,N_5181,N_7854);
or U10677 (N_10677,N_7686,N_7597);
xor U10678 (N_10678,N_9517,N_5731);
nand U10679 (N_10679,N_5679,N_7931);
nor U10680 (N_10680,N_6725,N_7566);
or U10681 (N_10681,N_5763,N_7762);
nand U10682 (N_10682,N_9505,N_5310);
nand U10683 (N_10683,N_6446,N_9951);
or U10684 (N_10684,N_7135,N_8280);
xor U10685 (N_10685,N_6255,N_5819);
nor U10686 (N_10686,N_6196,N_7351);
xor U10687 (N_10687,N_9360,N_8120);
or U10688 (N_10688,N_9864,N_7765);
xnor U10689 (N_10689,N_6854,N_5654);
nor U10690 (N_10690,N_7473,N_6143);
nor U10691 (N_10691,N_8747,N_8176);
and U10692 (N_10692,N_5984,N_7123);
nor U10693 (N_10693,N_8499,N_7821);
and U10694 (N_10694,N_5202,N_9011);
or U10695 (N_10695,N_6133,N_7766);
nand U10696 (N_10696,N_7699,N_6333);
or U10697 (N_10697,N_8593,N_8932);
nor U10698 (N_10698,N_9921,N_5007);
and U10699 (N_10699,N_9832,N_9077);
nor U10700 (N_10700,N_7324,N_5103);
nand U10701 (N_10701,N_7474,N_7770);
xor U10702 (N_10702,N_5341,N_7632);
and U10703 (N_10703,N_7417,N_8224);
and U10704 (N_10704,N_8629,N_5497);
or U10705 (N_10705,N_5170,N_9868);
and U10706 (N_10706,N_5166,N_6183);
nor U10707 (N_10707,N_9703,N_6689);
nand U10708 (N_10708,N_5338,N_5299);
nand U10709 (N_10709,N_9721,N_7582);
and U10710 (N_10710,N_8789,N_8074);
or U10711 (N_10711,N_9271,N_9722);
nand U10712 (N_10712,N_5530,N_6223);
and U10713 (N_10713,N_5405,N_7794);
nor U10714 (N_10714,N_6782,N_6862);
nor U10715 (N_10715,N_9930,N_7365);
nor U10716 (N_10716,N_8368,N_5769);
and U10717 (N_10717,N_8720,N_8771);
xnor U10718 (N_10718,N_6972,N_6340);
or U10719 (N_10719,N_8416,N_9587);
and U10720 (N_10720,N_6654,N_9210);
or U10721 (N_10721,N_8531,N_6105);
nand U10722 (N_10722,N_9349,N_5875);
or U10723 (N_10723,N_5237,N_8482);
nand U10724 (N_10724,N_9968,N_7354);
nor U10725 (N_10725,N_8354,N_9892);
nor U10726 (N_10726,N_6578,N_9130);
nor U10727 (N_10727,N_7583,N_6707);
or U10728 (N_10728,N_5019,N_7001);
and U10729 (N_10729,N_6199,N_7628);
xnor U10730 (N_10730,N_9631,N_6488);
xnor U10731 (N_10731,N_8820,N_9133);
nand U10732 (N_10732,N_8502,N_6409);
xor U10733 (N_10733,N_8915,N_7523);
nor U10734 (N_10734,N_8462,N_9809);
nor U10735 (N_10735,N_9314,N_5486);
nand U10736 (N_10736,N_8383,N_5598);
nand U10737 (N_10737,N_5011,N_7483);
or U10738 (N_10738,N_6215,N_8223);
xnor U10739 (N_10739,N_6761,N_6168);
xor U10740 (N_10740,N_5594,N_8693);
nand U10741 (N_10741,N_9429,N_8270);
and U10742 (N_10742,N_5262,N_6967);
nor U10743 (N_10743,N_7830,N_9455);
nor U10744 (N_10744,N_7393,N_7580);
and U10745 (N_10745,N_7102,N_9040);
xor U10746 (N_10746,N_7889,N_7169);
nor U10747 (N_10747,N_8374,N_5292);
and U10748 (N_10748,N_9364,N_5284);
nand U10749 (N_10749,N_6759,N_8538);
nor U10750 (N_10750,N_8155,N_9766);
nor U10751 (N_10751,N_9562,N_9980);
and U10752 (N_10752,N_7106,N_6772);
nor U10753 (N_10753,N_5595,N_9818);
xnor U10754 (N_10754,N_5150,N_9224);
nor U10755 (N_10755,N_7120,N_9475);
nor U10756 (N_10756,N_6865,N_8876);
xnor U10757 (N_10757,N_5487,N_7937);
nand U10758 (N_10758,N_8574,N_8207);
nand U10759 (N_10759,N_8780,N_7588);
nor U10760 (N_10760,N_7860,N_6526);
nand U10761 (N_10761,N_6181,N_7302);
nor U10762 (N_10762,N_5670,N_9117);
nand U10763 (N_10763,N_6166,N_9577);
nor U10764 (N_10764,N_9537,N_8839);
and U10765 (N_10765,N_8080,N_8265);
and U10766 (N_10766,N_7577,N_9874);
nor U10767 (N_10767,N_7734,N_8194);
or U10768 (N_10768,N_8940,N_7573);
xor U10769 (N_10769,N_7944,N_7341);
nor U10770 (N_10770,N_8609,N_7401);
xor U10771 (N_10771,N_5609,N_7391);
xnor U10772 (N_10772,N_5273,N_5477);
or U10773 (N_10773,N_9828,N_7675);
and U10774 (N_10774,N_8760,N_7340);
or U10775 (N_10775,N_8414,N_6476);
and U10776 (N_10776,N_6365,N_5221);
or U10777 (N_10777,N_5123,N_5537);
nor U10778 (N_10778,N_7418,N_8678);
and U10779 (N_10779,N_5631,N_7117);
nor U10780 (N_10780,N_9183,N_6984);
nand U10781 (N_10781,N_5139,N_5219);
and U10782 (N_10782,N_9819,N_5488);
or U10783 (N_10783,N_9617,N_9757);
nand U10784 (N_10784,N_9408,N_9820);
nor U10785 (N_10785,N_6868,N_8396);
nor U10786 (N_10786,N_6610,N_5775);
or U10787 (N_10787,N_8973,N_9629);
and U10788 (N_10788,N_9526,N_8981);
and U10789 (N_10789,N_6653,N_6558);
or U10790 (N_10790,N_9287,N_6336);
and U10791 (N_10791,N_9144,N_6912);
or U10792 (N_10792,N_6903,N_6518);
nand U10793 (N_10793,N_8882,N_7730);
and U10794 (N_10794,N_7372,N_7669);
nor U10795 (N_10795,N_6792,N_5970);
nor U10796 (N_10796,N_9507,N_9070);
or U10797 (N_10797,N_8555,N_8062);
xnor U10798 (N_10798,N_9068,N_8783);
or U10799 (N_10799,N_6329,N_5882);
nor U10800 (N_10800,N_6553,N_7055);
nor U10801 (N_10801,N_8162,N_9079);
xnor U10802 (N_10802,N_8551,N_6289);
nor U10803 (N_10803,N_8626,N_7795);
and U10804 (N_10804,N_9218,N_8533);
or U10805 (N_10805,N_9064,N_9982);
nand U10806 (N_10806,N_7684,N_7723);
and U10807 (N_10807,N_5079,N_8329);
xnor U10808 (N_10808,N_6091,N_6987);
xor U10809 (N_10809,N_6517,N_7429);
and U10810 (N_10810,N_5873,N_7318);
nand U10811 (N_10811,N_7800,N_6901);
and U10812 (N_10812,N_9304,N_5891);
and U10813 (N_10813,N_5899,N_6068);
nand U10814 (N_10814,N_7612,N_7880);
and U10815 (N_10815,N_8987,N_5469);
or U10816 (N_10816,N_6320,N_8628);
nand U10817 (N_10817,N_5161,N_5217);
and U10818 (N_10818,N_8599,N_7692);
or U10819 (N_10819,N_6109,N_8553);
xor U10820 (N_10820,N_5677,N_7366);
nor U10821 (N_10821,N_6780,N_8946);
nand U10822 (N_10822,N_7693,N_6343);
nor U10823 (N_10823,N_7805,N_8230);
and U10824 (N_10824,N_7964,N_7553);
nor U10825 (N_10825,N_7244,N_9199);
or U10826 (N_10826,N_6608,N_7320);
and U10827 (N_10827,N_5980,N_7004);
or U10828 (N_10828,N_6830,N_7808);
xnor U10829 (N_10829,N_6104,N_6900);
nor U10830 (N_10830,N_6419,N_8081);
xnor U10831 (N_10831,N_5260,N_9197);
and U10832 (N_10832,N_5934,N_7008);
or U10833 (N_10833,N_6313,N_5065);
nand U10834 (N_10834,N_6974,N_6810);
nor U10835 (N_10835,N_6354,N_5951);
nor U10836 (N_10836,N_6844,N_6560);
nand U10837 (N_10837,N_6688,N_8541);
nand U10838 (N_10838,N_9801,N_5056);
nor U10839 (N_10839,N_6245,N_6281);
or U10840 (N_10840,N_6161,N_7859);
and U10841 (N_10841,N_8854,N_8157);
xor U10842 (N_10842,N_9223,N_9052);
and U10843 (N_10843,N_6845,N_7312);
nor U10844 (N_10844,N_5927,N_8147);
xor U10845 (N_10845,N_5696,N_7082);
nand U10846 (N_10846,N_8749,N_7510);
nand U10847 (N_10847,N_9641,N_9634);
nor U10848 (N_10848,N_5117,N_9229);
xor U10849 (N_10849,N_7498,N_7867);
xor U10850 (N_10850,N_6117,N_7869);
or U10851 (N_10851,N_8419,N_7264);
nor U10852 (N_10852,N_7392,N_9462);
nand U10853 (N_10853,N_6675,N_8921);
nor U10854 (N_10854,N_6208,N_9249);
nor U10855 (N_10855,N_5905,N_6049);
nor U10856 (N_10856,N_6052,N_9933);
or U10857 (N_10857,N_7355,N_5979);
nand U10858 (N_10858,N_9715,N_9454);
xnor U10859 (N_10859,N_6394,N_6144);
xnor U10860 (N_10860,N_8545,N_7558);
nor U10861 (N_10861,N_8637,N_8408);
xor U10862 (N_10862,N_9756,N_9233);
nor U10863 (N_10863,N_9204,N_6767);
xnor U10864 (N_10864,N_9277,N_6108);
nand U10865 (N_10865,N_9296,N_8879);
nor U10866 (N_10866,N_7296,N_9489);
nand U10867 (N_10867,N_6531,N_8580);
nor U10868 (N_10868,N_9791,N_5085);
or U10869 (N_10869,N_6489,N_8428);
nor U10870 (N_10870,N_6802,N_8158);
and U10871 (N_10871,N_8446,N_9348);
nand U10872 (N_10872,N_9193,N_8591);
xor U10873 (N_10873,N_7020,N_5896);
and U10874 (N_10874,N_5032,N_7480);
or U10875 (N_10875,N_5585,N_9467);
xor U10876 (N_10876,N_5391,N_6884);
xor U10877 (N_10877,N_7295,N_5339);
nor U10878 (N_10878,N_8901,N_6736);
and U10879 (N_10879,N_9125,N_9706);
nor U10880 (N_10880,N_5801,N_8923);
nand U10881 (N_10881,N_9793,N_9644);
xnor U10882 (N_10882,N_6482,N_7409);
and U10883 (N_10883,N_8153,N_6544);
nor U10884 (N_10884,N_7847,N_8225);
or U10885 (N_10885,N_8397,N_8311);
nand U10886 (N_10886,N_8263,N_7084);
and U10887 (N_10887,N_6190,N_8307);
xor U10888 (N_10888,N_8166,N_6067);
and U10889 (N_10889,N_6236,N_8690);
and U10890 (N_10890,N_7007,N_6428);
nor U10891 (N_10891,N_8868,N_7060);
and U10892 (N_10892,N_9115,N_9876);
and U10893 (N_10893,N_9808,N_5021);
xor U10894 (N_10894,N_9387,N_5510);
or U10895 (N_10895,N_8704,N_7657);
nand U10896 (N_10896,N_7536,N_8740);
or U10897 (N_10897,N_6648,N_6632);
xnor U10898 (N_10898,N_7208,N_6670);
nand U10899 (N_10899,N_6729,N_7339);
nand U10900 (N_10900,N_5180,N_8534);
xnor U10901 (N_10901,N_7526,N_8409);
nor U10902 (N_10902,N_6220,N_7024);
nor U10903 (N_10903,N_8537,N_8085);
xnor U10904 (N_10904,N_8680,N_9640);
xor U10905 (N_10905,N_9269,N_7773);
nor U10906 (N_10906,N_8219,N_7286);
and U10907 (N_10907,N_6390,N_9046);
xnor U10908 (N_10908,N_7724,N_6630);
and U10909 (N_10909,N_5675,N_5113);
nand U10910 (N_10910,N_5372,N_7961);
nor U10911 (N_10911,N_5479,N_8506);
and U10912 (N_10912,N_9535,N_6000);
nor U10913 (N_10913,N_9362,N_6756);
xnor U10914 (N_10914,N_6726,N_7028);
xor U10915 (N_10915,N_5820,N_8909);
or U10916 (N_10916,N_6421,N_8031);
nand U10917 (N_10917,N_9321,N_9278);
and U10918 (N_10918,N_6009,N_9155);
and U10919 (N_10919,N_7647,N_5962);
or U10920 (N_10920,N_8552,N_9324);
or U10921 (N_10921,N_5157,N_5798);
nor U10922 (N_10922,N_9840,N_9575);
and U10923 (N_10923,N_9632,N_5717);
or U10924 (N_10924,N_7138,N_7206);
nand U10925 (N_10925,N_5088,N_7449);
xnor U10926 (N_10926,N_9967,N_9678);
nor U10927 (N_10927,N_9493,N_7262);
xor U10928 (N_10928,N_7427,N_6991);
or U10929 (N_10929,N_7740,N_7717);
or U10930 (N_10930,N_5992,N_5985);
or U10931 (N_10931,N_8172,N_9162);
or U10932 (N_10932,N_5833,N_5792);
and U10933 (N_10933,N_5901,N_5616);
nor U10934 (N_10934,N_6111,N_5757);
and U10935 (N_10935,N_8817,N_7277);
nand U10936 (N_10936,N_5697,N_7174);
or U10937 (N_10937,N_8261,N_9424);
xnor U10938 (N_10938,N_7620,N_9614);
or U10939 (N_10939,N_5132,N_8867);
nand U10940 (N_10940,N_9041,N_9529);
or U10941 (N_10941,N_9363,N_8767);
and U10942 (N_10942,N_5038,N_5728);
nor U10943 (N_10943,N_6054,N_9409);
xor U10944 (N_10944,N_7199,N_9351);
xor U10945 (N_10945,N_9400,N_8112);
xor U10946 (N_10946,N_7349,N_8421);
xnor U10947 (N_10947,N_9316,N_5028);
xnor U10948 (N_10948,N_9112,N_6268);
and U10949 (N_10949,N_5006,N_8812);
and U10950 (N_10950,N_5536,N_9014);
and U10951 (N_10951,N_9890,N_9177);
xnor U10952 (N_10952,N_6892,N_5869);
xnor U10953 (N_10953,N_5187,N_5519);
nor U10954 (N_10954,N_7997,N_6396);
nor U10955 (N_10955,N_5197,N_9275);
or U10956 (N_10956,N_7966,N_5266);
or U10957 (N_10957,N_7791,N_9404);
and U10958 (N_10958,N_9460,N_9423);
and U10959 (N_10959,N_7919,N_7705);
nor U10960 (N_10960,N_9603,N_5719);
and U10961 (N_10961,N_5704,N_9297);
nand U10962 (N_10962,N_7499,N_8467);
nor U10963 (N_10963,N_7528,N_8028);
nor U10964 (N_10964,N_7397,N_8804);
nor U10965 (N_10965,N_6092,N_9086);
nand U10966 (N_10966,N_6011,N_8245);
and U10967 (N_10967,N_8430,N_8285);
or U10968 (N_10968,N_6693,N_5323);
nand U10969 (N_10969,N_7041,N_9227);
or U10970 (N_10970,N_7959,N_9761);
nand U10971 (N_10971,N_7949,N_9983);
nand U10972 (N_10972,N_8348,N_8936);
xnor U10973 (N_10973,N_6047,N_5087);
or U10974 (N_10974,N_5200,N_8827);
nor U10975 (N_10975,N_9028,N_7737);
and U10976 (N_10976,N_6678,N_5475);
xor U10977 (N_10977,N_9570,N_6981);
xnor U10978 (N_10978,N_5040,N_8937);
nand U10979 (N_10979,N_5461,N_9906);
nor U10980 (N_10980,N_7776,N_6346);
nand U10981 (N_10981,N_9384,N_8567);
nand U10982 (N_10982,N_5244,N_9927);
nand U10983 (N_10983,N_8459,N_9099);
and U10984 (N_10984,N_6747,N_9985);
xnor U10985 (N_10985,N_5830,N_5272);
nor U10986 (N_10986,N_9251,N_7660);
nand U10987 (N_10987,N_6605,N_7995);
and U10988 (N_10988,N_7785,N_8914);
or U10989 (N_10989,N_7279,N_6557);
or U10990 (N_10990,N_7259,N_8297);
xor U10991 (N_10991,N_7046,N_9619);
nand U10992 (N_10992,N_9571,N_5306);
nor U10993 (N_10993,N_7171,N_8717);
xnor U10994 (N_10994,N_6820,N_7204);
nand U10995 (N_10995,N_9555,N_6521);
xor U10996 (N_10996,N_5650,N_7238);
nand U10997 (N_10997,N_8370,N_8004);
xnor U10998 (N_10998,N_5653,N_7088);
and U10999 (N_10999,N_8231,N_8588);
or U11000 (N_11000,N_5222,N_9669);
or U11001 (N_11001,N_5282,N_5351);
and U11002 (N_11002,N_5098,N_5131);
nor U11003 (N_11003,N_7789,N_6121);
and U11004 (N_11004,N_6555,N_6254);
xor U11005 (N_11005,N_6455,N_9545);
and U11006 (N_11006,N_6506,N_5039);
nor U11007 (N_11007,N_5186,N_8549);
or U11008 (N_11008,N_5593,N_6007);
nor U11009 (N_11009,N_9392,N_9994);
and U11010 (N_11010,N_7078,N_6376);
nand U11011 (N_11011,N_7333,N_6204);
and U11012 (N_11012,N_7932,N_6611);
nor U11013 (N_11013,N_8208,N_5629);
and U11014 (N_11014,N_7530,N_7453);
xor U11015 (N_11015,N_7011,N_6647);
nand U11016 (N_11016,N_8958,N_9690);
nand U11017 (N_11017,N_9434,N_9601);
nor U11018 (N_11018,N_6870,N_8856);
and U11019 (N_11019,N_6279,N_8661);
xnor U11020 (N_11020,N_8405,N_8595);
or U11021 (N_11021,N_9021,N_6720);
nor U11022 (N_11022,N_9894,N_9789);
xnor U11023 (N_11023,N_6122,N_8980);
nor U11024 (N_11024,N_9290,N_7742);
xnor U11025 (N_11025,N_9464,N_8407);
and U11026 (N_11026,N_7247,N_9962);
and U11027 (N_11027,N_9612,N_9857);
nand U11028 (N_11028,N_6487,N_7343);
xor U11029 (N_11029,N_5233,N_5572);
or U11030 (N_11030,N_5440,N_8048);
nand U11031 (N_11031,N_8560,N_7991);
and U11032 (N_11032,N_8264,N_7538);
nor U11033 (N_11033,N_5733,N_5740);
xor U11034 (N_11034,N_7212,N_6926);
nand U11035 (N_11035,N_8795,N_8753);
and U11036 (N_11036,N_7844,N_6996);
nand U11037 (N_11037,N_8432,N_9020);
nor U11038 (N_11038,N_6021,N_6469);
or U11039 (N_11039,N_6551,N_9139);
nand U11040 (N_11040,N_5956,N_9327);
or U11041 (N_11041,N_6434,N_6359);
nand U11042 (N_11042,N_7513,N_9242);
or U11043 (N_11043,N_5773,N_5688);
or U11044 (N_11044,N_6478,N_7442);
nor U11045 (N_11045,N_8511,N_9171);
nor U11046 (N_11046,N_5379,N_5971);
and U11047 (N_11047,N_7764,N_9699);
and U11048 (N_11048,N_9399,N_7631);
and U11049 (N_11049,N_5363,N_7909);
nor U11050 (N_11050,N_6699,N_5551);
nor U11051 (N_11051,N_7683,N_5964);
or U11052 (N_11052,N_6944,N_6513);
nor U11053 (N_11053,N_5225,N_6988);
and U11054 (N_11054,N_6812,N_7774);
nor U11055 (N_11055,N_6613,N_6408);
xnor U11056 (N_11056,N_9624,N_9729);
and U11057 (N_11057,N_9652,N_9657);
xor U11058 (N_11058,N_7903,N_5952);
nand U11059 (N_11059,N_7154,N_9751);
nor U11060 (N_11060,N_5349,N_9679);
and U11061 (N_11061,N_7189,N_9333);
or U11062 (N_11062,N_6382,N_5277);
nand U11063 (N_11063,N_7076,N_6591);
nor U11064 (N_11064,N_6650,N_8666);
and U11065 (N_11065,N_6690,N_9302);
nand U11066 (N_11066,N_6515,N_5287);
xnor U11067 (N_11067,N_9260,N_9257);
or U11068 (N_11068,N_6740,N_8257);
and U11069 (N_11069,N_9274,N_6749);
nand U11070 (N_11070,N_7452,N_5526);
nand U11071 (N_11071,N_8394,N_6939);
nor U11072 (N_11072,N_9939,N_8347);
or U11073 (N_11073,N_7304,N_6392);
xnor U11074 (N_11074,N_8040,N_6858);
nand U11075 (N_11075,N_6350,N_7404);
nand U11076 (N_11076,N_7912,N_5662);
nor U11077 (N_11077,N_9220,N_5490);
nor U11078 (N_11078,N_6001,N_6766);
nand U11079 (N_11079,N_8631,N_6156);
and U11080 (N_11080,N_5652,N_9731);
and U11081 (N_11081,N_8950,N_9628);
xnor U11082 (N_11082,N_9518,N_7939);
nor U11083 (N_11083,N_6559,N_6964);
nor U11084 (N_11084,N_6044,N_9289);
and U11085 (N_11085,N_9389,N_6556);
nand U11086 (N_11086,N_7243,N_9131);
or U11087 (N_11087,N_8360,N_8933);
and U11088 (N_11088,N_9329,N_9500);
xnor U11089 (N_11089,N_6588,N_9385);
nand U11090 (N_11090,N_6058,N_9711);
nor U11091 (N_11091,N_7574,N_5963);
nand U11092 (N_11092,N_9009,N_7828);
nand U11093 (N_11093,N_6075,N_7042);
nand U11094 (N_11094,N_6537,N_5313);
xnor U11095 (N_11095,N_9437,N_8963);
xnor U11096 (N_11096,N_8340,N_6923);
or U11097 (N_11097,N_9769,N_5004);
nor U11098 (N_11098,N_9241,N_7825);
and U11099 (N_11099,N_8328,N_5581);
xor U11100 (N_11100,N_6050,N_5218);
and U11101 (N_11101,N_7383,N_9554);
and U11102 (N_11102,N_9932,N_5878);
nand U11103 (N_11103,N_7462,N_6261);
nor U11104 (N_11104,N_6696,N_9450);
and U11105 (N_11105,N_5080,N_6867);
and U11106 (N_11106,N_7256,N_8871);
nor U11107 (N_11107,N_5022,N_5432);
nand U11108 (N_11108,N_9005,N_7375);
or U11109 (N_11109,N_8109,N_9595);
and U11110 (N_11110,N_5566,N_5877);
xor U11111 (N_11111,N_6965,N_8058);
and U11112 (N_11112,N_5245,N_7518);
and U11113 (N_11113,N_7984,N_7682);
nor U11114 (N_11114,N_7400,N_5257);
or U11115 (N_11115,N_9497,N_6023);
nand U11116 (N_11116,N_7936,N_8691);
xnor U11117 (N_11117,N_9418,N_5543);
nand U11118 (N_11118,N_9149,N_8813);
nor U11119 (N_11119,N_6801,N_8410);
xnor U11120 (N_11120,N_7438,N_9668);
xor U11121 (N_11121,N_8445,N_6292);
nand U11122 (N_11122,N_9540,N_9458);
nand U11123 (N_11123,N_9284,N_9949);
or U11124 (N_11124,N_5433,N_7748);
xnor U11125 (N_11125,N_8038,N_6384);
nor U11126 (N_11126,N_8220,N_7218);
nor U11127 (N_11127,N_9971,N_8212);
nor U11128 (N_11128,N_6682,N_6936);
or U11129 (N_11129,N_8608,N_6825);
and U11130 (N_11130,N_9664,N_5871);
and U11131 (N_11131,N_5141,N_7215);
nand U11132 (N_11132,N_7947,N_9401);
nand U11133 (N_11133,N_9402,N_5724);
nand U11134 (N_11134,N_9063,N_9051);
or U11135 (N_11135,N_7626,N_8483);
nor U11136 (N_11136,N_8507,N_8337);
or U11137 (N_11137,N_5527,N_8072);
nor U11138 (N_11138,N_7361,N_8113);
nand U11139 (N_11139,N_6096,N_8727);
and U11140 (N_11140,N_7406,N_9986);
nor U11141 (N_11141,N_6288,N_6457);
and U11142 (N_11142,N_7472,N_6230);
or U11143 (N_11143,N_9067,N_8137);
nor U11144 (N_11144,N_8050,N_8259);
or U11145 (N_11145,N_6229,N_5493);
or U11146 (N_11146,N_7756,N_9851);
and U11147 (N_11147,N_7595,N_8234);
and U11148 (N_11148,N_7158,N_7183);
nand U11149 (N_11149,N_5780,N_9797);
and U11150 (N_11150,N_8577,N_5455);
nor U11151 (N_11151,N_9096,N_9232);
and U11152 (N_11152,N_7668,N_9120);
xor U11153 (N_11153,N_6335,N_7527);
or U11154 (N_11154,N_9156,N_9499);
and U11155 (N_11155,N_9767,N_6994);
nor U11156 (N_11156,N_5438,N_9594);
nand U11157 (N_11157,N_7922,N_6885);
nor U11158 (N_11158,N_7958,N_9071);
xnor U11159 (N_11159,N_7951,N_6898);
xor U11160 (N_11160,N_6193,N_6202);
nand U11161 (N_11161,N_5782,N_6201);
xor U11162 (N_11162,N_5659,N_6719);
and U11163 (N_11163,N_5851,N_8939);
nand U11164 (N_11164,N_6293,N_8250);
nor U11165 (N_11165,N_8872,N_5239);
nand U11166 (N_11166,N_8175,N_9548);
nand U11167 (N_11167,N_6314,N_9977);
nor U11168 (N_11168,N_9771,N_8066);
nand U11169 (N_11169,N_6045,N_5926);
nor U11170 (N_11170,N_9313,N_6226);
and U11171 (N_11171,N_5375,N_6377);
nor U11172 (N_11172,N_6534,N_9212);
and U11173 (N_11173,N_6318,N_9380);
nor U11174 (N_11174,N_7619,N_7178);
nor U11175 (N_11175,N_6406,N_9536);
nand U11176 (N_11176,N_5790,N_5070);
xnor U11177 (N_11177,N_7665,N_6791);
xor U11178 (N_11178,N_9520,N_6807);
nor U11179 (N_11179,N_7035,N_5271);
and U11180 (N_11180,N_8173,N_9775);
and U11181 (N_11181,N_9674,N_9936);
and U11182 (N_11182,N_8586,N_9109);
xor U11183 (N_11183,N_6962,N_5590);
nand U11184 (N_11184,N_9192,N_5541);
or U11185 (N_11185,N_9752,N_9730);
or U11186 (N_11186,N_9733,N_6623);
or U11187 (N_11187,N_8885,N_8334);
xor U11188 (N_11188,N_9116,N_9428);
nand U11189 (N_11189,N_6456,N_9853);
nand U11190 (N_11190,N_6755,N_5977);
or U11191 (N_11191,N_9369,N_9610);
xnor U11192 (N_11192,N_8540,N_7232);
xor U11193 (N_11193,N_6441,N_9701);
nor U11194 (N_11194,N_8030,N_6407);
or U11195 (N_11195,N_7410,N_9058);
nand U11196 (N_11196,N_8395,N_9474);
nor U11197 (N_11197,N_6724,N_5789);
xnor U11198 (N_11198,N_6664,N_7021);
nand U11199 (N_11199,N_6828,N_9234);
and U11200 (N_11200,N_7677,N_5442);
or U11201 (N_11201,N_6149,N_5613);
nand U11202 (N_11202,N_9984,N_8890);
nor U11203 (N_11203,N_7225,N_6118);
nor U11204 (N_11204,N_9480,N_9154);
nand U11205 (N_11205,N_9317,N_6547);
nor U11206 (N_11206,N_7698,N_9148);
or U11207 (N_11207,N_6003,N_9273);
nor U11208 (N_11208,N_8734,N_7570);
and U11209 (N_11209,N_9330,N_6093);
nand U11210 (N_11210,N_9185,N_7522);
nor U11211 (N_11211,N_5159,N_9543);
nor U11212 (N_11212,N_6298,N_7036);
xnor U11213 (N_11213,N_5242,N_5548);
and U11214 (N_11214,N_5993,N_6386);
xor U11215 (N_11215,N_9169,N_8156);
or U11216 (N_11216,N_9916,N_9104);
or U11217 (N_11217,N_5274,N_9891);
and U11218 (N_11218,N_5164,N_7755);
or U11219 (N_11219,N_5243,N_7456);
nor U11220 (N_11220,N_8014,N_8617);
nand U11221 (N_11221,N_5953,N_5987);
and U11222 (N_11222,N_6307,N_7839);
nor U11223 (N_11223,N_6909,N_7287);
or U11224 (N_11224,N_9433,N_5054);
and U11225 (N_11225,N_5194,N_7803);
nand U11226 (N_11226,N_8547,N_5404);
or U11227 (N_11227,N_6617,N_6661);
and U11228 (N_11228,N_8473,N_9336);
nor U11229 (N_11229,N_8849,N_8049);
and U11230 (N_11230,N_5447,N_6634);
and U11231 (N_11231,N_9725,N_9566);
nand U11232 (N_11232,N_6366,N_8755);
nor U11233 (N_11233,N_8619,N_7714);
or U11234 (N_11234,N_6573,N_8215);
xnor U11235 (N_11235,N_5315,N_9636);
nand U11236 (N_11236,N_8232,N_5231);
or U11237 (N_11237,N_5835,N_7086);
xnor U11238 (N_11238,N_9581,N_7289);
or U11239 (N_11239,N_9033,N_9686);
nor U11240 (N_11240,N_8736,N_5610);
xnor U11241 (N_11241,N_7627,N_6250);
or U11242 (N_11242,N_5533,N_5886);
or U11243 (N_11243,N_7985,N_9838);
nand U11244 (N_11244,N_8016,N_8135);
xnor U11245 (N_11245,N_7873,N_7362);
or U11246 (N_11246,N_8891,N_6224);
and U11247 (N_11247,N_6262,N_8406);
xnor U11248 (N_11248,N_6692,N_8938);
nor U11249 (N_11249,N_6789,N_6816);
nand U11250 (N_11250,N_9782,N_8054);
and U11251 (N_11251,N_5110,N_7405);
or U11252 (N_11252,N_9538,N_5421);
nor U11253 (N_11253,N_5191,N_6191);
nor U11254 (N_11254,N_6533,N_6673);
and U11255 (N_11255,N_5208,N_5436);
nor U11256 (N_11256,N_6800,N_7614);
and U11257 (N_11257,N_8222,N_6454);
xnor U11258 (N_11258,N_8277,N_8989);
and U11259 (N_11259,N_9975,N_8491);
nand U11260 (N_11260,N_7702,N_7989);
nand U11261 (N_11261,N_9696,N_9776);
xor U11262 (N_11262,N_8929,N_6027);
and U11263 (N_11263,N_5579,N_9206);
and U11264 (N_11264,N_8344,N_8454);
and U11265 (N_11265,N_6508,N_8241);
and U11266 (N_11266,N_9083,N_8475);
nand U11267 (N_11267,N_5204,N_7851);
and U11268 (N_11268,N_8039,N_9988);
and U11269 (N_11269,N_6598,N_9947);
nor U11270 (N_11270,N_5135,N_6140);
nor U11271 (N_11271,N_5518,N_7388);
or U11272 (N_11272,N_5994,N_6157);
or U11273 (N_11273,N_6561,N_5286);
nand U11274 (N_11274,N_9110,N_8917);
nand U11275 (N_11275,N_7679,N_6203);
nor U11276 (N_11276,N_6160,N_7778);
nand U11277 (N_11277,N_8443,N_8659);
and U11278 (N_11278,N_8841,N_7314);
xor U11279 (N_11279,N_6503,N_9207);
xnor U11280 (N_11280,N_8333,N_5950);
and U11281 (N_11281,N_9990,N_7080);
nor U11282 (N_11282,N_8450,N_5503);
and U11283 (N_11283,N_6847,N_7978);
nand U11284 (N_11284,N_8185,N_5776);
nand U11285 (N_11285,N_7820,N_8345);
nor U11286 (N_11286,N_5069,N_9100);
and U11287 (N_11287,N_7226,N_5057);
nand U11288 (N_11288,N_8437,N_9461);
nor U11289 (N_11289,N_6728,N_8584);
and U11290 (N_11290,N_6507,N_6540);
nor U11291 (N_11291,N_9406,N_8228);
or U11292 (N_11292,N_7446,N_7251);
nor U11293 (N_11293,N_5564,N_9050);
or U11294 (N_11294,N_7796,N_7697);
nand U11295 (N_11295,N_5190,N_8613);
nand U11296 (N_11296,N_7716,N_7152);
or U11297 (N_11297,N_8115,N_6897);
xor U11298 (N_11298,N_9527,N_7034);
xor U11299 (N_11299,N_8104,N_8464);
and U11300 (N_11300,N_8444,N_8705);
nand U11301 (N_11301,N_7298,N_5718);
and U11302 (N_11302,N_8576,N_7114);
and U11303 (N_11303,N_7294,N_8682);
nor U11304 (N_11304,N_6727,N_6852);
nand U11305 (N_11305,N_5636,N_8144);
or U11306 (N_11306,N_6660,N_5883);
nor U11307 (N_11307,N_7168,N_7611);
and U11308 (N_11308,N_5001,N_7268);
and U11309 (N_11309,N_6322,N_8886);
xor U11310 (N_11310,N_9707,N_8242);
or U11311 (N_11311,N_7470,N_7548);
xnor U11312 (N_11312,N_9623,N_7562);
and U11313 (N_11313,N_8474,N_6600);
xor U11314 (N_11314,N_7003,N_8401);
nand U11315 (N_11315,N_5400,N_9176);
or U11316 (N_11316,N_9383,N_8434);
nor U11317 (N_11317,N_6405,N_6977);
and U11318 (N_11318,N_7224,N_8468);
nand U11319 (N_11319,N_6015,N_9365);
nor U11320 (N_11320,N_8088,N_6437);
xnor U11321 (N_11321,N_9547,N_7050);
xor U11322 (N_11322,N_9236,N_5327);
nand U11323 (N_11323,N_8105,N_5743);
or U11324 (N_11324,N_6918,N_8192);
nor U11325 (N_11325,N_8633,N_8931);
nor U11326 (N_11326,N_9753,N_5807);
nand U11327 (N_11327,N_6364,N_9559);
nand U11328 (N_11328,N_7585,N_8011);
nor U11329 (N_11329,N_6423,N_6252);
and U11330 (N_11330,N_9739,N_7534);
nor U11331 (N_11331,N_7190,N_7010);
and U11332 (N_11332,N_6920,N_5768);
and U11333 (N_11333,N_5424,N_7896);
and U11334 (N_11334,N_5796,N_6950);
and U11335 (N_11335,N_7636,N_5967);
xnor U11336 (N_11336,N_6905,N_7112);
and U11337 (N_11337,N_8883,N_8379);
nand U11338 (N_11338,N_9209,N_5943);
nor U11339 (N_11339,N_5109,N_5555);
xnor U11340 (N_11340,N_7508,N_6301);
nor U11341 (N_11341,N_6587,N_8102);
or U11342 (N_11342,N_8075,N_5589);
and U11343 (N_11343,N_9007,N_5671);
xor U11344 (N_11344,N_8853,N_6165);
or U11345 (N_11345,N_9795,N_7758);
and U11346 (N_11346,N_7555,N_6460);
nor U11347 (N_11347,N_5168,N_7145);
xor U11348 (N_11348,N_7954,N_8884);
or U11349 (N_11349,N_6085,N_8530);
or U11350 (N_11350,N_5802,N_6797);
xor U11351 (N_11351,N_9395,N_6522);
nor U11352 (N_11352,N_8791,N_6877);
nand U11353 (N_11353,N_7713,N_8785);
or U11354 (N_11354,N_9430,N_9059);
xor U11355 (N_11355,N_7425,N_8388);
xor U11356 (N_11356,N_8303,N_8657);
xor U11357 (N_11357,N_8187,N_6086);
xnor U11358 (N_11358,N_7023,N_9966);
nor U11359 (N_11359,N_5999,N_5005);
xor U11360 (N_11360,N_8398,N_9862);
xor U11361 (N_11361,N_8240,N_5326);
xnor U11362 (N_11362,N_9334,N_8309);
and U11363 (N_11363,N_7385,N_7240);
nand U11364 (N_11364,N_6880,N_7198);
xor U11365 (N_11365,N_9780,N_5837);
and U11366 (N_11366,N_5337,N_9098);
or U11367 (N_11367,N_9606,N_9533);
nand U11368 (N_11368,N_6387,N_6754);
xnor U11369 (N_11369,N_9940,N_5687);
xnor U11370 (N_11370,N_5249,N_5736);
nand U11371 (N_11371,N_9661,N_8907);
and U11372 (N_11372,N_9457,N_6061);
xor U11373 (N_11373,N_9025,N_5361);
nor U11374 (N_11374,N_9226,N_7487);
or U11375 (N_11375,N_7940,N_5557);
xnor U11376 (N_11376,N_8427,N_6211);
xor U11377 (N_11377,N_7594,N_5325);
nand U11378 (N_11378,N_6345,N_6112);
or U11379 (N_11379,N_8179,N_5699);
or U11380 (N_11380,N_7177,N_9298);
or U11381 (N_11381,N_8248,N_6357);
xor U11382 (N_11382,N_5051,N_8316);
and U11383 (N_11383,N_5265,N_6200);
nor U11384 (N_11384,N_5026,N_7797);
or U11385 (N_11385,N_9807,N_8960);
nand U11386 (N_11386,N_6938,N_5791);
nand U11387 (N_11387,N_8546,N_8729);
or U11388 (N_11388,N_6979,N_8019);
xnor U11389 (N_11389,N_5111,N_9225);
nor U11390 (N_11390,N_5809,N_7861);
nand U11391 (N_11391,N_8322,N_8376);
nor U11392 (N_11392,N_7664,N_7358);
or U11393 (N_11393,N_9010,N_7162);
nand U11394 (N_11394,N_5599,N_5220);
nor U11395 (N_11395,N_8964,N_5995);
or U11396 (N_11396,N_5184,N_5797);
and U11397 (N_11397,N_7382,N_7000);
and U11398 (N_11398,N_8903,N_6921);
and U11399 (N_11399,N_6372,N_7942);
or U11400 (N_11400,N_6219,N_8870);
xor U11401 (N_11401,N_5036,N_8296);
xnor U11402 (N_11402,N_5165,N_6297);
xor U11403 (N_11403,N_5745,N_8969);
nand U11404 (N_11404,N_8221,N_9145);
xnor U11405 (N_11405,N_7130,N_7887);
xnor U11406 (N_11406,N_8535,N_9448);
xor U11407 (N_11407,N_6764,N_5591);
nor U11408 (N_11408,N_5415,N_8614);
nand U11409 (N_11409,N_8070,N_8034);
xor U11410 (N_11410,N_8233,N_6228);
nand U11411 (N_11411,N_8196,N_6945);
nand U11412 (N_11412,N_5983,N_7902);
nor U11413 (N_11413,N_5806,N_6251);
nor U11414 (N_11414,N_9486,N_5092);
or U11415 (N_11415,N_6065,N_5946);
nor U11416 (N_11416,N_5407,N_7885);
nand U11417 (N_11417,N_5991,N_9926);
nand U11418 (N_11418,N_6787,N_6426);
or U11419 (N_11419,N_7486,N_5263);
nand U11420 (N_11420,N_5390,N_7618);
or U11421 (N_11421,N_7249,N_9732);
or U11422 (N_11422,N_8006,N_5781);
nand U11423 (N_11423,N_7188,N_6706);
and U11424 (N_11424,N_9230,N_9481);
xor U11425 (N_11425,N_9716,N_8371);
nor U11426 (N_11426,N_5464,N_6929);
and U11427 (N_11427,N_8452,N_6260);
or U11428 (N_11428,N_9748,N_7833);
and U11429 (N_11429,N_7210,N_6657);
nand U11430 (N_11430,N_6817,N_7514);
or U11431 (N_11431,N_7235,N_9196);
nor U11432 (N_11432,N_7875,N_7288);
xor U11433 (N_11433,N_9453,N_6099);
nor U11434 (N_11434,N_9773,N_9783);
or U11435 (N_11435,N_7257,N_7201);
nor U11436 (N_11436,N_9216,N_5439);
and U11437 (N_11437,N_6147,N_9905);
or U11438 (N_11438,N_5817,N_5176);
nand U11439 (N_11439,N_9413,N_5506);
nor U11440 (N_11440,N_6859,N_8701);
and U11441 (N_11441,N_9366,N_6338);
xnor U11442 (N_11442,N_9995,N_9913);
and U11443 (N_11443,N_9180,N_9738);
nand U11444 (N_11444,N_7635,N_5573);
and U11445 (N_11445,N_8488,N_8315);
xor U11446 (N_11446,N_8837,N_5414);
xor U11447 (N_11447,N_5914,N_5815);
or U11448 (N_11448,N_5966,N_5990);
or U11449 (N_11449,N_7306,N_7767);
xnor U11450 (N_11450,N_9993,N_9893);
nand U11451 (N_11451,N_6803,N_9938);
and U11452 (N_11452,N_9792,N_7890);
nand U11453 (N_11453,N_6597,N_8822);
xnor U11454 (N_11454,N_6539,N_8425);
xnor U11455 (N_11455,N_8082,N_5546);
or U11456 (N_11456,N_6087,N_7603);
xnor U11457 (N_11457,N_8605,N_9060);
xor U11458 (N_11458,N_8097,N_7956);
xnor U11459 (N_11459,N_6295,N_5694);
and U11460 (N_11460,N_8456,N_5753);
nor U11461 (N_11461,N_9266,N_6928);
nor U11462 (N_11462,N_7493,N_8357);
nor U11463 (N_11463,N_5340,N_9579);
nor U11464 (N_11464,N_7542,N_7278);
nor U11465 (N_11465,N_6286,N_8286);
and U11466 (N_11466,N_8611,N_6309);
or U11467 (N_11467,N_5335,N_6129);
or U11468 (N_11468,N_8325,N_8479);
xor U11469 (N_11469,N_7781,N_6463);
and U11470 (N_11470,N_8850,N_9618);
or U11471 (N_11471,N_9080,N_9607);
and U11472 (N_11472,N_5823,N_5000);
or U11473 (N_11473,N_6039,N_5729);
and U11474 (N_11474,N_7654,N_9511);
nor U11475 (N_11475,N_6369,N_7641);
or U11476 (N_11476,N_9709,N_8136);
or U11477 (N_11477,N_9279,N_9082);
xor U11478 (N_11478,N_5648,N_5958);
and U11479 (N_11479,N_9946,N_6399);
nand U11480 (N_11480,N_5378,N_8198);
or U11481 (N_11481,N_7194,N_8673);
xor U11482 (N_11482,N_6625,N_8442);
or U11483 (N_11483,N_6494,N_7402);
nor U11484 (N_11484,N_5238,N_6638);
nor U11485 (N_11485,N_5732,N_9487);
nand U11486 (N_11486,N_7160,N_5099);
xor U11487 (N_11487,N_8625,N_9479);
nand U11488 (N_11488,N_8505,N_5199);
nand U11489 (N_11489,N_7267,N_7786);
or U11490 (N_11490,N_6134,N_7403);
or U11491 (N_11491,N_9749,N_5210);
and U11492 (N_11492,N_9043,N_6563);
or U11493 (N_11493,N_9915,N_5854);
or U11494 (N_11494,N_5267,N_6980);
nand U11495 (N_11495,N_6733,N_7575);
and U11496 (N_11496,N_7416,N_9959);
nand U11497 (N_11497,N_9616,N_9998);
nand U11498 (N_11498,N_5360,N_8496);
xnor U11499 (N_11499,N_8578,N_8160);
and U11500 (N_11500,N_5029,N_8304);
xnor U11501 (N_11501,N_8781,N_7056);
and U11502 (N_11502,N_8008,N_7598);
xnor U11503 (N_11503,N_7637,N_8400);
nor U11504 (N_11504,N_7323,N_5023);
xnor U11505 (N_11505,N_6005,N_8985);
xnor U11506 (N_11506,N_8204,N_5127);
nor U11507 (N_11507,N_9881,N_5268);
and U11508 (N_11508,N_8745,N_5517);
nor U11509 (N_11509,N_5516,N_8579);
and U11510 (N_11510,N_6774,N_6132);
and U11511 (N_11511,N_6940,N_9643);
and U11512 (N_11512,N_7090,N_9889);
and U11513 (N_11513,N_8077,N_9823);
xor U11514 (N_11514,N_7599,N_6917);
and U11515 (N_11515,N_7685,N_5215);
or U11516 (N_11516,N_6429,N_5232);
or U11517 (N_11517,N_7051,N_5147);
nor U11518 (N_11518,N_5852,N_7460);
nor U11519 (N_11519,N_8087,N_8477);
xnor U11520 (N_11520,N_7311,N_9267);
nand U11521 (N_11521,N_7926,N_7049);
or U11522 (N_11522,N_6358,N_7772);
xor U11523 (N_11523,N_7211,N_5142);
xnor U11524 (N_11524,N_8686,N_7408);
or U11525 (N_11525,N_6170,N_6057);
nand U11526 (N_11526,N_6031,N_9508);
or U11527 (N_11527,N_9525,N_7129);
or U11528 (N_11528,N_6002,N_8894);
nor U11529 (N_11529,N_5642,N_8372);
nor U11530 (N_11530,N_5682,N_5010);
nor U11531 (N_11531,N_7325,N_7134);
xor U11532 (N_11532,N_8380,N_6713);
nor U11533 (N_11533,N_8094,N_7141);
or U11534 (N_11534,N_9502,N_5531);
or U11535 (N_11535,N_5874,N_7466);
and U11536 (N_11536,N_8992,N_7798);
nor U11537 (N_11537,N_5255,N_7689);
and U11538 (N_11538,N_8802,N_8708);
or U11539 (N_11539,N_7420,N_6040);
nor U11540 (N_11540,N_5845,N_8644);
and U11541 (N_11541,N_6516,N_6287);
nand U11542 (N_11542,N_9585,N_6836);
or U11543 (N_11543,N_7031,N_6130);
or U11544 (N_11544,N_5576,N_7337);
xnor U11545 (N_11545,N_7814,N_7317);
or U11546 (N_11546,N_9659,N_8926);
xor U11547 (N_11547,N_5133,N_8321);
and U11548 (N_11548,N_5419,N_5177);
and U11549 (N_11549,N_8182,N_8152);
xor U11550 (N_11550,N_9127,N_7622);
xnor U11551 (N_11551,N_5842,N_7992);
or U11552 (N_11552,N_8902,N_8148);
nor U11553 (N_11553,N_6528,N_8787);
nand U11554 (N_11554,N_9161,N_9902);
xor U11555 (N_11555,N_9066,N_5622);
nor U11556 (N_11556,N_8596,N_6235);
and U11557 (N_11557,N_7132,N_6685);
nand U11558 (N_11558,N_9419,N_5294);
and U11559 (N_11559,N_8161,N_6448);
xor U11560 (N_11560,N_7927,N_6773);
and U11561 (N_11561,N_5224,N_9740);
xor U11562 (N_11562,N_8526,N_8466);
and U11563 (N_11563,N_7882,N_6276);
and U11564 (N_11564,N_8833,N_5655);
or U11565 (N_11565,N_5575,N_5163);
and U11566 (N_11566,N_5663,N_7589);
nand U11567 (N_11567,N_7941,N_7137);
and U11568 (N_11568,N_8125,N_5201);
or U11569 (N_11569,N_5114,N_7245);
or U11570 (N_11570,N_6548,N_8896);
xor U11571 (N_11571,N_5571,N_7371);
nor U11572 (N_11572,N_8140,N_5828);
and U11573 (N_11573,N_6546,N_8324);
xnor U11574 (N_11574,N_7062,N_5795);
and U11575 (N_11575,N_7052,N_6554);
and U11576 (N_11576,N_8495,N_8145);
xnor U11577 (N_11577,N_5665,N_5412);
xor U11578 (N_11578,N_6019,N_7072);
or U11579 (N_11579,N_8209,N_6037);
nand U11580 (N_11580,N_6095,N_9001);
or U11581 (N_11581,N_9821,N_5925);
nand U11582 (N_11582,N_6827,N_7650);
xnor U11583 (N_11583,N_8518,N_6856);
nor U11584 (N_11584,N_6832,N_6025);
and U11585 (N_11585,N_8561,N_6947);
xnor U11586 (N_11586,N_7495,N_9941);
nand U11587 (N_11587,N_6480,N_9779);
or U11588 (N_11588,N_5314,N_7999);
or U11589 (N_11589,N_9541,N_6447);
xor U11590 (N_11590,N_7363,N_7469);
nand U11591 (N_11591,N_8447,N_7116);
and U11592 (N_11592,N_7572,N_7866);
nor U11593 (N_11593,N_7281,N_7590);
nor U11594 (N_11594,N_8211,N_9880);
and U11595 (N_11595,N_9834,N_9443);
or U11596 (N_11596,N_9655,N_9372);
or U11597 (N_11597,N_8021,N_5978);
or U11598 (N_11598,N_7384,N_6734);
xnor U11599 (N_11599,N_7559,N_8974);
or U11600 (N_11600,N_9087,N_5465);
or U11601 (N_11601,N_7173,N_8851);
or U11602 (N_11602,N_5392,N_9925);
nand U11603 (N_11603,N_9182,N_7606);
nor U11604 (N_11604,N_8900,N_5884);
and U11605 (N_11605,N_6265,N_7176);
and U11606 (N_11606,N_8059,N_8971);
or U11607 (N_11607,N_9465,N_9501);
xnor U11608 (N_11608,N_7353,N_5735);
or U11609 (N_11609,N_9960,N_6381);
or U11610 (N_11610,N_7591,N_6198);
nand U11611 (N_11611,N_9320,N_6363);
and U11612 (N_11612,N_8217,N_8554);
xor U11613 (N_11613,N_6089,N_8634);
and U11614 (N_11614,N_5664,N_8808);
and U11615 (N_11615,N_9405,N_8620);
nand U11616 (N_11616,N_5368,N_5916);
nand U11617 (N_11617,N_8977,N_9865);
or U11618 (N_11618,N_7728,N_6355);
and U11619 (N_11619,N_9621,N_7516);
nor U11620 (N_11620,N_8091,N_9954);
nor U11621 (N_11621,N_7690,N_7827);
nand U11622 (N_11622,N_9215,N_6090);
nor U11623 (N_11623,N_5831,N_7246);
or U11624 (N_11624,N_9213,N_6714);
xor U11625 (N_11625,N_9746,N_7760);
xnor U11626 (N_11626,N_9425,N_6341);
or U11627 (N_11627,N_5588,N_8045);
xor U11628 (N_11628,N_7857,N_6841);
nand U11629 (N_11629,N_6778,N_8095);
xnor U11630 (N_11630,N_5126,N_7810);
or U11631 (N_11631,N_8823,N_5887);
and U11632 (N_11632,N_8471,N_8536);
and U11633 (N_11633,N_9914,N_7261);
nand U11634 (N_11634,N_5354,N_5861);
or U11635 (N_11635,N_6571,N_7037);
or U11636 (N_11636,N_5420,N_7236);
nand U11637 (N_11637,N_8117,N_7097);
xor U11638 (N_11638,N_5902,N_5844);
xnor U11639 (N_11639,N_8572,N_5399);
and U11640 (N_11640,N_9829,N_9469);
nor U11641 (N_11641,N_5348,N_6395);
xor U11642 (N_11642,N_6367,N_8676);
and U11643 (N_11643,N_8494,N_9672);
nand U11644 (N_11644,N_7933,N_7920);
or U11645 (N_11645,N_6762,N_6153);
nor U11646 (N_11646,N_6779,N_5350);
or U11647 (N_11647,N_6815,N_7661);
and U11648 (N_11648,N_6837,N_6687);
xor U11649 (N_11649,N_5766,N_5138);
nor U11650 (N_11650,N_9611,N_6621);
nor U11651 (N_11651,N_6115,N_7596);
nor U11652 (N_11652,N_5331,N_9157);
or U11653 (N_11653,N_8268,N_8924);
xnor U11654 (N_11654,N_6790,N_6992);
and U11655 (N_11655,N_6659,N_9439);
xor U11656 (N_11656,N_8956,N_9268);
nand U11657 (N_11657,N_9463,N_8227);
nor U11658 (N_11658,N_5090,N_7150);
nand U11659 (N_11659,N_9309,N_9231);
nor U11660 (N_11660,N_5917,N_5499);
or U11661 (N_11661,N_6082,N_9942);
nor U11662 (N_11662,N_8604,N_8440);
nand U11663 (N_11663,N_6924,N_8669);
xor U11664 (N_11664,N_5071,N_5909);
nand U11665 (N_11665,N_9718,N_5756);
and U11666 (N_11666,N_9513,N_7908);
and U11667 (N_11667,N_9534,N_5082);
and U11668 (N_11668,N_5784,N_7014);
nand U11669 (N_11669,N_6575,N_6271);
and U11670 (N_11670,N_8319,N_6500);
nor U11671 (N_11671,N_7531,N_5596);
nand U11672 (N_11672,N_7695,N_5169);
nor U11673 (N_11673,N_5342,N_7545);
nor U11674 (N_11674,N_9057,N_9955);
nor U11675 (N_11675,N_6347,N_5106);
nor U11676 (N_11676,N_9074,N_8339);
nor U11677 (N_11677,N_9583,N_8015);
nor U11678 (N_11678,N_5597,N_9589);
xor U11679 (N_11679,N_7263,N_7330);
nor U11680 (N_11680,N_8893,N_8469);
or U11681 (N_11681,N_8716,N_7451);
xnor U11682 (N_11682,N_9214,N_6615);
xor U11683 (N_11683,N_5774,N_9604);
or U11684 (N_11684,N_9065,N_9129);
xnor U11685 (N_11685,N_9432,N_7193);
nand U11686 (N_11686,N_7308,N_9519);
or U11687 (N_11687,N_7292,N_9367);
and U11688 (N_11688,N_5411,N_7709);
nand U11689 (N_11689,N_6214,N_9910);
nand U11690 (N_11690,N_6103,N_9539);
xnor U11691 (N_11691,N_7468,N_6834);
or U11692 (N_11692,N_8943,N_5730);
nand U11693 (N_11693,N_6349,N_6633);
nor U11694 (N_11694,N_9445,N_6440);
or U11695 (N_11695,N_9143,N_6481);
nand U11696 (N_11696,N_7649,N_6174);
xnor U11697 (N_11697,N_6146,N_9957);
xnor U11698 (N_11698,N_7560,N_6371);
nor U11699 (N_11699,N_6222,N_6691);
or U11700 (N_11700,N_7313,N_9798);
nor U11701 (N_11701,N_9907,N_6197);
nand U11702 (N_11702,N_7759,N_9549);
and U11703 (N_11703,N_7993,N_8920);
or U11704 (N_11704,N_5318,N_9160);
and U11705 (N_11705,N_7858,N_9386);
and U11706 (N_11706,N_9352,N_8947);
and U11707 (N_11707,N_9512,N_9523);
or U11708 (N_11708,N_7436,N_8895);
nor U11709 (N_11709,N_7197,N_5705);
nand U11710 (N_11710,N_5681,N_5975);
nor U11711 (N_11711,N_5760,N_7846);
and U11712 (N_11712,N_5933,N_8848);
nor U11713 (N_11713,N_6186,N_5153);
xor U11714 (N_11714,N_9673,N_8528);
or U11715 (N_11715,N_5804,N_6809);
nand U11716 (N_11716,N_9846,N_5547);
xor U11717 (N_11717,N_8308,N_6315);
nor U11718 (N_11718,N_9847,N_9613);
xor U11719 (N_11719,N_5808,N_9306);
or U11720 (N_11720,N_8953,N_9506);
or U11721 (N_11721,N_6799,N_6106);
nand U11722 (N_11722,N_9414,N_9719);
or U11723 (N_11723,N_8544,N_7222);
or U11724 (N_11724,N_8413,N_8188);
nor U11725 (N_11725,N_9270,N_7061);
nor U11726 (N_11726,N_6552,N_6221);
nor U11727 (N_11727,N_9191,N_7447);
or U11728 (N_11728,N_7181,N_6098);
nand U11729 (N_11729,N_7445,N_8624);
and U11730 (N_11730,N_7549,N_5737);
xor U11731 (N_11731,N_6620,N_6330);
and U11732 (N_11732,N_6128,N_6443);
nand U11733 (N_11733,N_6110,N_5119);
and U11734 (N_11734,N_6566,N_8778);
and U11735 (N_11735,N_5091,N_7054);
xnor U11736 (N_11736,N_6300,N_5366);
and U11737 (N_11737,N_6860,N_6081);
and U11738 (N_11738,N_6311,N_5470);
nor U11739 (N_11739,N_6094,N_7387);
and U11740 (N_11740,N_7481,N_7394);
xor U11741 (N_11741,N_7057,N_8718);
xnor U11742 (N_11742,N_6785,N_9075);
nor U11743 (N_11743,N_5872,N_6145);
nand U11744 (N_11744,N_5302,N_7432);
or U11745 (N_11745,N_9217,N_6063);
xor U11746 (N_11746,N_5291,N_7584);
xor U11747 (N_11747,N_6652,N_7022);
or U11748 (N_11748,N_6246,N_8492);
xnor U11749 (N_11749,N_7477,N_7332);
xor U11750 (N_11750,N_8905,N_8470);
nor U11751 (N_11751,N_9091,N_8190);
xnor U11752 (N_11752,N_5550,N_9305);
nor U11753 (N_11753,N_7441,N_5848);
nor U11754 (N_11754,N_6182,N_7398);
nand U11755 (N_11755,N_8167,N_6239);
xor U11756 (N_11756,N_6491,N_9426);
or U11757 (N_11757,N_9491,N_8796);
nor U11758 (N_11758,N_6866,N_9567);
and U11759 (N_11759,N_7207,N_6915);
and U11760 (N_11760,N_6998,N_5538);
and U11761 (N_11761,N_5930,N_5894);
and U11762 (N_11762,N_8999,N_5647);
nand U11763 (N_11763,N_5738,N_9708);
and U11764 (N_11764,N_8327,N_5463);
nor U11765 (N_11765,N_7565,N_5920);
nand U11766 (N_11766,N_8942,N_8485);
nand U11767 (N_11767,N_6583,N_7754);
nand U11768 (N_11768,N_8994,N_9436);
xnor U11769 (N_11769,N_6062,N_6499);
and U11770 (N_11770,N_9036,N_6619);
nand U11771 (N_11771,N_9361,N_6822);
xor U11772 (N_11772,N_5063,N_6523);
or U11773 (N_11773,N_8965,N_8384);
or U11774 (N_11774,N_9684,N_5765);
nor U11775 (N_11775,N_6959,N_9344);
xor U11776 (N_11776,N_8149,N_8417);
and U11777 (N_11777,N_8635,N_6422);
nor U11778 (N_11778,N_7607,N_8864);
nand U11779 (N_11779,N_5278,N_6282);
nor U11780 (N_11780,N_7040,N_8563);
xor U11781 (N_11781,N_6818,N_9747);
or U11782 (N_11782,N_9653,N_8706);
xor U11783 (N_11783,N_9292,N_6708);
nor U11784 (N_11784,N_9972,N_9542);
nor U11785 (N_11785,N_8351,N_5094);
nor U11786 (N_11786,N_7505,N_6665);
nor U11787 (N_11787,N_6277,N_8642);
and U11788 (N_11788,N_7704,N_5156);
and U11789 (N_11789,N_5171,N_6046);
nor U11790 (N_11790,N_5148,N_9887);
nand U11791 (N_11791,N_9263,N_5942);
nand U11792 (N_11792,N_9085,N_6192);
and U11793 (N_11793,N_6097,N_5523);
and U11794 (N_11794,N_7741,N_9550);
nand U11795 (N_11795,N_7015,N_6269);
nand U11796 (N_11796,N_6325,N_9391);
nor U11797 (N_11797,N_6676,N_8527);
xnor U11798 (N_11798,N_6334,N_9190);
and U11799 (N_11799,N_9635,N_9179);
nand U11800 (N_11800,N_9811,N_6879);
and U11801 (N_11801,N_7601,N_5185);
xnor U11802 (N_11802,N_7930,N_7439);
nand U11803 (N_11803,N_8639,N_7166);
xnor U11804 (N_11804,N_9189,N_8367);
xor U11805 (N_11805,N_5206,N_7893);
nand U11806 (N_11806,N_6072,N_6721);
and U11807 (N_11807,N_9787,N_9976);
xnor U11808 (N_11808,N_5932,N_7817);
xnor U11809 (N_11809,N_8811,N_6814);
xnor U11810 (N_11810,N_7813,N_9837);
and U11811 (N_11811,N_6233,N_8260);
and U11812 (N_11812,N_5241,N_5124);
and U11813 (N_11813,N_8480,N_8830);
nand U11814 (N_11814,N_9843,N_7904);
nor U11815 (N_11815,N_9836,N_5725);
nor U11816 (N_11816,N_8711,N_8129);
and U11817 (N_11817,N_6028,N_8816);
nand U11818 (N_11818,N_7093,N_5473);
or U11819 (N_11819,N_6032,N_8203);
or U11820 (N_11820,N_5558,N_7835);
xor U11821 (N_11821,N_5305,N_7164);
xnor U11822 (N_11822,N_9956,N_9379);
or U11823 (N_11823,N_5720,N_8312);
and U11824 (N_11824,N_5352,N_8184);
and U11825 (N_11825,N_9256,N_8838);
xor U11826 (N_11826,N_8065,N_9638);
xor U11827 (N_11827,N_5761,N_7422);
nor U11828 (N_11828,N_6017,N_5880);
and U11829 (N_11829,N_5410,N_9393);
xnor U11830 (N_11830,N_6943,N_9909);
nand U11831 (N_11831,N_6425,N_8558);
or U11832 (N_11832,N_9097,N_7569);
nand U11833 (N_11833,N_7026,N_9311);
and U11834 (N_11834,N_9187,N_6467);
and U11835 (N_11835,N_7787,N_5207);
xnor U11836 (N_11836,N_5686,N_5229);
or U11837 (N_11837,N_6432,N_7905);
or U11838 (N_11838,N_6744,N_7687);
nand U11839 (N_11839,N_5700,N_5466);
xor U11840 (N_11840,N_7970,N_7883);
xnor U11841 (N_11841,N_9030,N_6483);
or U11842 (N_11842,N_9561,N_7979);
or U11843 (N_11843,N_9264,N_5923);
nor U11844 (N_11844,N_6995,N_5105);
or U11845 (N_11845,N_7144,N_8857);
nand U11846 (N_11846,N_6730,N_6210);
nor U11847 (N_11847,N_7965,N_8653);
or U11848 (N_11848,N_5638,N_7529);
or U11849 (N_11849,N_9849,N_6241);
or U11850 (N_11850,N_8681,N_7069);
nand U11851 (N_11851,N_6018,N_6776);
xor U11852 (N_11852,N_6258,N_8197);
or U11853 (N_11853,N_8517,N_9710);
and U11854 (N_11854,N_5003,N_9341);
and U11855 (N_11855,N_7609,N_6016);
and U11856 (N_11856,N_6151,N_9815);
xnor U11857 (N_11857,N_8053,N_9870);
nand U11858 (N_11858,N_8281,N_9119);
or U11859 (N_11859,N_8689,N_7066);
nor U11860 (N_11860,N_7769,N_7906);
nor U11861 (N_11861,N_9411,N_5134);
nor U11862 (N_11862,N_9737,N_7179);
or U11863 (N_11863,N_9410,N_8598);
xor U11864 (N_11864,N_6893,N_5818);
nor U11865 (N_11865,N_5121,N_5554);
and U11866 (N_11866,N_6253,N_5068);
nor U11867 (N_11867,N_8244,N_9338);
nand U11868 (N_11868,N_6894,N_6234);
nand U11869 (N_11869,N_6374,N_8029);
or U11870 (N_11870,N_6312,N_6294);
xnor U11871 (N_11871,N_8284,N_9412);
and U11872 (N_11872,N_7544,N_6100);
or U11873 (N_11873,N_5924,N_7131);
nor U11874 (N_11874,N_6339,N_8769);
nand U11875 (N_11875,N_5129,N_8834);
and U11876 (N_11876,N_5401,N_6568);
nand U11877 (N_11877,N_6189,N_8399);
or U11878 (N_11878,N_7750,N_5968);
xnor U11879 (N_11879,N_7379,N_7651);
xnor U11880 (N_11880,N_9252,N_6084);
and U11881 (N_11881,N_5075,N_5198);
or U11882 (N_11882,N_6786,N_7953);
nor U11883 (N_11883,N_7680,N_7645);
xor U11884 (N_11884,N_7881,N_9863);
and U11885 (N_11885,N_5173,N_9911);
nor U11886 (N_11886,N_8306,N_8191);
or U11887 (N_11887,N_6626,N_5767);
nand U11888 (N_11888,N_7342,N_5444);
and U11889 (N_11889,N_7016,N_5437);
and U11890 (N_11890,N_8068,N_9827);
or U11891 (N_11891,N_7747,N_7519);
xor U11892 (N_11892,N_8861,N_6543);
nor U11893 (N_11893,N_6304,N_7891);
nor U11894 (N_11894,N_6933,N_7148);
nor U11895 (N_11895,N_5778,N_5374);
nand U11896 (N_11896,N_7254,N_9328);
nor U11897 (N_11897,N_6008,N_9483);
nand U11898 (N_11898,N_6212,N_8362);
xnor U11899 (N_11899,N_6163,N_9044);
and U11900 (N_11900,N_5988,N_5913);
nand U11901 (N_11901,N_5788,N_8174);
nand U11902 (N_11902,N_8314,N_8845);
or U11903 (N_11903,N_7662,N_6445);
nand U11904 (N_11904,N_5162,N_5183);
nor U11905 (N_11905,N_5602,N_9531);
and U11906 (N_11906,N_9016,N_9720);
nor U11907 (N_11907,N_7633,N_8709);
nor U11908 (N_11908,N_7571,N_6042);
xnor U11909 (N_11909,N_6698,N_8594);
and U11910 (N_11910,N_5500,N_5406);
and U11911 (N_11911,N_6821,N_5035);
nand U11912 (N_11912,N_7142,N_5167);
nor U11913 (N_11913,N_7368,N_8361);
or U11914 (N_11914,N_5047,N_8762);
nand U11915 (N_11915,N_7146,N_7547);
nor U11916 (N_11916,N_7107,N_7360);
xor U11917 (N_11917,N_9675,N_8955);
and U11918 (N_11918,N_8874,N_9451);
xnor U11919 (N_11919,N_7535,N_5018);
xor U11920 (N_11920,N_5633,N_9403);
and U11921 (N_11921,N_9092,N_8520);
or U11922 (N_11922,N_8134,N_5712);
or U11923 (N_11923,N_6162,N_8247);
xnor U11924 (N_11924,N_9568,N_6401);
xor U11925 (N_11925,N_6410,N_6014);
and U11926 (N_11926,N_6022,N_6051);
nand U11927 (N_11927,N_7659,N_9244);
nand U11928 (N_11928,N_7615,N_6538);
xnor U11929 (N_11929,N_6536,N_6275);
or U11930 (N_11930,N_7721,N_8213);
or U11931 (N_11931,N_5462,N_5929);
or U11932 (N_11932,N_9593,N_9598);
or U11933 (N_11933,N_6158,N_6666);
or U11934 (N_11934,N_7229,N_7334);
nand U11935 (N_11935,N_5938,N_8881);
and U11936 (N_11936,N_7563,N_5285);
nand U11937 (N_11937,N_7133,N_9627);
and U11938 (N_11938,N_9122,N_5522);
xor U11939 (N_11939,N_6709,N_7802);
nor U11940 (N_11940,N_8251,N_7806);
or U11941 (N_11941,N_5104,N_6524);
or U11942 (N_11942,N_8646,N_7783);
xnor U11943 (N_11943,N_7745,N_5881);
nand U11944 (N_11944,N_6804,N_6360);
nand U11945 (N_11945,N_5073,N_5847);
xor U11946 (N_11946,N_9758,N_6891);
nand U11947 (N_11947,N_7623,N_8181);
xnor U11948 (N_11948,N_7917,N_5772);
nand U11949 (N_11949,N_6474,N_8562);
and U11950 (N_11950,N_9573,N_9255);
xor U11951 (N_11951,N_7602,N_7743);
xor U11952 (N_11952,N_7331,N_7537);
nor U11953 (N_11953,N_7497,N_7111);
nor U11954 (N_11954,N_7196,N_7064);
nand U11955 (N_11955,N_5965,N_6123);
nand U11956 (N_11956,N_8702,N_6205);
or U11957 (N_11957,N_9805,N_6722);
nor U11958 (N_11958,N_8846,N_6291);
or U11959 (N_11959,N_5673,N_7463);
and U11960 (N_11960,N_5308,N_7546);
nor U11961 (N_11961,N_6272,N_6352);
nand U11962 (N_11962,N_8460,N_7826);
nand U11963 (N_11963,N_6209,N_9964);
or U11964 (N_11964,N_6257,N_6264);
and U11965 (N_11965,N_7768,N_9456);
xor U11966 (N_11966,N_7399,N_5667);
nand U11967 (N_11967,N_9564,N_7005);
nor U11968 (N_11968,N_6177,N_9558);
and U11969 (N_11969,N_7963,N_6490);
and U11970 (N_11970,N_7336,N_6752);
or U11971 (N_11971,N_9124,N_9602);
nor U11972 (N_11972,N_9002,N_8532);
nor U11973 (N_11973,N_9934,N_5427);
xnor U11974 (N_11974,N_8060,N_8843);
xor U11975 (N_11975,N_5037,N_5086);
nand U11976 (N_11976,N_5580,N_5076);
or U11977 (N_11977,N_5863,N_8772);
nand U11978 (N_11978,N_9858,N_8967);
or U11979 (N_11979,N_6465,N_9854);
nor U11980 (N_11980,N_8832,N_7888);
xor U11981 (N_11981,N_9671,N_9444);
xor U11982 (N_11982,N_7666,N_7707);
nor U11983 (N_11983,N_6564,N_9438);
or U11984 (N_11984,N_7444,N_9873);
xor U11985 (N_11985,N_9291,N_5024);
nor U11986 (N_11986,N_5253,N_6680);
xnor U11987 (N_11987,N_7099,N_8025);
or U11988 (N_11988,N_9322,N_5276);
nor U11989 (N_11989,N_8819,N_7898);
xnor U11990 (N_11990,N_8829,N_8866);
xnor U11991 (N_11991,N_7838,N_6207);
or U11992 (N_11992,N_6655,N_9178);
nand U11993 (N_11993,N_7359,N_5658);
and U11994 (N_11994,N_6961,N_5422);
xor U11995 (N_11995,N_7195,N_7643);
xnor U11996 (N_11996,N_8116,N_8287);
nand U11997 (N_11997,N_8515,N_7233);
and U11998 (N_11998,N_5050,N_7811);
xnor U11999 (N_11999,N_9103,N_7892);
xor U12000 (N_12000,N_7793,N_6353);
nand U12001 (N_12001,N_5535,N_5501);
or U12002 (N_12002,N_8597,N_6542);
xnor U12003 (N_12003,N_9728,N_5290);
and U12004 (N_12004,N_9835,N_8707);
xnor U12005 (N_12005,N_6658,N_8171);
or U12006 (N_12006,N_7012,N_7009);
nand U12007 (N_12007,N_7945,N_7815);
nor U12008 (N_12008,N_7613,N_5014);
and U12009 (N_12009,N_6424,N_8289);
and U12010 (N_12010,N_6248,N_7850);
xnor U12011 (N_12011,N_8692,N_5957);
or U12012 (N_12012,N_6842,N_9908);
or U12013 (N_12013,N_6737,N_9622);
nand U12014 (N_12014,N_5582,N_6993);
or U12015 (N_12015,N_9586,N_9608);
nor U12016 (N_12016,N_5812,N_6274);
nor U12017 (N_12017,N_9151,N_8764);
and U12018 (N_12018,N_8737,N_5755);
nand U12019 (N_12019,N_5722,N_6875);
nand U12020 (N_12020,N_6125,N_5498);
nor U12021 (N_12021,N_6290,N_8064);
nor U12022 (N_12022,N_7376,N_9165);
nor U12023 (N_12023,N_8824,N_6179);
nand U12024 (N_12024,N_9923,N_7087);
and U12025 (N_12025,N_9691,N_7870);
and U12026 (N_12026,N_7836,N_9090);
and U12027 (N_12027,N_6671,N_5384);
xor U12028 (N_12028,N_7381,N_7720);
nor U12029 (N_12029,N_7809,N_5931);
and U12030 (N_12030,N_9670,N_5505);
nand U12031 (N_12031,N_8124,N_6798);
nand U12032 (N_12032,N_8237,N_7711);
nand U12033 (N_12033,N_6574,N_6585);
xor U12034 (N_12034,N_5605,N_5542);
nor U12035 (N_12035,N_9280,N_8238);
and U12036 (N_12036,N_7746,N_6718);
or U12037 (N_12037,N_5343,N_7159);
nor U12038 (N_12038,N_8998,N_9974);
xnor U12039 (N_12039,N_9072,N_8096);
xor U12040 (N_12040,N_6227,N_6036);
nand U12041 (N_12041,N_9374,N_5560);
and U12042 (N_12042,N_9888,N_9142);
nand U12043 (N_12043,N_9741,N_5330);
nor U12044 (N_12044,N_9201,N_8670);
xnor U12045 (N_12045,N_5612,N_5911);
nor U12046 (N_12046,N_6495,N_6284);
or U12047 (N_12047,N_6142,N_8356);
nand U12048 (N_12048,N_6855,N_7454);
and U12049 (N_12049,N_6612,N_5521);
or U12050 (N_12050,N_6768,N_7600);
or U12051 (N_12051,N_6101,N_6572);
xnor U12052 (N_12052,N_7255,N_7075);
nor U12053 (N_12053,N_8889,N_8523);
xnor U12054 (N_12054,N_9174,N_9029);
or U12055 (N_12055,N_5821,N_6590);
nor U12056 (N_12056,N_5716,N_5524);
and U12057 (N_12057,N_6076,N_9597);
nand U12058 (N_12058,N_9626,N_7032);
nor U12059 (N_12059,N_9697,N_5824);
nor U12060 (N_12060,N_9200,N_5747);
nand U12061 (N_12061,N_8836,N_6030);
nand U12062 (N_12062,N_8710,N_5709);
nand U12063 (N_12063,N_9810,N_7045);
xnor U12064 (N_12064,N_5888,N_9844);
or U12065 (N_12065,N_7303,N_5710);
nor U12066 (N_12066,N_6302,N_8381);
nor U12067 (N_12067,N_9871,N_5288);
nand U12068 (N_12068,N_9705,N_5102);
nand U12069 (N_12069,N_7328,N_7960);
or U12070 (N_12070,N_7118,N_7461);
nand U12071 (N_12071,N_6041,N_6819);
or U12072 (N_12072,N_5744,N_7013);
or U12073 (N_12073,N_8993,N_6492);
or U12074 (N_12074,N_5508,N_7935);
nand U12075 (N_12075,N_6904,N_9503);
or U12076 (N_12076,N_5431,N_8043);
xnor U12077 (N_12077,N_5120,N_7038);
and U12078 (N_12078,N_8369,N_5060);
and U12079 (N_12079,N_7955,N_7644);
nor U12080 (N_12080,N_7415,N_6973);
nand U12081 (N_12081,N_6976,N_6308);
and U12082 (N_12082,N_6266,N_8799);
nand U12083 (N_12083,N_8756,N_9625);
xor U12084 (N_12084,N_5879,N_5637);
nor U12085 (N_12085,N_9681,N_5295);
or U12086 (N_12086,N_9032,N_7621);
and U12087 (N_12087,N_7484,N_8051);
xnor U12088 (N_12088,N_8826,N_7172);
nand U12089 (N_12089,N_7843,N_8922);
and U12090 (N_12090,N_8353,N_5713);
xor U12091 (N_12091,N_5639,N_6911);
and U12092 (N_12092,N_9897,N_9113);
or U12093 (N_12093,N_6941,N_6704);
xnor U12094 (N_12094,N_6055,N_6584);
and U12095 (N_12095,N_5403,N_8860);
xor U12096 (N_12096,N_7214,N_6433);
nor U12097 (N_12097,N_5734,N_6717);
nor U12098 (N_12098,N_7948,N_8273);
and U12099 (N_12099,N_8641,N_9992);
nand U12100 (N_12100,N_6479,N_5192);
and U12101 (N_12101,N_7083,N_8665);
or U12102 (N_12102,N_8831,N_7237);
and U12103 (N_12103,N_5935,N_5843);
or U12104 (N_12104,N_5259,N_7517);
or U12105 (N_12105,N_7033,N_5620);
nand U12106 (N_12106,N_6083,N_5604);
xnor U12107 (N_12107,N_7918,N_8663);
xnor U12108 (N_12108,N_5097,N_5727);
nor U12109 (N_12109,N_5783,N_8037);
or U12110 (N_12110,N_5188,N_9315);
or U12111 (N_12111,N_5136,N_6978);
or U12112 (N_12112,N_5095,N_6594);
and U12113 (N_12113,N_5578,N_5785);
and U12114 (N_12114,N_7101,N_5534);
nand U12115 (N_12115,N_8404,N_8254);
nor U12116 (N_12116,N_8564,N_6711);
and U12117 (N_12117,N_9295,N_9687);
nand U12118 (N_12118,N_8424,N_9885);
nand U12119 (N_12119,N_6071,N_8887);
or U12120 (N_12120,N_8671,N_9677);
nor U12121 (N_12121,N_9435,N_6644);
xnor U12122 (N_12122,N_7775,N_6385);
nor U12123 (N_12123,N_9442,N_6849);
nand U12124 (N_12124,N_9667,N_6006);
and U12125 (N_12125,N_9772,N_7431);
xor U12126 (N_12126,N_6126,N_5540);
nor U12127 (N_12127,N_9259,N_8193);
or U12128 (N_12128,N_6997,N_9167);
nand U12129 (N_12129,N_9928,N_9134);
xnor U12130 (N_12130,N_7234,N_8493);
nor U12131 (N_12131,N_9332,N_7841);
nand U12132 (N_12132,N_8655,N_5034);
or U12133 (N_12133,N_5839,N_6710);
nor U12134 (N_12134,N_5373,N_7485);
or U12135 (N_12135,N_5714,N_9712);
and U12136 (N_12136,N_6813,N_7465);
nor U12137 (N_12137,N_7260,N_5346);
or U12138 (N_12138,N_7350,N_6124);
nor U12139 (N_12139,N_8411,N_5013);
xor U12140 (N_12140,N_9826,N_5382);
xnor U12141 (N_12141,N_8239,N_6393);
nand U12142 (N_12142,N_9114,N_9026);
nand U12143 (N_12143,N_5656,N_8878);
nor U12144 (N_12144,N_5607,N_6899);
xnor U12145 (N_12145,N_8550,N_6602);
or U12146 (N_12146,N_5614,N_7494);
nor U12147 (N_12147,N_8957,N_5347);
xnor U12148 (N_12148,N_6545,N_6468);
nand U12149 (N_12149,N_9883,N_8790);
or U12150 (N_12150,N_5048,N_9228);
xor U12151 (N_12151,N_9146,N_9778);
nor U12152 (N_12152,N_6840,N_6635);
xnor U12153 (N_12153,N_8331,N_6932);
and U12154 (N_12154,N_7103,N_9768);
nor U12155 (N_12155,N_6745,N_7128);
or U12156 (N_12156,N_5193,N_5976);
or U12157 (N_12157,N_5779,N_6960);
and U12158 (N_12158,N_8996,N_5269);
nand U12159 (N_12159,N_8100,N_7048);
xnor U12160 (N_12160,N_7967,N_5509);
and U12161 (N_12161,N_7309,N_5723);
nor U12162 (N_12162,N_5367,N_9663);
xor U12163 (N_12163,N_8121,N_8962);
xnor U12164 (N_12164,N_6449,N_5515);
or U12165 (N_12165,N_9326,N_8770);
and U12166 (N_12166,N_5279,N_8919);
nand U12167 (N_12167,N_8656,N_9494);
or U12168 (N_12168,N_5544,N_8026);
nand U12169 (N_12169,N_8700,N_9135);
nand U12170 (N_12170,N_9528,N_5974);
and U12171 (N_12171,N_9355,N_5041);
xnor U12172 (N_12172,N_8373,N_5908);
nor U12173 (N_12173,N_9061,N_5152);
nor U12174 (N_12174,N_7576,N_9895);
nand U12175 (N_12175,N_5759,N_9899);
or U12176 (N_12176,N_6541,N_6629);
and U12177 (N_12177,N_9996,N_9563);
xnor U12178 (N_12178,N_7710,N_9253);
xnor U12179 (N_12179,N_9685,N_8959);
or U12180 (N_12180,N_8246,N_8168);
xnor U12181 (N_12181,N_5031,N_5870);
nor U12182 (N_12182,N_6020,N_5669);
xnor U12183 (N_12183,N_5474,N_6283);
and U12184 (N_12184,N_6344,N_8632);
nand U12185 (N_12185,N_5441,N_6519);
xor U12186 (N_12186,N_6640,N_8945);
xor U12187 (N_12187,N_6697,N_9978);
or U12188 (N_12188,N_7816,N_7539);
xor U12189 (N_12189,N_5693,N_7749);
nor U12190 (N_12190,N_8364,N_5426);
nor U12191 (N_12191,N_6069,N_8044);
xor U12192 (N_12192,N_8258,N_9950);
xnor U12193 (N_12193,N_7688,N_5081);
and U12194 (N_12194,N_5258,N_9553);
and U12195 (N_12195,N_9376,N_6576);
xnor U12196 (N_12196,N_7507,N_9170);
xor U12197 (N_12197,N_8916,N_9164);
and U12198 (N_12198,N_7482,N_6631);
xnor U12199 (N_12199,N_7983,N_8970);
and U12200 (N_12200,N_8003,N_5947);
or U12201 (N_12201,N_5989,N_9665);
or U12202 (N_12202,N_8602,N_9695);
nor U12203 (N_12203,N_9642,N_6686);
nor U12204 (N_12204,N_7282,N_7630);
and U12205 (N_12205,N_7283,N_9698);
nor U12206 (N_12206,N_6148,N_5618);
xor U12207 (N_12207,N_7475,N_8650);
or U12208 (N_12208,N_6194,N_7733);
and U12209 (N_12209,N_8055,N_6525);
nand U12210 (N_12210,N_7186,N_5922);
and U12211 (N_12211,N_6731,N_7165);
nand U12212 (N_12212,N_9337,N_6902);
xnor U12213 (N_12213,N_7305,N_5386);
and U12214 (N_12214,N_8252,N_5096);
and U12215 (N_12215,N_6438,N_6783);
nand U12216 (N_12216,N_7834,N_9390);
and U12217 (N_12217,N_9331,N_5484);
or U12218 (N_12218,N_8825,N_5393);
nand U12219 (N_12219,N_9800,N_6851);
nand U12220 (N_12220,N_5434,N_5416);
or U12221 (N_12221,N_8310,N_5912);
and U12222 (N_12222,N_8151,N_6247);
nor U12223 (N_12223,N_9744,N_9546);
xnor U12224 (N_12224,N_9688,N_9812);
and U12225 (N_12225,N_7338,N_8402);
xor U12226 (N_12226,N_6171,N_9615);
or U12227 (N_12227,N_5910,N_8592);
nand U12228 (N_12228,N_8623,N_8256);
nand U12229 (N_12229,N_6305,N_8585);
and U12230 (N_12230,N_5972,N_9357);
nand U12231 (N_12231,N_6285,N_8668);
nand U12232 (N_12232,N_5624,N_7878);
nor U12233 (N_12233,N_9003,N_9848);
nand U12234 (N_12234,N_8741,N_7155);
and U12235 (N_12235,N_8013,N_6527);
or U12236 (N_12236,N_5814,N_9094);
and U12237 (N_12237,N_7271,N_8509);
and U12238 (N_12238,N_5539,N_7634);
or U12239 (N_12239,N_9991,N_7550);
nor U12240 (N_12240,N_8658,N_7476);
nor U12241 (N_12241,N_9639,N_6927);
or U12242 (N_12242,N_5301,N_7344);
and U12243 (N_12243,N_7437,N_5100);
xnor U12244 (N_12244,N_8036,N_7900);
nor U12245 (N_12245,N_6637,N_6362);
nor U12246 (N_12246,N_5179,N_6567);
nand U12247 (N_12247,N_5840,N_8226);
or U12248 (N_12248,N_6848,N_6999);
nor U12249 (N_12249,N_8683,N_8275);
and U12250 (N_12250,N_6914,N_8455);
or U12251 (N_12251,N_5246,N_8991);
xnor U12252 (N_12252,N_5495,N_5799);
nor U12253 (N_12253,N_6589,N_7104);
nand U12254 (N_12254,N_9944,N_9055);
nand U12255 (N_12255,N_9961,N_9620);
nor U12256 (N_12256,N_8677,N_9447);
nand U12257 (N_12257,N_5154,N_9308);
xnor U12258 (N_12258,N_7543,N_7642);
or U12259 (N_12259,N_7067,N_8782);
or U12260 (N_12260,N_6116,N_8792);
or U12261 (N_12261,N_8018,N_9785);
nor U12262 (N_12262,N_9482,N_6881);
nand U12263 (N_12263,N_6188,N_9202);
nor U12264 (N_12264,N_8742,N_8423);
and U12265 (N_12265,N_6238,N_6732);
nor U12266 (N_12266,N_7065,N_8001);
nor U12267 (N_12267,N_8660,N_9093);
and U12268 (N_12268,N_8283,N_7884);
and U12269 (N_12269,N_8195,N_9416);
nand U12270 (N_12270,N_6102,N_7500);
nor U12271 (N_12271,N_5504,N_9283);
xnor U12272 (N_12272,N_9053,N_6270);
or U12273 (N_12273,N_8412,N_5826);
nor U12274 (N_12274,N_8332,N_6948);
and U12275 (N_12275,N_6833,N_8949);
and U12276 (N_12276,N_8118,N_6466);
nand U12277 (N_12277,N_7223,N_5298);
or U12278 (N_12278,N_9963,N_7974);
nor U12279 (N_12279,N_6889,N_9446);
xnor U12280 (N_12280,N_7701,N_9294);
and U12281 (N_12281,N_6324,N_9794);
and U12282 (N_12282,N_7996,N_5182);
nand U12283 (N_12283,N_7175,N_5178);
and U12284 (N_12284,N_6968,N_8032);
nor U12285 (N_12285,N_5216,N_8293);
or U12286 (N_12286,N_8688,N_5750);
xnor U12287 (N_12287,N_7269,N_5945);
or U12288 (N_12288,N_7840,N_7119);
and U12289 (N_12289,N_7098,N_8218);
xnor U12290 (N_12290,N_7819,N_7678);
and U12291 (N_12291,N_9394,N_6702);
xor U12292 (N_12292,N_8786,N_8318);
nor U12293 (N_12293,N_9490,N_8393);
nor U12294 (N_12294,N_5020,N_7091);
nand U12295 (N_12295,N_5413,N_6172);
xor U12296 (N_12296,N_7681,N_7182);
or U12297 (N_12297,N_6319,N_6753);
and U12298 (N_12298,N_8697,N_8139);
and U12299 (N_12299,N_7285,N_8723);
nand U12300 (N_12300,N_5370,N_7329);
and U12301 (N_12301,N_8744,N_5928);
xor U12302 (N_12302,N_9237,N_7610);
and U12303 (N_12303,N_6505,N_6035);
nand U12304 (N_12304,N_5643,N_7319);
xor U12305 (N_12305,N_7291,N_9816);
and U12306 (N_12306,N_9222,N_8648);
or U12307 (N_12307,N_9912,N_6436);
or U12308 (N_12308,N_9459,N_8122);
and U12309 (N_12309,N_6957,N_8313);
nand U12310 (N_12310,N_9246,N_8803);
or U12311 (N_12311,N_5491,N_7837);
nor U12312 (N_12312,N_5467,N_9515);
nor U12313 (N_12313,N_5903,N_5482);
nor U12314 (N_12314,N_6649,N_9637);
nand U12315 (N_12315,N_5394,N_9018);
or U12316 (N_12316,N_5471,N_7871);
nor U12317 (N_12317,N_7726,N_5130);
xor U12318 (N_12318,N_6624,N_8035);
nand U12319 (N_12319,N_7975,N_7592);
xnor U12320 (N_12320,N_5627,N_8654);
xnor U12321 (N_12321,N_5435,N_9524);
or U12322 (N_12322,N_5460,N_5649);
and U12323 (N_12323,N_9935,N_8484);
xnor U12324 (N_12324,N_9370,N_6185);
and U12325 (N_12325,N_5867,N_7845);
nor U12326 (N_12326,N_9203,N_7149);
nand U12327 (N_12327,N_7346,N_9488);
nand U12328 (N_12328,N_8084,N_7252);
and U12329 (N_12329,N_8573,N_5494);
nand U12330 (N_12330,N_9917,N_6864);
and U12331 (N_12331,N_9654,N_5045);
nor U12332 (N_12332,N_7782,N_7512);
xnor U12333 (N_12333,N_7413,N_8365);
xnor U12334 (N_12334,N_7275,N_5937);
nor U12335 (N_12335,N_7804,N_5064);
nor U12336 (N_12336,N_5619,N_9580);
nor U12337 (N_12337,N_9221,N_9472);
and U12338 (N_12338,N_9727,N_8020);
nor U12339 (N_12339,N_8712,N_7593);
or U12340 (N_12340,N_9163,N_8478);
and U12341 (N_12341,N_9521,N_5365);
nand U12342 (N_12342,N_8621,N_9245);
or U12343 (N_12343,N_9108,N_9240);
nor U12344 (N_12344,N_6824,N_5827);
nor U12345 (N_12345,N_9353,N_6618);
xor U12346 (N_12346,N_7216,N_5640);
and U12347 (N_12347,N_8119,N_7374);
nor U12348 (N_12348,N_5936,N_8169);
xnor U12349 (N_12349,N_6869,N_5480);
nor U12350 (N_12350,N_8349,N_8131);
xnor U12351 (N_12351,N_7694,N_5376);
xor U12352 (N_12352,N_7691,N_7221);
or U12353 (N_12353,N_7525,N_8835);
nand U12354 (N_12354,N_7297,N_7217);
nor U12355 (N_12355,N_8806,N_8266);
and U12356 (N_12356,N_9958,N_9006);
or U12357 (N_12357,N_7616,N_6391);
nand U12358 (N_12358,N_5230,N_5356);
nand U12359 (N_12359,N_9158,N_5062);
and U12360 (N_12360,N_5002,N_6388);
nand U12361 (N_12361,N_5532,N_5628);
nand U12362 (N_12362,N_7818,N_5529);
and U12363 (N_12363,N_5428,N_8852);
or U12364 (N_12364,N_6989,N_6195);
or U12365 (N_12365,N_9683,N_6908);
and U12366 (N_12366,N_6750,N_7924);
nand U12367 (N_12367,N_5009,N_9397);
xor U12368 (N_12368,N_7203,N_8099);
nor U12369 (N_12369,N_5708,N_7899);
xor U12370 (N_12370,N_5587,N_5055);
nor U12371 (N_12371,N_6606,N_9293);
nor U12372 (N_12372,N_8110,N_9421);
nor U12373 (N_12373,N_8107,N_5059);
nor U12374 (N_12374,N_9879,N_6580);
nand U12375 (N_12375,N_6206,N_7874);
or U12376 (N_12376,N_5692,N_8647);
and U12377 (N_12377,N_5362,N_5707);
xnor U12378 (N_12378,N_5569,N_7639);
or U12379 (N_12379,N_8757,N_5451);
and U12380 (N_12380,N_6861,N_6060);
or U12381 (N_12381,N_9473,N_7209);
and U12382 (N_12382,N_5565,N_9692);
xor U12383 (N_12383,N_9105,N_5666);
and U12384 (N_12384,N_5281,N_5553);
xnor U12385 (N_12385,N_5381,N_7266);
nand U12386 (N_12386,N_9373,N_7327);
or U12387 (N_12387,N_6788,N_6378);
nand U12388 (N_12388,N_5454,N_5635);
or U12389 (N_12389,N_8108,N_6176);
xor U12390 (N_12390,N_5450,N_5939);
nand U12391 (N_12391,N_7925,N_9922);
and U12392 (N_12392,N_6969,N_7848);
and U12393 (N_12393,N_7751,N_5520);
and U12394 (N_12394,N_7440,N_6131);
nand U12395 (N_12395,N_8472,N_5856);
and U12396 (N_12396,N_8569,N_7110);
nor U12397 (N_12397,N_7357,N_6326);
xor U12398 (N_12398,N_8751,N_9132);
nor U12399 (N_12399,N_5316,N_5695);
nand U12400 (N_12400,N_7725,N_9004);
or U12401 (N_12401,N_6843,N_6887);
nor U12402 (N_12402,N_8229,N_8840);
xnor U12403 (N_12403,N_8699,N_9017);
or U12404 (N_12404,N_8733,N_7604);
and U12405 (N_12405,N_5690,N_5918);
or U12406 (N_12406,N_8912,N_8694);
or U12407 (N_12407,N_9238,N_5270);
nor U12408 (N_12408,N_5128,N_7100);
nor U12409 (N_12409,N_9662,N_6681);
nand U12410 (N_12410,N_9903,N_9346);
xnor U12411 (N_12411,N_9997,N_9788);
nor U12412 (N_12412,N_7646,N_7739);
nor U12413 (N_12413,N_9970,N_5417);
and U12414 (N_12414,N_6956,N_9282);
and U12415 (N_12415,N_9693,N_5388);
xnor U12416 (N_12416,N_5771,N_5247);
or U12417 (N_12417,N_6120,N_8302);
nand U12418 (N_12418,N_9973,N_8904);
nor U12419 (N_12419,N_5303,N_6569);
xnor U12420 (N_12420,N_7929,N_8041);
or U12421 (N_12421,N_7467,N_6549);
nor U12422 (N_12422,N_7448,N_7829);
nor U12423 (N_12423,N_8735,N_5357);
and U12424 (N_12424,N_6187,N_5329);
nand U12425 (N_12425,N_9509,N_8183);
and U12426 (N_12426,N_5549,N_6373);
xnor U12427 (N_12427,N_8784,N_7017);
nor U12428 (N_12428,N_5746,N_5369);
and U12429 (N_12429,N_7170,N_7736);
xnor U12430 (N_12430,N_8719,N_7950);
or U12431 (N_12431,N_9557,N_9599);
xor U12432 (N_12432,N_8461,N_9211);
and U12433 (N_12433,N_9544,N_9896);
and U12434 (N_12434,N_9335,N_8236);
nor U12435 (N_12435,N_9123,N_8448);
xnor U12436 (N_12436,N_6501,N_8763);
nor U12437 (N_12437,N_7502,N_6498);
nand U12438 (N_12438,N_9872,N_9102);
or U12439 (N_12439,N_5296,N_5646);
or U12440 (N_12440,N_9485,N_6477);
and U12441 (N_12441,N_6913,N_6356);
nand U12442 (N_12442,N_6805,N_5577);
nor U12443 (N_12443,N_5012,N_7722);
nor U12444 (N_12444,N_7121,N_9760);
nand U12445 (N_12445,N_6794,N_9195);
nor U12446 (N_12446,N_8326,N_8422);
nand U12447 (N_12447,N_7914,N_6636);
nor U12448 (N_12448,N_6835,N_7962);
xor U12449 (N_12449,N_9869,N_5353);
xnor U12450 (N_12450,N_6243,N_5834);
and U12451 (N_12451,N_8352,N_8128);
xnor U12452 (N_12452,N_7503,N_6218);
nor U12453 (N_12453,N_8042,N_8279);
nor U12454 (N_12454,N_5213,N_5668);
and U12455 (N_12455,N_6674,N_8818);
xnor U12456 (N_12456,N_9786,N_6963);
nand U12457 (N_12457,N_8721,N_9845);
nor U12458 (N_12458,N_9038,N_6570);
nand U12459 (N_12459,N_9258,N_5683);
or U12460 (N_12460,N_9901,N_5320);
nor U12461 (N_12461,N_6925,N_8017);
or U12462 (N_12462,N_7928,N_8731);
nor U12463 (N_12463,N_9303,N_8391);
nor U12464 (N_12464,N_8086,N_5275);
or U12465 (N_12465,N_5203,N_5143);
nor U12466 (N_12466,N_5803,N_5122);
xor U12467 (N_12467,N_5093,N_9656);
and U12468 (N_12468,N_8863,N_7853);
xnor U12469 (N_12469,N_8132,N_8743);
nor U12470 (N_12470,N_8010,N_8603);
nand U12471 (N_12471,N_9307,N_5146);
nor U12472 (N_12472,N_8559,N_6107);
or U12473 (N_12473,N_8858,N_8375);
or U12474 (N_12474,N_8127,N_9034);
and U12475 (N_12475,N_5996,N_8696);
nor U12476 (N_12476,N_5137,N_7579);
nand U12477 (N_12477,N_8516,N_9861);
nand U12478 (N_12478,N_8458,N_8759);
xnor U12479 (N_12479,N_7185,N_5568);
and U12480 (N_12480,N_5396,N_5701);
nor U12481 (N_12481,N_9689,N_6669);
or U12482 (N_12482,N_7895,N_7969);
or U12483 (N_12483,N_9173,N_5397);
and U12484 (N_12484,N_7761,N_9781);
or U12485 (N_12485,N_8908,N_9790);
nor U12486 (N_12486,N_5857,N_6930);
xnor U12487 (N_12487,N_5333,N_9590);
and U12488 (N_12488,N_8570,N_5227);
nand U12489 (N_12489,N_5195,N_9343);
nor U12490 (N_12490,N_9578,N_9877);
xnor U12491 (N_12491,N_6781,N_8975);
or U12492 (N_12492,N_7763,N_7943);
nand U12493 (N_12493,N_7105,N_8355);
xnor U12494 (N_12494,N_7373,N_6299);
nor U12495 (N_12495,N_6486,N_8027);
nor U12496 (N_12496,N_5468,N_6758);
xor U12497 (N_12497,N_5898,N_9172);
nand U12498 (N_12498,N_8910,N_8490);
nand U12499 (N_12499,N_6066,N_9510);
and U12500 (N_12500,N_9533,N_9519);
xnor U12501 (N_12501,N_5281,N_8381);
or U12502 (N_12502,N_5495,N_9840);
or U12503 (N_12503,N_6567,N_9219);
and U12504 (N_12504,N_8157,N_5154);
and U12505 (N_12505,N_6765,N_8698);
xnor U12506 (N_12506,N_5180,N_7276);
xor U12507 (N_12507,N_8022,N_7377);
or U12508 (N_12508,N_5504,N_8801);
nand U12509 (N_12509,N_5263,N_9195);
and U12510 (N_12510,N_7918,N_9889);
xnor U12511 (N_12511,N_8305,N_7188);
or U12512 (N_12512,N_5587,N_5935);
and U12513 (N_12513,N_8914,N_9809);
and U12514 (N_12514,N_8495,N_7286);
and U12515 (N_12515,N_7364,N_6638);
or U12516 (N_12516,N_8571,N_8761);
or U12517 (N_12517,N_7279,N_6361);
nor U12518 (N_12518,N_7700,N_7838);
nand U12519 (N_12519,N_8736,N_5604);
or U12520 (N_12520,N_6709,N_5964);
xor U12521 (N_12521,N_7499,N_8019);
nand U12522 (N_12522,N_5476,N_8499);
xor U12523 (N_12523,N_5635,N_8286);
nor U12524 (N_12524,N_9304,N_9640);
or U12525 (N_12525,N_6409,N_8993);
xor U12526 (N_12526,N_5051,N_6351);
and U12527 (N_12527,N_9007,N_7803);
or U12528 (N_12528,N_6833,N_9446);
or U12529 (N_12529,N_6374,N_8415);
nand U12530 (N_12530,N_9545,N_7660);
nor U12531 (N_12531,N_5708,N_8537);
and U12532 (N_12532,N_7685,N_5642);
xnor U12533 (N_12533,N_8094,N_5147);
nor U12534 (N_12534,N_8048,N_5818);
nor U12535 (N_12535,N_9455,N_9354);
or U12536 (N_12536,N_8012,N_8341);
or U12537 (N_12537,N_7983,N_7736);
nand U12538 (N_12538,N_9576,N_7994);
and U12539 (N_12539,N_7183,N_9070);
nand U12540 (N_12540,N_8391,N_6299);
nor U12541 (N_12541,N_8654,N_5526);
nand U12542 (N_12542,N_8833,N_7791);
and U12543 (N_12543,N_6902,N_9909);
nand U12544 (N_12544,N_6343,N_6587);
nor U12545 (N_12545,N_9795,N_8215);
nor U12546 (N_12546,N_7210,N_5618);
or U12547 (N_12547,N_5609,N_5905);
or U12548 (N_12548,N_7960,N_5778);
and U12549 (N_12549,N_5231,N_8642);
nand U12550 (N_12550,N_6074,N_7062);
or U12551 (N_12551,N_8150,N_6899);
and U12552 (N_12552,N_8050,N_9970);
nand U12553 (N_12553,N_5421,N_9603);
xnor U12554 (N_12554,N_7500,N_8018);
nand U12555 (N_12555,N_5283,N_7830);
nor U12556 (N_12556,N_8230,N_6123);
or U12557 (N_12557,N_7256,N_8329);
or U12558 (N_12558,N_9354,N_5403);
nand U12559 (N_12559,N_6090,N_6023);
or U12560 (N_12560,N_6424,N_5958);
nor U12561 (N_12561,N_5122,N_8212);
nor U12562 (N_12562,N_8837,N_6348);
and U12563 (N_12563,N_5667,N_7560);
and U12564 (N_12564,N_6740,N_9503);
nor U12565 (N_12565,N_6751,N_9269);
and U12566 (N_12566,N_7258,N_6698);
xnor U12567 (N_12567,N_8731,N_6908);
or U12568 (N_12568,N_9822,N_6874);
nand U12569 (N_12569,N_8425,N_9589);
or U12570 (N_12570,N_6449,N_5935);
nand U12571 (N_12571,N_7649,N_7093);
nor U12572 (N_12572,N_8852,N_5192);
nor U12573 (N_12573,N_8037,N_9891);
nand U12574 (N_12574,N_6295,N_7425);
nand U12575 (N_12575,N_8113,N_5620);
nor U12576 (N_12576,N_5614,N_5847);
and U12577 (N_12577,N_5812,N_8802);
nor U12578 (N_12578,N_7701,N_9488);
and U12579 (N_12579,N_7008,N_6867);
or U12580 (N_12580,N_5689,N_7828);
xnor U12581 (N_12581,N_7868,N_5035);
xnor U12582 (N_12582,N_9632,N_9455);
nand U12583 (N_12583,N_9598,N_9185);
xnor U12584 (N_12584,N_9566,N_9249);
xor U12585 (N_12585,N_6314,N_7183);
xnor U12586 (N_12586,N_8781,N_9482);
xor U12587 (N_12587,N_6675,N_8679);
nand U12588 (N_12588,N_6730,N_8470);
or U12589 (N_12589,N_6276,N_7416);
and U12590 (N_12590,N_9587,N_5565);
and U12591 (N_12591,N_5921,N_6113);
nand U12592 (N_12592,N_6702,N_5741);
or U12593 (N_12593,N_5475,N_7836);
xnor U12594 (N_12594,N_6619,N_8541);
xor U12595 (N_12595,N_8075,N_7911);
or U12596 (N_12596,N_7375,N_9858);
nor U12597 (N_12597,N_8048,N_7247);
nand U12598 (N_12598,N_9360,N_7619);
nor U12599 (N_12599,N_9109,N_8397);
xor U12600 (N_12600,N_5774,N_6870);
or U12601 (N_12601,N_5233,N_5497);
xor U12602 (N_12602,N_8271,N_9597);
or U12603 (N_12603,N_8609,N_9372);
and U12604 (N_12604,N_6590,N_7261);
and U12605 (N_12605,N_7886,N_7402);
xnor U12606 (N_12606,N_6124,N_8421);
xnor U12607 (N_12607,N_6708,N_8193);
or U12608 (N_12608,N_9250,N_9596);
nor U12609 (N_12609,N_5289,N_5936);
xnor U12610 (N_12610,N_5397,N_9708);
xor U12611 (N_12611,N_8290,N_9866);
or U12612 (N_12612,N_6946,N_8085);
and U12613 (N_12613,N_9117,N_8328);
or U12614 (N_12614,N_7508,N_9349);
nand U12615 (N_12615,N_9879,N_6114);
or U12616 (N_12616,N_9631,N_8955);
nand U12617 (N_12617,N_9691,N_5935);
nor U12618 (N_12618,N_8698,N_6313);
and U12619 (N_12619,N_8131,N_6051);
nand U12620 (N_12620,N_6887,N_7213);
or U12621 (N_12621,N_6005,N_5034);
nor U12622 (N_12622,N_9966,N_9462);
or U12623 (N_12623,N_5184,N_9983);
nand U12624 (N_12624,N_5944,N_6229);
nor U12625 (N_12625,N_8193,N_8409);
or U12626 (N_12626,N_9927,N_7365);
nor U12627 (N_12627,N_5849,N_6270);
and U12628 (N_12628,N_8219,N_9701);
and U12629 (N_12629,N_7493,N_7244);
or U12630 (N_12630,N_9931,N_9133);
and U12631 (N_12631,N_9123,N_9446);
xor U12632 (N_12632,N_6465,N_8347);
xor U12633 (N_12633,N_7666,N_9001);
nand U12634 (N_12634,N_6204,N_6068);
xnor U12635 (N_12635,N_9265,N_6904);
nand U12636 (N_12636,N_9500,N_8574);
and U12637 (N_12637,N_5103,N_5372);
nand U12638 (N_12638,N_8324,N_7446);
nand U12639 (N_12639,N_8173,N_5392);
or U12640 (N_12640,N_6306,N_5665);
or U12641 (N_12641,N_6594,N_8675);
and U12642 (N_12642,N_8081,N_7789);
nor U12643 (N_12643,N_9276,N_8344);
nor U12644 (N_12644,N_5061,N_7029);
xor U12645 (N_12645,N_7311,N_8134);
or U12646 (N_12646,N_7168,N_9302);
or U12647 (N_12647,N_5399,N_9236);
xor U12648 (N_12648,N_6506,N_6159);
or U12649 (N_12649,N_8875,N_6589);
nor U12650 (N_12650,N_9930,N_6702);
nand U12651 (N_12651,N_8239,N_8821);
nand U12652 (N_12652,N_9752,N_8006);
xnor U12653 (N_12653,N_5002,N_5733);
or U12654 (N_12654,N_8520,N_7871);
xnor U12655 (N_12655,N_5461,N_9989);
nor U12656 (N_12656,N_6018,N_6074);
xor U12657 (N_12657,N_5286,N_5376);
nand U12658 (N_12658,N_8717,N_8624);
xor U12659 (N_12659,N_8983,N_9093);
or U12660 (N_12660,N_5136,N_7118);
nor U12661 (N_12661,N_7357,N_6166);
nor U12662 (N_12662,N_9322,N_5435);
xnor U12663 (N_12663,N_5715,N_7131);
xnor U12664 (N_12664,N_8597,N_6695);
nand U12665 (N_12665,N_5627,N_8183);
nand U12666 (N_12666,N_6497,N_6835);
or U12667 (N_12667,N_8146,N_9318);
and U12668 (N_12668,N_6264,N_6910);
and U12669 (N_12669,N_5040,N_7823);
xnor U12670 (N_12670,N_5362,N_7101);
xnor U12671 (N_12671,N_9150,N_7976);
and U12672 (N_12672,N_6755,N_7345);
nand U12673 (N_12673,N_9699,N_6588);
or U12674 (N_12674,N_9136,N_7994);
nor U12675 (N_12675,N_7022,N_5899);
xnor U12676 (N_12676,N_7606,N_6562);
nor U12677 (N_12677,N_7811,N_5062);
and U12678 (N_12678,N_7821,N_9887);
nand U12679 (N_12679,N_5268,N_6448);
or U12680 (N_12680,N_9585,N_6535);
nand U12681 (N_12681,N_5602,N_9637);
and U12682 (N_12682,N_9464,N_7685);
or U12683 (N_12683,N_7410,N_5984);
or U12684 (N_12684,N_7230,N_6535);
xnor U12685 (N_12685,N_5536,N_5891);
or U12686 (N_12686,N_5295,N_9717);
nand U12687 (N_12687,N_8804,N_5812);
nand U12688 (N_12688,N_5206,N_7180);
nand U12689 (N_12689,N_5700,N_9901);
or U12690 (N_12690,N_9619,N_6686);
xnor U12691 (N_12691,N_9589,N_6776);
or U12692 (N_12692,N_7137,N_7639);
or U12693 (N_12693,N_5813,N_8515);
or U12694 (N_12694,N_9089,N_7630);
and U12695 (N_12695,N_6876,N_9058);
nand U12696 (N_12696,N_7434,N_5611);
nor U12697 (N_12697,N_6334,N_9448);
and U12698 (N_12698,N_7305,N_5252);
xor U12699 (N_12699,N_6640,N_7939);
nand U12700 (N_12700,N_6167,N_7848);
and U12701 (N_12701,N_7124,N_6388);
nand U12702 (N_12702,N_7010,N_6805);
or U12703 (N_12703,N_6701,N_7752);
nor U12704 (N_12704,N_5824,N_6426);
and U12705 (N_12705,N_5133,N_6886);
nand U12706 (N_12706,N_9443,N_7766);
xor U12707 (N_12707,N_8673,N_6091);
and U12708 (N_12708,N_9673,N_9643);
or U12709 (N_12709,N_9677,N_8784);
xor U12710 (N_12710,N_6941,N_7826);
nor U12711 (N_12711,N_6808,N_5904);
or U12712 (N_12712,N_8646,N_9119);
nand U12713 (N_12713,N_8540,N_7895);
and U12714 (N_12714,N_7959,N_5966);
xnor U12715 (N_12715,N_9656,N_8669);
xor U12716 (N_12716,N_9307,N_8385);
nor U12717 (N_12717,N_7076,N_7888);
nand U12718 (N_12718,N_8149,N_5269);
nor U12719 (N_12719,N_6131,N_7205);
xor U12720 (N_12720,N_5015,N_7118);
xnor U12721 (N_12721,N_7586,N_8769);
nor U12722 (N_12722,N_7392,N_8276);
and U12723 (N_12723,N_5426,N_6635);
nor U12724 (N_12724,N_8603,N_7045);
nor U12725 (N_12725,N_5616,N_9405);
or U12726 (N_12726,N_8250,N_9999);
nor U12727 (N_12727,N_5088,N_5589);
nor U12728 (N_12728,N_5327,N_6364);
nor U12729 (N_12729,N_9644,N_8777);
or U12730 (N_12730,N_8266,N_7383);
nor U12731 (N_12731,N_5007,N_5792);
nor U12732 (N_12732,N_8017,N_5472);
xor U12733 (N_12733,N_6218,N_9699);
nand U12734 (N_12734,N_7651,N_5084);
or U12735 (N_12735,N_6752,N_8300);
and U12736 (N_12736,N_6518,N_8747);
and U12737 (N_12737,N_5323,N_8708);
or U12738 (N_12738,N_9487,N_9844);
xnor U12739 (N_12739,N_8253,N_7307);
and U12740 (N_12740,N_5071,N_6059);
nor U12741 (N_12741,N_5889,N_9058);
or U12742 (N_12742,N_6325,N_9178);
or U12743 (N_12743,N_5398,N_7357);
xnor U12744 (N_12744,N_8593,N_8993);
nand U12745 (N_12745,N_7525,N_9336);
nand U12746 (N_12746,N_5377,N_6345);
nand U12747 (N_12747,N_5671,N_8324);
or U12748 (N_12748,N_8409,N_7040);
or U12749 (N_12749,N_6106,N_8452);
or U12750 (N_12750,N_8595,N_7576);
and U12751 (N_12751,N_9382,N_5256);
and U12752 (N_12752,N_9003,N_6125);
or U12753 (N_12753,N_6392,N_5049);
nand U12754 (N_12754,N_7353,N_7168);
nand U12755 (N_12755,N_8651,N_5546);
nand U12756 (N_12756,N_5484,N_7094);
and U12757 (N_12757,N_8890,N_6507);
nand U12758 (N_12758,N_6001,N_5242);
or U12759 (N_12759,N_7641,N_8151);
xnor U12760 (N_12760,N_6441,N_7107);
nor U12761 (N_12761,N_7240,N_6647);
nor U12762 (N_12762,N_9554,N_7111);
nand U12763 (N_12763,N_5649,N_9354);
xnor U12764 (N_12764,N_5481,N_5553);
nor U12765 (N_12765,N_8828,N_5255);
and U12766 (N_12766,N_5109,N_7108);
and U12767 (N_12767,N_6501,N_7409);
nor U12768 (N_12768,N_5468,N_6541);
and U12769 (N_12769,N_9585,N_9054);
or U12770 (N_12770,N_8761,N_7626);
and U12771 (N_12771,N_7473,N_6972);
and U12772 (N_12772,N_6427,N_7345);
nand U12773 (N_12773,N_9785,N_7623);
and U12774 (N_12774,N_8761,N_9800);
xor U12775 (N_12775,N_8516,N_9495);
and U12776 (N_12776,N_7743,N_6920);
xor U12777 (N_12777,N_5224,N_9689);
nand U12778 (N_12778,N_7828,N_6682);
nor U12779 (N_12779,N_7790,N_5547);
or U12780 (N_12780,N_7194,N_5112);
or U12781 (N_12781,N_8557,N_9503);
nand U12782 (N_12782,N_8209,N_7115);
nand U12783 (N_12783,N_9465,N_6359);
and U12784 (N_12784,N_9071,N_6187);
or U12785 (N_12785,N_7586,N_9262);
xor U12786 (N_12786,N_7503,N_6355);
and U12787 (N_12787,N_8208,N_7385);
xor U12788 (N_12788,N_6285,N_6071);
nand U12789 (N_12789,N_5169,N_7522);
nand U12790 (N_12790,N_7796,N_5491);
nand U12791 (N_12791,N_7085,N_9399);
nand U12792 (N_12792,N_8409,N_5407);
xnor U12793 (N_12793,N_5507,N_8294);
nand U12794 (N_12794,N_5949,N_6205);
nor U12795 (N_12795,N_8812,N_9891);
and U12796 (N_12796,N_9847,N_9987);
nand U12797 (N_12797,N_7416,N_9944);
or U12798 (N_12798,N_5236,N_8410);
or U12799 (N_12799,N_7331,N_9062);
xnor U12800 (N_12800,N_8762,N_8684);
and U12801 (N_12801,N_8863,N_9958);
or U12802 (N_12802,N_8692,N_9921);
and U12803 (N_12803,N_8146,N_8249);
and U12804 (N_12804,N_7830,N_5210);
or U12805 (N_12805,N_9911,N_6438);
or U12806 (N_12806,N_8735,N_6045);
xor U12807 (N_12807,N_8706,N_7136);
xnor U12808 (N_12808,N_6568,N_9883);
and U12809 (N_12809,N_8965,N_8488);
xor U12810 (N_12810,N_5436,N_8949);
or U12811 (N_12811,N_7052,N_9728);
or U12812 (N_12812,N_7653,N_7031);
and U12813 (N_12813,N_7964,N_5067);
or U12814 (N_12814,N_5920,N_5450);
xnor U12815 (N_12815,N_7745,N_6157);
xor U12816 (N_12816,N_7890,N_6942);
and U12817 (N_12817,N_9364,N_7699);
nor U12818 (N_12818,N_6806,N_9469);
nor U12819 (N_12819,N_9367,N_7518);
nand U12820 (N_12820,N_8003,N_6849);
xnor U12821 (N_12821,N_8768,N_5345);
xor U12822 (N_12822,N_7173,N_7143);
xnor U12823 (N_12823,N_6925,N_9448);
nand U12824 (N_12824,N_6604,N_6585);
xor U12825 (N_12825,N_6416,N_7861);
and U12826 (N_12826,N_7821,N_6036);
and U12827 (N_12827,N_7987,N_8352);
xnor U12828 (N_12828,N_6868,N_9681);
or U12829 (N_12829,N_8496,N_8732);
nor U12830 (N_12830,N_8956,N_9809);
nand U12831 (N_12831,N_6227,N_6706);
xnor U12832 (N_12832,N_5505,N_9644);
xnor U12833 (N_12833,N_7585,N_7270);
and U12834 (N_12834,N_8866,N_6214);
nor U12835 (N_12835,N_6107,N_8015);
xor U12836 (N_12836,N_5327,N_8430);
nand U12837 (N_12837,N_6539,N_7760);
and U12838 (N_12838,N_6793,N_8621);
nand U12839 (N_12839,N_5765,N_9148);
or U12840 (N_12840,N_8323,N_7155);
or U12841 (N_12841,N_8290,N_9858);
xor U12842 (N_12842,N_9559,N_7990);
and U12843 (N_12843,N_5214,N_6744);
and U12844 (N_12844,N_5642,N_8991);
xnor U12845 (N_12845,N_9429,N_6495);
and U12846 (N_12846,N_8085,N_8058);
nand U12847 (N_12847,N_7956,N_6125);
and U12848 (N_12848,N_6801,N_6062);
and U12849 (N_12849,N_5299,N_9670);
or U12850 (N_12850,N_8009,N_6794);
or U12851 (N_12851,N_6955,N_7936);
or U12852 (N_12852,N_9742,N_5900);
nand U12853 (N_12853,N_7802,N_6280);
nor U12854 (N_12854,N_7141,N_9461);
nand U12855 (N_12855,N_8264,N_9778);
or U12856 (N_12856,N_8023,N_9634);
and U12857 (N_12857,N_7274,N_9901);
or U12858 (N_12858,N_7140,N_9997);
nor U12859 (N_12859,N_8353,N_8020);
and U12860 (N_12860,N_8481,N_9212);
nand U12861 (N_12861,N_9558,N_8788);
xor U12862 (N_12862,N_5161,N_8737);
xor U12863 (N_12863,N_6846,N_9683);
xnor U12864 (N_12864,N_9592,N_8317);
nor U12865 (N_12865,N_7535,N_5248);
nand U12866 (N_12866,N_6992,N_6335);
and U12867 (N_12867,N_9023,N_6928);
nand U12868 (N_12868,N_8044,N_8473);
xnor U12869 (N_12869,N_5966,N_8054);
nor U12870 (N_12870,N_6326,N_8041);
nor U12871 (N_12871,N_9941,N_8402);
nand U12872 (N_12872,N_6030,N_6855);
nand U12873 (N_12873,N_9044,N_8014);
nand U12874 (N_12874,N_8664,N_6084);
or U12875 (N_12875,N_7655,N_6839);
nand U12876 (N_12876,N_9549,N_8544);
nor U12877 (N_12877,N_8544,N_8305);
and U12878 (N_12878,N_6033,N_6982);
nand U12879 (N_12879,N_6532,N_6762);
nor U12880 (N_12880,N_7492,N_6387);
xor U12881 (N_12881,N_8429,N_8921);
nor U12882 (N_12882,N_8099,N_9664);
nand U12883 (N_12883,N_6172,N_9917);
and U12884 (N_12884,N_8158,N_9668);
or U12885 (N_12885,N_9480,N_9202);
or U12886 (N_12886,N_6436,N_8828);
or U12887 (N_12887,N_7810,N_6620);
nor U12888 (N_12888,N_5468,N_7891);
xor U12889 (N_12889,N_7254,N_8833);
and U12890 (N_12890,N_8560,N_7089);
nor U12891 (N_12891,N_9706,N_5496);
or U12892 (N_12892,N_7994,N_5299);
nor U12893 (N_12893,N_8593,N_9773);
and U12894 (N_12894,N_8606,N_9240);
and U12895 (N_12895,N_5709,N_5316);
nor U12896 (N_12896,N_9825,N_5241);
nor U12897 (N_12897,N_5306,N_8204);
and U12898 (N_12898,N_8913,N_9827);
or U12899 (N_12899,N_6529,N_5381);
and U12900 (N_12900,N_6899,N_9533);
or U12901 (N_12901,N_9234,N_5167);
and U12902 (N_12902,N_9735,N_8032);
or U12903 (N_12903,N_9218,N_8042);
nand U12904 (N_12904,N_5012,N_6246);
xor U12905 (N_12905,N_7440,N_7546);
nand U12906 (N_12906,N_9160,N_8114);
xor U12907 (N_12907,N_7254,N_9269);
xor U12908 (N_12908,N_5119,N_7843);
nand U12909 (N_12909,N_6441,N_6471);
nor U12910 (N_12910,N_7807,N_8603);
nor U12911 (N_12911,N_7089,N_5524);
nor U12912 (N_12912,N_6242,N_9532);
and U12913 (N_12913,N_9894,N_6767);
nand U12914 (N_12914,N_8193,N_6610);
or U12915 (N_12915,N_5709,N_8509);
and U12916 (N_12916,N_8061,N_5966);
nand U12917 (N_12917,N_7446,N_5508);
and U12918 (N_12918,N_6883,N_6415);
nor U12919 (N_12919,N_5329,N_9275);
nor U12920 (N_12920,N_8476,N_7536);
or U12921 (N_12921,N_6081,N_5927);
and U12922 (N_12922,N_9817,N_8324);
or U12923 (N_12923,N_5973,N_9581);
and U12924 (N_12924,N_5088,N_9771);
xor U12925 (N_12925,N_7689,N_5767);
and U12926 (N_12926,N_5360,N_9438);
and U12927 (N_12927,N_5008,N_6772);
nor U12928 (N_12928,N_7173,N_6107);
or U12929 (N_12929,N_7610,N_6589);
nor U12930 (N_12930,N_9874,N_8835);
xor U12931 (N_12931,N_7340,N_8449);
nor U12932 (N_12932,N_8448,N_6482);
or U12933 (N_12933,N_7335,N_7066);
nor U12934 (N_12934,N_9546,N_6045);
or U12935 (N_12935,N_7797,N_5572);
or U12936 (N_12936,N_8202,N_6178);
and U12937 (N_12937,N_6119,N_8047);
or U12938 (N_12938,N_5159,N_7944);
or U12939 (N_12939,N_5274,N_9554);
and U12940 (N_12940,N_7778,N_6928);
and U12941 (N_12941,N_5800,N_8942);
and U12942 (N_12942,N_9308,N_5408);
nand U12943 (N_12943,N_5519,N_8298);
nand U12944 (N_12944,N_9289,N_6617);
and U12945 (N_12945,N_7011,N_7188);
nand U12946 (N_12946,N_9944,N_5971);
or U12947 (N_12947,N_7254,N_7075);
nand U12948 (N_12948,N_9284,N_5435);
and U12949 (N_12949,N_7530,N_7499);
nand U12950 (N_12950,N_6751,N_5733);
and U12951 (N_12951,N_6386,N_5546);
or U12952 (N_12952,N_5685,N_8878);
nand U12953 (N_12953,N_6652,N_6308);
nand U12954 (N_12954,N_6246,N_6885);
and U12955 (N_12955,N_7552,N_7249);
nand U12956 (N_12956,N_8372,N_8238);
xor U12957 (N_12957,N_9733,N_9671);
nor U12958 (N_12958,N_8809,N_8162);
and U12959 (N_12959,N_9955,N_8452);
xor U12960 (N_12960,N_6913,N_7468);
xnor U12961 (N_12961,N_9170,N_8459);
xnor U12962 (N_12962,N_7942,N_6647);
or U12963 (N_12963,N_6770,N_5253);
nand U12964 (N_12964,N_7587,N_7202);
nor U12965 (N_12965,N_7482,N_8237);
nand U12966 (N_12966,N_5982,N_7150);
and U12967 (N_12967,N_5013,N_5435);
nor U12968 (N_12968,N_7826,N_7965);
nor U12969 (N_12969,N_8045,N_6694);
or U12970 (N_12970,N_7327,N_8831);
or U12971 (N_12971,N_9267,N_5940);
nor U12972 (N_12972,N_8751,N_5692);
or U12973 (N_12973,N_9106,N_8810);
or U12974 (N_12974,N_9608,N_6989);
xor U12975 (N_12975,N_8225,N_6023);
nand U12976 (N_12976,N_5832,N_8377);
nand U12977 (N_12977,N_7080,N_7533);
and U12978 (N_12978,N_6697,N_5063);
nand U12979 (N_12979,N_7355,N_9746);
and U12980 (N_12980,N_7955,N_7987);
xor U12981 (N_12981,N_6908,N_7507);
or U12982 (N_12982,N_9681,N_5402);
or U12983 (N_12983,N_9234,N_6554);
or U12984 (N_12984,N_6234,N_6622);
xnor U12985 (N_12985,N_6091,N_7571);
nand U12986 (N_12986,N_9255,N_9226);
or U12987 (N_12987,N_7642,N_6733);
and U12988 (N_12988,N_5793,N_6274);
nand U12989 (N_12989,N_8233,N_5552);
nand U12990 (N_12990,N_5654,N_8943);
or U12991 (N_12991,N_9712,N_9203);
and U12992 (N_12992,N_7584,N_7109);
nand U12993 (N_12993,N_9782,N_9377);
xor U12994 (N_12994,N_6535,N_7328);
xnor U12995 (N_12995,N_6339,N_5837);
nor U12996 (N_12996,N_5293,N_9142);
and U12997 (N_12997,N_7221,N_9399);
and U12998 (N_12998,N_9672,N_5302);
and U12999 (N_12999,N_9018,N_9718);
nand U13000 (N_13000,N_6138,N_7017);
xor U13001 (N_13001,N_7907,N_5827);
nor U13002 (N_13002,N_9513,N_5486);
nand U13003 (N_13003,N_5695,N_6593);
nand U13004 (N_13004,N_6304,N_9121);
or U13005 (N_13005,N_6769,N_9545);
and U13006 (N_13006,N_9977,N_5413);
or U13007 (N_13007,N_9574,N_9422);
xor U13008 (N_13008,N_7403,N_9568);
or U13009 (N_13009,N_7215,N_5404);
xnor U13010 (N_13010,N_7472,N_9442);
or U13011 (N_13011,N_7211,N_6806);
nand U13012 (N_13012,N_8555,N_7851);
or U13013 (N_13013,N_6507,N_8707);
nor U13014 (N_13014,N_5583,N_8200);
nor U13015 (N_13015,N_6599,N_8114);
or U13016 (N_13016,N_7624,N_8362);
and U13017 (N_13017,N_8305,N_9859);
or U13018 (N_13018,N_6174,N_7001);
or U13019 (N_13019,N_7431,N_5109);
nand U13020 (N_13020,N_8042,N_6220);
nor U13021 (N_13021,N_6699,N_6503);
nor U13022 (N_13022,N_5549,N_9399);
and U13023 (N_13023,N_6208,N_9324);
nor U13024 (N_13024,N_9797,N_5244);
nor U13025 (N_13025,N_5078,N_9519);
and U13026 (N_13026,N_8850,N_9909);
xor U13027 (N_13027,N_5664,N_8005);
and U13028 (N_13028,N_8614,N_5575);
nor U13029 (N_13029,N_6005,N_5497);
or U13030 (N_13030,N_7245,N_6956);
or U13031 (N_13031,N_6399,N_8964);
and U13032 (N_13032,N_8785,N_6320);
or U13033 (N_13033,N_5835,N_5023);
nand U13034 (N_13034,N_6357,N_5247);
and U13035 (N_13035,N_9914,N_8662);
xor U13036 (N_13036,N_7220,N_8958);
nand U13037 (N_13037,N_6414,N_6275);
and U13038 (N_13038,N_6416,N_8589);
xor U13039 (N_13039,N_7192,N_6526);
nand U13040 (N_13040,N_5571,N_9515);
and U13041 (N_13041,N_7059,N_7794);
and U13042 (N_13042,N_7974,N_8334);
xnor U13043 (N_13043,N_9501,N_9092);
or U13044 (N_13044,N_5018,N_8371);
and U13045 (N_13045,N_6382,N_7188);
nor U13046 (N_13046,N_9151,N_8929);
xnor U13047 (N_13047,N_9103,N_5528);
nand U13048 (N_13048,N_7547,N_7160);
nor U13049 (N_13049,N_7683,N_5987);
and U13050 (N_13050,N_8766,N_7423);
xor U13051 (N_13051,N_6496,N_5891);
or U13052 (N_13052,N_6026,N_5580);
nand U13053 (N_13053,N_9622,N_7177);
nor U13054 (N_13054,N_9520,N_5645);
nand U13055 (N_13055,N_8718,N_8083);
and U13056 (N_13056,N_7772,N_6446);
and U13057 (N_13057,N_7755,N_5899);
xor U13058 (N_13058,N_7772,N_5638);
nand U13059 (N_13059,N_7216,N_6956);
xor U13060 (N_13060,N_7819,N_7305);
xor U13061 (N_13061,N_5860,N_7277);
xnor U13062 (N_13062,N_7908,N_6917);
and U13063 (N_13063,N_5938,N_8378);
or U13064 (N_13064,N_7131,N_8878);
and U13065 (N_13065,N_6214,N_9887);
xor U13066 (N_13066,N_8511,N_8049);
nor U13067 (N_13067,N_7963,N_8897);
nand U13068 (N_13068,N_9731,N_8890);
nor U13069 (N_13069,N_6939,N_9692);
nand U13070 (N_13070,N_6114,N_7827);
nand U13071 (N_13071,N_9938,N_5231);
xnor U13072 (N_13072,N_5995,N_6400);
xor U13073 (N_13073,N_6522,N_8501);
nor U13074 (N_13074,N_8048,N_8340);
xnor U13075 (N_13075,N_9164,N_6178);
nand U13076 (N_13076,N_8044,N_7921);
and U13077 (N_13077,N_7432,N_8460);
or U13078 (N_13078,N_7948,N_8860);
and U13079 (N_13079,N_8878,N_8858);
xor U13080 (N_13080,N_5972,N_5802);
or U13081 (N_13081,N_6534,N_5673);
and U13082 (N_13082,N_5184,N_7501);
nor U13083 (N_13083,N_5424,N_6639);
and U13084 (N_13084,N_5585,N_7616);
xnor U13085 (N_13085,N_8702,N_5692);
nand U13086 (N_13086,N_7881,N_7922);
and U13087 (N_13087,N_6667,N_9047);
nand U13088 (N_13088,N_5002,N_6497);
or U13089 (N_13089,N_6959,N_9633);
nand U13090 (N_13090,N_8915,N_9418);
nand U13091 (N_13091,N_7953,N_5206);
and U13092 (N_13092,N_7939,N_8083);
nor U13093 (N_13093,N_8753,N_8324);
nor U13094 (N_13094,N_8563,N_5676);
xor U13095 (N_13095,N_5819,N_5722);
and U13096 (N_13096,N_6466,N_7873);
xnor U13097 (N_13097,N_9269,N_7419);
or U13098 (N_13098,N_5886,N_9484);
and U13099 (N_13099,N_5048,N_9835);
and U13100 (N_13100,N_9867,N_7255);
or U13101 (N_13101,N_5974,N_8026);
or U13102 (N_13102,N_9002,N_8166);
and U13103 (N_13103,N_5960,N_7206);
xnor U13104 (N_13104,N_9452,N_7534);
xnor U13105 (N_13105,N_7165,N_7342);
nor U13106 (N_13106,N_6266,N_5994);
xnor U13107 (N_13107,N_9804,N_6906);
nor U13108 (N_13108,N_8951,N_7761);
and U13109 (N_13109,N_9512,N_5978);
nor U13110 (N_13110,N_6844,N_8903);
nor U13111 (N_13111,N_6851,N_8600);
nor U13112 (N_13112,N_5763,N_6270);
or U13113 (N_13113,N_8358,N_5231);
or U13114 (N_13114,N_5155,N_5368);
xnor U13115 (N_13115,N_8180,N_9532);
nand U13116 (N_13116,N_8916,N_5828);
or U13117 (N_13117,N_8224,N_9216);
xnor U13118 (N_13118,N_9649,N_9767);
xnor U13119 (N_13119,N_5438,N_5499);
nand U13120 (N_13120,N_5648,N_6278);
and U13121 (N_13121,N_7413,N_9912);
nand U13122 (N_13122,N_6081,N_9505);
xor U13123 (N_13123,N_8853,N_5667);
or U13124 (N_13124,N_9691,N_8800);
xnor U13125 (N_13125,N_5419,N_6630);
xnor U13126 (N_13126,N_8778,N_8528);
xnor U13127 (N_13127,N_5910,N_9829);
or U13128 (N_13128,N_9733,N_9157);
xor U13129 (N_13129,N_5137,N_6929);
nand U13130 (N_13130,N_9419,N_5073);
or U13131 (N_13131,N_6814,N_9811);
xor U13132 (N_13132,N_5589,N_8434);
nor U13133 (N_13133,N_9828,N_5999);
and U13134 (N_13134,N_8723,N_6688);
nor U13135 (N_13135,N_8471,N_6850);
and U13136 (N_13136,N_8016,N_6927);
and U13137 (N_13137,N_6888,N_8847);
xor U13138 (N_13138,N_8488,N_6353);
xor U13139 (N_13139,N_7347,N_9758);
and U13140 (N_13140,N_6387,N_6499);
and U13141 (N_13141,N_7993,N_6001);
or U13142 (N_13142,N_7444,N_5262);
nor U13143 (N_13143,N_6348,N_6106);
and U13144 (N_13144,N_8652,N_5652);
or U13145 (N_13145,N_7511,N_6310);
or U13146 (N_13146,N_8596,N_8073);
xnor U13147 (N_13147,N_9837,N_6102);
and U13148 (N_13148,N_6040,N_6389);
xor U13149 (N_13149,N_7676,N_8865);
or U13150 (N_13150,N_5034,N_7014);
nand U13151 (N_13151,N_5995,N_7443);
or U13152 (N_13152,N_9575,N_6813);
nor U13153 (N_13153,N_9664,N_6334);
and U13154 (N_13154,N_6758,N_5836);
nand U13155 (N_13155,N_8899,N_5853);
or U13156 (N_13156,N_9211,N_8503);
nor U13157 (N_13157,N_5617,N_7275);
nand U13158 (N_13158,N_6844,N_6999);
nand U13159 (N_13159,N_9975,N_8741);
xor U13160 (N_13160,N_7271,N_7626);
nor U13161 (N_13161,N_9487,N_6952);
nand U13162 (N_13162,N_7686,N_9038);
nor U13163 (N_13163,N_7523,N_7163);
and U13164 (N_13164,N_9411,N_8908);
nand U13165 (N_13165,N_9331,N_8673);
xor U13166 (N_13166,N_9868,N_8849);
xnor U13167 (N_13167,N_7648,N_6812);
nor U13168 (N_13168,N_5942,N_7792);
xnor U13169 (N_13169,N_7809,N_9958);
or U13170 (N_13170,N_6364,N_5271);
xor U13171 (N_13171,N_5155,N_6960);
or U13172 (N_13172,N_9737,N_5454);
or U13173 (N_13173,N_5730,N_8360);
or U13174 (N_13174,N_8933,N_7202);
nor U13175 (N_13175,N_9542,N_6952);
nor U13176 (N_13176,N_6455,N_5614);
or U13177 (N_13177,N_6445,N_5897);
and U13178 (N_13178,N_9087,N_5162);
nand U13179 (N_13179,N_5416,N_8206);
xor U13180 (N_13180,N_7540,N_8595);
xnor U13181 (N_13181,N_7999,N_6371);
xor U13182 (N_13182,N_5445,N_8338);
and U13183 (N_13183,N_7636,N_7974);
and U13184 (N_13184,N_6657,N_9858);
xor U13185 (N_13185,N_6326,N_8211);
or U13186 (N_13186,N_5046,N_8277);
nor U13187 (N_13187,N_5058,N_9341);
or U13188 (N_13188,N_9359,N_8436);
xor U13189 (N_13189,N_7827,N_9150);
nand U13190 (N_13190,N_8915,N_8237);
or U13191 (N_13191,N_6031,N_6255);
and U13192 (N_13192,N_9991,N_7614);
or U13193 (N_13193,N_9402,N_7874);
or U13194 (N_13194,N_9233,N_7969);
nand U13195 (N_13195,N_6250,N_5901);
xor U13196 (N_13196,N_9010,N_8508);
xnor U13197 (N_13197,N_8225,N_7050);
xor U13198 (N_13198,N_6408,N_8441);
and U13199 (N_13199,N_6256,N_8414);
or U13200 (N_13200,N_7136,N_8423);
nor U13201 (N_13201,N_9313,N_5664);
or U13202 (N_13202,N_5487,N_6951);
and U13203 (N_13203,N_7955,N_8327);
nand U13204 (N_13204,N_9505,N_5390);
and U13205 (N_13205,N_7704,N_9955);
or U13206 (N_13206,N_5099,N_5160);
nor U13207 (N_13207,N_5785,N_8124);
xnor U13208 (N_13208,N_8760,N_6993);
xnor U13209 (N_13209,N_8623,N_9102);
nand U13210 (N_13210,N_7006,N_8949);
or U13211 (N_13211,N_8522,N_9143);
and U13212 (N_13212,N_6796,N_8455);
nor U13213 (N_13213,N_8350,N_5227);
nor U13214 (N_13214,N_8725,N_8851);
nor U13215 (N_13215,N_7368,N_7469);
and U13216 (N_13216,N_6301,N_8115);
or U13217 (N_13217,N_7425,N_8718);
xor U13218 (N_13218,N_6887,N_6603);
nor U13219 (N_13219,N_7569,N_7976);
nand U13220 (N_13220,N_7895,N_7058);
xor U13221 (N_13221,N_9093,N_6442);
nor U13222 (N_13222,N_5964,N_8371);
nor U13223 (N_13223,N_8081,N_5586);
xnor U13224 (N_13224,N_6732,N_8259);
xnor U13225 (N_13225,N_7489,N_5993);
and U13226 (N_13226,N_5656,N_7346);
or U13227 (N_13227,N_7491,N_8921);
or U13228 (N_13228,N_5344,N_6530);
xnor U13229 (N_13229,N_5150,N_9206);
nor U13230 (N_13230,N_8728,N_5999);
nand U13231 (N_13231,N_6387,N_6892);
nor U13232 (N_13232,N_7067,N_5273);
or U13233 (N_13233,N_5791,N_7704);
xor U13234 (N_13234,N_5859,N_5110);
and U13235 (N_13235,N_7695,N_8912);
or U13236 (N_13236,N_5209,N_9886);
xnor U13237 (N_13237,N_5798,N_7231);
xnor U13238 (N_13238,N_5938,N_8791);
and U13239 (N_13239,N_5759,N_5607);
and U13240 (N_13240,N_5601,N_5208);
nor U13241 (N_13241,N_6020,N_8437);
or U13242 (N_13242,N_9158,N_6490);
xnor U13243 (N_13243,N_5458,N_8593);
nor U13244 (N_13244,N_5238,N_6978);
xor U13245 (N_13245,N_5568,N_6296);
and U13246 (N_13246,N_9895,N_5894);
or U13247 (N_13247,N_9564,N_6688);
and U13248 (N_13248,N_6965,N_6319);
nor U13249 (N_13249,N_6686,N_8562);
nand U13250 (N_13250,N_7652,N_9784);
xor U13251 (N_13251,N_9236,N_7795);
nand U13252 (N_13252,N_8459,N_7485);
nor U13253 (N_13253,N_8781,N_7620);
nor U13254 (N_13254,N_5946,N_9196);
xor U13255 (N_13255,N_5004,N_9391);
xnor U13256 (N_13256,N_9973,N_5101);
or U13257 (N_13257,N_5907,N_7864);
xor U13258 (N_13258,N_9428,N_5110);
or U13259 (N_13259,N_8886,N_5636);
xor U13260 (N_13260,N_7299,N_8933);
nand U13261 (N_13261,N_8342,N_7362);
xor U13262 (N_13262,N_7294,N_9181);
xor U13263 (N_13263,N_6915,N_8306);
and U13264 (N_13264,N_7942,N_6645);
or U13265 (N_13265,N_9730,N_7966);
nand U13266 (N_13266,N_5446,N_6958);
xor U13267 (N_13267,N_9975,N_7337);
nor U13268 (N_13268,N_8896,N_6718);
nor U13269 (N_13269,N_8684,N_5647);
and U13270 (N_13270,N_6836,N_7776);
or U13271 (N_13271,N_7416,N_6017);
xor U13272 (N_13272,N_9494,N_6525);
xor U13273 (N_13273,N_8622,N_5189);
nor U13274 (N_13274,N_5062,N_8140);
and U13275 (N_13275,N_6368,N_6496);
nand U13276 (N_13276,N_5542,N_7509);
xor U13277 (N_13277,N_8974,N_9771);
and U13278 (N_13278,N_5230,N_7968);
nand U13279 (N_13279,N_8548,N_9378);
and U13280 (N_13280,N_8822,N_5656);
and U13281 (N_13281,N_9534,N_8724);
nor U13282 (N_13282,N_6181,N_5725);
xnor U13283 (N_13283,N_8874,N_5875);
nor U13284 (N_13284,N_8188,N_5278);
and U13285 (N_13285,N_8716,N_9113);
nand U13286 (N_13286,N_5599,N_6684);
and U13287 (N_13287,N_7103,N_5096);
nand U13288 (N_13288,N_8375,N_8015);
or U13289 (N_13289,N_8209,N_7865);
nand U13290 (N_13290,N_5555,N_6862);
xor U13291 (N_13291,N_6672,N_6554);
nor U13292 (N_13292,N_8445,N_7618);
or U13293 (N_13293,N_9377,N_7911);
or U13294 (N_13294,N_5080,N_8637);
nand U13295 (N_13295,N_6716,N_7199);
and U13296 (N_13296,N_7346,N_5752);
or U13297 (N_13297,N_8709,N_7011);
or U13298 (N_13298,N_8835,N_9059);
nor U13299 (N_13299,N_5133,N_9815);
or U13300 (N_13300,N_9507,N_5246);
xor U13301 (N_13301,N_7578,N_8488);
nor U13302 (N_13302,N_7203,N_9305);
nand U13303 (N_13303,N_5182,N_7849);
or U13304 (N_13304,N_8666,N_5762);
nor U13305 (N_13305,N_6693,N_5309);
nor U13306 (N_13306,N_7454,N_8303);
and U13307 (N_13307,N_9007,N_7638);
or U13308 (N_13308,N_8571,N_9570);
or U13309 (N_13309,N_7957,N_8347);
or U13310 (N_13310,N_5970,N_6977);
or U13311 (N_13311,N_5438,N_8831);
or U13312 (N_13312,N_9018,N_8439);
xor U13313 (N_13313,N_5501,N_9332);
xor U13314 (N_13314,N_9287,N_9289);
nor U13315 (N_13315,N_9061,N_5416);
nand U13316 (N_13316,N_8631,N_5655);
xnor U13317 (N_13317,N_8519,N_8787);
xor U13318 (N_13318,N_6294,N_6048);
xor U13319 (N_13319,N_5661,N_6905);
and U13320 (N_13320,N_8694,N_6843);
nor U13321 (N_13321,N_7303,N_8209);
xnor U13322 (N_13322,N_7493,N_5573);
xnor U13323 (N_13323,N_5600,N_7012);
or U13324 (N_13324,N_9249,N_7122);
nand U13325 (N_13325,N_9536,N_7072);
and U13326 (N_13326,N_7404,N_9277);
or U13327 (N_13327,N_7803,N_9091);
nor U13328 (N_13328,N_6861,N_9218);
nor U13329 (N_13329,N_8772,N_5141);
or U13330 (N_13330,N_5626,N_5571);
or U13331 (N_13331,N_9236,N_9642);
or U13332 (N_13332,N_8708,N_8390);
and U13333 (N_13333,N_8881,N_6877);
xnor U13334 (N_13334,N_5044,N_9600);
xnor U13335 (N_13335,N_6629,N_8779);
nand U13336 (N_13336,N_6349,N_5609);
nand U13337 (N_13337,N_8613,N_9586);
nand U13338 (N_13338,N_9546,N_8660);
xnor U13339 (N_13339,N_5323,N_8692);
or U13340 (N_13340,N_5283,N_6699);
nand U13341 (N_13341,N_9016,N_8212);
or U13342 (N_13342,N_5314,N_8070);
and U13343 (N_13343,N_6013,N_5465);
nand U13344 (N_13344,N_6581,N_5332);
nor U13345 (N_13345,N_7618,N_8054);
or U13346 (N_13346,N_5531,N_6517);
xor U13347 (N_13347,N_6904,N_5364);
and U13348 (N_13348,N_5292,N_7918);
nor U13349 (N_13349,N_8411,N_8917);
and U13350 (N_13350,N_8338,N_5294);
or U13351 (N_13351,N_7168,N_6389);
xnor U13352 (N_13352,N_7133,N_6697);
or U13353 (N_13353,N_7536,N_6216);
nor U13354 (N_13354,N_5037,N_9486);
and U13355 (N_13355,N_9010,N_6220);
or U13356 (N_13356,N_6712,N_6893);
xor U13357 (N_13357,N_6137,N_9339);
or U13358 (N_13358,N_8671,N_9392);
xor U13359 (N_13359,N_8283,N_7016);
nor U13360 (N_13360,N_6178,N_8746);
nor U13361 (N_13361,N_5271,N_6202);
and U13362 (N_13362,N_7824,N_6228);
nand U13363 (N_13363,N_5370,N_8564);
nand U13364 (N_13364,N_8210,N_6087);
or U13365 (N_13365,N_5453,N_6035);
nand U13366 (N_13366,N_9023,N_5213);
xor U13367 (N_13367,N_8328,N_8023);
nor U13368 (N_13368,N_7742,N_6341);
xnor U13369 (N_13369,N_7782,N_6203);
and U13370 (N_13370,N_7827,N_6863);
nand U13371 (N_13371,N_9294,N_6475);
and U13372 (N_13372,N_7961,N_9411);
or U13373 (N_13373,N_5936,N_5013);
xnor U13374 (N_13374,N_9440,N_7637);
nand U13375 (N_13375,N_7342,N_8968);
and U13376 (N_13376,N_9474,N_7847);
nor U13377 (N_13377,N_6358,N_5429);
nor U13378 (N_13378,N_9854,N_6589);
nand U13379 (N_13379,N_9584,N_8666);
or U13380 (N_13380,N_6667,N_7393);
or U13381 (N_13381,N_7090,N_7228);
or U13382 (N_13382,N_7882,N_5854);
nand U13383 (N_13383,N_5113,N_5955);
nand U13384 (N_13384,N_7943,N_5354);
and U13385 (N_13385,N_9444,N_8761);
nor U13386 (N_13386,N_8400,N_6072);
xnor U13387 (N_13387,N_6440,N_7867);
and U13388 (N_13388,N_6897,N_7959);
xor U13389 (N_13389,N_5159,N_9280);
or U13390 (N_13390,N_8113,N_8227);
and U13391 (N_13391,N_7682,N_7812);
nand U13392 (N_13392,N_6100,N_5948);
nand U13393 (N_13393,N_6732,N_5988);
or U13394 (N_13394,N_7780,N_6486);
and U13395 (N_13395,N_9860,N_8911);
or U13396 (N_13396,N_9422,N_5085);
nor U13397 (N_13397,N_7176,N_9693);
nor U13398 (N_13398,N_6396,N_7795);
xor U13399 (N_13399,N_9442,N_9445);
and U13400 (N_13400,N_5048,N_7319);
and U13401 (N_13401,N_9876,N_9133);
or U13402 (N_13402,N_8637,N_8762);
nand U13403 (N_13403,N_5316,N_9855);
or U13404 (N_13404,N_5419,N_5603);
nor U13405 (N_13405,N_8692,N_8665);
and U13406 (N_13406,N_6569,N_9675);
nor U13407 (N_13407,N_7810,N_5524);
or U13408 (N_13408,N_8877,N_8446);
nand U13409 (N_13409,N_7691,N_7099);
or U13410 (N_13410,N_9985,N_8741);
and U13411 (N_13411,N_8282,N_6128);
xnor U13412 (N_13412,N_6036,N_8585);
nand U13413 (N_13413,N_8614,N_5163);
or U13414 (N_13414,N_8942,N_6432);
and U13415 (N_13415,N_7869,N_8580);
and U13416 (N_13416,N_5509,N_6855);
nand U13417 (N_13417,N_6086,N_9881);
or U13418 (N_13418,N_9622,N_7254);
nand U13419 (N_13419,N_9132,N_6712);
and U13420 (N_13420,N_8899,N_7619);
nand U13421 (N_13421,N_8438,N_5336);
nand U13422 (N_13422,N_7592,N_6721);
or U13423 (N_13423,N_7480,N_8807);
nand U13424 (N_13424,N_8221,N_6890);
nand U13425 (N_13425,N_7770,N_5148);
xor U13426 (N_13426,N_6495,N_9657);
or U13427 (N_13427,N_8635,N_7155);
nand U13428 (N_13428,N_8971,N_5035);
nand U13429 (N_13429,N_8771,N_8325);
nand U13430 (N_13430,N_7777,N_9311);
xor U13431 (N_13431,N_9872,N_9012);
nand U13432 (N_13432,N_9132,N_9492);
and U13433 (N_13433,N_7058,N_7216);
xnor U13434 (N_13434,N_7384,N_7624);
xor U13435 (N_13435,N_8612,N_5815);
or U13436 (N_13436,N_5408,N_9812);
xnor U13437 (N_13437,N_6951,N_9345);
nand U13438 (N_13438,N_9867,N_7773);
xnor U13439 (N_13439,N_5256,N_9277);
and U13440 (N_13440,N_9974,N_9730);
xor U13441 (N_13441,N_6894,N_8362);
nor U13442 (N_13442,N_7938,N_8654);
or U13443 (N_13443,N_8961,N_5095);
nand U13444 (N_13444,N_8963,N_7967);
nand U13445 (N_13445,N_6051,N_6558);
xnor U13446 (N_13446,N_6690,N_9361);
nor U13447 (N_13447,N_9366,N_7447);
xor U13448 (N_13448,N_7250,N_8743);
or U13449 (N_13449,N_8980,N_5250);
and U13450 (N_13450,N_8270,N_8170);
and U13451 (N_13451,N_6659,N_7538);
nor U13452 (N_13452,N_5911,N_5211);
xnor U13453 (N_13453,N_6623,N_6284);
and U13454 (N_13454,N_6633,N_9544);
and U13455 (N_13455,N_6502,N_8602);
or U13456 (N_13456,N_8058,N_8570);
nand U13457 (N_13457,N_6241,N_9951);
nand U13458 (N_13458,N_9721,N_6561);
or U13459 (N_13459,N_8288,N_6148);
or U13460 (N_13460,N_5401,N_9028);
nor U13461 (N_13461,N_5725,N_9834);
nor U13462 (N_13462,N_6042,N_5803);
nor U13463 (N_13463,N_7843,N_6025);
or U13464 (N_13464,N_9291,N_9029);
nand U13465 (N_13465,N_5987,N_8959);
xor U13466 (N_13466,N_6553,N_8743);
nand U13467 (N_13467,N_7217,N_5936);
xor U13468 (N_13468,N_7209,N_5578);
and U13469 (N_13469,N_6369,N_9131);
xnor U13470 (N_13470,N_7135,N_6546);
and U13471 (N_13471,N_9686,N_5628);
nor U13472 (N_13472,N_7673,N_6214);
or U13473 (N_13473,N_5253,N_8072);
xnor U13474 (N_13474,N_6985,N_9447);
xnor U13475 (N_13475,N_9105,N_5797);
nand U13476 (N_13476,N_8655,N_8296);
nand U13477 (N_13477,N_9922,N_5299);
and U13478 (N_13478,N_6147,N_5074);
nand U13479 (N_13479,N_8586,N_8577);
and U13480 (N_13480,N_9115,N_6112);
nand U13481 (N_13481,N_7035,N_5656);
xor U13482 (N_13482,N_7643,N_5294);
and U13483 (N_13483,N_7337,N_6738);
or U13484 (N_13484,N_8546,N_7401);
nor U13485 (N_13485,N_8208,N_6187);
xor U13486 (N_13486,N_5807,N_9222);
nand U13487 (N_13487,N_6344,N_7320);
xor U13488 (N_13488,N_6985,N_5560);
or U13489 (N_13489,N_8020,N_7393);
and U13490 (N_13490,N_7959,N_8385);
nand U13491 (N_13491,N_6955,N_7201);
nand U13492 (N_13492,N_5357,N_7320);
or U13493 (N_13493,N_8302,N_6599);
xor U13494 (N_13494,N_6361,N_7474);
nand U13495 (N_13495,N_6245,N_8428);
nand U13496 (N_13496,N_9024,N_7729);
or U13497 (N_13497,N_5660,N_8347);
xor U13498 (N_13498,N_8999,N_9221);
or U13499 (N_13499,N_9907,N_8228);
xnor U13500 (N_13500,N_5761,N_5478);
nor U13501 (N_13501,N_6397,N_5359);
xnor U13502 (N_13502,N_6243,N_6395);
and U13503 (N_13503,N_9002,N_5502);
and U13504 (N_13504,N_9378,N_7008);
and U13505 (N_13505,N_5388,N_5262);
nand U13506 (N_13506,N_9881,N_5312);
xor U13507 (N_13507,N_6939,N_8477);
and U13508 (N_13508,N_7823,N_6421);
nor U13509 (N_13509,N_6068,N_6820);
nor U13510 (N_13510,N_8126,N_6232);
and U13511 (N_13511,N_7163,N_6265);
or U13512 (N_13512,N_7347,N_5302);
and U13513 (N_13513,N_9425,N_8928);
xnor U13514 (N_13514,N_5032,N_5124);
nor U13515 (N_13515,N_5988,N_7806);
nor U13516 (N_13516,N_6290,N_5283);
nand U13517 (N_13517,N_8742,N_9248);
nor U13518 (N_13518,N_7928,N_9409);
nand U13519 (N_13519,N_8301,N_7296);
nor U13520 (N_13520,N_6450,N_8978);
nand U13521 (N_13521,N_5228,N_9605);
nand U13522 (N_13522,N_6332,N_5117);
nand U13523 (N_13523,N_5526,N_7292);
or U13524 (N_13524,N_8779,N_7951);
nor U13525 (N_13525,N_9464,N_5915);
or U13526 (N_13526,N_5776,N_9626);
or U13527 (N_13527,N_7148,N_8562);
xor U13528 (N_13528,N_8619,N_8311);
xor U13529 (N_13529,N_6364,N_9074);
or U13530 (N_13530,N_5198,N_8987);
nand U13531 (N_13531,N_8858,N_9779);
xnor U13532 (N_13532,N_8433,N_9534);
nand U13533 (N_13533,N_6270,N_7270);
or U13534 (N_13534,N_5324,N_8821);
or U13535 (N_13535,N_7233,N_9179);
nor U13536 (N_13536,N_8401,N_6710);
or U13537 (N_13537,N_7071,N_5341);
nand U13538 (N_13538,N_6853,N_8914);
or U13539 (N_13539,N_8672,N_8025);
and U13540 (N_13540,N_6050,N_9469);
and U13541 (N_13541,N_9713,N_7545);
nand U13542 (N_13542,N_9349,N_6713);
nand U13543 (N_13543,N_9853,N_9238);
nand U13544 (N_13544,N_7587,N_5387);
and U13545 (N_13545,N_6497,N_5079);
or U13546 (N_13546,N_5279,N_6004);
and U13547 (N_13547,N_9062,N_7716);
nand U13548 (N_13548,N_9388,N_5140);
or U13549 (N_13549,N_5305,N_9760);
and U13550 (N_13550,N_6914,N_9605);
or U13551 (N_13551,N_8591,N_7382);
nand U13552 (N_13552,N_7583,N_7372);
xor U13553 (N_13553,N_6006,N_9408);
and U13554 (N_13554,N_7796,N_8814);
nor U13555 (N_13555,N_7738,N_7788);
or U13556 (N_13556,N_5176,N_9589);
nor U13557 (N_13557,N_8240,N_5340);
nor U13558 (N_13558,N_5763,N_8331);
or U13559 (N_13559,N_9504,N_9982);
and U13560 (N_13560,N_7597,N_9251);
nor U13561 (N_13561,N_5466,N_5729);
xnor U13562 (N_13562,N_6367,N_6216);
or U13563 (N_13563,N_6197,N_8959);
or U13564 (N_13564,N_7532,N_7514);
nand U13565 (N_13565,N_8265,N_6888);
or U13566 (N_13566,N_8304,N_5561);
nand U13567 (N_13567,N_9398,N_5101);
nand U13568 (N_13568,N_8565,N_9376);
and U13569 (N_13569,N_7517,N_7821);
xor U13570 (N_13570,N_9938,N_9095);
nor U13571 (N_13571,N_7388,N_9698);
nor U13572 (N_13572,N_9649,N_6613);
nand U13573 (N_13573,N_6845,N_8458);
nor U13574 (N_13574,N_7742,N_9224);
or U13575 (N_13575,N_6319,N_5681);
and U13576 (N_13576,N_8213,N_5893);
nand U13577 (N_13577,N_6675,N_9943);
and U13578 (N_13578,N_7476,N_5554);
nor U13579 (N_13579,N_8404,N_7243);
xnor U13580 (N_13580,N_5776,N_7555);
nor U13581 (N_13581,N_6978,N_8092);
and U13582 (N_13582,N_9845,N_9022);
and U13583 (N_13583,N_9772,N_7858);
or U13584 (N_13584,N_7338,N_7788);
nor U13585 (N_13585,N_9868,N_6562);
and U13586 (N_13586,N_5334,N_5565);
nand U13587 (N_13587,N_5449,N_9475);
xor U13588 (N_13588,N_8916,N_9683);
nor U13589 (N_13589,N_5060,N_8554);
and U13590 (N_13590,N_7325,N_9775);
nor U13591 (N_13591,N_7030,N_6316);
xnor U13592 (N_13592,N_5802,N_9856);
or U13593 (N_13593,N_6620,N_6910);
or U13594 (N_13594,N_5623,N_7128);
or U13595 (N_13595,N_7685,N_6067);
xor U13596 (N_13596,N_8171,N_8615);
and U13597 (N_13597,N_6801,N_5598);
or U13598 (N_13598,N_7896,N_8905);
nand U13599 (N_13599,N_7463,N_5879);
or U13600 (N_13600,N_7839,N_7738);
xnor U13601 (N_13601,N_8738,N_9977);
and U13602 (N_13602,N_5306,N_9038);
nor U13603 (N_13603,N_7275,N_5314);
nor U13604 (N_13604,N_9395,N_9650);
xor U13605 (N_13605,N_8028,N_6688);
or U13606 (N_13606,N_9028,N_8598);
xnor U13607 (N_13607,N_7948,N_6484);
or U13608 (N_13608,N_5587,N_9943);
or U13609 (N_13609,N_9773,N_6898);
nand U13610 (N_13610,N_6578,N_6376);
and U13611 (N_13611,N_6020,N_9291);
nor U13612 (N_13612,N_7773,N_5832);
nand U13613 (N_13613,N_9350,N_7746);
nor U13614 (N_13614,N_9043,N_7310);
or U13615 (N_13615,N_8479,N_7299);
xnor U13616 (N_13616,N_8955,N_8086);
nand U13617 (N_13617,N_9729,N_7324);
or U13618 (N_13618,N_5438,N_6164);
nor U13619 (N_13619,N_6796,N_6615);
nand U13620 (N_13620,N_8204,N_6909);
nand U13621 (N_13621,N_5447,N_9316);
xor U13622 (N_13622,N_6280,N_5326);
xnor U13623 (N_13623,N_9603,N_9686);
xor U13624 (N_13624,N_8420,N_7495);
xnor U13625 (N_13625,N_6740,N_7300);
and U13626 (N_13626,N_7301,N_9354);
or U13627 (N_13627,N_7240,N_7690);
nand U13628 (N_13628,N_6778,N_5197);
nand U13629 (N_13629,N_7814,N_7461);
xor U13630 (N_13630,N_8336,N_6800);
nor U13631 (N_13631,N_7474,N_5752);
nand U13632 (N_13632,N_6847,N_5543);
xor U13633 (N_13633,N_8763,N_7829);
xor U13634 (N_13634,N_7750,N_9792);
and U13635 (N_13635,N_5430,N_8566);
nand U13636 (N_13636,N_7528,N_9393);
nand U13637 (N_13637,N_6153,N_7919);
nor U13638 (N_13638,N_6187,N_6812);
nand U13639 (N_13639,N_5668,N_8315);
nand U13640 (N_13640,N_5267,N_9440);
xor U13641 (N_13641,N_8407,N_5203);
nand U13642 (N_13642,N_8524,N_6721);
xor U13643 (N_13643,N_9738,N_5920);
or U13644 (N_13644,N_9778,N_7330);
xnor U13645 (N_13645,N_9738,N_9484);
xnor U13646 (N_13646,N_6016,N_6426);
and U13647 (N_13647,N_5615,N_7121);
or U13648 (N_13648,N_7962,N_5511);
and U13649 (N_13649,N_8813,N_5677);
nor U13650 (N_13650,N_6480,N_6281);
nor U13651 (N_13651,N_7894,N_9865);
nand U13652 (N_13652,N_7455,N_6522);
nand U13653 (N_13653,N_8436,N_7984);
xnor U13654 (N_13654,N_7065,N_9293);
or U13655 (N_13655,N_5239,N_9652);
or U13656 (N_13656,N_9102,N_9532);
or U13657 (N_13657,N_5680,N_5015);
or U13658 (N_13658,N_9202,N_7992);
xor U13659 (N_13659,N_7036,N_7325);
or U13660 (N_13660,N_7195,N_5964);
and U13661 (N_13661,N_5843,N_6672);
xor U13662 (N_13662,N_9541,N_8643);
xnor U13663 (N_13663,N_9634,N_9439);
xnor U13664 (N_13664,N_8800,N_8934);
xor U13665 (N_13665,N_6516,N_9586);
nand U13666 (N_13666,N_8201,N_6038);
nor U13667 (N_13667,N_8756,N_9408);
xnor U13668 (N_13668,N_5159,N_5647);
or U13669 (N_13669,N_7781,N_6923);
xor U13670 (N_13670,N_5201,N_5262);
and U13671 (N_13671,N_8548,N_9643);
nand U13672 (N_13672,N_8429,N_6401);
nor U13673 (N_13673,N_5561,N_6843);
nand U13674 (N_13674,N_8331,N_7679);
nand U13675 (N_13675,N_9906,N_9564);
and U13676 (N_13676,N_8623,N_7172);
nor U13677 (N_13677,N_6724,N_6245);
nor U13678 (N_13678,N_9557,N_5621);
xor U13679 (N_13679,N_5741,N_7065);
nand U13680 (N_13680,N_9162,N_9284);
and U13681 (N_13681,N_7434,N_9070);
nor U13682 (N_13682,N_7557,N_9380);
and U13683 (N_13683,N_7588,N_7208);
and U13684 (N_13684,N_9462,N_8592);
or U13685 (N_13685,N_9045,N_7412);
nor U13686 (N_13686,N_5457,N_8719);
xor U13687 (N_13687,N_8068,N_5845);
nor U13688 (N_13688,N_8502,N_5155);
and U13689 (N_13689,N_7980,N_9464);
nand U13690 (N_13690,N_8089,N_8616);
or U13691 (N_13691,N_9540,N_7951);
and U13692 (N_13692,N_6127,N_5182);
or U13693 (N_13693,N_9734,N_5786);
and U13694 (N_13694,N_9600,N_9419);
nor U13695 (N_13695,N_5627,N_6246);
xnor U13696 (N_13696,N_7594,N_5875);
xor U13697 (N_13697,N_6836,N_6258);
nor U13698 (N_13698,N_6369,N_5458);
and U13699 (N_13699,N_8380,N_9138);
nand U13700 (N_13700,N_7342,N_8328);
nor U13701 (N_13701,N_5406,N_6785);
and U13702 (N_13702,N_9457,N_5371);
and U13703 (N_13703,N_6657,N_8483);
and U13704 (N_13704,N_5786,N_9494);
nor U13705 (N_13705,N_9002,N_7116);
nand U13706 (N_13706,N_9790,N_8023);
nand U13707 (N_13707,N_5263,N_8697);
and U13708 (N_13708,N_5422,N_9650);
nand U13709 (N_13709,N_5151,N_5325);
and U13710 (N_13710,N_5811,N_7164);
and U13711 (N_13711,N_8737,N_8671);
or U13712 (N_13712,N_9229,N_7748);
nor U13713 (N_13713,N_8510,N_7968);
or U13714 (N_13714,N_8856,N_7692);
or U13715 (N_13715,N_7781,N_7394);
xor U13716 (N_13716,N_5477,N_6612);
nor U13717 (N_13717,N_9424,N_5973);
nor U13718 (N_13718,N_6412,N_6405);
or U13719 (N_13719,N_5384,N_7533);
and U13720 (N_13720,N_5220,N_9881);
or U13721 (N_13721,N_5103,N_6429);
nand U13722 (N_13722,N_8012,N_6516);
nor U13723 (N_13723,N_9560,N_8509);
xnor U13724 (N_13724,N_6217,N_7670);
and U13725 (N_13725,N_9386,N_9876);
or U13726 (N_13726,N_5298,N_9939);
or U13727 (N_13727,N_6465,N_6640);
xnor U13728 (N_13728,N_9358,N_8072);
nand U13729 (N_13729,N_9156,N_9869);
or U13730 (N_13730,N_6861,N_7895);
nor U13731 (N_13731,N_7024,N_9604);
nor U13732 (N_13732,N_9993,N_5148);
or U13733 (N_13733,N_5340,N_7928);
or U13734 (N_13734,N_6920,N_9451);
or U13735 (N_13735,N_8870,N_6820);
nand U13736 (N_13736,N_6793,N_7112);
or U13737 (N_13737,N_7743,N_8637);
xnor U13738 (N_13738,N_9494,N_7161);
and U13739 (N_13739,N_9235,N_5036);
and U13740 (N_13740,N_8600,N_6468);
nand U13741 (N_13741,N_7923,N_6805);
and U13742 (N_13742,N_5390,N_9151);
or U13743 (N_13743,N_7732,N_5419);
xor U13744 (N_13744,N_8719,N_6346);
nand U13745 (N_13745,N_7959,N_5123);
xnor U13746 (N_13746,N_8675,N_8824);
nand U13747 (N_13747,N_8057,N_8104);
or U13748 (N_13748,N_5680,N_9154);
nor U13749 (N_13749,N_8099,N_7305);
nor U13750 (N_13750,N_9430,N_6009);
or U13751 (N_13751,N_7489,N_7197);
nand U13752 (N_13752,N_8081,N_9276);
and U13753 (N_13753,N_8722,N_9870);
or U13754 (N_13754,N_5930,N_6715);
nand U13755 (N_13755,N_7372,N_9709);
or U13756 (N_13756,N_8538,N_9947);
or U13757 (N_13757,N_9190,N_8438);
and U13758 (N_13758,N_6087,N_7461);
xnor U13759 (N_13759,N_9092,N_6548);
and U13760 (N_13760,N_9651,N_5904);
xnor U13761 (N_13761,N_7589,N_7598);
or U13762 (N_13762,N_5769,N_5113);
xnor U13763 (N_13763,N_9643,N_8095);
and U13764 (N_13764,N_7294,N_6994);
xnor U13765 (N_13765,N_7337,N_5044);
nor U13766 (N_13766,N_7248,N_7218);
or U13767 (N_13767,N_9353,N_5470);
xnor U13768 (N_13768,N_5019,N_5981);
nor U13769 (N_13769,N_7593,N_6548);
nor U13770 (N_13770,N_7190,N_9317);
or U13771 (N_13771,N_9308,N_7737);
nor U13772 (N_13772,N_6329,N_6306);
and U13773 (N_13773,N_6425,N_6249);
and U13774 (N_13774,N_8879,N_6344);
or U13775 (N_13775,N_8784,N_9534);
and U13776 (N_13776,N_8864,N_8201);
nand U13777 (N_13777,N_9309,N_9555);
or U13778 (N_13778,N_7786,N_7243);
and U13779 (N_13779,N_6493,N_7049);
and U13780 (N_13780,N_5966,N_7642);
and U13781 (N_13781,N_9866,N_6966);
and U13782 (N_13782,N_7875,N_7550);
nor U13783 (N_13783,N_5118,N_7476);
xnor U13784 (N_13784,N_9271,N_7785);
nand U13785 (N_13785,N_8615,N_6678);
and U13786 (N_13786,N_7144,N_6781);
nand U13787 (N_13787,N_6904,N_8638);
xnor U13788 (N_13788,N_7380,N_9922);
or U13789 (N_13789,N_5308,N_7430);
and U13790 (N_13790,N_8315,N_6462);
nor U13791 (N_13791,N_5232,N_9536);
nor U13792 (N_13792,N_8532,N_8423);
nand U13793 (N_13793,N_9204,N_7351);
or U13794 (N_13794,N_6935,N_6658);
or U13795 (N_13795,N_7889,N_5846);
xnor U13796 (N_13796,N_7873,N_5469);
or U13797 (N_13797,N_5914,N_8640);
xor U13798 (N_13798,N_8606,N_9342);
or U13799 (N_13799,N_9748,N_9331);
or U13800 (N_13800,N_6402,N_8682);
nor U13801 (N_13801,N_9637,N_7266);
and U13802 (N_13802,N_8332,N_9483);
xor U13803 (N_13803,N_9402,N_5214);
nand U13804 (N_13804,N_6398,N_6911);
or U13805 (N_13805,N_5832,N_9081);
and U13806 (N_13806,N_8239,N_8855);
and U13807 (N_13807,N_7584,N_5558);
nor U13808 (N_13808,N_7343,N_9193);
xnor U13809 (N_13809,N_9397,N_7712);
and U13810 (N_13810,N_7044,N_6800);
nor U13811 (N_13811,N_6470,N_9785);
nand U13812 (N_13812,N_9688,N_6221);
nand U13813 (N_13813,N_9431,N_9596);
nand U13814 (N_13814,N_5180,N_5803);
nand U13815 (N_13815,N_7809,N_6934);
nand U13816 (N_13816,N_6931,N_9022);
nand U13817 (N_13817,N_8265,N_5716);
xnor U13818 (N_13818,N_9546,N_9422);
nand U13819 (N_13819,N_9321,N_9440);
nand U13820 (N_13820,N_6210,N_5397);
and U13821 (N_13821,N_9884,N_6779);
and U13822 (N_13822,N_5309,N_8020);
and U13823 (N_13823,N_8351,N_9693);
and U13824 (N_13824,N_6117,N_5423);
or U13825 (N_13825,N_5543,N_7202);
xnor U13826 (N_13826,N_8944,N_7215);
or U13827 (N_13827,N_6906,N_5727);
or U13828 (N_13828,N_5813,N_6236);
nor U13829 (N_13829,N_8674,N_5414);
or U13830 (N_13830,N_6428,N_5219);
and U13831 (N_13831,N_8626,N_7310);
or U13832 (N_13832,N_9670,N_8029);
xor U13833 (N_13833,N_8635,N_8952);
xnor U13834 (N_13834,N_5413,N_5510);
nand U13835 (N_13835,N_7274,N_8420);
nand U13836 (N_13836,N_9768,N_6000);
and U13837 (N_13837,N_8477,N_8651);
or U13838 (N_13838,N_9263,N_9417);
xor U13839 (N_13839,N_8562,N_7853);
nor U13840 (N_13840,N_7848,N_5001);
xnor U13841 (N_13841,N_9348,N_9971);
xor U13842 (N_13842,N_5476,N_5472);
xnor U13843 (N_13843,N_7395,N_7786);
nor U13844 (N_13844,N_5755,N_8591);
or U13845 (N_13845,N_9442,N_8189);
xor U13846 (N_13846,N_5473,N_6560);
or U13847 (N_13847,N_5559,N_8353);
or U13848 (N_13848,N_6017,N_5521);
nor U13849 (N_13849,N_8840,N_7860);
nor U13850 (N_13850,N_6921,N_8084);
and U13851 (N_13851,N_7130,N_5555);
or U13852 (N_13852,N_6463,N_7767);
xnor U13853 (N_13853,N_7198,N_7650);
nor U13854 (N_13854,N_6262,N_6112);
and U13855 (N_13855,N_9429,N_7491);
xnor U13856 (N_13856,N_7675,N_9420);
or U13857 (N_13857,N_6422,N_7516);
or U13858 (N_13858,N_5210,N_8512);
and U13859 (N_13859,N_5353,N_6200);
nor U13860 (N_13860,N_6816,N_5100);
nor U13861 (N_13861,N_5917,N_8295);
or U13862 (N_13862,N_5233,N_7974);
xnor U13863 (N_13863,N_5845,N_8746);
nor U13864 (N_13864,N_9550,N_5059);
xor U13865 (N_13865,N_6729,N_6333);
or U13866 (N_13866,N_7411,N_6924);
and U13867 (N_13867,N_7170,N_6164);
and U13868 (N_13868,N_6802,N_9541);
or U13869 (N_13869,N_9918,N_7208);
and U13870 (N_13870,N_6794,N_6623);
nand U13871 (N_13871,N_8154,N_6441);
xor U13872 (N_13872,N_5536,N_9470);
xor U13873 (N_13873,N_9451,N_9780);
nor U13874 (N_13874,N_5510,N_8168);
xor U13875 (N_13875,N_5032,N_9058);
xnor U13876 (N_13876,N_6452,N_7513);
nand U13877 (N_13877,N_5029,N_9445);
and U13878 (N_13878,N_7306,N_5557);
xor U13879 (N_13879,N_6733,N_6312);
xor U13880 (N_13880,N_8841,N_8130);
nand U13881 (N_13881,N_5871,N_9143);
nand U13882 (N_13882,N_7158,N_6610);
nor U13883 (N_13883,N_5504,N_7799);
nand U13884 (N_13884,N_6377,N_8063);
and U13885 (N_13885,N_7257,N_9323);
nand U13886 (N_13886,N_5396,N_6949);
nand U13887 (N_13887,N_9563,N_5460);
xor U13888 (N_13888,N_6188,N_6642);
nor U13889 (N_13889,N_5246,N_5573);
and U13890 (N_13890,N_9367,N_8912);
nor U13891 (N_13891,N_9475,N_9977);
nand U13892 (N_13892,N_6928,N_8815);
nor U13893 (N_13893,N_5315,N_7660);
or U13894 (N_13894,N_5172,N_6757);
and U13895 (N_13895,N_6562,N_8801);
or U13896 (N_13896,N_7924,N_5886);
xor U13897 (N_13897,N_8626,N_7760);
nand U13898 (N_13898,N_5620,N_8414);
or U13899 (N_13899,N_6155,N_8845);
nand U13900 (N_13900,N_9563,N_7574);
nand U13901 (N_13901,N_6129,N_7839);
or U13902 (N_13902,N_5281,N_7276);
xor U13903 (N_13903,N_7420,N_5695);
xnor U13904 (N_13904,N_9433,N_5615);
xor U13905 (N_13905,N_6186,N_7587);
nand U13906 (N_13906,N_9909,N_8557);
nor U13907 (N_13907,N_8277,N_9196);
and U13908 (N_13908,N_8036,N_6753);
and U13909 (N_13909,N_8521,N_8457);
or U13910 (N_13910,N_9145,N_8298);
and U13911 (N_13911,N_8525,N_5393);
or U13912 (N_13912,N_8774,N_7136);
and U13913 (N_13913,N_9420,N_8170);
nor U13914 (N_13914,N_6406,N_6405);
and U13915 (N_13915,N_5024,N_8717);
nor U13916 (N_13916,N_6732,N_7059);
or U13917 (N_13917,N_5006,N_5043);
or U13918 (N_13918,N_6350,N_8023);
and U13919 (N_13919,N_8041,N_8390);
and U13920 (N_13920,N_8931,N_6765);
or U13921 (N_13921,N_9749,N_5752);
or U13922 (N_13922,N_7561,N_9692);
and U13923 (N_13923,N_5111,N_5579);
nor U13924 (N_13924,N_6917,N_9525);
and U13925 (N_13925,N_6736,N_5556);
and U13926 (N_13926,N_6157,N_7960);
or U13927 (N_13927,N_5383,N_9553);
nand U13928 (N_13928,N_5449,N_9792);
xor U13929 (N_13929,N_7532,N_7055);
nand U13930 (N_13930,N_8904,N_7419);
and U13931 (N_13931,N_7536,N_8483);
nor U13932 (N_13932,N_5801,N_9152);
and U13933 (N_13933,N_5901,N_7478);
and U13934 (N_13934,N_5251,N_9561);
nor U13935 (N_13935,N_8333,N_5576);
or U13936 (N_13936,N_8297,N_6850);
and U13937 (N_13937,N_8665,N_8313);
and U13938 (N_13938,N_5647,N_9119);
xnor U13939 (N_13939,N_9143,N_9367);
or U13940 (N_13940,N_6967,N_7131);
xnor U13941 (N_13941,N_6732,N_9906);
nor U13942 (N_13942,N_8935,N_7250);
nand U13943 (N_13943,N_8293,N_5825);
xor U13944 (N_13944,N_5240,N_6659);
nor U13945 (N_13945,N_7153,N_6788);
xnor U13946 (N_13946,N_6175,N_6450);
xnor U13947 (N_13947,N_6399,N_7245);
nor U13948 (N_13948,N_5128,N_6694);
or U13949 (N_13949,N_9078,N_7063);
xnor U13950 (N_13950,N_9906,N_6080);
xnor U13951 (N_13951,N_9153,N_8690);
or U13952 (N_13952,N_6244,N_6545);
or U13953 (N_13953,N_5192,N_8305);
and U13954 (N_13954,N_8491,N_6666);
and U13955 (N_13955,N_8443,N_5807);
nand U13956 (N_13956,N_5797,N_5352);
nor U13957 (N_13957,N_7494,N_8362);
nor U13958 (N_13958,N_7913,N_8611);
or U13959 (N_13959,N_9817,N_9504);
nor U13960 (N_13960,N_7238,N_6046);
and U13961 (N_13961,N_6014,N_8719);
nor U13962 (N_13962,N_6312,N_5715);
xnor U13963 (N_13963,N_5317,N_7137);
nand U13964 (N_13964,N_5874,N_7909);
and U13965 (N_13965,N_9550,N_7748);
xor U13966 (N_13966,N_9901,N_6950);
nor U13967 (N_13967,N_9659,N_7319);
xor U13968 (N_13968,N_6581,N_5623);
nor U13969 (N_13969,N_8764,N_7312);
nand U13970 (N_13970,N_8652,N_6526);
xor U13971 (N_13971,N_8286,N_5802);
nor U13972 (N_13972,N_6959,N_8933);
nand U13973 (N_13973,N_9734,N_6544);
nor U13974 (N_13974,N_8374,N_5683);
nand U13975 (N_13975,N_9654,N_6018);
or U13976 (N_13976,N_5758,N_7985);
nand U13977 (N_13977,N_7410,N_8107);
xnor U13978 (N_13978,N_7602,N_5086);
xnor U13979 (N_13979,N_5377,N_6525);
xor U13980 (N_13980,N_8994,N_7625);
nor U13981 (N_13981,N_7065,N_7117);
and U13982 (N_13982,N_8044,N_5933);
or U13983 (N_13983,N_9741,N_9389);
and U13984 (N_13984,N_8488,N_7024);
or U13985 (N_13985,N_8541,N_8745);
or U13986 (N_13986,N_6162,N_8214);
or U13987 (N_13987,N_8876,N_6985);
xor U13988 (N_13988,N_8651,N_6124);
nand U13989 (N_13989,N_8656,N_8648);
and U13990 (N_13990,N_8117,N_7981);
or U13991 (N_13991,N_5881,N_6120);
xor U13992 (N_13992,N_8928,N_7772);
and U13993 (N_13993,N_9326,N_7405);
nor U13994 (N_13994,N_7466,N_8678);
xor U13995 (N_13995,N_7065,N_6900);
nor U13996 (N_13996,N_6735,N_8635);
xor U13997 (N_13997,N_5419,N_9722);
and U13998 (N_13998,N_9231,N_8648);
nor U13999 (N_13999,N_8894,N_7755);
nand U14000 (N_14000,N_9307,N_8686);
xor U14001 (N_14001,N_7054,N_7455);
nand U14002 (N_14002,N_9759,N_6440);
or U14003 (N_14003,N_8845,N_6434);
nand U14004 (N_14004,N_6646,N_7573);
nor U14005 (N_14005,N_5683,N_5551);
nand U14006 (N_14006,N_8629,N_6966);
or U14007 (N_14007,N_5126,N_9616);
nor U14008 (N_14008,N_7693,N_7372);
xnor U14009 (N_14009,N_6985,N_9477);
xnor U14010 (N_14010,N_6704,N_5289);
nor U14011 (N_14011,N_8894,N_7859);
nor U14012 (N_14012,N_8100,N_9681);
nor U14013 (N_14013,N_5040,N_7309);
nand U14014 (N_14014,N_5798,N_5767);
and U14015 (N_14015,N_5094,N_7610);
nor U14016 (N_14016,N_5965,N_6169);
nor U14017 (N_14017,N_9652,N_8439);
nor U14018 (N_14018,N_8640,N_9705);
or U14019 (N_14019,N_5472,N_5385);
nor U14020 (N_14020,N_5923,N_6552);
nor U14021 (N_14021,N_6402,N_9881);
xnor U14022 (N_14022,N_9959,N_8781);
xor U14023 (N_14023,N_5544,N_7652);
and U14024 (N_14024,N_6302,N_9800);
nor U14025 (N_14025,N_5381,N_5711);
nand U14026 (N_14026,N_7138,N_9050);
nor U14027 (N_14027,N_7272,N_6375);
or U14028 (N_14028,N_6418,N_7253);
and U14029 (N_14029,N_8313,N_5287);
nor U14030 (N_14030,N_5761,N_6068);
xor U14031 (N_14031,N_9953,N_8981);
nor U14032 (N_14032,N_8111,N_6962);
nand U14033 (N_14033,N_7851,N_9707);
or U14034 (N_14034,N_5439,N_9810);
xnor U14035 (N_14035,N_6072,N_8942);
nand U14036 (N_14036,N_8169,N_5909);
nand U14037 (N_14037,N_9084,N_7939);
or U14038 (N_14038,N_9374,N_8779);
nand U14039 (N_14039,N_8442,N_6823);
and U14040 (N_14040,N_6219,N_9380);
or U14041 (N_14041,N_6232,N_6189);
or U14042 (N_14042,N_8945,N_6184);
nor U14043 (N_14043,N_7339,N_7392);
or U14044 (N_14044,N_5469,N_7559);
and U14045 (N_14045,N_5196,N_5550);
and U14046 (N_14046,N_9155,N_8826);
nand U14047 (N_14047,N_9207,N_5211);
nand U14048 (N_14048,N_8943,N_8126);
nor U14049 (N_14049,N_7113,N_8962);
or U14050 (N_14050,N_7335,N_9195);
and U14051 (N_14051,N_6852,N_6794);
nand U14052 (N_14052,N_8334,N_9184);
and U14053 (N_14053,N_8187,N_6885);
nor U14054 (N_14054,N_5401,N_6492);
nand U14055 (N_14055,N_5770,N_8630);
nand U14056 (N_14056,N_7821,N_5530);
nand U14057 (N_14057,N_6718,N_8230);
xor U14058 (N_14058,N_7839,N_8153);
nand U14059 (N_14059,N_5176,N_6060);
xor U14060 (N_14060,N_6629,N_9291);
xor U14061 (N_14061,N_5727,N_8767);
and U14062 (N_14062,N_7291,N_7298);
xor U14063 (N_14063,N_8915,N_9346);
or U14064 (N_14064,N_7476,N_9203);
or U14065 (N_14065,N_5065,N_6057);
and U14066 (N_14066,N_9873,N_8091);
xor U14067 (N_14067,N_7661,N_8056);
xor U14068 (N_14068,N_5781,N_5694);
xnor U14069 (N_14069,N_9553,N_6740);
or U14070 (N_14070,N_7431,N_7292);
and U14071 (N_14071,N_5795,N_6267);
or U14072 (N_14072,N_6372,N_9946);
and U14073 (N_14073,N_9949,N_8499);
and U14074 (N_14074,N_7170,N_8852);
xnor U14075 (N_14075,N_6124,N_8891);
or U14076 (N_14076,N_9684,N_6333);
nand U14077 (N_14077,N_9909,N_6287);
and U14078 (N_14078,N_6595,N_7154);
and U14079 (N_14079,N_9305,N_9414);
and U14080 (N_14080,N_9657,N_8957);
xnor U14081 (N_14081,N_8921,N_5978);
and U14082 (N_14082,N_5974,N_7754);
nor U14083 (N_14083,N_9530,N_7162);
or U14084 (N_14084,N_8384,N_6399);
or U14085 (N_14085,N_5182,N_6653);
xor U14086 (N_14086,N_9294,N_8802);
nor U14087 (N_14087,N_7804,N_7025);
nand U14088 (N_14088,N_6901,N_8281);
xor U14089 (N_14089,N_6462,N_8376);
and U14090 (N_14090,N_9146,N_6139);
xor U14091 (N_14091,N_6657,N_7133);
nor U14092 (N_14092,N_5512,N_7879);
nand U14093 (N_14093,N_6731,N_9536);
nor U14094 (N_14094,N_6774,N_6972);
xor U14095 (N_14095,N_5683,N_5234);
nor U14096 (N_14096,N_9225,N_8001);
nor U14097 (N_14097,N_5088,N_6293);
and U14098 (N_14098,N_5555,N_8699);
nand U14099 (N_14099,N_7076,N_9826);
nor U14100 (N_14100,N_5567,N_6889);
and U14101 (N_14101,N_8572,N_8809);
or U14102 (N_14102,N_7403,N_6569);
xor U14103 (N_14103,N_6745,N_6037);
and U14104 (N_14104,N_7876,N_6122);
nor U14105 (N_14105,N_8750,N_9363);
nand U14106 (N_14106,N_7600,N_8311);
xnor U14107 (N_14107,N_7052,N_9337);
nor U14108 (N_14108,N_7422,N_8261);
or U14109 (N_14109,N_8229,N_6968);
nand U14110 (N_14110,N_5233,N_8352);
or U14111 (N_14111,N_6602,N_5174);
or U14112 (N_14112,N_9533,N_8050);
xor U14113 (N_14113,N_9191,N_8975);
nor U14114 (N_14114,N_7302,N_7184);
nor U14115 (N_14115,N_8351,N_7579);
xnor U14116 (N_14116,N_9886,N_5814);
and U14117 (N_14117,N_5877,N_6088);
nor U14118 (N_14118,N_7862,N_9055);
xnor U14119 (N_14119,N_8948,N_5487);
or U14120 (N_14120,N_8038,N_8299);
nor U14121 (N_14121,N_9628,N_8764);
or U14122 (N_14122,N_8513,N_8529);
nor U14123 (N_14123,N_6519,N_6049);
xnor U14124 (N_14124,N_7371,N_7380);
or U14125 (N_14125,N_7999,N_9934);
xnor U14126 (N_14126,N_6989,N_7825);
and U14127 (N_14127,N_6727,N_8142);
or U14128 (N_14128,N_7461,N_9668);
xor U14129 (N_14129,N_7881,N_8442);
and U14130 (N_14130,N_7780,N_9797);
nand U14131 (N_14131,N_6065,N_5435);
xor U14132 (N_14132,N_9059,N_7346);
nor U14133 (N_14133,N_9065,N_8572);
xor U14134 (N_14134,N_9597,N_7907);
xor U14135 (N_14135,N_6174,N_9472);
nand U14136 (N_14136,N_6392,N_6389);
or U14137 (N_14137,N_9086,N_8588);
nand U14138 (N_14138,N_8056,N_6353);
or U14139 (N_14139,N_6687,N_8321);
xnor U14140 (N_14140,N_7223,N_5095);
or U14141 (N_14141,N_5585,N_6936);
or U14142 (N_14142,N_5368,N_6826);
and U14143 (N_14143,N_6448,N_6185);
or U14144 (N_14144,N_7856,N_8497);
nand U14145 (N_14145,N_6215,N_7490);
xor U14146 (N_14146,N_9049,N_6902);
or U14147 (N_14147,N_5539,N_9462);
nand U14148 (N_14148,N_6907,N_7037);
xor U14149 (N_14149,N_8718,N_6315);
and U14150 (N_14150,N_8930,N_7364);
xor U14151 (N_14151,N_5455,N_9183);
or U14152 (N_14152,N_8379,N_5789);
xnor U14153 (N_14153,N_8419,N_8724);
xnor U14154 (N_14154,N_5054,N_6576);
or U14155 (N_14155,N_9729,N_6764);
nor U14156 (N_14156,N_7169,N_9682);
or U14157 (N_14157,N_5215,N_8620);
xnor U14158 (N_14158,N_6965,N_7825);
nand U14159 (N_14159,N_7308,N_8111);
xor U14160 (N_14160,N_8220,N_7732);
nor U14161 (N_14161,N_8096,N_9810);
or U14162 (N_14162,N_7391,N_9088);
nand U14163 (N_14163,N_9506,N_5580);
nor U14164 (N_14164,N_8454,N_8559);
nor U14165 (N_14165,N_9275,N_8096);
nor U14166 (N_14166,N_6900,N_7229);
nor U14167 (N_14167,N_7796,N_6279);
nand U14168 (N_14168,N_8413,N_6395);
nor U14169 (N_14169,N_7142,N_9021);
xor U14170 (N_14170,N_5185,N_6315);
nand U14171 (N_14171,N_8366,N_6197);
nand U14172 (N_14172,N_7482,N_7004);
nand U14173 (N_14173,N_5002,N_8289);
and U14174 (N_14174,N_8926,N_7275);
or U14175 (N_14175,N_7760,N_6055);
and U14176 (N_14176,N_9933,N_8566);
or U14177 (N_14177,N_7215,N_5410);
or U14178 (N_14178,N_9911,N_5387);
xor U14179 (N_14179,N_7422,N_6869);
and U14180 (N_14180,N_9645,N_5543);
nand U14181 (N_14181,N_9473,N_8293);
and U14182 (N_14182,N_8416,N_7983);
nor U14183 (N_14183,N_6286,N_8450);
xor U14184 (N_14184,N_9808,N_7396);
xnor U14185 (N_14185,N_9462,N_9344);
nor U14186 (N_14186,N_8485,N_5820);
nor U14187 (N_14187,N_9754,N_7542);
nor U14188 (N_14188,N_6383,N_7654);
or U14189 (N_14189,N_7623,N_7113);
or U14190 (N_14190,N_6871,N_7115);
or U14191 (N_14191,N_5908,N_5017);
nand U14192 (N_14192,N_6260,N_8859);
xor U14193 (N_14193,N_7127,N_7990);
or U14194 (N_14194,N_7282,N_6096);
xnor U14195 (N_14195,N_7484,N_7901);
nor U14196 (N_14196,N_7612,N_8049);
xor U14197 (N_14197,N_9105,N_8226);
xor U14198 (N_14198,N_5029,N_6366);
nand U14199 (N_14199,N_9404,N_7933);
xor U14200 (N_14200,N_5966,N_6270);
xnor U14201 (N_14201,N_6366,N_9514);
nand U14202 (N_14202,N_9082,N_9295);
and U14203 (N_14203,N_6534,N_7434);
or U14204 (N_14204,N_8213,N_8573);
and U14205 (N_14205,N_5200,N_8403);
and U14206 (N_14206,N_7415,N_5249);
nor U14207 (N_14207,N_7067,N_7755);
nand U14208 (N_14208,N_6981,N_5130);
and U14209 (N_14209,N_7610,N_5593);
and U14210 (N_14210,N_5178,N_7468);
nor U14211 (N_14211,N_9675,N_7158);
nand U14212 (N_14212,N_8155,N_8768);
or U14213 (N_14213,N_7615,N_6373);
nand U14214 (N_14214,N_7103,N_9024);
xor U14215 (N_14215,N_7133,N_5765);
nor U14216 (N_14216,N_6222,N_5174);
nor U14217 (N_14217,N_9221,N_7018);
or U14218 (N_14218,N_8627,N_7845);
or U14219 (N_14219,N_8566,N_5461);
nand U14220 (N_14220,N_5989,N_8952);
xor U14221 (N_14221,N_7358,N_6336);
xnor U14222 (N_14222,N_8963,N_6814);
nor U14223 (N_14223,N_7304,N_5960);
nor U14224 (N_14224,N_9499,N_5926);
and U14225 (N_14225,N_5552,N_8084);
xnor U14226 (N_14226,N_6529,N_7879);
or U14227 (N_14227,N_6766,N_8540);
nor U14228 (N_14228,N_6197,N_5735);
and U14229 (N_14229,N_6211,N_9188);
or U14230 (N_14230,N_7121,N_8529);
and U14231 (N_14231,N_9654,N_5795);
xnor U14232 (N_14232,N_8991,N_6115);
or U14233 (N_14233,N_7328,N_5940);
nand U14234 (N_14234,N_9349,N_6271);
and U14235 (N_14235,N_5067,N_8014);
nand U14236 (N_14236,N_7403,N_8206);
nor U14237 (N_14237,N_9723,N_8881);
xnor U14238 (N_14238,N_9509,N_8560);
nor U14239 (N_14239,N_8737,N_5237);
xor U14240 (N_14240,N_8840,N_6725);
or U14241 (N_14241,N_5666,N_8696);
xor U14242 (N_14242,N_5340,N_6605);
nor U14243 (N_14243,N_5253,N_9066);
nand U14244 (N_14244,N_6426,N_5462);
nor U14245 (N_14245,N_5103,N_6806);
nand U14246 (N_14246,N_6629,N_9680);
nand U14247 (N_14247,N_8250,N_5096);
nand U14248 (N_14248,N_9168,N_6171);
or U14249 (N_14249,N_9447,N_7186);
xnor U14250 (N_14250,N_6498,N_6983);
nor U14251 (N_14251,N_7380,N_7263);
nand U14252 (N_14252,N_6777,N_7849);
nand U14253 (N_14253,N_5445,N_5999);
and U14254 (N_14254,N_9722,N_5960);
nor U14255 (N_14255,N_9075,N_9344);
and U14256 (N_14256,N_5242,N_7234);
and U14257 (N_14257,N_6319,N_7985);
nor U14258 (N_14258,N_8582,N_5664);
or U14259 (N_14259,N_8856,N_7722);
nor U14260 (N_14260,N_5234,N_7996);
xor U14261 (N_14261,N_7105,N_8414);
and U14262 (N_14262,N_8803,N_9106);
xor U14263 (N_14263,N_7829,N_6584);
or U14264 (N_14264,N_6513,N_8317);
or U14265 (N_14265,N_7222,N_9182);
and U14266 (N_14266,N_7702,N_7182);
or U14267 (N_14267,N_8730,N_8043);
nand U14268 (N_14268,N_6845,N_6033);
and U14269 (N_14269,N_9391,N_6430);
nand U14270 (N_14270,N_6342,N_9707);
nand U14271 (N_14271,N_5984,N_7925);
nand U14272 (N_14272,N_5694,N_6545);
nor U14273 (N_14273,N_5698,N_9727);
or U14274 (N_14274,N_6392,N_7649);
and U14275 (N_14275,N_8562,N_8470);
or U14276 (N_14276,N_7510,N_7080);
nand U14277 (N_14277,N_7636,N_7332);
xnor U14278 (N_14278,N_9723,N_8035);
xor U14279 (N_14279,N_5825,N_8712);
or U14280 (N_14280,N_7065,N_7336);
and U14281 (N_14281,N_7556,N_6692);
and U14282 (N_14282,N_9839,N_8568);
xor U14283 (N_14283,N_6870,N_7560);
nor U14284 (N_14284,N_5372,N_5935);
nand U14285 (N_14285,N_8459,N_5588);
or U14286 (N_14286,N_8130,N_6610);
nand U14287 (N_14287,N_6881,N_7384);
or U14288 (N_14288,N_5740,N_9510);
or U14289 (N_14289,N_5851,N_9717);
nor U14290 (N_14290,N_8491,N_6856);
nor U14291 (N_14291,N_8227,N_7316);
nor U14292 (N_14292,N_5110,N_6246);
xnor U14293 (N_14293,N_7454,N_5818);
and U14294 (N_14294,N_8387,N_6176);
xor U14295 (N_14295,N_8495,N_5628);
nor U14296 (N_14296,N_7629,N_8950);
nand U14297 (N_14297,N_7451,N_7582);
nand U14298 (N_14298,N_5264,N_6616);
and U14299 (N_14299,N_6971,N_6554);
and U14300 (N_14300,N_5465,N_7042);
nand U14301 (N_14301,N_9302,N_6286);
and U14302 (N_14302,N_5782,N_8527);
nor U14303 (N_14303,N_9664,N_9550);
nor U14304 (N_14304,N_9506,N_8782);
and U14305 (N_14305,N_8629,N_7978);
or U14306 (N_14306,N_8509,N_9962);
nor U14307 (N_14307,N_8847,N_9598);
nand U14308 (N_14308,N_9593,N_9319);
nand U14309 (N_14309,N_5435,N_8410);
or U14310 (N_14310,N_6418,N_5462);
or U14311 (N_14311,N_8611,N_8773);
or U14312 (N_14312,N_8974,N_5441);
nand U14313 (N_14313,N_9917,N_7604);
nor U14314 (N_14314,N_7842,N_8086);
and U14315 (N_14315,N_7254,N_6735);
and U14316 (N_14316,N_6974,N_6202);
or U14317 (N_14317,N_8159,N_6594);
xnor U14318 (N_14318,N_5444,N_5030);
or U14319 (N_14319,N_6195,N_5659);
xnor U14320 (N_14320,N_7370,N_7778);
nand U14321 (N_14321,N_7578,N_7136);
nor U14322 (N_14322,N_9996,N_8612);
xor U14323 (N_14323,N_5694,N_5058);
and U14324 (N_14324,N_9847,N_5194);
xor U14325 (N_14325,N_5632,N_9949);
and U14326 (N_14326,N_5306,N_8861);
nand U14327 (N_14327,N_9123,N_5737);
nand U14328 (N_14328,N_5488,N_6490);
nor U14329 (N_14329,N_8036,N_6946);
nor U14330 (N_14330,N_8568,N_6509);
nor U14331 (N_14331,N_6698,N_9970);
nor U14332 (N_14332,N_6981,N_6747);
or U14333 (N_14333,N_7843,N_6609);
nand U14334 (N_14334,N_5710,N_7063);
and U14335 (N_14335,N_6787,N_8424);
xnor U14336 (N_14336,N_7748,N_7148);
nand U14337 (N_14337,N_5220,N_7076);
and U14338 (N_14338,N_5804,N_6049);
or U14339 (N_14339,N_9770,N_8242);
and U14340 (N_14340,N_7995,N_6993);
and U14341 (N_14341,N_7725,N_8453);
and U14342 (N_14342,N_9681,N_5320);
nand U14343 (N_14343,N_6906,N_6791);
nand U14344 (N_14344,N_9268,N_6553);
nand U14345 (N_14345,N_8265,N_9940);
xnor U14346 (N_14346,N_8167,N_6872);
xor U14347 (N_14347,N_7327,N_8604);
nand U14348 (N_14348,N_9104,N_9796);
or U14349 (N_14349,N_8727,N_9050);
nand U14350 (N_14350,N_5459,N_5664);
xnor U14351 (N_14351,N_8903,N_6960);
nand U14352 (N_14352,N_5849,N_9856);
xnor U14353 (N_14353,N_6871,N_5016);
nor U14354 (N_14354,N_9053,N_5865);
or U14355 (N_14355,N_8841,N_7863);
nor U14356 (N_14356,N_6009,N_8159);
nand U14357 (N_14357,N_7039,N_5787);
nand U14358 (N_14358,N_8487,N_6311);
and U14359 (N_14359,N_8354,N_7206);
nor U14360 (N_14360,N_7925,N_6499);
or U14361 (N_14361,N_7328,N_9430);
and U14362 (N_14362,N_8422,N_8379);
nand U14363 (N_14363,N_5503,N_9859);
nor U14364 (N_14364,N_7225,N_9050);
nand U14365 (N_14365,N_6721,N_7604);
xnor U14366 (N_14366,N_5571,N_7564);
nor U14367 (N_14367,N_7514,N_7766);
nand U14368 (N_14368,N_5194,N_5340);
nand U14369 (N_14369,N_7338,N_5867);
xor U14370 (N_14370,N_8377,N_6200);
or U14371 (N_14371,N_5932,N_9735);
nand U14372 (N_14372,N_6668,N_7699);
nand U14373 (N_14373,N_9483,N_7256);
nand U14374 (N_14374,N_6946,N_5436);
nor U14375 (N_14375,N_7809,N_8746);
and U14376 (N_14376,N_7900,N_8972);
or U14377 (N_14377,N_9379,N_5477);
or U14378 (N_14378,N_6864,N_5369);
and U14379 (N_14379,N_6190,N_7050);
xor U14380 (N_14380,N_5078,N_9942);
xnor U14381 (N_14381,N_7492,N_5140);
and U14382 (N_14382,N_6352,N_8171);
nand U14383 (N_14383,N_9631,N_6450);
nand U14384 (N_14384,N_5976,N_6353);
xnor U14385 (N_14385,N_7928,N_8459);
xor U14386 (N_14386,N_7600,N_7661);
xor U14387 (N_14387,N_6404,N_5060);
or U14388 (N_14388,N_7627,N_6324);
nor U14389 (N_14389,N_6109,N_6997);
xor U14390 (N_14390,N_5411,N_9179);
or U14391 (N_14391,N_5958,N_6527);
and U14392 (N_14392,N_8370,N_7279);
nand U14393 (N_14393,N_5884,N_8243);
xnor U14394 (N_14394,N_6516,N_7134);
nor U14395 (N_14395,N_6846,N_5688);
xnor U14396 (N_14396,N_5358,N_5399);
xnor U14397 (N_14397,N_6999,N_8431);
nor U14398 (N_14398,N_7888,N_8957);
and U14399 (N_14399,N_8644,N_6356);
nor U14400 (N_14400,N_8457,N_6678);
xor U14401 (N_14401,N_8844,N_9844);
nand U14402 (N_14402,N_8936,N_9455);
nand U14403 (N_14403,N_5913,N_7296);
nand U14404 (N_14404,N_5085,N_6523);
xor U14405 (N_14405,N_6059,N_9628);
and U14406 (N_14406,N_7851,N_8117);
xor U14407 (N_14407,N_5631,N_6653);
nor U14408 (N_14408,N_9084,N_6441);
xor U14409 (N_14409,N_8166,N_6711);
and U14410 (N_14410,N_9898,N_5621);
nand U14411 (N_14411,N_5652,N_5798);
nor U14412 (N_14412,N_8951,N_8956);
nand U14413 (N_14413,N_6706,N_9998);
xor U14414 (N_14414,N_8133,N_7648);
nor U14415 (N_14415,N_7755,N_8188);
xnor U14416 (N_14416,N_9897,N_8560);
or U14417 (N_14417,N_7109,N_7168);
xor U14418 (N_14418,N_8331,N_9489);
xor U14419 (N_14419,N_6787,N_8301);
xor U14420 (N_14420,N_5249,N_9102);
and U14421 (N_14421,N_8209,N_7679);
nor U14422 (N_14422,N_9727,N_9515);
or U14423 (N_14423,N_9009,N_8804);
and U14424 (N_14424,N_6618,N_5513);
nand U14425 (N_14425,N_5869,N_9066);
nand U14426 (N_14426,N_9318,N_7181);
nor U14427 (N_14427,N_8704,N_7856);
or U14428 (N_14428,N_5256,N_5542);
xor U14429 (N_14429,N_7901,N_9891);
xor U14430 (N_14430,N_9325,N_8891);
nor U14431 (N_14431,N_8877,N_7513);
nand U14432 (N_14432,N_8178,N_7661);
or U14433 (N_14433,N_6694,N_7666);
and U14434 (N_14434,N_5038,N_8524);
nand U14435 (N_14435,N_9829,N_9286);
or U14436 (N_14436,N_5358,N_5187);
and U14437 (N_14437,N_8939,N_9646);
xor U14438 (N_14438,N_8722,N_5633);
and U14439 (N_14439,N_6151,N_8805);
nor U14440 (N_14440,N_8801,N_5518);
or U14441 (N_14441,N_8189,N_5352);
nand U14442 (N_14442,N_5750,N_6851);
nand U14443 (N_14443,N_7352,N_6076);
xor U14444 (N_14444,N_7472,N_5436);
xor U14445 (N_14445,N_9113,N_9920);
or U14446 (N_14446,N_6729,N_5705);
or U14447 (N_14447,N_8224,N_7145);
nor U14448 (N_14448,N_8965,N_9445);
xnor U14449 (N_14449,N_9247,N_7012);
or U14450 (N_14450,N_5361,N_8381);
xnor U14451 (N_14451,N_7074,N_6923);
and U14452 (N_14452,N_5290,N_9165);
xnor U14453 (N_14453,N_5963,N_7935);
and U14454 (N_14454,N_6521,N_6994);
or U14455 (N_14455,N_8720,N_9637);
xnor U14456 (N_14456,N_5670,N_9601);
nor U14457 (N_14457,N_7092,N_7876);
xor U14458 (N_14458,N_9035,N_5653);
nand U14459 (N_14459,N_8736,N_8677);
or U14460 (N_14460,N_9864,N_7169);
nor U14461 (N_14461,N_5552,N_6663);
or U14462 (N_14462,N_7386,N_6936);
xnor U14463 (N_14463,N_5237,N_8476);
nand U14464 (N_14464,N_9849,N_9082);
nand U14465 (N_14465,N_5297,N_7793);
xnor U14466 (N_14466,N_8674,N_7734);
xnor U14467 (N_14467,N_8461,N_7915);
or U14468 (N_14468,N_5604,N_8228);
nand U14469 (N_14469,N_7860,N_8584);
and U14470 (N_14470,N_8083,N_5146);
nor U14471 (N_14471,N_9496,N_7093);
and U14472 (N_14472,N_6965,N_8393);
xnor U14473 (N_14473,N_6914,N_9897);
nand U14474 (N_14474,N_5780,N_8170);
and U14475 (N_14475,N_6863,N_7488);
or U14476 (N_14476,N_5200,N_6058);
nand U14477 (N_14477,N_6153,N_5518);
xor U14478 (N_14478,N_8789,N_7028);
xor U14479 (N_14479,N_9813,N_5620);
xnor U14480 (N_14480,N_6680,N_7009);
and U14481 (N_14481,N_9937,N_9601);
or U14482 (N_14482,N_5175,N_7851);
nand U14483 (N_14483,N_5737,N_8855);
xnor U14484 (N_14484,N_6969,N_6721);
xnor U14485 (N_14485,N_9686,N_9465);
xor U14486 (N_14486,N_8891,N_7486);
or U14487 (N_14487,N_6126,N_6723);
or U14488 (N_14488,N_9798,N_8091);
nand U14489 (N_14489,N_9087,N_5373);
nor U14490 (N_14490,N_9639,N_8848);
and U14491 (N_14491,N_9042,N_7395);
or U14492 (N_14492,N_5988,N_5123);
or U14493 (N_14493,N_9678,N_6385);
nor U14494 (N_14494,N_5554,N_7955);
nor U14495 (N_14495,N_7580,N_9059);
xnor U14496 (N_14496,N_6186,N_5017);
and U14497 (N_14497,N_7006,N_8804);
nor U14498 (N_14498,N_5083,N_8929);
nor U14499 (N_14499,N_6137,N_9917);
and U14500 (N_14500,N_7333,N_5962);
nor U14501 (N_14501,N_9049,N_8966);
and U14502 (N_14502,N_8327,N_9891);
nor U14503 (N_14503,N_7406,N_9503);
or U14504 (N_14504,N_5948,N_7108);
nor U14505 (N_14505,N_9832,N_7753);
nor U14506 (N_14506,N_8804,N_6716);
and U14507 (N_14507,N_9889,N_8901);
nor U14508 (N_14508,N_9755,N_7708);
and U14509 (N_14509,N_7258,N_5840);
or U14510 (N_14510,N_5102,N_7130);
nand U14511 (N_14511,N_9880,N_7751);
nor U14512 (N_14512,N_6188,N_6544);
nor U14513 (N_14513,N_6235,N_5607);
nand U14514 (N_14514,N_5715,N_9900);
or U14515 (N_14515,N_6361,N_5713);
xnor U14516 (N_14516,N_6024,N_8788);
and U14517 (N_14517,N_6723,N_7265);
nor U14518 (N_14518,N_8068,N_6715);
nand U14519 (N_14519,N_7150,N_9367);
nand U14520 (N_14520,N_8012,N_5906);
and U14521 (N_14521,N_6275,N_9985);
xor U14522 (N_14522,N_5925,N_9847);
nand U14523 (N_14523,N_5138,N_5967);
and U14524 (N_14524,N_9781,N_9764);
or U14525 (N_14525,N_8350,N_8157);
nor U14526 (N_14526,N_5318,N_9439);
or U14527 (N_14527,N_7549,N_7623);
nand U14528 (N_14528,N_6666,N_7057);
or U14529 (N_14529,N_7869,N_8193);
or U14530 (N_14530,N_9199,N_7430);
nand U14531 (N_14531,N_8020,N_7632);
or U14532 (N_14532,N_5213,N_5642);
or U14533 (N_14533,N_8745,N_9317);
or U14534 (N_14534,N_5228,N_7184);
nor U14535 (N_14535,N_6303,N_8867);
and U14536 (N_14536,N_8073,N_6613);
nor U14537 (N_14537,N_5362,N_9391);
xor U14538 (N_14538,N_5775,N_7429);
nand U14539 (N_14539,N_9434,N_5570);
or U14540 (N_14540,N_5663,N_7047);
nand U14541 (N_14541,N_9639,N_9518);
and U14542 (N_14542,N_6272,N_7051);
nor U14543 (N_14543,N_9960,N_8836);
xor U14544 (N_14544,N_7671,N_5916);
or U14545 (N_14545,N_5023,N_8864);
xor U14546 (N_14546,N_6083,N_9859);
nor U14547 (N_14547,N_8416,N_7406);
nor U14548 (N_14548,N_7546,N_8433);
nand U14549 (N_14549,N_7674,N_8969);
nand U14550 (N_14550,N_8891,N_7744);
nor U14551 (N_14551,N_8268,N_6118);
xor U14552 (N_14552,N_9392,N_7603);
nand U14553 (N_14553,N_7815,N_7864);
xnor U14554 (N_14554,N_9864,N_5219);
and U14555 (N_14555,N_8004,N_8119);
or U14556 (N_14556,N_7921,N_9251);
and U14557 (N_14557,N_9098,N_7019);
xor U14558 (N_14558,N_5953,N_9702);
and U14559 (N_14559,N_7746,N_6791);
nor U14560 (N_14560,N_9793,N_8789);
and U14561 (N_14561,N_8038,N_8694);
nand U14562 (N_14562,N_7004,N_6248);
nand U14563 (N_14563,N_6499,N_8267);
nor U14564 (N_14564,N_8613,N_8492);
and U14565 (N_14565,N_9710,N_9749);
or U14566 (N_14566,N_9469,N_7969);
and U14567 (N_14567,N_5764,N_7262);
and U14568 (N_14568,N_5352,N_5056);
and U14569 (N_14569,N_6627,N_8645);
nand U14570 (N_14570,N_9026,N_8667);
and U14571 (N_14571,N_8400,N_8789);
xor U14572 (N_14572,N_6015,N_7153);
xor U14573 (N_14573,N_8752,N_9355);
nand U14574 (N_14574,N_8675,N_6790);
or U14575 (N_14575,N_5541,N_7603);
and U14576 (N_14576,N_5909,N_9384);
nor U14577 (N_14577,N_9244,N_6147);
nor U14578 (N_14578,N_8396,N_6585);
and U14579 (N_14579,N_5586,N_9203);
and U14580 (N_14580,N_7014,N_8162);
and U14581 (N_14581,N_5256,N_6694);
nor U14582 (N_14582,N_5096,N_6469);
nand U14583 (N_14583,N_5604,N_7754);
nand U14584 (N_14584,N_5261,N_5742);
nand U14585 (N_14585,N_6260,N_5718);
and U14586 (N_14586,N_5348,N_5086);
xor U14587 (N_14587,N_9559,N_8866);
and U14588 (N_14588,N_7597,N_5690);
xor U14589 (N_14589,N_5206,N_6596);
and U14590 (N_14590,N_9004,N_9729);
or U14591 (N_14591,N_9343,N_8563);
and U14592 (N_14592,N_6954,N_5062);
xor U14593 (N_14593,N_5687,N_6950);
nor U14594 (N_14594,N_6494,N_6253);
nor U14595 (N_14595,N_8587,N_6522);
xnor U14596 (N_14596,N_7124,N_8824);
nand U14597 (N_14597,N_5615,N_7680);
nor U14598 (N_14598,N_8931,N_6591);
nor U14599 (N_14599,N_6703,N_5268);
and U14600 (N_14600,N_5746,N_7322);
nor U14601 (N_14601,N_5580,N_5329);
nand U14602 (N_14602,N_7664,N_7356);
and U14603 (N_14603,N_9874,N_8229);
nor U14604 (N_14604,N_6041,N_8138);
nand U14605 (N_14605,N_6119,N_8340);
xnor U14606 (N_14606,N_8724,N_7864);
or U14607 (N_14607,N_9690,N_5306);
and U14608 (N_14608,N_8052,N_9747);
xnor U14609 (N_14609,N_9603,N_8527);
nor U14610 (N_14610,N_8295,N_6612);
or U14611 (N_14611,N_7711,N_9822);
or U14612 (N_14612,N_9883,N_5170);
and U14613 (N_14613,N_5811,N_6818);
nand U14614 (N_14614,N_8022,N_5143);
xor U14615 (N_14615,N_8987,N_5453);
nand U14616 (N_14616,N_9983,N_9280);
nor U14617 (N_14617,N_9486,N_6970);
xnor U14618 (N_14618,N_6295,N_7940);
and U14619 (N_14619,N_7105,N_7688);
and U14620 (N_14620,N_7801,N_8903);
xor U14621 (N_14621,N_7730,N_8963);
nand U14622 (N_14622,N_8891,N_7346);
nor U14623 (N_14623,N_9697,N_8061);
xnor U14624 (N_14624,N_6304,N_6257);
or U14625 (N_14625,N_8178,N_9507);
and U14626 (N_14626,N_9577,N_5786);
or U14627 (N_14627,N_7145,N_6883);
nor U14628 (N_14628,N_5204,N_9529);
nor U14629 (N_14629,N_7692,N_8308);
or U14630 (N_14630,N_7082,N_8603);
nand U14631 (N_14631,N_7859,N_7793);
or U14632 (N_14632,N_7299,N_5034);
nor U14633 (N_14633,N_6429,N_8510);
and U14634 (N_14634,N_5869,N_9932);
nor U14635 (N_14635,N_8165,N_5596);
xnor U14636 (N_14636,N_8583,N_7477);
or U14637 (N_14637,N_8507,N_9793);
nor U14638 (N_14638,N_6640,N_9321);
or U14639 (N_14639,N_9842,N_8821);
and U14640 (N_14640,N_6078,N_8429);
or U14641 (N_14641,N_8329,N_5243);
or U14642 (N_14642,N_6036,N_6235);
or U14643 (N_14643,N_5792,N_6433);
and U14644 (N_14644,N_7144,N_8495);
and U14645 (N_14645,N_8469,N_6377);
nor U14646 (N_14646,N_8603,N_8021);
xnor U14647 (N_14647,N_9744,N_6134);
nor U14648 (N_14648,N_6172,N_9553);
and U14649 (N_14649,N_7111,N_9465);
xor U14650 (N_14650,N_6334,N_5990);
nand U14651 (N_14651,N_7231,N_6809);
nand U14652 (N_14652,N_5529,N_7145);
and U14653 (N_14653,N_6452,N_6391);
nor U14654 (N_14654,N_8196,N_7840);
and U14655 (N_14655,N_6162,N_6335);
nand U14656 (N_14656,N_6022,N_9806);
and U14657 (N_14657,N_5915,N_8777);
nand U14658 (N_14658,N_7730,N_9024);
and U14659 (N_14659,N_7121,N_8669);
xor U14660 (N_14660,N_7129,N_7287);
nor U14661 (N_14661,N_6921,N_8448);
or U14662 (N_14662,N_7527,N_5487);
nand U14663 (N_14663,N_8970,N_8499);
or U14664 (N_14664,N_9424,N_6511);
nand U14665 (N_14665,N_9919,N_9537);
nor U14666 (N_14666,N_8408,N_6602);
nand U14667 (N_14667,N_9783,N_8377);
or U14668 (N_14668,N_7313,N_9759);
and U14669 (N_14669,N_8721,N_5349);
xor U14670 (N_14670,N_8891,N_5211);
nor U14671 (N_14671,N_8711,N_8271);
and U14672 (N_14672,N_6881,N_5648);
and U14673 (N_14673,N_7368,N_6166);
nor U14674 (N_14674,N_8606,N_8076);
and U14675 (N_14675,N_9507,N_7744);
nor U14676 (N_14676,N_7315,N_8662);
and U14677 (N_14677,N_5332,N_5613);
nor U14678 (N_14678,N_8956,N_6825);
xor U14679 (N_14679,N_6522,N_9433);
and U14680 (N_14680,N_9959,N_5721);
nor U14681 (N_14681,N_8934,N_9144);
and U14682 (N_14682,N_5923,N_6112);
nor U14683 (N_14683,N_7582,N_5344);
nor U14684 (N_14684,N_8679,N_5455);
or U14685 (N_14685,N_7493,N_7708);
and U14686 (N_14686,N_9989,N_9946);
nor U14687 (N_14687,N_6190,N_6979);
nand U14688 (N_14688,N_9433,N_7702);
nand U14689 (N_14689,N_5885,N_9781);
and U14690 (N_14690,N_9512,N_5069);
or U14691 (N_14691,N_8951,N_9724);
nor U14692 (N_14692,N_6508,N_5792);
and U14693 (N_14693,N_6671,N_7369);
and U14694 (N_14694,N_6834,N_9825);
or U14695 (N_14695,N_5387,N_5189);
xnor U14696 (N_14696,N_6387,N_9657);
and U14697 (N_14697,N_7204,N_7854);
xnor U14698 (N_14698,N_5440,N_8075);
nand U14699 (N_14699,N_9817,N_8298);
nor U14700 (N_14700,N_5926,N_5545);
and U14701 (N_14701,N_6277,N_8008);
nor U14702 (N_14702,N_7516,N_5643);
nor U14703 (N_14703,N_9228,N_6407);
xnor U14704 (N_14704,N_5439,N_9275);
xor U14705 (N_14705,N_9322,N_8983);
nor U14706 (N_14706,N_7970,N_6686);
nand U14707 (N_14707,N_6990,N_6671);
nand U14708 (N_14708,N_9814,N_7498);
xor U14709 (N_14709,N_6288,N_5441);
xor U14710 (N_14710,N_7063,N_5639);
nor U14711 (N_14711,N_9293,N_9926);
nand U14712 (N_14712,N_5252,N_6824);
or U14713 (N_14713,N_5443,N_8008);
xor U14714 (N_14714,N_7939,N_9249);
xor U14715 (N_14715,N_7167,N_6519);
and U14716 (N_14716,N_8170,N_9913);
xnor U14717 (N_14717,N_6488,N_6713);
nor U14718 (N_14718,N_9420,N_7173);
xor U14719 (N_14719,N_7437,N_7665);
xnor U14720 (N_14720,N_8272,N_7338);
and U14721 (N_14721,N_9142,N_6532);
nor U14722 (N_14722,N_7508,N_8478);
nand U14723 (N_14723,N_6854,N_8904);
nand U14724 (N_14724,N_7184,N_9394);
nor U14725 (N_14725,N_6398,N_8070);
xor U14726 (N_14726,N_6600,N_9678);
and U14727 (N_14727,N_5648,N_9791);
and U14728 (N_14728,N_7923,N_5248);
and U14729 (N_14729,N_6459,N_9667);
nand U14730 (N_14730,N_8797,N_9691);
nand U14731 (N_14731,N_5417,N_9297);
or U14732 (N_14732,N_8107,N_8038);
nor U14733 (N_14733,N_5453,N_9948);
nor U14734 (N_14734,N_5062,N_8020);
xor U14735 (N_14735,N_8832,N_6298);
xor U14736 (N_14736,N_5963,N_9569);
or U14737 (N_14737,N_5949,N_6551);
nand U14738 (N_14738,N_7196,N_9764);
and U14739 (N_14739,N_8078,N_5819);
or U14740 (N_14740,N_5859,N_9313);
xor U14741 (N_14741,N_5855,N_9524);
xnor U14742 (N_14742,N_6292,N_7787);
nand U14743 (N_14743,N_9118,N_7222);
nand U14744 (N_14744,N_6850,N_8159);
nor U14745 (N_14745,N_7400,N_5507);
and U14746 (N_14746,N_6507,N_8093);
nand U14747 (N_14747,N_5544,N_6712);
nor U14748 (N_14748,N_9893,N_6228);
xor U14749 (N_14749,N_5216,N_8541);
or U14750 (N_14750,N_7884,N_9702);
xnor U14751 (N_14751,N_8528,N_5955);
nor U14752 (N_14752,N_8503,N_6399);
xor U14753 (N_14753,N_5039,N_8767);
and U14754 (N_14754,N_8272,N_5217);
nand U14755 (N_14755,N_8006,N_7250);
nor U14756 (N_14756,N_9385,N_8951);
xor U14757 (N_14757,N_8334,N_7647);
and U14758 (N_14758,N_9549,N_8818);
and U14759 (N_14759,N_9843,N_5891);
nand U14760 (N_14760,N_8518,N_8605);
or U14761 (N_14761,N_9449,N_7470);
xnor U14762 (N_14762,N_7978,N_8803);
xnor U14763 (N_14763,N_7277,N_6760);
nor U14764 (N_14764,N_7178,N_8938);
xor U14765 (N_14765,N_9988,N_6505);
nand U14766 (N_14766,N_8049,N_6484);
nand U14767 (N_14767,N_7774,N_8239);
nor U14768 (N_14768,N_7558,N_8574);
xnor U14769 (N_14769,N_8584,N_6984);
and U14770 (N_14770,N_9482,N_6166);
nand U14771 (N_14771,N_7587,N_8649);
or U14772 (N_14772,N_6567,N_7019);
nand U14773 (N_14773,N_6873,N_6510);
nor U14774 (N_14774,N_7618,N_5969);
and U14775 (N_14775,N_8745,N_6451);
nand U14776 (N_14776,N_7329,N_8131);
and U14777 (N_14777,N_8339,N_8690);
nor U14778 (N_14778,N_7231,N_8849);
nor U14779 (N_14779,N_9119,N_9972);
or U14780 (N_14780,N_8940,N_7104);
xor U14781 (N_14781,N_6910,N_6245);
xnor U14782 (N_14782,N_7912,N_9690);
xnor U14783 (N_14783,N_6681,N_8219);
nor U14784 (N_14784,N_8453,N_9257);
and U14785 (N_14785,N_6809,N_6032);
nand U14786 (N_14786,N_5932,N_6581);
nand U14787 (N_14787,N_9002,N_8568);
nor U14788 (N_14788,N_9881,N_7877);
nand U14789 (N_14789,N_8652,N_5620);
and U14790 (N_14790,N_7494,N_6831);
xor U14791 (N_14791,N_6026,N_8041);
nor U14792 (N_14792,N_7671,N_6235);
or U14793 (N_14793,N_6107,N_7175);
xor U14794 (N_14794,N_5261,N_6031);
nor U14795 (N_14795,N_7826,N_8092);
nand U14796 (N_14796,N_8978,N_9557);
or U14797 (N_14797,N_5017,N_6726);
xnor U14798 (N_14798,N_7194,N_7615);
nand U14799 (N_14799,N_9104,N_5944);
or U14800 (N_14800,N_5760,N_8243);
nor U14801 (N_14801,N_6376,N_5694);
xnor U14802 (N_14802,N_7286,N_9247);
or U14803 (N_14803,N_7954,N_6996);
nand U14804 (N_14804,N_7327,N_7744);
or U14805 (N_14805,N_8209,N_7658);
nand U14806 (N_14806,N_5932,N_9903);
xnor U14807 (N_14807,N_7588,N_6552);
or U14808 (N_14808,N_6908,N_6537);
xor U14809 (N_14809,N_6813,N_7891);
xor U14810 (N_14810,N_9627,N_7991);
nor U14811 (N_14811,N_9721,N_5830);
and U14812 (N_14812,N_7639,N_7894);
or U14813 (N_14813,N_8964,N_6136);
xnor U14814 (N_14814,N_9465,N_9265);
nand U14815 (N_14815,N_9281,N_7558);
nand U14816 (N_14816,N_5160,N_7954);
nor U14817 (N_14817,N_9977,N_7023);
xnor U14818 (N_14818,N_8260,N_6363);
and U14819 (N_14819,N_5769,N_5980);
nand U14820 (N_14820,N_8942,N_5610);
nor U14821 (N_14821,N_5512,N_6302);
or U14822 (N_14822,N_8256,N_9997);
nand U14823 (N_14823,N_6315,N_6737);
xnor U14824 (N_14824,N_8967,N_8499);
nor U14825 (N_14825,N_6227,N_8514);
nor U14826 (N_14826,N_5478,N_7476);
and U14827 (N_14827,N_8211,N_8128);
or U14828 (N_14828,N_7931,N_9853);
xnor U14829 (N_14829,N_6740,N_8859);
or U14830 (N_14830,N_8776,N_9021);
and U14831 (N_14831,N_8034,N_6758);
or U14832 (N_14832,N_8341,N_9117);
nor U14833 (N_14833,N_6206,N_9178);
xnor U14834 (N_14834,N_7002,N_6502);
or U14835 (N_14835,N_9445,N_8925);
nand U14836 (N_14836,N_6630,N_5116);
or U14837 (N_14837,N_5714,N_8959);
or U14838 (N_14838,N_5547,N_5965);
nand U14839 (N_14839,N_6277,N_6956);
nor U14840 (N_14840,N_5013,N_7701);
xnor U14841 (N_14841,N_7456,N_5318);
nor U14842 (N_14842,N_8364,N_8099);
or U14843 (N_14843,N_6755,N_8530);
and U14844 (N_14844,N_7842,N_9667);
nor U14845 (N_14845,N_5358,N_9817);
or U14846 (N_14846,N_8951,N_8056);
nand U14847 (N_14847,N_7453,N_9317);
and U14848 (N_14848,N_6509,N_5208);
nand U14849 (N_14849,N_5196,N_5875);
xnor U14850 (N_14850,N_5397,N_6425);
or U14851 (N_14851,N_5747,N_8299);
or U14852 (N_14852,N_6070,N_7373);
xnor U14853 (N_14853,N_7979,N_8975);
or U14854 (N_14854,N_5808,N_5902);
xnor U14855 (N_14855,N_7517,N_9717);
nor U14856 (N_14856,N_6739,N_9849);
nand U14857 (N_14857,N_8463,N_5165);
and U14858 (N_14858,N_7838,N_5762);
nand U14859 (N_14859,N_6638,N_6479);
nor U14860 (N_14860,N_6375,N_7359);
and U14861 (N_14861,N_9017,N_5978);
xor U14862 (N_14862,N_6044,N_8243);
nand U14863 (N_14863,N_9691,N_6234);
xnor U14864 (N_14864,N_6089,N_7293);
xor U14865 (N_14865,N_6367,N_7012);
or U14866 (N_14866,N_9204,N_6796);
nor U14867 (N_14867,N_5625,N_7069);
and U14868 (N_14868,N_9287,N_8122);
nand U14869 (N_14869,N_7486,N_5668);
nor U14870 (N_14870,N_8652,N_6639);
xor U14871 (N_14871,N_7795,N_6071);
nand U14872 (N_14872,N_6036,N_7531);
or U14873 (N_14873,N_8287,N_7454);
nand U14874 (N_14874,N_8970,N_8354);
or U14875 (N_14875,N_7920,N_5407);
or U14876 (N_14876,N_7241,N_5032);
xor U14877 (N_14877,N_9922,N_5694);
and U14878 (N_14878,N_7122,N_5772);
nor U14879 (N_14879,N_8446,N_8980);
and U14880 (N_14880,N_8460,N_9922);
and U14881 (N_14881,N_9189,N_5314);
and U14882 (N_14882,N_7337,N_6436);
xor U14883 (N_14883,N_6870,N_6191);
nand U14884 (N_14884,N_9940,N_8050);
and U14885 (N_14885,N_8334,N_8307);
nor U14886 (N_14886,N_9953,N_9866);
and U14887 (N_14887,N_8358,N_6385);
and U14888 (N_14888,N_6805,N_5688);
nand U14889 (N_14889,N_6653,N_8278);
nor U14890 (N_14890,N_5983,N_7324);
and U14891 (N_14891,N_5291,N_9999);
xnor U14892 (N_14892,N_8244,N_6097);
xnor U14893 (N_14893,N_8157,N_5510);
and U14894 (N_14894,N_5329,N_6283);
nor U14895 (N_14895,N_9077,N_7323);
or U14896 (N_14896,N_6148,N_6263);
nor U14897 (N_14897,N_5282,N_9631);
nand U14898 (N_14898,N_5937,N_7527);
and U14899 (N_14899,N_5227,N_5650);
nand U14900 (N_14900,N_8636,N_6064);
or U14901 (N_14901,N_6555,N_7942);
xnor U14902 (N_14902,N_5876,N_7343);
or U14903 (N_14903,N_5711,N_6024);
nor U14904 (N_14904,N_6839,N_6694);
nand U14905 (N_14905,N_8790,N_9816);
or U14906 (N_14906,N_7301,N_7926);
xor U14907 (N_14907,N_9000,N_8422);
nor U14908 (N_14908,N_9541,N_9084);
or U14909 (N_14909,N_8466,N_5359);
nand U14910 (N_14910,N_5054,N_9608);
nand U14911 (N_14911,N_9091,N_7414);
xnor U14912 (N_14912,N_7996,N_9507);
and U14913 (N_14913,N_8960,N_8809);
nor U14914 (N_14914,N_9412,N_8575);
and U14915 (N_14915,N_7718,N_8017);
nor U14916 (N_14916,N_5316,N_6305);
xor U14917 (N_14917,N_5260,N_8648);
nor U14918 (N_14918,N_9355,N_7014);
nor U14919 (N_14919,N_8208,N_8986);
or U14920 (N_14920,N_6224,N_9103);
xor U14921 (N_14921,N_6868,N_9109);
nand U14922 (N_14922,N_6088,N_9092);
xor U14923 (N_14923,N_7065,N_9331);
nor U14924 (N_14924,N_7398,N_5989);
and U14925 (N_14925,N_9457,N_7242);
xor U14926 (N_14926,N_9824,N_9053);
or U14927 (N_14927,N_6242,N_7434);
nand U14928 (N_14928,N_9122,N_9925);
and U14929 (N_14929,N_5781,N_8661);
xor U14930 (N_14930,N_8600,N_6071);
nor U14931 (N_14931,N_8456,N_6231);
and U14932 (N_14932,N_8040,N_9955);
or U14933 (N_14933,N_8532,N_5832);
nand U14934 (N_14934,N_8613,N_6140);
xor U14935 (N_14935,N_6619,N_9786);
or U14936 (N_14936,N_9744,N_5279);
or U14937 (N_14937,N_9176,N_9024);
nor U14938 (N_14938,N_6798,N_6647);
nor U14939 (N_14939,N_8653,N_9298);
and U14940 (N_14940,N_8317,N_7203);
or U14941 (N_14941,N_6967,N_6360);
nor U14942 (N_14942,N_8280,N_9306);
and U14943 (N_14943,N_7836,N_5914);
nor U14944 (N_14944,N_8963,N_8283);
or U14945 (N_14945,N_5228,N_6083);
or U14946 (N_14946,N_5406,N_7663);
and U14947 (N_14947,N_8404,N_6917);
xnor U14948 (N_14948,N_6801,N_5524);
nand U14949 (N_14949,N_8875,N_8276);
or U14950 (N_14950,N_8453,N_5899);
nand U14951 (N_14951,N_5816,N_6803);
or U14952 (N_14952,N_8385,N_8280);
xor U14953 (N_14953,N_8591,N_5426);
xor U14954 (N_14954,N_9976,N_6735);
xnor U14955 (N_14955,N_8904,N_5313);
and U14956 (N_14956,N_6913,N_6920);
nand U14957 (N_14957,N_7989,N_5318);
nand U14958 (N_14958,N_9987,N_5421);
nand U14959 (N_14959,N_6480,N_6269);
xor U14960 (N_14960,N_5144,N_7249);
nand U14961 (N_14961,N_5451,N_8601);
or U14962 (N_14962,N_9586,N_8975);
and U14963 (N_14963,N_6492,N_5529);
nand U14964 (N_14964,N_8721,N_7657);
nand U14965 (N_14965,N_9022,N_9021);
xnor U14966 (N_14966,N_5717,N_5144);
xor U14967 (N_14967,N_7830,N_7908);
nor U14968 (N_14968,N_7400,N_8711);
and U14969 (N_14969,N_6025,N_8701);
xnor U14970 (N_14970,N_6530,N_6016);
nand U14971 (N_14971,N_8463,N_9825);
nor U14972 (N_14972,N_6896,N_7880);
and U14973 (N_14973,N_5971,N_9584);
or U14974 (N_14974,N_7233,N_6190);
nor U14975 (N_14975,N_8363,N_6966);
nand U14976 (N_14976,N_9958,N_8135);
or U14977 (N_14977,N_7581,N_8686);
nand U14978 (N_14978,N_7162,N_9249);
xor U14979 (N_14979,N_9243,N_9434);
nand U14980 (N_14980,N_9454,N_9922);
xor U14981 (N_14981,N_5456,N_5818);
or U14982 (N_14982,N_7423,N_6325);
nor U14983 (N_14983,N_9802,N_6838);
xnor U14984 (N_14984,N_6459,N_7489);
and U14985 (N_14985,N_9575,N_8459);
nand U14986 (N_14986,N_5481,N_5116);
or U14987 (N_14987,N_9639,N_9197);
xor U14988 (N_14988,N_5354,N_8036);
nor U14989 (N_14989,N_9784,N_9717);
xnor U14990 (N_14990,N_9700,N_9774);
and U14991 (N_14991,N_5857,N_8115);
nor U14992 (N_14992,N_9241,N_8278);
nand U14993 (N_14993,N_7971,N_7232);
nand U14994 (N_14994,N_9458,N_8481);
nand U14995 (N_14995,N_9907,N_6139);
and U14996 (N_14996,N_7914,N_7903);
or U14997 (N_14997,N_7830,N_5057);
xnor U14998 (N_14998,N_5578,N_7449);
and U14999 (N_14999,N_5991,N_6624);
xnor U15000 (N_15000,N_10713,N_13815);
xor U15001 (N_15001,N_14785,N_14373);
or U15002 (N_15002,N_13533,N_11670);
xor U15003 (N_15003,N_10574,N_12771);
xor U15004 (N_15004,N_13126,N_12184);
or U15005 (N_15005,N_12324,N_10876);
xnor U15006 (N_15006,N_13922,N_10421);
or U15007 (N_15007,N_14669,N_10431);
or U15008 (N_15008,N_14722,N_14989);
xnor U15009 (N_15009,N_13301,N_11780);
nor U15010 (N_15010,N_14371,N_14942);
and U15011 (N_15011,N_14774,N_12294);
and U15012 (N_15012,N_10850,N_11635);
and U15013 (N_15013,N_10372,N_11575);
and U15014 (N_15014,N_11485,N_10238);
nand U15015 (N_15015,N_10654,N_14219);
nor U15016 (N_15016,N_14132,N_14603);
and U15017 (N_15017,N_10236,N_12461);
xor U15018 (N_15018,N_10323,N_11545);
nand U15019 (N_15019,N_14453,N_14519);
or U15020 (N_15020,N_13620,N_13544);
nor U15021 (N_15021,N_12232,N_11756);
and U15022 (N_15022,N_13887,N_11494);
and U15023 (N_15023,N_12208,N_11304);
and U15024 (N_15024,N_11006,N_12080);
xor U15025 (N_15025,N_14059,N_12648);
and U15026 (N_15026,N_11112,N_12941);
nand U15027 (N_15027,N_13600,N_14849);
or U15028 (N_15028,N_13347,N_11057);
nand U15029 (N_15029,N_11283,N_10561);
or U15030 (N_15030,N_10439,N_10247);
xnor U15031 (N_15031,N_11521,N_13291);
xnor U15032 (N_15032,N_14437,N_12172);
nor U15033 (N_15033,N_14225,N_13538);
and U15034 (N_15034,N_12198,N_11370);
and U15035 (N_15035,N_14996,N_12818);
xnor U15036 (N_15036,N_12051,N_12511);
xnor U15037 (N_15037,N_10605,N_12246);
or U15038 (N_15038,N_10956,N_10181);
xnor U15039 (N_15039,N_12234,N_13860);
nor U15040 (N_15040,N_14995,N_14833);
xor U15041 (N_15041,N_14843,N_11888);
xor U15042 (N_15042,N_13574,N_10933);
nor U15043 (N_15043,N_10278,N_12591);
xnor U15044 (N_15044,N_11622,N_14697);
nand U15045 (N_15045,N_10827,N_14736);
xnor U15046 (N_15046,N_13254,N_14422);
or U15047 (N_15047,N_10808,N_14546);
xnor U15048 (N_15048,N_14513,N_11335);
xnor U15049 (N_15049,N_10169,N_11506);
xor U15050 (N_15050,N_12154,N_14004);
or U15051 (N_15051,N_14465,N_13270);
xor U15052 (N_15052,N_11799,N_10538);
nor U15053 (N_15053,N_11072,N_10925);
and U15054 (N_15054,N_12054,N_14290);
nand U15055 (N_15055,N_14881,N_14742);
xnor U15056 (N_15056,N_11765,N_12245);
xor U15057 (N_15057,N_10168,N_11679);
and U15058 (N_15058,N_10893,N_12380);
nor U15059 (N_15059,N_10855,N_12560);
nor U15060 (N_15060,N_14951,N_11994);
or U15061 (N_15061,N_12181,N_13409);
nand U15062 (N_15062,N_10902,N_12578);
xor U15063 (N_15063,N_11712,N_10687);
and U15064 (N_15064,N_11873,N_14585);
nor U15065 (N_15065,N_10601,N_11911);
nor U15066 (N_15066,N_10977,N_14434);
and U15067 (N_15067,N_14700,N_14845);
nor U15068 (N_15068,N_11464,N_10949);
nand U15069 (N_15069,N_10979,N_11022);
xor U15070 (N_15070,N_10491,N_11499);
xnor U15071 (N_15071,N_12641,N_12185);
xnor U15072 (N_15072,N_12371,N_11204);
or U15073 (N_15073,N_12488,N_13774);
and U15074 (N_15074,N_11559,N_11916);
and U15075 (N_15075,N_11385,N_12233);
nor U15076 (N_15076,N_10381,N_14897);
or U15077 (N_15077,N_12948,N_13666);
xnor U15078 (N_15078,N_12748,N_11656);
xnor U15079 (N_15079,N_10974,N_13144);
and U15080 (N_15080,N_10283,N_14027);
nand U15081 (N_15081,N_14285,N_11353);
or U15082 (N_15082,N_11946,N_14433);
nand U15083 (N_15083,N_11035,N_13532);
and U15084 (N_15084,N_14076,N_14760);
and U15085 (N_15085,N_10208,N_13726);
nor U15086 (N_15086,N_11746,N_14092);
nor U15087 (N_15087,N_14918,N_13374);
xor U15088 (N_15088,N_11801,N_10055);
xor U15089 (N_15089,N_11044,N_11291);
nand U15090 (N_15090,N_12375,N_11583);
nand U15091 (N_15091,N_10680,N_10034);
xor U15092 (N_15092,N_13388,N_14958);
or U15093 (N_15093,N_11252,N_13548);
xnor U15094 (N_15094,N_10670,N_11382);
or U15095 (N_15095,N_12250,N_10694);
nand U15096 (N_15096,N_11984,N_14956);
nor U15097 (N_15097,N_13528,N_14087);
and U15098 (N_15098,N_14895,N_14628);
nand U15099 (N_15099,N_10139,N_14034);
nand U15100 (N_15100,N_14738,N_11964);
nor U15101 (N_15101,N_10269,N_12601);
and U15102 (N_15102,N_10768,N_13603);
nor U15103 (N_15103,N_10820,N_14477);
nor U15104 (N_15104,N_13673,N_14043);
xor U15105 (N_15105,N_10194,N_11699);
or U15106 (N_15106,N_10607,N_12997);
xnor U15107 (N_15107,N_10767,N_14035);
xor U15108 (N_15108,N_14348,N_13503);
xor U15109 (N_15109,N_12792,N_12118);
nor U15110 (N_15110,N_11373,N_13688);
or U15111 (N_15111,N_13809,N_12483);
and U15112 (N_15112,N_14349,N_13236);
nor U15113 (N_15113,N_13235,N_13753);
and U15114 (N_15114,N_13911,N_11560);
nor U15115 (N_15115,N_10683,N_10301);
nand U15116 (N_15116,N_14495,N_12244);
nand U15117 (N_15117,N_14049,N_10839);
nand U15118 (N_15118,N_10866,N_13054);
or U15119 (N_15119,N_11748,N_11923);
and U15120 (N_15120,N_10412,N_10100);
nor U15121 (N_15121,N_14478,N_14795);
or U15122 (N_15122,N_13466,N_13734);
nand U15123 (N_15123,N_11609,N_11488);
nand U15124 (N_15124,N_11033,N_11692);
xnor U15125 (N_15125,N_10882,N_14379);
xnor U15126 (N_15126,N_11973,N_13178);
nand U15127 (N_15127,N_11932,N_14636);
and U15128 (N_15128,N_13875,N_10463);
nand U15129 (N_15129,N_11685,N_13523);
xor U15130 (N_15130,N_14862,N_12078);
nand U15131 (N_15131,N_11008,N_10591);
nand U15132 (N_15132,N_14124,N_14028);
and U15133 (N_15133,N_11358,N_11403);
xnor U15134 (N_15134,N_11000,N_12799);
or U15135 (N_15135,N_12654,N_11844);
or U15136 (N_15136,N_10122,N_11711);
nor U15137 (N_15137,N_13959,N_10216);
nor U15138 (N_15138,N_12343,N_14852);
xnor U15139 (N_15139,N_12366,N_12123);
and U15140 (N_15140,N_11238,N_11982);
xnor U15141 (N_15141,N_12254,N_12721);
and U15142 (N_15142,N_14014,N_12731);
and U15143 (N_15143,N_13190,N_10916);
nor U15144 (N_15144,N_14982,N_14428);
nand U15145 (N_15145,N_10110,N_10059);
nor U15146 (N_15146,N_14611,N_14113);
and U15147 (N_15147,N_10415,N_12551);
nand U15148 (N_15148,N_13246,N_10316);
nand U15149 (N_15149,N_13589,N_12664);
and U15150 (N_15150,N_14330,N_13304);
xor U15151 (N_15151,N_10281,N_11914);
nor U15152 (N_15152,N_12336,N_12262);
or U15153 (N_15153,N_11438,N_13970);
xor U15154 (N_15154,N_10815,N_10420);
xor U15155 (N_15155,N_13325,N_14719);
nor U15156 (N_15156,N_12061,N_12588);
nand U15157 (N_15157,N_10470,N_11338);
nand U15158 (N_15158,N_10403,N_14621);
nor U15159 (N_15159,N_11881,N_14073);
xor U15160 (N_15160,N_14333,N_10520);
nand U15161 (N_15161,N_13316,N_10273);
nand U15162 (N_15162,N_10571,N_12943);
nand U15163 (N_15163,N_13307,N_13816);
or U15164 (N_15164,N_14528,N_10478);
xor U15165 (N_15165,N_13442,N_10954);
and U15166 (N_15166,N_12173,N_14165);
or U15167 (N_15167,N_11846,N_14788);
xnor U15168 (N_15168,N_13718,N_10417);
xnor U15169 (N_15169,N_12758,N_11715);
nor U15170 (N_15170,N_10096,N_10159);
xnor U15171 (N_15171,N_12691,N_13955);
or U15172 (N_15172,N_11056,N_12710);
nand U15173 (N_15173,N_10896,N_10294);
nand U15174 (N_15174,N_13559,N_13396);
nand U15175 (N_15175,N_12940,N_10353);
nor U15176 (N_15176,N_10393,N_13974);
and U15177 (N_15177,N_10277,N_13111);
nor U15178 (N_15178,N_13663,N_13473);
or U15179 (N_15179,N_14518,N_12044);
nor U15180 (N_15180,N_13892,N_14872);
or U15181 (N_15181,N_13188,N_12686);
and U15182 (N_15182,N_12919,N_12155);
xor U15183 (N_15183,N_14311,N_11917);
and U15184 (N_15184,N_11629,N_13822);
nor U15185 (N_15185,N_13381,N_10518);
nor U15186 (N_15186,N_12117,N_13091);
and U15187 (N_15187,N_14575,N_13963);
xnor U15188 (N_15188,N_10540,N_13013);
nor U15189 (N_15189,N_13711,N_11132);
nor U15190 (N_15190,N_14684,N_10928);
nand U15191 (N_15191,N_11228,N_11834);
or U15192 (N_15192,N_14990,N_13321);
nand U15193 (N_15193,N_14119,N_13329);
or U15194 (N_15194,N_13365,N_10483);
nor U15195 (N_15195,N_13370,N_10813);
nand U15196 (N_15196,N_14935,N_10743);
and U15197 (N_15197,N_11084,N_10148);
or U15198 (N_15198,N_11927,N_12162);
or U15199 (N_15199,N_10380,N_13668);
nor U15200 (N_15200,N_13098,N_10618);
nor U15201 (N_15201,N_13707,N_12190);
nor U15202 (N_15202,N_12222,N_14058);
and U15203 (N_15203,N_13938,N_12410);
xnor U15204 (N_15204,N_12287,N_14095);
xor U15205 (N_15205,N_14279,N_12150);
and U15206 (N_15206,N_14765,N_10600);
nor U15207 (N_15207,N_14509,N_13817);
nor U15208 (N_15208,N_11139,N_12901);
nor U15209 (N_15209,N_13170,N_13171);
nand U15210 (N_15210,N_13040,N_10230);
or U15211 (N_15211,N_11096,N_11552);
nor U15212 (N_15212,N_10073,N_13501);
nand U15213 (N_15213,N_10578,N_13750);
or U15214 (N_15214,N_14046,N_13036);
or U15215 (N_15215,N_13217,N_14790);
or U15216 (N_15216,N_10461,N_14824);
nor U15217 (N_15217,N_12963,N_11413);
nor U15218 (N_15218,N_12216,N_13653);
or U15219 (N_15219,N_11406,N_12482);
and U15220 (N_15220,N_13848,N_14713);
xor U15221 (N_15221,N_13529,N_10061);
and U15222 (N_15222,N_13279,N_13695);
xnor U15223 (N_15223,N_14754,N_14159);
nand U15224 (N_15224,N_13818,N_11101);
and U15225 (N_15225,N_10496,N_10919);
xor U15226 (N_15226,N_13511,N_10634);
xnor U15227 (N_15227,N_14925,N_12021);
xnor U15228 (N_15228,N_13919,N_12019);
nand U15229 (N_15229,N_12097,N_14751);
and U15230 (N_15230,N_10394,N_12533);
nand U15231 (N_15231,N_11002,N_14067);
and U15232 (N_15232,N_14018,N_14410);
and U15233 (N_15233,N_13696,N_14604);
xnor U15234 (N_15234,N_12487,N_11613);
nor U15235 (N_15235,N_11165,N_10682);
xnor U15236 (N_15236,N_13803,N_14031);
nor U15237 (N_15237,N_14226,N_10632);
nand U15238 (N_15238,N_11273,N_12740);
xor U15239 (N_15239,N_14761,N_10130);
or U15240 (N_15240,N_13748,N_12831);
nand U15241 (N_15241,N_10414,N_10488);
nand U15242 (N_15242,N_14566,N_11543);
or U15243 (N_15243,N_10458,N_11160);
nor U15244 (N_15244,N_10543,N_11179);
nand U15245 (N_15245,N_12773,N_14454);
and U15246 (N_15246,N_10526,N_12703);
and U15247 (N_15247,N_10486,N_13865);
nand U15248 (N_15248,N_10377,N_14971);
nand U15249 (N_15249,N_10806,N_13593);
xnor U15250 (N_15250,N_13904,N_10057);
nor U15251 (N_15251,N_14642,N_11354);
nand U15252 (N_15252,N_10756,N_13915);
and U15253 (N_15253,N_10923,N_11151);
and U15254 (N_15254,N_12841,N_12678);
nand U15255 (N_15255,N_10881,N_13450);
nand U15256 (N_15256,N_12443,N_14666);
or U15257 (N_15257,N_11071,N_12679);
nor U15258 (N_15258,N_10026,N_10580);
nand U15259 (N_15259,N_14402,N_11300);
nand U15260 (N_15260,N_11038,N_11890);
nor U15261 (N_15261,N_11810,N_10691);
or U15262 (N_15262,N_11965,N_13678);
nand U15263 (N_15263,N_10755,N_11872);
xor U15264 (N_15264,N_12301,N_14419);
or U15265 (N_15265,N_10615,N_11297);
and U15266 (N_15266,N_11152,N_14040);
xnor U15267 (N_15267,N_14405,N_14056);
or U15268 (N_15268,N_13512,N_12376);
xor U15269 (N_15269,N_14111,N_10209);
nand U15270 (N_15270,N_14679,N_10892);
xor U15271 (N_15271,N_14266,N_12379);
and U15272 (N_15272,N_11563,N_13759);
or U15273 (N_15273,N_14134,N_10089);
xnor U15274 (N_15274,N_13801,N_14414);
xor U15275 (N_15275,N_12252,N_13319);
nor U15276 (N_15276,N_12354,N_12474);
nor U15277 (N_15277,N_14471,N_13861);
nor U15278 (N_15278,N_11538,N_12439);
or U15279 (N_15279,N_10142,N_11732);
nor U15280 (N_15280,N_12409,N_12018);
xnor U15281 (N_15281,N_13941,N_11417);
xnor U15282 (N_15282,N_10706,N_14607);
and U15283 (N_15283,N_10473,N_12204);
nand U15284 (N_15284,N_12001,N_11404);
nand U15285 (N_15285,N_12899,N_12689);
nor U15286 (N_15286,N_14401,N_14701);
xor U15287 (N_15287,N_14120,N_11637);
and U15288 (N_15288,N_10986,N_12647);
or U15289 (N_15289,N_12312,N_13084);
nand U15290 (N_15290,N_13104,N_10685);
nand U15291 (N_15291,N_12256,N_10443);
nor U15292 (N_15292,N_12039,N_11533);
nor U15293 (N_15293,N_10118,N_11752);
and U15294 (N_15294,N_14517,N_14818);
xnor U15295 (N_15295,N_11540,N_13835);
xnor U15296 (N_15296,N_10966,N_12913);
xnor U15297 (N_15297,N_11663,N_10964);
nor U15298 (N_15298,N_10645,N_11856);
nor U15299 (N_15299,N_13619,N_12258);
nand U15300 (N_15300,N_12548,N_12055);
nor U15301 (N_15301,N_14933,N_14118);
or U15302 (N_15302,N_11673,N_12413);
xnor U15303 (N_15303,N_14823,N_14562);
xnor U15304 (N_15304,N_14888,N_11241);
nor U15305 (N_15305,N_10853,N_11524);
xnor U15306 (N_15306,N_14292,N_12263);
nand U15307 (N_15307,N_14389,N_12856);
nand U15308 (N_15308,N_11742,N_14875);
or U15309 (N_15309,N_12833,N_14681);
nor U15310 (N_15310,N_11725,N_11761);
or U15311 (N_15311,N_12920,N_11860);
nand U15312 (N_15312,N_11630,N_12574);
nor U15313 (N_15313,N_11651,N_12036);
nor U15314 (N_15314,N_14456,N_13960);
and U15315 (N_15315,N_13315,N_10708);
xnor U15316 (N_15316,N_14949,N_12728);
nor U15317 (N_15317,N_14984,N_11850);
and U15318 (N_15318,N_12669,N_11749);
or U15319 (N_15319,N_11526,N_10516);
nor U15320 (N_15320,N_11040,N_12772);
xnor U15321 (N_15321,N_13741,N_10287);
and U15322 (N_15322,N_10418,N_10707);
nand U15323 (N_15323,N_10132,N_10886);
or U15324 (N_15324,N_10400,N_14705);
xnor U15325 (N_15325,N_12670,N_10738);
nand U15326 (N_15326,N_10782,N_10195);
or U15327 (N_15327,N_10482,N_14190);
nor U15328 (N_15328,N_11050,N_13041);
or U15329 (N_15329,N_12300,N_14116);
and U15330 (N_15330,N_14408,N_10941);
and U15331 (N_15331,N_11664,N_10157);
xor U15332 (N_15332,N_14153,N_13356);
nor U15333 (N_15333,N_14934,N_13928);
or U15334 (N_15334,N_10199,N_10432);
or U15335 (N_15335,N_13527,N_10981);
nand U15336 (N_15336,N_11350,N_13326);
nor U15337 (N_15337,N_14457,N_13049);
and U15338 (N_15338,N_14084,N_10428);
nor U15339 (N_15339,N_11420,N_11633);
xor U15340 (N_15340,N_14157,N_10052);
or U15341 (N_15341,N_11076,N_11119);
nor U15342 (N_15342,N_11792,N_12674);
nor U15343 (N_15343,N_12690,N_10335);
nor U15344 (N_15344,N_14128,N_13193);
nand U15345 (N_15345,N_11808,N_10533);
and U15346 (N_15346,N_11694,N_10416);
nor U15347 (N_15347,N_13514,N_12730);
nand U15348 (N_15348,N_11220,N_11416);
xnor U15349 (N_15349,N_14294,N_12497);
nand U15350 (N_15350,N_10668,N_13612);
nand U15351 (N_15351,N_12210,N_11396);
xnor U15352 (N_15352,N_10006,N_11796);
nand U15353 (N_15353,N_13335,N_12192);
nor U15354 (N_15354,N_14491,N_13830);
xnor U15355 (N_15355,N_11012,N_11318);
or U15356 (N_15356,N_13027,N_12267);
xnor U15357 (N_15357,N_13089,N_10865);
or U15358 (N_15358,N_10565,N_14846);
and U15359 (N_15359,N_12053,N_14920);
nor U15360 (N_15360,N_10185,N_14099);
and U15361 (N_15361,N_14343,N_10555);
and U15362 (N_15362,N_11938,N_10289);
xnor U15363 (N_15363,N_11547,N_10655);
nor U15364 (N_15364,N_10003,N_13447);
nand U15365 (N_15365,N_14924,N_11230);
nand U15366 (N_15366,N_14556,N_11546);
or U15367 (N_15367,N_11014,N_13539);
xnor U15368 (N_15368,N_14325,N_10930);
or U15369 (N_15369,N_13605,N_14310);
xnor U15370 (N_15370,N_14199,N_12992);
xor U15371 (N_15371,N_13004,N_10807);
and U15372 (N_15372,N_13278,N_11996);
and U15373 (N_15373,N_13758,N_13588);
xnor U15374 (N_15374,N_10440,N_11989);
nand U15375 (N_15375,N_12939,N_13761);
nand U15376 (N_15376,N_12741,N_12709);
xnor U15377 (N_15377,N_13011,N_12017);
xnor U15378 (N_15378,N_11047,N_14071);
nand U15379 (N_15379,N_10550,N_12951);
and U15380 (N_15380,N_14616,N_14623);
and U15381 (N_15381,N_11723,N_13127);
nand U15382 (N_15382,N_12701,N_11489);
xnor U15383 (N_15383,N_14201,N_13106);
xor U15384 (N_15384,N_12535,N_14555);
nand U15385 (N_15385,N_10429,N_10279);
nor U15386 (N_15386,N_12594,N_14619);
nand U15387 (N_15387,N_10369,N_11019);
nor U15388 (N_15388,N_11753,N_14388);
or U15389 (N_15389,N_11958,N_13449);
nand U15390 (N_15390,N_11631,N_10542);
nor U15391 (N_15391,N_10237,N_10485);
nand U15392 (N_15392,N_13419,N_12149);
and U15393 (N_15393,N_13059,N_14740);
nand U15394 (N_15394,N_14867,N_12255);
nand U15395 (N_15395,N_12978,N_12512);
or U15396 (N_15396,N_11829,N_10628);
nand U15397 (N_15397,N_13039,N_14228);
or U15398 (N_15398,N_10261,N_14955);
nor U15399 (N_15399,N_11561,N_14024);
or U15400 (N_15400,N_14857,N_10757);
and U15401 (N_15401,N_12692,N_10180);
and U15402 (N_15402,N_10164,N_12115);
and U15403 (N_15403,N_13251,N_10354);
or U15404 (N_15404,N_11730,N_14677);
or U15405 (N_15405,N_10252,N_10218);
nand U15406 (N_15406,N_12420,N_11594);
or U15407 (N_15407,N_13080,N_12937);
nand U15408 (N_15408,N_12981,N_11457);
nor U15409 (N_15409,N_12361,N_12297);
nand U15410 (N_15410,N_14552,N_10450);
or U15411 (N_15411,N_11149,N_13375);
nor U15412 (N_15412,N_13926,N_11477);
nor U15413 (N_15413,N_11628,N_13780);
xor U15414 (N_15414,N_13068,N_14727);
nand U15415 (N_15415,N_11103,N_13191);
nand U15416 (N_15416,N_12194,N_14144);
xnor U15417 (N_15417,N_13853,N_12119);
nor U15418 (N_15418,N_12127,N_10135);
and U15419 (N_15419,N_13614,N_13979);
or U15420 (N_15420,N_12604,N_12851);
xnor U15421 (N_15421,N_11310,N_14561);
nor U15422 (N_15422,N_13789,N_13704);
or U15423 (N_15423,N_12809,N_12368);
xor U15424 (N_15424,N_11871,N_10346);
xor U15425 (N_15425,N_12201,N_13585);
nand U15426 (N_15426,N_11997,N_14794);
nand U15427 (N_15427,N_14468,N_11210);
xor U15428 (N_15428,N_13231,N_14635);
nor U15429 (N_15429,N_10868,N_13159);
nand U15430 (N_15430,N_14185,N_10326);
nor U15431 (N_15431,N_10737,N_11407);
or U15432 (N_15432,N_14103,N_13754);
and U15433 (N_15433,N_12737,N_12337);
xnor U15434 (N_15434,N_14251,N_12342);
or U15435 (N_15435,N_14976,N_12849);
xor U15436 (N_15436,N_12935,N_11317);
nand U15437 (N_15437,N_10812,N_10894);
nand U15438 (N_15438,N_12933,N_11323);
or U15439 (N_15439,N_14278,N_10976);
and U15440 (N_15440,N_13681,N_13147);
nor U15441 (N_15441,N_11313,N_10641);
and U15442 (N_15442,N_14182,N_13889);
xor U15443 (N_15443,N_11777,N_12016);
nand U15444 (N_15444,N_13516,N_13716);
xor U15445 (N_15445,N_14932,N_14902);
nand U15446 (N_15446,N_13458,N_11471);
nand U15447 (N_15447,N_12553,N_10290);
nand U15448 (N_15448,N_13829,N_10616);
or U15449 (N_15449,N_11024,N_13694);
nor U15450 (N_15450,N_13196,N_13459);
and U15451 (N_15451,N_13289,N_10253);
or U15452 (N_15452,N_11470,N_10501);
and U15453 (N_15453,N_14931,N_14704);
and U15454 (N_15454,N_11527,N_13766);
nor U15455 (N_15455,N_10733,N_10465);
or U15456 (N_15456,N_10085,N_10444);
nand U15457 (N_15457,N_14717,N_13500);
nor U15458 (N_15458,N_11919,N_10386);
and U15459 (N_15459,N_10529,N_13160);
or U15460 (N_15460,N_10872,N_13699);
and U15461 (N_15461,N_11088,N_13738);
and U15462 (N_15462,N_13406,N_14654);
nor U15463 (N_15463,N_13903,N_14022);
nor U15464 (N_15464,N_11361,N_12713);
nor U15465 (N_15465,N_12542,N_13317);
and U15466 (N_15466,N_14238,N_10936);
nand U15467 (N_15467,N_12481,N_14590);
nor U15468 (N_15468,N_14193,N_12429);
nor U15469 (N_15469,N_11556,N_10714);
and U15470 (N_15470,N_13859,N_11140);
nor U15471 (N_15471,N_13932,N_12893);
and U15472 (N_15472,N_12695,N_14156);
nor U15473 (N_15473,N_13491,N_11430);
and U15474 (N_15474,N_11897,N_14001);
nand U15475 (N_15475,N_10811,N_13705);
xor U15476 (N_15476,N_10536,N_12335);
nand U15477 (N_15477,N_12663,N_13925);
or U15478 (N_15478,N_13854,N_13725);
nor U15479 (N_15479,N_10051,N_12789);
nor U15480 (N_15480,N_12635,N_11514);
or U15481 (N_15481,N_10398,N_12526);
and U15482 (N_15482,N_10291,N_14596);
nand U15483 (N_15483,N_13475,N_11697);
or U15484 (N_15484,N_13224,N_10134);
or U15485 (N_15485,N_10462,N_13845);
nor U15486 (N_15486,N_14516,N_11943);
nor U15487 (N_15487,N_14406,N_10763);
xnor U15488 (N_15488,N_14338,N_14687);
or U15489 (N_15489,N_11678,N_11005);
or U15490 (N_15490,N_14724,N_13713);
nor U15491 (N_15491,N_13402,N_12897);
nor U15492 (N_15492,N_10679,N_11447);
xnor U15493 (N_15493,N_10293,N_14339);
or U15494 (N_15494,N_14905,N_12105);
or U15495 (N_15495,N_10623,N_14577);
nor U15496 (N_15496,N_10970,N_10385);
nand U15497 (N_15497,N_13985,N_12259);
and U15498 (N_15498,N_14879,N_10748);
or U15499 (N_15499,N_14960,N_12870);
or U15500 (N_15500,N_11223,N_11311);
xnor U15501 (N_15501,N_11926,N_13023);
or U15502 (N_15502,N_11900,N_13804);
nand U15503 (N_15503,N_13868,N_11383);
and U15504 (N_15504,N_14661,N_13720);
and U15505 (N_15505,N_11840,N_12166);
xnor U15506 (N_15506,N_13430,N_12791);
or U15507 (N_15507,N_11733,N_11516);
nor U15508 (N_15508,N_10370,N_13542);
xor U15509 (N_15509,N_12008,N_14126);
nand U15510 (N_15510,N_11827,N_13714);
or U15511 (N_15511,N_11154,N_14466);
xor U15512 (N_15512,N_14626,N_10614);
nor U15513 (N_15513,N_14476,N_14364);
or U15514 (N_15514,N_14685,N_11879);
nand U15515 (N_15515,N_10728,N_13006);
xnor U15516 (N_15516,N_10065,N_11921);
nor U15517 (N_15517,N_13670,N_14921);
or U15518 (N_15518,N_11295,N_11500);
nor U15519 (N_15519,N_11388,N_10031);
and U15520 (N_15520,N_14360,N_12108);
nand U15521 (N_15521,N_13141,N_11617);
nor U15522 (N_15522,N_11141,N_11137);
nor U15523 (N_15523,N_14211,N_13571);
or U15524 (N_15524,N_10307,N_11128);
xnor U15525 (N_15525,N_10907,N_10720);
nand U15526 (N_15526,N_10532,N_13031);
and U15527 (N_15527,N_12824,N_13177);
nor U15528 (N_15528,N_12459,N_10722);
nor U15529 (N_15529,N_12332,N_11113);
nor U15530 (N_15530,N_13608,N_13881);
nor U15531 (N_15531,N_14316,N_12011);
xor U15532 (N_15532,N_10711,N_11876);
nand U15533 (N_15533,N_13826,N_14273);
or U15534 (N_15534,N_13556,N_12006);
or U15535 (N_15535,N_12177,N_10171);
and U15536 (N_15536,N_14568,N_14438);
xnor U15537 (N_15537,N_12145,N_13820);
xor U15538 (N_15538,N_12666,N_10310);
nand U15539 (N_15539,N_11728,N_12473);
or U15540 (N_15540,N_11026,N_14377);
nand U15541 (N_15541,N_14579,N_11785);
xnor U15542 (N_15542,N_12161,N_13703);
xnor U15543 (N_15543,N_11276,N_12094);
or U15544 (N_15544,N_11493,N_14385);
xor U15545 (N_15545,N_10397,N_11719);
or U15546 (N_15546,N_10226,N_14652);
xor U15547 (N_15547,N_12872,N_10619);
or U15548 (N_15548,N_12584,N_10384);
nand U15549 (N_15549,N_11551,N_10363);
nand U15550 (N_15550,N_14362,N_14336);
and U15551 (N_15551,N_13808,N_11087);
xnor U15552 (N_15552,N_13138,N_14538);
xnor U15553 (N_15553,N_14836,N_12508);
nand U15554 (N_15554,N_14231,N_10043);
nor U15555 (N_15555,N_14985,N_10522);
nand U15556 (N_15556,N_10248,N_12203);
nand U15557 (N_15557,N_14646,N_14368);
or U15558 (N_15558,N_10260,N_13427);
and U15559 (N_15559,N_14253,N_12549);
xor U15560 (N_15560,N_11875,N_11757);
nand U15561 (N_15561,N_14630,N_13524);
and U15562 (N_15562,N_14841,N_12756);
and U15563 (N_15563,N_11476,N_10544);
xnor U15564 (N_15564,N_13775,N_14322);
or U15565 (N_15565,N_14638,N_10200);
or U15566 (N_15566,N_12066,N_10911);
nor U15567 (N_15567,N_14572,N_12100);
xnor U15568 (N_15568,N_14007,N_10696);
and U15569 (N_15569,N_14009,N_12662);
nand U15570 (N_15570,N_11597,N_11261);
or U15571 (N_15571,N_10880,N_10197);
and U15572 (N_15572,N_13546,N_12527);
nand U15573 (N_15573,N_12480,N_10257);
nand U15574 (N_15574,N_10351,N_12502);
and U15575 (N_15575,N_12885,N_14502);
or U15576 (N_15576,N_10092,N_10837);
xor U15577 (N_15577,N_13950,N_10490);
xnor U15578 (N_15578,N_14557,N_13998);
nor U15579 (N_15579,N_10929,N_12676);
and U15580 (N_15580,N_10495,N_13674);
and U15581 (N_15581,N_11845,N_13969);
nor U15582 (N_15582,N_14649,N_13210);
nand U15583 (N_15583,N_11479,N_12048);
or U15584 (N_15584,N_10007,N_12496);
and U15585 (N_15585,N_14531,N_11331);
nor U15586 (N_15586,N_12349,N_11409);
or U15587 (N_15587,N_11842,N_10531);
nor U15588 (N_15588,N_14909,N_13807);
or U15589 (N_15589,N_13743,N_10022);
or U15590 (N_15590,N_11783,N_13272);
and U15591 (N_15591,N_14163,N_12426);
xor U15592 (N_15592,N_12164,N_12843);
or U15593 (N_15593,N_12993,N_12133);
or U15594 (N_15594,N_10285,N_12165);
nand U15595 (N_15595,N_13504,N_14524);
nand U15596 (N_15596,N_13438,N_13461);
or U15597 (N_15597,N_11522,N_14770);
nor U15598 (N_15598,N_11999,N_12842);
xnor U15599 (N_15599,N_13625,N_14098);
and U15600 (N_15600,N_10249,N_12076);
and U15601 (N_15601,N_12921,N_12815);
nand U15602 (N_15602,N_12945,N_14622);
xnor U15603 (N_15603,N_14768,N_12002);
and U15604 (N_15604,N_10201,N_13487);
nand U15605 (N_15605,N_13420,N_12859);
and U15606 (N_15606,N_14030,N_14643);
and U15607 (N_15607,N_10579,N_14615);
and U15608 (N_15608,N_11389,N_14106);
xnor U15609 (N_15609,N_14672,N_11573);
and U15610 (N_15610,N_11445,N_14822);
xnor U15611 (N_15611,N_14329,N_11429);
and U15612 (N_15612,N_12698,N_14678);
xor U15613 (N_15613,N_11991,N_12029);
nor U15614 (N_15614,N_10479,N_13185);
and U15615 (N_15615,N_13592,N_12453);
xor U15616 (N_15616,N_10572,N_14334);
nor U15617 (N_15617,N_11111,N_14464);
nor U15618 (N_15618,N_10505,N_10947);
nand U15619 (N_15619,N_11588,N_11838);
nor U15620 (N_15620,N_13099,N_12583);
or U15621 (N_15621,N_13944,N_10503);
nor U15622 (N_15622,N_11463,N_13194);
or U15623 (N_15623,N_11131,N_12273);
and U15624 (N_15624,N_13186,N_10072);
nor U15625 (N_15625,N_12506,N_14057);
and U15626 (N_15626,N_11062,N_14928);
xor U15627 (N_15627,N_10740,N_11650);
nor U15628 (N_15628,N_11078,N_13570);
and U15629 (N_15629,N_14798,N_11041);
nor U15630 (N_15630,N_12529,N_13093);
nand U15631 (N_15631,N_12458,N_14299);
or U15632 (N_15632,N_12682,N_14634);
xor U15633 (N_15633,N_10869,N_11557);
xor U15634 (N_15634,N_10651,N_14247);
and U15635 (N_15635,N_12520,N_11755);
and U15636 (N_15636,N_11030,N_13631);
xor U15637 (N_15637,N_13214,N_14158);
xnor U15638 (N_15638,N_14617,N_13480);
nor U15639 (N_15639,N_10700,N_10545);
nand U15640 (N_15640,N_12930,N_11334);
and U15641 (N_15641,N_10321,N_10235);
xnor U15642 (N_15642,N_11536,N_13519);
xnor U15643 (N_15643,N_14224,N_14271);
and U15644 (N_15644,N_14187,N_14961);
xor U15645 (N_15645,N_12652,N_13584);
xor U15646 (N_15646,N_13869,N_13494);
and U15647 (N_15647,N_10425,N_10998);
and U15648 (N_15648,N_10116,N_11599);
xor U15649 (N_15649,N_10802,N_10192);
and U15650 (N_15650,N_13824,N_10456);
and U15651 (N_15651,N_10534,N_10039);
nor U15652 (N_15652,N_11959,N_14694);
nand U15653 (N_15653,N_12460,N_13479);
xor U15654 (N_15654,N_11212,N_11720);
nand U15655 (N_15655,N_10856,N_11978);
or U15656 (N_15656,N_10829,N_13692);
nor U15657 (N_15657,N_11272,N_10358);
nor U15658 (N_15658,N_11836,N_10701);
xnor U15659 (N_15659,N_10863,N_12347);
and U15660 (N_15660,N_11641,N_14758);
nor U15661 (N_15661,N_10282,N_13771);
nor U15662 (N_15662,N_11768,N_11544);
nor U15663 (N_15663,N_13935,N_13227);
xor U15664 (N_15664,N_14730,N_13263);
nand U15665 (N_15665,N_11754,N_13206);
and U15666 (N_15666,N_11963,N_13318);
xnor U15667 (N_15667,N_12310,N_14176);
nor U15668 (N_15668,N_13081,N_10438);
nand U15669 (N_15669,N_14523,N_12186);
nor U15670 (N_15670,N_10141,N_12821);
nand U15671 (N_15671,N_10013,N_12786);
nor U15672 (N_15672,N_13189,N_13685);
or U15673 (N_15673,N_14302,N_11899);
and U15674 (N_15674,N_10915,N_10365);
or U15675 (N_15675,N_12656,N_13783);
xor U15676 (N_15676,N_12720,N_12767);
and U15677 (N_15677,N_10087,N_10175);
or U15678 (N_15678,N_10405,N_10681);
nor U15679 (N_15679,N_11655,N_10952);
nand U15680 (N_15680,N_11893,N_14010);
nor U15681 (N_15681,N_12725,N_12178);
nand U15682 (N_15682,N_13072,N_12450);
nand U15683 (N_15683,N_12622,N_10268);
and U15684 (N_15684,N_11983,N_10189);
and U15685 (N_15685,N_11010,N_12614);
and U15686 (N_15686,N_12522,N_11267);
xor U15687 (N_15687,N_13154,N_10786);
and U15688 (N_15688,N_13526,N_11672);
nor U15689 (N_15689,N_10922,N_11814);
and U15690 (N_15690,N_12341,N_13680);
or U15691 (N_15691,N_13287,N_10554);
and U15692 (N_15692,N_11461,N_14693);
nand U15693 (N_15693,N_13443,N_11639);
or U15694 (N_15694,N_14847,N_10005);
nor U15695 (N_15695,N_13078,N_12314);
or U15696 (N_15696,N_11758,N_14501);
or U15697 (N_15697,N_12829,N_14150);
or U15698 (N_15698,N_14479,N_13618);
and U15699 (N_15699,N_13306,N_10844);
xnor U15700 (N_15700,N_12638,N_14023);
nor U15701 (N_15701,N_13910,N_10914);
nand U15702 (N_15702,N_11608,N_13882);
nor U15703 (N_15703,N_12278,N_10338);
or U15704 (N_15704,N_10048,N_13371);
nor U15705 (N_15705,N_14441,N_12093);
nor U15706 (N_15706,N_11634,N_10008);
and U15707 (N_15707,N_12440,N_13878);
xor U15708 (N_15708,N_13996,N_13435);
xnor U15709 (N_15709,N_10727,N_10675);
xnor U15710 (N_15710,N_13565,N_10090);
nor U15711 (N_15711,N_10136,N_13880);
or U15712 (N_15712,N_10012,N_14455);
or U15713 (N_15713,N_12983,N_12547);
xnor U15714 (N_15714,N_13742,N_10360);
and U15715 (N_15715,N_12753,N_12918);
xor U15716 (N_15716,N_10454,N_13242);
nand U15717 (N_15717,N_10347,N_10311);
and U15718 (N_15718,N_12783,N_13876);
or U15719 (N_15719,N_10732,N_11474);
nand U15720 (N_15720,N_10620,N_14830);
xor U15721 (N_15721,N_12706,N_13408);
xor U15722 (N_15722,N_14032,N_12131);
or U15723 (N_15723,N_14383,N_12009);
xor U15724 (N_15724,N_11190,N_10742);
nor U15725 (N_15725,N_13643,N_11427);
or U15726 (N_15726,N_11001,N_11214);
xnor U15727 (N_15727,N_11198,N_13852);
or U15728 (N_15728,N_13439,N_10938);
or U15729 (N_15729,N_12365,N_14355);
and U15730 (N_15730,N_10703,N_13667);
and U15731 (N_15731,N_10686,N_14392);
or U15732 (N_15732,N_12064,N_11219);
and U15733 (N_15733,N_11760,N_10661);
or U15734 (N_15734,N_12033,N_11433);
xnor U15735 (N_15735,N_10801,N_14232);
and U15736 (N_15736,N_12451,N_12632);
or U15737 (N_15737,N_13228,N_14240);
or U15738 (N_15738,N_14668,N_12477);
nand U15739 (N_15739,N_12214,N_13407);
or U15740 (N_15740,N_13811,N_11045);
nand U15741 (N_15741,N_14537,N_12505);
and U15742 (N_15742,N_11554,N_10202);
nor U15743 (N_15743,N_13945,N_14250);
or U15744 (N_15744,N_10514,N_14397);
nor U15745 (N_15745,N_10138,N_11104);
or U15746 (N_15746,N_10847,N_10630);
nand U15747 (N_15747,N_12081,N_13069);
or U15748 (N_15748,N_13038,N_10948);
xor U15749 (N_15749,N_14815,N_13380);
and U15750 (N_15750,N_10355,N_11595);
and U15751 (N_15751,N_10984,N_13295);
nand U15752 (N_15752,N_12412,N_12971);
nor U15753 (N_15753,N_14171,N_10067);
or U15754 (N_15754,N_10076,N_12757);
or U15755 (N_15755,N_14123,N_12911);
and U15756 (N_15756,N_14994,N_13465);
and U15757 (N_15757,N_13472,N_11346);
or U15758 (N_15758,N_11831,N_13042);
or U15759 (N_15759,N_10587,N_13795);
and U15760 (N_15760,N_10599,N_10071);
nand U15761 (N_15761,N_10017,N_13508);
or U15762 (N_15762,N_11735,N_13812);
and U15763 (N_15763,N_14551,N_12677);
nor U15764 (N_15764,N_10702,N_11689);
or U15765 (N_15765,N_11150,N_13587);
xor U15766 (N_15766,N_12590,N_13292);
or U15767 (N_15767,N_11004,N_11867);
nand U15768 (N_15768,N_12456,N_14204);
nor U15769 (N_15769,N_12914,N_14003);
nand U15770 (N_15770,N_11270,N_13386);
or U15771 (N_15771,N_11703,N_12860);
xnor U15772 (N_15772,N_11886,N_13702);
nor U15773 (N_15773,N_13432,N_12869);
or U15774 (N_15774,N_10564,N_11189);
and U15775 (N_15775,N_10824,N_14564);
nand U15776 (N_15776,N_13989,N_10019);
nand U15777 (N_15777,N_11110,N_13684);
nand U15778 (N_15778,N_11738,N_14194);
xnor U15779 (N_15779,N_10140,N_11822);
nand U15780 (N_15780,N_10303,N_12858);
xor U15781 (N_15781,N_13558,N_12261);
nand U15782 (N_15782,N_13906,N_11042);
or U15783 (N_15783,N_14096,N_14445);
nand U15784 (N_15784,N_12098,N_13256);
xnor U15785 (N_15785,N_11442,N_13708);
and U15786 (N_15786,N_12953,N_13364);
xor U15787 (N_15787,N_10000,N_12472);
nand U15788 (N_15788,N_14313,N_14718);
nand U15789 (N_15789,N_12043,N_11509);
xor U15790 (N_15790,N_13103,N_12257);
xnor U15791 (N_15791,N_12279,N_14482);
xnor U15792 (N_15792,N_10395,N_11803);
and U15793 (N_15793,N_12065,N_11467);
nand U15794 (N_15794,N_14733,N_11710);
nor U15795 (N_15795,N_10436,N_10642);
nand U15796 (N_15796,N_13965,N_11194);
and U15797 (N_15797,N_10375,N_12694);
nor U15798 (N_15798,N_12820,N_11883);
nor U15799 (N_15799,N_14753,N_10776);
nand U15800 (N_15800,N_11604,N_14016);
xnor U15801 (N_15801,N_11788,N_11316);
and U15802 (N_15802,N_14151,N_10819);
xnor U15803 (N_15803,N_13448,N_10459);
nor U15804 (N_15804,N_14281,N_12374);
nand U15805 (N_15805,N_11349,N_13021);
nand U15806 (N_15806,N_14143,N_11640);
or U15807 (N_15807,N_10809,N_13161);
or U15808 (N_15808,N_11903,N_12193);
nor U15809 (N_15809,N_13143,N_13284);
xnor U15810 (N_15810,N_13247,N_12738);
nor U15811 (N_15811,N_10741,N_12800);
nand U15812 (N_15812,N_10577,N_11158);
nand U15813 (N_15813,N_12571,N_13719);
xnor U15814 (N_15814,N_14653,N_14398);
nand U15815 (N_15815,N_14988,N_13333);
or U15816 (N_15816,N_13946,N_12968);
or U15817 (N_15817,N_11052,N_14496);
and U15818 (N_15818,N_13416,N_11607);
xor U15819 (N_15819,N_14964,N_14312);
or U15820 (N_15820,N_13166,N_14763);
or U15821 (N_15821,N_14062,N_14597);
and U15822 (N_15822,N_11369,N_11987);
nand U15823 (N_15823,N_13896,N_14610);
or U15824 (N_15824,N_10978,N_12582);
and U15825 (N_15825,N_11015,N_14169);
or U15826 (N_15826,N_14651,N_10441);
nand U15827 (N_15827,N_11954,N_13382);
or U15828 (N_15828,N_14354,N_14337);
xnor U15829 (N_15829,N_10993,N_14246);
xor U15830 (N_15830,N_11507,N_14806);
or U15831 (N_15831,N_11936,N_10753);
or U15832 (N_15832,N_12345,N_11186);
or U15833 (N_15833,N_11611,N_12229);
xnor U15834 (N_15834,N_12646,N_14946);
nand U15835 (N_15835,N_12402,N_12422);
nor U15836 (N_15836,N_12625,N_12956);
nor U15837 (N_15837,N_12847,N_11623);
xor U15838 (N_15838,N_12736,N_14069);
nand U15839 (N_15839,N_12629,N_11234);
xnor U15840 (N_15840,N_13151,N_11671);
xor U15841 (N_15841,N_10791,N_14569);
nor U15842 (N_15842,N_11049,N_12363);
xor U15843 (N_15843,N_14584,N_13894);
nand U15844 (N_15844,N_13654,N_13182);
xor U15845 (N_15845,N_12433,N_12712);
or U15846 (N_15846,N_12928,N_14142);
nand U15847 (N_15847,N_12762,N_11161);
nand U15848 (N_15848,N_13180,N_13444);
or U15849 (N_15849,N_10666,N_12236);
nand U15850 (N_15850,N_10752,N_14282);
and U15851 (N_15851,N_13568,N_14764);
xor U15852 (N_15852,N_11390,N_10699);
nand U15853 (N_15853,N_10212,N_14966);
or U15854 (N_15854,N_13920,N_14089);
or U15855 (N_15855,N_12340,N_11122);
nor U15856 (N_15856,N_10609,N_14655);
or U15857 (N_15857,N_13455,N_13262);
nand U15858 (N_15858,N_12239,N_13744);
xnor U15859 (N_15859,N_12969,N_10280);
xnor U15860 (N_15860,N_14825,N_13604);
or U15861 (N_15861,N_12724,N_14940);
or U15862 (N_15862,N_11776,N_14184);
and U15863 (N_15863,N_10830,N_12147);
nand U15864 (N_15864,N_14745,N_10477);
or U15865 (N_15865,N_13413,N_12769);
and U15866 (N_15866,N_10025,N_13513);
nand U15867 (N_15867,N_14870,N_14854);
nand U15868 (N_15868,N_12946,N_12538);
nand U15869 (N_15869,N_14341,N_14769);
nand U15870 (N_15870,N_11518,N_13735);
and U15871 (N_15871,N_12389,N_10083);
or U15872 (N_15872,N_14987,N_10590);
xnor U15873 (N_15873,N_13125,N_10760);
nor U15874 (N_15874,N_11074,N_13639);
or U15875 (N_15875,N_11115,N_14460);
nand U15876 (N_15876,N_11393,N_14221);
nand U15877 (N_15877,N_13650,N_11011);
xor U15878 (N_15878,N_13924,N_12248);
nand U15879 (N_15879,N_12806,N_13153);
nor U15880 (N_15880,N_14624,N_12812);
nor U15881 (N_15881,N_10749,N_12082);
nand U15882 (N_15882,N_11969,N_11193);
nor U15883 (N_15883,N_10232,N_12593);
and U15884 (N_15884,N_11525,N_13602);
nand U15885 (N_15885,N_14699,N_12823);
nand U15886 (N_15886,N_13297,N_12853);
nor U15887 (N_15887,N_14793,N_14691);
and U15888 (N_15888,N_13441,N_12546);
or U15889 (N_15889,N_13058,N_10445);
nand U15890 (N_15890,N_10213,N_10848);
nand U15891 (N_15891,N_13348,N_10049);
nand U15892 (N_15892,N_14647,N_10611);
nor U15893 (N_15893,N_12922,N_13721);
nor U15894 (N_15894,N_10300,N_10982);
nand U15895 (N_15895,N_11647,N_11060);
or U15896 (N_15896,N_11855,N_10927);
xor U15897 (N_15897,N_11929,N_14627);
and U15898 (N_15898,N_10508,N_13712);
or U15899 (N_15899,N_14832,N_12388);
nand U15900 (N_15900,N_13359,N_10790);
or U15901 (N_15901,N_11708,N_10960);
nor U15902 (N_15902,N_14952,N_11682);
xnor U15903 (N_15903,N_12565,N_12156);
nand U15904 (N_15904,N_12822,N_11450);
xnor U15905 (N_15905,N_11144,N_14712);
and U15906 (N_15906,N_12597,N_13372);
and U15907 (N_15907,N_14662,N_13505);
and U15908 (N_15908,N_11286,N_10126);
nor U15909 (N_15909,N_13064,N_11163);
xnor U15910 (N_15910,N_12468,N_13662);
xnor U15911 (N_15911,N_10324,N_14080);
or U15912 (N_15912,N_13165,N_10342);
or U15913 (N_15913,N_14506,N_11878);
xor U15914 (N_15914,N_13756,N_13813);
xnor U15915 (N_15915,N_12318,N_10305);
and U15916 (N_15916,N_14412,N_14461);
nand U15917 (N_15917,N_12839,N_13145);
nor U15918 (N_15918,N_14510,N_13362);
and U15919 (N_15919,N_14970,N_10818);
nand U15920 (N_15920,N_14692,N_10079);
nand U15921 (N_15921,N_11377,N_10913);
or U15922 (N_15922,N_10362,N_13831);
or U15923 (N_15923,N_14307,N_11580);
and U15924 (N_15924,N_13395,N_13112);
nor U15925 (N_15925,N_10210,N_13799);
nor U15926 (N_15926,N_11426,N_12942);
or U15927 (N_15927,N_13334,N_11727);
nor U15928 (N_15928,N_12657,N_10299);
nor U15929 (N_15929,N_14805,N_12031);
and U15930 (N_15930,N_12445,N_10155);
nor U15931 (N_15931,N_12357,N_11907);
and U15932 (N_15932,N_13077,N_11884);
nor U15933 (N_15933,N_13632,N_14515);
nand U15934 (N_15934,N_13997,N_10028);
or U15935 (N_15935,N_12364,N_10357);
and U15936 (N_15936,N_11988,N_12878);
and U15937 (N_15937,N_10078,N_10144);
or U15938 (N_15938,N_11397,N_14511);
nand U15939 (N_15939,N_14554,N_13342);
nand U15940 (N_15940,N_14529,N_14780);
or U15941 (N_15941,N_10524,N_12323);
xor U15942 (N_15942,N_11098,N_14420);
xor U15943 (N_15943,N_10953,N_13978);
or U15944 (N_15944,N_11055,N_13390);
xor U15945 (N_15945,N_11809,N_13097);
xnor U15946 (N_15946,N_13198,N_11698);
xor U15947 (N_15947,N_11986,N_10004);
nor U15948 (N_15948,N_14130,N_14417);
nor U15949 (N_15949,N_11660,N_11534);
xor U15950 (N_15950,N_12755,N_10530);
and U15951 (N_15951,N_10243,N_11466);
and U15952 (N_15952,N_13727,N_12382);
nand U15953 (N_15953,N_13757,N_14039);
xor U15954 (N_15954,N_13793,N_10521);
or U15955 (N_15955,N_12727,N_11700);
nor U15956 (N_15956,N_13636,N_14732);
nand U15957 (N_15957,N_11705,N_11368);
or U15958 (N_15958,N_11408,N_13498);
xor U15959 (N_15959,N_10775,N_10095);
and U15960 (N_15960,N_13590,N_14077);
nand U15961 (N_15961,N_12355,N_14814);
and U15962 (N_15962,N_12296,N_11209);
and U15963 (N_15963,N_12970,N_13293);
or U15964 (N_15964,N_10191,N_13821);
and U15965 (N_15965,N_10263,N_10426);
or U15966 (N_15966,N_12982,N_12621);
nor U15967 (N_15967,N_14592,N_13740);
xnor U15968 (N_15968,N_14787,N_11498);
or U15969 (N_15969,N_13252,N_10640);
nand U15970 (N_15970,N_11502,N_10793);
and U15971 (N_15971,N_10724,N_13661);
nor U15972 (N_15972,N_12627,N_13634);
and U15973 (N_15973,N_10217,N_13858);
and U15974 (N_15974,N_10382,N_10566);
nand U15975 (N_15975,N_13129,N_13509);
and U15976 (N_15976,N_13693,N_14242);
nand U15977 (N_15977,N_14580,N_14327);
and U15978 (N_15978,N_13230,N_14962);
and U15979 (N_15979,N_12881,N_10875);
xnor U15980 (N_15980,N_11066,N_13730);
xnor U15981 (N_15981,N_11279,N_11868);
or U15982 (N_15982,N_10822,N_10990);
or U15983 (N_15983,N_14541,N_10671);
nor U15984 (N_15984,N_11555,N_12749);
nand U15985 (N_15985,N_10449,N_13522);
or U15986 (N_15986,N_13842,N_10206);
xnor U15987 (N_15987,N_12544,N_11744);
nor U15988 (N_15988,N_12868,N_10376);
xnor U15989 (N_15989,N_14489,N_11441);
xnor U15990 (N_15990,N_14807,N_14520);
xnor U15991 (N_15991,N_10489,N_12260);
xor U15992 (N_15992,N_11771,N_11106);
and U15993 (N_15993,N_12085,N_12083);
or U15994 (N_15994,N_11195,N_12438);
xor U15995 (N_15995,N_11870,N_11857);
or U15996 (N_15996,N_11109,N_10871);
nand U15997 (N_15997,N_13016,N_11263);
or U15998 (N_15998,N_12465,N_12803);
or U15999 (N_15999,N_12137,N_14664);
nand U16000 (N_16000,N_11774,N_12566);
or U16001 (N_16001,N_11636,N_12517);
or U16002 (N_16002,N_10633,N_10066);
nor U16003 (N_16003,N_12780,N_14026);
or U16004 (N_16004,N_12532,N_13723);
nand U16005 (N_16005,N_11747,N_13032);
nor U16006 (N_16006,N_10211,N_14012);
xnor U16007 (N_16007,N_12475,N_11789);
nor U16008 (N_16008,N_12863,N_13257);
and U16009 (N_16009,N_14136,N_11439);
and U16010 (N_16010,N_11891,N_12224);
and U16011 (N_16011,N_12867,N_12950);
or U16012 (N_16012,N_10153,N_13253);
nor U16013 (N_16013,N_10475,N_14581);
or U16014 (N_16014,N_14085,N_13785);
and U16015 (N_16015,N_12463,N_11759);
nor U16016 (N_16016,N_11456,N_11736);
xor U16017 (N_16017,N_12132,N_11646);
nand U16018 (N_16018,N_14472,N_11869);
nor U16019 (N_16019,N_11704,N_12618);
nor U16020 (N_16020,N_10419,N_11400);
xor U16021 (N_16021,N_14162,N_12299);
or U16022 (N_16022,N_13581,N_13739);
and U16023 (N_16023,N_13288,N_10961);
xor U16024 (N_16024,N_10864,N_10734);
or U16025 (N_16025,N_12158,N_14663);
nand U16026 (N_16026,N_14166,N_12142);
xnor U16027 (N_16027,N_10241,N_12900);
nor U16028 (N_16028,N_12887,N_11437);
and U16029 (N_16029,N_14944,N_11081);
and U16030 (N_16030,N_13116,N_14800);
nor U16031 (N_16031,N_14869,N_10772);
and U16032 (N_16032,N_10563,N_13490);
xnor U16033 (N_16033,N_10918,N_13484);
or U16034 (N_16034,N_14303,N_14345);
nor U16035 (N_16035,N_11902,N_12391);
nor U16036 (N_16036,N_10797,N_11079);
nor U16037 (N_16037,N_11365,N_12134);
nand U16038 (N_16038,N_10383,N_13354);
or U16039 (N_16039,N_12620,N_10705);
xnor U16040 (N_16040,N_12096,N_10971);
or U16041 (N_16041,N_14620,N_11075);
nand U16042 (N_16042,N_10650,N_11553);
nand U16043 (N_16043,N_11157,N_13271);
or U16044 (N_16044,N_14233,N_14323);
or U16045 (N_16045,N_12667,N_10364);
nor U16046 (N_16046,N_13624,N_12228);
or U16047 (N_16047,N_12005,N_13222);
nand U16048 (N_16048,N_11099,N_11668);
or U16049 (N_16049,N_10643,N_12428);
nor U16050 (N_16050,N_14588,N_13350);
or U16051 (N_16051,N_11935,N_11652);
nor U16052 (N_16052,N_12286,N_10537);
xor U16053 (N_16053,N_10674,N_12855);
nand U16054 (N_16054,N_12892,N_12015);
and U16055 (N_16055,N_11933,N_13572);
and U16056 (N_16056,N_12160,N_10256);
and U16057 (N_16057,N_14821,N_13499);
xor U16058 (N_16058,N_13535,N_11848);
nor U16059 (N_16059,N_11453,N_10015);
nand U16060 (N_16060,N_14884,N_13563);
xnor U16061 (N_16061,N_11094,N_13676);
and U16062 (N_16062,N_11950,N_12714);
nor U16063 (N_16063,N_14483,N_13951);
or U16064 (N_16064,N_11250,N_12910);
nor U16065 (N_16065,N_12325,N_12275);
xor U16066 (N_16066,N_11255,N_13898);
xnor U16067 (N_16067,N_14429,N_10091);
or U16068 (N_16068,N_12671,N_11199);
nand U16069 (N_16069,N_14152,N_12673);
xnor U16070 (N_16070,N_11065,N_11481);
nand U16071 (N_16071,N_13168,N_12027);
nand U16072 (N_16072,N_13412,N_12489);
nor U16073 (N_16073,N_10594,N_13417);
xor U16074 (N_16074,N_12333,N_10246);
or U16075 (N_16075,N_13644,N_11155);
nand U16076 (N_16076,N_11515,N_10904);
nand U16077 (N_16077,N_11866,N_14114);
xor U16078 (N_16078,N_12075,N_13917);
nor U16079 (N_16079,N_14521,N_13392);
and U16080 (N_16080,N_14488,N_11603);
nor U16081 (N_16081,N_14188,N_14074);
nor U16082 (N_16082,N_11352,N_11366);
nor U16083 (N_16083,N_13610,N_11253);
and U16084 (N_16084,N_10128,N_14101);
nor U16085 (N_16085,N_14264,N_10359);
or U16086 (N_16086,N_14808,N_13550);
xnor U16087 (N_16087,N_11779,N_13462);
nand U16088 (N_16088,N_12628,N_13836);
or U16089 (N_16089,N_12170,N_14365);
nor U16090 (N_16090,N_14094,N_10295);
or U16091 (N_16091,N_14775,N_10391);
nor U16092 (N_16092,N_13173,N_11203);
or U16093 (N_16093,N_13311,N_13096);
nor U16094 (N_16094,N_13949,N_10709);
or U16095 (N_16095,N_10547,N_10215);
and U16096 (N_16096,N_10487,N_14214);
nor U16097 (N_16097,N_12509,N_13179);
nand U16098 (N_16098,N_10551,N_13690);
xnor U16099 (N_16099,N_12253,N_12188);
or U16100 (N_16100,N_13689,N_10963);
nand U16101 (N_16101,N_12592,N_12060);
and U16102 (N_16102,N_14418,N_11483);
nor U16103 (N_16103,N_13502,N_14395);
xnor U16104 (N_16104,N_12486,N_10942);
nand U16105 (N_16105,N_14848,N_14558);
nand U16106 (N_16106,N_10149,N_14573);
or U16107 (N_16107,N_12020,N_10658);
xor U16108 (N_16108,N_11874,N_10946);
or U16109 (N_16109,N_14503,N_12864);
xor U16110 (N_16110,N_12545,N_13152);
and U16111 (N_16111,N_12788,N_12405);
xor U16112 (N_16112,N_10131,N_10040);
nand U16113 (N_16113,N_14025,N_13094);
or U16114 (N_16114,N_14759,N_13102);
nand U16115 (N_16115,N_12240,N_11529);
and U16116 (N_16116,N_11530,N_10715);
nand U16117 (N_16117,N_13706,N_10114);
xnor U16118 (N_16118,N_12655,N_14695);
and U16119 (N_16119,N_13747,N_10988);
xor U16120 (N_16120,N_12298,N_10081);
nor U16121 (N_16121,N_13934,N_13140);
nor U16122 (N_16122,N_13343,N_13645);
xor U16123 (N_16123,N_11410,N_10313);
xor U16124 (N_16124,N_11211,N_14801);
xnor U16125 (N_16125,N_12759,N_12124);
and U16126 (N_16126,N_12808,N_12176);
nand U16127 (N_16127,N_10225,N_13167);
or U16128 (N_16128,N_11278,N_12399);
nor U16129 (N_16129,N_12810,N_11182);
and U16130 (N_16130,N_11431,N_10889);
nor U16131 (N_16131,N_14550,N_13648);
nor U16132 (N_16132,N_10188,N_10784);
nor U16133 (N_16133,N_14771,N_11566);
or U16134 (N_16134,N_14522,N_11398);
nand U16135 (N_16135,N_10451,N_10825);
xnor U16136 (N_16136,N_12350,N_12977);
and U16137 (N_16137,N_10446,N_12086);
and U16138 (N_16138,N_11343,N_13672);
xnor U16139 (N_16139,N_14186,N_11188);
nand U16140 (N_16140,N_13971,N_13579);
nand U16141 (N_16141,N_10766,N_13872);
xor U16142 (N_16142,N_13276,N_14631);
or U16143 (N_16143,N_12745,N_13005);
or U16144 (N_16144,N_13897,N_10991);
and U16145 (N_16145,N_12972,N_13445);
and U16146 (N_16146,N_11882,N_14858);
or U16147 (N_16147,N_10387,N_14644);
xnor U16148 (N_16148,N_14842,N_13936);
xnor U16149 (N_16149,N_11582,N_13008);
nand U16150 (N_16150,N_13373,N_11224);
nor U16151 (N_16151,N_14260,N_12903);
nor U16152 (N_16152,N_12739,N_12122);
nor U16153 (N_16153,N_13671,N_13065);
nor U16154 (N_16154,N_13033,N_14320);
nor U16155 (N_16155,N_14399,N_14784);
nand U16156 (N_16156,N_11357,N_12798);
or U16157 (N_16157,N_12328,N_10719);
nand U16158 (N_16158,N_10798,N_10325);
nand U16159 (N_16159,N_10069,N_10348);
nor U16160 (N_16160,N_14050,N_13208);
nand U16161 (N_16161,N_12726,N_11918);
nand U16162 (N_16162,N_14696,N_11472);
and U16163 (N_16163,N_10318,N_14177);
xnor U16164 (N_16164,N_14369,N_13067);
nor U16165 (N_16165,N_11657,N_13956);
or U16166 (N_16166,N_11605,N_14589);
nor U16167 (N_16167,N_13204,N_11282);
xor U16168 (N_16168,N_10094,N_11215);
or U16169 (N_16169,N_10411,N_11232);
and U16170 (N_16170,N_10939,N_10684);
nor U16171 (N_16171,N_11620,N_13383);
and U16172 (N_16172,N_11289,N_10525);
or U16173 (N_16173,N_14708,N_10585);
or U16174 (N_16174,N_13806,N_10660);
xor U16175 (N_16175,N_14749,N_13120);
and U16176 (N_16176,N_12894,N_13195);
xor U16177 (N_16177,N_10920,N_10975);
nand U16178 (N_16178,N_11895,N_14683);
nor U16179 (N_16179,N_11764,N_12976);
xor U16180 (N_16180,N_14108,N_10170);
or U16181 (N_16181,N_11955,N_13916);
and U16182 (N_16182,N_13192,N_14161);
nor U16183 (N_16183,N_14110,N_11669);
and U16184 (N_16184,N_10744,N_11460);
or U16185 (N_16185,N_12959,N_13902);
or U16186 (N_16186,N_13506,N_14887);
and U16187 (N_16187,N_11942,N_11051);
nor U16188 (N_16188,N_14378,N_12091);
nand U16189 (N_16189,N_12014,N_11290);
nor U16190 (N_16190,N_10646,N_13244);
or U16191 (N_16191,N_13150,N_14249);
nand U16192 (N_16192,N_13942,N_14967);
or U16193 (N_16193,N_10044,N_13309);
nand U16194 (N_16194,N_12206,N_11130);
or U16195 (N_16195,N_10361,N_14492);
or U16196 (N_16196,N_13424,N_12052);
xor U16197 (N_16197,N_12381,N_14838);
nand U16198 (N_16198,N_14442,N_14196);
and U16199 (N_16199,N_10553,N_14291);
or U16200 (N_16200,N_13700,N_14725);
xnor U16201 (N_16201,N_14435,N_10492);
and U16202 (N_16202,N_14748,N_13765);
nor U16203 (N_16203,N_12639,N_12890);
or U16204 (N_16204,N_13669,N_11244);
and U16205 (N_16205,N_14998,N_10423);
nand U16206 (N_16206,N_12906,N_10466);
nand U16207 (N_16207,N_10220,N_14601);
nand U16208 (N_16208,N_12171,N_12411);
nand U16209 (N_16209,N_12837,N_12114);
xor U16210 (N_16210,N_13322,N_10464);
and U16211 (N_16211,N_10924,N_12163);
and U16212 (N_16212,N_10024,N_11032);
xor U16213 (N_16213,N_14937,N_10644);
nor U16214 (N_16214,N_10373,N_11183);
or U16215 (N_16215,N_10452,N_12866);
nand U16216 (N_16216,N_12238,N_13088);
or U16217 (N_16217,N_11925,N_12125);
nand U16218 (N_16218,N_14553,N_11858);
nand U16219 (N_16219,N_10950,N_10649);
and U16220 (N_16220,N_13947,N_14230);
and U16221 (N_16221,N_11037,N_10622);
nor U16222 (N_16222,N_13035,N_10697);
nor U16223 (N_16223,N_13397,N_12896);
xor U16224 (N_16224,N_11292,N_12493);
and U16225 (N_16225,N_13176,N_12290);
nand U16226 (N_16226,N_12073,N_11977);
xnor U16227 (N_16227,N_13873,N_11567);
nor U16228 (N_16228,N_11362,N_10371);
and U16229 (N_16229,N_14449,N_13710);
nor U16230 (N_16230,N_12598,N_11440);
nand U16231 (N_16231,N_10573,N_11386);
nor U16232 (N_16232,N_10286,N_12103);
xor U16233 (N_16233,N_10379,N_11976);
nor U16234 (N_16234,N_11680,N_12175);
and U16235 (N_16235,N_12912,N_12209);
xor U16236 (N_16236,N_14512,N_12424);
xnor U16237 (N_16237,N_12313,N_14586);
nand U16238 (N_16238,N_13855,N_14786);
xnor U16239 (N_16239,N_12431,N_13486);
xnor U16240 (N_16240,N_12554,N_13857);
nand U16241 (N_16241,N_14474,N_11542);
nand U16242 (N_16242,N_11702,N_14469);
or U16243 (N_16243,N_14305,N_12467);
and U16244 (N_16244,N_11328,N_14900);
xor U16245 (N_16245,N_14079,N_14532);
xor U16246 (N_16246,N_11394,N_11448);
xnor U16247 (N_16247,N_14332,N_14295);
and U16248 (N_16248,N_12558,N_10845);
and U16249 (N_16249,N_14254,N_11523);
nor U16250 (N_16250,N_11061,N_11778);
xnor U16251 (N_16251,N_14140,N_13787);
nor U16252 (N_16252,N_13389,N_12521);
nand U16253 (N_16253,N_12242,N_12151);
nand U16254 (N_16254,N_14008,N_13261);
nand U16255 (N_16255,N_11913,N_11569);
and U16256 (N_16256,N_13531,N_13079);
xnor U16257 (N_16257,N_11028,N_12587);
nor U16258 (N_16258,N_11729,N_12661);
and U16259 (N_16259,N_14965,N_10063);
xnor U16260 (N_16260,N_11207,N_13573);
xnor U16261 (N_16261,N_10617,N_11979);
nor U16262 (N_16262,N_10497,N_10739);
nor U16263 (N_16263,N_10716,N_14986);
nor U16264 (N_16264,N_11816,N_10895);
nand U16265 (N_16265,N_13867,N_13075);
or U16266 (N_16266,N_12500,N_11830);
or U16267 (N_16267,N_11475,N_10402);
xor U16268 (N_16268,N_13431,N_14894);
or U16269 (N_16269,N_11274,N_12845);
xnor U16270 (N_16270,N_12025,N_12631);
or U16271 (N_16271,N_11915,N_11138);
and U16272 (N_16272,N_13404,N_12747);
xor U16273 (N_16273,N_13819,N_12403);
and U16274 (N_16274,N_11091,N_13336);
or U16275 (N_16275,N_13169,N_14432);
and U16276 (N_16276,N_12653,N_12507);
nand U16277 (N_16277,N_11136,N_12359);
nand U16278 (N_16278,N_14578,N_10255);
nor U16279 (N_16279,N_10861,N_13731);
nor U16280 (N_16280,N_10502,N_11171);
and U16281 (N_16281,N_12732,N_12572);
and U16282 (N_16282,N_14146,N_10736);
nand U16283 (N_16283,N_12718,N_11908);
nor U16284 (N_16284,N_10626,N_12559);
xnor U16285 (N_16285,N_12770,N_13988);
and U16286 (N_16286,N_13209,N_12949);
nor U16287 (N_16287,N_12032,N_12321);
nand U16288 (N_16288,N_11621,N_10374);
nand U16289 (N_16289,N_14129,N_11772);
xnor U16290 (N_16290,N_11240,N_14953);
nand U16291 (N_16291,N_11107,N_10879);
nor U16292 (N_16292,N_12840,N_13237);
xnor U16293 (N_16293,N_10656,N_14915);
nor U16294 (N_16294,N_14197,N_12936);
xnor U16295 (N_16295,N_11490,N_12570);
nor U16296 (N_16296,N_12514,N_14781);
and U16297 (N_16297,N_14384,N_12857);
or U16298 (N_16298,N_10507,N_10669);
nand U16299 (N_16299,N_14860,N_12987);
nor U16300 (N_16300,N_13991,N_10002);
and U16301 (N_16301,N_14234,N_12291);
or U16302 (N_16302,N_12619,N_11889);
nor U16303 (N_16303,N_10583,N_11549);
nor U16304 (N_16304,N_13717,N_14287);
nor U16305 (N_16305,N_12235,N_11415);
and U16306 (N_16306,N_13617,N_10329);
nor U16307 (N_16307,N_10730,N_14301);
xor U16308 (N_16308,N_10108,N_14926);
and U16309 (N_16309,N_11363,N_13784);
and U16310 (N_16310,N_11380,N_13940);
xor U16311 (N_16311,N_10228,N_13086);
xor U16312 (N_16312,N_14766,N_10133);
xnor U16313 (N_16313,N_13163,N_13677);
or U16314 (N_16314,N_12804,N_12923);
or U16315 (N_16315,N_13495,N_13745);
and U16316 (N_16316,N_12130,N_13467);
xnor U16317 (N_16317,N_11570,N_10343);
nand U16318 (N_16318,N_14314,N_12729);
and U16319 (N_16319,N_12967,N_12401);
xor U16320 (N_16320,N_10598,N_14183);
nand U16321 (N_16321,N_11018,N_12649);
nor U16322 (N_16322,N_10506,N_11146);
nand U16323 (N_16323,N_11435,N_14160);
nor U16324 (N_16324,N_13131,N_10762);
nand U16325 (N_16325,N_13652,N_13598);
nand U16326 (N_16326,N_10203,N_10535);
nor U16327 (N_16327,N_11852,N_14812);
and U16328 (N_16328,N_11287,N_14487);
and U16329 (N_16329,N_12665,N_13265);
or U16330 (N_16330,N_14127,N_12603);
and U16331 (N_16331,N_14413,N_12777);
and U16332 (N_16332,N_10957,N_12271);
and U16333 (N_16333,N_13729,N_12353);
xnor U16334 (N_16334,N_11436,N_13948);
nor U16335 (N_16335,N_12464,N_12781);
nand U16336 (N_16336,N_12986,N_10112);
or U16337 (N_16337,N_11718,N_11412);
xnor U16338 (N_16338,N_10795,N_12251);
nand U16339 (N_16339,N_14698,N_11374);
and U16340 (N_16340,N_14783,N_12476);
or U16341 (N_16341,N_11714,N_12817);
nand U16342 (N_16342,N_12633,N_12696);
xor U16343 (N_16343,N_12430,N_14876);
nor U16344 (N_16344,N_12955,N_12785);
nand U16345 (N_16345,N_10921,N_13656);
xnor U16346 (N_16346,N_11548,N_12764);
nand U16347 (N_16347,N_13267,N_13525);
nor U16348 (N_16348,N_13355,N_13537);
or U16349 (N_16349,N_12221,N_13266);
or U16350 (N_16350,N_14618,N_13883);
or U16351 (N_16351,N_12697,N_14133);
nor U16352 (N_16352,N_14535,N_13629);
and U16353 (N_16353,N_14072,N_12494);
nor U16354 (N_16354,N_10011,N_10833);
and U16355 (N_16355,N_10874,N_11821);
and U16356 (N_16356,N_14716,N_10337);
nor U16357 (N_16357,N_12962,N_12106);
xor U16358 (N_16358,N_10898,N_12087);
xor U16359 (N_16359,N_14755,N_11218);
xnor U16360 (N_16360,N_10546,N_10677);
and U16361 (N_16361,N_10604,N_14409);
xor U16362 (N_16362,N_11245,N_12908);
nor U16363 (N_16363,N_14563,N_14690);
nor U16364 (N_16364,N_11372,N_11371);
nor U16365 (N_16365,N_14792,N_12356);
or U16366 (N_16366,N_11462,N_13515);
xor U16367 (N_16367,N_14021,N_10689);
xnor U16368 (N_16368,N_10001,N_12605);
or U16369 (N_16369,N_12205,N_12360);
nor U16370 (N_16370,N_11265,N_10569);
nand U16371 (N_16371,N_10746,N_13248);
nand U16372 (N_16372,N_10214,N_11909);
and U16373 (N_16373,N_11940,N_11092);
nor U16374 (N_16374,N_14063,N_11645);
nor U16375 (N_16375,N_11319,N_13085);
nor U16376 (N_16376,N_11805,N_10731);
nor U16377 (N_16377,N_11329,N_10427);
xnor U16378 (N_16378,N_11421,N_13599);
nand U16379 (N_16379,N_13376,N_11342);
and U16380 (N_16380,N_11627,N_13299);
and U16381 (N_16381,N_10494,N_12174);
xor U16382 (N_16382,N_14376,N_10264);
nand U16383 (N_16383,N_14497,N_10945);
nor U16384 (N_16384,N_10250,N_13401);
or U16385 (N_16385,N_12580,N_14452);
and U16386 (N_16386,N_13015,N_10764);
nand U16387 (N_16387,N_11054,N_14436);
or U16388 (N_16388,N_13805,N_11480);
or U16389 (N_16389,N_13975,N_14866);
xnor U16390 (N_16390,N_12685,N_14048);
xor U16391 (N_16391,N_13122,N_12478);
or U16392 (N_16392,N_13339,N_12828);
xor U16393 (N_16393,N_11333,N_14536);
or U16394 (N_16394,N_10832,N_13092);
and U16395 (N_16395,N_14044,N_12491);
nor U16396 (N_16396,N_14547,N_12760);
and U16397 (N_16397,N_14141,N_11434);
nand U16398 (N_16398,N_10653,N_14359);
or U16399 (N_16399,N_10102,N_12965);
or U16400 (N_16400,N_12003,N_13313);
or U16401 (N_16401,N_11446,N_11906);
or U16402 (N_16402,N_13591,N_10146);
nand U16403 (N_16403,N_13659,N_11579);
nor U16404 (N_16404,N_11023,N_13623);
nor U16405 (N_16405,N_11674,N_12283);
and U16406 (N_16406,N_13877,N_10266);
or U16407 (N_16407,N_10828,N_14064);
xor U16408 (N_16408,N_14977,N_13802);
or U16409 (N_16409,N_14086,N_13282);
nor U16410 (N_16410,N_13615,N_12681);
nor U16411 (N_16411,N_10859,N_14723);
nor U16412 (N_16412,N_13124,N_13767);
nor U16413 (N_16413,N_11007,N_13108);
xnor U16414 (N_16414,N_13215,N_13243);
xor U16415 (N_16415,N_10912,N_13468);
and U16416 (N_16416,N_14803,N_12168);
and U16417 (N_16417,N_14633,N_11231);
nand U16418 (N_16418,N_14425,N_10349);
nand U16419 (N_16419,N_14485,N_10430);
and U16420 (N_16420,N_10816,N_14109);
nand U16421 (N_16421,N_11644,N_13586);
xor U16422 (N_16422,N_10493,N_13601);
nor U16423 (N_16423,N_10513,N_14545);
nor U16424 (N_16424,N_14346,N_13277);
xor U16425 (N_16425,N_14632,N_10903);
xor U16426 (N_16426,N_11677,N_10899);
and U16427 (N_16427,N_11201,N_11344);
nor U16428 (N_16428,N_12875,N_14324);
or U16429 (N_16429,N_11782,N_13183);
nor U16430 (N_16430,N_13918,N_11469);
or U16431 (N_16431,N_10070,N_13139);
xnor U16432 (N_16432,N_10333,N_13110);
and U16433 (N_16433,N_14102,N_12268);
or U16434 (N_16434,N_14463,N_14274);
and U16435 (N_16435,N_12650,N_11320);
and U16436 (N_16436,N_13627,N_10447);
xnor U16437 (N_16437,N_11124,N_13113);
or U16438 (N_16438,N_13943,N_14239);
and U16439 (N_16439,N_12436,N_10672);
nand U16440 (N_16440,N_10664,N_12138);
xor U16441 (N_16441,N_14802,N_12092);
and U16442 (N_16442,N_12470,N_13394);
nor U16443 (N_16443,N_11642,N_12519);
xnor U16444 (N_16444,N_14367,N_12827);
nand U16445 (N_16445,N_13367,N_13203);
or U16446 (N_16446,N_13837,N_12796);
and U16447 (N_16447,N_10320,N_11399);
nand U16448 (N_16448,N_12700,N_14215);
nand U16449 (N_16449,N_13923,N_12088);
or U16450 (N_16450,N_11296,N_12295);
nor U16451 (N_16451,N_13164,N_14347);
xnor U16452 (N_16452,N_14744,N_14149);
and U16453 (N_16453,N_12469,N_10906);
xor U16454 (N_16454,N_12556,N_11941);
nand U16455 (N_16455,N_12022,N_11593);
and U16456 (N_16456,N_14480,N_11327);
or U16457 (N_16457,N_14430,N_14930);
or U16458 (N_16458,N_11293,N_13422);
nor U16459 (N_16459,N_10951,N_13385);
and U16460 (N_16460,N_13769,N_10327);
nor U16461 (N_16461,N_10127,N_13478);
and U16462 (N_16462,N_12607,N_11225);
and U16463 (N_16463,N_13218,N_12711);
nor U16464 (N_16464,N_12344,N_14342);
and U16465 (N_16465,N_11832,N_13320);
nor U16466 (N_16466,N_11306,N_11745);
nand U16467 (N_16467,N_11425,N_13798);
nor U16468 (N_16468,N_13597,N_10336);
nand U16469 (N_16469,N_14047,N_14131);
or U16470 (N_16470,N_12961,N_14711);
nand U16471 (N_16471,N_14606,N_11695);
and U16472 (N_16472,N_10962,N_10166);
nand U16473 (N_16473,N_10940,N_12985);
nor U16474 (N_16474,N_10931,N_12958);
nand U16475 (N_16475,N_13328,N_12049);
or U16476 (N_16476,N_11517,N_12811);
and U16477 (N_16477,N_11133,N_14599);
nand U16478 (N_16478,N_12067,N_11168);
and U16479 (N_16479,N_13879,N_10229);
xnor U16480 (N_16480,N_12660,N_11892);
nand U16481 (N_16481,N_14356,N_14178);
nand U16482 (N_16482,N_13751,N_12292);
nand U16483 (N_16483,N_11016,N_14403);
or U16484 (N_16484,N_11541,N_11877);
xnor U16485 (N_16485,N_14075,N_12994);
xnor U16486 (N_16486,N_13967,N_14813);
xor U16487 (N_16487,N_14703,N_13814);
or U16488 (N_16488,N_10042,N_10435);
or U16489 (N_16489,N_12423,N_10054);
nand U16490 (N_16490,N_14682,N_11501);
nand U16491 (N_16491,N_12854,N_11843);
nor U16492 (N_16492,N_11375,N_14370);
xnor U16493 (N_16493,N_13772,N_12882);
and U16494 (N_16494,N_14809,N_13982);
and U16495 (N_16495,N_13162,N_12852);
or U16496 (N_16496,N_14212,N_13338);
and U16497 (N_16497,N_13469,N_10147);
or U16498 (N_16498,N_14871,N_14268);
nor U16499 (N_16499,N_14208,N_10143);
nand U16500 (N_16500,N_10659,N_11418);
or U16501 (N_16501,N_12419,N_10987);
nor U16502 (N_16502,N_14734,N_11861);
or U16503 (N_16503,N_11401,N_12895);
nand U16504 (N_16504,N_12708,N_12613);
nor U16505 (N_16505,N_10968,N_11129);
nand U16506 (N_16506,N_12111,N_13305);
and U16507 (N_16507,N_14283,N_12113);
xor U16508 (N_16508,N_14475,N_12452);
nor U16509 (N_16509,N_10515,N_11235);
and U16510 (N_16510,N_10448,N_10106);
and U16511 (N_16511,N_10636,N_11134);
xor U16512 (N_16512,N_13543,N_11795);
and U16513 (N_16513,N_14543,N_14055);
nor U16514 (N_16514,N_13939,N_13737);
nor U16515 (N_16515,N_12684,N_12834);
nand U16516 (N_16516,N_12112,N_13175);
and U16517 (N_16517,N_11807,N_13022);
nand U16518 (N_16518,N_10814,N_14213);
and U16519 (N_16519,N_13310,N_12282);
xnor U16520 (N_16520,N_14051,N_14750);
nand U16521 (N_16521,N_13361,N_13137);
xor U16522 (N_16522,N_10511,N_11819);
and U16523 (N_16523,N_11473,N_11268);
xor U16524 (N_16524,N_10137,N_14837);
nand U16525 (N_16525,N_10517,N_12045);
xnor U16526 (N_16526,N_12455,N_13838);
nand U16527 (N_16527,N_12836,N_12595);
and U16528 (N_16528,N_11034,N_12157);
xnor U16529 (N_16529,N_11381,N_14899);
and U16530 (N_16530,N_11288,N_14625);
nor U16531 (N_16531,N_11455,N_14289);
nand U16532 (N_16532,N_13964,N_10510);
xnor U16533 (N_16533,N_13576,N_12449);
nor U16534 (N_16534,N_13324,N_14443);
nand U16535 (N_16535,N_13794,N_13980);
or U16536 (N_16536,N_12352,N_10667);
nor U16537 (N_16537,N_11793,N_11048);
xor U16538 (N_16538,N_13158,N_10366);
and U16539 (N_16539,N_14416,N_14865);
nor U16540 (N_16540,N_14591,N_13353);
or U16541 (N_16541,N_14756,N_13987);
or U16542 (N_16542,N_14261,N_12421);
nor U16543 (N_16543,N_10480,N_13452);
nor U16544 (N_16544,N_13534,N_13551);
and U16545 (N_16545,N_13063,N_13043);
nand U16546 (N_16546,N_11085,N_13200);
xnor U16547 (N_16547,N_14172,N_10408);
and U16548 (N_16548,N_11787,N_10973);
nor U16549 (N_16549,N_11376,N_14941);
or U16550 (N_16550,N_11205,N_10983);
and U16551 (N_16551,N_14706,N_10721);
nor U16552 (N_16552,N_11975,N_14216);
nor U16553 (N_16553,N_13728,N_13954);
and U16554 (N_16554,N_12485,N_14947);
and U16555 (N_16555,N_10826,N_10309);
xor U16556 (N_16556,N_14288,N_12448);
xor U16557 (N_16557,N_12034,N_10862);
and U16558 (N_16558,N_10109,N_11930);
or U16559 (N_16559,N_10638,N_11707);
nor U16560 (N_16560,N_13864,N_11854);
and U16561 (N_16561,N_12418,N_14936);
or U16562 (N_16562,N_11592,N_14583);
nor U16563 (N_16563,N_10870,N_10101);
nand U16564 (N_16564,N_11781,N_11451);
xor U16565 (N_16565,N_12579,N_10965);
xor U16566 (N_16566,N_12733,N_14386);
nand U16567 (N_16567,N_11800,N_14029);
nor U16568 (N_16568,N_12358,N_13851);
or U16569 (N_16569,N_10854,N_14206);
or U16570 (N_16570,N_14526,N_11968);
and U16571 (N_16571,N_13421,N_12373);
and U16572 (N_16572,N_14978,N_12059);
and U16573 (N_16573,N_14534,N_13557);
nand U16574 (N_16574,N_10997,N_10312);
nand U16575 (N_16575,N_13239,N_12035);
nand U16576 (N_16576,N_13028,N_11108);
xnor U16577 (N_16577,N_10780,N_10999);
or U16578 (N_16578,N_14011,N_12585);
xor U16579 (N_16579,N_10224,N_11750);
nand U16580 (N_16580,N_13555,N_13212);
nand U16581 (N_16581,N_14498,N_10723);
xnor U16582 (N_16582,N_11233,N_10560);
xnor U16583 (N_16583,N_12999,N_11120);
and U16584 (N_16584,N_13128,N_12995);
nand U16585 (N_16585,N_11321,N_11658);
or U16586 (N_16586,N_10735,N_12988);
or U16587 (N_16587,N_14826,N_14180);
nor U16588 (N_16588,N_10222,N_11284);
xor U16589 (N_16589,N_14829,N_14366);
nand U16590 (N_16590,N_13607,N_11135);
nand U16591 (N_16591,N_11666,N_11606);
or U16592 (N_16592,N_12408,N_10350);
nand U16593 (N_16593,N_14256,N_13977);
nand U16594 (N_16594,N_10219,N_11452);
nand U16595 (N_16595,N_14893,N_14205);
xor U16596 (N_16596,N_12540,N_13781);
nand U16597 (N_16597,N_13791,N_12101);
xor U16598 (N_16598,N_12144,N_14702);
nor U16599 (N_16599,N_11766,N_10334);
and U16600 (N_16600,N_14613,N_12768);
nor U16601 (N_16601,N_10759,N_13312);
or U16602 (N_16602,N_13470,N_11070);
nand U16603 (N_16603,N_10038,N_10804);
nand U16604 (N_16604,N_13913,N_12735);
nand U16605 (N_16605,N_13400,N_12644);
or U16606 (N_16606,N_12787,N_11299);
or U16607 (N_16607,N_11828,N_14148);
nor U16608 (N_16608,N_11813,N_10676);
nand U16609 (N_16609,N_13213,N_13642);
xnor U16610 (N_16610,N_13331,N_10328);
nand U16611 (N_16611,N_14721,N_12264);
nand U16612 (N_16612,N_14507,N_10779);
xnor U16613 (N_16613,N_11961,N_13933);
or U16614 (N_16614,N_10834,N_13554);
xor U16615 (N_16615,N_10322,N_11326);
and U16616 (N_16616,N_14053,N_14400);
nor U16617 (N_16617,N_11612,N_11281);
xnor U16618 (N_16618,N_11740,N_14276);
and U16619 (N_16619,N_12743,N_12196);
nor U16620 (N_16620,N_12704,N_14641);
nor U16621 (N_16621,N_13411,N_10254);
nand U16622 (N_16622,N_11315,N_12746);
nand U16623 (N_16623,N_10173,N_10883);
and U16624 (N_16624,N_12089,N_13281);
and U16625 (N_16625,N_11114,N_11082);
and U16626 (N_16626,N_13930,N_12575);
and U16627 (N_16627,N_12805,N_13567);
and U16628 (N_16628,N_14810,N_11176);
xnor U16629 (N_16629,N_14317,N_10315);
and U16630 (N_16630,N_11737,N_14493);
xnor U16631 (N_16631,N_14298,N_14423);
xor U16632 (N_16632,N_10985,N_13074);
xor U16633 (N_16633,N_10453,N_14304);
nand U16634 (N_16634,N_13833,N_11863);
xnor U16635 (N_16635,N_14486,N_13029);
nor U16636 (N_16636,N_13269,N_13405);
xor U16637 (N_16637,N_14959,N_14877);
or U16638 (N_16638,N_11266,N_13202);
nand U16639 (N_16639,N_14906,N_13114);
xnor U16640 (N_16640,N_11332,N_14407);
xor U16641 (N_16641,N_11459,N_10469);
xnor U16642 (N_16642,N_11482,N_11027);
nor U16643 (N_16643,N_13007,N_13453);
and U16644 (N_16644,N_14499,N_13647);
and U16645 (N_16645,N_14154,N_12576);
nand U16646 (N_16646,N_11309,N_13314);
nand U16647 (N_16647,N_13832,N_11905);
or U16648 (N_16648,N_13483,N_10603);
or U16649 (N_16649,N_10306,N_10205);
nor U16650 (N_16650,N_11247,N_13220);
or U16651 (N_16651,N_12322,N_11564);
xnor U16652 (N_16652,N_11688,N_12510);
xor U16653 (N_16653,N_12281,N_11585);
nor U16654 (N_16654,N_13418,N_13446);
nand U16655 (N_16655,N_10712,N_13895);
nand U16656 (N_16656,N_13037,N_14070);
nand U16657 (N_16657,N_11142,N_14189);
and U16658 (N_16658,N_14444,N_12623);
xor U16659 (N_16659,N_10227,N_10158);
nand U16660 (N_16660,N_12610,N_10272);
xor U16661 (N_16661,N_10010,N_10678);
nor U16662 (N_16662,N_11345,N_12984);
or U16663 (N_16663,N_11166,N_12050);
or U16664 (N_16664,N_10773,N_14735);
nand U16665 (N_16665,N_11341,N_14357);
or U16666 (N_16666,N_13308,N_12564);
nor U16667 (N_16667,N_13773,N_11021);
nand U16668 (N_16668,N_11069,N_13637);
nand U16669 (N_16669,N_14318,N_13134);
and U16670 (N_16670,N_10196,N_13609);
or U16671 (N_16671,N_10846,N_14945);
or U16672 (N_16672,N_14037,N_14340);
xnor U16673 (N_16673,N_12074,N_12616);
nor U16674 (N_16674,N_11077,N_12763);
or U16675 (N_16675,N_12651,N_11880);
nand U16676 (N_16676,N_13492,N_12182);
xnor U16677 (N_16677,N_10107,N_14657);
and U16678 (N_16678,N_10584,N_10557);
or U16679 (N_16679,N_13156,N_13024);
and U16680 (N_16680,N_10330,N_10980);
nand U16681 (N_16681,N_11960,N_14300);
nor U16682 (N_16682,N_12169,N_14675);
and U16683 (N_16683,N_10027,N_11528);
or U16684 (N_16684,N_13181,N_11302);
nor U16685 (N_16685,N_11053,N_11105);
or U16686 (N_16686,N_11865,N_12754);
nand U16687 (N_16687,N_13841,N_12879);
nor U16688 (N_16688,N_12302,N_11063);
nand U16689 (N_16689,N_12680,N_10093);
nor U16690 (N_16690,N_13763,N_11945);
nor U16691 (N_16691,N_12274,N_11143);
and U16692 (N_16692,N_10367,N_12990);
xor U16693 (N_16693,N_12393,N_13460);
nor U16694 (N_16694,N_13009,N_14856);
nand U16695 (N_16695,N_12938,N_12231);
nand U16696 (N_16696,N_10688,N_12457);
xnor U16697 (N_16697,N_12693,N_10817);
or U16698 (N_16698,N_14321,N_12802);
nor U16699 (N_16699,N_11931,N_10190);
nor U16700 (N_16700,N_13521,N_13025);
nand U16701 (N_16701,N_14726,N_14083);
and U16702 (N_16702,N_10637,N_11495);
nor U16703 (N_16703,N_11348,N_10298);
xor U16704 (N_16704,N_11713,N_11497);
and U16705 (N_16705,N_10404,N_10726);
nor U16706 (N_16706,N_14078,N_14540);
and U16707 (N_16707,N_13135,N_12599);
and U16708 (N_16708,N_10341,N_13630);
or U16709 (N_16709,N_11242,N_10593);
and U16710 (N_16710,N_13010,N_12390);
nand U16711 (N_16711,N_13101,N_10433);
or U16712 (N_16712,N_11837,N_11009);
nor U16713 (N_16713,N_14954,N_13493);
or U16714 (N_16714,N_10177,N_10851);
nand U16715 (N_16715,N_12525,N_14542);
nand U16716 (N_16716,N_10761,N_13403);
or U16717 (N_16717,N_12825,N_11423);
and U16718 (N_16718,N_10204,N_12960);
xnor U16719 (N_16719,N_12442,N_13583);
nor U16720 (N_16720,N_13219,N_11147);
or U16721 (N_16721,N_10718,N_12658);
or U16722 (N_16722,N_13123,N_13921);
xor U16723 (N_16723,N_11763,N_14593);
and U16724 (N_16724,N_11256,N_11667);
xor U16725 (N_16725,N_14828,N_12095);
xnor U16726 (N_16726,N_11046,N_10331);
and U16727 (N_16727,N_13633,N_11170);
nand U16728 (N_16728,N_12041,N_14451);
and U16729 (N_16729,N_13464,N_13368);
and U16730 (N_16730,N_12784,N_14863);
or U16731 (N_16731,N_13423,N_11402);
and U16732 (N_16732,N_12766,N_11003);
nor U16733 (N_16733,N_13083,N_13259);
and U16734 (N_16734,N_14602,N_11581);
or U16735 (N_16735,N_14889,N_12752);
and U16736 (N_16736,N_14259,N_14571);
and U16737 (N_16737,N_12007,N_13119);
xnor U16738 (N_16738,N_12687,N_11202);
nand U16739 (N_16739,N_10777,N_14673);
nand U16740 (N_16740,N_13885,N_12744);
nor U16741 (N_16741,N_11167,N_10972);
nor U16742 (N_16742,N_13562,N_10662);
xnor U16743 (N_16743,N_12615,N_13207);
nor U16744 (N_16744,N_11200,N_14680);
nand U16745 (N_16745,N_14296,N_10098);
xor U16746 (N_16746,N_10842,N_14582);
and U16747 (N_16747,N_11126,N_14560);
or U16748 (N_16748,N_13828,N_14229);
and U16749 (N_16749,N_11384,N_14372);
nor U16750 (N_16750,N_12826,N_13323);
or U16751 (N_16751,N_11853,N_10481);
nor U16752 (N_16752,N_10897,N_12563);
nor U16753 (N_16753,N_11802,N_10104);
or U16754 (N_16754,N_13755,N_11254);
xor U16755 (N_16755,N_10476,N_14983);
or U16756 (N_16756,N_14670,N_12397);
nand U16757 (N_16757,N_12794,N_12207);
or U16758 (N_16758,N_13566,N_10799);
and U16759 (N_16759,N_13900,N_11340);
xor U16760 (N_16760,N_10943,N_13788);
nor U16761 (N_16761,N_11153,N_10084);
xnor U16762 (N_16762,N_11080,N_13352);
or U16763 (N_16763,N_14878,N_12634);
nand U16764 (N_16764,N_11013,N_14637);
and U16765 (N_16765,N_14374,N_12116);
and U16766 (N_16766,N_11550,N_10045);
or U16767 (N_16767,N_14202,N_10407);
nand U16768 (N_16768,N_13294,N_12396);
or U16769 (N_16769,N_10221,N_13839);
or U16770 (N_16770,N_14859,N_10695);
nor U16771 (N_16771,N_14851,N_11762);
and U16772 (N_16772,N_14811,N_14910);
xnor U16773 (N_16773,N_13912,N_12865);
xnor U16774 (N_16774,N_11444,N_10124);
or U16775 (N_16775,N_12905,N_11901);
or U16776 (N_16776,N_14991,N_13825);
or U16777 (N_16777,N_10317,N_13622);
xor U16778 (N_16778,N_12630,N_12058);
or U16779 (N_16779,N_13995,N_12416);
and U16780 (N_16780,N_13888,N_12266);
nand U16781 (N_16781,N_12782,N_12394);
nor U16782 (N_16782,N_11654,N_14816);
nor U16783 (N_16783,N_10056,N_10413);
nand U16784 (N_16784,N_10390,N_14671);
and U16785 (N_16785,N_11601,N_14728);
or U16786 (N_16786,N_10352,N_13984);
and U16787 (N_16787,N_11097,N_10606);
nand U16788 (N_16788,N_11920,N_13863);
or U16789 (N_16789,N_13847,N_10186);
and U16790 (N_16790,N_14831,N_10062);
nand U16791 (N_16791,N_12707,N_12761);
nor U16792 (N_16792,N_10556,N_11537);
xnor U16793 (N_16793,N_14308,N_12383);
and U16794 (N_16794,N_13810,N_13047);
and U16795 (N_16795,N_13976,N_12369);
nand U16796 (N_16796,N_11043,N_13100);
or U16797 (N_16797,N_13109,N_11432);
or U16798 (N_16798,N_10690,N_12189);
xnor U16799 (N_16799,N_12876,N_10877);
or U16800 (N_16800,N_13377,N_12284);
nor U16801 (N_16801,N_12501,N_10401);
nand U16802 (N_16802,N_11724,N_12947);
or U16803 (N_16803,N_14975,N_10060);
and U16804 (N_16804,N_13366,N_10717);
xor U16805 (N_16805,N_12523,N_12272);
or U16806 (N_16806,N_14514,N_11972);
nand U16807 (N_16807,N_10284,N_10296);
nand U16808 (N_16808,N_11562,N_12276);
nand U16809 (N_16809,N_12319,N_11519);
and U16810 (N_16810,N_14352,N_10276);
nand U16811 (N_16811,N_11598,N_14277);
nand U16812 (N_16812,N_12513,N_10558);
nand U16813 (N_16813,N_12427,N_10499);
and U16814 (N_16814,N_12534,N_12980);
nand U16815 (N_16815,N_13249,N_14350);
nor U16816 (N_16816,N_14923,N_12877);
nor U16817 (N_16817,N_13786,N_14381);
and U16818 (N_16818,N_13646,N_14265);
and U16819 (N_16819,N_11511,N_10119);
nand U16820 (N_16820,N_12964,N_14258);
or U16821 (N_16821,N_13937,N_11734);
and U16822 (N_16822,N_12417,N_11031);
and U16823 (N_16823,N_12227,N_13782);
or U16824 (N_16824,N_12110,N_14576);
and U16825 (N_16825,N_12285,N_12612);
xnor U16826 (N_16826,N_11360,N_11675);
nand U16827 (N_16827,N_12699,N_13962);
nand U16828 (N_16828,N_12557,N_13477);
nor U16829 (N_16829,N_14494,N_12850);
and U16830 (N_16830,N_13034,N_13746);
nand U16831 (N_16831,N_10123,N_13536);
or U16832 (N_16832,N_10648,N_12531);
xor U16833 (N_16833,N_11823,N_12404);
nor U16834 (N_16834,N_14939,N_14145);
or U16835 (N_16835,N_13931,N_10588);
xor U16836 (N_16836,N_13223,N_14907);
xor U16837 (N_16837,N_11773,N_14244);
xnor U16838 (N_16838,N_11090,N_14782);
or U16839 (N_16839,N_12848,N_10193);
nand U16840 (N_16840,N_14912,N_12991);
nor U16841 (N_16841,N_12370,N_11449);
xnor U16842 (N_16842,N_14227,N_10223);
xor U16843 (N_16843,N_11102,N_10068);
nand U16844 (N_16844,N_10969,N_14387);
nand U16845 (N_16845,N_10500,N_13778);
nor U16846 (N_16846,N_10125,N_12326);
nor U16847 (N_16847,N_14045,N_13992);
nor U16848 (N_16848,N_14015,N_14088);
or U16849 (N_16849,N_12561,N_12645);
nand U16850 (N_16850,N_10831,N_11910);
or U16851 (N_16851,N_12715,N_10917);
and U16852 (N_16852,N_11826,N_10244);
or U16853 (N_16853,N_12931,N_10053);
xor U16854 (N_16854,N_14269,N_13649);
nand U16855 (N_16855,N_11116,N_11957);
nor U16856 (N_16856,N_12197,N_11337);
or U16857 (N_16857,N_12524,N_13914);
xnor U16858 (N_16858,N_14901,N_11769);
nor U16859 (N_16859,N_12195,N_11392);
nand U16860 (N_16860,N_14527,N_14688);
nand U16861 (N_16861,N_10996,N_13691);
and U16862 (N_16862,N_13482,N_14255);
and U16863 (N_16863,N_10967,N_11280);
and U16864 (N_16864,N_12884,N_12139);
or U16865 (N_16865,N_12293,N_10086);
nor U16866 (N_16866,N_10033,N_10233);
or U16867 (N_16867,N_13908,N_14948);
nand U16868 (N_16868,N_12378,N_10841);
nor U16869 (N_16869,N_11683,N_11364);
nand U16870 (N_16870,N_11993,N_12329);
nand U16871 (N_16871,N_13957,N_12277);
and U16872 (N_16872,N_12814,N_10935);
nand U16873 (N_16873,N_13425,N_14125);
and U16874 (N_16874,N_13549,N_14548);
nand U16875 (N_16875,N_10297,N_13638);
nand U16876 (N_16876,N_11073,N_10467);
nor U16877 (N_16877,N_10934,N_14504);
nand U16878 (N_16878,N_13358,N_12577);
nand U16879 (N_16879,N_13226,N_14839);
or U16880 (N_16880,N_11864,N_12327);
xnor U16881 (N_16881,N_12063,N_10624);
or U16882 (N_16882,N_11686,N_14164);
nand U16883 (N_16883,N_13517,N_14796);
and U16884 (N_16884,N_13606,N_11632);
or U16885 (N_16885,N_10783,N_14013);
xnor U16886 (N_16886,N_12503,N_10388);
and U16887 (N_16887,N_10302,N_12573);
nand U16888 (N_16888,N_11478,N_14218);
nand U16889 (N_16889,N_13061,N_12975);
xnor U16890 (N_16890,N_12107,N_11590);
and U16891 (N_16891,N_14752,N_10944);
nand U16892 (N_16892,N_14710,N_11992);
nand U16893 (N_16893,N_12026,N_11790);
and U16894 (N_16894,N_11275,N_13142);
nor U16895 (N_16895,N_13440,N_12090);
nor U16896 (N_16896,N_11359,N_13800);
nor U16897 (N_16897,N_11610,N_12071);
nor U16898 (N_16898,N_13020,N_13245);
and U16899 (N_16899,N_11953,N_13701);
nand U16900 (N_16900,N_11676,N_13117);
and U16901 (N_16901,N_12600,N_14938);
xnor U16902 (N_16902,N_14587,N_11862);
and U16903 (N_16903,N_11487,N_11619);
nand U16904 (N_16904,N_12028,N_12143);
and U16905 (N_16905,N_11835,N_13349);
nor U16906 (N_16906,N_14855,N_13332);
and U16907 (N_16907,N_12213,N_13174);
nor U16908 (N_16908,N_10885,N_10020);
xnor U16909 (N_16909,N_12602,N_10099);
xor U16910 (N_16910,N_11818,N_13779);
nand U16911 (N_16911,N_13398,N_11691);
xnor U16912 (N_16912,N_13018,N_12434);
and U16913 (N_16913,N_12226,N_14241);
nor U16914 (N_16914,N_14393,N_11159);
nand U16915 (N_16915,N_13547,N_13302);
or U16916 (N_16916,N_11236,N_12723);
and U16917 (N_16917,N_10843,N_10356);
nor U16918 (N_16918,N_13454,N_11944);
and U16919 (N_16919,N_11859,N_11998);
nor U16920 (N_16920,N_10575,N_11226);
nand U16921 (N_16921,N_14791,N_11324);
and U16922 (N_16922,N_10021,N_11424);
xor U16923 (N_16923,N_13953,N_13050);
and U16924 (N_16924,N_13136,N_12062);
nor U16925 (N_16925,N_14174,N_12569);
xnor U16926 (N_16926,N_14973,N_12386);
nand U16927 (N_16927,N_12609,N_11786);
xor U16928 (N_16928,N_10803,N_10064);
nand U16929 (N_16929,N_10474,N_11239);
nand U16930 (N_16930,N_13862,N_12917);
or U16931 (N_16931,N_11770,N_14415);
nor U16932 (N_16932,N_14262,N_14648);
nand U16933 (N_16933,N_14138,N_12215);
nor U16934 (N_16934,N_14121,N_13330);
nor U16935 (N_16935,N_13927,N_14396);
and U16936 (N_16936,N_10424,N_11173);
nor U16937 (N_16937,N_14490,N_12068);
and U16938 (N_16938,N_13886,N_12338);
nand U16939 (N_16939,N_13762,N_10009);
xor U16940 (N_16940,N_12288,N_14891);
and U16941 (N_16941,N_10582,N_14883);
nand U16942 (N_16942,N_12303,N_11741);
nand U16943 (N_16943,N_10018,N_14929);
nand U16944 (N_16944,N_13679,N_10840);
and U16945 (N_16945,N_10528,N_11661);
nand U16946 (N_16946,N_11428,N_14898);
xor U16947 (N_16947,N_13118,N_11118);
or U16948 (N_16948,N_12832,N_11187);
or U16949 (N_16949,N_10498,N_14000);
xor U16950 (N_16950,N_12289,N_14267);
and U16951 (N_16951,N_13850,N_14421);
nand U16952 (N_16952,N_14595,N_13749);
nand U16953 (N_16953,N_13682,N_10639);
xor U16954 (N_16954,N_11833,N_11378);
xnor U16955 (N_16955,N_11990,N_11743);
and U16956 (N_16956,N_14038,N_13000);
and U16957 (N_16957,N_12444,N_10161);
and U16958 (N_16958,N_14173,N_14908);
nor U16959 (N_16959,N_10442,N_13952);
or U16960 (N_16960,N_11172,N_13983);
or U16961 (N_16961,N_12904,N_13275);
or U16962 (N_16962,N_13796,N_12567);
nand U16963 (N_16963,N_14500,N_10995);
and U16964 (N_16964,N_11067,N_10608);
xor U16965 (N_16965,N_10410,N_12425);
nor U16966 (N_16966,N_10567,N_14886);
or U16967 (N_16967,N_10041,N_10602);
nand U16968 (N_16968,N_10262,N_14979);
nor U16969 (N_16969,N_12830,N_14659);
and U16970 (N_16970,N_13048,N_11089);
nand U16971 (N_16971,N_11716,N_13736);
nor U16972 (N_16972,N_11587,N_12915);
xor U16973 (N_16973,N_12637,N_12916);
nand U16974 (N_16974,N_13087,N_14943);
nand U16975 (N_16975,N_14957,N_11260);
nor U16976 (N_16976,N_14731,N_13541);
or U16977 (N_16977,N_10046,N_12702);
nor U16978 (N_16978,N_10625,N_11486);
or U16979 (N_16979,N_11058,N_12838);
and U16980 (N_16980,N_14207,N_13485);
and U16981 (N_16981,N_13268,N_13823);
nand U16982 (N_16982,N_10319,N_14981);
or U16983 (N_16983,N_12129,N_11379);
and U16984 (N_16984,N_12530,N_11696);
and U16985 (N_16985,N_10314,N_13415);
nor U16986 (N_16986,N_11894,N_10597);
nor U16987 (N_16987,N_10568,N_11221);
nor U16988 (N_16988,N_12466,N_14922);
or U16989 (N_16989,N_13575,N_10860);
and U16990 (N_16990,N_13264,N_13437);
and U16991 (N_16991,N_10787,N_11885);
or U16992 (N_16992,N_10162,N_12883);
xor U16993 (N_16993,N_11922,N_11325);
or U16994 (N_16994,N_14817,N_14508);
and U16995 (N_16995,N_13149,N_13026);
nor U16996 (N_16996,N_12484,N_14331);
nor U16997 (N_16997,N_10275,N_12797);
and U16998 (N_16998,N_14882,N_14358);
nor U16999 (N_16999,N_14777,N_14328);
nand U17000 (N_17000,N_10647,N_11967);
nand U17001 (N_17001,N_11285,N_11812);
and U17002 (N_17002,N_13621,N_10163);
nor U17003 (N_17003,N_13360,N_10292);
and U17004 (N_17004,N_11956,N_13233);
nor U17005 (N_17005,N_12415,N_14614);
xnor U17006 (N_17006,N_12617,N_14715);
or U17007 (N_17007,N_13046,N_12716);
nand U17008 (N_17008,N_14605,N_11643);
xnor U17009 (N_17009,N_13843,N_10265);
nor U17010 (N_17010,N_13540,N_13777);
and U17011 (N_17011,N_12471,N_14608);
nand U17012 (N_17012,N_11505,N_11584);
and U17013 (N_17013,N_11468,N_12528);
nand U17014 (N_17014,N_12414,N_13518);
nand U17015 (N_17015,N_12888,N_14091);
and U17016 (N_17016,N_12846,N_10115);
nand U17017 (N_17017,N_14203,N_12932);
or U17018 (N_17018,N_13471,N_12249);
nand U17019 (N_17019,N_14033,N_13457);
nor U17020 (N_17020,N_10992,N_12966);
nor U17021 (N_17021,N_13060,N_11411);
nor U17022 (N_17022,N_12218,N_13463);
nor U17023 (N_17023,N_10891,N_14835);
or U17024 (N_17024,N_13520,N_12040);
xnor U17025 (N_17025,N_11229,N_14567);
and U17026 (N_17026,N_13057,N_14263);
nand U17027 (N_17027,N_11237,N_14391);
nor U17028 (N_17028,N_11948,N_10769);
or U17029 (N_17029,N_10621,N_10409);
nand U17030 (N_17030,N_12589,N_13792);
and U17031 (N_17031,N_11924,N_11618);
xor U17032 (N_17032,N_13434,N_13760);
and U17033 (N_17033,N_12372,N_14840);
and U17034 (N_17034,N_12000,N_13628);
xor U17035 (N_17035,N_14065,N_12010);
and U17036 (N_17036,N_12675,N_14439);
xor U17037 (N_17037,N_13157,N_12056);
xnor U17038 (N_17038,N_12734,N_12779);
nor U17039 (N_17039,N_14081,N_11180);
and U17040 (N_17040,N_12230,N_12492);
and U17041 (N_17041,N_11539,N_10245);
nand U17042 (N_17042,N_11243,N_13283);
or U17043 (N_17043,N_12543,N_12046);
xnor U17044 (N_17044,N_14950,N_12515);
nand U17045 (N_17045,N_14658,N_13722);
nor U17046 (N_17046,N_13146,N_10562);
and U17047 (N_17047,N_11520,N_13545);
nand U17048 (N_17048,N_10512,N_13683);
and U17049 (N_17049,N_14963,N_12886);
nand U17050 (N_17050,N_11017,N_13451);
or U17051 (N_17051,N_13994,N_11298);
or U17052 (N_17052,N_13132,N_11036);
and U17053 (N_17053,N_11068,N_14297);
nand U17054 (N_17054,N_14914,N_11934);
nor U17055 (N_17055,N_11249,N_13616);
nand U17056 (N_17056,N_11162,N_10867);
or U17057 (N_17057,N_10852,N_14911);
nand U17058 (N_17058,N_12909,N_12398);
nor U17059 (N_17059,N_13410,N_11825);
nand U17060 (N_17060,N_14820,N_11059);
xor U17061 (N_17061,N_12307,N_11443);
and U17062 (N_17062,N_12146,N_12683);
nor U17063 (N_17063,N_14827,N_10378);
nor U17064 (N_17064,N_13090,N_10596);
and U17065 (N_17065,N_11294,N_10082);
nor U17066 (N_17066,N_12309,N_14179);
and U17067 (N_17067,N_13510,N_12454);
and U17068 (N_17068,N_10771,N_12668);
nand U17069 (N_17069,N_12030,N_13003);
nand U17070 (N_17070,N_11722,N_10150);
nand U17071 (N_17071,N_13972,N_14819);
xor U17072 (N_17072,N_11259,N_10239);
nor U17073 (N_17073,N_11751,N_12104);
nor U17074 (N_17074,N_14235,N_11145);
xor U17075 (N_17075,N_13216,N_14525);
nor U17076 (N_17076,N_11898,N_11177);
or U17077 (N_17077,N_11794,N_11653);
and U17078 (N_17078,N_13596,N_12346);
nand U17079 (N_17079,N_12717,N_12871);
and U17080 (N_17080,N_14544,N_11117);
xor U17081 (N_17081,N_11980,N_12304);
nand U17082 (N_17082,N_12153,N_13582);
nand U17083 (N_17083,N_10901,N_12047);
and U17084 (N_17084,N_11638,N_13664);
and U17085 (N_17085,N_14799,N_14834);
nor U17086 (N_17086,N_13238,N_12722);
nor U17087 (N_17087,N_11962,N_10657);
and U17088 (N_17088,N_12504,N_12385);
xor U17089 (N_17089,N_10849,N_10888);
nand U17090 (N_17090,N_12606,N_10156);
or U17091 (N_17091,N_11784,N_10729);
or U17092 (N_17092,N_10184,N_13280);
nor U17093 (N_17093,N_11981,N_10304);
xnor U17094 (N_17094,N_12269,N_12891);
xor U17095 (N_17095,N_13560,N_14720);
nor U17096 (N_17096,N_13569,N_11312);
nand U17097 (N_17097,N_11970,N_10910);
nand U17098 (N_17098,N_13387,N_11336);
nand U17099 (N_17099,N_11125,N_12407);
and U17100 (N_17100,N_10576,N_14424);
nand U17101 (N_17101,N_12462,N_12079);
xor U17102 (N_17102,N_14280,N_10559);
nor U17103 (N_17103,N_10592,N_12844);
nand U17104 (N_17104,N_14629,N_11614);
nor U17105 (N_17105,N_14252,N_10389);
and U17106 (N_17106,N_12120,N_14041);
nor U17107 (N_17107,N_13488,N_13657);
nand U17108 (N_17108,N_14068,N_14904);
xnor U17109 (N_17109,N_11806,N_14861);
nand U17110 (N_17110,N_12889,N_10955);
nand U17111 (N_17111,N_11512,N_14450);
nor U17112 (N_17112,N_13250,N_14195);
and U17113 (N_17113,N_13901,N_14776);
nand U17114 (N_17114,N_10240,N_11847);
xor U17115 (N_17115,N_12305,N_11277);
xnor U17116 (N_17116,N_12392,N_14375);
and U17117 (N_17117,N_13993,N_13070);
xor U17118 (N_17118,N_12400,N_10758);
or U17119 (N_17119,N_14533,N_13133);
nand U17120 (N_17120,N_14082,N_14066);
and U17121 (N_17121,N_11206,N_13073);
or U17122 (N_17122,N_10959,N_12626);
and U17123 (N_17123,N_12624,N_11174);
or U17124 (N_17124,N_10838,N_10251);
and U17125 (N_17125,N_10751,N_13379);
nor U17126 (N_17126,N_11271,N_13973);
and U17127 (N_17127,N_14530,N_14257);
and U17128 (N_17128,N_13298,N_10570);
xnor U17129 (N_17129,N_13205,N_10258);
xnor U17130 (N_17130,N_14209,N_11531);
and U17131 (N_17131,N_12807,N_10267);
or U17132 (N_17132,N_10595,N_13697);
xnor U17133 (N_17133,N_14913,N_10887);
and U17134 (N_17134,N_11181,N_14674);
nand U17135 (N_17135,N_12742,N_12705);
and U17136 (N_17136,N_14112,N_12813);
or U17137 (N_17137,N_13968,N_11841);
xor U17138 (N_17138,N_12077,N_12957);
nand U17139 (N_17139,N_12596,N_14147);
nor U17140 (N_17140,N_14974,N_14353);
or U17141 (N_17141,N_14844,N_10259);
nor U17142 (N_17142,N_14789,N_14002);
nor U17143 (N_17143,N_10725,N_14100);
or U17144 (N_17144,N_11307,N_12367);
and U17145 (N_17145,N_13378,N_13474);
xor U17146 (N_17146,N_14380,N_12084);
or U17147 (N_17147,N_11681,N_14917);
and U17148 (N_17148,N_14054,N_13327);
and U17149 (N_17149,N_14746,N_10080);
and U17150 (N_17150,N_11387,N_14484);
nand U17151 (N_17151,N_13229,N_14762);
nor U17152 (N_17152,N_10519,N_14446);
or U17153 (N_17153,N_11192,N_13626);
or U17154 (N_17154,N_14042,N_11532);
or U17155 (N_17155,N_10058,N_13391);
and U17156 (N_17156,N_13715,N_11591);
xor U17157 (N_17157,N_12447,N_10613);
nor U17158 (N_17158,N_10926,N_11339);
nor U17159 (N_17159,N_12643,N_13578);
or U17160 (N_17160,N_11572,N_10035);
and U17161 (N_17161,N_13062,N_14217);
and U17162 (N_17162,N_14036,N_10878);
nor U17163 (N_17163,N_14447,N_13187);
or U17164 (N_17164,N_11262,N_14440);
nor U17165 (N_17165,N_10437,N_13481);
or U17166 (N_17166,N_12536,N_14210);
or U17167 (N_17167,N_12109,N_12102);
xnor U17168 (N_17168,N_11217,N_13507);
nor U17169 (N_17169,N_10778,N_14892);
xnor U17170 (N_17170,N_14574,N_13733);
nand U17171 (N_17171,N_13530,N_11535);
and U17172 (N_17172,N_10023,N_11356);
nor U17173 (N_17173,N_10693,N_12934);
nand U17174 (N_17174,N_14105,N_10050);
and U17175 (N_17175,N_14853,N_10399);
xnor U17176 (N_17176,N_12237,N_11739);
xor U17177 (N_17177,N_12211,N_10332);
or U17178 (N_17178,N_10270,N_13346);
nor U17179 (N_17179,N_12395,N_10154);
nor U17180 (N_17180,N_13115,N_10805);
and U17181 (N_17181,N_11164,N_10673);
and U17182 (N_17182,N_14061,N_11951);
xor U17183 (N_17183,N_10610,N_13986);
or U17184 (N_17184,N_10873,N_11693);
nor U17185 (N_17185,N_14639,N_12873);
or U17186 (N_17186,N_14689,N_12568);
nand U17187 (N_17187,N_11626,N_11020);
or U17188 (N_17188,N_13752,N_12320);
or U17189 (N_17189,N_10117,N_13580);
and U17190 (N_17190,N_12765,N_10652);
nand U17191 (N_17191,N_13561,N_14448);
and U17192 (N_17192,N_10589,N_12974);
nor U17193 (N_17193,N_12306,N_10909);
nand U17194 (N_17194,N_12490,N_12973);
or U17195 (N_17195,N_10745,N_11767);
or U17196 (N_17196,N_12954,N_10457);
nand U17197 (N_17197,N_14972,N_14104);
and U17198 (N_17198,N_12406,N_10422);
nand U17199 (N_17199,N_14284,N_14344);
and U17200 (N_17200,N_10014,N_14874);
or U17201 (N_17201,N_11322,N_10396);
and U17202 (N_17202,N_11465,N_14243);
nor U17203 (N_17203,N_13225,N_10234);
or U17204 (N_17204,N_12902,N_14005);
and U17205 (N_17205,N_13105,N_11971);
nand U17206 (N_17206,N_12880,N_11600);
or U17207 (N_17207,N_13221,N_14565);
or U17208 (N_17208,N_10434,N_10183);
xnor U17209 (N_17209,N_14181,N_13764);
or U17210 (N_17210,N_11127,N_10937);
nand U17211 (N_17211,N_11659,N_11191);
xor U17212 (N_17212,N_12835,N_11684);
xor U17213 (N_17213,N_12384,N_11422);
and U17214 (N_17214,N_11798,N_14968);
xor U17215 (N_17215,N_13076,N_11586);
and U17216 (N_17216,N_11625,N_13641);
xnor U17217 (N_17217,N_13274,N_14248);
or U17218 (N_17218,N_14549,N_13260);
or U17219 (N_17219,N_11121,N_10821);
or U17220 (N_17220,N_11939,N_12581);
nor U17221 (N_17221,N_14778,N_12552);
or U17222 (N_17222,N_12793,N_14757);
nand U17223 (N_17223,N_13258,N_14167);
and U17224 (N_17224,N_10612,N_11596);
xor U17225 (N_17225,N_12126,N_10789);
and U17226 (N_17226,N_14470,N_14223);
nor U17227 (N_17227,N_10792,N_10120);
xor U17228 (N_17228,N_11995,N_11811);
and U17229 (N_17229,N_11086,N_13341);
xor U17230 (N_17230,N_14570,N_11904);
and U17231 (N_17231,N_12362,N_12141);
or U17232 (N_17232,N_11314,N_12013);
nor U17233 (N_17233,N_11896,N_14220);
xnor U17234 (N_17234,N_14868,N_12219);
or U17235 (N_17235,N_10032,N_11815);
nand U17236 (N_17236,N_14286,N_12148);
nand U17237 (N_17237,N_13849,N_14737);
and U17238 (N_17238,N_12280,N_12135);
and U17239 (N_17239,N_13184,N_11887);
nand U17240 (N_17240,N_11458,N_12331);
nor U17241 (N_17241,N_11308,N_10794);
nand U17242 (N_17242,N_10692,N_13095);
and U17243 (N_17243,N_12012,N_13155);
or U17244 (N_17244,N_10823,N_12979);
nand U17245 (N_17245,N_10800,N_14390);
nor U17246 (N_17246,N_12387,N_14237);
nand U17247 (N_17247,N_10663,N_12672);
xor U17248 (N_17248,N_12925,N_11454);
and U17249 (N_17249,N_13966,N_11414);
and U17250 (N_17250,N_10765,N_13201);
and U17251 (N_17251,N_12136,N_11093);
and U17252 (N_17252,N_14873,N_11269);
and U17253 (N_17253,N_12069,N_12187);
nand U17254 (N_17254,N_11347,N_11185);
and U17255 (N_17255,N_14382,N_14192);
xor U17256 (N_17256,N_14459,N_13017);
xor U17257 (N_17257,N_13234,N_13651);
or U17258 (N_17258,N_12241,N_10029);
nor U17259 (N_17259,N_12499,N_14319);
xnor U17260 (N_17260,N_14656,N_13665);
nor U17261 (N_17261,N_10785,N_13958);
nand U17262 (N_17262,N_10905,N_14326);
xnor U17263 (N_17263,N_14714,N_10111);
and U17264 (N_17264,N_12179,N_13426);
nand U17265 (N_17265,N_11169,N_12432);
nand U17266 (N_17266,N_10509,N_12435);
nand U17267 (N_17267,N_10368,N_10231);
nor U17268 (N_17268,N_12996,N_14481);
or U17269 (N_17269,N_13834,N_13429);
nor U17270 (N_17270,N_10455,N_11330);
nor U17271 (N_17271,N_13827,N_10075);
or U17272 (N_17272,N_13351,N_11851);
nor U17273 (N_17273,N_12778,N_11726);
nand U17274 (N_17274,N_11839,N_14115);
nor U17275 (N_17275,N_10198,N_12751);
nand U17276 (N_17276,N_12057,N_11123);
or U17277 (N_17277,N_12944,N_13012);
nor U17278 (N_17278,N_13436,N_11952);
and U17279 (N_17279,N_11568,N_13732);
nand U17280 (N_17280,N_13001,N_12167);
xnor U17281 (N_17281,N_11947,N_14155);
or U17282 (N_17282,N_10176,N_13286);
or U17283 (N_17283,N_11419,N_14992);
or U17284 (N_17284,N_12907,N_14293);
or U17285 (N_17285,N_12217,N_13044);
or U17286 (N_17286,N_13241,N_11248);
and U17287 (N_17287,N_12334,N_12927);
or U17288 (N_17288,N_12719,N_14097);
nor U17289 (N_17289,N_13776,N_11648);
or U17290 (N_17290,N_12330,N_12659);
nand U17291 (N_17291,N_14729,N_10308);
or U17292 (N_17292,N_10207,N_13433);
or U17293 (N_17293,N_11804,N_10074);
and U17294 (N_17294,N_11251,N_14236);
or U17295 (N_17295,N_10635,N_11649);
and U17296 (N_17296,N_10541,N_13660);
nand U17297 (N_17297,N_11504,N_14747);
nand U17298 (N_17298,N_10340,N_12441);
nand U17299 (N_17299,N_13066,N_12128);
or U17300 (N_17300,N_12223,N_11264);
and U17301 (N_17301,N_12220,N_10581);
nor U17302 (N_17302,N_11624,N_11496);
nor U17303 (N_17303,N_12774,N_11578);
nand U17304 (N_17304,N_11706,N_14275);
and U17305 (N_17305,N_12072,N_10344);
xnor U17306 (N_17306,N_11257,N_12611);
or U17307 (N_17307,N_14107,N_11974);
and U17308 (N_17308,N_11602,N_14093);
nand U17309 (N_17309,N_12037,N_11513);
or U17310 (N_17310,N_13899,N_12042);
nor U17311 (N_17311,N_12225,N_11687);
nor U17312 (N_17312,N_14175,N_13002);
xor U17313 (N_17313,N_13384,N_10097);
nor U17314 (N_17314,N_14645,N_11491);
nand U17315 (N_17315,N_11395,N_12816);
or U17316 (N_17316,N_13357,N_11731);
and U17317 (N_17317,N_11928,N_12998);
or U17318 (N_17318,N_13290,N_12121);
nand U17319 (N_17319,N_13870,N_14864);
xnor U17320 (N_17320,N_12024,N_12541);
nor U17321 (N_17321,N_14919,N_12212);
and U17322 (N_17322,N_10774,N_12924);
and U17323 (N_17323,N_13071,N_10472);
nor U17324 (N_17324,N_14804,N_11301);
xor U17325 (N_17325,N_10030,N_12070);
or U17326 (N_17326,N_14117,N_11367);
xor U17327 (N_17327,N_14135,N_11484);
nor U17328 (N_17328,N_14779,N_10271);
xor U17329 (N_17329,N_12351,N_10242);
nand U17330 (N_17330,N_10549,N_14020);
nand U17331 (N_17331,N_11216,N_10781);
nand U17332 (N_17332,N_11227,N_14709);
nor U17333 (N_17333,N_11222,N_13337);
nand U17334 (N_17334,N_10179,N_11985);
nand U17335 (N_17335,N_12929,N_10274);
xnor U17336 (N_17336,N_10165,N_11246);
and U17337 (N_17337,N_10288,N_12586);
nor U17338 (N_17338,N_12539,N_13999);
xor U17339 (N_17339,N_13199,N_13797);
nand U17340 (N_17340,N_11508,N_13553);
or U17341 (N_17341,N_14168,N_13303);
nor U17342 (N_17342,N_13273,N_11355);
and U17343 (N_17343,N_13577,N_10629);
nand U17344 (N_17344,N_13476,N_14612);
nor U17345 (N_17345,N_11849,N_13197);
xnor U17346 (N_17346,N_12316,N_14600);
or U17347 (N_17347,N_10932,N_12308);
nor U17348 (N_17348,N_10152,N_14139);
nor U17349 (N_17349,N_13052,N_14594);
nor U17350 (N_17350,N_10172,N_13856);
or U17351 (N_17351,N_11095,N_10994);
xor U17352 (N_17352,N_14270,N_10857);
or U17353 (N_17353,N_10908,N_14767);
nand U17354 (N_17354,N_12099,N_14361);
nand U17355 (N_17355,N_13686,N_12265);
nand U17356 (N_17356,N_12775,N_14426);
or U17357 (N_17357,N_13990,N_11717);
or U17358 (N_17358,N_13345,N_14137);
or U17359 (N_17359,N_10586,N_11100);
nor U17360 (N_17360,N_12159,N_13393);
nor U17361 (N_17361,N_11391,N_11351);
or U17362 (N_17362,N_10345,N_14351);
and U17363 (N_17363,N_14969,N_14505);
nor U17364 (N_17364,N_12180,N_13891);
nand U17365 (N_17365,N_14773,N_13428);
and U17366 (N_17366,N_11503,N_11966);
or U17367 (N_17367,N_14122,N_11775);
nor U17368 (N_17368,N_11039,N_13640);
or U17369 (N_17369,N_11615,N_13594);
nand U17370 (N_17370,N_13635,N_10527);
nand U17371 (N_17371,N_14927,N_12801);
nand U17372 (N_17372,N_11156,N_12874);
or U17373 (N_17373,N_13929,N_12140);
nor U17374 (N_17374,N_10747,N_10835);
and U17375 (N_17375,N_10187,N_11196);
and U17376 (N_17376,N_11148,N_12152);
nor U17377 (N_17377,N_10036,N_12518);
nand U17378 (N_17378,N_14850,N_12348);
nor U17379 (N_17379,N_10121,N_12562);
xnor U17380 (N_17380,N_12688,N_14222);
xor U17381 (N_17381,N_12183,N_13790);
nand U17382 (N_17382,N_13846,N_13611);
or U17383 (N_17383,N_11949,N_10750);
nand U17384 (N_17384,N_12790,N_14394);
and U17385 (N_17385,N_13211,N_12023);
or U17386 (N_17386,N_12640,N_14880);
nand U17387 (N_17387,N_10810,N_12862);
and U17388 (N_17388,N_10167,N_13045);
and U17389 (N_17389,N_12247,N_13698);
nand U17390 (N_17390,N_13613,N_14006);
nor U17391 (N_17391,N_10047,N_13055);
xnor U17392 (N_17392,N_14741,N_13107);
or U17393 (N_17393,N_13874,N_12038);
nor U17394 (N_17394,N_10631,N_13909);
xor U17395 (N_17395,N_10339,N_10077);
xor U17396 (N_17396,N_11303,N_10129);
nand U17397 (N_17397,N_13285,N_10504);
and U17398 (N_17398,N_13399,N_13658);
or U17399 (N_17399,N_13030,N_14903);
or U17400 (N_17400,N_13655,N_12200);
nand U17401 (N_17401,N_11175,N_13840);
nand U17402 (N_17402,N_11690,N_12642);
and U17403 (N_17403,N_10174,N_10471);
xor U17404 (N_17404,N_13300,N_14198);
nor U17405 (N_17405,N_11083,N_10890);
nand U17406 (N_17406,N_11571,N_14306);
xnor U17407 (N_17407,N_11576,N_12377);
and U17408 (N_17408,N_13130,N_11589);
xnor U17409 (N_17409,N_14017,N_14431);
and U17410 (N_17410,N_12776,N_14980);
and U17411 (N_17411,N_11817,N_14060);
or U17412 (N_17412,N_14665,N_10145);
xnor U17413 (N_17413,N_14999,N_14427);
xnor U17414 (N_17414,N_12311,N_11305);
xor U17415 (N_17415,N_10392,N_12608);
or U17416 (N_17416,N_13844,N_14640);
or U17417 (N_17417,N_12537,N_11721);
or U17418 (N_17418,N_14458,N_13019);
and U17419 (N_17419,N_13340,N_14676);
and U17420 (N_17420,N_13051,N_13456);
xnor U17421 (N_17421,N_14052,N_14707);
and U17422 (N_17422,N_13255,N_13768);
and U17423 (N_17423,N_11064,N_11025);
or U17424 (N_17424,N_10698,N_14309);
nor U17425 (N_17425,N_13981,N_10796);
or U17426 (N_17426,N_10468,N_10836);
or U17427 (N_17427,N_12317,N_12339);
and U17428 (N_17428,N_14916,N_10016);
and U17429 (N_17429,N_13595,N_14890);
or U17430 (N_17430,N_12479,N_14739);
xnor U17431 (N_17431,N_10539,N_13172);
nor U17432 (N_17432,N_14272,N_13148);
nand U17433 (N_17433,N_12989,N_13082);
nand U17434 (N_17434,N_12315,N_14598);
or U17435 (N_17435,N_11791,N_14772);
nand U17436 (N_17436,N_12437,N_13240);
and U17437 (N_17437,N_12270,N_14539);
xnor U17438 (N_17438,N_11662,N_10754);
xor U17439 (N_17439,N_13497,N_10182);
and U17440 (N_17440,N_14473,N_14467);
or U17441 (N_17441,N_12495,N_10178);
nor U17442 (N_17442,N_14090,N_14191);
nand U17443 (N_17443,N_13414,N_10460);
xnor U17444 (N_17444,N_11178,N_10484);
nor U17445 (N_17445,N_10105,N_14245);
nor U17446 (N_17446,N_14335,N_14743);
or U17447 (N_17447,N_11665,N_10770);
nor U17448 (N_17448,N_10406,N_14885);
nor U17449 (N_17449,N_11558,N_11213);
nand U17450 (N_17450,N_11701,N_12795);
and U17451 (N_17451,N_10858,N_12750);
nor U17452 (N_17452,N_14019,N_13961);
and U17453 (N_17453,N_10900,N_12191);
nand U17454 (N_17454,N_12636,N_10151);
and U17455 (N_17455,N_11258,N_11937);
and U17456 (N_17456,N_12926,N_14609);
nor U17457 (N_17457,N_12861,N_13893);
and U17458 (N_17458,N_13363,N_14462);
nand U17459 (N_17459,N_14667,N_14315);
and U17460 (N_17460,N_12243,N_13890);
nand U17461 (N_17461,N_12199,N_10788);
xnor U17462 (N_17462,N_13866,N_14411);
nand U17463 (N_17463,N_14686,N_13296);
or U17464 (N_17464,N_12498,N_10113);
xnor U17465 (N_17465,N_10160,N_10523);
nand U17466 (N_17466,N_13232,N_10710);
xnor U17467 (N_17467,N_11197,N_13675);
nand U17468 (N_17468,N_12819,N_13552);
and U17469 (N_17469,N_10958,N_12004);
and U17470 (N_17470,N_11709,N_13871);
and U17471 (N_17471,N_12516,N_13770);
nor U17472 (N_17472,N_11820,N_13496);
or U17473 (N_17473,N_14404,N_10989);
and U17474 (N_17474,N_13687,N_11208);
nor U17475 (N_17475,N_14363,N_13369);
nand U17476 (N_17476,N_10103,N_14993);
nor U17477 (N_17477,N_10884,N_11510);
nor U17478 (N_17478,N_11824,N_12202);
nor U17479 (N_17479,N_11577,N_13489);
nor U17480 (N_17480,N_11616,N_13907);
or U17481 (N_17481,N_11492,N_14997);
and U17482 (N_17482,N_11405,N_10704);
nor U17483 (N_17483,N_11565,N_14797);
nor U17484 (N_17484,N_14896,N_10548);
nand U17485 (N_17485,N_13053,N_12898);
and U17486 (N_17486,N_10088,N_13056);
or U17487 (N_17487,N_10552,N_13344);
and U17488 (N_17488,N_13014,N_12952);
xnor U17489 (N_17489,N_11912,N_13905);
or U17490 (N_17490,N_12446,N_11574);
and U17491 (N_17491,N_13884,N_10665);
nand U17492 (N_17492,N_12555,N_14200);
or U17493 (N_17493,N_13121,N_10037);
and U17494 (N_17494,N_13724,N_11797);
nand U17495 (N_17495,N_14170,N_12550);
and U17496 (N_17496,N_13709,N_13564);
nor U17497 (N_17497,N_11184,N_14559);
nand U17498 (N_17498,N_14660,N_10627);
or U17499 (N_17499,N_14650,N_11029);
xnor U17500 (N_17500,N_13138,N_11820);
nor U17501 (N_17501,N_14708,N_13430);
nand U17502 (N_17502,N_12393,N_11843);
and U17503 (N_17503,N_14605,N_13563);
nand U17504 (N_17504,N_14582,N_13817);
or U17505 (N_17505,N_13035,N_14934);
and U17506 (N_17506,N_13741,N_12465);
xor U17507 (N_17507,N_10106,N_11435);
and U17508 (N_17508,N_12163,N_13272);
nor U17509 (N_17509,N_10741,N_13404);
and U17510 (N_17510,N_11128,N_14754);
or U17511 (N_17511,N_14415,N_14259);
xnor U17512 (N_17512,N_13076,N_13100);
or U17513 (N_17513,N_14824,N_12265);
or U17514 (N_17514,N_14776,N_11518);
nand U17515 (N_17515,N_12699,N_12031);
and U17516 (N_17516,N_10719,N_11689);
nor U17517 (N_17517,N_14860,N_11348);
and U17518 (N_17518,N_10264,N_13591);
nand U17519 (N_17519,N_10520,N_11584);
xnor U17520 (N_17520,N_10777,N_14327);
and U17521 (N_17521,N_13231,N_12807);
xor U17522 (N_17522,N_14544,N_10862);
and U17523 (N_17523,N_12828,N_13807);
and U17524 (N_17524,N_12718,N_14918);
and U17525 (N_17525,N_13911,N_11548);
xor U17526 (N_17526,N_14331,N_10872);
or U17527 (N_17527,N_14321,N_10940);
xnor U17528 (N_17528,N_10483,N_11410);
xor U17529 (N_17529,N_12430,N_10011);
and U17530 (N_17530,N_12645,N_12668);
and U17531 (N_17531,N_13544,N_11926);
nor U17532 (N_17532,N_10964,N_14029);
nor U17533 (N_17533,N_13775,N_13002);
nand U17534 (N_17534,N_12850,N_11177);
nand U17535 (N_17535,N_10811,N_12172);
or U17536 (N_17536,N_13654,N_12428);
nand U17537 (N_17537,N_11250,N_13265);
nor U17538 (N_17538,N_12676,N_10495);
xor U17539 (N_17539,N_10814,N_11822);
or U17540 (N_17540,N_12325,N_14750);
or U17541 (N_17541,N_12380,N_10324);
xor U17542 (N_17542,N_12373,N_11806);
and U17543 (N_17543,N_11075,N_12429);
and U17544 (N_17544,N_10127,N_14884);
or U17545 (N_17545,N_13629,N_14990);
or U17546 (N_17546,N_10816,N_12668);
nand U17547 (N_17547,N_10109,N_14248);
nand U17548 (N_17548,N_10382,N_11842);
nand U17549 (N_17549,N_11500,N_11849);
nor U17550 (N_17550,N_12728,N_11076);
xnor U17551 (N_17551,N_12936,N_10693);
nor U17552 (N_17552,N_11362,N_10640);
nand U17553 (N_17553,N_10303,N_13087);
nand U17554 (N_17554,N_11650,N_14632);
xnor U17555 (N_17555,N_11377,N_11394);
nand U17556 (N_17556,N_13550,N_11274);
nand U17557 (N_17557,N_14450,N_14828);
and U17558 (N_17558,N_13966,N_11856);
xor U17559 (N_17559,N_14038,N_13787);
or U17560 (N_17560,N_10084,N_12625);
nor U17561 (N_17561,N_14436,N_14882);
nand U17562 (N_17562,N_12253,N_14875);
or U17563 (N_17563,N_13633,N_12242);
nand U17564 (N_17564,N_10152,N_14195);
nor U17565 (N_17565,N_12307,N_11368);
nor U17566 (N_17566,N_11134,N_11308);
nor U17567 (N_17567,N_12284,N_13557);
nand U17568 (N_17568,N_13747,N_11088);
nor U17569 (N_17569,N_10740,N_11377);
xnor U17570 (N_17570,N_11986,N_13015);
or U17571 (N_17571,N_12485,N_12662);
xnor U17572 (N_17572,N_13987,N_14235);
nand U17573 (N_17573,N_11949,N_11299);
and U17574 (N_17574,N_12006,N_10561);
nand U17575 (N_17575,N_13985,N_13670);
nand U17576 (N_17576,N_12457,N_11295);
xnor U17577 (N_17577,N_13236,N_12909);
nor U17578 (N_17578,N_11690,N_10820);
xnor U17579 (N_17579,N_11537,N_13942);
nor U17580 (N_17580,N_13878,N_13781);
or U17581 (N_17581,N_14096,N_11817);
nand U17582 (N_17582,N_10321,N_14434);
nor U17583 (N_17583,N_12500,N_13461);
nor U17584 (N_17584,N_14056,N_14498);
and U17585 (N_17585,N_13760,N_13645);
and U17586 (N_17586,N_12794,N_10412);
or U17587 (N_17587,N_11201,N_10937);
and U17588 (N_17588,N_11432,N_10195);
nor U17589 (N_17589,N_13915,N_12680);
or U17590 (N_17590,N_13125,N_12288);
or U17591 (N_17591,N_13463,N_14865);
xor U17592 (N_17592,N_10024,N_14433);
nand U17593 (N_17593,N_12831,N_10234);
and U17594 (N_17594,N_13705,N_12399);
nor U17595 (N_17595,N_14898,N_10663);
nor U17596 (N_17596,N_10618,N_13936);
xnor U17597 (N_17597,N_12603,N_12318);
nor U17598 (N_17598,N_10323,N_10333);
xnor U17599 (N_17599,N_10414,N_13767);
xnor U17600 (N_17600,N_13171,N_12638);
and U17601 (N_17601,N_14961,N_14740);
and U17602 (N_17602,N_14337,N_14848);
xor U17603 (N_17603,N_14371,N_11035);
or U17604 (N_17604,N_14662,N_14803);
xnor U17605 (N_17605,N_12276,N_10128);
or U17606 (N_17606,N_12001,N_12235);
nand U17607 (N_17607,N_12385,N_12193);
and U17608 (N_17608,N_12018,N_14690);
or U17609 (N_17609,N_11913,N_12448);
xor U17610 (N_17610,N_12945,N_10413);
nor U17611 (N_17611,N_10693,N_10397);
nor U17612 (N_17612,N_10930,N_12720);
nor U17613 (N_17613,N_13688,N_11955);
and U17614 (N_17614,N_12775,N_14280);
and U17615 (N_17615,N_10083,N_13220);
or U17616 (N_17616,N_13190,N_10188);
or U17617 (N_17617,N_13605,N_10048);
nand U17618 (N_17618,N_10523,N_13368);
nor U17619 (N_17619,N_12539,N_10707);
and U17620 (N_17620,N_11130,N_14489);
nor U17621 (N_17621,N_14270,N_11184);
nor U17622 (N_17622,N_12266,N_14041);
xnor U17623 (N_17623,N_10285,N_13060);
xnor U17624 (N_17624,N_14876,N_11951);
xnor U17625 (N_17625,N_11558,N_11548);
xor U17626 (N_17626,N_12576,N_11818);
or U17627 (N_17627,N_11409,N_14407);
nor U17628 (N_17628,N_12424,N_13431);
nor U17629 (N_17629,N_12361,N_12493);
and U17630 (N_17630,N_10927,N_14076);
xor U17631 (N_17631,N_11804,N_12588);
or U17632 (N_17632,N_11497,N_12324);
xor U17633 (N_17633,N_10056,N_12261);
nor U17634 (N_17634,N_11905,N_14351);
or U17635 (N_17635,N_12910,N_14697);
xor U17636 (N_17636,N_11405,N_14051);
and U17637 (N_17637,N_10559,N_12402);
and U17638 (N_17638,N_13830,N_11496);
nor U17639 (N_17639,N_13857,N_12436);
nor U17640 (N_17640,N_11719,N_13220);
and U17641 (N_17641,N_10053,N_11704);
or U17642 (N_17642,N_11503,N_11018);
nor U17643 (N_17643,N_11104,N_10901);
and U17644 (N_17644,N_10102,N_14193);
nor U17645 (N_17645,N_12580,N_10619);
and U17646 (N_17646,N_12058,N_12215);
xnor U17647 (N_17647,N_13300,N_12575);
nor U17648 (N_17648,N_13365,N_14339);
and U17649 (N_17649,N_10487,N_12219);
xor U17650 (N_17650,N_13563,N_12849);
or U17651 (N_17651,N_14998,N_10476);
xor U17652 (N_17652,N_11802,N_14920);
or U17653 (N_17653,N_14218,N_11916);
nor U17654 (N_17654,N_10696,N_11001);
or U17655 (N_17655,N_11076,N_14974);
nor U17656 (N_17656,N_13377,N_14556);
or U17657 (N_17657,N_14972,N_12022);
or U17658 (N_17658,N_11540,N_11770);
or U17659 (N_17659,N_14740,N_14028);
and U17660 (N_17660,N_10272,N_11704);
and U17661 (N_17661,N_12185,N_10397);
nand U17662 (N_17662,N_13189,N_13845);
nor U17663 (N_17663,N_11580,N_14850);
nand U17664 (N_17664,N_12982,N_10387);
and U17665 (N_17665,N_14153,N_13983);
xnor U17666 (N_17666,N_11485,N_13613);
or U17667 (N_17667,N_13048,N_13556);
and U17668 (N_17668,N_12773,N_13397);
or U17669 (N_17669,N_11218,N_12623);
or U17670 (N_17670,N_14553,N_11244);
xnor U17671 (N_17671,N_13067,N_13353);
nand U17672 (N_17672,N_14218,N_11053);
nand U17673 (N_17673,N_14821,N_12152);
and U17674 (N_17674,N_11316,N_13163);
nand U17675 (N_17675,N_10250,N_12362);
nor U17676 (N_17676,N_13217,N_10313);
or U17677 (N_17677,N_11453,N_11586);
xnor U17678 (N_17678,N_11524,N_11354);
or U17679 (N_17679,N_11879,N_11062);
nand U17680 (N_17680,N_13396,N_12117);
and U17681 (N_17681,N_11667,N_11101);
xor U17682 (N_17682,N_10961,N_13991);
nand U17683 (N_17683,N_11614,N_10695);
nor U17684 (N_17684,N_13249,N_13138);
nor U17685 (N_17685,N_11455,N_14316);
or U17686 (N_17686,N_12688,N_10620);
and U17687 (N_17687,N_11702,N_11860);
xor U17688 (N_17688,N_13637,N_11738);
and U17689 (N_17689,N_10464,N_12628);
nand U17690 (N_17690,N_12365,N_12148);
nor U17691 (N_17691,N_13077,N_14985);
and U17692 (N_17692,N_11192,N_10353);
and U17693 (N_17693,N_10188,N_13032);
nor U17694 (N_17694,N_10699,N_11536);
or U17695 (N_17695,N_14343,N_13152);
nand U17696 (N_17696,N_11359,N_11353);
and U17697 (N_17697,N_12290,N_10407);
or U17698 (N_17698,N_12738,N_14898);
or U17699 (N_17699,N_12109,N_14841);
nor U17700 (N_17700,N_12542,N_11891);
nand U17701 (N_17701,N_12616,N_10586);
and U17702 (N_17702,N_12808,N_12212);
nand U17703 (N_17703,N_11553,N_11225);
and U17704 (N_17704,N_11276,N_11197);
nand U17705 (N_17705,N_12484,N_11566);
nor U17706 (N_17706,N_11931,N_14830);
and U17707 (N_17707,N_14632,N_13533);
or U17708 (N_17708,N_13121,N_14086);
nand U17709 (N_17709,N_13844,N_14637);
and U17710 (N_17710,N_14487,N_14420);
xnor U17711 (N_17711,N_14185,N_13640);
xor U17712 (N_17712,N_11274,N_10245);
nand U17713 (N_17713,N_12668,N_11521);
nand U17714 (N_17714,N_12247,N_13730);
nor U17715 (N_17715,N_12344,N_10136);
or U17716 (N_17716,N_13010,N_12504);
nand U17717 (N_17717,N_11161,N_12279);
or U17718 (N_17718,N_14852,N_11900);
nor U17719 (N_17719,N_10202,N_10684);
xnor U17720 (N_17720,N_13410,N_11690);
and U17721 (N_17721,N_11231,N_11623);
xnor U17722 (N_17722,N_14434,N_12091);
and U17723 (N_17723,N_10356,N_12631);
or U17724 (N_17724,N_10184,N_13766);
or U17725 (N_17725,N_14824,N_11515);
or U17726 (N_17726,N_11591,N_14166);
and U17727 (N_17727,N_14803,N_13225);
nand U17728 (N_17728,N_14301,N_13917);
or U17729 (N_17729,N_12746,N_13731);
and U17730 (N_17730,N_12643,N_10521);
nor U17731 (N_17731,N_10856,N_11862);
and U17732 (N_17732,N_13431,N_11197);
or U17733 (N_17733,N_12334,N_12765);
xor U17734 (N_17734,N_11582,N_14334);
nor U17735 (N_17735,N_14265,N_14632);
and U17736 (N_17736,N_10005,N_13835);
xor U17737 (N_17737,N_11866,N_13309);
xnor U17738 (N_17738,N_10850,N_12575);
nor U17739 (N_17739,N_12384,N_10389);
xnor U17740 (N_17740,N_13138,N_12962);
xor U17741 (N_17741,N_14735,N_12681);
nand U17742 (N_17742,N_13641,N_12932);
nand U17743 (N_17743,N_10263,N_10183);
and U17744 (N_17744,N_14789,N_10118);
and U17745 (N_17745,N_11014,N_11166);
and U17746 (N_17746,N_11817,N_14205);
or U17747 (N_17747,N_11853,N_14067);
nor U17748 (N_17748,N_10995,N_10811);
and U17749 (N_17749,N_13820,N_10092);
nand U17750 (N_17750,N_10647,N_14597);
xnor U17751 (N_17751,N_14176,N_11963);
and U17752 (N_17752,N_14583,N_11263);
and U17753 (N_17753,N_11546,N_12544);
nor U17754 (N_17754,N_11433,N_10903);
or U17755 (N_17755,N_10080,N_10715);
nand U17756 (N_17756,N_14448,N_12065);
xor U17757 (N_17757,N_14133,N_14796);
or U17758 (N_17758,N_14525,N_10640);
xnor U17759 (N_17759,N_13211,N_10235);
nand U17760 (N_17760,N_12765,N_14133);
nand U17761 (N_17761,N_14111,N_11849);
and U17762 (N_17762,N_10059,N_11141);
nor U17763 (N_17763,N_11451,N_13804);
and U17764 (N_17764,N_12730,N_13279);
nor U17765 (N_17765,N_14896,N_11185);
nand U17766 (N_17766,N_12545,N_10172);
nand U17767 (N_17767,N_13419,N_12409);
nor U17768 (N_17768,N_14146,N_14967);
and U17769 (N_17769,N_10472,N_13708);
or U17770 (N_17770,N_10328,N_11928);
xor U17771 (N_17771,N_12490,N_13565);
nor U17772 (N_17772,N_13231,N_11682);
or U17773 (N_17773,N_14240,N_14756);
nand U17774 (N_17774,N_13687,N_11124);
nand U17775 (N_17775,N_12808,N_13115);
nor U17776 (N_17776,N_14322,N_12361);
nor U17777 (N_17777,N_10471,N_10173);
or U17778 (N_17778,N_13768,N_11588);
or U17779 (N_17779,N_12520,N_14173);
nor U17780 (N_17780,N_11070,N_11356);
xnor U17781 (N_17781,N_13340,N_10939);
xor U17782 (N_17782,N_11155,N_11636);
nand U17783 (N_17783,N_14173,N_14835);
nor U17784 (N_17784,N_10538,N_11081);
and U17785 (N_17785,N_12517,N_12281);
nand U17786 (N_17786,N_12467,N_11532);
or U17787 (N_17787,N_13609,N_10618);
nor U17788 (N_17788,N_10923,N_14991);
xor U17789 (N_17789,N_11494,N_14699);
nor U17790 (N_17790,N_11304,N_13151);
xnor U17791 (N_17791,N_13990,N_12220);
nand U17792 (N_17792,N_12739,N_14247);
and U17793 (N_17793,N_12471,N_10614);
nand U17794 (N_17794,N_14629,N_10311);
xor U17795 (N_17795,N_11072,N_13797);
xnor U17796 (N_17796,N_12267,N_10460);
nor U17797 (N_17797,N_14796,N_13178);
nand U17798 (N_17798,N_13843,N_14099);
xnor U17799 (N_17799,N_11829,N_13385);
or U17800 (N_17800,N_14127,N_10941);
nor U17801 (N_17801,N_12239,N_13459);
or U17802 (N_17802,N_14636,N_12019);
nor U17803 (N_17803,N_13619,N_14531);
or U17804 (N_17804,N_11880,N_13641);
nor U17805 (N_17805,N_10114,N_14593);
or U17806 (N_17806,N_12253,N_10761);
xnor U17807 (N_17807,N_13888,N_10608);
nand U17808 (N_17808,N_11529,N_14341);
nor U17809 (N_17809,N_10442,N_13175);
and U17810 (N_17810,N_11084,N_14489);
nor U17811 (N_17811,N_14052,N_13150);
nor U17812 (N_17812,N_13741,N_10452);
xnor U17813 (N_17813,N_12215,N_12121);
nand U17814 (N_17814,N_13170,N_11705);
and U17815 (N_17815,N_14227,N_11513);
nand U17816 (N_17816,N_12883,N_10539);
nand U17817 (N_17817,N_10397,N_14867);
xor U17818 (N_17818,N_13152,N_13625);
nand U17819 (N_17819,N_13638,N_14078);
and U17820 (N_17820,N_11781,N_12057);
nor U17821 (N_17821,N_10680,N_11292);
xor U17822 (N_17822,N_13765,N_10020);
nand U17823 (N_17823,N_11199,N_12445);
and U17824 (N_17824,N_13406,N_14919);
xnor U17825 (N_17825,N_14259,N_10972);
and U17826 (N_17826,N_12434,N_14861);
nor U17827 (N_17827,N_10538,N_14749);
nand U17828 (N_17828,N_10649,N_11301);
nor U17829 (N_17829,N_13236,N_10378);
xor U17830 (N_17830,N_12270,N_10125);
and U17831 (N_17831,N_13977,N_11606);
or U17832 (N_17832,N_11330,N_10035);
and U17833 (N_17833,N_14034,N_11718);
xor U17834 (N_17834,N_10415,N_10095);
or U17835 (N_17835,N_12500,N_12707);
nor U17836 (N_17836,N_10956,N_13473);
or U17837 (N_17837,N_13972,N_10158);
or U17838 (N_17838,N_13126,N_12789);
nor U17839 (N_17839,N_10613,N_10784);
nand U17840 (N_17840,N_10864,N_13392);
and U17841 (N_17841,N_14759,N_13315);
xnor U17842 (N_17842,N_11604,N_14215);
nand U17843 (N_17843,N_13195,N_13562);
and U17844 (N_17844,N_13516,N_13230);
nor U17845 (N_17845,N_12193,N_10050);
and U17846 (N_17846,N_14159,N_13594);
or U17847 (N_17847,N_12661,N_11005);
xor U17848 (N_17848,N_14078,N_14956);
nor U17849 (N_17849,N_12761,N_11704);
nand U17850 (N_17850,N_12380,N_12322);
or U17851 (N_17851,N_14214,N_11274);
xor U17852 (N_17852,N_10223,N_14668);
and U17853 (N_17853,N_12962,N_11675);
nor U17854 (N_17854,N_13447,N_10590);
nor U17855 (N_17855,N_10802,N_14336);
xor U17856 (N_17856,N_13636,N_14326);
and U17857 (N_17857,N_14633,N_14535);
nor U17858 (N_17858,N_13439,N_13004);
nor U17859 (N_17859,N_12525,N_14338);
xor U17860 (N_17860,N_11179,N_10883);
and U17861 (N_17861,N_13894,N_12613);
xor U17862 (N_17862,N_10207,N_14969);
nand U17863 (N_17863,N_14212,N_14310);
nor U17864 (N_17864,N_11419,N_10683);
nor U17865 (N_17865,N_14075,N_10236);
or U17866 (N_17866,N_13114,N_14028);
or U17867 (N_17867,N_11687,N_10536);
and U17868 (N_17868,N_13682,N_10995);
xnor U17869 (N_17869,N_14067,N_10174);
and U17870 (N_17870,N_11986,N_10619);
nor U17871 (N_17871,N_14973,N_13916);
or U17872 (N_17872,N_13185,N_10220);
and U17873 (N_17873,N_11055,N_11767);
or U17874 (N_17874,N_14391,N_10939);
and U17875 (N_17875,N_10555,N_13670);
and U17876 (N_17876,N_10546,N_12726);
and U17877 (N_17877,N_11471,N_12923);
xnor U17878 (N_17878,N_10253,N_11285);
nand U17879 (N_17879,N_10611,N_14005);
nor U17880 (N_17880,N_13323,N_13944);
or U17881 (N_17881,N_12462,N_11695);
xor U17882 (N_17882,N_13109,N_14444);
xor U17883 (N_17883,N_14026,N_13292);
nor U17884 (N_17884,N_12069,N_11318);
nor U17885 (N_17885,N_10358,N_13361);
and U17886 (N_17886,N_11142,N_13186);
and U17887 (N_17887,N_11927,N_10490);
nor U17888 (N_17888,N_11622,N_13968);
nand U17889 (N_17889,N_11947,N_10386);
nor U17890 (N_17890,N_12254,N_10072);
xnor U17891 (N_17891,N_11198,N_10934);
nor U17892 (N_17892,N_11821,N_12609);
nand U17893 (N_17893,N_13926,N_10492);
and U17894 (N_17894,N_14629,N_12855);
nand U17895 (N_17895,N_10183,N_11688);
and U17896 (N_17896,N_10333,N_13156);
nand U17897 (N_17897,N_13344,N_12371);
nor U17898 (N_17898,N_11698,N_13963);
nor U17899 (N_17899,N_10617,N_14240);
nand U17900 (N_17900,N_12125,N_10975);
nand U17901 (N_17901,N_14149,N_13545);
nand U17902 (N_17902,N_14751,N_14628);
nor U17903 (N_17903,N_10168,N_10010);
or U17904 (N_17904,N_13372,N_11270);
nand U17905 (N_17905,N_14157,N_13810);
xnor U17906 (N_17906,N_13768,N_14955);
or U17907 (N_17907,N_12013,N_13724);
and U17908 (N_17908,N_12111,N_10452);
nor U17909 (N_17909,N_11567,N_10367);
nor U17910 (N_17910,N_11252,N_10708);
or U17911 (N_17911,N_14265,N_14365);
nor U17912 (N_17912,N_13923,N_10885);
and U17913 (N_17913,N_11976,N_12371);
and U17914 (N_17914,N_10534,N_14962);
or U17915 (N_17915,N_12979,N_10174);
and U17916 (N_17916,N_14803,N_11581);
and U17917 (N_17917,N_10048,N_12906);
nor U17918 (N_17918,N_10076,N_13169);
nand U17919 (N_17919,N_12232,N_10491);
and U17920 (N_17920,N_14876,N_12135);
nand U17921 (N_17921,N_12144,N_10606);
or U17922 (N_17922,N_12171,N_11833);
or U17923 (N_17923,N_10968,N_10874);
nand U17924 (N_17924,N_10468,N_13788);
nand U17925 (N_17925,N_12940,N_13347);
nor U17926 (N_17926,N_10863,N_13276);
xnor U17927 (N_17927,N_14414,N_10575);
xor U17928 (N_17928,N_11203,N_13408);
or U17929 (N_17929,N_13942,N_13961);
xnor U17930 (N_17930,N_13808,N_14612);
and U17931 (N_17931,N_13726,N_11312);
nand U17932 (N_17932,N_10245,N_13847);
nand U17933 (N_17933,N_14855,N_13810);
nor U17934 (N_17934,N_11001,N_14491);
nand U17935 (N_17935,N_12388,N_10493);
and U17936 (N_17936,N_12311,N_14006);
nor U17937 (N_17937,N_11524,N_13812);
nor U17938 (N_17938,N_14929,N_14913);
and U17939 (N_17939,N_10722,N_12197);
or U17940 (N_17940,N_11867,N_14363);
nand U17941 (N_17941,N_13756,N_13991);
and U17942 (N_17942,N_11905,N_14495);
xnor U17943 (N_17943,N_11928,N_14323);
or U17944 (N_17944,N_12861,N_14508);
and U17945 (N_17945,N_14151,N_11377);
nor U17946 (N_17946,N_14361,N_11252);
nor U17947 (N_17947,N_12317,N_10487);
nor U17948 (N_17948,N_11563,N_10908);
and U17949 (N_17949,N_13596,N_10810);
nand U17950 (N_17950,N_14849,N_12001);
nor U17951 (N_17951,N_11007,N_13420);
nor U17952 (N_17952,N_12805,N_10930);
nand U17953 (N_17953,N_13547,N_10954);
or U17954 (N_17954,N_11343,N_11541);
or U17955 (N_17955,N_11911,N_12339);
nand U17956 (N_17956,N_11069,N_12741);
nand U17957 (N_17957,N_14916,N_11228);
nor U17958 (N_17958,N_13470,N_12480);
nand U17959 (N_17959,N_14573,N_14677);
or U17960 (N_17960,N_11533,N_14411);
or U17961 (N_17961,N_14121,N_11895);
xnor U17962 (N_17962,N_10380,N_14429);
and U17963 (N_17963,N_13074,N_11571);
xnor U17964 (N_17964,N_14038,N_10152);
nor U17965 (N_17965,N_10104,N_13244);
nand U17966 (N_17966,N_11262,N_12388);
and U17967 (N_17967,N_10138,N_12656);
xnor U17968 (N_17968,N_13127,N_10981);
and U17969 (N_17969,N_13736,N_14381);
and U17970 (N_17970,N_14455,N_11920);
nand U17971 (N_17971,N_12096,N_10134);
nand U17972 (N_17972,N_12933,N_10368);
nand U17973 (N_17973,N_11679,N_11071);
and U17974 (N_17974,N_10744,N_12966);
xor U17975 (N_17975,N_10074,N_12961);
and U17976 (N_17976,N_12138,N_12559);
or U17977 (N_17977,N_10445,N_12921);
nor U17978 (N_17978,N_11153,N_13683);
nand U17979 (N_17979,N_10112,N_12630);
nand U17980 (N_17980,N_13646,N_13928);
nor U17981 (N_17981,N_10936,N_11774);
nor U17982 (N_17982,N_10623,N_14335);
xnor U17983 (N_17983,N_12671,N_12119);
nand U17984 (N_17984,N_12466,N_12738);
nor U17985 (N_17985,N_13584,N_11640);
xnor U17986 (N_17986,N_13137,N_12952);
nor U17987 (N_17987,N_13260,N_12905);
or U17988 (N_17988,N_10603,N_14523);
and U17989 (N_17989,N_10760,N_10130);
xor U17990 (N_17990,N_14082,N_14169);
nor U17991 (N_17991,N_10063,N_11295);
nor U17992 (N_17992,N_12844,N_14237);
nor U17993 (N_17993,N_12664,N_10209);
nand U17994 (N_17994,N_12738,N_12918);
xor U17995 (N_17995,N_11063,N_10423);
or U17996 (N_17996,N_12779,N_12306);
or U17997 (N_17997,N_11014,N_13253);
xnor U17998 (N_17998,N_13493,N_11291);
nor U17999 (N_17999,N_14202,N_11896);
xnor U18000 (N_18000,N_12742,N_11538);
nand U18001 (N_18001,N_12076,N_10368);
or U18002 (N_18002,N_14073,N_13876);
xnor U18003 (N_18003,N_12163,N_10935);
nor U18004 (N_18004,N_13995,N_11960);
xor U18005 (N_18005,N_12932,N_13041);
or U18006 (N_18006,N_10412,N_11608);
nor U18007 (N_18007,N_14621,N_10306);
nand U18008 (N_18008,N_12146,N_14439);
or U18009 (N_18009,N_12744,N_10995);
xnor U18010 (N_18010,N_14055,N_11071);
nor U18011 (N_18011,N_12022,N_13721);
or U18012 (N_18012,N_11387,N_11243);
nor U18013 (N_18013,N_11795,N_13221);
and U18014 (N_18014,N_10003,N_12669);
xnor U18015 (N_18015,N_13977,N_10108);
or U18016 (N_18016,N_13091,N_10656);
nor U18017 (N_18017,N_14245,N_14144);
or U18018 (N_18018,N_14149,N_13272);
nor U18019 (N_18019,N_14940,N_14411);
and U18020 (N_18020,N_12973,N_14132);
nand U18021 (N_18021,N_11328,N_13263);
or U18022 (N_18022,N_13027,N_10033);
xnor U18023 (N_18023,N_10644,N_12826);
nor U18024 (N_18024,N_10149,N_11111);
nor U18025 (N_18025,N_10560,N_11288);
nand U18026 (N_18026,N_13958,N_11956);
or U18027 (N_18027,N_10983,N_14648);
or U18028 (N_18028,N_13104,N_13867);
and U18029 (N_18029,N_11424,N_12957);
xor U18030 (N_18030,N_11220,N_11278);
nor U18031 (N_18031,N_12212,N_11341);
nand U18032 (N_18032,N_11622,N_13255);
or U18033 (N_18033,N_12587,N_14625);
nor U18034 (N_18034,N_11288,N_11314);
or U18035 (N_18035,N_11797,N_13931);
or U18036 (N_18036,N_10241,N_12244);
and U18037 (N_18037,N_12889,N_14130);
nor U18038 (N_18038,N_14806,N_10387);
nand U18039 (N_18039,N_14028,N_10332);
nand U18040 (N_18040,N_14568,N_12642);
xnor U18041 (N_18041,N_11195,N_14962);
or U18042 (N_18042,N_11473,N_13365);
and U18043 (N_18043,N_12428,N_14541);
xor U18044 (N_18044,N_11716,N_13794);
nor U18045 (N_18045,N_12387,N_10729);
xor U18046 (N_18046,N_10385,N_11611);
nor U18047 (N_18047,N_13577,N_14591);
xor U18048 (N_18048,N_10726,N_13795);
xor U18049 (N_18049,N_10054,N_11224);
xnor U18050 (N_18050,N_13701,N_14241);
and U18051 (N_18051,N_11545,N_10774);
and U18052 (N_18052,N_10519,N_14814);
nor U18053 (N_18053,N_11036,N_14430);
xor U18054 (N_18054,N_13299,N_10343);
or U18055 (N_18055,N_13380,N_10268);
or U18056 (N_18056,N_13241,N_11850);
nand U18057 (N_18057,N_11285,N_11307);
nor U18058 (N_18058,N_13512,N_13370);
and U18059 (N_18059,N_13757,N_12342);
or U18060 (N_18060,N_14115,N_10170);
and U18061 (N_18061,N_10081,N_13992);
nand U18062 (N_18062,N_14555,N_12136);
nand U18063 (N_18063,N_13314,N_13976);
and U18064 (N_18064,N_14991,N_13534);
and U18065 (N_18065,N_12847,N_10821);
and U18066 (N_18066,N_11389,N_11736);
xor U18067 (N_18067,N_14190,N_12739);
nand U18068 (N_18068,N_13287,N_10896);
nor U18069 (N_18069,N_14018,N_10398);
or U18070 (N_18070,N_13111,N_14221);
nand U18071 (N_18071,N_11632,N_10324);
xor U18072 (N_18072,N_10379,N_11148);
and U18073 (N_18073,N_13436,N_10675);
nor U18074 (N_18074,N_12339,N_12157);
nand U18075 (N_18075,N_14990,N_12252);
xnor U18076 (N_18076,N_13426,N_14864);
xnor U18077 (N_18077,N_12517,N_14858);
nand U18078 (N_18078,N_12391,N_14249);
nor U18079 (N_18079,N_10666,N_10064);
nand U18080 (N_18080,N_13831,N_14403);
or U18081 (N_18081,N_10125,N_10465);
or U18082 (N_18082,N_11369,N_11063);
and U18083 (N_18083,N_13162,N_10469);
xor U18084 (N_18084,N_11650,N_14559);
or U18085 (N_18085,N_10462,N_12219);
and U18086 (N_18086,N_13496,N_14985);
nand U18087 (N_18087,N_13481,N_11635);
xor U18088 (N_18088,N_10081,N_12076);
xnor U18089 (N_18089,N_10824,N_12202);
nor U18090 (N_18090,N_10042,N_12739);
or U18091 (N_18091,N_12277,N_11303);
and U18092 (N_18092,N_12883,N_10112);
xor U18093 (N_18093,N_14826,N_13011);
and U18094 (N_18094,N_10636,N_10504);
nand U18095 (N_18095,N_11409,N_11077);
or U18096 (N_18096,N_14022,N_10876);
nand U18097 (N_18097,N_12573,N_12409);
nor U18098 (N_18098,N_14279,N_14304);
nand U18099 (N_18099,N_12272,N_10126);
and U18100 (N_18100,N_10695,N_12944);
and U18101 (N_18101,N_10429,N_13091);
nor U18102 (N_18102,N_13886,N_10101);
and U18103 (N_18103,N_13246,N_10199);
and U18104 (N_18104,N_13492,N_12354);
xor U18105 (N_18105,N_12875,N_12420);
xnor U18106 (N_18106,N_10554,N_11326);
nand U18107 (N_18107,N_13806,N_10441);
nor U18108 (N_18108,N_13671,N_13551);
and U18109 (N_18109,N_14343,N_12528);
and U18110 (N_18110,N_14243,N_11269);
and U18111 (N_18111,N_14748,N_10272);
or U18112 (N_18112,N_12048,N_11519);
nor U18113 (N_18113,N_11756,N_14355);
nor U18114 (N_18114,N_14065,N_14068);
and U18115 (N_18115,N_12734,N_12920);
or U18116 (N_18116,N_10994,N_11576);
nor U18117 (N_18117,N_13891,N_13910);
nor U18118 (N_18118,N_14682,N_13828);
and U18119 (N_18119,N_10770,N_10835);
and U18120 (N_18120,N_13609,N_10925);
nand U18121 (N_18121,N_12662,N_11762);
nand U18122 (N_18122,N_11451,N_12845);
xor U18123 (N_18123,N_10088,N_13766);
nand U18124 (N_18124,N_11138,N_11652);
or U18125 (N_18125,N_10399,N_10269);
xor U18126 (N_18126,N_14433,N_10732);
nand U18127 (N_18127,N_14507,N_10297);
or U18128 (N_18128,N_11762,N_10780);
or U18129 (N_18129,N_11522,N_10506);
nor U18130 (N_18130,N_11744,N_12160);
nor U18131 (N_18131,N_12196,N_11254);
and U18132 (N_18132,N_14983,N_11962);
nor U18133 (N_18133,N_12431,N_10420);
or U18134 (N_18134,N_14167,N_14219);
xnor U18135 (N_18135,N_10664,N_12677);
xnor U18136 (N_18136,N_10859,N_11673);
or U18137 (N_18137,N_10201,N_12291);
or U18138 (N_18138,N_13479,N_11548);
xnor U18139 (N_18139,N_10036,N_12278);
nand U18140 (N_18140,N_12825,N_14810);
or U18141 (N_18141,N_12233,N_13101);
nand U18142 (N_18142,N_10049,N_14787);
nand U18143 (N_18143,N_13494,N_11274);
nand U18144 (N_18144,N_11879,N_10130);
nor U18145 (N_18145,N_11978,N_10194);
and U18146 (N_18146,N_14310,N_12427);
or U18147 (N_18147,N_12802,N_13709);
nor U18148 (N_18148,N_12910,N_12989);
or U18149 (N_18149,N_13679,N_12939);
and U18150 (N_18150,N_10931,N_12827);
and U18151 (N_18151,N_14926,N_14487);
and U18152 (N_18152,N_10413,N_12325);
or U18153 (N_18153,N_10406,N_10995);
xnor U18154 (N_18154,N_13547,N_10672);
and U18155 (N_18155,N_12301,N_10226);
nand U18156 (N_18156,N_11100,N_10826);
and U18157 (N_18157,N_13325,N_12760);
or U18158 (N_18158,N_13885,N_11890);
xor U18159 (N_18159,N_11006,N_12337);
and U18160 (N_18160,N_12076,N_11334);
or U18161 (N_18161,N_10588,N_10168);
xor U18162 (N_18162,N_10556,N_14077);
xor U18163 (N_18163,N_12891,N_13553);
and U18164 (N_18164,N_12226,N_14255);
nor U18165 (N_18165,N_14377,N_13819);
or U18166 (N_18166,N_12418,N_11245);
and U18167 (N_18167,N_14440,N_13723);
xor U18168 (N_18168,N_12267,N_13278);
nand U18169 (N_18169,N_10478,N_12916);
and U18170 (N_18170,N_12295,N_11155);
xnor U18171 (N_18171,N_12817,N_13867);
or U18172 (N_18172,N_12511,N_13050);
xor U18173 (N_18173,N_11446,N_12983);
xor U18174 (N_18174,N_11376,N_11195);
and U18175 (N_18175,N_11797,N_13391);
and U18176 (N_18176,N_11110,N_13126);
or U18177 (N_18177,N_12237,N_14019);
and U18178 (N_18178,N_11165,N_11570);
or U18179 (N_18179,N_10776,N_10328);
nor U18180 (N_18180,N_12569,N_10934);
and U18181 (N_18181,N_10680,N_10267);
nand U18182 (N_18182,N_12488,N_12546);
or U18183 (N_18183,N_12445,N_14267);
nand U18184 (N_18184,N_10728,N_11749);
nand U18185 (N_18185,N_14757,N_10260);
nor U18186 (N_18186,N_14211,N_10919);
and U18187 (N_18187,N_11585,N_10671);
or U18188 (N_18188,N_11873,N_14215);
and U18189 (N_18189,N_14038,N_12737);
nand U18190 (N_18190,N_12659,N_12787);
xor U18191 (N_18191,N_10102,N_14107);
or U18192 (N_18192,N_14047,N_11703);
or U18193 (N_18193,N_12208,N_13385);
nor U18194 (N_18194,N_11992,N_14156);
nand U18195 (N_18195,N_11804,N_13616);
or U18196 (N_18196,N_12710,N_13532);
or U18197 (N_18197,N_12074,N_11862);
or U18198 (N_18198,N_10750,N_12023);
or U18199 (N_18199,N_10933,N_12980);
xnor U18200 (N_18200,N_10405,N_13328);
and U18201 (N_18201,N_12281,N_12096);
xnor U18202 (N_18202,N_10480,N_12742);
or U18203 (N_18203,N_10935,N_13194);
or U18204 (N_18204,N_14232,N_13392);
or U18205 (N_18205,N_12409,N_11998);
nand U18206 (N_18206,N_14034,N_12001);
or U18207 (N_18207,N_13364,N_13905);
nor U18208 (N_18208,N_11509,N_13966);
or U18209 (N_18209,N_10818,N_10378);
xnor U18210 (N_18210,N_10261,N_13846);
or U18211 (N_18211,N_13166,N_10348);
and U18212 (N_18212,N_10142,N_11108);
nand U18213 (N_18213,N_11912,N_14904);
xor U18214 (N_18214,N_12478,N_11925);
nand U18215 (N_18215,N_10488,N_14004);
nand U18216 (N_18216,N_12747,N_10775);
and U18217 (N_18217,N_10728,N_12683);
nand U18218 (N_18218,N_10331,N_11045);
nor U18219 (N_18219,N_10643,N_10554);
or U18220 (N_18220,N_12266,N_10339);
nand U18221 (N_18221,N_12170,N_12009);
nor U18222 (N_18222,N_13005,N_13877);
nand U18223 (N_18223,N_13332,N_10109);
xor U18224 (N_18224,N_12607,N_10804);
nor U18225 (N_18225,N_11928,N_13962);
xnor U18226 (N_18226,N_14407,N_11813);
nand U18227 (N_18227,N_11593,N_11558);
and U18228 (N_18228,N_13346,N_14315);
nor U18229 (N_18229,N_14000,N_12355);
xor U18230 (N_18230,N_14606,N_14019);
nand U18231 (N_18231,N_14935,N_11985);
nor U18232 (N_18232,N_11994,N_13917);
and U18233 (N_18233,N_10141,N_12883);
or U18234 (N_18234,N_14416,N_14479);
xnor U18235 (N_18235,N_10421,N_10161);
and U18236 (N_18236,N_13875,N_10723);
nand U18237 (N_18237,N_10367,N_13269);
and U18238 (N_18238,N_10319,N_12841);
and U18239 (N_18239,N_13697,N_10197);
and U18240 (N_18240,N_12373,N_13787);
xor U18241 (N_18241,N_13171,N_11751);
and U18242 (N_18242,N_10735,N_11047);
xnor U18243 (N_18243,N_14416,N_10565);
and U18244 (N_18244,N_11615,N_14933);
nand U18245 (N_18245,N_13082,N_14271);
nor U18246 (N_18246,N_10096,N_13780);
and U18247 (N_18247,N_12138,N_10762);
nor U18248 (N_18248,N_12071,N_11798);
or U18249 (N_18249,N_13521,N_13335);
xor U18250 (N_18250,N_13869,N_11262);
or U18251 (N_18251,N_12801,N_12336);
xnor U18252 (N_18252,N_12828,N_11518);
and U18253 (N_18253,N_13430,N_14268);
nand U18254 (N_18254,N_12323,N_14915);
nand U18255 (N_18255,N_12963,N_13405);
or U18256 (N_18256,N_11653,N_14062);
nor U18257 (N_18257,N_14520,N_11038);
or U18258 (N_18258,N_11319,N_12547);
and U18259 (N_18259,N_11082,N_14938);
xnor U18260 (N_18260,N_14702,N_10390);
nor U18261 (N_18261,N_12983,N_14184);
xor U18262 (N_18262,N_12367,N_12932);
and U18263 (N_18263,N_10981,N_14470);
nor U18264 (N_18264,N_13247,N_13619);
xnor U18265 (N_18265,N_12686,N_14933);
nor U18266 (N_18266,N_14787,N_10218);
or U18267 (N_18267,N_13852,N_13337);
and U18268 (N_18268,N_10490,N_12598);
and U18269 (N_18269,N_14226,N_11711);
nand U18270 (N_18270,N_13419,N_10393);
nand U18271 (N_18271,N_10291,N_10888);
xnor U18272 (N_18272,N_13757,N_14830);
nand U18273 (N_18273,N_10113,N_11770);
or U18274 (N_18274,N_11085,N_13791);
nand U18275 (N_18275,N_12120,N_13919);
and U18276 (N_18276,N_13233,N_14807);
and U18277 (N_18277,N_13784,N_12797);
nor U18278 (N_18278,N_12275,N_10988);
xor U18279 (N_18279,N_11441,N_12180);
and U18280 (N_18280,N_13613,N_12104);
and U18281 (N_18281,N_14859,N_12670);
xnor U18282 (N_18282,N_11265,N_11240);
nand U18283 (N_18283,N_14574,N_13767);
nand U18284 (N_18284,N_11063,N_12031);
and U18285 (N_18285,N_12353,N_11026);
and U18286 (N_18286,N_12278,N_12316);
nand U18287 (N_18287,N_13352,N_11304);
nor U18288 (N_18288,N_12386,N_13578);
xnor U18289 (N_18289,N_13568,N_13345);
xnor U18290 (N_18290,N_10075,N_14649);
and U18291 (N_18291,N_11686,N_12696);
and U18292 (N_18292,N_12709,N_12687);
nor U18293 (N_18293,N_12313,N_13300);
or U18294 (N_18294,N_13419,N_10545);
nor U18295 (N_18295,N_12147,N_11424);
xnor U18296 (N_18296,N_11988,N_13797);
and U18297 (N_18297,N_13675,N_14792);
or U18298 (N_18298,N_12699,N_11786);
xnor U18299 (N_18299,N_13324,N_10802);
and U18300 (N_18300,N_14319,N_10988);
and U18301 (N_18301,N_10467,N_11830);
nor U18302 (N_18302,N_11286,N_11931);
or U18303 (N_18303,N_10559,N_14796);
and U18304 (N_18304,N_10914,N_14897);
nand U18305 (N_18305,N_10471,N_13902);
or U18306 (N_18306,N_11741,N_10305);
and U18307 (N_18307,N_12551,N_12104);
or U18308 (N_18308,N_11024,N_11504);
and U18309 (N_18309,N_10601,N_14681);
xnor U18310 (N_18310,N_14040,N_10179);
and U18311 (N_18311,N_10001,N_10620);
nor U18312 (N_18312,N_14553,N_12317);
xnor U18313 (N_18313,N_10140,N_14976);
nor U18314 (N_18314,N_12939,N_10216);
nor U18315 (N_18315,N_11395,N_10831);
xor U18316 (N_18316,N_13152,N_10072);
and U18317 (N_18317,N_11420,N_10423);
and U18318 (N_18318,N_13659,N_10473);
and U18319 (N_18319,N_12944,N_10150);
and U18320 (N_18320,N_11572,N_13268);
xor U18321 (N_18321,N_13125,N_14038);
xnor U18322 (N_18322,N_12870,N_12982);
nand U18323 (N_18323,N_14953,N_12902);
nor U18324 (N_18324,N_13716,N_13785);
nor U18325 (N_18325,N_13422,N_10895);
or U18326 (N_18326,N_13578,N_10964);
or U18327 (N_18327,N_12295,N_11017);
nand U18328 (N_18328,N_12348,N_14319);
nand U18329 (N_18329,N_14796,N_13269);
and U18330 (N_18330,N_12076,N_12141);
or U18331 (N_18331,N_10804,N_14459);
xnor U18332 (N_18332,N_12099,N_14892);
nand U18333 (N_18333,N_12809,N_10947);
and U18334 (N_18334,N_10955,N_12407);
xnor U18335 (N_18335,N_12680,N_14395);
or U18336 (N_18336,N_14346,N_11901);
xnor U18337 (N_18337,N_14810,N_10522);
nor U18338 (N_18338,N_14378,N_11636);
nand U18339 (N_18339,N_10243,N_12920);
xnor U18340 (N_18340,N_12591,N_12453);
nand U18341 (N_18341,N_10431,N_14229);
nor U18342 (N_18342,N_11750,N_11398);
xor U18343 (N_18343,N_10904,N_13097);
or U18344 (N_18344,N_13424,N_10747);
or U18345 (N_18345,N_13220,N_12744);
and U18346 (N_18346,N_11231,N_12701);
and U18347 (N_18347,N_10991,N_14169);
nand U18348 (N_18348,N_13927,N_13163);
or U18349 (N_18349,N_11390,N_11011);
or U18350 (N_18350,N_12605,N_13804);
and U18351 (N_18351,N_12513,N_13613);
nand U18352 (N_18352,N_11583,N_14082);
or U18353 (N_18353,N_14657,N_13517);
or U18354 (N_18354,N_10689,N_12129);
and U18355 (N_18355,N_11515,N_11954);
nand U18356 (N_18356,N_14052,N_13148);
nor U18357 (N_18357,N_10935,N_13023);
nor U18358 (N_18358,N_14659,N_14652);
nand U18359 (N_18359,N_13979,N_14637);
xnor U18360 (N_18360,N_12113,N_13892);
xnor U18361 (N_18361,N_11546,N_10640);
or U18362 (N_18362,N_13882,N_12557);
or U18363 (N_18363,N_11451,N_10104);
xor U18364 (N_18364,N_13140,N_13322);
and U18365 (N_18365,N_12473,N_11975);
and U18366 (N_18366,N_11217,N_12834);
or U18367 (N_18367,N_11334,N_10115);
xnor U18368 (N_18368,N_11310,N_13810);
nor U18369 (N_18369,N_12135,N_11278);
xnor U18370 (N_18370,N_14195,N_10568);
and U18371 (N_18371,N_11102,N_11684);
nor U18372 (N_18372,N_13843,N_11151);
nand U18373 (N_18373,N_13536,N_12996);
nand U18374 (N_18374,N_13065,N_13649);
nor U18375 (N_18375,N_14332,N_11807);
nor U18376 (N_18376,N_13941,N_14086);
or U18377 (N_18377,N_14022,N_13475);
nand U18378 (N_18378,N_10632,N_13020);
nand U18379 (N_18379,N_14972,N_10671);
and U18380 (N_18380,N_12917,N_11907);
nor U18381 (N_18381,N_11490,N_12457);
nor U18382 (N_18382,N_10010,N_13766);
nor U18383 (N_18383,N_14728,N_11871);
nor U18384 (N_18384,N_14191,N_10931);
nor U18385 (N_18385,N_13712,N_12178);
nand U18386 (N_18386,N_12495,N_11763);
nand U18387 (N_18387,N_11762,N_13717);
xnor U18388 (N_18388,N_11567,N_13107);
xnor U18389 (N_18389,N_14794,N_12614);
or U18390 (N_18390,N_14522,N_14268);
nand U18391 (N_18391,N_12307,N_14524);
nand U18392 (N_18392,N_12629,N_12601);
xor U18393 (N_18393,N_14880,N_12431);
or U18394 (N_18394,N_14776,N_12479);
nand U18395 (N_18395,N_13691,N_14013);
or U18396 (N_18396,N_12268,N_13006);
and U18397 (N_18397,N_11291,N_13617);
or U18398 (N_18398,N_10470,N_10727);
nand U18399 (N_18399,N_10371,N_13127);
nand U18400 (N_18400,N_14492,N_14366);
nor U18401 (N_18401,N_11765,N_13552);
nand U18402 (N_18402,N_12422,N_13082);
nor U18403 (N_18403,N_11605,N_13495);
and U18404 (N_18404,N_11394,N_10475);
nor U18405 (N_18405,N_10306,N_14533);
nand U18406 (N_18406,N_14540,N_12613);
xnor U18407 (N_18407,N_12432,N_12685);
xnor U18408 (N_18408,N_12629,N_13014);
and U18409 (N_18409,N_14516,N_10497);
or U18410 (N_18410,N_12679,N_13031);
xnor U18411 (N_18411,N_12292,N_13209);
xor U18412 (N_18412,N_10602,N_10630);
nor U18413 (N_18413,N_14293,N_14582);
nand U18414 (N_18414,N_10207,N_11718);
nand U18415 (N_18415,N_10774,N_11373);
nor U18416 (N_18416,N_14256,N_11586);
nor U18417 (N_18417,N_13080,N_12827);
xnor U18418 (N_18418,N_14484,N_12335);
xor U18419 (N_18419,N_13412,N_14436);
xnor U18420 (N_18420,N_10260,N_14369);
or U18421 (N_18421,N_14202,N_14379);
xnor U18422 (N_18422,N_12067,N_11300);
or U18423 (N_18423,N_13233,N_12180);
xnor U18424 (N_18424,N_14288,N_14605);
and U18425 (N_18425,N_14452,N_11649);
nor U18426 (N_18426,N_12962,N_11410);
nand U18427 (N_18427,N_13685,N_11434);
nand U18428 (N_18428,N_13440,N_13606);
or U18429 (N_18429,N_13164,N_12773);
nor U18430 (N_18430,N_10756,N_10915);
nand U18431 (N_18431,N_11258,N_12184);
nand U18432 (N_18432,N_10741,N_12257);
and U18433 (N_18433,N_12620,N_10688);
nand U18434 (N_18434,N_14355,N_14688);
nand U18435 (N_18435,N_13406,N_13644);
nor U18436 (N_18436,N_14317,N_14660);
or U18437 (N_18437,N_11795,N_14521);
nand U18438 (N_18438,N_13647,N_10616);
and U18439 (N_18439,N_12192,N_13568);
nor U18440 (N_18440,N_14683,N_12635);
nor U18441 (N_18441,N_11285,N_13162);
xor U18442 (N_18442,N_11313,N_11259);
nor U18443 (N_18443,N_14968,N_14944);
and U18444 (N_18444,N_12554,N_12814);
or U18445 (N_18445,N_10623,N_10273);
or U18446 (N_18446,N_12032,N_11787);
nand U18447 (N_18447,N_12901,N_10869);
or U18448 (N_18448,N_13825,N_14822);
or U18449 (N_18449,N_10732,N_14943);
and U18450 (N_18450,N_10035,N_12811);
nand U18451 (N_18451,N_14382,N_12678);
nor U18452 (N_18452,N_13999,N_11497);
and U18453 (N_18453,N_12985,N_12845);
nand U18454 (N_18454,N_14744,N_12321);
and U18455 (N_18455,N_12163,N_10542);
or U18456 (N_18456,N_11608,N_13327);
or U18457 (N_18457,N_11471,N_13405);
xor U18458 (N_18458,N_13684,N_12978);
nand U18459 (N_18459,N_12627,N_14784);
nor U18460 (N_18460,N_13679,N_11705);
and U18461 (N_18461,N_13088,N_11036);
xnor U18462 (N_18462,N_13156,N_13458);
and U18463 (N_18463,N_12884,N_11874);
xnor U18464 (N_18464,N_10864,N_14077);
or U18465 (N_18465,N_11370,N_14116);
nor U18466 (N_18466,N_13517,N_11337);
nand U18467 (N_18467,N_14853,N_14276);
xnor U18468 (N_18468,N_10584,N_11827);
or U18469 (N_18469,N_14204,N_11392);
nor U18470 (N_18470,N_13956,N_11149);
nor U18471 (N_18471,N_14807,N_14454);
and U18472 (N_18472,N_13577,N_11475);
nand U18473 (N_18473,N_11443,N_14802);
nand U18474 (N_18474,N_10226,N_10971);
nor U18475 (N_18475,N_14777,N_13690);
and U18476 (N_18476,N_14107,N_14108);
nand U18477 (N_18477,N_14776,N_12697);
or U18478 (N_18478,N_14078,N_12561);
or U18479 (N_18479,N_14553,N_14762);
and U18480 (N_18480,N_13464,N_11734);
xor U18481 (N_18481,N_12583,N_12067);
nor U18482 (N_18482,N_13678,N_11444);
nor U18483 (N_18483,N_14550,N_14794);
nor U18484 (N_18484,N_14982,N_13119);
nand U18485 (N_18485,N_11695,N_11554);
nand U18486 (N_18486,N_11002,N_14365);
nand U18487 (N_18487,N_13642,N_10060);
or U18488 (N_18488,N_14760,N_12719);
and U18489 (N_18489,N_14425,N_14483);
or U18490 (N_18490,N_13492,N_14581);
xnor U18491 (N_18491,N_14512,N_11543);
nor U18492 (N_18492,N_14070,N_11196);
xor U18493 (N_18493,N_11721,N_10030);
and U18494 (N_18494,N_12746,N_11299);
xnor U18495 (N_18495,N_11523,N_13812);
and U18496 (N_18496,N_13670,N_10674);
nor U18497 (N_18497,N_11687,N_11219);
nor U18498 (N_18498,N_10099,N_10379);
xor U18499 (N_18499,N_10022,N_10065);
xor U18500 (N_18500,N_10222,N_13607);
or U18501 (N_18501,N_11358,N_11189);
or U18502 (N_18502,N_14524,N_11964);
nand U18503 (N_18503,N_13823,N_13375);
and U18504 (N_18504,N_12587,N_13081);
or U18505 (N_18505,N_11617,N_13295);
nor U18506 (N_18506,N_12904,N_12619);
or U18507 (N_18507,N_12058,N_12526);
nor U18508 (N_18508,N_12816,N_12840);
and U18509 (N_18509,N_10122,N_12107);
and U18510 (N_18510,N_12895,N_12479);
xor U18511 (N_18511,N_10408,N_13475);
or U18512 (N_18512,N_10598,N_10111);
or U18513 (N_18513,N_11431,N_13294);
nor U18514 (N_18514,N_14227,N_12714);
xnor U18515 (N_18515,N_14246,N_14038);
xnor U18516 (N_18516,N_10763,N_10592);
xnor U18517 (N_18517,N_13245,N_11967);
xor U18518 (N_18518,N_11180,N_10278);
nor U18519 (N_18519,N_13631,N_14727);
and U18520 (N_18520,N_11172,N_12157);
and U18521 (N_18521,N_12677,N_10263);
and U18522 (N_18522,N_10757,N_11490);
and U18523 (N_18523,N_12100,N_12001);
or U18524 (N_18524,N_14454,N_12031);
or U18525 (N_18525,N_14842,N_11015);
nor U18526 (N_18526,N_12292,N_10184);
nand U18527 (N_18527,N_12814,N_14124);
and U18528 (N_18528,N_11980,N_10699);
or U18529 (N_18529,N_14594,N_11067);
and U18530 (N_18530,N_13237,N_13333);
and U18531 (N_18531,N_13166,N_13983);
nand U18532 (N_18532,N_10015,N_11715);
and U18533 (N_18533,N_12417,N_12741);
nand U18534 (N_18534,N_12045,N_14893);
xnor U18535 (N_18535,N_11034,N_13221);
nor U18536 (N_18536,N_10627,N_10741);
xnor U18537 (N_18537,N_10578,N_12633);
xnor U18538 (N_18538,N_12005,N_11391);
or U18539 (N_18539,N_12803,N_14339);
or U18540 (N_18540,N_12052,N_14740);
nor U18541 (N_18541,N_12803,N_14723);
xnor U18542 (N_18542,N_13381,N_12732);
nand U18543 (N_18543,N_14837,N_11444);
xor U18544 (N_18544,N_14319,N_10961);
nor U18545 (N_18545,N_11612,N_12515);
nor U18546 (N_18546,N_12886,N_10005);
nor U18547 (N_18547,N_10863,N_12641);
and U18548 (N_18548,N_14280,N_13308);
nand U18549 (N_18549,N_10303,N_12675);
and U18550 (N_18550,N_12801,N_14470);
and U18551 (N_18551,N_14460,N_11139);
or U18552 (N_18552,N_12173,N_12972);
and U18553 (N_18553,N_13059,N_13429);
xnor U18554 (N_18554,N_10118,N_11188);
or U18555 (N_18555,N_12448,N_12994);
nand U18556 (N_18556,N_11030,N_10267);
or U18557 (N_18557,N_13173,N_10034);
or U18558 (N_18558,N_11381,N_11759);
and U18559 (N_18559,N_12173,N_10434);
or U18560 (N_18560,N_12058,N_12075);
nand U18561 (N_18561,N_11660,N_11761);
and U18562 (N_18562,N_10585,N_11078);
nor U18563 (N_18563,N_14707,N_14488);
and U18564 (N_18564,N_13121,N_13334);
and U18565 (N_18565,N_11556,N_11217);
nor U18566 (N_18566,N_11867,N_12355);
and U18567 (N_18567,N_12785,N_13692);
nor U18568 (N_18568,N_14028,N_10509);
and U18569 (N_18569,N_12971,N_12276);
nor U18570 (N_18570,N_13386,N_11751);
xor U18571 (N_18571,N_11131,N_13956);
xor U18572 (N_18572,N_13519,N_12277);
nor U18573 (N_18573,N_13583,N_10814);
and U18574 (N_18574,N_14251,N_12069);
nor U18575 (N_18575,N_12654,N_11727);
xnor U18576 (N_18576,N_11848,N_10072);
nand U18577 (N_18577,N_13941,N_13461);
xor U18578 (N_18578,N_14085,N_13847);
and U18579 (N_18579,N_14804,N_13623);
nand U18580 (N_18580,N_10345,N_13355);
xor U18581 (N_18581,N_14089,N_14399);
xnor U18582 (N_18582,N_14566,N_13402);
nor U18583 (N_18583,N_11632,N_10797);
or U18584 (N_18584,N_13745,N_14102);
or U18585 (N_18585,N_11061,N_10712);
xnor U18586 (N_18586,N_13783,N_14603);
and U18587 (N_18587,N_10007,N_12953);
nor U18588 (N_18588,N_13698,N_14573);
and U18589 (N_18589,N_12981,N_11925);
and U18590 (N_18590,N_13252,N_10111);
xor U18591 (N_18591,N_11242,N_14275);
and U18592 (N_18592,N_11528,N_13569);
xnor U18593 (N_18593,N_11702,N_14172);
nand U18594 (N_18594,N_14812,N_11686);
nor U18595 (N_18595,N_11147,N_12373);
nor U18596 (N_18596,N_13370,N_14301);
nand U18597 (N_18597,N_10600,N_10330);
and U18598 (N_18598,N_13348,N_12028);
or U18599 (N_18599,N_10536,N_11384);
xor U18600 (N_18600,N_10749,N_11765);
and U18601 (N_18601,N_13795,N_12071);
nor U18602 (N_18602,N_14547,N_10045);
nor U18603 (N_18603,N_10464,N_11573);
nand U18604 (N_18604,N_10391,N_13017);
or U18605 (N_18605,N_12424,N_10431);
nand U18606 (N_18606,N_13423,N_10868);
nand U18607 (N_18607,N_14726,N_12564);
or U18608 (N_18608,N_11874,N_11039);
xnor U18609 (N_18609,N_11352,N_13401);
nand U18610 (N_18610,N_14601,N_10053);
nor U18611 (N_18611,N_10767,N_10677);
nor U18612 (N_18612,N_12642,N_12529);
and U18613 (N_18613,N_10527,N_11507);
xor U18614 (N_18614,N_12819,N_13438);
and U18615 (N_18615,N_13607,N_13054);
or U18616 (N_18616,N_12767,N_11524);
nor U18617 (N_18617,N_11570,N_11688);
xnor U18618 (N_18618,N_14026,N_10589);
nor U18619 (N_18619,N_12429,N_10279);
or U18620 (N_18620,N_10923,N_13844);
or U18621 (N_18621,N_10753,N_10531);
and U18622 (N_18622,N_13108,N_12263);
nor U18623 (N_18623,N_14878,N_11386);
nor U18624 (N_18624,N_12374,N_10129);
or U18625 (N_18625,N_14106,N_14534);
and U18626 (N_18626,N_11835,N_11555);
nor U18627 (N_18627,N_13040,N_11501);
nand U18628 (N_18628,N_13051,N_10378);
and U18629 (N_18629,N_11223,N_12605);
xnor U18630 (N_18630,N_11237,N_13300);
xnor U18631 (N_18631,N_10073,N_14124);
and U18632 (N_18632,N_11394,N_10611);
or U18633 (N_18633,N_10792,N_10389);
and U18634 (N_18634,N_14549,N_12369);
nor U18635 (N_18635,N_13855,N_12768);
or U18636 (N_18636,N_12229,N_11225);
and U18637 (N_18637,N_11437,N_10163);
or U18638 (N_18638,N_12261,N_12686);
or U18639 (N_18639,N_11911,N_12251);
xor U18640 (N_18640,N_10914,N_13056);
and U18641 (N_18641,N_13797,N_13008);
and U18642 (N_18642,N_10127,N_12518);
and U18643 (N_18643,N_14191,N_12004);
xnor U18644 (N_18644,N_13845,N_13732);
nor U18645 (N_18645,N_10183,N_10399);
nor U18646 (N_18646,N_10772,N_13456);
nand U18647 (N_18647,N_11148,N_11946);
xor U18648 (N_18648,N_12029,N_11953);
and U18649 (N_18649,N_11254,N_11977);
nor U18650 (N_18650,N_14046,N_10188);
nand U18651 (N_18651,N_10087,N_12991);
nand U18652 (N_18652,N_12866,N_10814);
xor U18653 (N_18653,N_13220,N_10927);
xnor U18654 (N_18654,N_14720,N_12667);
nand U18655 (N_18655,N_14942,N_11306);
and U18656 (N_18656,N_10459,N_13059);
nand U18657 (N_18657,N_14596,N_11619);
nor U18658 (N_18658,N_11896,N_12058);
nand U18659 (N_18659,N_12675,N_13289);
nand U18660 (N_18660,N_13909,N_13774);
or U18661 (N_18661,N_10320,N_11283);
and U18662 (N_18662,N_14066,N_11223);
nor U18663 (N_18663,N_11485,N_14763);
xor U18664 (N_18664,N_12827,N_13648);
nor U18665 (N_18665,N_14063,N_10922);
nand U18666 (N_18666,N_13415,N_10603);
xnor U18667 (N_18667,N_14508,N_13706);
and U18668 (N_18668,N_13768,N_11487);
nor U18669 (N_18669,N_11481,N_13471);
and U18670 (N_18670,N_13088,N_13192);
nor U18671 (N_18671,N_14416,N_10411);
and U18672 (N_18672,N_11456,N_12366);
or U18673 (N_18673,N_13835,N_12036);
nand U18674 (N_18674,N_10825,N_10996);
and U18675 (N_18675,N_14805,N_10240);
or U18676 (N_18676,N_12812,N_12485);
xnor U18677 (N_18677,N_14443,N_14483);
and U18678 (N_18678,N_12510,N_11131);
or U18679 (N_18679,N_10531,N_10701);
nor U18680 (N_18680,N_11951,N_12685);
nand U18681 (N_18681,N_12954,N_12563);
xor U18682 (N_18682,N_14345,N_10488);
and U18683 (N_18683,N_10886,N_12972);
or U18684 (N_18684,N_10049,N_10058);
nor U18685 (N_18685,N_10054,N_10471);
or U18686 (N_18686,N_14324,N_13248);
or U18687 (N_18687,N_14070,N_12673);
and U18688 (N_18688,N_11582,N_10479);
and U18689 (N_18689,N_14527,N_13559);
or U18690 (N_18690,N_14897,N_13070);
and U18691 (N_18691,N_10622,N_13902);
nor U18692 (N_18692,N_10714,N_10821);
nor U18693 (N_18693,N_10509,N_13217);
or U18694 (N_18694,N_13028,N_12075);
or U18695 (N_18695,N_12575,N_12110);
nand U18696 (N_18696,N_10186,N_10443);
xor U18697 (N_18697,N_11942,N_11770);
xor U18698 (N_18698,N_12436,N_12831);
nor U18699 (N_18699,N_14378,N_14333);
nor U18700 (N_18700,N_12787,N_11918);
nor U18701 (N_18701,N_10780,N_13190);
or U18702 (N_18702,N_10925,N_12859);
and U18703 (N_18703,N_14291,N_13368);
or U18704 (N_18704,N_12323,N_10920);
and U18705 (N_18705,N_11214,N_10579);
or U18706 (N_18706,N_12818,N_11867);
and U18707 (N_18707,N_10815,N_10760);
or U18708 (N_18708,N_10273,N_10822);
nor U18709 (N_18709,N_13407,N_12291);
nand U18710 (N_18710,N_12400,N_12251);
xnor U18711 (N_18711,N_13434,N_14456);
nor U18712 (N_18712,N_14503,N_10932);
nor U18713 (N_18713,N_12127,N_11422);
or U18714 (N_18714,N_10306,N_13066);
nand U18715 (N_18715,N_12668,N_12508);
xnor U18716 (N_18716,N_11441,N_14131);
nand U18717 (N_18717,N_13380,N_11584);
nor U18718 (N_18718,N_11717,N_11627);
and U18719 (N_18719,N_14418,N_11411);
and U18720 (N_18720,N_13511,N_10551);
xnor U18721 (N_18721,N_12095,N_11345);
xnor U18722 (N_18722,N_13418,N_12124);
nand U18723 (N_18723,N_11378,N_14672);
nand U18724 (N_18724,N_13784,N_11795);
nor U18725 (N_18725,N_11871,N_14770);
nand U18726 (N_18726,N_11722,N_12689);
xor U18727 (N_18727,N_13576,N_12171);
xnor U18728 (N_18728,N_12251,N_11192);
or U18729 (N_18729,N_13883,N_14105);
xor U18730 (N_18730,N_13536,N_14518);
xor U18731 (N_18731,N_10142,N_14481);
nor U18732 (N_18732,N_14929,N_11184);
nor U18733 (N_18733,N_11070,N_11827);
xor U18734 (N_18734,N_14238,N_11703);
nand U18735 (N_18735,N_14367,N_13735);
xnor U18736 (N_18736,N_11398,N_14397);
or U18737 (N_18737,N_10610,N_11545);
nand U18738 (N_18738,N_12527,N_13897);
nand U18739 (N_18739,N_10409,N_14690);
and U18740 (N_18740,N_11573,N_10885);
xnor U18741 (N_18741,N_10328,N_12401);
nor U18742 (N_18742,N_11466,N_10227);
xor U18743 (N_18743,N_11873,N_14014);
xnor U18744 (N_18744,N_10913,N_14273);
xnor U18745 (N_18745,N_13097,N_11552);
xor U18746 (N_18746,N_11495,N_12902);
xor U18747 (N_18747,N_11173,N_14717);
and U18748 (N_18748,N_12295,N_12549);
xnor U18749 (N_18749,N_14364,N_12793);
nor U18750 (N_18750,N_11368,N_14452);
nand U18751 (N_18751,N_11718,N_11411);
nor U18752 (N_18752,N_11026,N_14543);
nand U18753 (N_18753,N_11160,N_14822);
xor U18754 (N_18754,N_11941,N_14546);
nand U18755 (N_18755,N_11287,N_11648);
or U18756 (N_18756,N_13032,N_13340);
xor U18757 (N_18757,N_11128,N_13686);
xor U18758 (N_18758,N_14599,N_12647);
nor U18759 (N_18759,N_13305,N_13400);
nand U18760 (N_18760,N_11166,N_11592);
nor U18761 (N_18761,N_10798,N_14380);
and U18762 (N_18762,N_11641,N_14867);
nor U18763 (N_18763,N_12272,N_14831);
or U18764 (N_18764,N_14256,N_12257);
or U18765 (N_18765,N_14873,N_14073);
and U18766 (N_18766,N_12537,N_11670);
or U18767 (N_18767,N_10297,N_11296);
nor U18768 (N_18768,N_10751,N_11027);
nor U18769 (N_18769,N_12713,N_11868);
and U18770 (N_18770,N_11632,N_10207);
nand U18771 (N_18771,N_11591,N_12767);
and U18772 (N_18772,N_11784,N_13818);
nor U18773 (N_18773,N_12895,N_11164);
and U18774 (N_18774,N_11530,N_13169);
and U18775 (N_18775,N_10886,N_12553);
xor U18776 (N_18776,N_14697,N_12323);
xor U18777 (N_18777,N_14323,N_13362);
nand U18778 (N_18778,N_10591,N_12062);
and U18779 (N_18779,N_12142,N_10599);
xnor U18780 (N_18780,N_14324,N_10472);
nor U18781 (N_18781,N_10704,N_13239);
or U18782 (N_18782,N_14308,N_12210);
nor U18783 (N_18783,N_12099,N_12576);
xor U18784 (N_18784,N_12260,N_14890);
and U18785 (N_18785,N_10889,N_12111);
xnor U18786 (N_18786,N_12052,N_14786);
and U18787 (N_18787,N_12799,N_11501);
xnor U18788 (N_18788,N_13314,N_13655);
xor U18789 (N_18789,N_13128,N_14559);
and U18790 (N_18790,N_14576,N_14318);
xnor U18791 (N_18791,N_12586,N_13859);
nor U18792 (N_18792,N_10183,N_13612);
or U18793 (N_18793,N_14413,N_12742);
nor U18794 (N_18794,N_12842,N_14322);
xor U18795 (N_18795,N_11446,N_14376);
and U18796 (N_18796,N_11987,N_12999);
xnor U18797 (N_18797,N_14118,N_11325);
and U18798 (N_18798,N_10268,N_13345);
xor U18799 (N_18799,N_11174,N_12758);
and U18800 (N_18800,N_10155,N_11130);
nor U18801 (N_18801,N_13794,N_13071);
and U18802 (N_18802,N_12233,N_11492);
nor U18803 (N_18803,N_10480,N_14471);
nor U18804 (N_18804,N_11479,N_13474);
or U18805 (N_18805,N_14672,N_12107);
and U18806 (N_18806,N_10512,N_10223);
nand U18807 (N_18807,N_12776,N_11163);
and U18808 (N_18808,N_11597,N_11817);
or U18809 (N_18809,N_14419,N_10557);
nand U18810 (N_18810,N_12925,N_10709);
xor U18811 (N_18811,N_14985,N_14414);
xor U18812 (N_18812,N_14860,N_10303);
and U18813 (N_18813,N_10170,N_13842);
or U18814 (N_18814,N_11086,N_12326);
xnor U18815 (N_18815,N_14850,N_12742);
xor U18816 (N_18816,N_12042,N_14438);
and U18817 (N_18817,N_14331,N_14309);
nand U18818 (N_18818,N_12754,N_11131);
nor U18819 (N_18819,N_14500,N_10179);
nand U18820 (N_18820,N_12563,N_12327);
and U18821 (N_18821,N_11515,N_11424);
xor U18822 (N_18822,N_10141,N_10430);
or U18823 (N_18823,N_14150,N_10493);
nand U18824 (N_18824,N_10523,N_12520);
and U18825 (N_18825,N_14425,N_10213);
and U18826 (N_18826,N_10684,N_13461);
or U18827 (N_18827,N_13760,N_14902);
or U18828 (N_18828,N_12224,N_14743);
or U18829 (N_18829,N_10155,N_14032);
or U18830 (N_18830,N_11652,N_13254);
nand U18831 (N_18831,N_10422,N_11490);
or U18832 (N_18832,N_14705,N_12370);
and U18833 (N_18833,N_11569,N_10431);
nand U18834 (N_18834,N_11832,N_14918);
xnor U18835 (N_18835,N_11681,N_14240);
nor U18836 (N_18836,N_14266,N_11530);
xor U18837 (N_18837,N_12238,N_14215);
or U18838 (N_18838,N_13247,N_14321);
or U18839 (N_18839,N_13565,N_12459);
or U18840 (N_18840,N_14658,N_11577);
nand U18841 (N_18841,N_14356,N_12173);
and U18842 (N_18842,N_14654,N_13245);
and U18843 (N_18843,N_12324,N_14903);
nand U18844 (N_18844,N_14711,N_10429);
and U18845 (N_18845,N_13339,N_10635);
and U18846 (N_18846,N_10313,N_12424);
nand U18847 (N_18847,N_14365,N_13257);
and U18848 (N_18848,N_12502,N_12852);
nor U18849 (N_18849,N_11032,N_13245);
or U18850 (N_18850,N_13936,N_13022);
or U18851 (N_18851,N_11487,N_13769);
or U18852 (N_18852,N_10002,N_14238);
xor U18853 (N_18853,N_11771,N_12189);
and U18854 (N_18854,N_12074,N_10432);
nor U18855 (N_18855,N_12243,N_14374);
nor U18856 (N_18856,N_14362,N_13042);
xnor U18857 (N_18857,N_10186,N_11659);
or U18858 (N_18858,N_12901,N_13333);
nand U18859 (N_18859,N_13073,N_12228);
nand U18860 (N_18860,N_13049,N_10430);
or U18861 (N_18861,N_13218,N_11222);
nand U18862 (N_18862,N_13133,N_13800);
nor U18863 (N_18863,N_12204,N_12490);
nand U18864 (N_18864,N_14238,N_13745);
or U18865 (N_18865,N_14010,N_14638);
nand U18866 (N_18866,N_13396,N_12425);
xnor U18867 (N_18867,N_12074,N_13522);
nor U18868 (N_18868,N_12398,N_10261);
or U18869 (N_18869,N_12713,N_10006);
and U18870 (N_18870,N_11336,N_12179);
nor U18871 (N_18871,N_12727,N_11932);
nand U18872 (N_18872,N_12298,N_10843);
or U18873 (N_18873,N_14623,N_13937);
or U18874 (N_18874,N_13616,N_10815);
xor U18875 (N_18875,N_14995,N_10590);
and U18876 (N_18876,N_10603,N_13384);
nor U18877 (N_18877,N_13191,N_13955);
nand U18878 (N_18878,N_10937,N_14691);
nand U18879 (N_18879,N_11665,N_12322);
xnor U18880 (N_18880,N_12994,N_13434);
nand U18881 (N_18881,N_13196,N_11602);
nand U18882 (N_18882,N_13276,N_11754);
nand U18883 (N_18883,N_13241,N_14923);
nor U18884 (N_18884,N_11280,N_12392);
and U18885 (N_18885,N_13852,N_12570);
xor U18886 (N_18886,N_10074,N_12838);
or U18887 (N_18887,N_11890,N_14426);
xor U18888 (N_18888,N_13385,N_11966);
or U18889 (N_18889,N_12793,N_12245);
nand U18890 (N_18890,N_13192,N_14941);
nor U18891 (N_18891,N_12593,N_14992);
or U18892 (N_18892,N_13291,N_12387);
nor U18893 (N_18893,N_10208,N_12807);
nor U18894 (N_18894,N_14633,N_11000);
nand U18895 (N_18895,N_13326,N_10094);
nand U18896 (N_18896,N_11371,N_10054);
nand U18897 (N_18897,N_12260,N_11103);
xnor U18898 (N_18898,N_12200,N_11103);
nor U18899 (N_18899,N_14637,N_14654);
or U18900 (N_18900,N_13809,N_10432);
nor U18901 (N_18901,N_12170,N_10329);
and U18902 (N_18902,N_10188,N_12285);
xor U18903 (N_18903,N_14330,N_14352);
and U18904 (N_18904,N_12507,N_13256);
nand U18905 (N_18905,N_10528,N_13654);
nand U18906 (N_18906,N_13166,N_10511);
nand U18907 (N_18907,N_12475,N_14221);
nand U18908 (N_18908,N_12331,N_11944);
and U18909 (N_18909,N_14108,N_10036);
nand U18910 (N_18910,N_13004,N_11824);
nor U18911 (N_18911,N_10466,N_10983);
and U18912 (N_18912,N_12831,N_14939);
nor U18913 (N_18913,N_10775,N_12302);
or U18914 (N_18914,N_13548,N_11110);
nand U18915 (N_18915,N_13613,N_10269);
or U18916 (N_18916,N_11597,N_13707);
xnor U18917 (N_18917,N_13873,N_11006);
xor U18918 (N_18918,N_13038,N_12083);
xor U18919 (N_18919,N_14779,N_10827);
or U18920 (N_18920,N_10468,N_12976);
nor U18921 (N_18921,N_13989,N_12943);
and U18922 (N_18922,N_12998,N_13849);
nand U18923 (N_18923,N_12654,N_14581);
xor U18924 (N_18924,N_13463,N_13627);
and U18925 (N_18925,N_10662,N_14792);
and U18926 (N_18926,N_11635,N_10535);
or U18927 (N_18927,N_10104,N_14444);
nor U18928 (N_18928,N_11162,N_11208);
and U18929 (N_18929,N_12996,N_11747);
xor U18930 (N_18930,N_11975,N_12278);
xnor U18931 (N_18931,N_14835,N_11604);
and U18932 (N_18932,N_10164,N_12803);
xnor U18933 (N_18933,N_13226,N_13157);
or U18934 (N_18934,N_12567,N_13606);
or U18935 (N_18935,N_13347,N_14305);
and U18936 (N_18936,N_10888,N_12794);
nand U18937 (N_18937,N_10716,N_11187);
and U18938 (N_18938,N_14300,N_10188);
xnor U18939 (N_18939,N_14604,N_11717);
nor U18940 (N_18940,N_12926,N_14462);
nor U18941 (N_18941,N_12074,N_11601);
nand U18942 (N_18942,N_12329,N_14675);
xnor U18943 (N_18943,N_13208,N_14729);
xor U18944 (N_18944,N_12139,N_14958);
xnor U18945 (N_18945,N_13061,N_13977);
or U18946 (N_18946,N_13755,N_14518);
and U18947 (N_18947,N_11809,N_10545);
or U18948 (N_18948,N_13084,N_10230);
or U18949 (N_18949,N_12954,N_14464);
xor U18950 (N_18950,N_13171,N_12042);
nor U18951 (N_18951,N_11662,N_12201);
and U18952 (N_18952,N_13792,N_12688);
and U18953 (N_18953,N_14799,N_12801);
nand U18954 (N_18954,N_12221,N_14586);
and U18955 (N_18955,N_11656,N_13721);
and U18956 (N_18956,N_13165,N_10476);
and U18957 (N_18957,N_10994,N_12159);
or U18958 (N_18958,N_13796,N_13651);
xor U18959 (N_18959,N_10113,N_13807);
nor U18960 (N_18960,N_11977,N_12786);
and U18961 (N_18961,N_11301,N_12515);
nand U18962 (N_18962,N_13697,N_10826);
xor U18963 (N_18963,N_12167,N_11048);
and U18964 (N_18964,N_11160,N_13402);
nand U18965 (N_18965,N_10398,N_12830);
and U18966 (N_18966,N_10426,N_11665);
or U18967 (N_18967,N_13985,N_10709);
nand U18968 (N_18968,N_10629,N_11171);
nor U18969 (N_18969,N_14872,N_11558);
or U18970 (N_18970,N_11161,N_11398);
xnor U18971 (N_18971,N_11874,N_11467);
xnor U18972 (N_18972,N_14807,N_13366);
xor U18973 (N_18973,N_11388,N_11600);
nor U18974 (N_18974,N_11642,N_10553);
and U18975 (N_18975,N_11029,N_14569);
nor U18976 (N_18976,N_13143,N_13816);
or U18977 (N_18977,N_14292,N_12116);
xnor U18978 (N_18978,N_14747,N_12208);
or U18979 (N_18979,N_13017,N_12233);
or U18980 (N_18980,N_12274,N_13015);
or U18981 (N_18981,N_14003,N_11738);
xor U18982 (N_18982,N_10668,N_13810);
nand U18983 (N_18983,N_13822,N_11829);
and U18984 (N_18984,N_14137,N_11261);
and U18985 (N_18985,N_11085,N_13972);
and U18986 (N_18986,N_11505,N_11506);
and U18987 (N_18987,N_14512,N_13231);
xnor U18988 (N_18988,N_10048,N_12040);
nor U18989 (N_18989,N_11402,N_13842);
xor U18990 (N_18990,N_11118,N_11960);
nand U18991 (N_18991,N_13553,N_11172);
nor U18992 (N_18992,N_11030,N_10411);
xor U18993 (N_18993,N_13123,N_13550);
nand U18994 (N_18994,N_10875,N_11605);
or U18995 (N_18995,N_12029,N_12374);
nand U18996 (N_18996,N_13570,N_11486);
xnor U18997 (N_18997,N_10036,N_13076);
xnor U18998 (N_18998,N_13723,N_12697);
or U18999 (N_18999,N_12851,N_10269);
nand U19000 (N_19000,N_12383,N_12320);
nand U19001 (N_19001,N_12022,N_12246);
and U19002 (N_19002,N_10035,N_12092);
nand U19003 (N_19003,N_14396,N_10296);
xnor U19004 (N_19004,N_13641,N_10312);
nand U19005 (N_19005,N_14153,N_13762);
and U19006 (N_19006,N_12856,N_11906);
or U19007 (N_19007,N_13249,N_12744);
and U19008 (N_19008,N_13265,N_10680);
xor U19009 (N_19009,N_11259,N_11326);
nor U19010 (N_19010,N_11953,N_14448);
nor U19011 (N_19011,N_11371,N_10154);
and U19012 (N_19012,N_12521,N_11550);
nand U19013 (N_19013,N_11087,N_14130);
xor U19014 (N_19014,N_10624,N_13186);
or U19015 (N_19015,N_10323,N_13265);
nor U19016 (N_19016,N_11748,N_12727);
nor U19017 (N_19017,N_10144,N_14611);
or U19018 (N_19018,N_14820,N_12669);
and U19019 (N_19019,N_10641,N_10096);
or U19020 (N_19020,N_10629,N_13198);
xnor U19021 (N_19021,N_13048,N_12208);
and U19022 (N_19022,N_12130,N_11412);
or U19023 (N_19023,N_11017,N_12883);
nand U19024 (N_19024,N_14698,N_12163);
or U19025 (N_19025,N_11927,N_12075);
nor U19026 (N_19026,N_10883,N_14420);
and U19027 (N_19027,N_10692,N_10508);
xor U19028 (N_19028,N_13385,N_13089);
nor U19029 (N_19029,N_11672,N_13535);
or U19030 (N_19030,N_11833,N_14262);
or U19031 (N_19031,N_12922,N_10584);
xor U19032 (N_19032,N_12020,N_11501);
nor U19033 (N_19033,N_10690,N_14175);
or U19034 (N_19034,N_14989,N_13288);
nand U19035 (N_19035,N_10315,N_10056);
nand U19036 (N_19036,N_12761,N_13944);
nand U19037 (N_19037,N_14457,N_13786);
and U19038 (N_19038,N_11963,N_12994);
xor U19039 (N_19039,N_14215,N_14411);
nand U19040 (N_19040,N_13780,N_14527);
nand U19041 (N_19041,N_13673,N_14596);
nand U19042 (N_19042,N_14993,N_11782);
and U19043 (N_19043,N_12681,N_13255);
and U19044 (N_19044,N_12397,N_11793);
xnor U19045 (N_19045,N_13802,N_10045);
nor U19046 (N_19046,N_13458,N_14462);
xor U19047 (N_19047,N_10469,N_11416);
and U19048 (N_19048,N_10351,N_11810);
or U19049 (N_19049,N_11609,N_13503);
nand U19050 (N_19050,N_11424,N_11436);
and U19051 (N_19051,N_14156,N_11875);
or U19052 (N_19052,N_12812,N_14461);
and U19053 (N_19053,N_12996,N_11886);
nor U19054 (N_19054,N_13936,N_13596);
or U19055 (N_19055,N_14278,N_14178);
nand U19056 (N_19056,N_10617,N_10455);
xnor U19057 (N_19057,N_10970,N_11116);
nand U19058 (N_19058,N_14265,N_12983);
nor U19059 (N_19059,N_12012,N_10651);
or U19060 (N_19060,N_11756,N_10186);
or U19061 (N_19061,N_12428,N_12993);
and U19062 (N_19062,N_13719,N_10064);
or U19063 (N_19063,N_12877,N_11542);
or U19064 (N_19064,N_14897,N_12089);
and U19065 (N_19065,N_11663,N_14498);
or U19066 (N_19066,N_12215,N_13081);
nor U19067 (N_19067,N_12030,N_11778);
and U19068 (N_19068,N_14922,N_10397);
and U19069 (N_19069,N_14062,N_10986);
nand U19070 (N_19070,N_10958,N_11206);
nor U19071 (N_19071,N_11180,N_13662);
nand U19072 (N_19072,N_11894,N_14150);
nand U19073 (N_19073,N_11798,N_10191);
and U19074 (N_19074,N_11140,N_10863);
xnor U19075 (N_19075,N_13265,N_12711);
and U19076 (N_19076,N_12748,N_10968);
xor U19077 (N_19077,N_12157,N_10025);
or U19078 (N_19078,N_10545,N_11380);
and U19079 (N_19079,N_12064,N_12908);
nor U19080 (N_19080,N_10033,N_10654);
nand U19081 (N_19081,N_10487,N_12839);
xnor U19082 (N_19082,N_11032,N_11667);
nand U19083 (N_19083,N_14632,N_10304);
nor U19084 (N_19084,N_11706,N_13312);
and U19085 (N_19085,N_13997,N_11920);
and U19086 (N_19086,N_12551,N_14080);
nand U19087 (N_19087,N_13671,N_10888);
nand U19088 (N_19088,N_13292,N_11034);
and U19089 (N_19089,N_11887,N_13600);
or U19090 (N_19090,N_10894,N_11449);
and U19091 (N_19091,N_13029,N_10627);
nand U19092 (N_19092,N_11174,N_10714);
or U19093 (N_19093,N_12450,N_14567);
nand U19094 (N_19094,N_13280,N_10650);
and U19095 (N_19095,N_14399,N_14752);
and U19096 (N_19096,N_11250,N_13492);
nand U19097 (N_19097,N_13969,N_14025);
nor U19098 (N_19098,N_14792,N_12268);
and U19099 (N_19099,N_11455,N_13745);
or U19100 (N_19100,N_13622,N_11783);
or U19101 (N_19101,N_11285,N_13206);
nand U19102 (N_19102,N_13700,N_13733);
or U19103 (N_19103,N_13741,N_13160);
xor U19104 (N_19104,N_12948,N_11606);
xor U19105 (N_19105,N_14698,N_12225);
nor U19106 (N_19106,N_14805,N_11095);
nand U19107 (N_19107,N_13558,N_11043);
and U19108 (N_19108,N_10692,N_13763);
xnor U19109 (N_19109,N_12114,N_11212);
xor U19110 (N_19110,N_13176,N_14924);
nor U19111 (N_19111,N_12100,N_10776);
xnor U19112 (N_19112,N_10610,N_11792);
nor U19113 (N_19113,N_13115,N_11601);
and U19114 (N_19114,N_13204,N_12731);
nor U19115 (N_19115,N_10275,N_12453);
or U19116 (N_19116,N_10163,N_10722);
or U19117 (N_19117,N_13781,N_13617);
xor U19118 (N_19118,N_14865,N_13671);
nand U19119 (N_19119,N_10074,N_13493);
and U19120 (N_19120,N_14835,N_10430);
and U19121 (N_19121,N_10682,N_12855);
nand U19122 (N_19122,N_11055,N_12116);
nor U19123 (N_19123,N_12289,N_11858);
nand U19124 (N_19124,N_13880,N_14743);
nor U19125 (N_19125,N_12947,N_13616);
nand U19126 (N_19126,N_14519,N_14038);
xor U19127 (N_19127,N_14686,N_11058);
or U19128 (N_19128,N_14326,N_11554);
and U19129 (N_19129,N_12406,N_10850);
xor U19130 (N_19130,N_10745,N_14738);
nor U19131 (N_19131,N_14061,N_14149);
or U19132 (N_19132,N_12759,N_10080);
xor U19133 (N_19133,N_11788,N_12601);
nor U19134 (N_19134,N_14355,N_11302);
nand U19135 (N_19135,N_13455,N_12425);
or U19136 (N_19136,N_12803,N_10595);
nand U19137 (N_19137,N_11147,N_14747);
nor U19138 (N_19138,N_13409,N_11436);
and U19139 (N_19139,N_10509,N_12309);
or U19140 (N_19140,N_11761,N_14388);
xnor U19141 (N_19141,N_10736,N_11774);
nand U19142 (N_19142,N_13917,N_13846);
or U19143 (N_19143,N_14345,N_11019);
nor U19144 (N_19144,N_14363,N_14996);
xor U19145 (N_19145,N_13352,N_13955);
and U19146 (N_19146,N_12635,N_11632);
or U19147 (N_19147,N_11396,N_11430);
nand U19148 (N_19148,N_12066,N_13177);
or U19149 (N_19149,N_12359,N_12549);
and U19150 (N_19150,N_10039,N_13554);
or U19151 (N_19151,N_13745,N_12607);
xor U19152 (N_19152,N_13126,N_12065);
xor U19153 (N_19153,N_11093,N_11642);
and U19154 (N_19154,N_14726,N_11603);
or U19155 (N_19155,N_14311,N_10262);
xnor U19156 (N_19156,N_13576,N_13858);
nor U19157 (N_19157,N_14822,N_12524);
nor U19158 (N_19158,N_13178,N_14562);
nor U19159 (N_19159,N_11346,N_13997);
and U19160 (N_19160,N_14561,N_12934);
or U19161 (N_19161,N_11989,N_10489);
nand U19162 (N_19162,N_10930,N_14628);
or U19163 (N_19163,N_13647,N_14146);
nand U19164 (N_19164,N_14326,N_11855);
nand U19165 (N_19165,N_14208,N_13594);
or U19166 (N_19166,N_13062,N_11946);
xnor U19167 (N_19167,N_12309,N_11386);
xnor U19168 (N_19168,N_12709,N_10503);
nand U19169 (N_19169,N_10417,N_13788);
or U19170 (N_19170,N_14013,N_14657);
or U19171 (N_19171,N_12854,N_11114);
or U19172 (N_19172,N_11366,N_11855);
xnor U19173 (N_19173,N_13673,N_12184);
xor U19174 (N_19174,N_11435,N_10775);
nand U19175 (N_19175,N_14805,N_10705);
or U19176 (N_19176,N_14730,N_12935);
xor U19177 (N_19177,N_12555,N_14034);
or U19178 (N_19178,N_10191,N_11502);
xor U19179 (N_19179,N_13352,N_11315);
nand U19180 (N_19180,N_13401,N_13258);
nand U19181 (N_19181,N_12758,N_14376);
nand U19182 (N_19182,N_11845,N_12334);
nand U19183 (N_19183,N_14196,N_10713);
xor U19184 (N_19184,N_12580,N_11557);
or U19185 (N_19185,N_13798,N_12762);
xnor U19186 (N_19186,N_13664,N_13597);
or U19187 (N_19187,N_11768,N_14693);
xor U19188 (N_19188,N_11495,N_13250);
nor U19189 (N_19189,N_13874,N_10249);
nand U19190 (N_19190,N_14473,N_11597);
nand U19191 (N_19191,N_10882,N_11357);
or U19192 (N_19192,N_13544,N_10327);
nand U19193 (N_19193,N_13602,N_14170);
nand U19194 (N_19194,N_10390,N_12969);
xor U19195 (N_19195,N_14792,N_10191);
and U19196 (N_19196,N_12733,N_11952);
nand U19197 (N_19197,N_13419,N_12911);
and U19198 (N_19198,N_12049,N_11311);
xor U19199 (N_19199,N_10521,N_13877);
or U19200 (N_19200,N_10588,N_10101);
nor U19201 (N_19201,N_14373,N_14884);
or U19202 (N_19202,N_10563,N_14274);
nand U19203 (N_19203,N_10269,N_11237);
xor U19204 (N_19204,N_12311,N_10541);
or U19205 (N_19205,N_14420,N_13922);
xor U19206 (N_19206,N_10597,N_14580);
xor U19207 (N_19207,N_12111,N_10813);
nor U19208 (N_19208,N_13578,N_10236);
nor U19209 (N_19209,N_13134,N_13551);
and U19210 (N_19210,N_12262,N_12873);
nand U19211 (N_19211,N_14833,N_10609);
xor U19212 (N_19212,N_10888,N_12115);
xor U19213 (N_19213,N_14992,N_14686);
nor U19214 (N_19214,N_11205,N_11397);
nand U19215 (N_19215,N_14516,N_11109);
or U19216 (N_19216,N_10017,N_11868);
xor U19217 (N_19217,N_13943,N_14928);
or U19218 (N_19218,N_14358,N_12520);
xor U19219 (N_19219,N_11879,N_14541);
or U19220 (N_19220,N_13033,N_12122);
and U19221 (N_19221,N_12924,N_14528);
and U19222 (N_19222,N_13514,N_14279);
nor U19223 (N_19223,N_14936,N_14550);
or U19224 (N_19224,N_12015,N_11837);
or U19225 (N_19225,N_10734,N_14629);
nor U19226 (N_19226,N_12453,N_14390);
or U19227 (N_19227,N_13937,N_11526);
xor U19228 (N_19228,N_10530,N_13671);
nor U19229 (N_19229,N_10456,N_13770);
or U19230 (N_19230,N_12645,N_11560);
nor U19231 (N_19231,N_14665,N_11247);
nor U19232 (N_19232,N_10953,N_12673);
nand U19233 (N_19233,N_14454,N_11605);
xnor U19234 (N_19234,N_13508,N_10313);
and U19235 (N_19235,N_12184,N_11447);
xnor U19236 (N_19236,N_11797,N_11021);
xor U19237 (N_19237,N_12120,N_14661);
or U19238 (N_19238,N_14231,N_10622);
and U19239 (N_19239,N_13803,N_11301);
xor U19240 (N_19240,N_13206,N_14359);
xor U19241 (N_19241,N_14132,N_10822);
nor U19242 (N_19242,N_12652,N_13788);
xor U19243 (N_19243,N_10060,N_13499);
or U19244 (N_19244,N_10886,N_11376);
xor U19245 (N_19245,N_13780,N_14198);
nand U19246 (N_19246,N_12792,N_11280);
xnor U19247 (N_19247,N_13633,N_10169);
or U19248 (N_19248,N_10577,N_10288);
nand U19249 (N_19249,N_10458,N_10390);
nand U19250 (N_19250,N_13867,N_12569);
or U19251 (N_19251,N_13679,N_10217);
and U19252 (N_19252,N_13704,N_10281);
xor U19253 (N_19253,N_13178,N_13318);
nor U19254 (N_19254,N_14852,N_11292);
nand U19255 (N_19255,N_10876,N_11195);
nand U19256 (N_19256,N_14896,N_10563);
and U19257 (N_19257,N_10153,N_10786);
nand U19258 (N_19258,N_12771,N_12485);
or U19259 (N_19259,N_14663,N_14046);
xor U19260 (N_19260,N_13667,N_14979);
xor U19261 (N_19261,N_12906,N_14332);
nor U19262 (N_19262,N_10216,N_13780);
and U19263 (N_19263,N_13113,N_13017);
nor U19264 (N_19264,N_12111,N_12602);
nor U19265 (N_19265,N_13773,N_11823);
or U19266 (N_19266,N_13302,N_10351);
xor U19267 (N_19267,N_13016,N_10390);
nand U19268 (N_19268,N_10794,N_11230);
and U19269 (N_19269,N_14176,N_13813);
nor U19270 (N_19270,N_10099,N_11931);
nand U19271 (N_19271,N_10346,N_11746);
or U19272 (N_19272,N_11357,N_11021);
or U19273 (N_19273,N_10777,N_14698);
or U19274 (N_19274,N_11187,N_10392);
nor U19275 (N_19275,N_11228,N_12263);
nor U19276 (N_19276,N_12781,N_14925);
xor U19277 (N_19277,N_13363,N_12431);
xnor U19278 (N_19278,N_13183,N_12643);
or U19279 (N_19279,N_12391,N_11413);
and U19280 (N_19280,N_12949,N_11786);
nand U19281 (N_19281,N_14440,N_11623);
and U19282 (N_19282,N_13425,N_14871);
or U19283 (N_19283,N_12902,N_13811);
or U19284 (N_19284,N_14226,N_11604);
or U19285 (N_19285,N_14663,N_12221);
and U19286 (N_19286,N_11194,N_13372);
and U19287 (N_19287,N_14190,N_10624);
xor U19288 (N_19288,N_14265,N_14317);
xnor U19289 (N_19289,N_12536,N_11634);
xor U19290 (N_19290,N_12350,N_14907);
or U19291 (N_19291,N_10362,N_11986);
and U19292 (N_19292,N_10712,N_10187);
xnor U19293 (N_19293,N_14425,N_14731);
and U19294 (N_19294,N_12631,N_10299);
and U19295 (N_19295,N_10017,N_10115);
nand U19296 (N_19296,N_10056,N_14623);
or U19297 (N_19297,N_10625,N_12145);
or U19298 (N_19298,N_10386,N_11159);
xor U19299 (N_19299,N_13271,N_11870);
nand U19300 (N_19300,N_10257,N_11369);
or U19301 (N_19301,N_11503,N_14244);
or U19302 (N_19302,N_14796,N_14031);
or U19303 (N_19303,N_14667,N_11203);
nand U19304 (N_19304,N_12618,N_11754);
xor U19305 (N_19305,N_11827,N_10017);
and U19306 (N_19306,N_13590,N_12723);
xor U19307 (N_19307,N_12000,N_11207);
xor U19308 (N_19308,N_12255,N_14404);
xor U19309 (N_19309,N_12374,N_13932);
nor U19310 (N_19310,N_12381,N_14235);
or U19311 (N_19311,N_12819,N_13207);
or U19312 (N_19312,N_11392,N_14462);
nor U19313 (N_19313,N_11509,N_12206);
or U19314 (N_19314,N_13721,N_14601);
nor U19315 (N_19315,N_14463,N_13105);
nand U19316 (N_19316,N_11331,N_11361);
or U19317 (N_19317,N_13853,N_11504);
xor U19318 (N_19318,N_13985,N_11202);
xor U19319 (N_19319,N_12183,N_10732);
nor U19320 (N_19320,N_12726,N_10745);
nand U19321 (N_19321,N_14578,N_13300);
or U19322 (N_19322,N_14381,N_14726);
and U19323 (N_19323,N_13670,N_11674);
xnor U19324 (N_19324,N_10579,N_14994);
or U19325 (N_19325,N_12310,N_10179);
and U19326 (N_19326,N_11736,N_10682);
or U19327 (N_19327,N_11850,N_14996);
nand U19328 (N_19328,N_14812,N_13741);
and U19329 (N_19329,N_13168,N_14355);
nand U19330 (N_19330,N_11148,N_11546);
xor U19331 (N_19331,N_13686,N_10688);
and U19332 (N_19332,N_14755,N_11340);
or U19333 (N_19333,N_13501,N_13010);
nor U19334 (N_19334,N_11022,N_11668);
nor U19335 (N_19335,N_12868,N_10605);
nor U19336 (N_19336,N_13002,N_12135);
xnor U19337 (N_19337,N_13609,N_14469);
xnor U19338 (N_19338,N_10921,N_12971);
or U19339 (N_19339,N_14544,N_11920);
nand U19340 (N_19340,N_11563,N_14862);
xor U19341 (N_19341,N_10994,N_11112);
nor U19342 (N_19342,N_10541,N_10650);
nor U19343 (N_19343,N_14671,N_12500);
and U19344 (N_19344,N_14820,N_10922);
and U19345 (N_19345,N_11880,N_14149);
or U19346 (N_19346,N_14043,N_13636);
and U19347 (N_19347,N_12514,N_14374);
or U19348 (N_19348,N_14729,N_11039);
nand U19349 (N_19349,N_11191,N_10806);
xnor U19350 (N_19350,N_12620,N_11928);
and U19351 (N_19351,N_13878,N_14844);
and U19352 (N_19352,N_11107,N_10481);
or U19353 (N_19353,N_13565,N_10506);
and U19354 (N_19354,N_13869,N_14516);
nor U19355 (N_19355,N_14295,N_14780);
or U19356 (N_19356,N_11579,N_11645);
and U19357 (N_19357,N_14572,N_10457);
nor U19358 (N_19358,N_14700,N_14499);
nor U19359 (N_19359,N_12213,N_10367);
nor U19360 (N_19360,N_14151,N_10872);
nand U19361 (N_19361,N_11612,N_13337);
nor U19362 (N_19362,N_11971,N_14857);
and U19363 (N_19363,N_13246,N_13541);
nand U19364 (N_19364,N_12917,N_14765);
or U19365 (N_19365,N_14793,N_13835);
nand U19366 (N_19366,N_12069,N_11786);
xor U19367 (N_19367,N_10896,N_12240);
nand U19368 (N_19368,N_12368,N_12515);
xor U19369 (N_19369,N_14978,N_14972);
xor U19370 (N_19370,N_14378,N_11681);
or U19371 (N_19371,N_11003,N_10753);
xnor U19372 (N_19372,N_14489,N_13013);
nor U19373 (N_19373,N_10336,N_14928);
nor U19374 (N_19374,N_12282,N_12909);
or U19375 (N_19375,N_10208,N_13217);
nand U19376 (N_19376,N_13826,N_14179);
or U19377 (N_19377,N_11829,N_14041);
nand U19378 (N_19378,N_11637,N_12751);
and U19379 (N_19379,N_10350,N_11024);
xor U19380 (N_19380,N_11942,N_14305);
xor U19381 (N_19381,N_12227,N_11751);
xor U19382 (N_19382,N_10418,N_14029);
nor U19383 (N_19383,N_11754,N_11847);
nor U19384 (N_19384,N_10976,N_11233);
nand U19385 (N_19385,N_14732,N_10469);
or U19386 (N_19386,N_12690,N_11356);
or U19387 (N_19387,N_11682,N_12631);
xnor U19388 (N_19388,N_14170,N_11035);
and U19389 (N_19389,N_10888,N_13256);
nand U19390 (N_19390,N_10841,N_10153);
xor U19391 (N_19391,N_10422,N_12683);
nor U19392 (N_19392,N_14589,N_13941);
xor U19393 (N_19393,N_12522,N_11907);
or U19394 (N_19394,N_13516,N_12278);
nand U19395 (N_19395,N_13078,N_12066);
or U19396 (N_19396,N_12623,N_14143);
nor U19397 (N_19397,N_11364,N_11043);
or U19398 (N_19398,N_12175,N_12517);
nor U19399 (N_19399,N_13577,N_10642);
or U19400 (N_19400,N_13747,N_13494);
xor U19401 (N_19401,N_12631,N_14916);
and U19402 (N_19402,N_14962,N_12235);
or U19403 (N_19403,N_13340,N_10991);
nand U19404 (N_19404,N_11812,N_10561);
or U19405 (N_19405,N_12917,N_13322);
xnor U19406 (N_19406,N_11007,N_10317);
or U19407 (N_19407,N_10956,N_13673);
xor U19408 (N_19408,N_14400,N_14759);
xor U19409 (N_19409,N_13553,N_12271);
nor U19410 (N_19410,N_11259,N_14285);
nand U19411 (N_19411,N_14500,N_13798);
nand U19412 (N_19412,N_10730,N_10374);
or U19413 (N_19413,N_10834,N_12863);
and U19414 (N_19414,N_12871,N_10179);
or U19415 (N_19415,N_10951,N_11140);
and U19416 (N_19416,N_12119,N_13692);
or U19417 (N_19417,N_11817,N_11007);
xor U19418 (N_19418,N_12662,N_12942);
or U19419 (N_19419,N_11320,N_11444);
nand U19420 (N_19420,N_10748,N_13080);
or U19421 (N_19421,N_13873,N_11525);
nor U19422 (N_19422,N_13709,N_14406);
xnor U19423 (N_19423,N_13480,N_12326);
nor U19424 (N_19424,N_14626,N_11470);
and U19425 (N_19425,N_14483,N_13002);
or U19426 (N_19426,N_10060,N_14408);
xor U19427 (N_19427,N_10139,N_12668);
or U19428 (N_19428,N_13881,N_11980);
xnor U19429 (N_19429,N_10354,N_10319);
and U19430 (N_19430,N_13322,N_11127);
nand U19431 (N_19431,N_13432,N_10216);
nand U19432 (N_19432,N_14824,N_12737);
and U19433 (N_19433,N_12388,N_12528);
xnor U19434 (N_19434,N_10787,N_11004);
xor U19435 (N_19435,N_11990,N_12511);
nor U19436 (N_19436,N_10617,N_12676);
or U19437 (N_19437,N_14315,N_11988);
and U19438 (N_19438,N_14570,N_14580);
nand U19439 (N_19439,N_14263,N_13609);
xnor U19440 (N_19440,N_14581,N_11234);
nor U19441 (N_19441,N_10476,N_11540);
or U19442 (N_19442,N_10618,N_11756);
nor U19443 (N_19443,N_11984,N_12502);
nand U19444 (N_19444,N_10214,N_10213);
or U19445 (N_19445,N_13778,N_10173);
xnor U19446 (N_19446,N_13364,N_14975);
nor U19447 (N_19447,N_11120,N_12890);
nand U19448 (N_19448,N_12547,N_12525);
xor U19449 (N_19449,N_10919,N_14904);
or U19450 (N_19450,N_10817,N_13593);
xor U19451 (N_19451,N_14759,N_12657);
xnor U19452 (N_19452,N_12428,N_11742);
nor U19453 (N_19453,N_11226,N_11803);
nand U19454 (N_19454,N_13412,N_10139);
and U19455 (N_19455,N_13794,N_10890);
xor U19456 (N_19456,N_12586,N_10084);
or U19457 (N_19457,N_12950,N_12118);
nor U19458 (N_19458,N_12009,N_11082);
or U19459 (N_19459,N_14440,N_11852);
and U19460 (N_19460,N_10144,N_13547);
nand U19461 (N_19461,N_13230,N_10575);
xor U19462 (N_19462,N_13221,N_13169);
and U19463 (N_19463,N_12606,N_12745);
xnor U19464 (N_19464,N_13401,N_10135);
nand U19465 (N_19465,N_13414,N_11184);
or U19466 (N_19466,N_13110,N_10354);
nor U19467 (N_19467,N_12391,N_11072);
nor U19468 (N_19468,N_10787,N_13676);
and U19469 (N_19469,N_12569,N_10760);
nor U19470 (N_19470,N_13582,N_14899);
or U19471 (N_19471,N_11562,N_13233);
nor U19472 (N_19472,N_13910,N_10219);
or U19473 (N_19473,N_11781,N_13127);
xor U19474 (N_19474,N_14158,N_14337);
nand U19475 (N_19475,N_11152,N_13602);
or U19476 (N_19476,N_13116,N_14932);
or U19477 (N_19477,N_10801,N_14951);
or U19478 (N_19478,N_11132,N_10086);
nor U19479 (N_19479,N_14189,N_13826);
xnor U19480 (N_19480,N_11486,N_11330);
and U19481 (N_19481,N_12862,N_12047);
and U19482 (N_19482,N_14444,N_10865);
xnor U19483 (N_19483,N_10552,N_10081);
nor U19484 (N_19484,N_10715,N_11901);
nor U19485 (N_19485,N_14753,N_14169);
or U19486 (N_19486,N_10830,N_10114);
and U19487 (N_19487,N_13411,N_10710);
nand U19488 (N_19488,N_11366,N_10936);
nor U19489 (N_19489,N_10648,N_14739);
or U19490 (N_19490,N_13159,N_14505);
or U19491 (N_19491,N_12520,N_14674);
xnor U19492 (N_19492,N_14201,N_14644);
and U19493 (N_19493,N_11880,N_14501);
nand U19494 (N_19494,N_11341,N_13489);
nand U19495 (N_19495,N_12673,N_13485);
nand U19496 (N_19496,N_13385,N_11795);
and U19497 (N_19497,N_11946,N_13890);
or U19498 (N_19498,N_14857,N_13428);
or U19499 (N_19499,N_10925,N_10729);
nand U19500 (N_19500,N_13476,N_12588);
nor U19501 (N_19501,N_11063,N_13745);
xnor U19502 (N_19502,N_12608,N_13345);
and U19503 (N_19503,N_14504,N_14607);
nor U19504 (N_19504,N_13931,N_14731);
xnor U19505 (N_19505,N_11141,N_13279);
nand U19506 (N_19506,N_10420,N_11782);
nor U19507 (N_19507,N_11207,N_11362);
nand U19508 (N_19508,N_10299,N_11166);
xnor U19509 (N_19509,N_13832,N_14703);
or U19510 (N_19510,N_11605,N_10935);
nand U19511 (N_19511,N_12727,N_10185);
nand U19512 (N_19512,N_14072,N_14835);
xor U19513 (N_19513,N_14520,N_11990);
nor U19514 (N_19514,N_14931,N_11143);
or U19515 (N_19515,N_13762,N_12031);
or U19516 (N_19516,N_12899,N_11709);
or U19517 (N_19517,N_10552,N_12701);
xor U19518 (N_19518,N_13141,N_12887);
or U19519 (N_19519,N_13367,N_10228);
nand U19520 (N_19520,N_12315,N_11988);
and U19521 (N_19521,N_14550,N_12862);
or U19522 (N_19522,N_13008,N_10518);
or U19523 (N_19523,N_12800,N_12160);
or U19524 (N_19524,N_10463,N_13336);
nand U19525 (N_19525,N_14945,N_12010);
nand U19526 (N_19526,N_10632,N_12301);
nor U19527 (N_19527,N_14637,N_11870);
or U19528 (N_19528,N_14122,N_10150);
nor U19529 (N_19529,N_12566,N_12585);
xnor U19530 (N_19530,N_14300,N_12683);
xnor U19531 (N_19531,N_13582,N_12132);
nand U19532 (N_19532,N_11413,N_14311);
xor U19533 (N_19533,N_12259,N_14510);
xor U19534 (N_19534,N_10693,N_14996);
or U19535 (N_19535,N_11285,N_13497);
or U19536 (N_19536,N_12087,N_10010);
or U19537 (N_19537,N_13068,N_11022);
nand U19538 (N_19538,N_11491,N_12606);
nor U19539 (N_19539,N_14807,N_11528);
or U19540 (N_19540,N_12547,N_14227);
nor U19541 (N_19541,N_12636,N_12178);
nand U19542 (N_19542,N_10625,N_13978);
or U19543 (N_19543,N_14882,N_13088);
nor U19544 (N_19544,N_13021,N_11219);
xor U19545 (N_19545,N_14535,N_10668);
or U19546 (N_19546,N_12422,N_10148);
nand U19547 (N_19547,N_11780,N_13805);
nor U19548 (N_19548,N_10576,N_12533);
xor U19549 (N_19549,N_11912,N_14794);
or U19550 (N_19550,N_12614,N_11656);
or U19551 (N_19551,N_11304,N_10222);
nand U19552 (N_19552,N_12725,N_13278);
and U19553 (N_19553,N_11537,N_11000);
nand U19554 (N_19554,N_11859,N_13885);
nand U19555 (N_19555,N_10013,N_13663);
or U19556 (N_19556,N_14718,N_12115);
nor U19557 (N_19557,N_11773,N_11926);
nor U19558 (N_19558,N_14077,N_12826);
xnor U19559 (N_19559,N_11096,N_14263);
xnor U19560 (N_19560,N_10682,N_11439);
nor U19561 (N_19561,N_11371,N_13048);
xor U19562 (N_19562,N_12702,N_11691);
or U19563 (N_19563,N_10215,N_14351);
or U19564 (N_19564,N_10699,N_13149);
xnor U19565 (N_19565,N_12709,N_12353);
xnor U19566 (N_19566,N_11498,N_11122);
nand U19567 (N_19567,N_11409,N_10874);
or U19568 (N_19568,N_14007,N_12433);
nand U19569 (N_19569,N_13316,N_11134);
and U19570 (N_19570,N_13618,N_12260);
and U19571 (N_19571,N_10531,N_10840);
or U19572 (N_19572,N_13762,N_14309);
nand U19573 (N_19573,N_11338,N_14412);
or U19574 (N_19574,N_12569,N_11207);
and U19575 (N_19575,N_10052,N_10871);
nor U19576 (N_19576,N_12576,N_11205);
nor U19577 (N_19577,N_11906,N_14972);
xnor U19578 (N_19578,N_10755,N_13419);
nor U19579 (N_19579,N_12735,N_12908);
nor U19580 (N_19580,N_12547,N_10638);
nand U19581 (N_19581,N_12300,N_14252);
and U19582 (N_19582,N_13371,N_10735);
or U19583 (N_19583,N_11652,N_14116);
nor U19584 (N_19584,N_14488,N_11888);
nand U19585 (N_19585,N_12789,N_12311);
nand U19586 (N_19586,N_13779,N_11054);
and U19587 (N_19587,N_14534,N_11292);
nor U19588 (N_19588,N_13684,N_13460);
nand U19589 (N_19589,N_13027,N_12573);
nand U19590 (N_19590,N_14823,N_10643);
nor U19591 (N_19591,N_14929,N_12062);
and U19592 (N_19592,N_14381,N_14130);
nor U19593 (N_19593,N_11122,N_10631);
xnor U19594 (N_19594,N_10739,N_11054);
nand U19595 (N_19595,N_14521,N_10714);
or U19596 (N_19596,N_14856,N_10624);
nor U19597 (N_19597,N_13359,N_13026);
and U19598 (N_19598,N_13087,N_14714);
or U19599 (N_19599,N_10493,N_12524);
xnor U19600 (N_19600,N_12071,N_10085);
nor U19601 (N_19601,N_12619,N_11249);
xor U19602 (N_19602,N_11787,N_12757);
xor U19603 (N_19603,N_14962,N_10816);
xor U19604 (N_19604,N_14146,N_13562);
or U19605 (N_19605,N_11524,N_13541);
nor U19606 (N_19606,N_10642,N_12182);
xnor U19607 (N_19607,N_14314,N_13100);
xnor U19608 (N_19608,N_11574,N_10524);
nor U19609 (N_19609,N_14891,N_12738);
nand U19610 (N_19610,N_14447,N_14351);
xnor U19611 (N_19611,N_12325,N_13831);
and U19612 (N_19612,N_12266,N_11459);
or U19613 (N_19613,N_14878,N_12959);
and U19614 (N_19614,N_14124,N_13654);
xor U19615 (N_19615,N_10342,N_12529);
nand U19616 (N_19616,N_13558,N_10860);
and U19617 (N_19617,N_11841,N_10324);
and U19618 (N_19618,N_13844,N_12219);
and U19619 (N_19619,N_10494,N_10598);
xnor U19620 (N_19620,N_13682,N_11726);
xnor U19621 (N_19621,N_11722,N_13104);
and U19622 (N_19622,N_11971,N_12848);
xnor U19623 (N_19623,N_10297,N_12360);
and U19624 (N_19624,N_12242,N_13837);
xor U19625 (N_19625,N_12028,N_12076);
and U19626 (N_19626,N_11962,N_11311);
xnor U19627 (N_19627,N_13932,N_12115);
xnor U19628 (N_19628,N_10028,N_13522);
or U19629 (N_19629,N_10328,N_13176);
nor U19630 (N_19630,N_12783,N_11565);
or U19631 (N_19631,N_12895,N_10460);
nor U19632 (N_19632,N_11880,N_13986);
nor U19633 (N_19633,N_13604,N_13498);
and U19634 (N_19634,N_11276,N_12058);
and U19635 (N_19635,N_10300,N_14414);
or U19636 (N_19636,N_10745,N_14225);
nand U19637 (N_19637,N_14626,N_10387);
nor U19638 (N_19638,N_14088,N_10934);
nor U19639 (N_19639,N_13941,N_12841);
nand U19640 (N_19640,N_13338,N_13231);
and U19641 (N_19641,N_14380,N_10609);
nor U19642 (N_19642,N_11597,N_13578);
or U19643 (N_19643,N_10655,N_10991);
nand U19644 (N_19644,N_10343,N_13476);
nor U19645 (N_19645,N_10379,N_11875);
or U19646 (N_19646,N_11974,N_12853);
or U19647 (N_19647,N_14547,N_12522);
nor U19648 (N_19648,N_14634,N_12726);
or U19649 (N_19649,N_10419,N_11375);
nand U19650 (N_19650,N_12322,N_12006);
nand U19651 (N_19651,N_12244,N_10526);
and U19652 (N_19652,N_12854,N_13895);
and U19653 (N_19653,N_13562,N_13199);
nand U19654 (N_19654,N_13461,N_14499);
xor U19655 (N_19655,N_11630,N_11504);
nor U19656 (N_19656,N_12994,N_10613);
and U19657 (N_19657,N_11083,N_14951);
or U19658 (N_19658,N_14468,N_14463);
and U19659 (N_19659,N_14733,N_14242);
or U19660 (N_19660,N_10750,N_10858);
or U19661 (N_19661,N_11358,N_10793);
or U19662 (N_19662,N_10064,N_14969);
nand U19663 (N_19663,N_10141,N_13419);
xnor U19664 (N_19664,N_13297,N_10648);
and U19665 (N_19665,N_14531,N_14167);
nand U19666 (N_19666,N_11643,N_11978);
and U19667 (N_19667,N_11457,N_14342);
nor U19668 (N_19668,N_10709,N_13335);
xnor U19669 (N_19669,N_10730,N_14397);
xnor U19670 (N_19670,N_10566,N_11985);
and U19671 (N_19671,N_12997,N_12696);
nor U19672 (N_19672,N_12838,N_14566);
or U19673 (N_19673,N_13623,N_14145);
and U19674 (N_19674,N_11043,N_14650);
xnor U19675 (N_19675,N_10036,N_11527);
nand U19676 (N_19676,N_12464,N_13290);
xnor U19677 (N_19677,N_12887,N_10450);
and U19678 (N_19678,N_12272,N_13650);
xor U19679 (N_19679,N_11597,N_10407);
or U19680 (N_19680,N_11239,N_12920);
nand U19681 (N_19681,N_10718,N_13340);
or U19682 (N_19682,N_10832,N_10550);
xor U19683 (N_19683,N_13331,N_10433);
xor U19684 (N_19684,N_12569,N_13007);
and U19685 (N_19685,N_10238,N_13501);
nor U19686 (N_19686,N_14974,N_13420);
nor U19687 (N_19687,N_11179,N_14141);
xor U19688 (N_19688,N_11449,N_12975);
nand U19689 (N_19689,N_13619,N_11624);
nand U19690 (N_19690,N_10742,N_10174);
and U19691 (N_19691,N_13566,N_13003);
and U19692 (N_19692,N_10217,N_10809);
nand U19693 (N_19693,N_10332,N_13291);
nor U19694 (N_19694,N_14295,N_13026);
or U19695 (N_19695,N_11580,N_10940);
nor U19696 (N_19696,N_11099,N_14765);
nand U19697 (N_19697,N_10292,N_10682);
nor U19698 (N_19698,N_13485,N_10880);
xor U19699 (N_19699,N_13859,N_12195);
xor U19700 (N_19700,N_12952,N_14158);
and U19701 (N_19701,N_10237,N_14204);
nand U19702 (N_19702,N_10467,N_11020);
nor U19703 (N_19703,N_10976,N_14764);
nand U19704 (N_19704,N_13977,N_12609);
nand U19705 (N_19705,N_10787,N_10054);
or U19706 (N_19706,N_12749,N_12568);
nor U19707 (N_19707,N_12615,N_14654);
xnor U19708 (N_19708,N_14185,N_11781);
and U19709 (N_19709,N_12394,N_10960);
or U19710 (N_19710,N_11694,N_13351);
xor U19711 (N_19711,N_13571,N_13992);
nand U19712 (N_19712,N_11669,N_13770);
nand U19713 (N_19713,N_11486,N_13743);
nor U19714 (N_19714,N_12499,N_14167);
or U19715 (N_19715,N_11413,N_11376);
nand U19716 (N_19716,N_13251,N_13439);
nor U19717 (N_19717,N_10768,N_11061);
or U19718 (N_19718,N_11955,N_13663);
nor U19719 (N_19719,N_12723,N_12965);
xor U19720 (N_19720,N_14708,N_10955);
or U19721 (N_19721,N_11523,N_11270);
xor U19722 (N_19722,N_10036,N_11431);
or U19723 (N_19723,N_13039,N_12896);
nor U19724 (N_19724,N_11163,N_14777);
nand U19725 (N_19725,N_13867,N_11060);
nor U19726 (N_19726,N_12687,N_12889);
nor U19727 (N_19727,N_14417,N_13323);
nor U19728 (N_19728,N_13448,N_14123);
xor U19729 (N_19729,N_13764,N_10590);
xnor U19730 (N_19730,N_12124,N_12530);
or U19731 (N_19731,N_12310,N_14951);
xnor U19732 (N_19732,N_11227,N_12321);
xnor U19733 (N_19733,N_14670,N_10148);
and U19734 (N_19734,N_13780,N_11583);
xor U19735 (N_19735,N_10212,N_14951);
nor U19736 (N_19736,N_12562,N_13047);
xor U19737 (N_19737,N_11745,N_12372);
or U19738 (N_19738,N_12079,N_12836);
nor U19739 (N_19739,N_10689,N_11393);
nor U19740 (N_19740,N_13414,N_11515);
and U19741 (N_19741,N_14860,N_12706);
or U19742 (N_19742,N_11250,N_13552);
nand U19743 (N_19743,N_14294,N_14952);
nand U19744 (N_19744,N_13393,N_10834);
nor U19745 (N_19745,N_14145,N_10668);
nor U19746 (N_19746,N_11383,N_12769);
xnor U19747 (N_19747,N_10596,N_14691);
or U19748 (N_19748,N_14508,N_10216);
or U19749 (N_19749,N_13989,N_14665);
xnor U19750 (N_19750,N_11093,N_13388);
xor U19751 (N_19751,N_12208,N_12309);
xor U19752 (N_19752,N_11126,N_10182);
nand U19753 (N_19753,N_10707,N_14119);
or U19754 (N_19754,N_10011,N_12589);
xnor U19755 (N_19755,N_13457,N_11238);
or U19756 (N_19756,N_12567,N_10807);
nor U19757 (N_19757,N_14242,N_14586);
or U19758 (N_19758,N_13130,N_11239);
and U19759 (N_19759,N_14758,N_13288);
or U19760 (N_19760,N_10232,N_13386);
and U19761 (N_19761,N_11906,N_10747);
nand U19762 (N_19762,N_10286,N_13861);
or U19763 (N_19763,N_14687,N_11760);
nand U19764 (N_19764,N_12497,N_10099);
nor U19765 (N_19765,N_14250,N_10138);
and U19766 (N_19766,N_10298,N_13031);
and U19767 (N_19767,N_10786,N_12352);
nor U19768 (N_19768,N_12755,N_10804);
xnor U19769 (N_19769,N_10694,N_12223);
xnor U19770 (N_19770,N_14962,N_12869);
or U19771 (N_19771,N_10652,N_10081);
and U19772 (N_19772,N_10946,N_13317);
xnor U19773 (N_19773,N_11931,N_13343);
nand U19774 (N_19774,N_10845,N_10617);
or U19775 (N_19775,N_13871,N_13552);
and U19776 (N_19776,N_10792,N_11826);
or U19777 (N_19777,N_10818,N_12249);
or U19778 (N_19778,N_13561,N_10899);
nor U19779 (N_19779,N_14182,N_10274);
nor U19780 (N_19780,N_13018,N_12360);
and U19781 (N_19781,N_13625,N_13560);
nor U19782 (N_19782,N_11370,N_12074);
and U19783 (N_19783,N_11733,N_12377);
nand U19784 (N_19784,N_12061,N_14517);
and U19785 (N_19785,N_13226,N_12035);
and U19786 (N_19786,N_12531,N_14531);
and U19787 (N_19787,N_11373,N_11717);
or U19788 (N_19788,N_14273,N_14633);
nor U19789 (N_19789,N_11446,N_13674);
nand U19790 (N_19790,N_10754,N_10404);
or U19791 (N_19791,N_10160,N_14309);
nand U19792 (N_19792,N_11889,N_11053);
xnor U19793 (N_19793,N_14005,N_13847);
and U19794 (N_19794,N_14570,N_10640);
or U19795 (N_19795,N_12655,N_14322);
and U19796 (N_19796,N_10608,N_10825);
or U19797 (N_19797,N_10335,N_10309);
or U19798 (N_19798,N_14468,N_14046);
or U19799 (N_19799,N_13534,N_12672);
and U19800 (N_19800,N_13309,N_14221);
xor U19801 (N_19801,N_13730,N_11408);
xor U19802 (N_19802,N_10867,N_13345);
xor U19803 (N_19803,N_10303,N_14821);
or U19804 (N_19804,N_11993,N_11774);
nor U19805 (N_19805,N_14872,N_13547);
nand U19806 (N_19806,N_10592,N_11352);
and U19807 (N_19807,N_14172,N_14373);
nor U19808 (N_19808,N_12084,N_13231);
nor U19809 (N_19809,N_12662,N_10706);
and U19810 (N_19810,N_12448,N_10383);
xnor U19811 (N_19811,N_11811,N_13746);
and U19812 (N_19812,N_10299,N_13754);
xor U19813 (N_19813,N_11491,N_14369);
or U19814 (N_19814,N_10552,N_11764);
or U19815 (N_19815,N_13764,N_12621);
or U19816 (N_19816,N_11443,N_12294);
nand U19817 (N_19817,N_10394,N_12512);
and U19818 (N_19818,N_10472,N_10445);
nand U19819 (N_19819,N_11633,N_14839);
and U19820 (N_19820,N_10545,N_13749);
nand U19821 (N_19821,N_10754,N_12168);
and U19822 (N_19822,N_12730,N_12316);
and U19823 (N_19823,N_12753,N_10177);
or U19824 (N_19824,N_12066,N_12824);
xnor U19825 (N_19825,N_14156,N_11655);
nand U19826 (N_19826,N_12809,N_10258);
and U19827 (N_19827,N_10034,N_13501);
nor U19828 (N_19828,N_13116,N_14073);
nor U19829 (N_19829,N_12293,N_11209);
nand U19830 (N_19830,N_13278,N_12465);
nor U19831 (N_19831,N_13602,N_12346);
and U19832 (N_19832,N_13074,N_14004);
or U19833 (N_19833,N_11738,N_10671);
and U19834 (N_19834,N_13087,N_13252);
nor U19835 (N_19835,N_12190,N_11580);
nand U19836 (N_19836,N_14522,N_12813);
xnor U19837 (N_19837,N_13716,N_10958);
nor U19838 (N_19838,N_14316,N_13369);
and U19839 (N_19839,N_10473,N_14404);
nand U19840 (N_19840,N_11916,N_12944);
and U19841 (N_19841,N_11305,N_10329);
xor U19842 (N_19842,N_12254,N_13763);
xnor U19843 (N_19843,N_10127,N_10308);
nand U19844 (N_19844,N_14786,N_10768);
or U19845 (N_19845,N_10225,N_11386);
xor U19846 (N_19846,N_11028,N_12022);
or U19847 (N_19847,N_13004,N_12028);
or U19848 (N_19848,N_11186,N_10501);
and U19849 (N_19849,N_10257,N_12875);
or U19850 (N_19850,N_11756,N_13536);
nor U19851 (N_19851,N_14781,N_11793);
xnor U19852 (N_19852,N_14810,N_14198);
nand U19853 (N_19853,N_14543,N_13884);
and U19854 (N_19854,N_13969,N_14754);
or U19855 (N_19855,N_10807,N_13646);
and U19856 (N_19856,N_10872,N_14982);
nor U19857 (N_19857,N_10918,N_10220);
xnor U19858 (N_19858,N_12375,N_13549);
nor U19859 (N_19859,N_10266,N_14050);
and U19860 (N_19860,N_10495,N_12040);
nand U19861 (N_19861,N_12384,N_11155);
xnor U19862 (N_19862,N_14892,N_10800);
nand U19863 (N_19863,N_10252,N_10702);
xnor U19864 (N_19864,N_11071,N_13837);
and U19865 (N_19865,N_11593,N_12830);
nor U19866 (N_19866,N_13569,N_11383);
and U19867 (N_19867,N_13278,N_11871);
and U19868 (N_19868,N_10185,N_12756);
or U19869 (N_19869,N_11592,N_13090);
nor U19870 (N_19870,N_10417,N_12285);
xnor U19871 (N_19871,N_14079,N_12103);
and U19872 (N_19872,N_10900,N_10241);
or U19873 (N_19873,N_12695,N_10508);
or U19874 (N_19874,N_12783,N_14467);
xor U19875 (N_19875,N_10066,N_11840);
and U19876 (N_19876,N_13740,N_10086);
nand U19877 (N_19877,N_14184,N_11787);
or U19878 (N_19878,N_11744,N_14299);
xor U19879 (N_19879,N_12122,N_12742);
or U19880 (N_19880,N_13288,N_11171);
or U19881 (N_19881,N_13750,N_12829);
nand U19882 (N_19882,N_10322,N_11882);
nand U19883 (N_19883,N_11510,N_11031);
nor U19884 (N_19884,N_12162,N_11850);
nor U19885 (N_19885,N_13280,N_12793);
nor U19886 (N_19886,N_10901,N_10962);
nor U19887 (N_19887,N_13094,N_11167);
and U19888 (N_19888,N_11264,N_11537);
or U19889 (N_19889,N_14252,N_13156);
and U19890 (N_19890,N_13787,N_12867);
and U19891 (N_19891,N_11936,N_14382);
xor U19892 (N_19892,N_12487,N_13704);
nor U19893 (N_19893,N_11145,N_10671);
nor U19894 (N_19894,N_11034,N_12330);
xor U19895 (N_19895,N_11972,N_11824);
xnor U19896 (N_19896,N_11211,N_12988);
nand U19897 (N_19897,N_10077,N_12449);
and U19898 (N_19898,N_10577,N_12384);
nor U19899 (N_19899,N_14407,N_14756);
nand U19900 (N_19900,N_13639,N_13769);
nor U19901 (N_19901,N_11473,N_13487);
nand U19902 (N_19902,N_13861,N_13929);
xnor U19903 (N_19903,N_13075,N_13626);
nand U19904 (N_19904,N_13099,N_13687);
and U19905 (N_19905,N_14724,N_12922);
and U19906 (N_19906,N_12570,N_13955);
or U19907 (N_19907,N_11253,N_13048);
xnor U19908 (N_19908,N_12457,N_13562);
or U19909 (N_19909,N_13625,N_12446);
or U19910 (N_19910,N_10996,N_10356);
and U19911 (N_19911,N_11658,N_10443);
and U19912 (N_19912,N_13903,N_13608);
and U19913 (N_19913,N_11977,N_10903);
xnor U19914 (N_19914,N_11439,N_10381);
nand U19915 (N_19915,N_10097,N_13886);
and U19916 (N_19916,N_10347,N_12836);
nand U19917 (N_19917,N_14890,N_14130);
nand U19918 (N_19918,N_13397,N_13356);
nor U19919 (N_19919,N_13432,N_11874);
and U19920 (N_19920,N_14037,N_10156);
and U19921 (N_19921,N_13934,N_11396);
nand U19922 (N_19922,N_10003,N_11573);
nand U19923 (N_19923,N_13920,N_11004);
xor U19924 (N_19924,N_12707,N_11284);
nand U19925 (N_19925,N_13762,N_11345);
nor U19926 (N_19926,N_12320,N_10702);
nand U19927 (N_19927,N_14104,N_14721);
xnor U19928 (N_19928,N_13948,N_12092);
xor U19929 (N_19929,N_12846,N_10525);
and U19930 (N_19930,N_14783,N_13802);
or U19931 (N_19931,N_13245,N_12734);
or U19932 (N_19932,N_10064,N_13700);
and U19933 (N_19933,N_13688,N_12716);
nand U19934 (N_19934,N_13097,N_14929);
xnor U19935 (N_19935,N_14657,N_10871);
or U19936 (N_19936,N_14510,N_13822);
nand U19937 (N_19937,N_10722,N_12067);
nor U19938 (N_19938,N_12350,N_10996);
xnor U19939 (N_19939,N_10328,N_12548);
or U19940 (N_19940,N_14171,N_14814);
nand U19941 (N_19941,N_10106,N_13864);
xnor U19942 (N_19942,N_10913,N_12694);
or U19943 (N_19943,N_12714,N_14606);
xnor U19944 (N_19944,N_13847,N_11119);
and U19945 (N_19945,N_12947,N_10719);
nor U19946 (N_19946,N_12239,N_10918);
or U19947 (N_19947,N_11369,N_13800);
xor U19948 (N_19948,N_12876,N_10099);
nand U19949 (N_19949,N_11291,N_11678);
and U19950 (N_19950,N_11749,N_13107);
nand U19951 (N_19951,N_10000,N_14192);
or U19952 (N_19952,N_13373,N_14290);
or U19953 (N_19953,N_10154,N_13644);
or U19954 (N_19954,N_10376,N_14119);
xnor U19955 (N_19955,N_12069,N_12347);
xor U19956 (N_19956,N_11947,N_10466);
and U19957 (N_19957,N_14117,N_13429);
xnor U19958 (N_19958,N_12259,N_10046);
and U19959 (N_19959,N_11090,N_14774);
xnor U19960 (N_19960,N_10643,N_13152);
nand U19961 (N_19961,N_12749,N_13968);
nand U19962 (N_19962,N_13126,N_14983);
nor U19963 (N_19963,N_10675,N_10338);
nand U19964 (N_19964,N_11023,N_11678);
and U19965 (N_19965,N_13281,N_13472);
nand U19966 (N_19966,N_14970,N_11466);
and U19967 (N_19967,N_12955,N_10558);
xnor U19968 (N_19968,N_11123,N_13866);
xnor U19969 (N_19969,N_12607,N_13823);
xnor U19970 (N_19970,N_12323,N_12982);
and U19971 (N_19971,N_10461,N_11025);
xnor U19972 (N_19972,N_11491,N_13347);
nand U19973 (N_19973,N_11628,N_13901);
or U19974 (N_19974,N_12476,N_13104);
or U19975 (N_19975,N_11222,N_11334);
or U19976 (N_19976,N_14651,N_13448);
xor U19977 (N_19977,N_11688,N_13648);
or U19978 (N_19978,N_10001,N_13897);
xor U19979 (N_19979,N_11667,N_12343);
or U19980 (N_19980,N_11442,N_11437);
or U19981 (N_19981,N_10338,N_10944);
xor U19982 (N_19982,N_14675,N_12438);
nand U19983 (N_19983,N_11988,N_10462);
nand U19984 (N_19984,N_12038,N_14982);
xor U19985 (N_19985,N_10640,N_10244);
and U19986 (N_19986,N_14528,N_12512);
xor U19987 (N_19987,N_11660,N_10226);
nor U19988 (N_19988,N_12967,N_14119);
nand U19989 (N_19989,N_14795,N_13301);
and U19990 (N_19990,N_13578,N_12295);
xnor U19991 (N_19991,N_11240,N_12744);
or U19992 (N_19992,N_11572,N_10923);
and U19993 (N_19993,N_12649,N_11002);
or U19994 (N_19994,N_12871,N_13578);
nor U19995 (N_19995,N_12887,N_12137);
nor U19996 (N_19996,N_11242,N_14645);
or U19997 (N_19997,N_14910,N_14656);
and U19998 (N_19998,N_10867,N_11683);
or U19999 (N_19999,N_12902,N_11271);
or U20000 (N_20000,N_19789,N_15547);
and U20001 (N_20001,N_16285,N_19764);
xnor U20002 (N_20002,N_15068,N_15165);
nand U20003 (N_20003,N_19360,N_18953);
or U20004 (N_20004,N_18960,N_18510);
nor U20005 (N_20005,N_19774,N_18162);
nand U20006 (N_20006,N_17959,N_15836);
and U20007 (N_20007,N_19129,N_19077);
nor U20008 (N_20008,N_18441,N_15881);
or U20009 (N_20009,N_16517,N_16498);
nor U20010 (N_20010,N_15059,N_15768);
nand U20011 (N_20011,N_18939,N_19311);
and U20012 (N_20012,N_16495,N_18318);
and U20013 (N_20013,N_17515,N_16863);
or U20014 (N_20014,N_16243,N_18155);
xnor U20015 (N_20015,N_16166,N_19771);
nor U20016 (N_20016,N_19744,N_16780);
nand U20017 (N_20017,N_17230,N_16855);
and U20018 (N_20018,N_18738,N_18357);
or U20019 (N_20019,N_18726,N_16689);
nor U20020 (N_20020,N_19784,N_16705);
nor U20021 (N_20021,N_15078,N_19341);
xnor U20022 (N_20022,N_18394,N_19811);
and U20023 (N_20023,N_17893,N_16029);
or U20024 (N_20024,N_17155,N_18687);
and U20025 (N_20025,N_16043,N_19816);
and U20026 (N_20026,N_17688,N_15957);
nand U20027 (N_20027,N_17575,N_16991);
or U20028 (N_20028,N_17557,N_16733);
nor U20029 (N_20029,N_16736,N_17775);
nand U20030 (N_20030,N_18782,N_15026);
nand U20031 (N_20031,N_18489,N_15590);
and U20032 (N_20032,N_19932,N_15344);
and U20033 (N_20033,N_15097,N_15446);
nand U20034 (N_20034,N_18376,N_16587);
xnor U20035 (N_20035,N_18134,N_16073);
and U20036 (N_20036,N_19503,N_19794);
or U20037 (N_20037,N_18469,N_17184);
nor U20038 (N_20038,N_16908,N_18429);
or U20039 (N_20039,N_17586,N_16239);
and U20040 (N_20040,N_19069,N_19025);
nand U20041 (N_20041,N_17530,N_19467);
nor U20042 (N_20042,N_16885,N_16819);
nand U20043 (N_20043,N_15003,N_15605);
or U20044 (N_20044,N_15997,N_15618);
and U20045 (N_20045,N_16936,N_15350);
nor U20046 (N_20046,N_16021,N_16115);
nand U20047 (N_20047,N_18360,N_17900);
nor U20048 (N_20048,N_19458,N_16737);
nand U20049 (N_20049,N_16844,N_16135);
and U20050 (N_20050,N_15405,N_17639);
xor U20051 (N_20051,N_19793,N_16762);
xor U20052 (N_20052,N_18600,N_17559);
or U20053 (N_20053,N_15540,N_19185);
xor U20054 (N_20054,N_17000,N_15480);
nor U20055 (N_20055,N_19868,N_18359);
xor U20056 (N_20056,N_19449,N_16236);
xnor U20057 (N_20057,N_18324,N_16169);
xor U20058 (N_20058,N_16856,N_18169);
xnor U20059 (N_20059,N_19248,N_19866);
and U20060 (N_20060,N_18408,N_17408);
and U20061 (N_20061,N_19551,N_18460);
nor U20062 (N_20062,N_17713,N_17794);
xor U20063 (N_20063,N_19756,N_16351);
nor U20064 (N_20064,N_16328,N_18455);
nor U20065 (N_20065,N_16866,N_17704);
xnor U20066 (N_20066,N_15439,N_19713);
and U20067 (N_20067,N_18284,N_18727);
xor U20068 (N_20068,N_15361,N_17881);
or U20069 (N_20069,N_15835,N_17728);
nor U20070 (N_20070,N_19613,N_18185);
and U20071 (N_20071,N_19590,N_16370);
and U20072 (N_20072,N_18728,N_16238);
nand U20073 (N_20073,N_16217,N_15409);
nor U20074 (N_20074,N_18900,N_17897);
nor U20075 (N_20075,N_18666,N_19751);
nand U20076 (N_20076,N_17473,N_15724);
xnor U20077 (N_20077,N_19254,N_15093);
or U20078 (N_20078,N_16375,N_15660);
nand U20079 (N_20079,N_18114,N_15573);
xnor U20080 (N_20080,N_18046,N_16838);
and U20081 (N_20081,N_16261,N_19451);
or U20082 (N_20082,N_18137,N_17654);
nor U20083 (N_20083,N_18299,N_19354);
or U20084 (N_20084,N_18679,N_16099);
or U20085 (N_20085,N_15688,N_17087);
xnor U20086 (N_20086,N_18436,N_19284);
xnor U20087 (N_20087,N_17187,N_18197);
or U20088 (N_20088,N_16227,N_19929);
and U20089 (N_20089,N_17287,N_17004);
and U20090 (N_20090,N_17103,N_16065);
nand U20091 (N_20091,N_16028,N_19967);
nor U20092 (N_20092,N_16276,N_18282);
and U20093 (N_20093,N_17052,N_15232);
xnor U20094 (N_20094,N_19469,N_17203);
nor U20095 (N_20095,N_16961,N_19170);
or U20096 (N_20096,N_17300,N_15918);
nor U20097 (N_20097,N_17862,N_19495);
or U20098 (N_20098,N_17263,N_18451);
or U20099 (N_20099,N_17924,N_19640);
nand U20100 (N_20100,N_15231,N_15914);
xnor U20101 (N_20101,N_17487,N_19285);
nor U20102 (N_20102,N_19265,N_17815);
and U20103 (N_20103,N_15150,N_16155);
and U20104 (N_20104,N_18854,N_18486);
xnor U20105 (N_20105,N_15579,N_15910);
and U20106 (N_20106,N_18266,N_17617);
or U20107 (N_20107,N_16806,N_16684);
nand U20108 (N_20108,N_17420,N_18423);
and U20109 (N_20109,N_19930,N_16042);
nand U20110 (N_20110,N_17185,N_15847);
nor U20111 (N_20111,N_16396,N_16342);
and U20112 (N_20112,N_19050,N_19300);
nand U20113 (N_20113,N_16251,N_16113);
nand U20114 (N_20114,N_15539,N_15456);
nor U20115 (N_20115,N_15025,N_16134);
or U20116 (N_20116,N_17196,N_17268);
xnor U20117 (N_20117,N_19320,N_16272);
nor U20118 (N_20118,N_15017,N_19507);
nand U20119 (N_20119,N_18024,N_19239);
xnor U20120 (N_20120,N_19044,N_19110);
nor U20121 (N_20121,N_16055,N_16526);
or U20122 (N_20122,N_16949,N_17072);
or U20123 (N_20123,N_15512,N_18615);
nand U20124 (N_20124,N_15988,N_18336);
xnor U20125 (N_20125,N_17279,N_17074);
or U20126 (N_20126,N_17429,N_19673);
xnor U20127 (N_20127,N_17751,N_19876);
and U20128 (N_20128,N_16117,N_17086);
xor U20129 (N_20129,N_16761,N_16559);
or U20130 (N_20130,N_15984,N_15535);
and U20131 (N_20131,N_18651,N_15533);
or U20132 (N_20132,N_19679,N_15657);
nor U20133 (N_20133,N_18287,N_19849);
nand U20134 (N_20134,N_18109,N_19213);
xor U20135 (N_20135,N_19063,N_16444);
xnor U20136 (N_20136,N_15457,N_19134);
nand U20137 (N_20137,N_19061,N_19571);
nor U20138 (N_20138,N_17038,N_16255);
xnor U20139 (N_20139,N_16241,N_15027);
xnor U20140 (N_20140,N_18749,N_19605);
or U20141 (N_20141,N_17333,N_17991);
and U20142 (N_20142,N_18541,N_19048);
nor U20143 (N_20143,N_17822,N_19954);
nor U20144 (N_20144,N_16112,N_15929);
or U20145 (N_20145,N_15073,N_18100);
and U20146 (N_20146,N_15321,N_18640);
nor U20147 (N_20147,N_15109,N_17289);
nor U20148 (N_20148,N_16367,N_15578);
xor U20149 (N_20149,N_19040,N_19216);
or U20150 (N_20150,N_15580,N_19323);
and U20151 (N_20151,N_18957,N_15705);
nand U20152 (N_20152,N_19095,N_19173);
and U20153 (N_20153,N_15875,N_16645);
xor U20154 (N_20154,N_18833,N_16363);
or U20155 (N_20155,N_19537,N_16466);
or U20156 (N_20156,N_19938,N_19135);
nand U20157 (N_20157,N_17440,N_18275);
and U20158 (N_20158,N_16044,N_19399);
or U20159 (N_20159,N_17765,N_17774);
or U20160 (N_20160,N_17217,N_18772);
nand U20161 (N_20161,N_19045,N_18081);
and U20162 (N_20162,N_18467,N_15346);
and U20163 (N_20163,N_15282,N_19970);
or U20164 (N_20164,N_16814,N_17883);
nor U20165 (N_20165,N_19096,N_19090);
or U20166 (N_20166,N_16574,N_19748);
and U20167 (N_20167,N_19066,N_16572);
xnor U20168 (N_20168,N_18249,N_17727);
xor U20169 (N_20169,N_15264,N_16932);
or U20170 (N_20170,N_15667,N_15091);
or U20171 (N_20171,N_15832,N_19690);
and U20172 (N_20172,N_19902,N_18334);
and U20173 (N_20173,N_18924,N_15906);
nor U20174 (N_20174,N_17489,N_16300);
nor U20175 (N_20175,N_17152,N_19710);
and U20176 (N_20176,N_18413,N_16626);
or U20177 (N_20177,N_17043,N_18444);
nor U20178 (N_20178,N_18618,N_19693);
and U20179 (N_20179,N_17042,N_18589);
nand U20180 (N_20180,N_18828,N_17288);
or U20181 (N_20181,N_17856,N_17030);
nor U20182 (N_20182,N_16054,N_18718);
nand U20183 (N_20183,N_17572,N_17051);
or U20184 (N_20184,N_15081,N_17672);
or U20185 (N_20185,N_19965,N_15101);
or U20186 (N_20186,N_19567,N_18810);
nor U20187 (N_20187,N_18926,N_16805);
and U20188 (N_20188,N_19945,N_16947);
nor U20189 (N_20189,N_19030,N_18977);
nand U20190 (N_20190,N_15257,N_16383);
or U20191 (N_20191,N_17968,N_16405);
nor U20192 (N_20192,N_15191,N_19892);
nand U20193 (N_20193,N_19994,N_15309);
nor U20194 (N_20194,N_17478,N_18497);
xnor U20195 (N_20195,N_18161,N_18396);
xor U20196 (N_20196,N_15725,N_17213);
xor U20197 (N_20197,N_15889,N_19648);
nand U20198 (N_20198,N_19149,N_16193);
nor U20199 (N_20199,N_18212,N_17120);
and U20200 (N_20200,N_18326,N_18530);
or U20201 (N_20201,N_15450,N_19009);
and U20202 (N_20202,N_19526,N_17026);
and U20203 (N_20203,N_18830,N_15461);
and U20204 (N_20204,N_16612,N_18381);
nand U20205 (N_20205,N_18919,N_16090);
xor U20206 (N_20206,N_16304,N_15124);
xnor U20207 (N_20207,N_18804,N_19980);
nor U20208 (N_20208,N_15103,N_15225);
nand U20209 (N_20209,N_18599,N_17148);
nor U20210 (N_20210,N_16260,N_18976);
xnor U20211 (N_20211,N_15712,N_15438);
xnor U20212 (N_20212,N_16870,N_15055);
and U20213 (N_20213,N_19934,N_17186);
or U20214 (N_20214,N_15287,N_17384);
or U20215 (N_20215,N_19806,N_15216);
and U20216 (N_20216,N_17522,N_17983);
xnor U20217 (N_20217,N_16017,N_16605);
xnor U20218 (N_20218,N_16075,N_15009);
or U20219 (N_20219,N_18079,N_16586);
xor U20220 (N_20220,N_15293,N_18860);
or U20221 (N_20221,N_16631,N_17491);
or U20222 (N_20222,N_19865,N_18290);
and U20223 (N_20223,N_19671,N_17464);
nor U20224 (N_20224,N_18914,N_16129);
and U20225 (N_20225,N_18215,N_16616);
xnor U20226 (N_20226,N_15599,N_19656);
nand U20227 (N_20227,N_17409,N_17861);
nand U20228 (N_20228,N_15779,N_16122);
and U20229 (N_20229,N_18567,N_15270);
or U20230 (N_20230,N_18598,N_17111);
and U20231 (N_20231,N_17484,N_15917);
nand U20232 (N_20232,N_18349,N_16168);
xor U20233 (N_20233,N_18179,N_16012);
nor U20234 (N_20234,N_18461,N_18412);
nor U20235 (N_20235,N_15715,N_15567);
or U20236 (N_20236,N_17339,N_15833);
nand U20237 (N_20237,N_16787,N_16333);
nor U20238 (N_20238,N_16533,N_15834);
nor U20239 (N_20239,N_16077,N_18377);
and U20240 (N_20240,N_15253,N_18094);
nand U20241 (N_20241,N_17432,N_17322);
or U20242 (N_20242,N_19001,N_15565);
and U20243 (N_20243,N_19260,N_17730);
nor U20244 (N_20244,N_19370,N_16837);
or U20245 (N_20245,N_15830,N_19487);
nor U20246 (N_20246,N_19888,N_18827);
nor U20247 (N_20247,N_16194,N_17054);
or U20248 (N_20248,N_19803,N_17700);
or U20249 (N_20249,N_19989,N_16311);
and U20250 (N_20250,N_17281,N_15925);
xor U20251 (N_20251,N_17175,N_17503);
nand U20252 (N_20252,N_16490,N_18934);
and U20253 (N_20253,N_19686,N_17819);
and U20254 (N_20254,N_19776,N_18335);
nand U20255 (N_20255,N_16690,N_19258);
nand U20256 (N_20256,N_16551,N_19624);
xnor U20257 (N_20257,N_15186,N_15358);
nor U20258 (N_20258,N_16110,N_17718);
and U20259 (N_20259,N_16822,N_16469);
nor U20260 (N_20260,N_15513,N_17130);
nand U20261 (N_20261,N_16182,N_15463);
and U20262 (N_20262,N_16195,N_18090);
or U20263 (N_20263,N_19661,N_17623);
and U20264 (N_20264,N_16357,N_19010);
xor U20265 (N_20265,N_18710,N_18233);
nand U20266 (N_20266,N_15699,N_18979);
nand U20267 (N_20267,N_16053,N_18871);
nand U20268 (N_20268,N_18040,N_16297);
and U20269 (N_20269,N_17467,N_16468);
nand U20270 (N_20270,N_17525,N_19805);
nor U20271 (N_20271,N_16512,N_18388);
xnor U20272 (N_20272,N_17675,N_19855);
nor U20273 (N_20273,N_17200,N_15728);
and U20274 (N_20274,N_18517,N_15639);
nand U20275 (N_20275,N_15710,N_18111);
or U20276 (N_20276,N_16753,N_16557);
nand U20277 (N_20277,N_17233,N_15864);
nor U20278 (N_20278,N_16389,N_19633);
xor U20279 (N_20279,N_16292,N_18339);
xnor U20280 (N_20280,N_19312,N_19915);
or U20281 (N_20281,N_18133,N_15490);
and U20282 (N_20282,N_16585,N_17461);
nor U20283 (N_20283,N_19197,N_17684);
or U20284 (N_20284,N_17466,N_15846);
or U20285 (N_20285,N_17443,N_19670);
and U20286 (N_20286,N_19502,N_15263);
and U20287 (N_20287,N_18125,N_18384);
nor U20288 (N_20288,N_16208,N_19293);
xor U20289 (N_20289,N_19400,N_15290);
or U20290 (N_20290,N_19801,N_19218);
nand U20291 (N_20291,N_17729,N_17039);
xnor U20292 (N_20292,N_19510,N_15709);
and U20293 (N_20293,N_17108,N_15067);
or U20294 (N_20294,N_19829,N_18855);
and U20295 (N_20295,N_17070,N_17075);
and U20296 (N_20296,N_17257,N_15804);
nand U20297 (N_20297,N_19772,N_18839);
nand U20298 (N_20298,N_18043,N_19576);
nor U20299 (N_20299,N_15288,N_15538);
and U20300 (N_20300,N_18617,N_19616);
nand U20301 (N_20301,N_18829,N_15992);
xnor U20302 (N_20302,N_15942,N_15410);
and U20303 (N_20303,N_18027,N_15951);
or U20304 (N_20304,N_16035,N_19523);
or U20305 (N_20305,N_16346,N_15423);
and U20306 (N_20306,N_19240,N_19421);
or U20307 (N_20307,N_18380,N_17243);
and U20308 (N_20308,N_17476,N_16069);
nand U20309 (N_20309,N_19442,N_15203);
xor U20310 (N_20310,N_18626,N_15492);
or U20311 (N_20311,N_17511,N_17320);
nand U20312 (N_20312,N_17437,N_16368);
xnor U20313 (N_20313,N_19128,N_19968);
xor U20314 (N_20314,N_18310,N_16659);
and U20315 (N_20315,N_19423,N_16985);
and U20316 (N_20316,N_18942,N_16066);
nand U20317 (N_20317,N_17643,N_16237);
or U20318 (N_20318,N_16886,N_17113);
xnor U20319 (N_20319,N_18945,N_17362);
nor U20320 (N_20320,N_19271,N_19292);
and U20321 (N_20321,N_18166,N_19575);
xor U20322 (N_20322,N_15129,N_16011);
and U20323 (N_20323,N_17829,N_19785);
nand U20324 (N_20324,N_17329,N_17386);
xnor U20325 (N_20325,N_15327,N_19739);
nor U20326 (N_20326,N_18389,N_15277);
nand U20327 (N_20327,N_16222,N_15395);
nand U20328 (N_20328,N_19610,N_15390);
and U20329 (N_20329,N_18099,N_18064);
xor U20330 (N_20330,N_17536,N_15175);
and U20331 (N_20331,N_15212,N_16421);
nand U20332 (N_20332,N_18563,N_18247);
and U20333 (N_20333,N_19543,N_19737);
and U20334 (N_20334,N_19018,N_19490);
and U20335 (N_20335,N_19908,N_19696);
nor U20336 (N_20336,N_19559,N_17207);
and U20337 (N_20337,N_19434,N_17543);
xor U20338 (N_20338,N_16016,N_18244);
nand U20339 (N_20339,N_17450,N_17926);
and U20340 (N_20340,N_15343,N_16515);
nor U20341 (N_20341,N_19205,N_16505);
xor U20342 (N_20342,N_16714,N_17598);
nor U20343 (N_20343,N_17297,N_19286);
nor U20344 (N_20344,N_18395,N_16253);
and U20345 (N_20345,N_19977,N_16442);
or U20346 (N_20346,N_18673,N_19741);
xnor U20347 (N_20347,N_16769,N_18462);
and U20348 (N_20348,N_15556,N_16820);
or U20349 (N_20349,N_17715,N_18083);
nor U20350 (N_20350,N_16470,N_18889);
or U20351 (N_20351,N_16731,N_17092);
xor U20352 (N_20352,N_16609,N_15963);
xor U20353 (N_20353,N_17341,N_18521);
or U20354 (N_20354,N_17949,N_15772);
or U20355 (N_20355,N_17622,N_17568);
nor U20356 (N_20356,N_17769,N_18753);
xnor U20357 (N_20357,N_16918,N_19719);
nand U20358 (N_20358,N_19669,N_15004);
nor U20359 (N_20359,N_18512,N_16177);
nor U20360 (N_20360,N_18262,N_19156);
nand U20361 (N_20361,N_15054,N_15482);
xnor U20362 (N_20362,N_17295,N_19296);
nand U20363 (N_20363,N_16931,N_16282);
or U20364 (N_20364,N_17671,N_15708);
or U20365 (N_20365,N_15069,N_16638);
nand U20366 (N_20366,N_19773,N_19005);
nand U20367 (N_20367,N_15105,N_16747);
xor U20368 (N_20368,N_19174,N_15912);
xnor U20369 (N_20369,N_18613,N_17451);
xnor U20370 (N_20370,N_19897,N_17911);
nand U20371 (N_20371,N_17331,N_18251);
nand U20372 (N_20372,N_18476,N_15958);
nand U20373 (N_20373,N_19450,N_17888);
xor U20374 (N_20374,N_18146,N_16211);
and U20375 (N_20375,N_18201,N_18021);
xor U20376 (N_20376,N_15615,N_17745);
and U20377 (N_20377,N_19767,N_19080);
nor U20378 (N_20378,N_17264,N_17789);
nor U20379 (N_20379,N_16547,N_19856);
nor U20380 (N_20380,N_15469,N_16473);
xor U20381 (N_20381,N_16732,N_18509);
and U20382 (N_20382,N_16330,N_17025);
or U20383 (N_20383,N_17833,N_19881);
and U20384 (N_20384,N_16589,N_19362);
nor U20385 (N_20385,N_18963,N_18695);
nand U20386 (N_20386,N_18165,N_19283);
xnor U20387 (N_20387,N_15620,N_15142);
or U20388 (N_20388,N_19081,N_19247);
nand U20389 (N_20389,N_17462,N_18824);
or U20390 (N_20390,N_18117,N_15933);
nor U20391 (N_20391,N_15800,N_18452);
and U20392 (N_20392,N_17285,N_19484);
nand U20393 (N_20393,N_18098,N_19879);
nor U20394 (N_20394,N_18226,N_17823);
or U20395 (N_20395,N_17371,N_18366);
xor U20396 (N_20396,N_19448,N_17270);
and U20397 (N_20397,N_17855,N_18999);
nor U20398 (N_20398,N_19058,N_18642);
and U20399 (N_20399,N_19603,N_16390);
nand U20400 (N_20400,N_17098,N_16104);
and U20401 (N_20401,N_18494,N_16789);
and U20402 (N_20402,N_19663,N_17212);
and U20403 (N_20403,N_19447,N_18204);
nor U20404 (N_20404,N_19899,N_15941);
and U20405 (N_20405,N_16451,N_17293);
xnor U20406 (N_20406,N_18536,N_16613);
or U20407 (N_20407,N_19665,N_16232);
nand U20408 (N_20408,N_18011,N_16800);
nor U20409 (N_20409,N_17758,N_15178);
or U20410 (N_20410,N_19532,N_19560);
or U20411 (N_20411,N_18566,N_16158);
nand U20412 (N_20412,N_18767,N_15525);
and U20413 (N_20413,N_17274,N_17685);
xnor U20414 (N_20414,N_16399,N_19883);
nor U20415 (N_20415,N_17766,N_18260);
nor U20416 (N_20416,N_17799,N_15966);
nor U20417 (N_20417,N_19319,N_18940);
xnor U20418 (N_20418,N_19735,N_15592);
nor U20419 (N_20419,N_15582,N_16951);
and U20420 (N_20420,N_18093,N_19652);
and U20421 (N_20421,N_18200,N_19092);
or U20422 (N_20422,N_15351,N_18097);
xor U20423 (N_20423,N_15137,N_18714);
and U20424 (N_20424,N_17402,N_17990);
xnor U20425 (N_20425,N_18082,N_16173);
and U20426 (N_20426,N_15119,N_19987);
or U20427 (N_20427,N_15738,N_16554);
or U20428 (N_20428,N_15892,N_18057);
nand U20429 (N_20429,N_15669,N_15862);
and U20430 (N_20430,N_16449,N_17428);
and U20431 (N_20431,N_16127,N_16565);
xor U20432 (N_20432,N_15495,N_18795);
nor U20433 (N_20433,N_17249,N_15707);
nor U20434 (N_20434,N_15817,N_16422);
nand U20435 (N_20435,N_15690,N_17225);
and U20436 (N_20436,N_18779,N_17050);
nor U20437 (N_20437,N_19723,N_18351);
nand U20438 (N_20438,N_18593,N_17697);
or U20439 (N_20439,N_18986,N_15882);
or U20440 (N_20440,N_18713,N_16461);
or U20441 (N_20441,N_17920,N_15701);
xor U20442 (N_20442,N_17520,N_18288);
or U20443 (N_20443,N_17974,N_17618);
xnor U20444 (N_20444,N_18263,N_18811);
nand U20445 (N_20445,N_19931,N_17076);
or U20446 (N_20446,N_19389,N_16114);
nand U20447 (N_20447,N_18978,N_16676);
xnor U20448 (N_20448,N_16150,N_19783);
nor U20449 (N_20449,N_17040,N_15447);
xor U20450 (N_20450,N_19409,N_19570);
nand U20451 (N_20451,N_16994,N_15507);
xnor U20452 (N_20452,N_15498,N_19390);
nand U20453 (N_20453,N_19179,N_16454);
xnor U20454 (N_20454,N_19355,N_18186);
xor U20455 (N_20455,N_16776,N_17492);
or U20456 (N_20456,N_18794,N_19426);
xnor U20457 (N_20457,N_16818,N_18692);
xnor U20458 (N_20458,N_16321,N_17146);
and U20459 (N_20459,N_16244,N_17997);
nand U20460 (N_20460,N_17360,N_16998);
nand U20461 (N_20461,N_19694,N_17967);
nand U20462 (N_20462,N_17865,N_17154);
nor U20463 (N_20463,N_19636,N_19678);
nand U20464 (N_20464,N_16051,N_16025);
and U20465 (N_20465,N_18411,N_18682);
nand U20466 (N_20466,N_16492,N_18591);
nor U20467 (N_20467,N_16190,N_15767);
and U20468 (N_20468,N_15559,N_16989);
and U20469 (N_20469,N_19078,N_18602);
nor U20470 (N_20470,N_15890,N_16520);
xnor U20471 (N_20471,N_16698,N_19138);
and U20472 (N_20472,N_19632,N_15534);
nand U20473 (N_20473,N_15784,N_18835);
or U20474 (N_20474,N_19943,N_18597);
and U20475 (N_20475,N_16446,N_19219);
nor U20476 (N_20476,N_17960,N_19022);
nor U20477 (N_20477,N_15776,N_18523);
nand U20478 (N_20478,N_16773,N_19113);
nand U20479 (N_20479,N_18048,N_18107);
and U20480 (N_20480,N_15801,N_16269);
and U20481 (N_20481,N_18070,N_15745);
or U20482 (N_20482,N_16435,N_17176);
nand U20483 (N_20483,N_17665,N_18437);
or U20484 (N_20484,N_17104,N_15653);
nand U20485 (N_20485,N_17452,N_15157);
and U20486 (N_20486,N_17242,N_19637);
xor U20487 (N_20487,N_18751,N_18876);
nor U20488 (N_20488,N_17223,N_16600);
and U20489 (N_20489,N_19795,N_19918);
nor U20490 (N_20490,N_17204,N_19591);
xnor U20491 (N_20491,N_19425,N_15064);
nand U20492 (N_20492,N_17015,N_16970);
xor U20493 (N_20493,N_17326,N_16892);
nor U20494 (N_20494,N_19211,N_17961);
or U20495 (N_20495,N_17147,N_17749);
or U20496 (N_20496,N_18343,N_15298);
nor U20497 (N_20497,N_17860,N_17899);
nor U20498 (N_20498,N_19208,N_16360);
and U20499 (N_20499,N_19734,N_18734);
xnor U20500 (N_20500,N_15421,N_19394);
nor U20501 (N_20501,N_17348,N_15062);
xor U20502 (N_20502,N_19659,N_16413);
nand U20503 (N_20503,N_15575,N_17215);
or U20504 (N_20504,N_19726,N_18701);
and U20505 (N_20505,N_19979,N_16081);
xnor U20506 (N_20506,N_16957,N_17741);
or U20507 (N_20507,N_18390,N_15985);
nand U20508 (N_20508,N_16229,N_16326);
nor U20509 (N_20509,N_16906,N_16325);
nor U20510 (N_20510,N_15995,N_19887);
nand U20511 (N_20511,N_17442,N_15655);
and U20512 (N_20512,N_18899,N_16428);
or U20513 (N_20513,N_19963,N_16535);
or U20514 (N_20514,N_18327,N_19736);
nand U20515 (N_20515,N_16270,N_18472);
or U20516 (N_20516,N_16700,N_16423);
or U20517 (N_20517,N_15118,N_18585);
nor U20518 (N_20518,N_17621,N_16096);
and U20519 (N_20519,N_19891,N_18502);
and U20520 (N_20520,N_16704,N_17009);
or U20521 (N_20521,N_19026,N_19190);
nor U20522 (N_20522,N_18672,N_17194);
nand U20523 (N_20523,N_18344,N_18239);
xnor U20524 (N_20524,N_16827,N_15496);
and U20525 (N_20525,N_16485,N_17722);
or U20526 (N_20526,N_18652,N_15549);
xor U20527 (N_20527,N_19952,N_18101);
nand U20528 (N_20528,N_16106,N_19295);
xor U20529 (N_20529,N_17832,N_16322);
and U20530 (N_20530,N_15029,N_18034);
and U20531 (N_20531,N_16808,N_15065);
nand U20532 (N_20532,N_15299,N_17309);
or U20533 (N_20533,N_17034,N_19530);
or U20534 (N_20534,N_15747,N_19015);
nor U20535 (N_20535,N_19422,N_16577);
nor U20536 (N_20536,N_18328,N_15260);
or U20537 (N_20537,N_18549,N_19972);
and U20538 (N_20538,N_19322,N_15827);
and U20539 (N_20539,N_16472,N_18685);
xnor U20540 (N_20540,N_16040,N_17301);
nor U20541 (N_20541,N_18931,N_18294);
xor U20542 (N_20542,N_19701,N_15070);
and U20543 (N_20543,N_15824,N_15842);
or U20544 (N_20544,N_17397,N_19384);
and U20545 (N_20545,N_18202,N_19778);
nor U20546 (N_20546,N_19545,N_18500);
and U20547 (N_20547,N_18121,N_17493);
nor U20548 (N_20548,N_17554,N_16266);
nand U20549 (N_20549,N_16358,N_19290);
nand U20550 (N_20550,N_15671,N_16507);
or U20551 (N_20551,N_16909,N_15603);
or U20552 (N_20552,N_18746,N_19168);
nor U20553 (N_20553,N_16201,N_15007);
or U20554 (N_20554,N_19222,N_18709);
nor U20555 (N_20555,N_18910,N_15718);
nor U20556 (N_20556,N_17781,N_15053);
and U20557 (N_20557,N_16356,N_15074);
nand U20558 (N_20558,N_16763,N_18501);
and U20559 (N_20559,N_17998,N_19352);
or U20560 (N_20560,N_19137,N_16474);
nor U20561 (N_20561,N_17065,N_19895);
nor U20562 (N_20562,N_19099,N_18329);
and U20563 (N_20563,N_15588,N_17118);
and U20564 (N_20564,N_19574,N_15553);
or U20565 (N_20565,N_16691,N_15355);
or U20566 (N_20566,N_16530,N_19315);
and U20567 (N_20567,N_18927,N_17754);
nor U20568 (N_20568,N_19131,N_15713);
nor U20569 (N_20569,N_17680,N_17534);
and U20570 (N_20570,N_15609,N_19792);
nand U20571 (N_20571,N_17648,N_16031);
and U20572 (N_20572,N_15952,N_16807);
and U20573 (N_20573,N_19821,N_16802);
or U20574 (N_20574,N_18571,N_16569);
nand U20575 (N_20575,N_17825,N_17434);
nand U20576 (N_20576,N_18921,N_17993);
and U20577 (N_20577,N_16597,N_15694);
and U20578 (N_20578,N_16527,N_15477);
and U20579 (N_20579,N_17963,N_18551);
or U20580 (N_20580,N_15189,N_18990);
or U20581 (N_20581,N_15312,N_17699);
xnor U20582 (N_20582,N_19453,N_19430);
or U20583 (N_20583,N_18374,N_18657);
and U20584 (N_20584,N_17506,N_15262);
and U20585 (N_20585,N_19521,N_17321);
xnor U20586 (N_20586,N_16196,N_19905);
nor U20587 (N_20587,N_16639,N_16063);
or U20588 (N_20588,N_15094,N_15362);
xor U20589 (N_20589,N_15673,N_15570);
or U20590 (N_20590,N_15646,N_19599);
xor U20591 (N_20591,N_15080,N_18891);
nor U20592 (N_20592,N_16729,N_17306);
or U20593 (N_20593,N_16362,N_17595);
and U20594 (N_20594,N_19003,N_18798);
and U20595 (N_20595,N_16192,N_16878);
nor U20596 (N_20596,N_18844,N_15940);
and U20597 (N_20597,N_18789,N_18995);
xnor U20598 (N_20598,N_17439,N_15812);
nor U20599 (N_20599,N_16552,N_15978);
nor U20600 (N_20600,N_18320,N_15219);
xnor U20601 (N_20601,N_16944,N_18177);
or U20602 (N_20602,N_19781,N_18153);
or U20603 (N_20603,N_19330,N_17711);
xor U20604 (N_20604,N_19374,N_15944);
nand U20605 (N_20605,N_15744,N_19380);
and U20606 (N_20606,N_19207,N_18401);
or U20607 (N_20607,N_19615,N_16102);
nand U20608 (N_20608,N_17918,N_16912);
nand U20609 (N_20609,N_19765,N_19120);
xor U20610 (N_20610,N_15751,N_18837);
nand U20611 (N_20611,N_19985,N_15683);
nand U20612 (N_20612,N_17017,N_19962);
xnor U20613 (N_20613,N_16412,N_18893);
nor U20614 (N_20614,N_18514,N_15894);
or U20615 (N_20615,N_15179,N_16420);
xnor U20616 (N_20616,N_16873,N_18834);
and U20617 (N_20617,N_18866,N_15964);
xnor U20618 (N_20618,N_16480,N_19332);
nand U20619 (N_20619,N_18143,N_17922);
xnor U20620 (N_20620,N_17182,N_16476);
xor U20621 (N_20621,N_18688,N_19424);
nor U20622 (N_20622,N_18151,N_19587);
and U20623 (N_20623,N_15135,N_17539);
or U20624 (N_20624,N_15205,N_15937);
nand U20625 (N_20625,N_16189,N_16607);
nand U20626 (N_20626,N_17143,N_18558);
nand U20627 (N_20627,N_15823,N_15612);
nor U20628 (N_20628,N_15122,N_15340);
or U20629 (N_20629,N_15759,N_19921);
and U20630 (N_20630,N_19706,N_15286);
xnor U20631 (N_20631,N_18880,N_17019);
nor U20632 (N_20632,N_18577,N_16397);
and U20633 (N_20633,N_18628,N_16022);
nor U20634 (N_20634,N_18907,N_16228);
nand U20635 (N_20635,N_17078,N_16543);
xnor U20636 (N_20636,N_17517,N_19578);
and U20637 (N_20637,N_19976,N_18974);
or U20638 (N_20638,N_16347,N_17366);
or U20639 (N_20639,N_17142,N_18105);
and U20640 (N_20640,N_19655,N_17873);
xor U20641 (N_20641,N_15023,N_17299);
nand U20642 (N_20642,N_19998,N_17724);
or U20643 (N_20643,N_18207,N_15829);
xnor U20644 (N_20644,N_19702,N_18885);
nand U20645 (N_20645,N_16137,N_18524);
nand U20646 (N_20646,N_15140,N_19102);
nand U20647 (N_20647,N_17115,N_17073);
nor U20648 (N_20648,N_19850,N_16256);
or U20649 (N_20649,N_19491,N_18498);
and U20650 (N_20650,N_17791,N_19847);
nor U20651 (N_20651,N_16717,N_15419);
nor U20652 (N_20652,N_16078,N_16525);
nand U20653 (N_20653,N_16414,N_18474);
or U20654 (N_20654,N_17468,N_15562);
or U20655 (N_20655,N_18248,N_17469);
xnor U20656 (N_20656,N_19863,N_17705);
nor U20657 (N_20657,N_15872,N_16294);
nand U20658 (N_20658,N_15153,N_16561);
or U20659 (N_20659,N_15084,N_15434);
nand U20660 (N_20660,N_15485,N_15627);
xor U20661 (N_20661,N_15893,N_16488);
nand U20662 (N_20662,N_18039,N_17198);
and U20663 (N_20663,N_17939,N_18721);
and U20664 (N_20664,N_15611,N_17071);
nand U20665 (N_20665,N_16034,N_16313);
nand U20666 (N_20666,N_16199,N_18637);
or U20667 (N_20667,N_17008,N_15628);
nor U20668 (N_20668,N_15459,N_19035);
and U20669 (N_20669,N_19367,N_19628);
nor U20670 (N_20670,N_18647,N_15316);
nand U20671 (N_20671,N_18886,N_17294);
nor U20672 (N_20672,N_19172,N_16783);
nor U20673 (N_20673,N_17112,N_19715);
xor U20674 (N_20674,N_15857,N_19504);
nand U20675 (N_20675,N_17677,N_19871);
nor U20676 (N_20676,N_18668,N_19834);
nor U20677 (N_20677,N_18430,N_15594);
nand U20678 (N_20678,N_16694,N_15195);
nand U20679 (N_20679,N_17129,N_16164);
nand U20680 (N_20680,N_17653,N_19681);
xnor U20681 (N_20681,N_19501,N_17337);
or U20682 (N_20682,N_18821,N_15196);
or U20683 (N_20683,N_18050,N_17166);
xor U20684 (N_20684,N_15380,N_18731);
nand U20685 (N_20685,N_19088,N_18755);
and U20686 (N_20686,N_17364,N_16982);
xor U20687 (N_20687,N_19631,N_16738);
xor U20688 (N_20688,N_17080,N_17061);
xor U20689 (N_20689,N_18973,N_18254);
nor U20690 (N_20690,N_19171,N_15167);
nor U20691 (N_20691,N_17770,N_15662);
and U20692 (N_20692,N_19186,N_19711);
xnor U20693 (N_20693,N_17921,N_18160);
xnor U20694 (N_20694,N_17095,N_17752);
nand U20695 (N_20695,N_18980,N_16867);
nor U20696 (N_20696,N_16529,N_15953);
and U20697 (N_20697,N_16157,N_17445);
nand U20698 (N_20698,N_19123,N_17325);
xnor U20699 (N_20699,N_18610,N_18302);
nor U20700 (N_20700,N_17889,N_17958);
nor U20701 (N_20701,N_18190,N_17691);
xor U20702 (N_20702,N_19697,N_17497);
nand U20703 (N_20703,N_18892,N_17940);
or U20704 (N_20704,N_18601,N_19547);
nor U20705 (N_20705,N_16301,N_18962);
xnor U20706 (N_20706,N_18132,N_15274);
nand U20707 (N_20707,N_15337,N_16275);
and U20708 (N_20708,N_15733,N_18991);
and U20709 (N_20709,N_15481,N_16828);
and U20710 (N_20710,N_16224,N_17391);
or U20711 (N_20711,N_17626,N_16916);
nor U20712 (N_20712,N_19083,N_19133);
nand U20713 (N_20713,N_16245,N_16352);
nand U20714 (N_20714,N_16992,N_16436);
nor U20715 (N_20715,N_16359,N_18743);
and U20716 (N_20716,N_16979,N_16746);
nor U20717 (N_20717,N_15519,N_19667);
and U20718 (N_20718,N_19760,N_15414);
and U20719 (N_20719,N_16558,N_15313);
xor U20720 (N_20720,N_18658,N_19775);
and U20721 (N_20721,N_18744,N_18382);
and U20722 (N_20722,N_19465,N_15033);
or U20723 (N_20723,N_18781,N_19791);
nor U20724 (N_20724,N_16080,N_17472);
nor U20725 (N_20725,N_17116,N_15675);
nor U20726 (N_20726,N_16430,N_16152);
or U20727 (N_20727,N_19860,N_17999);
nand U20728 (N_20728,N_16424,N_15867);
nor U20729 (N_20729,N_18386,N_16836);
nand U20730 (N_20730,N_19177,N_17844);
xor U20731 (N_20731,N_19704,N_15374);
or U20732 (N_20732,N_17251,N_15422);
or U20733 (N_20733,N_16457,N_16392);
xor U20734 (N_20734,N_16688,N_17028);
xor U20735 (N_20735,N_17347,N_19826);
xor U20736 (N_20736,N_19786,N_18869);
nand U20737 (N_20737,N_18587,N_19446);
nand U20738 (N_20738,N_17119,N_18550);
nor U20739 (N_20739,N_18482,N_19812);
or U20740 (N_20740,N_16398,N_19750);
and U20741 (N_20741,N_16929,N_15291);
xor U20742 (N_20742,N_16439,N_17839);
xnor U20743 (N_20743,N_16832,N_19452);
nor U20744 (N_20744,N_15051,N_15404);
nor U20745 (N_20745,N_18592,N_15483);
and U20746 (N_20746,N_17419,N_18378);
nand U20747 (N_20747,N_19869,N_15602);
and U20748 (N_20748,N_17415,N_19141);
nor U20749 (N_20749,N_16212,N_19071);
or U20750 (N_20750,N_15787,N_16086);
xnor U20751 (N_20751,N_18645,N_19483);
nor U20752 (N_20752,N_18434,N_19196);
xor U20753 (N_20753,N_17843,N_18449);
and U20754 (N_20754,N_16898,N_17374);
nand U20755 (N_20755,N_17721,N_16871);
nand U20756 (N_20756,N_17738,N_15222);
nand U20757 (N_20757,N_17310,N_18506);
and U20758 (N_20758,N_15468,N_15182);
nor U20759 (N_20759,N_18752,N_16254);
and U20760 (N_20760,N_18898,N_19901);
nor U20761 (N_20761,N_19658,N_17660);
nand U20762 (N_20762,N_18199,N_19960);
and U20763 (N_20763,N_16664,N_15143);
nand U20764 (N_20764,N_18629,N_17720);
nand U20765 (N_20765,N_17526,N_18641);
or U20766 (N_20766,N_15160,N_15401);
and U20767 (N_20767,N_19721,N_15896);
nor U20768 (N_20768,N_15991,N_16934);
nor U20769 (N_20769,N_15428,N_15529);
and U20770 (N_20770,N_16489,N_15255);
and U20771 (N_20771,N_16312,N_19224);
nand U20772 (N_20772,N_17624,N_16945);
or U20773 (N_20773,N_15561,N_15304);
xnor U20774 (N_20774,N_18946,N_17734);
xnor U20775 (N_20775,N_17657,N_15994);
or U20776 (N_20776,N_16203,N_16721);
nand U20777 (N_20777,N_17659,N_16981);
and U20778 (N_20778,N_18557,N_17094);
or U20779 (N_20779,N_15740,N_19489);
or U20780 (N_20780,N_18771,N_15443);
xnor U20781 (N_20781,N_19480,N_16540);
nand U20782 (N_20782,N_16162,N_19558);
xor U20783 (N_20783,N_19411,N_16518);
or U20784 (N_20784,N_19947,N_17954);
or U20785 (N_20785,N_16880,N_18913);
nor U20786 (N_20786,N_17267,N_19289);
xnor U20787 (N_20787,N_16642,N_16513);
or U20788 (N_20788,N_18220,N_19340);
or U20789 (N_20789,N_19992,N_19109);
or U20790 (N_20790,N_19520,N_17385);
or U20791 (N_20791,N_16378,N_15661);
nor U20792 (N_20792,N_18580,N_15735);
and U20793 (N_20793,N_19552,N_15546);
xor U20794 (N_20794,N_18292,N_16650);
or U20795 (N_20795,N_18801,N_17845);
xor U20796 (N_20796,N_18948,N_15214);
xnor U20797 (N_20797,N_15451,N_16772);
nor U20798 (N_20798,N_18067,N_16184);
or U20799 (N_20799,N_15541,N_19766);
and U20800 (N_20800,N_15757,N_19823);
nand U20801 (N_20801,N_16937,N_17591);
and U20802 (N_20802,N_18717,N_15858);
xor U20803 (N_20803,N_18438,N_19269);
nand U20804 (N_20804,N_15235,N_17037);
xor U20805 (N_20805,N_16741,N_18606);
xnor U20806 (N_20806,N_15162,N_16450);
nand U20807 (N_20807,N_18515,N_19562);
nor U20808 (N_20808,N_19391,N_15075);
nor U20809 (N_20809,N_17149,N_15790);
or U20810 (N_20810,N_18295,N_15887);
xnor U20811 (N_20811,N_15976,N_17917);
and U20812 (N_20812,N_19182,N_16987);
and U20813 (N_20813,N_16580,N_17782);
nand U20814 (N_20814,N_18393,N_16477);
nand U20815 (N_20815,N_16893,N_18918);
and U20816 (N_20816,N_18983,N_16136);
and U20817 (N_20817,N_15782,N_19572);
xor U20818 (N_20818,N_15018,N_15144);
nand U20819 (N_20819,N_17016,N_15852);
nand U20820 (N_20820,N_17079,N_15014);
nand U20821 (N_20821,N_16662,N_15853);
nand U20822 (N_20822,N_18475,N_17060);
nor U20823 (N_20823,N_15859,N_19476);
nand U20824 (N_20824,N_19627,N_18022);
xor U20825 (N_20825,N_16966,N_17454);
xnor U20826 (N_20826,N_17361,N_18542);
or U20827 (N_20827,N_18938,N_18904);
nor U20828 (N_20828,N_16858,N_17353);
or U20829 (N_20829,N_19975,N_15335);
or U20830 (N_20830,N_17638,N_19512);
xor U20831 (N_20831,N_18157,N_18228);
nand U20832 (N_20832,N_15425,N_17027);
or U20833 (N_20833,N_15980,N_17795);
and U20834 (N_20834,N_19481,N_17663);
and U20835 (N_20835,N_19822,N_19420);
or U20836 (N_20836,N_17163,N_16921);
or U20837 (N_20837,N_15973,N_17059);
and U20838 (N_20838,N_15325,N_17252);
xor U20839 (N_20839,N_19351,N_18759);
xnor U20840 (N_20840,N_15831,N_18841);
or U20841 (N_20841,N_18737,N_18929);
xnor U20842 (N_20842,N_15112,N_17646);
xnor U20843 (N_20843,N_17788,N_17001);
nand U20844 (N_20844,N_16381,N_17532);
and U20845 (N_20845,N_18951,N_16088);
xor U20846 (N_20846,N_16443,N_15159);
or U20847 (N_20847,N_16438,N_18347);
xor U20848 (N_20848,N_16845,N_15798);
nand U20849 (N_20849,N_16617,N_18035);
nor U20850 (N_20850,N_17914,N_16248);
or U20851 (N_20851,N_15352,N_17537);
and U20852 (N_20852,N_18192,N_18236);
and U20853 (N_20853,N_19376,N_18783);
nor U20854 (N_20854,N_17710,N_16978);
nand U20855 (N_20855,N_19561,N_18852);
nor U20856 (N_20856,N_19692,N_15695);
or U20857 (N_20857,N_16897,N_16286);
xor U20858 (N_20858,N_17636,N_17498);
or U20859 (N_20859,N_18769,N_16955);
nor U20860 (N_20860,N_15096,N_17919);
nand U20861 (N_20861,N_16720,N_15596);
and U20862 (N_20862,N_16277,N_19220);
nand U20863 (N_20863,N_16973,N_17985);
and U20864 (N_20864,N_18154,N_19272);
or U20865 (N_20865,N_17286,N_18397);
nand U20866 (N_20866,N_18609,N_15020);
or U20867 (N_20867,N_19275,N_15900);
nand U20868 (N_20868,N_17712,N_18322);
nand U20869 (N_20869,N_17193,N_18819);
xnor U20870 (N_20870,N_18554,N_18756);
and U20871 (N_20871,N_19714,N_16952);
nand U20872 (N_20872,N_16584,N_18796);
nand U20873 (N_20873,N_19335,N_19163);
xor U20874 (N_20874,N_18069,N_17927);
and U20875 (N_20875,N_16343,N_19799);
xnor U20876 (N_20876,N_17599,N_17367);
or U20877 (N_20877,N_16782,N_17857);
xor U20878 (N_20878,N_17036,N_19361);
nand U20879 (N_20879,N_17241,N_18198);
nand U20880 (N_20880,N_15474,N_19933);
or U20881 (N_20881,N_18778,N_18144);
nor U20882 (N_20882,N_15161,N_19907);
nor U20883 (N_20883,N_17161,N_17227);
nor U20884 (N_20884,N_15783,N_16281);
nor U20885 (N_20885,N_19890,N_19236);
or U20886 (N_20886,N_19956,N_19200);
xnor U20887 (N_20887,N_16777,N_18865);
and U20888 (N_20888,N_18242,N_18061);
and U20889 (N_20889,N_17836,N_17846);
xor U20890 (N_20890,N_16583,N_17424);
nand U20891 (N_20891,N_17222,N_19824);
nand U20892 (N_20892,N_16877,N_17514);
and U20893 (N_20893,N_16553,N_17790);
or U20894 (N_20894,N_15458,N_16209);
or U20895 (N_20895,N_15622,N_19014);
nor U20896 (N_20896,N_15810,N_17746);
and U20897 (N_20897,N_16813,N_19841);
nor U20898 (N_20898,N_16250,N_15001);
and U20899 (N_20899,N_19103,N_17664);
and U20900 (N_20900,N_18319,N_17527);
nand U20901 (N_20901,N_16904,N_15015);
and U20902 (N_20902,N_16756,N_16309);
nor U20903 (N_20903,N_15249,N_17303);
nand U20904 (N_20904,N_19722,N_15147);
xor U20905 (N_20905,N_16464,N_19046);
and U20906 (N_20906,N_17499,N_16914);
and U20907 (N_20907,N_16999,N_17218);
nor U20908 (N_20908,N_16234,N_15868);
and U20909 (N_20909,N_18768,N_16582);
nand U20910 (N_20910,N_18576,N_18315);
xor U20911 (N_20911,N_16917,N_17316);
and U20912 (N_20912,N_19687,N_17551);
nand U20913 (N_20913,N_17645,N_18042);
nand U20914 (N_20914,N_15531,N_18806);
and U20915 (N_20915,N_19780,N_18446);
and U20916 (N_20916,N_15032,N_17913);
or U20917 (N_20917,N_19712,N_16154);
or U20918 (N_20918,N_17937,N_19935);
and U20919 (N_20919,N_17135,N_15926);
and U20920 (N_20920,N_17879,N_16739);
xnor U20921 (N_20921,N_18433,N_17496);
nor U20922 (N_20922,N_16133,N_19232);
xnor U20923 (N_20923,N_15658,N_19230);
nand U20924 (N_20924,N_15982,N_18856);
xnor U20925 (N_20925,N_17929,N_18345);
nand U20926 (N_20926,N_19032,N_19259);
or U20927 (N_20927,N_15849,N_16524);
xnor U20928 (N_20928,N_18791,N_15110);
or U20929 (N_20929,N_17633,N_16939);
and U20930 (N_20930,N_18255,N_16188);
and U20931 (N_20931,N_18608,N_19203);
or U20932 (N_20932,N_17045,N_19255);
nand U20933 (N_20933,N_15047,N_16009);
xor U20934 (N_20934,N_19238,N_16842);
nor U20935 (N_20935,N_18634,N_15731);
and U20936 (N_20936,N_18422,N_15895);
nand U20937 (N_20937,N_19527,N_19534);
nor U20938 (N_20938,N_15814,N_16602);
and U20939 (N_20939,N_17516,N_16674);
and U20940 (N_20940,N_19500,N_19012);
nor U20941 (N_20941,N_19708,N_17719);
xor U20942 (N_20942,N_18520,N_15281);
and U20943 (N_20943,N_17797,N_17523);
nand U20944 (N_20944,N_19796,N_15123);
and U20945 (N_20945,N_18964,N_19126);
xnor U20946 (N_20946,N_15489,N_15292);
xor U20947 (N_20947,N_15330,N_19233);
nand U20948 (N_20948,N_15138,N_15785);
or U20949 (N_20949,N_19325,N_15442);
nand U20950 (N_20950,N_19486,N_18159);
and U20951 (N_20951,N_18552,N_15663);
xnor U20952 (N_20952,N_16785,N_17368);
or U20953 (N_20953,N_16323,N_17673);
or U20954 (N_20954,N_16015,N_16064);
nor U20955 (N_20955,N_15502,N_16740);
and U20956 (N_20956,N_18604,N_15742);
or U20957 (N_20957,N_17945,N_17359);
or U20958 (N_20958,N_17931,N_19608);
or U20959 (N_20959,N_18142,N_16432);
xnor U20960 (N_20960,N_16504,N_15839);
nor U20961 (N_20961,N_18659,N_15218);
xnor U20962 (N_20962,N_17737,N_19579);
nor U20963 (N_20963,N_19245,N_19654);
nand U20964 (N_20964,N_15114,N_18969);
xor U20965 (N_20965,N_15107,N_15871);
xor U20966 (N_20966,N_15363,N_15907);
xor U20967 (N_20967,N_16202,N_17261);
and U20968 (N_20968,N_15795,N_18888);
xnor U20969 (N_20969,N_16372,N_16588);
or U20970 (N_20970,N_15430,N_19538);
and U20971 (N_20971,N_15237,N_15347);
xor U20972 (N_20972,N_15656,N_19730);
nor U20973 (N_20973,N_15883,N_18002);
nand U20974 (N_20974,N_18158,N_16848);
nor U20975 (N_20975,N_17803,N_19474);
and U20976 (N_20976,N_19235,N_15387);
nand U20977 (N_20977,N_16735,N_19742);
or U20978 (N_20978,N_18944,N_18440);
nand U20979 (N_20979,N_19350,N_19981);
or U20980 (N_20980,N_18987,N_17604);
nand U20981 (N_20981,N_19583,N_19611);
nor U20982 (N_20982,N_17315,N_15674);
or U20983 (N_20983,N_17023,N_16935);
nor U20984 (N_20984,N_15698,N_19584);
nor U20985 (N_20985,N_15721,N_15524);
nand U20986 (N_20986,N_18763,N_16695);
nand U20987 (N_20987,N_16008,N_18403);
and U20988 (N_20988,N_19282,N_19460);
and U20989 (N_20989,N_17760,N_19073);
nor U20990 (N_20990,N_15727,N_18235);
xor U20991 (N_20991,N_19617,N_19705);
nand U20992 (N_20992,N_15071,N_16502);
nand U20993 (N_20993,N_18120,N_15644);
and U20994 (N_20994,N_15154,N_19147);
nor U20995 (N_20995,N_19151,N_16759);
xor U20996 (N_20996,N_16682,N_15113);
xor U20997 (N_20997,N_18754,N_16665);
xnor U20998 (N_20998,N_15909,N_17588);
nor U20999 (N_20999,N_17508,N_16247);
nand U21000 (N_21000,N_19955,N_16467);
and U21001 (N_21001,N_18671,N_17750);
xnor U21002 (N_21002,N_15623,N_17934);
and U21003 (N_21003,N_16591,N_19913);
or U21004 (N_21004,N_17966,N_17413);
nand U21005 (N_21005,N_19485,N_15163);
nor U21006 (N_21006,N_17878,N_19209);
and U21007 (N_21007,N_17311,N_15530);
nand U21008 (N_21008,N_17755,N_16335);
nor U21009 (N_21009,N_19995,N_16331);
xnor U21010 (N_21010,N_18210,N_19160);
and U21011 (N_21011,N_18073,N_18092);
or U21012 (N_21012,N_17807,N_18807);
and U21013 (N_21013,N_19581,N_16594);
nand U21014 (N_21014,N_19564,N_19839);
nor U21015 (N_21015,N_17345,N_17757);
nor U21016 (N_21016,N_16076,N_18194);
or U21017 (N_21017,N_17136,N_19835);
nor U21018 (N_21018,N_18303,N_16391);
nand U21019 (N_21019,N_16891,N_15046);
or U21020 (N_21020,N_17804,N_17500);
nor U21021 (N_21021,N_17615,N_15736);
nand U21022 (N_21022,N_17151,N_19851);
nor U21023 (N_21023,N_18972,N_18431);
nor U21024 (N_21024,N_16298,N_19518);
and U21025 (N_21025,N_15680,N_19136);
xnor U21026 (N_21026,N_15019,N_18553);
nor U21027 (N_21027,N_17047,N_15151);
nand U21028 (N_21028,N_17029,N_15088);
nand U21029 (N_21029,N_15475,N_15252);
and U21030 (N_21030,N_19231,N_16646);
nand U21031 (N_21031,N_18750,N_17674);
and U21032 (N_21032,N_19492,N_19326);
xnor U21033 (N_21033,N_17378,N_16895);
xor U21034 (N_21034,N_17122,N_17188);
and U21035 (N_21035,N_18428,N_17678);
nor U21036 (N_21036,N_15271,N_16221);
and U21037 (N_21037,N_17005,N_16388);
nor U21038 (N_21038,N_17180,N_17933);
or U21039 (N_21039,N_19864,N_15318);
and U21040 (N_21040,N_15946,N_19782);
and U21041 (N_21041,N_16429,N_18216);
xnor U21042 (N_21042,N_17370,N_16233);
xnor U21043 (N_21043,N_17179,N_18333);
or U21044 (N_21044,N_16680,N_17407);
nand U21045 (N_21045,N_16825,N_16634);
and U21046 (N_21046,N_16291,N_17133);
nor U21047 (N_21047,N_19732,N_16060);
xor U21048 (N_21048,N_18785,N_18383);
and U21049 (N_21049,N_18410,N_15719);
nor U21050 (N_21050,N_19886,N_18932);
and U21051 (N_21051,N_18676,N_16903);
nand U21052 (N_21052,N_17486,N_18029);
and U21053 (N_21053,N_19329,N_18548);
nor U21054 (N_21054,N_18447,N_19317);
nand U21055 (N_21055,N_16988,N_15949);
or U21056 (N_21056,N_17069,N_15460);
xor U21057 (N_21057,N_16943,N_19769);
xor U21058 (N_21058,N_17244,N_15928);
and U21059 (N_21059,N_17088,N_19550);
or U21060 (N_21060,N_17247,N_18484);
and U21061 (N_21061,N_16755,N_16417);
nor U21062 (N_21062,N_19790,N_17811);
nor U21063 (N_21063,N_19004,N_16849);
nand U21064 (N_21064,N_18400,N_15233);
nor U21065 (N_21065,N_18126,N_19844);
and U21066 (N_21066,N_17651,N_18712);
nand U21067 (N_21067,N_16899,N_16350);
and U21068 (N_21068,N_16890,N_16647);
nand U21069 (N_21069,N_18503,N_19443);
or U21070 (N_21070,N_19988,N_16874);
and U21071 (N_21071,N_17404,N_18491);
nor U21072 (N_21072,N_17976,N_15455);
xor U21073 (N_21073,N_19342,N_17658);
or U21074 (N_21074,N_16799,N_17826);
xor U21075 (N_21075,N_19127,N_16094);
nand U21076 (N_21076,N_19144,N_18681);
nand U21077 (N_21077,N_19942,N_15104);
and U21078 (N_21078,N_16941,N_15317);
nor U21079 (N_21079,N_17905,N_18663);
nor U21080 (N_21080,N_16632,N_17904);
nor U21081 (N_21081,N_18241,N_18572);
and U21082 (N_21082,N_16599,N_15509);
xor U21083 (N_21083,N_17125,N_19339);
and U21084 (N_21084,N_17256,N_15278);
and U21085 (N_21085,N_16954,N_19488);
nand U21086 (N_21086,N_16481,N_18952);
xor U21087 (N_21087,N_15415,N_16262);
xnor U21088 (N_21088,N_16798,N_19724);
and U21089 (N_21089,N_19226,N_17058);
nand U21090 (N_21090,N_15256,N_19241);
nor U21091 (N_21091,N_15986,N_15021);
or U21092 (N_21092,N_18012,N_15837);
and U21093 (N_21093,N_18621,N_17821);
xnor U21094 (N_21094,N_15861,N_17463);
and U21095 (N_21095,N_18594,N_16206);
nand U21096 (N_21096,N_19903,N_17110);
xnor U21097 (N_21097,N_19438,N_18379);
nand U21098 (N_21098,N_15297,N_19589);
and U21099 (N_21099,N_15636,N_16374);
nand U21100 (N_21100,N_18387,N_18003);
xnor U21101 (N_21101,N_16653,N_18916);
or U21102 (N_21102,N_16259,N_18603);
nor U21103 (N_21103,N_15936,N_18293);
nand U21104 (N_21104,N_17481,N_15732);
xnor U21105 (N_21105,N_15634,N_18901);
nor U21106 (N_21106,N_19808,N_18847);
or U21107 (N_21107,N_16447,N_18285);
xnor U21108 (N_21108,N_16278,N_16623);
nor U21109 (N_21109,N_15813,N_17596);
nand U21110 (N_21110,N_17565,N_18209);
or U21111 (N_21111,N_15624,N_15356);
and U21112 (N_21112,N_17884,N_15170);
or U21113 (N_21113,N_15642,N_19062);
xor U21114 (N_21114,N_18304,N_15666);
nand U21115 (N_21115,N_17201,N_15384);
or U21116 (N_21116,N_16619,N_16083);
or U21117 (N_21117,N_19064,N_15217);
and U21118 (N_21118,N_17278,N_17507);
and U21119 (N_21119,N_19635,N_17117);
or U21120 (N_21120,N_18770,N_17987);
nand U21121 (N_21121,N_15454,N_18468);
and U21122 (N_21122,N_17834,N_18519);
and U21123 (N_21123,N_17938,N_19997);
and U21124 (N_21124,N_18532,N_16187);
and U21125 (N_21125,N_16089,N_16990);
nor U21126 (N_21126,N_19586,N_16426);
xor U21127 (N_21127,N_19522,N_16437);
and U21128 (N_21128,N_17880,N_18023);
or U21129 (N_21129,N_17909,N_15593);
and U21130 (N_21130,N_15999,N_18496);
xor U21131 (N_21131,N_18323,N_16026);
nor U21132 (N_21132,N_19508,N_19053);
xnor U21133 (N_21133,N_15417,N_15924);
xnor U21134 (N_21134,N_19287,N_15537);
xnor U21135 (N_21135,N_18808,N_19698);
and U21136 (N_21136,N_15532,N_17423);
and U21137 (N_21137,N_16754,N_16786);
xor U21138 (N_21138,N_19359,N_18526);
or U21139 (N_21139,N_17284,N_19588);
and U21140 (N_21140,N_16302,N_17886);
or U21141 (N_21141,N_15552,N_15311);
xnor U21142 (N_21142,N_17390,N_19919);
or U21143 (N_21143,N_16719,N_19878);
nor U21144 (N_21144,N_18538,N_19875);
or U21145 (N_21145,N_19779,N_16327);
nor U21146 (N_21146,N_16058,N_16062);
xnor U21147 (N_21147,N_15598,N_16596);
or U21148 (N_21148,N_17012,N_15572);
xnor U21149 (N_21149,N_19630,N_17817);
nor U21150 (N_21150,N_18905,N_17485);
nor U21151 (N_21151,N_18180,N_18638);
nand U21152 (N_21152,N_15983,N_17369);
xnor U21153 (N_21153,N_16462,N_15904);
xnor U21154 (N_21154,N_15960,N_17896);
nor U21155 (N_21155,N_18708,N_16857);
nand U21156 (N_21156,N_16334,N_16165);
nor U21157 (N_21157,N_17328,N_19301);
or U21158 (N_21158,N_15659,N_18562);
nor U21159 (N_21159,N_18301,N_17389);
xnor U21160 (N_21160,N_19418,N_17915);
and U21161 (N_21161,N_18761,N_16453);
and U21162 (N_21162,N_18836,N_17733);
and U21163 (N_21163,N_15396,N_18758);
nor U21164 (N_21164,N_19819,N_19911);
and U21165 (N_21165,N_17965,N_18049);
or U21166 (N_21166,N_19770,N_18677);
nand U21167 (N_21167,N_18309,N_15838);
or U21168 (N_21168,N_18136,N_15373);
nand U21169 (N_21169,N_16085,N_16865);
xnor U21170 (N_21170,N_18044,N_18465);
and U21171 (N_21171,N_18665,N_18481);
or U21172 (N_21172,N_15484,N_18072);
nand U21173 (N_21173,N_18661,N_16853);
and U21174 (N_21174,N_19397,N_17635);
nor U21175 (N_21175,N_17132,N_15510);
nand U21176 (N_21176,N_19318,N_18875);
and U21177 (N_21177,N_15777,N_17901);
nor U21178 (N_21178,N_17475,N_16751);
and U21179 (N_21179,N_19119,N_19951);
xnor U21180 (N_21180,N_17372,N_18902);
nor U21181 (N_21181,N_19900,N_19836);
nor U21182 (N_21182,N_18656,N_18488);
xnor U21183 (N_21183,N_16167,N_19405);
xor U21184 (N_21184,N_18217,N_16303);
xnor U21185 (N_21185,N_18321,N_18947);
and U21186 (N_21186,N_17171,N_18409);
nor U21187 (N_21187,N_16980,N_16907);
and U21188 (N_21188,N_17951,N_16339);
and U21189 (N_21189,N_19304,N_15187);
nand U21190 (N_21190,N_17510,N_17955);
or U21191 (N_21191,N_18715,N_19910);
and U21192 (N_21192,N_15497,N_15213);
xnor U21193 (N_21193,N_19445,N_16851);
nor U21194 (N_21194,N_17314,N_19274);
nor U21195 (N_21195,N_16149,N_15251);
xor U21196 (N_21196,N_19904,N_15515);
xor U21197 (N_21197,N_15600,N_15766);
xor U21198 (N_21198,N_17169,N_15246);
and U21199 (N_21199,N_19327,N_17533);
xnor U21200 (N_21200,N_19515,N_16748);
xnor U21201 (N_21201,N_17928,N_17031);
nor U21202 (N_21202,N_17662,N_16215);
and U21203 (N_21203,N_15797,N_16213);
xnor U21204 (N_21204,N_18355,N_16207);
nor U21205 (N_21205,N_17637,N_18473);
nor U21206 (N_21206,N_18561,N_15505);
nand U21207 (N_21207,N_16531,N_18031);
and U21208 (N_21208,N_18492,N_19983);
or U21209 (N_21209,N_17093,N_19195);
nor U21210 (N_21210,N_17425,N_19433);
and U21211 (N_21211,N_17731,N_17853);
nand U21212 (N_21212,N_17982,N_19029);
nand U21213 (N_21213,N_19193,N_17453);
or U21214 (N_21214,N_19105,N_19720);
and U21215 (N_21215,N_16750,N_16010);
nor U21216 (N_21216,N_17890,N_19978);
and U21217 (N_21217,N_19065,N_18308);
nor U21218 (N_21218,N_19067,N_16288);
nand U21219 (N_21219,N_15793,N_16147);
nand U21220 (N_21220,N_15433,N_18843);
nor U21221 (N_21221,N_19188,N_15465);
xnor U21222 (N_21222,N_17560,N_15324);
and U21223 (N_21223,N_19234,N_19516);
or U21224 (N_21224,N_17354,N_17650);
xnor U21225 (N_21225,N_15756,N_18719);
nand U21226 (N_21226,N_15243,N_17181);
or U21227 (N_21227,N_17696,N_16163);
xnor U21228 (N_21228,N_16306,N_18148);
xnor U21229 (N_21229,N_16622,N_18193);
and U21230 (N_21230,N_19820,N_19675);
nand U21231 (N_21231,N_19920,N_15635);
and U21232 (N_21232,N_17334,N_19288);
and U21233 (N_21233,N_15651,N_18711);
or U21234 (N_21234,N_16896,N_16757);
nor U21235 (N_21235,N_19825,N_16859);
nand U21236 (N_21236,N_17379,N_17265);
nand U21237 (N_21237,N_18646,N_18147);
nand U21238 (N_21238,N_15548,N_17590);
nand U21239 (N_21239,N_19021,N_16726);
nand U21240 (N_21240,N_17365,N_18909);
nand U21241 (N_21241,N_19703,N_15915);
nor U21242 (N_21242,N_15360,N_19279);
and U21243 (N_21243,N_15494,N_15342);
and U21244 (N_21244,N_16320,N_15045);
nor U21245 (N_21245,N_16536,N_17932);
or U21246 (N_21246,N_15626,N_16677);
xor U21247 (N_21247,N_19478,N_15765);
or U21248 (N_21248,N_17165,N_19740);
nor U21249 (N_21249,N_15672,N_17099);
or U21250 (N_21250,N_18607,N_15571);
xor U21251 (N_21251,N_18966,N_17195);
nand U21252 (N_21252,N_19257,N_19914);
or U21253 (N_21253,N_19169,N_16004);
and U21254 (N_21254,N_17101,N_17566);
and U21255 (N_21255,N_16002,N_16458);
and U21256 (N_21256,N_16793,N_17620);
nand U21257 (N_21257,N_17607,N_19093);
or U21258 (N_21258,N_18281,N_18221);
and U21259 (N_21259,N_15411,N_19996);
or U21260 (N_21260,N_17308,N_19112);
nor U21261 (N_21261,N_18780,N_17502);
nor U21262 (N_21262,N_17756,N_17702);
or U21263 (N_21263,N_19402,N_16993);
and U21264 (N_21264,N_19034,N_15200);
nor U21265 (N_21265,N_19387,N_19262);
nand U21266 (N_21266,N_18163,N_15645);
nor U21267 (N_21267,N_19870,N_16220);
or U21268 (N_21268,N_18988,N_18001);
nor U21269 (N_21269,N_16191,N_16496);
nand U21270 (N_21270,N_15305,N_19038);
or U21271 (N_21271,N_15763,N_17869);
and U21272 (N_21272,N_16835,N_19606);
or U21273 (N_21273,N_18191,N_15353);
nand U21274 (N_21274,N_17209,N_17894);
or U21275 (N_21275,N_18189,N_19115);
nor U21276 (N_21276,N_15934,N_16815);
or U21277 (N_21277,N_19152,N_16332);
and U21278 (N_21278,N_15227,N_17813);
nor U21279 (N_21279,N_15650,N_18777);
and U21280 (N_21280,N_18495,N_16790);
and U21281 (N_21281,N_15752,N_17842);
nand U21282 (N_21282,N_17302,N_16635);
or U21283 (N_21283,N_15471,N_19716);
nand U21284 (N_21284,N_18660,N_15402);
xnor U21285 (N_21285,N_19297,N_17714);
and U21286 (N_21286,N_16669,N_19243);
and U21287 (N_21287,N_16930,N_19041);
nand U21288 (N_21288,N_15848,N_16226);
nor U21289 (N_21289,N_15462,N_16708);
nor U21290 (N_21290,N_16218,N_15050);
nor U21291 (N_21291,N_17603,N_16651);
xor U21292 (N_21292,N_15039,N_17141);
and U21293 (N_21293,N_19444,N_16864);
xnor U21294 (N_21294,N_19143,N_18006);
or U21295 (N_21295,N_17573,N_17283);
or U21296 (N_21296,N_18203,N_19086);
nor U21297 (N_21297,N_15493,N_18135);
xnor U21298 (N_21298,N_18416,N_17022);
or U21299 (N_21299,N_15022,N_18747);
and U21300 (N_21300,N_15987,N_17344);
nor U21301 (N_21301,N_19140,N_16824);
and U21302 (N_21302,N_17726,N_18005);
xnor U21303 (N_21303,N_19626,N_16564);
nand U21304 (N_21304,N_17840,N_15863);
or U21305 (N_21305,N_18635,N_16811);
and U21306 (N_21306,N_16534,N_18846);
nor U21307 (N_21307,N_18662,N_19302);
or U21308 (N_21308,N_19316,N_15268);
or U21309 (N_21309,N_15136,N_17418);
xor U21310 (N_21310,N_18800,N_19331);
or U21311 (N_21311,N_15604,N_17084);
or U21312 (N_21312,N_16107,N_15517);
nor U21313 (N_21313,N_17989,N_19815);
and U21314 (N_21314,N_18872,N_16734);
nand U21315 (N_21315,N_18089,N_18056);
or U21316 (N_21316,N_15607,N_19454);
nor U21317 (N_21317,N_19563,N_19104);
and U21318 (N_21318,N_17438,N_17891);
nand U21319 (N_21319,N_19000,N_15880);
nor U21320 (N_21320,N_18000,N_19338);
nand U21321 (N_21321,N_17907,N_16562);
nand U21322 (N_21322,N_15366,N_18178);
nor U21323 (N_21323,N_19085,N_18252);
or U21324 (N_21324,N_15487,N_16030);
nor U21325 (N_21325,N_16427,N_16693);
nand U21326 (N_21326,N_17197,N_17538);
nor U21327 (N_21327,N_18528,N_19940);
nand U21328 (N_21328,N_19072,N_15574);
nor U21329 (N_21329,N_16709,N_18622);
xnor U21330 (N_21330,N_15377,N_15319);
xnor U21331 (N_21331,N_15467,N_18337);
xor U21332 (N_21332,N_17483,N_17126);
nor U21333 (N_21333,N_18776,N_17703);
and U21334 (N_21334,N_16604,N_17743);
nand U21335 (N_21335,N_19928,N_18998);
nor U21336 (N_21336,N_18691,N_18129);
and U21337 (N_21337,N_19356,N_16019);
and U21338 (N_21338,N_19358,N_19682);
xnor U21339 (N_21339,N_19019,N_15294);
nand U21340 (N_21340,N_18078,N_18123);
xor U21341 (N_21341,N_17417,N_18933);
and U21342 (N_21342,N_19738,N_19969);
and U21343 (N_21343,N_16795,N_15267);
and U21344 (N_21344,N_15008,N_15764);
or U21345 (N_21345,N_18724,N_18368);
or U21346 (N_21346,N_18230,N_19201);
xor U21347 (N_21347,N_17363,N_16911);
nor U21348 (N_21348,N_19176,N_18464);
nand U21349 (N_21349,N_18703,N_18895);
nand U21350 (N_21350,N_18176,N_17576);
nor U21351 (N_21351,N_16511,N_17298);
nand U21352 (N_21352,N_18565,N_17831);
and U21353 (N_21353,N_15273,N_15185);
nand U21354 (N_21354,N_19178,N_19212);
nand U21355 (N_21355,N_17627,N_16508);
nand U21356 (N_21356,N_19310,N_17107);
nand U21357 (N_21357,N_18522,N_15155);
nand U21358 (N_21358,N_16345,N_15648);
or U21359 (N_21359,N_18036,N_18704);
xor U21360 (N_21360,N_19609,N_19596);
nor U21361 (N_21361,N_18427,N_18612);
nor U21362 (N_21362,N_18487,N_18967);
or U21363 (N_21363,N_17102,N_16713);
nand U21364 (N_21364,N_18689,N_16959);
or U21365 (N_21365,N_16235,N_15969);
and U21366 (N_21366,N_15146,N_17083);
nand U21367 (N_21367,N_19416,N_18307);
xnor U21368 (N_21368,N_16570,N_17992);
xnor U21369 (N_21369,N_16125,N_18356);
xnor U21370 (N_21370,N_16455,N_17057);
or U21371 (N_21371,N_17082,N_16925);
and U21372 (N_21372,N_16523,N_16046);
xor U21373 (N_21373,N_15393,N_16532);
nor U21374 (N_21374,N_19333,N_19535);
nand U21375 (N_21375,N_18958,N_16771);
nor U21376 (N_21376,N_15723,N_17317);
xor U21377 (N_21377,N_15132,N_18013);
and U21378 (N_21378,N_15825,N_19641);
nand U21379 (N_21379,N_16625,N_15584);
and U21380 (N_21380,N_16678,N_18269);
nor U21381 (N_21381,N_17375,N_18188);
nor U21382 (N_21382,N_17376,N_19666);
nand U21383 (N_21383,N_17090,N_15792);
or U21384 (N_21384,N_19961,N_19181);
nand U21385 (N_21385,N_19117,N_18859);
xnor U21386 (N_21386,N_16571,N_16927);
nand U21387 (N_21387,N_16541,N_19964);
nand U21388 (N_21388,N_17342,N_19225);
or U21389 (N_21389,N_19642,N_16672);
xnor U21390 (N_21390,N_16482,N_17545);
or U21391 (N_21391,N_18365,N_15431);
xor U21392 (N_21392,N_17400,N_15079);
xor U21393 (N_21393,N_18582,N_17410);
nand U21394 (N_21394,N_15621,N_19644);
and U21395 (N_21395,N_15226,N_17158);
xnor U21396 (N_21396,N_19569,N_19727);
and U21397 (N_21397,N_18707,N_19761);
or U21398 (N_21398,N_15499,N_18019);
and U21399 (N_21399,N_15389,N_18363);
nor U21400 (N_21400,N_19202,N_18975);
or U21401 (N_21401,N_19699,N_17818);
or U21402 (N_21402,N_16655,N_15874);
and U21403 (N_21403,N_19519,N_18218);
xor U21404 (N_21404,N_18015,N_16131);
xor U21405 (N_21405,N_18845,N_17946);
nand U21406 (N_21406,N_17003,N_16965);
nand U21407 (N_21407,N_16249,N_17980);
or U21408 (N_21408,N_15630,N_19108);
or U21409 (N_21409,N_16590,N_17097);
or U21410 (N_21410,N_15866,N_15544);
nor U21411 (N_21411,N_17064,N_19691);
or U21412 (N_21412,N_19846,N_16506);
nand U21413 (N_21413,N_18906,N_19439);
nor U21414 (N_21414,N_15331,N_18735);
nand U21415 (N_21415,N_17121,N_16274);
and U21416 (N_21416,N_17273,N_17972);
and U21417 (N_21417,N_17495,N_19555);
nand U21418 (N_21418,N_15938,N_18283);
xnor U21419 (N_21419,N_18928,N_18881);
nand U21420 (N_21420,N_15691,N_18256);
nand U21421 (N_21421,N_17587,N_15174);
nor U21422 (N_21422,N_19959,N_19473);
nor U21423 (N_21423,N_16071,N_15173);
xor U21424 (N_21424,N_16148,N_17941);
nor U21425 (N_21425,N_17332,N_19237);
nand U21426 (N_21426,N_18270,N_19114);
and U21427 (N_21427,N_17226,N_17796);
nor U21428 (N_21428,N_19798,N_18417);
and U21429 (N_21429,N_17168,N_19215);
or U21430 (N_21430,N_15700,N_18187);
nand U21431 (N_21431,N_19922,N_17625);
or U21432 (N_21432,N_17676,N_16140);
xnor U21433 (N_21433,N_17153,N_18485);
nand U21434 (N_21434,N_18332,N_17561);
xnor U21435 (N_21435,N_19278,N_15711);
and U21436 (N_21436,N_18511,N_16816);
nand U21437 (N_21437,N_19828,N_15637);
nand U21438 (N_21438,N_18253,N_18448);
xnor U21439 (N_21439,N_16986,N_17096);
nor U21440 (N_21440,N_16132,N_18699);
xnor U21441 (N_21441,N_18316,N_17852);
and U21442 (N_21442,N_16465,N_17100);
nor U21443 (N_21443,N_15754,N_19167);
and U21444 (N_21444,N_16197,N_18588);
xor U21445 (N_21445,N_15303,N_19228);
nor U21446 (N_21446,N_17304,N_17235);
nand U21447 (N_21447,N_17916,N_17501);
nand U21448 (N_21448,N_15931,N_17032);
xor U21449 (N_21449,N_18222,N_18115);
nand U21450 (N_21450,N_16707,N_15254);
or U21451 (N_21451,N_19553,N_19459);
or U21452 (N_21452,N_16876,N_16910);
nand U21453 (N_21453,N_17668,N_16528);
or U21454 (N_21454,N_16821,N_15407);
or U21455 (N_21455,N_19917,N_18873);
and U21456 (N_21456,N_15746,N_19948);
xor U21457 (N_21457,N_17399,N_15152);
xor U21458 (N_21458,N_18867,N_16491);
and U21459 (N_21459,N_16385,N_19464);
nand U21460 (N_21460,N_16084,N_18265);
xnor U21461 (N_21461,N_16369,N_19707);
and U21462 (N_21462,N_16794,N_19646);
xor U21463 (N_21463,N_18341,N_15307);
xor U21464 (N_21464,N_16057,N_15879);
and U21465 (N_21465,N_18361,N_15720);
and U21466 (N_21466,N_17205,N_19427);
xor U21467 (N_21467,N_16310,N_16287);
nor U21468 (N_21468,N_17277,N_16621);
and U21469 (N_21469,N_15328,N_16341);
nand U21470 (N_21470,N_15749,N_15753);
xor U21471 (N_21471,N_17140,N_19153);
nor U21472 (N_21472,N_17156,N_16730);
or U21473 (N_21473,N_16566,N_17649);
nor U21474 (N_21474,N_16252,N_15184);
xor U21475 (N_21475,N_18432,N_18298);
or U21476 (N_21476,N_15905,N_16614);
or U21477 (N_21477,N_18545,N_16744);
xor U21478 (N_21478,N_19273,N_18130);
nor U21479 (N_21479,N_17254,N_19889);
nor U21480 (N_21480,N_15223,N_19068);
and U21481 (N_21481,N_15927,N_16550);
nor U21482 (N_21482,N_15038,N_19651);
and U21483 (N_21483,N_19845,N_17144);
nor U21484 (N_21484,N_16379,N_17824);
and U21485 (N_21485,N_15697,N_19813);
nand U21486 (N_21486,N_15416,N_19392);
nor U21487 (N_21487,N_19937,N_16975);
xnor U21488 (N_21488,N_18250,N_16463);
nand U21489 (N_21489,N_18300,N_15692);
nor U21490 (N_21490,N_18234,N_19091);
nor U21491 (N_21491,N_15500,N_15750);
nor U21492 (N_21492,N_18398,N_19027);
nor U21493 (N_21493,N_17902,N_15211);
nor U21494 (N_21494,N_15878,N_16415);
nand U21495 (N_21495,N_18733,N_16176);
nand U21496 (N_21496,N_16404,N_15840);
or U21497 (N_21497,N_18453,N_18809);
and U21498 (N_21498,N_16036,N_16185);
nand U21499 (N_21499,N_17046,N_15028);
xnor U21500 (N_21500,N_15791,N_17239);
and U21501 (N_21501,N_18258,N_15181);
xor U21502 (N_21502,N_15365,N_19880);
nand U21503 (N_21503,N_19403,N_15397);
nand U21504 (N_21504,N_18174,N_15899);
xnor U21505 (N_21505,N_17091,N_19802);
and U21506 (N_21506,N_15117,N_15632);
nor U21507 (N_21507,N_16317,N_19011);
nand U21508 (N_21508,N_16329,N_19683);
nand U21509 (N_21509,N_16796,N_16760);
nor U21510 (N_21510,N_19971,N_17435);
nand U21511 (N_21511,N_16223,N_19493);
and U21512 (N_21512,N_18052,N_17870);
nor U21513 (N_21513,N_16143,N_16214);
or U21514 (N_21514,N_15974,N_17105);
nor U21515 (N_21515,N_19381,N_19529);
and U21516 (N_21516,N_16068,N_19437);
xnor U21517 (N_21517,N_15076,N_16778);
nand U21518 (N_21518,N_15796,N_18694);
and U21519 (N_21519,N_19122,N_16108);
xnor U21520 (N_21520,N_18595,N_16997);
xor U21521 (N_21521,N_16268,N_15086);
nand U21522 (N_21522,N_19840,N_18992);
or U21523 (N_21523,N_16000,N_19189);
nor U21524 (N_21524,N_15399,N_19884);
and U21525 (N_21525,N_16174,N_15780);
xnor U21526 (N_21526,N_15210,N_16884);
or U21527 (N_21527,N_17521,N_17835);
or U21528 (N_21528,N_16180,N_16862);
xnor U21529 (N_21529,N_17892,N_17276);
and U21530 (N_21530,N_16745,N_16349);
xnor U21531 (N_21531,N_16950,N_19461);
nand U21532 (N_21532,N_18670,N_18196);
nand U21533 (N_21533,N_15016,N_18385);
and U21534 (N_21534,N_17035,N_17996);
or U21535 (N_21535,N_15955,N_17541);
nor U21536 (N_21536,N_15441,N_19357);
or U21537 (N_21537,N_16963,N_18102);
xor U21538 (N_21538,N_15625,N_17546);
or U21539 (N_21539,N_16576,N_15193);
nor U21540 (N_21540,N_17850,N_15945);
nand U21541 (N_21541,N_15920,N_19204);
nand U21542 (N_21542,N_19059,N_19843);
xor U21543 (N_21543,N_19183,N_16109);
nor U21544 (N_21544,N_17291,N_17053);
or U21545 (N_21545,N_17258,N_18407);
or U21546 (N_21546,N_17800,N_15613);
xnor U21547 (N_21547,N_18897,N_15194);
nor U21548 (N_21548,N_16377,N_17647);
or U21549 (N_21549,N_15098,N_15822);
nor U21550 (N_21550,N_18537,N_18095);
nand U21551 (N_21551,N_16995,N_15368);
nand U21552 (N_21552,N_17614,N_15506);
and U21553 (N_21553,N_16151,N_16615);
or U21554 (N_21554,N_15761,N_17540);
or U21555 (N_21555,N_18624,N_16711);
nand U21556 (N_21556,N_15276,N_17238);
nand U21557 (N_21557,N_18544,N_16996);
and U21558 (N_21558,N_18858,N_17049);
and U21559 (N_21559,N_19455,N_18568);
and U21560 (N_21560,N_17335,N_18868);
or U21561 (N_21561,N_15250,N_17358);
nand U21562 (N_21562,N_18118,N_19525);
or U21563 (N_21563,N_18392,N_17259);
nor U21564 (N_21564,N_18208,N_17509);
nor U21565 (N_21565,N_19511,N_17898);
and U21566 (N_21566,N_15464,N_19159);
nor U21567 (N_21567,N_17172,N_17160);
or U21568 (N_21568,N_19375,N_18150);
and U21569 (N_21569,N_15819,N_17652);
xnor U21570 (N_21570,N_15608,N_16510);
nor U21571 (N_21571,N_16384,N_15372);
or U21572 (N_21572,N_16724,N_17957);
xor U21573 (N_21573,N_15998,N_15557);
nand U21574 (N_21574,N_18219,N_19898);
and U21575 (N_21575,N_18903,N_17137);
or U21576 (N_21576,N_17106,N_18418);
xor U21577 (N_21577,N_19893,N_18077);
or U21578 (N_21578,N_17020,N_18935);
nand U21579 (N_21579,N_17549,N_15236);
nand U21580 (N_21580,N_15188,N_19214);
and U21581 (N_21581,N_19539,N_16440);
xor U21582 (N_21582,N_18723,N_15856);
nor U21583 (N_21583,N_15737,N_15876);
nor U21584 (N_21584,N_16120,N_18788);
nand U21585 (N_21585,N_18119,N_17885);
and U21586 (N_21586,N_16846,N_17693);
nand U21587 (N_21587,N_18113,N_15554);
and U21588 (N_21588,N_15357,N_19157);
or U21589 (N_21589,N_16087,N_18325);
nand U21590 (N_21590,N_19533,N_19471);
xor U21591 (N_21591,N_18669,N_19365);
and U21592 (N_21592,N_16598,N_18038);
and U21593 (N_21593,N_17403,N_17709);
nor U21594 (N_21594,N_16098,N_17953);
nor U21595 (N_21595,N_17355,N_18352);
xnor U21596 (N_21596,N_17669,N_17882);
nor U21597 (N_21597,N_15228,N_15962);
nor U21598 (N_21598,N_16033,N_15770);
or U21599 (N_21599,N_16686,N_15595);
nor U21600 (N_21600,N_16056,N_15803);
xnor U21601 (N_21601,N_19227,N_15398);
nand U21602 (N_21602,N_16624,N_17240);
nand U21603 (N_21603,N_18369,N_15716);
nand U21604 (N_21604,N_17600,N_17208);
and U21605 (N_21605,N_18225,N_15169);
nand U21606 (N_21606,N_16542,N_15845);
or U21607 (N_21607,N_15371,N_17441);
xor U21608 (N_21608,N_18183,N_17806);
xnor U21609 (N_21609,N_17446,N_16606);
nor U21610 (N_21610,N_18786,N_19306);
nand U21611 (N_21611,N_16459,N_18706);
nand U21612 (N_21612,N_19506,N_15145);
nand U21613 (N_21613,N_17553,N_15816);
xor U21614 (N_21614,N_19674,N_18680);
and U21615 (N_21615,N_19184,N_16258);
xnor U21616 (N_21616,N_18276,N_18740);
or U21617 (N_21617,N_15518,N_15106);
and U21618 (N_21618,N_17935,N_18456);
nand U21619 (N_21619,N_17759,N_17793);
nor U21620 (N_21620,N_16595,N_19368);
or U21621 (N_21621,N_15436,N_18030);
and U21622 (N_21622,N_15686,N_15283);
nor U21623 (N_21623,N_15248,N_19194);
nand U21624 (N_21624,N_17925,N_16340);
nor U21625 (N_21625,N_15315,N_19223);
and U21626 (N_21626,N_17571,N_18168);
nor U21627 (N_21627,N_16831,N_19242);
xor U21628 (N_21628,N_19517,N_16003);
nand U21629 (N_21629,N_17859,N_18684);
nand U21630 (N_21630,N_17518,N_17430);
xnor U21631 (N_21631,N_15550,N_15036);
nand U21632 (N_21632,N_18955,N_18450);
or U21633 (N_21633,N_16840,N_15449);
xor U21634 (N_21634,N_15077,N_17550);
and U21635 (N_21635,N_18459,N_15678);
xor U21636 (N_21636,N_16797,N_15922);
and U21637 (N_21637,N_16681,N_18075);
nor U21638 (N_21638,N_17838,N_15197);
xnor U21639 (N_21639,N_19600,N_17318);
nor U21640 (N_21640,N_19281,N_15730);
and U21641 (N_21641,N_17801,N_17255);
nor U21642 (N_21642,N_18857,N_16509);
xnor U21643 (N_21643,N_15043,N_19180);
xor U21644 (N_21644,N_17426,N_16924);
nor U21645 (N_21645,N_15166,N_19946);
and U21646 (N_21646,N_19668,N_17827);
or U21647 (N_21647,N_19582,N_18850);
xor U21648 (N_21648,N_17505,N_17081);
xor U21649 (N_21649,N_18274,N_17307);
xor U21650 (N_21650,N_17210,N_17055);
and U21651 (N_21651,N_16144,N_17392);
nand U21652 (N_21652,N_15420,N_15042);
nand U21653 (N_21653,N_17336,N_17373);
or U21654 (N_21654,N_19074,N_17798);
and U21655 (N_21655,N_18296,N_16142);
or U21656 (N_21656,N_17814,N_18803);
or U21657 (N_21657,N_15472,N_18504);
xnor U21658 (N_21658,N_16159,N_15336);
nand U21659 (N_21659,N_17574,N_19762);
or U21660 (N_21660,N_16400,N_15566);
nor U21661 (N_21661,N_15190,N_18471);
xnor U21662 (N_21662,N_15308,N_16974);
or U21663 (N_21663,N_17717,N_17577);
nor U21664 (N_21664,N_19807,N_15689);
nor U21665 (N_21665,N_17849,N_16179);
or U21666 (N_21666,N_19601,N_16364);
xor U21667 (N_21667,N_17018,N_18745);
xnor U21668 (N_21668,N_18268,N_15241);
nand U21669 (N_21669,N_16460,N_17173);
nor U21670 (N_21670,N_15726,N_16630);
and U21671 (N_21671,N_19276,N_16843);
and U21672 (N_21672,N_18426,N_18033);
nand U21673 (N_21673,N_15762,N_18271);
and U21674 (N_21674,N_18442,N_19927);
and U21675 (N_21675,N_16097,N_17569);
or U21676 (N_21676,N_18923,N_19540);
xor U21677 (N_21677,N_19685,N_15448);
and U21678 (N_21678,N_17837,N_16770);
xnor U21679 (N_21679,N_17044,N_16663);
and U21680 (N_21680,N_17761,N_17848);
nand U21681 (N_21681,N_18559,N_18091);
and U21682 (N_21682,N_17221,N_18569);
nor U21683 (N_21683,N_17679,N_17742);
and U21684 (N_21684,N_15208,N_17162);
nand U21685 (N_21685,N_17744,N_15807);
nand U21686 (N_21686,N_18424,N_18443);
nor U21687 (N_21687,N_16419,N_19363);
nor U21688 (N_21688,N_19294,N_16628);
xor U21689 (N_21689,N_18853,N_18103);
nand U21690 (N_21690,N_15108,N_19124);
xor U21691 (N_21691,N_18211,N_16882);
or U21692 (N_21692,N_17772,N_17666);
nand U21693 (N_21693,N_16344,N_18840);
nor U21694 (N_21694,N_19007,N_17535);
xnor U21695 (N_21695,N_15130,N_17296);
nor U21696 (N_21696,N_16082,N_18140);
xor U21697 (N_21697,N_15131,N_18797);
nand U21698 (N_21698,N_15082,N_17748);
nor U21699 (N_21699,N_16608,N_15668);
nand U21700 (N_21700,N_17583,N_18616);
or U21701 (N_21701,N_16673,N_15589);
nand U21702 (N_21702,N_19852,N_17178);
nor U21703 (N_21703,N_16926,N_16758);
nor U21704 (N_21704,N_17455,N_19470);
or U21705 (N_21705,N_16581,N_17183);
nor U21706 (N_21706,N_18068,N_17944);
or U21707 (N_21707,N_19106,N_17670);
nand U21708 (N_21708,N_17820,N_15238);
or U21709 (N_21709,N_15873,N_17192);
nand U21710 (N_21710,N_18224,N_18479);
xor U21711 (N_21711,N_18556,N_17382);
nor U21712 (N_21712,N_18257,N_15597);
nand U21713 (N_21713,N_17405,N_17984);
and U21714 (N_21714,N_17634,N_15403);
or U21715 (N_21715,N_18742,N_16728);
and U21716 (N_21716,N_18104,N_19162);
xor U21717 (N_21717,N_17139,N_18838);
nand U21718 (N_21718,N_15569,N_15811);
nor U21719 (N_21719,N_15908,N_16953);
and U21720 (N_21720,N_19494,N_18539);
or U21721 (N_21721,N_15568,N_18884);
or U21722 (N_21722,N_16830,N_17986);
xor U21723 (N_21723,N_17962,N_17950);
and U21724 (N_21724,N_16308,N_17547);
nor U21725 (N_21725,N_19953,N_16984);
nor U21726 (N_21726,N_18018,N_17753);
or U21727 (N_21727,N_16743,N_16293);
nor U21728 (N_21728,N_19872,N_15470);
nor U21729 (N_21729,N_15523,N_18581);
or U21730 (N_21730,N_18167,N_16406);
nand U21731 (N_21731,N_16231,N_18614);
nand U21732 (N_21732,N_17851,N_15967);
or U21733 (N_21733,N_15301,N_16007);
or U21734 (N_21734,N_15844,N_17641);
and U21735 (N_21735,N_18574,N_16425);
xor U21736 (N_21736,N_17157,N_16103);
and U21737 (N_21737,N_15820,N_15939);
nor U21738 (N_21738,N_16376,N_17488);
and U21739 (N_21739,N_16416,N_19877);
nand U21740 (N_21740,N_18116,N_15125);
and U21741 (N_21741,N_18954,N_18937);
and U21742 (N_21742,N_16644,N_16039);
nor U21743 (N_21743,N_19936,N_16640);
nand U21744 (N_21744,N_16620,N_17272);
and U21745 (N_21745,N_19466,N_19614);
nand U21746 (N_21746,N_19548,N_15543);
nor U21747 (N_21747,N_17930,N_18863);
nor U21748 (N_21748,N_19664,N_15828);
xnor U21749 (N_21749,N_18579,N_17330);
nand U21750 (N_21750,N_17189,N_15932);
xor U21751 (N_21751,N_17504,N_16337);
xor U21752 (N_21752,N_17319,N_17010);
and U21753 (N_21753,N_15386,N_15041);
xor U21754 (N_21754,N_15220,N_19974);
nor U21755 (N_21755,N_15486,N_17692);
nor U21756 (N_21756,N_17948,N_17231);
and U21757 (N_21757,N_15240,N_18648);
or U21758 (N_21758,N_16766,N_16273);
nor U21759 (N_21759,N_17943,N_17229);
xor U21760 (N_21760,N_17594,N_17416);
nor U21761 (N_21761,N_18025,N_15440);
or U21762 (N_21762,N_19505,N_19999);
nand U21763 (N_21763,N_15965,N_15601);
or U21764 (N_21764,N_17401,N_18149);
nor U21765 (N_21765,N_19541,N_19842);
and U21766 (N_21766,N_15230,N_16774);
nor U21767 (N_21767,N_18722,N_19949);
xnor U21768 (N_21768,N_15851,N_15058);
xor U21769 (N_21769,N_18625,N_19680);
and U21770 (N_21770,N_19413,N_15139);
and U21771 (N_21771,N_15558,N_17942);
and U21772 (N_21772,N_16410,N_15326);
nand U21773 (N_21773,N_15320,N_15289);
nor U21774 (N_21774,N_15348,N_19187);
xor U21775 (N_21775,N_16411,N_18636);
or U21776 (N_21776,N_17716,N_17033);
and U21777 (N_21777,N_16305,N_15610);
xnor U21778 (N_21778,N_18822,N_16479);
xor U21779 (N_21779,N_17191,N_18439);
nor U21780 (N_21780,N_19244,N_19882);
nor U21781 (N_21781,N_19731,N_16001);
nand U21782 (N_21782,N_15591,N_16448);
nor U21783 (N_21783,N_17024,N_19787);
nand U21784 (N_21784,N_17584,N_18289);
nand U21785 (N_21785,N_15972,N_18086);
or U21786 (N_21786,N_16101,N_16610);
nor U21787 (N_21787,N_18989,N_19650);
or U21788 (N_21788,N_19146,N_19280);
or U21789 (N_21789,N_19643,N_15099);
xor U21790 (N_21790,N_18633,N_18620);
nand U21791 (N_21791,N_18623,N_16723);
nor U21792 (N_21792,N_19251,N_19428);
and U21793 (N_21793,N_17282,N_15341);
xnor U21794 (N_21794,N_15748,N_18564);
and U21795 (N_21795,N_16781,N_15134);
xor U21796 (N_21796,N_19395,N_18649);
and U21797 (N_21797,N_19161,N_18088);
xnor U21798 (N_21798,N_18152,N_17124);
xor U21799 (N_21799,N_15581,N_19155);
and U21800 (N_21800,N_15128,N_19598);
nand U21801 (N_21801,N_15133,N_18372);
nand U21802 (N_21802,N_19192,N_18493);
nand U21803 (N_21803,N_17773,N_17947);
and U21804 (N_21804,N_16854,N_18096);
nor U21805 (N_21805,N_15542,N_16968);
xor U21806 (N_21806,N_16183,N_16225);
or U21807 (N_21807,N_19991,N_15204);
xnor U21808 (N_21808,N_19536,N_16545);
nor U21809 (N_21809,N_18478,N_18818);
nand U21810 (N_21810,N_16141,N_16494);
xnor U21811 (N_21811,N_18466,N_16627);
and U21812 (N_21812,N_18032,N_18644);
nand U21813 (N_21813,N_16948,N_17687);
nand U21814 (N_21814,N_15935,N_16641);
xor U21815 (N_21815,N_19383,N_19833);
xnor U21816 (N_21816,N_16263,N_19695);
xor U21817 (N_21817,N_18084,N_18632);
or U21818 (N_21818,N_19749,N_16265);
nand U21819 (N_21819,N_19042,N_15322);
xor U21820 (N_21820,N_17513,N_18667);
or U21821 (N_21821,N_17969,N_19984);
xnor U21822 (N_21822,N_16567,N_17220);
nand U21823 (N_21823,N_18700,N_16637);
and U21824 (N_21824,N_16969,N_17338);
nor U21825 (N_21825,N_16267,N_18535);
nand U21826 (N_21826,N_19549,N_18124);
or U21827 (N_21827,N_16722,N_19344);
xor U21828 (N_21828,N_18419,N_16050);
xor U21829 (N_21829,N_19116,N_19874);
xnor U21830 (N_21830,N_16922,N_16578);
nor U21831 (N_21831,N_17975,N_18278);
and U21832 (N_21832,N_17067,N_16387);
and U21833 (N_21833,N_18415,N_15855);
or U21834 (N_21834,N_18405,N_15011);
and U21835 (N_21835,N_18261,N_16555);
nor U21836 (N_21836,N_18879,N_17708);
and U21837 (N_21837,N_16696,N_18683);
or U21838 (N_21838,N_16296,N_16556);
and U21839 (N_21839,N_19542,N_18943);
nor U21840 (N_21840,N_19565,N_16059);
nor U21841 (N_21841,N_15413,N_19441);
nand U21842 (N_21842,N_19909,N_18080);
or U21843 (N_21843,N_15734,N_16271);
and U21844 (N_21844,N_18993,N_18041);
nor U21845 (N_21845,N_18981,N_18028);
xnor U21846 (N_21846,N_16546,N_18787);
or U21847 (N_21847,N_15006,N_17248);
xor U21848 (N_21848,N_18399,N_18518);
nand U21849 (N_21849,N_18861,N_19386);
or U21850 (N_21850,N_18748,N_16649);
xor U21851 (N_21851,N_16699,N_18342);
nand U21852 (N_21852,N_18805,N_17655);
nand U21853 (N_21853,N_16037,N_15418);
or U21854 (N_21854,N_18920,N_17763);
and U21855 (N_21855,N_16718,N_18490);
nand U21856 (N_21856,N_18793,N_17783);
nand U21857 (N_21857,N_18087,N_17260);
or U21858 (N_21858,N_17979,N_19101);
nand U21859 (N_21859,N_17350,N_19768);
xnor U21860 (N_21860,N_19797,N_18421);
and U21861 (N_21861,N_15526,N_15206);
or U21862 (N_21862,N_15901,N_18702);
nor U21863 (N_21863,N_18060,N_16499);
or U21864 (N_21864,N_16872,N_15171);
nand U21865 (N_21865,N_15551,N_18054);
nor U21866 (N_21866,N_15664,N_19343);
or U21867 (N_21867,N_19198,N_17642);
nor U21868 (N_21868,N_19436,N_17313);
or U21869 (N_21869,N_17077,N_16290);
xor U21870 (N_21870,N_17707,N_18286);
and U21871 (N_21871,N_17706,N_15703);
and U21872 (N_21872,N_17589,N_16666);
and U21873 (N_21873,N_19924,N_16801);
or U21874 (N_21874,N_19556,N_17381);
nor U21875 (N_21875,N_16257,N_18531);
xor U21876 (N_21876,N_15048,N_18414);
or U21877 (N_21877,N_16027,N_15616);
and U21878 (N_21878,N_17771,N_18071);
nand U21879 (N_21879,N_15930,N_15285);
or U21880 (N_21880,N_17978,N_19857);
nand U21881 (N_21881,N_19745,N_17973);
or U21882 (N_21882,N_15400,N_16501);
nor U21883 (N_21883,N_16875,N_16861);
nand U21884 (N_21884,N_17480,N_19017);
or U21885 (N_21885,N_19379,N_19941);
nand U21886 (N_21886,N_16493,N_18630);
nand U21887 (N_21887,N_16156,N_17723);
nand U21888 (N_21888,N_15665,N_16100);
nor U21889 (N_21889,N_15300,N_17864);
and U21890 (N_21890,N_18362,N_19619);
nor U21891 (N_21891,N_18741,N_17970);
or U21892 (N_21892,N_15488,N_15977);
nand U21893 (N_21893,N_17477,N_18010);
nor U21894 (N_21894,N_19728,N_15629);
xnor U21895 (N_21895,N_15247,N_18348);
nand U21896 (N_21896,N_15061,N_18425);
xnor U21897 (N_21897,N_19264,N_16124);
xor U21898 (N_21898,N_16373,N_15379);
xnor U21899 (N_21899,N_19412,N_15576);
and U21900 (N_21900,N_15921,N_16471);
nand U21901 (N_21901,N_17868,N_17906);
and U21902 (N_21902,N_19020,N_18259);
nand U21903 (N_21903,N_19916,N_17828);
and U21904 (N_21904,N_16380,N_19369);
xnor U21905 (N_21905,N_18890,N_15916);
nand U21906 (N_21906,N_19634,N_19479);
nand U21907 (N_21907,N_16938,N_15115);
or U21908 (N_21908,N_17444,N_17349);
and U21909 (N_21909,N_16889,N_17150);
xnor U21910 (N_21910,N_19573,N_19346);
and U21911 (N_21911,N_16683,N_17874);
or U21912 (N_21912,N_17266,N_18766);
nand U21913 (N_21913,N_15367,N_19033);
and U21914 (N_21914,N_16675,N_16500);
nand U21915 (N_21915,N_17608,N_15141);
nor U21916 (N_21916,N_16047,N_18575);
nand U21917 (N_21917,N_18686,N_17981);
nor U21918 (N_21918,N_19261,N_15180);
xor U21919 (N_21919,N_19662,N_19252);
nor U21920 (N_21920,N_16964,N_17875);
or U21921 (N_21921,N_19047,N_15000);
nor U21922 (N_21922,N_19763,N_16119);
or U21923 (N_21923,N_19150,N_15338);
xnor U21924 (N_21924,N_17245,N_17779);
nor U21925 (N_21925,N_16172,N_17695);
or U21926 (N_21926,N_16618,N_16382);
nor U21927 (N_21927,N_18420,N_17237);
and U21928 (N_21928,N_16354,N_17449);
nand U21929 (N_21929,N_16216,N_18619);
nor U21930 (N_21930,N_19079,N_19385);
and U21931 (N_21931,N_18371,N_19142);
or U21932 (N_21932,N_19817,N_18435);
xor U21933 (N_21933,N_19377,N_15869);
and U21934 (N_21934,N_16200,N_16487);
xor U21935 (N_21935,N_17164,N_16295);
and U21936 (N_21936,N_19070,N_17562);
nor U21937 (N_21937,N_15035,N_17632);
xnor U21938 (N_21938,N_16123,N_19060);
xor U21939 (N_21939,N_16072,N_19023);
nand U21940 (N_21940,N_15239,N_19462);
or U21941 (N_21941,N_18279,N_15638);
and U21942 (N_21942,N_17528,N_16967);
or U21943 (N_21943,N_15095,N_19747);
nor U21944 (N_21944,N_17610,N_17262);
xnor U21945 (N_21945,N_15201,N_19746);
or U21946 (N_21946,N_17479,N_16601);
nor U21947 (N_21947,N_17134,N_15066);
and U21948 (N_21948,N_17558,N_19002);
or U21949 (N_21949,N_16365,N_17346);
nand U21950 (N_21950,N_16307,N_16023);
nand U21951 (N_21951,N_15378,N_17482);
or U21952 (N_21952,N_18546,N_16860);
nand U21953 (N_21953,N_17681,N_18277);
or U21954 (N_21954,N_19777,N_19166);
xor U21955 (N_21955,N_15121,N_15102);
and U21956 (N_21956,N_16913,N_15092);
xnor U21957 (N_21957,N_17936,N_16371);
xnor U21958 (N_21958,N_16749,N_19986);
nand U21959 (N_21959,N_17867,N_18760);
and U21960 (N_21960,N_19990,N_17531);
nand U21961 (N_21961,N_15996,N_15435);
or U21962 (N_21962,N_17552,N_18982);
xor U21963 (N_21963,N_19217,N_15229);
or U21964 (N_21964,N_16093,N_18016);
and U21965 (N_21965,N_15272,N_19056);
or U21966 (N_21966,N_15148,N_18984);
nand U21967 (N_21967,N_19206,N_17174);
or U21968 (N_21968,N_19475,N_15947);
xnor U21969 (N_21969,N_17863,N_17206);
and U21970 (N_21970,N_19210,N_15979);
and U21971 (N_21971,N_15643,N_18173);
or U21972 (N_21972,N_15269,N_15354);
nand U21973 (N_21973,N_16283,N_16668);
and U21974 (N_21974,N_15560,N_15959);
and U21975 (N_21975,N_19514,N_19256);
nor U21976 (N_21976,N_19923,N_15453);
and U21977 (N_21977,N_15345,N_15424);
xor U21978 (N_21978,N_17808,N_17542);
and U21979 (N_21979,N_17387,N_17433);
xnor U21980 (N_21980,N_19253,N_18047);
nor U21981 (N_21981,N_15536,N_17414);
nor U21982 (N_21982,N_18074,N_17167);
and U21983 (N_21983,N_16850,N_18643);
nor U21984 (N_21984,N_15808,N_17580);
nand U21985 (N_21985,N_18915,N_19926);
and U21986 (N_21986,N_19089,N_18560);
and U21987 (N_21987,N_15806,N_17872);
xnor U21988 (N_21988,N_15479,N_15619);
and U21989 (N_21989,N_16116,N_18214);
and U21990 (N_21990,N_17841,N_17280);
nor U21991 (N_21991,N_15943,N_18525);
or U21992 (N_21992,N_18402,N_15968);
or U21993 (N_21993,N_18364,N_15478);
xnor U21994 (N_21994,N_19049,N_15100);
nor U21995 (N_21995,N_15805,N_15388);
and U21996 (N_21996,N_16839,N_19957);
nor U21997 (N_21997,N_16355,N_16687);
or U21998 (N_21998,N_18655,N_16521);
and U21999 (N_21999,N_15391,N_17447);
nor U22000 (N_22000,N_15429,N_19657);
xnor U22001 (N_22001,N_15183,N_15412);
and U22002 (N_22002,N_18792,N_17275);
xnor U22003 (N_22003,N_15259,N_17585);
nor U22004 (N_22004,N_18131,N_19229);
nand U22005 (N_22005,N_18037,N_15755);
nor U22006 (N_22006,N_16920,N_16219);
and U22007 (N_22007,N_16431,N_18527);
nand U22008 (N_22008,N_17448,N_15063);
xor U22009 (N_22009,N_16661,N_17630);
nor U22010 (N_22010,N_15323,N_16716);
nor U22011 (N_22011,N_16105,N_18110);
and U22012 (N_22012,N_16940,N_17177);
xor U22013 (N_22013,N_15245,N_17228);
and U22014 (N_22014,N_18008,N_19291);
or U22015 (N_22015,N_16775,N_16070);
nor U22016 (N_22016,N_17740,N_16752);
or U22017 (N_22017,N_16418,N_17395);
nand U22018 (N_22018,N_18172,N_17971);
nand U22019 (N_22019,N_16792,N_16052);
xor U22020 (N_22020,N_16660,N_16315);
nor U22021 (N_22021,N_19052,N_16905);
xnor U22022 (N_22022,N_16045,N_19804);
and U22023 (N_22023,N_16809,N_19689);
nand U22024 (N_22024,N_19336,N_15406);
xor U22025 (N_22025,N_17236,N_16702);
or U22026 (N_22026,N_18639,N_15060);
xnor U22027 (N_22027,N_15375,N_15049);
or U22028 (N_22028,N_16549,N_19121);
and U22029 (N_22029,N_16186,N_15491);
nand U22030 (N_22030,N_19544,N_18654);
and U22031 (N_22031,N_16246,N_15773);
nand U22032 (N_22032,N_18773,N_15332);
or U22033 (N_22033,N_15089,N_16452);
nor U22034 (N_22034,N_18985,N_15563);
xor U22035 (N_22035,N_16289,N_18716);
xor U22036 (N_22036,N_18547,N_18007);
or U22037 (N_22037,N_18583,N_18305);
nor U22038 (N_22038,N_15466,N_19373);
nand U22039 (N_22039,N_15885,N_17457);
nand U22040 (N_22040,N_18823,N_16657);
xnor U22041 (N_22041,N_17762,N_18968);
nor U22042 (N_22042,N_18457,N_19111);
nor U22043 (N_22043,N_15649,N_19528);
or U22044 (N_22044,N_19602,N_16768);
and U22045 (N_22045,N_18653,N_19618);
and U22046 (N_22046,N_19848,N_18238);
nand U22047 (N_22047,N_15923,N_18896);
nor U22048 (N_22048,N_19810,N_16338);
xor U22049 (N_22049,N_19396,N_15279);
or U22050 (N_22050,N_17802,N_16314);
nand U22051 (N_22051,N_18631,N_15221);
or U22052 (N_22052,N_15044,N_18815);
and U22053 (N_22053,N_16977,N_17048);
xor U22054 (N_22054,N_17876,N_17292);
nor U22055 (N_22055,N_15760,N_17062);
or U22056 (N_22056,N_15799,N_18831);
and U22057 (N_22057,N_16652,N_19894);
and U22058 (N_22058,N_19408,N_19016);
nand U22059 (N_22059,N_17698,N_16933);
nand U22060 (N_22060,N_17002,N_15302);
and U22061 (N_22061,N_16592,N_16679);
nor U22062 (N_22062,N_18922,N_15473);
and U22063 (N_22063,N_19973,N_18181);
xor U22064 (N_22064,N_18814,N_17421);
xnor U22065 (N_22065,N_17459,N_18085);
or U22066 (N_22066,N_15265,N_16847);
nor U22067 (N_22067,N_19800,N_19754);
nand U22068 (N_22068,N_18014,N_16242);
xor U22069 (N_22069,N_18908,N_17578);
nor U22070 (N_22070,N_17524,N_18965);
nand U22071 (N_22071,N_17956,N_17398);
nor U22072 (N_22072,N_16324,N_18106);
nand U22073 (N_22073,N_17767,N_16703);
or U22074 (N_22074,N_16812,N_17519);
xnor U22075 (N_22075,N_18206,N_15149);
or U22076 (N_22076,N_16573,N_15382);
nand U22077 (N_22077,N_16205,N_17597);
xor U22078 (N_22078,N_15826,N_16742);
or U22079 (N_22079,N_18338,N_15788);
or U22080 (N_22080,N_18004,N_17011);
and U22081 (N_22081,N_16928,N_18108);
or U22082 (N_22082,N_16575,N_18874);
and U22083 (N_22083,N_18128,N_17556);
xnor U22084 (N_22084,N_17458,N_15383);
xor U22085 (N_22085,N_18950,N_19378);
xor U22086 (N_22086,N_15587,N_17021);
or U22087 (N_22087,N_18573,N_18062);
xor U22088 (N_22088,N_17063,N_15349);
or U22089 (N_22089,N_15209,N_19314);
xnor U22090 (N_22090,N_17640,N_18997);
nand U22091 (N_22091,N_16210,N_18650);
xor U22092 (N_22092,N_18775,N_15202);
nand U22093 (N_22093,N_18483,N_15891);
and U22094 (N_22094,N_15369,N_15647);
or U22095 (N_22095,N_17411,N_15392);
xnor U22096 (N_22096,N_15802,N_17512);
and U22097 (N_22097,N_19858,N_19406);
and U22098 (N_22098,N_19419,N_19645);
and U22099 (N_22099,N_18813,N_17219);
or U22100 (N_22100,N_19008,N_15056);
xnor U22101 (N_22101,N_17305,N_16972);
xnor U22102 (N_22102,N_17232,N_19725);
and U22103 (N_22103,N_16403,N_18802);
nand U22104 (N_22104,N_16456,N_15717);
or U22105 (N_22105,N_19612,N_15741);
nand U22106 (N_22106,N_18570,N_19676);
xor U22107 (N_22107,N_15809,N_19307);
xnor U22108 (N_22108,N_18882,N_15774);
and U22109 (N_22109,N_17159,N_17810);
and U22110 (N_22110,N_17854,N_19165);
or U22111 (N_22111,N_15177,N_19623);
nor U22112 (N_22112,N_15284,N_16316);
or U22113 (N_22113,N_18959,N_19468);
nand U22114 (N_22114,N_18020,N_18291);
xnor U22115 (N_22115,N_15633,N_17131);
and U22116 (N_22116,N_18505,N_19431);
nor U22117 (N_22117,N_15886,N_17628);
and U22118 (N_22118,N_19743,N_19809);
xor U22119 (N_22119,N_16803,N_15381);
xor U22120 (N_22120,N_15087,N_18698);
nor U22121 (N_22121,N_17056,N_19308);
nand U22122 (N_22122,N_15052,N_16408);
and U22123 (N_22123,N_19531,N_18227);
or U22124 (N_22124,N_18367,N_17912);
nor U22125 (N_22125,N_19353,N_17784);
nor U22126 (N_22126,N_19036,N_15585);
and U22127 (N_22127,N_15030,N_17431);
xnor U22128 (N_22128,N_15503,N_15521);
or U22129 (N_22129,N_18862,N_16483);
xor U22130 (N_22130,N_19107,N_19366);
xor U22131 (N_22131,N_17356,N_17616);
xor U22132 (N_22132,N_18245,N_18877);
xor U22133 (N_22133,N_16817,N_16128);
nand U22134 (N_22134,N_17977,N_16900);
xor U22135 (N_22135,N_19417,N_17224);
or U22136 (N_22136,N_19324,N_19221);
and U22137 (N_22137,N_18697,N_16409);
or U22138 (N_22138,N_18063,N_18826);
xor U22139 (N_22139,N_18516,N_15057);
xnor U22140 (N_22140,N_15427,N_18058);
or U22141 (N_22141,N_18127,N_15850);
nand U22142 (N_22142,N_15606,N_15729);
and U22143 (N_22143,N_17739,N_15687);
nand U22144 (N_22144,N_19677,N_19684);
nor U22145 (N_22145,N_17785,N_19125);
nand U22146 (N_22146,N_16160,N_18971);
and U22147 (N_22147,N_16593,N_18765);
nor U22148 (N_22148,N_17805,N_16764);
nand U22149 (N_22149,N_18375,N_19051);
nor U22150 (N_22150,N_19818,N_18156);
nor U22151 (N_22151,N_15394,N_15426);
nand U22152 (N_22152,N_19154,N_16336);
and U22153 (N_22153,N_15706,N_19554);
or U22154 (N_22154,N_18240,N_19175);
xnor U22155 (N_22155,N_16161,N_16280);
xnor U22156 (N_22156,N_16942,N_16883);
or U22157 (N_22157,N_19191,N_19139);
nand U22158 (N_22158,N_18825,N_18508);
nor U22159 (N_22159,N_19566,N_18026);
nor U22160 (N_22160,N_18055,N_18507);
or U22161 (N_22161,N_15841,N_18373);
or U22162 (N_22162,N_15815,N_18112);
and U22163 (N_22163,N_15364,N_15511);
nor U22164 (N_22164,N_15258,N_18182);
xnor U22165 (N_22165,N_15888,N_19132);
xor U22166 (N_22166,N_19497,N_19277);
xor U22167 (N_22167,N_19410,N_15176);
nor U22168 (N_22168,N_17109,N_18820);
nor U22169 (N_22169,N_17601,N_18586);
xor U22170 (N_22170,N_19039,N_19054);
xnor U22171 (N_22171,N_16841,N_15989);
nor U22172 (N_22172,N_15794,N_17787);
or U22173 (N_22173,N_15527,N_16067);
nand U22174 (N_22174,N_16153,N_16005);
or U22175 (N_22175,N_17343,N_15504);
nand U22176 (N_22176,N_18596,N_17351);
nor U22177 (N_22177,N_16516,N_15786);
and U22178 (N_22178,N_18458,N_17383);
and U22179 (N_22179,N_18941,N_19896);
and U22180 (N_22180,N_16810,N_16514);
xor U22181 (N_22181,N_15743,N_15818);
nor U22182 (N_22182,N_15244,N_15156);
or U22183 (N_22183,N_17768,N_18790);
and U22184 (N_22184,N_16284,N_15085);
or U22185 (N_22185,N_17988,N_15614);
and U22186 (N_22186,N_17725,N_16894);
or U22187 (N_22187,N_19266,N_19939);
nor U22188 (N_22188,N_15339,N_18720);
nand U22189 (N_22189,N_16393,N_17747);
and U22190 (N_22190,N_19305,N_19524);
and U22191 (N_22191,N_16386,N_19595);
xnor U22192 (N_22192,N_17312,N_19885);
nand U22193 (N_22193,N_15172,N_17214);
or U22194 (N_22194,N_19513,N_19580);
and U22195 (N_22195,N_18849,N_18499);
nand U22196 (N_22196,N_16519,N_15854);
and U22197 (N_22197,N_16230,N_19755);
nand U22198 (N_22198,N_15911,N_16353);
nand U22199 (N_22199,N_18529,N_15681);
nor U22200 (N_22200,N_19873,N_17250);
or U22201 (N_22201,N_16656,N_17606);
or U22202 (N_22202,N_15333,N_15919);
or U22203 (N_22203,N_15126,N_16366);
or U22204 (N_22204,N_15445,N_19270);
nand U22205 (N_22205,N_18229,N_17211);
xor U22206 (N_22206,N_16126,N_15961);
nand U22207 (N_22207,N_18764,N_16198);
and U22208 (N_22208,N_18690,N_19013);
xnor U22209 (N_22209,N_18925,N_19966);
or U22210 (N_22210,N_19440,N_16445);
nor U22211 (N_22211,N_18065,N_17068);
nand U22212 (N_22212,N_15234,N_19577);
xnor U22213 (N_22213,N_19546,N_16013);
xnor U22214 (N_22214,N_16402,N_17388);
nor U22215 (N_22215,N_18590,N_19622);
and U22216 (N_22216,N_18961,N_16348);
nand U22217 (N_22217,N_19472,N_16497);
nor U22218 (N_22218,N_19349,N_15586);
xor U22219 (N_22219,N_19854,N_17812);
nand U22220 (N_22220,N_16919,N_18540);
or U22221 (N_22221,N_16956,N_19118);
or U22222 (N_22222,N_17427,N_19477);
nand U22223 (N_22223,N_17830,N_19164);
or U22224 (N_22224,N_15296,N_17357);
and U22225 (N_22225,N_17732,N_15654);
and U22226 (N_22226,N_17592,N_17694);
or U22227 (N_22227,N_16204,N_17786);
or U22228 (N_22228,N_18911,N_15516);
nand U22229 (N_22229,N_18736,N_15696);
nand U22230 (N_22230,N_15676,N_19557);
nand U22231 (N_22231,N_17619,N_16240);
or U22232 (N_22232,N_18864,N_18314);
xnor U22233 (N_22233,N_15950,N_17377);
and U22234 (N_22234,N_19084,N_17114);
xor U22235 (N_22235,N_15758,N_19709);
and U22236 (N_22236,N_18627,N_18076);
nor U22237 (N_22237,N_19585,N_16983);
nand U22238 (N_22238,N_17234,N_19372);
nor U22239 (N_22239,N_19076,N_19024);
and U22240 (N_22240,N_19788,N_17764);
or U22241 (N_22241,N_17895,N_17582);
or U22242 (N_22242,N_15005,N_17471);
or U22243 (N_22243,N_19649,N_16095);
or U22244 (N_22244,N_17465,N_18138);
xnor U22245 (N_22245,N_15437,N_17563);
and U22246 (N_22246,N_17290,N_18445);
nand U22247 (N_22247,N_15522,N_15306);
nor U22248 (N_22248,N_18842,N_18354);
and U22249 (N_22249,N_16394,N_16020);
nand U22250 (N_22250,N_17555,N_17682);
nand U22251 (N_22251,N_18996,N_18264);
and U22252 (N_22252,N_15385,N_19717);
or U22253 (N_22253,N_16701,N_17271);
or U22254 (N_22254,N_19435,N_16804);
nor U22255 (N_22255,N_15476,N_19718);
xor U22256 (N_22256,N_16170,N_19621);
or U22257 (N_22257,N_15704,N_18311);
xnor U22258 (N_22258,N_16484,N_18678);
nor U22259 (N_22259,N_19752,N_17667);
or U22260 (N_22260,N_19415,N_15083);
and U22261 (N_22261,N_16279,N_17995);
or U22262 (N_22262,N_15329,N_16407);
xor U22263 (N_22263,N_18330,N_16118);
and U22264 (N_22264,N_15640,N_16671);
and U22265 (N_22265,N_19620,N_15199);
and U22266 (N_22266,N_16441,N_18894);
xnor U22267 (N_22267,N_15870,N_18970);
xor U22268 (N_22268,N_16544,N_18936);
xnor U22269 (N_22269,N_15224,N_15631);
or U22270 (N_22270,N_16958,N_19055);
or U22271 (N_22271,N_15778,N_16522);
xnor U22272 (N_22272,N_16712,N_17396);
nor U22273 (N_22273,N_15670,N_19432);
nand U22274 (N_22274,N_19404,N_16478);
xor U22275 (N_22275,N_18584,N_16643);
nor U22276 (N_22276,N_15528,N_17202);
or U22277 (N_22277,N_15771,N_18675);
xnor U22278 (N_22278,N_18674,N_19263);
nor U22279 (N_22279,N_18870,N_15408);
and U22280 (N_22280,N_19830,N_18784);
or U22281 (N_22281,N_16079,N_18232);
nor U22282 (N_22282,N_18223,N_17123);
and U22283 (N_22283,N_17066,N_17456);
or U22284 (N_22284,N_19313,N_19733);
nand U22285 (N_22285,N_18887,N_19031);
nand U22286 (N_22286,N_15034,N_18533);
xnor U22287 (N_22287,N_19482,N_17436);
nand U22288 (N_22288,N_16548,N_19309);
nand U22289 (N_22289,N_15769,N_16852);
or U22290 (N_22290,N_18930,N_19456);
nand U22291 (N_22291,N_18555,N_19593);
nor U22292 (N_22292,N_19371,N_17629);
or U22293 (N_22293,N_17544,N_19148);
xor U22294 (N_22294,N_15865,N_18267);
nor U22295 (N_22295,N_15295,N_19639);
xnor U22296 (N_22296,N_18145,N_16032);
nand U22297 (N_22297,N_16667,N_15508);
xor U22298 (N_22298,N_18353,N_15897);
nand U22299 (N_22299,N_19867,N_16579);
or U22300 (N_22300,N_16685,N_15514);
and U22301 (N_22301,N_17246,N_16727);
nand U22302 (N_22302,N_16902,N_15970);
nand U22303 (N_22303,N_17923,N_18184);
and U22304 (N_22304,N_16946,N_17007);
or U22305 (N_22305,N_16178,N_18346);
xor U22306 (N_22306,N_16319,N_15261);
xnor U22307 (N_22307,N_15685,N_19457);
xnor U22308 (N_22308,N_16888,N_18817);
and U22309 (N_22309,N_18851,N_15310);
nor U22310 (N_22310,N_15376,N_18313);
xnor U22311 (N_22311,N_18912,N_19862);
and U22312 (N_22312,N_18956,N_17910);
and U22313 (N_22313,N_17816,N_16881);
nand U22314 (N_22314,N_15545,N_17908);
xor U22315 (N_22315,N_19334,N_19597);
and U22316 (N_22316,N_18237,N_17412);
or U22317 (N_22317,N_18774,N_15116);
and U22318 (N_22318,N_15975,N_16767);
xnor U22319 (N_22319,N_15215,N_15781);
nor U22320 (N_22320,N_15242,N_18017);
nor U22321 (N_22321,N_19382,N_16869);
and U22322 (N_22322,N_17394,N_18664);
and U22323 (N_22323,N_19853,N_16092);
xnor U22324 (N_22324,N_15981,N_15903);
xnor U22325 (N_22325,N_19568,N_16960);
nand U22326 (N_22326,N_17269,N_18513);
and U22327 (N_22327,N_15192,N_19672);
nand U22328 (N_22328,N_15031,N_19057);
or U22329 (N_22329,N_15789,N_16074);
xor U22330 (N_22330,N_17780,N_15722);
nor U22331 (N_22331,N_19496,N_15684);
xnor U22332 (N_22332,N_15444,N_16560);
xor U22333 (N_22333,N_18732,N_15877);
nand U22334 (N_22334,N_15275,N_19388);
nor U22335 (N_22335,N_15040,N_15913);
and U22336 (N_22336,N_18175,N_18994);
nor U22337 (N_22337,N_19499,N_17470);
xnor U22338 (N_22338,N_15652,N_19906);
nand U22339 (N_22339,N_19859,N_15012);
xnor U22340 (N_22340,N_17490,N_16692);
nand U22341 (N_22341,N_17529,N_15207);
or U22342 (N_22342,N_17089,N_17380);
or U22343 (N_22343,N_17887,N_17393);
nand U22344 (N_22344,N_19268,N_16868);
nand U22345 (N_22345,N_15314,N_19607);
nor U22346 (N_22346,N_18009,N_16633);
or U22347 (N_22347,N_18949,N_16121);
nand U22348 (N_22348,N_18213,N_19158);
or U22349 (N_22349,N_17605,N_16834);
or U22350 (N_22350,N_19982,N_18762);
nand U22351 (N_22351,N_16139,N_18317);
xnor U22352 (N_22352,N_17735,N_19660);
nand U22353 (N_22353,N_18273,N_15714);
xnor U22354 (N_22354,N_18848,N_15120);
xnor U22355 (N_22355,N_18141,N_15127);
or U22356 (N_22356,N_17041,N_18205);
xnor U22357 (N_22357,N_18812,N_17567);
nand U22358 (N_22358,N_16138,N_18195);
xnor U22359 (N_22359,N_15843,N_16629);
xnor U22360 (N_22360,N_15902,N_18340);
nor U22361 (N_22361,N_17494,N_17564);
nor U22362 (N_22362,N_15577,N_19348);
nand U22363 (N_22363,N_17190,N_15520);
or U22364 (N_22364,N_18477,N_16014);
and U22365 (N_22365,N_16538,N_19832);
nand U22366 (N_22366,N_16061,N_17406);
nor U22367 (N_22367,N_19759,N_17602);
nand U22368 (N_22368,N_16434,N_17127);
xnor U22369 (N_22369,N_17324,N_16887);
and U22370 (N_22370,N_18053,N_16833);
nand U22371 (N_22371,N_17736,N_16791);
nor U22372 (N_22372,N_18331,N_18578);
nor U22373 (N_22373,N_16784,N_19347);
or U22374 (N_22374,N_17611,N_17612);
nor U22375 (N_22375,N_17903,N_17656);
xnor U22376 (N_22376,N_18463,N_19498);
or U22377 (N_22377,N_16915,N_18404);
and U22378 (N_22378,N_19638,N_17701);
or U22379 (N_22379,N_15641,N_17686);
or U22380 (N_22380,N_16048,N_15501);
xor U22381 (N_22381,N_16091,N_16823);
nand U22382 (N_22382,N_19463,N_17138);
and U22383 (N_22383,N_16826,N_17323);
or U22384 (N_22384,N_19364,N_18729);
nand U22385 (N_22385,N_15617,N_17858);
nor U22386 (N_22386,N_15898,N_19097);
nand U22387 (N_22387,N_18739,N_15954);
or U22388 (N_22388,N_16611,N_18231);
nand U22389 (N_22389,N_15821,N_19246);
xor U22390 (N_22390,N_15168,N_16539);
nand U22391 (N_22391,N_15334,N_16788);
nand U22392 (N_22392,N_19043,N_19958);
xor U22393 (N_22393,N_19629,N_19321);
or U22394 (N_22394,N_19398,N_16041);
xnor U22395 (N_22395,N_19653,N_19298);
xnor U22396 (N_22396,N_19094,N_19861);
xor U22397 (N_22397,N_15775,N_16024);
nor U22398 (N_22398,N_18170,N_16971);
nand U22399 (N_22399,N_19647,N_16486);
and U22400 (N_22400,N_16361,N_19827);
xnor U22401 (N_22401,N_17809,N_15432);
or U22402 (N_22402,N_18171,N_16962);
nor U22403 (N_22403,N_16318,N_16018);
or U22404 (N_22404,N_17340,N_16111);
or U22405 (N_22405,N_17014,N_15948);
and U22406 (N_22406,N_15860,N_19944);
nor U22407 (N_22407,N_19729,N_15072);
nor U22408 (N_22408,N_18543,N_17847);
nand U22409 (N_22409,N_19912,N_16145);
or U22410 (N_22410,N_19299,N_18480);
nand U22411 (N_22411,N_15682,N_17994);
nor U22412 (N_22412,N_18705,N_19393);
nand U22413 (N_22413,N_15956,N_16725);
or U22414 (N_22414,N_18164,N_19814);
or U22415 (N_22415,N_18406,N_17145);
xor U22416 (N_22416,N_19757,N_19592);
nand U22417 (N_22417,N_17690,N_18370);
or U22418 (N_22418,N_16923,N_16181);
and U22419 (N_22419,N_18045,N_15198);
nor U22420 (N_22420,N_18799,N_19925);
nand U22421 (N_22421,N_19753,N_15555);
xnor U22422 (N_22422,N_16299,N_18470);
nor U22423 (N_22423,N_16658,N_16636);
and U22424 (N_22424,N_17776,N_17952);
xor U22425 (N_22425,N_16130,N_17579);
or U22426 (N_22426,N_15693,N_19429);
nor U22427 (N_22427,N_16603,N_15739);
and U22428 (N_22428,N_18454,N_17085);
or U22429 (N_22429,N_19688,N_17609);
nor U22430 (N_22430,N_15024,N_18297);
xor U22431 (N_22431,N_19950,N_17777);
nand U22432 (N_22432,N_17199,N_18878);
nand U22433 (N_22433,N_19700,N_19249);
and U22434 (N_22434,N_16433,N_16264);
xor U22435 (N_22435,N_19100,N_16715);
or U22436 (N_22436,N_17352,N_15452);
nand U22437 (N_22437,N_15111,N_19037);
or U22438 (N_22438,N_19006,N_15583);
or U22439 (N_22439,N_17460,N_18696);
nand U22440 (N_22440,N_15884,N_19250);
or U22441 (N_22441,N_17548,N_17661);
or U22442 (N_22442,N_18693,N_17216);
and U22443 (N_22443,N_16006,N_17877);
xnor U22444 (N_22444,N_17422,N_18272);
nand U22445 (N_22445,N_16503,N_19509);
nor U22446 (N_22446,N_18611,N_17683);
nand U22447 (N_22447,N_19345,N_16901);
or U22448 (N_22448,N_15037,N_19082);
xnor U22449 (N_22449,N_15090,N_19414);
and U22450 (N_22450,N_17474,N_16706);
or U22451 (N_22451,N_18280,N_15679);
xnor U22452 (N_22452,N_19028,N_17593);
nor U22453 (N_22453,N_18917,N_15359);
and U22454 (N_22454,N_18246,N_15010);
or U22455 (N_22455,N_16171,N_17871);
or U22456 (N_22456,N_19199,N_19098);
xnor U22457 (N_22457,N_16670,N_17613);
nor U22458 (N_22458,N_17170,N_19267);
xor U22459 (N_22459,N_18391,N_15971);
nand U22460 (N_22460,N_19837,N_17778);
or U22461 (N_22461,N_18358,N_16175);
xor U22462 (N_22462,N_18059,N_16765);
and U22463 (N_22463,N_19407,N_17581);
or U22464 (N_22464,N_18312,N_17570);
or U22465 (N_22465,N_16401,N_16038);
or U22466 (N_22466,N_18730,N_15002);
nor U22467 (N_22467,N_16829,N_16697);
or U22468 (N_22468,N_18122,N_15158);
xor U22469 (N_22469,N_19758,N_15013);
nand U22470 (N_22470,N_16648,N_18350);
xnor U22471 (N_22471,N_18051,N_16146);
nor U22472 (N_22472,N_19087,N_19130);
or U22473 (N_22473,N_15993,N_17006);
xor U22474 (N_22474,N_16976,N_16568);
nor U22475 (N_22475,N_16049,N_17792);
nor U22476 (N_22476,N_19401,N_18534);
nand U22477 (N_22477,N_15702,N_19625);
nor U22478 (N_22478,N_15266,N_18883);
and U22479 (N_22479,N_18816,N_18725);
xnor U22480 (N_22480,N_18306,N_19328);
nand U22481 (N_22481,N_19838,N_15564);
nand U22482 (N_22482,N_18757,N_19075);
and U22483 (N_22483,N_16879,N_19337);
xnor U22484 (N_22484,N_19831,N_17631);
xnor U22485 (N_22485,N_16395,N_16563);
or U22486 (N_22486,N_19604,N_15164);
xor U22487 (N_22487,N_17866,N_17689);
and U22488 (N_22488,N_19145,N_16710);
nand U22489 (N_22489,N_17128,N_19594);
nor U22490 (N_22490,N_18832,N_16654);
nand U22491 (N_22491,N_17327,N_18243);
nand U22492 (N_22492,N_15677,N_18139);
xnor U22493 (N_22493,N_17964,N_15370);
nand U22494 (N_22494,N_19993,N_18605);
nand U22495 (N_22495,N_16537,N_17013);
nand U22496 (N_22496,N_15990,N_19303);
and U22497 (N_22497,N_17253,N_15280);
and U22498 (N_22498,N_17644,N_16475);
nand U22499 (N_22499,N_18066,N_16779);
nor U22500 (N_22500,N_19316,N_19972);
nand U22501 (N_22501,N_16682,N_18673);
nor U22502 (N_22502,N_19185,N_19356);
nand U22503 (N_22503,N_15194,N_16256);
and U22504 (N_22504,N_17140,N_16982);
or U22505 (N_22505,N_19285,N_17470);
nor U22506 (N_22506,N_17422,N_18797);
and U22507 (N_22507,N_15186,N_19349);
nor U22508 (N_22508,N_19603,N_18590);
or U22509 (N_22509,N_19164,N_18025);
or U22510 (N_22510,N_16891,N_17084);
nor U22511 (N_22511,N_17449,N_19535);
nor U22512 (N_22512,N_16072,N_16810);
nor U22513 (N_22513,N_17281,N_19689);
nand U22514 (N_22514,N_19242,N_15505);
nor U22515 (N_22515,N_16540,N_19359);
xnor U22516 (N_22516,N_19659,N_17556);
or U22517 (N_22517,N_18880,N_18371);
or U22518 (N_22518,N_19034,N_15274);
xnor U22519 (N_22519,N_18644,N_18109);
nor U22520 (N_22520,N_15796,N_15918);
or U22521 (N_22521,N_18021,N_19882);
or U22522 (N_22522,N_15465,N_16590);
and U22523 (N_22523,N_15226,N_19557);
nand U22524 (N_22524,N_19151,N_18046);
or U22525 (N_22525,N_19324,N_17287);
xor U22526 (N_22526,N_18724,N_18947);
and U22527 (N_22527,N_17694,N_16901);
or U22528 (N_22528,N_19261,N_16903);
nand U22529 (N_22529,N_16441,N_15011);
nand U22530 (N_22530,N_18709,N_15653);
xor U22531 (N_22531,N_17497,N_18529);
and U22532 (N_22532,N_19891,N_18127);
nand U22533 (N_22533,N_19418,N_15987);
xnor U22534 (N_22534,N_17358,N_19968);
nand U22535 (N_22535,N_19664,N_17374);
nand U22536 (N_22536,N_18492,N_17866);
xnor U22537 (N_22537,N_18594,N_16540);
or U22538 (N_22538,N_17338,N_16524);
or U22539 (N_22539,N_19515,N_15536);
or U22540 (N_22540,N_15170,N_15839);
and U22541 (N_22541,N_17664,N_19206);
xnor U22542 (N_22542,N_17027,N_15012);
or U22543 (N_22543,N_16505,N_18008);
and U22544 (N_22544,N_18526,N_17616);
nand U22545 (N_22545,N_18118,N_17450);
or U22546 (N_22546,N_16230,N_16549);
xor U22547 (N_22547,N_17217,N_18315);
nand U22548 (N_22548,N_16962,N_18841);
nand U22549 (N_22549,N_17146,N_15682);
or U22550 (N_22550,N_17171,N_15105);
or U22551 (N_22551,N_19647,N_17486);
and U22552 (N_22552,N_17832,N_16771);
or U22553 (N_22553,N_15815,N_18871);
xor U22554 (N_22554,N_17011,N_18433);
and U22555 (N_22555,N_17000,N_18506);
nor U22556 (N_22556,N_15829,N_18808);
or U22557 (N_22557,N_18313,N_17232);
or U22558 (N_22558,N_17586,N_17030);
nor U22559 (N_22559,N_15442,N_16052);
xor U22560 (N_22560,N_16099,N_16505);
nor U22561 (N_22561,N_18190,N_19445);
or U22562 (N_22562,N_15225,N_17077);
nor U22563 (N_22563,N_18447,N_15531);
nor U22564 (N_22564,N_15264,N_16598);
or U22565 (N_22565,N_18894,N_16380);
nand U22566 (N_22566,N_18229,N_16102);
nand U22567 (N_22567,N_18391,N_17035);
or U22568 (N_22568,N_19003,N_19381);
nand U22569 (N_22569,N_16509,N_15276);
xor U22570 (N_22570,N_19697,N_18626);
nand U22571 (N_22571,N_18371,N_16793);
nand U22572 (N_22572,N_19049,N_18292);
nand U22573 (N_22573,N_15180,N_19348);
nand U22574 (N_22574,N_18405,N_18553);
xor U22575 (N_22575,N_17592,N_17291);
or U22576 (N_22576,N_16872,N_17535);
nor U22577 (N_22577,N_17867,N_16920);
xor U22578 (N_22578,N_15001,N_18550);
xnor U22579 (N_22579,N_18627,N_17030);
nand U22580 (N_22580,N_18726,N_19533);
and U22581 (N_22581,N_15673,N_15939);
nand U22582 (N_22582,N_18034,N_16448);
and U22583 (N_22583,N_16579,N_16498);
xnor U22584 (N_22584,N_16421,N_15035);
nor U22585 (N_22585,N_16068,N_17205);
or U22586 (N_22586,N_19639,N_19349);
or U22587 (N_22587,N_18971,N_19892);
and U22588 (N_22588,N_15143,N_16275);
or U22589 (N_22589,N_18211,N_18322);
or U22590 (N_22590,N_18861,N_17510);
nand U22591 (N_22591,N_19504,N_17065);
nor U22592 (N_22592,N_19263,N_16000);
nor U22593 (N_22593,N_16309,N_15460);
or U22594 (N_22594,N_16838,N_15090);
nand U22595 (N_22595,N_19503,N_19467);
nor U22596 (N_22596,N_19702,N_17017);
nand U22597 (N_22597,N_16200,N_17807);
xnor U22598 (N_22598,N_16769,N_19351);
nand U22599 (N_22599,N_16971,N_17982);
xor U22600 (N_22600,N_15972,N_17494);
nand U22601 (N_22601,N_18775,N_17824);
nor U22602 (N_22602,N_16393,N_16004);
nor U22603 (N_22603,N_19908,N_15790);
and U22604 (N_22604,N_16266,N_15538);
nand U22605 (N_22605,N_16464,N_18925);
xor U22606 (N_22606,N_18442,N_16855);
or U22607 (N_22607,N_18538,N_18704);
and U22608 (N_22608,N_16663,N_17055);
and U22609 (N_22609,N_15690,N_15148);
nand U22610 (N_22610,N_17335,N_18439);
or U22611 (N_22611,N_17246,N_16675);
or U22612 (N_22612,N_17243,N_16041);
nor U22613 (N_22613,N_15878,N_15053);
xor U22614 (N_22614,N_16745,N_18941);
nand U22615 (N_22615,N_15069,N_17385);
xnor U22616 (N_22616,N_16230,N_17643);
xor U22617 (N_22617,N_18701,N_18518);
nand U22618 (N_22618,N_16579,N_19040);
xor U22619 (N_22619,N_19696,N_19481);
and U22620 (N_22620,N_17528,N_17393);
nand U22621 (N_22621,N_15331,N_19827);
xor U22622 (N_22622,N_15989,N_15132);
nor U22623 (N_22623,N_17805,N_15743);
and U22624 (N_22624,N_19631,N_16448);
xnor U22625 (N_22625,N_15528,N_16303);
nand U22626 (N_22626,N_16793,N_17157);
and U22627 (N_22627,N_16521,N_15350);
or U22628 (N_22628,N_16915,N_18414);
and U22629 (N_22629,N_15372,N_18104);
nand U22630 (N_22630,N_19729,N_18088);
xor U22631 (N_22631,N_16475,N_18311);
and U22632 (N_22632,N_16829,N_16526);
and U22633 (N_22633,N_17780,N_17084);
or U22634 (N_22634,N_15422,N_15635);
or U22635 (N_22635,N_17275,N_18047);
or U22636 (N_22636,N_19045,N_17916);
nand U22637 (N_22637,N_16660,N_18331);
or U22638 (N_22638,N_17396,N_18597);
and U22639 (N_22639,N_18865,N_15362);
nand U22640 (N_22640,N_17011,N_19234);
xor U22641 (N_22641,N_19843,N_18050);
or U22642 (N_22642,N_15311,N_18720);
and U22643 (N_22643,N_15776,N_16466);
xor U22644 (N_22644,N_18010,N_19105);
and U22645 (N_22645,N_19576,N_18977);
xor U22646 (N_22646,N_15271,N_17339);
xor U22647 (N_22647,N_15931,N_19601);
or U22648 (N_22648,N_17798,N_15873);
nor U22649 (N_22649,N_15374,N_16142);
and U22650 (N_22650,N_18702,N_18024);
nand U22651 (N_22651,N_15020,N_16130);
or U22652 (N_22652,N_16405,N_19793);
xor U22653 (N_22653,N_19240,N_19214);
nor U22654 (N_22654,N_15934,N_17415);
nand U22655 (N_22655,N_18735,N_16044);
or U22656 (N_22656,N_16317,N_19172);
or U22657 (N_22657,N_15863,N_19792);
nand U22658 (N_22658,N_18785,N_19941);
xor U22659 (N_22659,N_15799,N_17145);
nand U22660 (N_22660,N_19425,N_15379);
or U22661 (N_22661,N_16944,N_18965);
or U22662 (N_22662,N_17104,N_18863);
nor U22663 (N_22663,N_17334,N_17946);
nor U22664 (N_22664,N_17834,N_17019);
xor U22665 (N_22665,N_15736,N_17663);
or U22666 (N_22666,N_17871,N_15842);
nand U22667 (N_22667,N_17226,N_18599);
xnor U22668 (N_22668,N_16616,N_15305);
nor U22669 (N_22669,N_16190,N_17430);
nand U22670 (N_22670,N_17513,N_16838);
and U22671 (N_22671,N_18881,N_15883);
or U22672 (N_22672,N_17995,N_17478);
nand U22673 (N_22673,N_18834,N_17821);
nor U22674 (N_22674,N_16013,N_17027);
xnor U22675 (N_22675,N_16235,N_18180);
nor U22676 (N_22676,N_18259,N_16420);
and U22677 (N_22677,N_16872,N_18079);
nor U22678 (N_22678,N_15693,N_16589);
or U22679 (N_22679,N_18018,N_17968);
or U22680 (N_22680,N_19093,N_19514);
xor U22681 (N_22681,N_17952,N_17187);
nand U22682 (N_22682,N_17627,N_19908);
nor U22683 (N_22683,N_16837,N_17653);
nand U22684 (N_22684,N_15584,N_19468);
nand U22685 (N_22685,N_19967,N_19538);
xor U22686 (N_22686,N_19227,N_19189);
nor U22687 (N_22687,N_19141,N_17862);
nand U22688 (N_22688,N_18057,N_18935);
nor U22689 (N_22689,N_15616,N_18866);
xnor U22690 (N_22690,N_16540,N_18320);
nor U22691 (N_22691,N_17493,N_15741);
or U22692 (N_22692,N_17253,N_16998);
nand U22693 (N_22693,N_18691,N_16153);
and U22694 (N_22694,N_16098,N_16819);
xor U22695 (N_22695,N_15990,N_18603);
nand U22696 (N_22696,N_19704,N_19492);
xor U22697 (N_22697,N_17350,N_15918);
or U22698 (N_22698,N_15571,N_17147);
and U22699 (N_22699,N_16628,N_19008);
nor U22700 (N_22700,N_17607,N_17275);
and U22701 (N_22701,N_15764,N_16907);
or U22702 (N_22702,N_19552,N_19644);
nand U22703 (N_22703,N_18580,N_17424);
or U22704 (N_22704,N_16805,N_15526);
nor U22705 (N_22705,N_15860,N_18072);
nand U22706 (N_22706,N_18372,N_15754);
or U22707 (N_22707,N_15689,N_15736);
nor U22708 (N_22708,N_18147,N_18978);
and U22709 (N_22709,N_16272,N_17720);
and U22710 (N_22710,N_17157,N_17912);
nand U22711 (N_22711,N_18480,N_15826);
and U22712 (N_22712,N_16276,N_19158);
nor U22713 (N_22713,N_16636,N_17184);
and U22714 (N_22714,N_19399,N_16032);
xor U22715 (N_22715,N_15618,N_18979);
nand U22716 (N_22716,N_15752,N_16155);
xnor U22717 (N_22717,N_17177,N_17345);
xnor U22718 (N_22718,N_16189,N_18676);
or U22719 (N_22719,N_19027,N_18834);
nor U22720 (N_22720,N_18356,N_17064);
or U22721 (N_22721,N_17908,N_15533);
xnor U22722 (N_22722,N_15218,N_19441);
xnor U22723 (N_22723,N_15843,N_17540);
and U22724 (N_22724,N_16561,N_18564);
nor U22725 (N_22725,N_18929,N_16822);
xnor U22726 (N_22726,N_16600,N_18649);
and U22727 (N_22727,N_18384,N_15871);
or U22728 (N_22728,N_17431,N_16114);
xor U22729 (N_22729,N_17759,N_18037);
and U22730 (N_22730,N_19559,N_16960);
or U22731 (N_22731,N_19552,N_16235);
nand U22732 (N_22732,N_16049,N_16606);
or U22733 (N_22733,N_18959,N_15086);
and U22734 (N_22734,N_18329,N_15881);
xor U22735 (N_22735,N_18261,N_15440);
nor U22736 (N_22736,N_17839,N_19781);
nor U22737 (N_22737,N_16369,N_19134);
nor U22738 (N_22738,N_18377,N_19567);
xor U22739 (N_22739,N_17272,N_18997);
nor U22740 (N_22740,N_17471,N_19714);
or U22741 (N_22741,N_19835,N_19424);
nand U22742 (N_22742,N_17681,N_15322);
and U22743 (N_22743,N_19410,N_18604);
nand U22744 (N_22744,N_16519,N_16466);
nand U22745 (N_22745,N_15607,N_17699);
nand U22746 (N_22746,N_18646,N_18752);
xnor U22747 (N_22747,N_18879,N_17944);
and U22748 (N_22748,N_17953,N_17284);
nor U22749 (N_22749,N_18890,N_18041);
nor U22750 (N_22750,N_17214,N_16640);
or U22751 (N_22751,N_18389,N_17747);
xnor U22752 (N_22752,N_16653,N_17038);
nor U22753 (N_22753,N_15296,N_16721);
nor U22754 (N_22754,N_15794,N_18291);
xor U22755 (N_22755,N_19564,N_16850);
nor U22756 (N_22756,N_18789,N_19822);
or U22757 (N_22757,N_18450,N_18220);
or U22758 (N_22758,N_18043,N_15317);
or U22759 (N_22759,N_15499,N_15478);
or U22760 (N_22760,N_18415,N_19805);
and U22761 (N_22761,N_18797,N_15755);
xnor U22762 (N_22762,N_16266,N_15288);
xnor U22763 (N_22763,N_19992,N_17443);
nand U22764 (N_22764,N_15338,N_15979);
nand U22765 (N_22765,N_19861,N_17641);
nand U22766 (N_22766,N_16786,N_16745);
xnor U22767 (N_22767,N_19455,N_15334);
or U22768 (N_22768,N_17017,N_16245);
xor U22769 (N_22769,N_18121,N_16784);
nor U22770 (N_22770,N_17985,N_19614);
and U22771 (N_22771,N_15126,N_16007);
or U22772 (N_22772,N_17908,N_17243);
nand U22773 (N_22773,N_15063,N_15944);
nand U22774 (N_22774,N_15748,N_16320);
or U22775 (N_22775,N_15073,N_19937);
or U22776 (N_22776,N_16899,N_17107);
and U22777 (N_22777,N_15456,N_15559);
or U22778 (N_22778,N_19239,N_15453);
nand U22779 (N_22779,N_19775,N_17923);
xor U22780 (N_22780,N_15883,N_19800);
and U22781 (N_22781,N_15733,N_19377);
or U22782 (N_22782,N_17974,N_19081);
or U22783 (N_22783,N_17206,N_17613);
xor U22784 (N_22784,N_15284,N_19185);
and U22785 (N_22785,N_18873,N_18244);
nand U22786 (N_22786,N_18605,N_19127);
nor U22787 (N_22787,N_18119,N_16793);
or U22788 (N_22788,N_17017,N_18007);
nor U22789 (N_22789,N_17854,N_17684);
and U22790 (N_22790,N_18219,N_17222);
nand U22791 (N_22791,N_19595,N_16171);
or U22792 (N_22792,N_15736,N_16133);
nand U22793 (N_22793,N_18184,N_16711);
nand U22794 (N_22794,N_15117,N_18637);
or U22795 (N_22795,N_16103,N_18820);
and U22796 (N_22796,N_17645,N_19531);
xor U22797 (N_22797,N_17666,N_18924);
nor U22798 (N_22798,N_18339,N_19080);
xor U22799 (N_22799,N_17444,N_16559);
and U22800 (N_22800,N_15152,N_15150);
nor U22801 (N_22801,N_18967,N_19266);
xnor U22802 (N_22802,N_18328,N_17531);
nor U22803 (N_22803,N_18810,N_16068);
xor U22804 (N_22804,N_15485,N_18436);
nor U22805 (N_22805,N_19070,N_15440);
or U22806 (N_22806,N_15723,N_19753);
nor U22807 (N_22807,N_16515,N_19694);
and U22808 (N_22808,N_17234,N_16524);
and U22809 (N_22809,N_18132,N_18161);
and U22810 (N_22810,N_16476,N_18909);
nor U22811 (N_22811,N_18791,N_17362);
nor U22812 (N_22812,N_18590,N_15277);
xnor U22813 (N_22813,N_15072,N_18678);
and U22814 (N_22814,N_17147,N_16469);
nor U22815 (N_22815,N_15444,N_19147);
or U22816 (N_22816,N_16779,N_16634);
or U22817 (N_22817,N_15037,N_19441);
or U22818 (N_22818,N_16203,N_18483);
nand U22819 (N_22819,N_18103,N_18877);
nor U22820 (N_22820,N_19543,N_16487);
and U22821 (N_22821,N_16564,N_17548);
and U22822 (N_22822,N_19211,N_16189);
nand U22823 (N_22823,N_19355,N_16497);
and U22824 (N_22824,N_17003,N_19777);
xnor U22825 (N_22825,N_19103,N_17808);
nand U22826 (N_22826,N_19091,N_15750);
nand U22827 (N_22827,N_19846,N_18060);
nand U22828 (N_22828,N_17634,N_15719);
xnor U22829 (N_22829,N_17636,N_17624);
xnor U22830 (N_22830,N_16688,N_15093);
nor U22831 (N_22831,N_18193,N_15236);
and U22832 (N_22832,N_17530,N_16510);
xnor U22833 (N_22833,N_19782,N_16619);
nor U22834 (N_22834,N_19574,N_18595);
xnor U22835 (N_22835,N_19688,N_15153);
and U22836 (N_22836,N_15998,N_17582);
or U22837 (N_22837,N_19032,N_19419);
nand U22838 (N_22838,N_18730,N_18981);
and U22839 (N_22839,N_18942,N_18036);
and U22840 (N_22840,N_19525,N_17459);
xnor U22841 (N_22841,N_15886,N_16800);
nand U22842 (N_22842,N_15866,N_17762);
or U22843 (N_22843,N_16395,N_15065);
nor U22844 (N_22844,N_15163,N_17191);
and U22845 (N_22845,N_16800,N_15829);
nand U22846 (N_22846,N_16701,N_19450);
xnor U22847 (N_22847,N_15732,N_15059);
nor U22848 (N_22848,N_15616,N_17874);
and U22849 (N_22849,N_19878,N_17401);
nand U22850 (N_22850,N_17905,N_17338);
and U22851 (N_22851,N_18907,N_17053);
nor U22852 (N_22852,N_15351,N_15237);
or U22853 (N_22853,N_17788,N_18469);
and U22854 (N_22854,N_19216,N_18640);
nor U22855 (N_22855,N_18174,N_19153);
nor U22856 (N_22856,N_18441,N_17725);
nand U22857 (N_22857,N_16349,N_16437);
or U22858 (N_22858,N_16854,N_19240);
and U22859 (N_22859,N_16373,N_18753);
xor U22860 (N_22860,N_16311,N_17912);
nand U22861 (N_22861,N_16226,N_18543);
nand U22862 (N_22862,N_17018,N_18728);
xor U22863 (N_22863,N_16748,N_16699);
xor U22864 (N_22864,N_18001,N_15897);
or U22865 (N_22865,N_18666,N_19372);
nor U22866 (N_22866,N_17444,N_15333);
xnor U22867 (N_22867,N_15042,N_16591);
nor U22868 (N_22868,N_18505,N_16325);
nor U22869 (N_22869,N_15950,N_18155);
and U22870 (N_22870,N_18236,N_17467);
nor U22871 (N_22871,N_17002,N_17819);
or U22872 (N_22872,N_18467,N_18872);
nor U22873 (N_22873,N_17641,N_18460);
nor U22874 (N_22874,N_17693,N_17448);
xnor U22875 (N_22875,N_18751,N_18859);
or U22876 (N_22876,N_15699,N_17507);
nor U22877 (N_22877,N_15057,N_15127);
nor U22878 (N_22878,N_18699,N_17567);
nor U22879 (N_22879,N_18958,N_15334);
nand U22880 (N_22880,N_17472,N_19192);
xnor U22881 (N_22881,N_17097,N_17211);
xnor U22882 (N_22882,N_16456,N_18434);
or U22883 (N_22883,N_15114,N_15651);
nand U22884 (N_22884,N_15342,N_16412);
nor U22885 (N_22885,N_15566,N_15726);
and U22886 (N_22886,N_18786,N_16575);
nor U22887 (N_22887,N_15834,N_16952);
nor U22888 (N_22888,N_18234,N_19060);
or U22889 (N_22889,N_17358,N_19316);
nor U22890 (N_22890,N_18489,N_19039);
xnor U22891 (N_22891,N_18174,N_16838);
xor U22892 (N_22892,N_18804,N_19386);
and U22893 (N_22893,N_17740,N_17234);
and U22894 (N_22894,N_18521,N_19734);
or U22895 (N_22895,N_19573,N_15147);
or U22896 (N_22896,N_17398,N_15005);
xor U22897 (N_22897,N_17371,N_18049);
or U22898 (N_22898,N_19727,N_19882);
nand U22899 (N_22899,N_16237,N_19633);
nand U22900 (N_22900,N_16733,N_17981);
nand U22901 (N_22901,N_19764,N_16641);
or U22902 (N_22902,N_15699,N_16686);
nor U22903 (N_22903,N_18883,N_19021);
xor U22904 (N_22904,N_17706,N_15219);
or U22905 (N_22905,N_18598,N_15188);
xnor U22906 (N_22906,N_15331,N_18308);
or U22907 (N_22907,N_18163,N_19314);
or U22908 (N_22908,N_17141,N_19434);
and U22909 (N_22909,N_16870,N_19646);
xor U22910 (N_22910,N_16392,N_16568);
xor U22911 (N_22911,N_16312,N_15864);
nand U22912 (N_22912,N_17338,N_17138);
or U22913 (N_22913,N_19812,N_19400);
and U22914 (N_22914,N_15712,N_16738);
nand U22915 (N_22915,N_16981,N_15156);
nand U22916 (N_22916,N_18849,N_18241);
nand U22917 (N_22917,N_17379,N_15148);
and U22918 (N_22918,N_18848,N_18052);
nor U22919 (N_22919,N_16015,N_19388);
and U22920 (N_22920,N_17522,N_17119);
or U22921 (N_22921,N_18476,N_19956);
xor U22922 (N_22922,N_19498,N_17228);
nand U22923 (N_22923,N_15805,N_18762);
xor U22924 (N_22924,N_15427,N_17991);
nand U22925 (N_22925,N_15844,N_17816);
or U22926 (N_22926,N_19354,N_18374);
xnor U22927 (N_22927,N_16811,N_19586);
xor U22928 (N_22928,N_16002,N_18178);
nand U22929 (N_22929,N_19617,N_16972);
xnor U22930 (N_22930,N_15326,N_18781);
xnor U22931 (N_22931,N_16440,N_16003);
xor U22932 (N_22932,N_15929,N_18900);
and U22933 (N_22933,N_19368,N_18815);
xnor U22934 (N_22934,N_18708,N_18253);
xnor U22935 (N_22935,N_15947,N_19987);
and U22936 (N_22936,N_17051,N_19320);
nor U22937 (N_22937,N_15665,N_16388);
nor U22938 (N_22938,N_17959,N_15119);
xor U22939 (N_22939,N_17082,N_15785);
and U22940 (N_22940,N_15826,N_19059);
and U22941 (N_22941,N_18250,N_17733);
or U22942 (N_22942,N_17757,N_19348);
nand U22943 (N_22943,N_19866,N_19127);
nor U22944 (N_22944,N_16759,N_17825);
xor U22945 (N_22945,N_19314,N_16495);
or U22946 (N_22946,N_16271,N_19249);
nor U22947 (N_22947,N_18436,N_18267);
nand U22948 (N_22948,N_18479,N_19282);
nor U22949 (N_22949,N_17433,N_15754);
nand U22950 (N_22950,N_17177,N_17602);
nor U22951 (N_22951,N_17561,N_17611);
or U22952 (N_22952,N_16750,N_17116);
or U22953 (N_22953,N_15805,N_18539);
and U22954 (N_22954,N_17554,N_17518);
nand U22955 (N_22955,N_18294,N_18073);
xnor U22956 (N_22956,N_19235,N_17044);
and U22957 (N_22957,N_15809,N_18506);
nand U22958 (N_22958,N_18525,N_17173);
and U22959 (N_22959,N_15586,N_17609);
nand U22960 (N_22960,N_15330,N_18862);
xnor U22961 (N_22961,N_17885,N_17641);
xor U22962 (N_22962,N_15182,N_17589);
nand U22963 (N_22963,N_16875,N_15104);
and U22964 (N_22964,N_15733,N_15852);
and U22965 (N_22965,N_15960,N_16436);
xor U22966 (N_22966,N_18351,N_17657);
nor U22967 (N_22967,N_15096,N_17372);
nor U22968 (N_22968,N_16241,N_16019);
nand U22969 (N_22969,N_18764,N_16312);
nand U22970 (N_22970,N_16277,N_19810);
nor U22971 (N_22971,N_17388,N_18600);
or U22972 (N_22972,N_19862,N_18678);
nor U22973 (N_22973,N_17683,N_18766);
xor U22974 (N_22974,N_17734,N_15845);
and U22975 (N_22975,N_19715,N_19033);
nand U22976 (N_22976,N_18692,N_19855);
and U22977 (N_22977,N_17601,N_17162);
nor U22978 (N_22978,N_18384,N_19770);
xor U22979 (N_22979,N_15075,N_19710);
nor U22980 (N_22980,N_18406,N_18706);
or U22981 (N_22981,N_18227,N_15471);
xor U22982 (N_22982,N_18580,N_16040);
or U22983 (N_22983,N_17831,N_16297);
nand U22984 (N_22984,N_17211,N_19052);
and U22985 (N_22985,N_16190,N_15888);
or U22986 (N_22986,N_18505,N_19605);
nand U22987 (N_22987,N_15786,N_18147);
xnor U22988 (N_22988,N_18191,N_16131);
nand U22989 (N_22989,N_19501,N_18062);
nor U22990 (N_22990,N_19071,N_17184);
nand U22991 (N_22991,N_16382,N_16741);
and U22992 (N_22992,N_17905,N_17200);
or U22993 (N_22993,N_16433,N_18755);
nor U22994 (N_22994,N_18950,N_18848);
or U22995 (N_22995,N_18122,N_18279);
nor U22996 (N_22996,N_15605,N_18141);
xnor U22997 (N_22997,N_16450,N_17665);
xor U22998 (N_22998,N_15617,N_17686);
and U22999 (N_22999,N_17564,N_17574);
and U23000 (N_23000,N_17862,N_16723);
or U23001 (N_23001,N_18825,N_17944);
xnor U23002 (N_23002,N_18443,N_16715);
or U23003 (N_23003,N_16001,N_19299);
and U23004 (N_23004,N_15094,N_18167);
nor U23005 (N_23005,N_17932,N_15990);
or U23006 (N_23006,N_16959,N_18605);
xnor U23007 (N_23007,N_19597,N_17180);
and U23008 (N_23008,N_17100,N_17064);
and U23009 (N_23009,N_18603,N_17090);
nor U23010 (N_23010,N_19544,N_17371);
or U23011 (N_23011,N_15993,N_15412);
nor U23012 (N_23012,N_16667,N_18236);
or U23013 (N_23013,N_19531,N_15544);
and U23014 (N_23014,N_17830,N_19078);
or U23015 (N_23015,N_18588,N_18128);
nand U23016 (N_23016,N_19654,N_17268);
or U23017 (N_23017,N_17480,N_16326);
nand U23018 (N_23018,N_19083,N_19641);
or U23019 (N_23019,N_19682,N_18853);
xnor U23020 (N_23020,N_19528,N_19111);
nor U23021 (N_23021,N_15416,N_18862);
nand U23022 (N_23022,N_18970,N_16153);
nand U23023 (N_23023,N_19527,N_19568);
nor U23024 (N_23024,N_17234,N_16130);
and U23025 (N_23025,N_16710,N_16055);
nand U23026 (N_23026,N_18976,N_16090);
and U23027 (N_23027,N_16558,N_15618);
and U23028 (N_23028,N_19564,N_16872);
and U23029 (N_23029,N_15352,N_17052);
and U23030 (N_23030,N_16103,N_18185);
nor U23031 (N_23031,N_17085,N_17683);
or U23032 (N_23032,N_17022,N_16447);
or U23033 (N_23033,N_16229,N_18550);
xnor U23034 (N_23034,N_17862,N_17588);
xnor U23035 (N_23035,N_17156,N_17448);
nand U23036 (N_23036,N_17556,N_18832);
nor U23037 (N_23037,N_19779,N_15580);
xor U23038 (N_23038,N_17581,N_17946);
xor U23039 (N_23039,N_17647,N_18107);
or U23040 (N_23040,N_16279,N_17766);
and U23041 (N_23041,N_18415,N_18359);
xnor U23042 (N_23042,N_18870,N_18495);
nand U23043 (N_23043,N_19665,N_16592);
xor U23044 (N_23044,N_15133,N_19682);
nor U23045 (N_23045,N_18470,N_16465);
or U23046 (N_23046,N_18872,N_15689);
nand U23047 (N_23047,N_19209,N_16928);
nand U23048 (N_23048,N_18986,N_15194);
nand U23049 (N_23049,N_16760,N_16978);
xnor U23050 (N_23050,N_16118,N_15187);
nor U23051 (N_23051,N_16458,N_17843);
and U23052 (N_23052,N_19013,N_18886);
nand U23053 (N_23053,N_17213,N_15118);
and U23054 (N_23054,N_17832,N_16248);
or U23055 (N_23055,N_18853,N_16184);
and U23056 (N_23056,N_18420,N_16610);
or U23057 (N_23057,N_15886,N_18017);
and U23058 (N_23058,N_19170,N_15099);
nor U23059 (N_23059,N_15727,N_16695);
and U23060 (N_23060,N_16160,N_15955);
xnor U23061 (N_23061,N_17188,N_16954);
xor U23062 (N_23062,N_16129,N_19536);
nor U23063 (N_23063,N_16204,N_18374);
and U23064 (N_23064,N_19079,N_15101);
or U23065 (N_23065,N_15293,N_18410);
xnor U23066 (N_23066,N_19630,N_16093);
nand U23067 (N_23067,N_15501,N_15376);
and U23068 (N_23068,N_16431,N_15762);
and U23069 (N_23069,N_19396,N_16220);
nor U23070 (N_23070,N_19232,N_18868);
and U23071 (N_23071,N_18114,N_19763);
nand U23072 (N_23072,N_17270,N_16238);
xnor U23073 (N_23073,N_18819,N_19495);
and U23074 (N_23074,N_17771,N_15656);
xnor U23075 (N_23075,N_19775,N_18104);
and U23076 (N_23076,N_15401,N_17882);
nand U23077 (N_23077,N_16681,N_19172);
nand U23078 (N_23078,N_15242,N_18148);
xnor U23079 (N_23079,N_15967,N_15879);
xor U23080 (N_23080,N_15875,N_19544);
nor U23081 (N_23081,N_18031,N_15286);
xnor U23082 (N_23082,N_16265,N_15576);
nand U23083 (N_23083,N_19520,N_15826);
and U23084 (N_23084,N_17813,N_19272);
nor U23085 (N_23085,N_18028,N_15865);
nor U23086 (N_23086,N_17352,N_15141);
nor U23087 (N_23087,N_18671,N_15408);
or U23088 (N_23088,N_18196,N_17322);
xnor U23089 (N_23089,N_15051,N_19070);
nand U23090 (N_23090,N_18117,N_15643);
and U23091 (N_23091,N_18503,N_17413);
or U23092 (N_23092,N_16380,N_17569);
or U23093 (N_23093,N_19507,N_19137);
xnor U23094 (N_23094,N_16138,N_15483);
or U23095 (N_23095,N_18273,N_17604);
or U23096 (N_23096,N_16294,N_19658);
xnor U23097 (N_23097,N_19095,N_19515);
nand U23098 (N_23098,N_18901,N_17046);
xnor U23099 (N_23099,N_19634,N_17103);
nand U23100 (N_23100,N_15323,N_18453);
and U23101 (N_23101,N_17110,N_16994);
and U23102 (N_23102,N_18632,N_19778);
xnor U23103 (N_23103,N_18163,N_15589);
nor U23104 (N_23104,N_16932,N_15623);
and U23105 (N_23105,N_18146,N_19813);
nor U23106 (N_23106,N_19366,N_16937);
and U23107 (N_23107,N_16938,N_16421);
and U23108 (N_23108,N_18032,N_15004);
nand U23109 (N_23109,N_19766,N_15211);
xor U23110 (N_23110,N_18435,N_19839);
nand U23111 (N_23111,N_15275,N_18643);
nor U23112 (N_23112,N_16376,N_18746);
nor U23113 (N_23113,N_16696,N_15490);
nor U23114 (N_23114,N_17066,N_15641);
or U23115 (N_23115,N_15505,N_16373);
nor U23116 (N_23116,N_16464,N_17130);
xor U23117 (N_23117,N_19179,N_17624);
nand U23118 (N_23118,N_17728,N_15289);
nor U23119 (N_23119,N_16415,N_15723);
nor U23120 (N_23120,N_15989,N_18581);
nor U23121 (N_23121,N_16924,N_17437);
xor U23122 (N_23122,N_18560,N_17868);
nor U23123 (N_23123,N_17886,N_15888);
or U23124 (N_23124,N_19691,N_18741);
and U23125 (N_23125,N_17851,N_15438);
nand U23126 (N_23126,N_15660,N_19816);
or U23127 (N_23127,N_16973,N_19670);
xnor U23128 (N_23128,N_19739,N_16093);
xnor U23129 (N_23129,N_16736,N_16319);
or U23130 (N_23130,N_15685,N_15181);
or U23131 (N_23131,N_16132,N_18295);
nor U23132 (N_23132,N_18829,N_15740);
and U23133 (N_23133,N_18850,N_18569);
nand U23134 (N_23134,N_16208,N_15215);
nand U23135 (N_23135,N_16611,N_15925);
nor U23136 (N_23136,N_18687,N_15447);
nor U23137 (N_23137,N_15596,N_16122);
and U23138 (N_23138,N_18692,N_15050);
nand U23139 (N_23139,N_15325,N_17935);
or U23140 (N_23140,N_17158,N_15955);
nor U23141 (N_23141,N_16728,N_16069);
xnor U23142 (N_23142,N_17276,N_18885);
or U23143 (N_23143,N_19094,N_19047);
xor U23144 (N_23144,N_16819,N_15386);
xor U23145 (N_23145,N_17601,N_15329);
and U23146 (N_23146,N_18705,N_16743);
or U23147 (N_23147,N_16938,N_19675);
xor U23148 (N_23148,N_18145,N_16354);
nand U23149 (N_23149,N_17428,N_19760);
and U23150 (N_23150,N_15827,N_18610);
nand U23151 (N_23151,N_19458,N_18084);
and U23152 (N_23152,N_16992,N_18005);
nand U23153 (N_23153,N_18952,N_15118);
or U23154 (N_23154,N_15441,N_17775);
and U23155 (N_23155,N_17193,N_18242);
nand U23156 (N_23156,N_16549,N_15319);
and U23157 (N_23157,N_17774,N_15126);
nand U23158 (N_23158,N_19338,N_17156);
and U23159 (N_23159,N_15193,N_16808);
nand U23160 (N_23160,N_19757,N_17442);
nand U23161 (N_23161,N_18489,N_18491);
and U23162 (N_23162,N_15133,N_17605);
xor U23163 (N_23163,N_18630,N_15935);
xnor U23164 (N_23164,N_15561,N_17971);
and U23165 (N_23165,N_19862,N_15817);
nand U23166 (N_23166,N_18333,N_18445);
and U23167 (N_23167,N_18747,N_19202);
or U23168 (N_23168,N_15364,N_19152);
xor U23169 (N_23169,N_15783,N_18428);
and U23170 (N_23170,N_16039,N_16007);
nand U23171 (N_23171,N_15808,N_17355);
nor U23172 (N_23172,N_19730,N_19851);
nand U23173 (N_23173,N_17945,N_16343);
or U23174 (N_23174,N_19437,N_15113);
or U23175 (N_23175,N_17929,N_19582);
or U23176 (N_23176,N_17573,N_18189);
and U23177 (N_23177,N_16009,N_19244);
nand U23178 (N_23178,N_19695,N_19956);
or U23179 (N_23179,N_17143,N_16184);
nor U23180 (N_23180,N_16460,N_15858);
nand U23181 (N_23181,N_15441,N_17979);
and U23182 (N_23182,N_19880,N_17765);
nand U23183 (N_23183,N_17445,N_18178);
or U23184 (N_23184,N_19647,N_15571);
and U23185 (N_23185,N_19045,N_19788);
xnor U23186 (N_23186,N_17297,N_15167);
nor U23187 (N_23187,N_19654,N_16343);
nand U23188 (N_23188,N_18173,N_19695);
xor U23189 (N_23189,N_18101,N_19344);
xor U23190 (N_23190,N_19386,N_17575);
xor U23191 (N_23191,N_17752,N_19667);
nor U23192 (N_23192,N_15156,N_18470);
or U23193 (N_23193,N_17111,N_19459);
nand U23194 (N_23194,N_16239,N_15117);
xnor U23195 (N_23195,N_18405,N_17811);
nand U23196 (N_23196,N_17264,N_17457);
nor U23197 (N_23197,N_15058,N_16676);
and U23198 (N_23198,N_19481,N_16776);
or U23199 (N_23199,N_18850,N_17813);
and U23200 (N_23200,N_17060,N_16967);
and U23201 (N_23201,N_15829,N_19856);
and U23202 (N_23202,N_16700,N_19989);
nand U23203 (N_23203,N_18070,N_16449);
or U23204 (N_23204,N_15851,N_15473);
nor U23205 (N_23205,N_18352,N_19312);
nor U23206 (N_23206,N_15456,N_16901);
nand U23207 (N_23207,N_15761,N_16983);
nor U23208 (N_23208,N_18776,N_18336);
nor U23209 (N_23209,N_15982,N_16606);
or U23210 (N_23210,N_16624,N_16426);
or U23211 (N_23211,N_15508,N_19456);
and U23212 (N_23212,N_18289,N_18770);
nand U23213 (N_23213,N_17539,N_16415);
and U23214 (N_23214,N_15149,N_17448);
or U23215 (N_23215,N_17668,N_17152);
or U23216 (N_23216,N_15295,N_16794);
or U23217 (N_23217,N_18057,N_17569);
nand U23218 (N_23218,N_18644,N_19286);
and U23219 (N_23219,N_17343,N_17751);
nand U23220 (N_23220,N_15869,N_16401);
xor U23221 (N_23221,N_19406,N_19001);
nand U23222 (N_23222,N_19665,N_18895);
or U23223 (N_23223,N_16663,N_16328);
or U23224 (N_23224,N_17156,N_16934);
nand U23225 (N_23225,N_16864,N_18230);
nand U23226 (N_23226,N_16934,N_16926);
nand U23227 (N_23227,N_19895,N_15368);
nand U23228 (N_23228,N_19455,N_17587);
and U23229 (N_23229,N_19846,N_17499);
nor U23230 (N_23230,N_16830,N_17989);
nand U23231 (N_23231,N_15382,N_17520);
nor U23232 (N_23232,N_19157,N_18328);
and U23233 (N_23233,N_19130,N_19404);
nand U23234 (N_23234,N_16354,N_18987);
and U23235 (N_23235,N_19371,N_17203);
xor U23236 (N_23236,N_18256,N_19704);
and U23237 (N_23237,N_17578,N_18471);
nor U23238 (N_23238,N_19884,N_18013);
nand U23239 (N_23239,N_19220,N_17553);
or U23240 (N_23240,N_19114,N_18696);
and U23241 (N_23241,N_17456,N_17606);
and U23242 (N_23242,N_17471,N_18979);
nor U23243 (N_23243,N_16424,N_19290);
and U23244 (N_23244,N_17252,N_19015);
nand U23245 (N_23245,N_16163,N_16956);
nor U23246 (N_23246,N_16263,N_18779);
or U23247 (N_23247,N_15661,N_19501);
or U23248 (N_23248,N_16169,N_18360);
and U23249 (N_23249,N_17355,N_19869);
nor U23250 (N_23250,N_18160,N_19979);
or U23251 (N_23251,N_15808,N_19044);
and U23252 (N_23252,N_15632,N_19420);
nor U23253 (N_23253,N_18947,N_18726);
nor U23254 (N_23254,N_17207,N_19989);
and U23255 (N_23255,N_15634,N_19902);
or U23256 (N_23256,N_15954,N_15895);
nand U23257 (N_23257,N_17554,N_17643);
or U23258 (N_23258,N_18604,N_19502);
and U23259 (N_23259,N_18979,N_16576);
nand U23260 (N_23260,N_16007,N_18396);
or U23261 (N_23261,N_15294,N_15431);
or U23262 (N_23262,N_17397,N_18742);
xor U23263 (N_23263,N_18738,N_17805);
xnor U23264 (N_23264,N_19906,N_15569);
and U23265 (N_23265,N_17489,N_16624);
xor U23266 (N_23266,N_19654,N_17541);
or U23267 (N_23267,N_18524,N_19035);
or U23268 (N_23268,N_16370,N_16120);
xor U23269 (N_23269,N_16000,N_18614);
nor U23270 (N_23270,N_19943,N_18497);
and U23271 (N_23271,N_18146,N_16035);
nor U23272 (N_23272,N_17749,N_17910);
nand U23273 (N_23273,N_16987,N_17415);
xnor U23274 (N_23274,N_17453,N_19031);
nor U23275 (N_23275,N_16880,N_19463);
nand U23276 (N_23276,N_15146,N_19126);
or U23277 (N_23277,N_19382,N_19654);
nand U23278 (N_23278,N_16870,N_16624);
and U23279 (N_23279,N_16426,N_16661);
and U23280 (N_23280,N_16308,N_18961);
xnor U23281 (N_23281,N_15997,N_19563);
or U23282 (N_23282,N_15583,N_16590);
and U23283 (N_23283,N_16874,N_16439);
xor U23284 (N_23284,N_15312,N_19891);
nand U23285 (N_23285,N_16570,N_19222);
xnor U23286 (N_23286,N_15689,N_15639);
or U23287 (N_23287,N_17723,N_18574);
and U23288 (N_23288,N_18030,N_16483);
and U23289 (N_23289,N_17318,N_19160);
nor U23290 (N_23290,N_15523,N_15977);
or U23291 (N_23291,N_15436,N_17814);
and U23292 (N_23292,N_17047,N_19013);
xnor U23293 (N_23293,N_16971,N_16921);
or U23294 (N_23294,N_16354,N_15392);
nor U23295 (N_23295,N_17649,N_18021);
or U23296 (N_23296,N_16186,N_16767);
or U23297 (N_23297,N_15492,N_19474);
nand U23298 (N_23298,N_18689,N_17120);
nor U23299 (N_23299,N_15195,N_17260);
or U23300 (N_23300,N_16458,N_19120);
and U23301 (N_23301,N_19390,N_19619);
or U23302 (N_23302,N_18280,N_15543);
nor U23303 (N_23303,N_16263,N_17798);
nand U23304 (N_23304,N_19507,N_17834);
nor U23305 (N_23305,N_18531,N_15655);
nand U23306 (N_23306,N_18885,N_15342);
or U23307 (N_23307,N_19613,N_18603);
nand U23308 (N_23308,N_18343,N_16648);
and U23309 (N_23309,N_15322,N_15111);
nand U23310 (N_23310,N_16126,N_18473);
nor U23311 (N_23311,N_19976,N_18859);
xnor U23312 (N_23312,N_18220,N_19872);
nand U23313 (N_23313,N_16261,N_15984);
nor U23314 (N_23314,N_18524,N_17526);
nand U23315 (N_23315,N_15338,N_17540);
or U23316 (N_23316,N_15939,N_16958);
nand U23317 (N_23317,N_19651,N_19539);
nor U23318 (N_23318,N_19748,N_15536);
and U23319 (N_23319,N_18750,N_16933);
nand U23320 (N_23320,N_17220,N_16779);
nand U23321 (N_23321,N_19275,N_15799);
nor U23322 (N_23322,N_15814,N_18204);
or U23323 (N_23323,N_15567,N_18218);
and U23324 (N_23324,N_18826,N_17500);
xnor U23325 (N_23325,N_18358,N_18074);
nand U23326 (N_23326,N_18739,N_18534);
nor U23327 (N_23327,N_18284,N_17754);
nand U23328 (N_23328,N_18807,N_18491);
nor U23329 (N_23329,N_15560,N_16733);
nor U23330 (N_23330,N_15993,N_19468);
nand U23331 (N_23331,N_19423,N_15300);
or U23332 (N_23332,N_19102,N_19836);
and U23333 (N_23333,N_15004,N_15096);
or U23334 (N_23334,N_15651,N_18781);
nand U23335 (N_23335,N_17724,N_19667);
or U23336 (N_23336,N_18229,N_15891);
xnor U23337 (N_23337,N_19681,N_17858);
nor U23338 (N_23338,N_16439,N_19852);
nor U23339 (N_23339,N_15258,N_16713);
or U23340 (N_23340,N_16207,N_18001);
or U23341 (N_23341,N_15052,N_18834);
xnor U23342 (N_23342,N_18436,N_15084);
nor U23343 (N_23343,N_18172,N_17026);
and U23344 (N_23344,N_16377,N_15243);
nor U23345 (N_23345,N_17051,N_17531);
and U23346 (N_23346,N_16848,N_19455);
or U23347 (N_23347,N_16053,N_19156);
nor U23348 (N_23348,N_15673,N_15785);
xor U23349 (N_23349,N_15723,N_19816);
nand U23350 (N_23350,N_15465,N_16325);
or U23351 (N_23351,N_17772,N_18250);
nand U23352 (N_23352,N_19763,N_15370);
nor U23353 (N_23353,N_18635,N_18789);
and U23354 (N_23354,N_17116,N_16343);
and U23355 (N_23355,N_15760,N_19866);
nand U23356 (N_23356,N_16413,N_17629);
xnor U23357 (N_23357,N_19113,N_19981);
nand U23358 (N_23358,N_19515,N_17916);
nand U23359 (N_23359,N_16812,N_15650);
nand U23360 (N_23360,N_16123,N_17721);
xor U23361 (N_23361,N_16946,N_15418);
xnor U23362 (N_23362,N_19986,N_16503);
nor U23363 (N_23363,N_18960,N_17114);
xor U23364 (N_23364,N_15856,N_16609);
xor U23365 (N_23365,N_16224,N_16738);
nand U23366 (N_23366,N_15619,N_15102);
or U23367 (N_23367,N_17157,N_15823);
and U23368 (N_23368,N_18614,N_15942);
or U23369 (N_23369,N_16328,N_16066);
or U23370 (N_23370,N_18334,N_15424);
and U23371 (N_23371,N_19814,N_17221);
nand U23372 (N_23372,N_16254,N_15453);
nor U23373 (N_23373,N_16707,N_16791);
nand U23374 (N_23374,N_19631,N_17944);
and U23375 (N_23375,N_17282,N_16381);
and U23376 (N_23376,N_18223,N_19620);
nor U23377 (N_23377,N_18540,N_17965);
xor U23378 (N_23378,N_17634,N_16771);
xor U23379 (N_23379,N_16882,N_18239);
or U23380 (N_23380,N_19755,N_18341);
or U23381 (N_23381,N_16803,N_17923);
or U23382 (N_23382,N_15949,N_16390);
nand U23383 (N_23383,N_18983,N_19086);
nor U23384 (N_23384,N_16089,N_17953);
xnor U23385 (N_23385,N_16220,N_15673);
nand U23386 (N_23386,N_19860,N_18081);
or U23387 (N_23387,N_16840,N_18672);
xnor U23388 (N_23388,N_19370,N_17382);
and U23389 (N_23389,N_15779,N_19571);
and U23390 (N_23390,N_18251,N_17342);
and U23391 (N_23391,N_19463,N_15599);
nor U23392 (N_23392,N_16101,N_17666);
or U23393 (N_23393,N_17244,N_19542);
nand U23394 (N_23394,N_15441,N_18653);
xnor U23395 (N_23395,N_16265,N_15837);
or U23396 (N_23396,N_16540,N_18204);
nor U23397 (N_23397,N_18536,N_18189);
xor U23398 (N_23398,N_17565,N_19253);
and U23399 (N_23399,N_18433,N_16379);
nor U23400 (N_23400,N_16759,N_16306);
xor U23401 (N_23401,N_17002,N_16688);
or U23402 (N_23402,N_16449,N_15934);
nor U23403 (N_23403,N_19630,N_15363);
and U23404 (N_23404,N_19173,N_17895);
or U23405 (N_23405,N_17745,N_19318);
or U23406 (N_23406,N_16929,N_19621);
nor U23407 (N_23407,N_18678,N_16230);
or U23408 (N_23408,N_16412,N_18240);
or U23409 (N_23409,N_19280,N_15437);
nand U23410 (N_23410,N_18417,N_19651);
and U23411 (N_23411,N_19240,N_18448);
nand U23412 (N_23412,N_16236,N_19061);
nand U23413 (N_23413,N_15211,N_19461);
and U23414 (N_23414,N_15566,N_17576);
nand U23415 (N_23415,N_19091,N_19894);
nand U23416 (N_23416,N_15149,N_17462);
and U23417 (N_23417,N_18505,N_19008);
or U23418 (N_23418,N_15985,N_16364);
xnor U23419 (N_23419,N_16090,N_19341);
and U23420 (N_23420,N_19448,N_15958);
nor U23421 (N_23421,N_15464,N_15630);
xor U23422 (N_23422,N_15881,N_15672);
and U23423 (N_23423,N_16505,N_16345);
xor U23424 (N_23424,N_17724,N_17011);
xnor U23425 (N_23425,N_16411,N_16409);
xor U23426 (N_23426,N_15143,N_16713);
or U23427 (N_23427,N_15964,N_19655);
nand U23428 (N_23428,N_18615,N_17907);
xnor U23429 (N_23429,N_18954,N_16221);
nand U23430 (N_23430,N_17764,N_18306);
or U23431 (N_23431,N_16235,N_16408);
or U23432 (N_23432,N_18653,N_19651);
nand U23433 (N_23433,N_17026,N_16751);
and U23434 (N_23434,N_18595,N_15340);
and U23435 (N_23435,N_18352,N_18765);
xnor U23436 (N_23436,N_17286,N_19917);
xor U23437 (N_23437,N_16745,N_15770);
nor U23438 (N_23438,N_18003,N_15107);
nand U23439 (N_23439,N_17896,N_18965);
nor U23440 (N_23440,N_16459,N_16800);
or U23441 (N_23441,N_16494,N_15737);
and U23442 (N_23442,N_17988,N_18451);
and U23443 (N_23443,N_18719,N_17250);
nor U23444 (N_23444,N_19348,N_17892);
or U23445 (N_23445,N_17268,N_18704);
and U23446 (N_23446,N_16617,N_17769);
nand U23447 (N_23447,N_15211,N_16067);
nor U23448 (N_23448,N_17206,N_15285);
and U23449 (N_23449,N_18973,N_15494);
and U23450 (N_23450,N_17228,N_17944);
nand U23451 (N_23451,N_19438,N_16398);
nand U23452 (N_23452,N_15109,N_18882);
nor U23453 (N_23453,N_17027,N_17454);
xnor U23454 (N_23454,N_16475,N_16782);
or U23455 (N_23455,N_17732,N_17297);
xnor U23456 (N_23456,N_15528,N_19244);
and U23457 (N_23457,N_15574,N_17555);
or U23458 (N_23458,N_19269,N_19948);
nand U23459 (N_23459,N_16454,N_16272);
or U23460 (N_23460,N_16783,N_18693);
xor U23461 (N_23461,N_16348,N_15745);
nand U23462 (N_23462,N_16099,N_16261);
nand U23463 (N_23463,N_19373,N_18033);
and U23464 (N_23464,N_19621,N_15670);
xor U23465 (N_23465,N_17784,N_18473);
nor U23466 (N_23466,N_19445,N_19366);
or U23467 (N_23467,N_18003,N_18629);
nand U23468 (N_23468,N_15294,N_18354);
or U23469 (N_23469,N_16856,N_18289);
xor U23470 (N_23470,N_17843,N_16397);
and U23471 (N_23471,N_18173,N_18399);
nor U23472 (N_23472,N_17267,N_15727);
nor U23473 (N_23473,N_18511,N_16853);
nor U23474 (N_23474,N_15199,N_16637);
nand U23475 (N_23475,N_19004,N_15880);
and U23476 (N_23476,N_18707,N_16065);
and U23477 (N_23477,N_17586,N_16981);
and U23478 (N_23478,N_15426,N_16870);
nand U23479 (N_23479,N_18594,N_16304);
xnor U23480 (N_23480,N_19953,N_17488);
nand U23481 (N_23481,N_16711,N_17158);
nand U23482 (N_23482,N_19716,N_18350);
nand U23483 (N_23483,N_18084,N_16546);
xor U23484 (N_23484,N_19313,N_18955);
nand U23485 (N_23485,N_16641,N_16769);
and U23486 (N_23486,N_19039,N_16877);
or U23487 (N_23487,N_16418,N_15170);
nor U23488 (N_23488,N_16662,N_17678);
nor U23489 (N_23489,N_15605,N_15830);
and U23490 (N_23490,N_18228,N_16228);
nor U23491 (N_23491,N_19795,N_18484);
and U23492 (N_23492,N_18886,N_16614);
or U23493 (N_23493,N_18287,N_19633);
and U23494 (N_23494,N_16234,N_18005);
and U23495 (N_23495,N_19201,N_19302);
nand U23496 (N_23496,N_16777,N_18735);
and U23497 (N_23497,N_19409,N_18284);
nand U23498 (N_23498,N_18642,N_15927);
xnor U23499 (N_23499,N_15909,N_19174);
and U23500 (N_23500,N_17588,N_16953);
or U23501 (N_23501,N_16688,N_17167);
or U23502 (N_23502,N_18899,N_19645);
nor U23503 (N_23503,N_15063,N_17756);
or U23504 (N_23504,N_19801,N_16640);
and U23505 (N_23505,N_15043,N_16449);
nand U23506 (N_23506,N_17015,N_19304);
nor U23507 (N_23507,N_17536,N_19613);
and U23508 (N_23508,N_17977,N_16086);
nor U23509 (N_23509,N_19891,N_16007);
nor U23510 (N_23510,N_17055,N_19629);
and U23511 (N_23511,N_15761,N_16774);
and U23512 (N_23512,N_15442,N_19121);
xor U23513 (N_23513,N_17189,N_16619);
and U23514 (N_23514,N_17073,N_19301);
xnor U23515 (N_23515,N_15835,N_18827);
nand U23516 (N_23516,N_19669,N_19917);
nand U23517 (N_23517,N_18539,N_19136);
or U23518 (N_23518,N_18251,N_19765);
and U23519 (N_23519,N_15878,N_16466);
nor U23520 (N_23520,N_16346,N_17718);
and U23521 (N_23521,N_16938,N_18329);
or U23522 (N_23522,N_15475,N_16826);
nand U23523 (N_23523,N_18601,N_17767);
and U23524 (N_23524,N_19838,N_19191);
and U23525 (N_23525,N_16184,N_19702);
xnor U23526 (N_23526,N_16078,N_15904);
xnor U23527 (N_23527,N_19081,N_19817);
and U23528 (N_23528,N_17963,N_15719);
nand U23529 (N_23529,N_17921,N_17161);
nor U23530 (N_23530,N_18093,N_17277);
nor U23531 (N_23531,N_19311,N_15744);
or U23532 (N_23532,N_18728,N_17802);
nor U23533 (N_23533,N_18052,N_18618);
nand U23534 (N_23534,N_17008,N_18991);
nand U23535 (N_23535,N_17527,N_16717);
nand U23536 (N_23536,N_18016,N_19586);
nor U23537 (N_23537,N_19673,N_15336);
nor U23538 (N_23538,N_15495,N_18522);
or U23539 (N_23539,N_17456,N_15762);
nor U23540 (N_23540,N_15239,N_16286);
xor U23541 (N_23541,N_16958,N_16457);
nor U23542 (N_23542,N_19089,N_19013);
nand U23543 (N_23543,N_16761,N_15397);
nand U23544 (N_23544,N_19832,N_18368);
nor U23545 (N_23545,N_16701,N_19393);
or U23546 (N_23546,N_17791,N_18649);
xor U23547 (N_23547,N_17217,N_17976);
xor U23548 (N_23548,N_17748,N_19395);
and U23549 (N_23549,N_18110,N_19114);
nand U23550 (N_23550,N_18914,N_17016);
xnor U23551 (N_23551,N_16802,N_19406);
and U23552 (N_23552,N_15211,N_19487);
and U23553 (N_23553,N_16790,N_18593);
and U23554 (N_23554,N_15707,N_16379);
and U23555 (N_23555,N_17532,N_16330);
and U23556 (N_23556,N_15421,N_17310);
xnor U23557 (N_23557,N_18395,N_18679);
nand U23558 (N_23558,N_19838,N_15457);
nand U23559 (N_23559,N_17961,N_16575);
xor U23560 (N_23560,N_15231,N_15009);
or U23561 (N_23561,N_15353,N_19817);
nor U23562 (N_23562,N_19411,N_17038);
or U23563 (N_23563,N_16291,N_17266);
or U23564 (N_23564,N_15144,N_19036);
nand U23565 (N_23565,N_18119,N_19776);
nand U23566 (N_23566,N_15778,N_18378);
and U23567 (N_23567,N_19947,N_18772);
or U23568 (N_23568,N_17423,N_16664);
and U23569 (N_23569,N_19554,N_17858);
nand U23570 (N_23570,N_16984,N_15557);
xnor U23571 (N_23571,N_16877,N_15185);
xor U23572 (N_23572,N_15174,N_15165);
and U23573 (N_23573,N_18445,N_18640);
nor U23574 (N_23574,N_15655,N_18977);
xnor U23575 (N_23575,N_19773,N_19349);
nor U23576 (N_23576,N_18495,N_18727);
or U23577 (N_23577,N_15073,N_15295);
xor U23578 (N_23578,N_19456,N_15065);
or U23579 (N_23579,N_17366,N_18306);
nand U23580 (N_23580,N_17296,N_16016);
or U23581 (N_23581,N_16125,N_19018);
and U23582 (N_23582,N_17088,N_17332);
or U23583 (N_23583,N_19518,N_18588);
nor U23584 (N_23584,N_19333,N_19562);
xnor U23585 (N_23585,N_15623,N_15309);
and U23586 (N_23586,N_16013,N_17388);
or U23587 (N_23587,N_16454,N_16987);
xnor U23588 (N_23588,N_17390,N_15820);
nor U23589 (N_23589,N_17556,N_17980);
and U23590 (N_23590,N_16481,N_15781);
xnor U23591 (N_23591,N_16196,N_16474);
nand U23592 (N_23592,N_19123,N_15977);
nand U23593 (N_23593,N_18878,N_18785);
and U23594 (N_23594,N_17244,N_15792);
nor U23595 (N_23595,N_17872,N_17206);
nor U23596 (N_23596,N_19980,N_15713);
or U23597 (N_23597,N_15118,N_15601);
xor U23598 (N_23598,N_15086,N_18435);
or U23599 (N_23599,N_18122,N_15527);
xor U23600 (N_23600,N_16192,N_18651);
and U23601 (N_23601,N_18390,N_18487);
xnor U23602 (N_23602,N_18746,N_16111);
nand U23603 (N_23603,N_19033,N_18628);
nand U23604 (N_23604,N_19748,N_17003);
nor U23605 (N_23605,N_18347,N_17728);
or U23606 (N_23606,N_17210,N_18724);
and U23607 (N_23607,N_16185,N_18371);
and U23608 (N_23608,N_15888,N_19086);
or U23609 (N_23609,N_19667,N_18235);
nor U23610 (N_23610,N_19745,N_15568);
nand U23611 (N_23611,N_15149,N_15955);
xnor U23612 (N_23612,N_18462,N_15418);
or U23613 (N_23613,N_15982,N_15065);
nand U23614 (N_23614,N_15519,N_16891);
nand U23615 (N_23615,N_18666,N_16030);
and U23616 (N_23616,N_16286,N_19521);
nor U23617 (N_23617,N_16043,N_19251);
xor U23618 (N_23618,N_16497,N_18685);
and U23619 (N_23619,N_19617,N_19576);
nor U23620 (N_23620,N_17485,N_17056);
or U23621 (N_23621,N_18746,N_18432);
xor U23622 (N_23622,N_15235,N_15172);
xnor U23623 (N_23623,N_15070,N_19003);
nor U23624 (N_23624,N_18816,N_18578);
nor U23625 (N_23625,N_18226,N_18185);
nand U23626 (N_23626,N_18981,N_18102);
xnor U23627 (N_23627,N_15816,N_16449);
or U23628 (N_23628,N_15026,N_17972);
or U23629 (N_23629,N_18075,N_17676);
nor U23630 (N_23630,N_16024,N_17533);
nand U23631 (N_23631,N_16733,N_17889);
and U23632 (N_23632,N_19901,N_18925);
or U23633 (N_23633,N_17922,N_17367);
or U23634 (N_23634,N_17824,N_19543);
nand U23635 (N_23635,N_15821,N_17687);
or U23636 (N_23636,N_19379,N_16580);
nand U23637 (N_23637,N_15474,N_17420);
or U23638 (N_23638,N_18936,N_19967);
or U23639 (N_23639,N_17697,N_19666);
and U23640 (N_23640,N_19221,N_18608);
xnor U23641 (N_23641,N_15903,N_17409);
xor U23642 (N_23642,N_18010,N_17986);
and U23643 (N_23643,N_17555,N_19690);
and U23644 (N_23644,N_16225,N_15311);
or U23645 (N_23645,N_17022,N_19580);
nor U23646 (N_23646,N_18625,N_18952);
xnor U23647 (N_23647,N_17115,N_19972);
xnor U23648 (N_23648,N_18461,N_16440);
xor U23649 (N_23649,N_16537,N_19959);
or U23650 (N_23650,N_19238,N_19193);
and U23651 (N_23651,N_18306,N_18336);
nand U23652 (N_23652,N_15880,N_17290);
or U23653 (N_23653,N_19859,N_18899);
and U23654 (N_23654,N_15350,N_16133);
nand U23655 (N_23655,N_18754,N_17759);
and U23656 (N_23656,N_18763,N_18865);
nor U23657 (N_23657,N_19931,N_16653);
nor U23658 (N_23658,N_15316,N_15950);
nor U23659 (N_23659,N_19544,N_17081);
and U23660 (N_23660,N_17092,N_15433);
xor U23661 (N_23661,N_16306,N_16958);
and U23662 (N_23662,N_16479,N_15295);
nor U23663 (N_23663,N_16221,N_17957);
nand U23664 (N_23664,N_19274,N_18545);
nor U23665 (N_23665,N_15196,N_15672);
nor U23666 (N_23666,N_18042,N_18298);
nand U23667 (N_23667,N_18902,N_18401);
and U23668 (N_23668,N_16795,N_19151);
or U23669 (N_23669,N_15245,N_16834);
and U23670 (N_23670,N_19805,N_19308);
nor U23671 (N_23671,N_17997,N_17505);
nor U23672 (N_23672,N_16521,N_16243);
or U23673 (N_23673,N_16156,N_19828);
nor U23674 (N_23674,N_18039,N_15756);
and U23675 (N_23675,N_15963,N_19547);
or U23676 (N_23676,N_15037,N_17808);
nand U23677 (N_23677,N_16960,N_17261);
xor U23678 (N_23678,N_16467,N_15481);
xnor U23679 (N_23679,N_19970,N_16045);
and U23680 (N_23680,N_15048,N_15645);
or U23681 (N_23681,N_15140,N_19185);
nor U23682 (N_23682,N_16804,N_16504);
nand U23683 (N_23683,N_16043,N_19789);
or U23684 (N_23684,N_18486,N_18303);
or U23685 (N_23685,N_18316,N_18331);
nor U23686 (N_23686,N_16060,N_17204);
and U23687 (N_23687,N_17348,N_16181);
nand U23688 (N_23688,N_16982,N_16891);
xnor U23689 (N_23689,N_17641,N_16868);
nor U23690 (N_23690,N_19674,N_17540);
nor U23691 (N_23691,N_16808,N_15582);
nand U23692 (N_23692,N_16667,N_15033);
nand U23693 (N_23693,N_18721,N_19721);
and U23694 (N_23694,N_16166,N_19386);
nor U23695 (N_23695,N_19324,N_18425);
xnor U23696 (N_23696,N_19455,N_19876);
nor U23697 (N_23697,N_18804,N_19169);
xor U23698 (N_23698,N_17155,N_18201);
and U23699 (N_23699,N_16896,N_18528);
nand U23700 (N_23700,N_19473,N_19814);
nand U23701 (N_23701,N_15485,N_16250);
nand U23702 (N_23702,N_18955,N_19355);
and U23703 (N_23703,N_15062,N_18291);
nand U23704 (N_23704,N_17885,N_16864);
and U23705 (N_23705,N_16180,N_17080);
or U23706 (N_23706,N_19849,N_17456);
nor U23707 (N_23707,N_17618,N_19573);
or U23708 (N_23708,N_17585,N_17857);
nor U23709 (N_23709,N_19107,N_19453);
nor U23710 (N_23710,N_18356,N_16808);
nor U23711 (N_23711,N_18839,N_19700);
nand U23712 (N_23712,N_19486,N_19121);
and U23713 (N_23713,N_17887,N_16800);
or U23714 (N_23714,N_19723,N_18825);
nand U23715 (N_23715,N_15558,N_19288);
and U23716 (N_23716,N_17025,N_19272);
and U23717 (N_23717,N_19844,N_19313);
nand U23718 (N_23718,N_15790,N_19422);
nor U23719 (N_23719,N_15842,N_15554);
nor U23720 (N_23720,N_15755,N_19558);
nor U23721 (N_23721,N_16859,N_16442);
and U23722 (N_23722,N_19705,N_19424);
and U23723 (N_23723,N_18779,N_18630);
nand U23724 (N_23724,N_18747,N_18058);
or U23725 (N_23725,N_19417,N_18654);
xnor U23726 (N_23726,N_16745,N_19628);
nor U23727 (N_23727,N_18790,N_15194);
or U23728 (N_23728,N_15754,N_19016);
or U23729 (N_23729,N_17559,N_17110);
and U23730 (N_23730,N_18856,N_15389);
nor U23731 (N_23731,N_18270,N_18824);
xor U23732 (N_23732,N_17666,N_16177);
nand U23733 (N_23733,N_16908,N_18789);
nand U23734 (N_23734,N_18277,N_19958);
or U23735 (N_23735,N_15760,N_19573);
and U23736 (N_23736,N_18104,N_16080);
nand U23737 (N_23737,N_18982,N_16734);
nand U23738 (N_23738,N_17916,N_19982);
xnor U23739 (N_23739,N_17334,N_16770);
and U23740 (N_23740,N_16314,N_15747);
xnor U23741 (N_23741,N_18539,N_17853);
or U23742 (N_23742,N_19713,N_17027);
nor U23743 (N_23743,N_16775,N_18287);
xor U23744 (N_23744,N_17241,N_17096);
and U23745 (N_23745,N_15267,N_19431);
and U23746 (N_23746,N_19642,N_16270);
xor U23747 (N_23747,N_16529,N_17158);
nor U23748 (N_23748,N_17029,N_15660);
and U23749 (N_23749,N_18577,N_16440);
nand U23750 (N_23750,N_15163,N_17800);
and U23751 (N_23751,N_17907,N_17686);
and U23752 (N_23752,N_15580,N_17467);
nand U23753 (N_23753,N_16444,N_17916);
or U23754 (N_23754,N_19078,N_16368);
xnor U23755 (N_23755,N_19123,N_16301);
or U23756 (N_23756,N_19002,N_18659);
nor U23757 (N_23757,N_17211,N_16877);
xor U23758 (N_23758,N_16764,N_16447);
or U23759 (N_23759,N_18037,N_15358);
nand U23760 (N_23760,N_16717,N_18082);
xnor U23761 (N_23761,N_17755,N_17133);
nor U23762 (N_23762,N_16553,N_17054);
xor U23763 (N_23763,N_18173,N_17917);
or U23764 (N_23764,N_15958,N_18342);
and U23765 (N_23765,N_16862,N_17155);
and U23766 (N_23766,N_18335,N_16183);
nand U23767 (N_23767,N_15621,N_19970);
nand U23768 (N_23768,N_18847,N_19318);
nand U23769 (N_23769,N_16679,N_17276);
nor U23770 (N_23770,N_15835,N_17975);
nor U23771 (N_23771,N_15470,N_18123);
nor U23772 (N_23772,N_19223,N_17168);
xor U23773 (N_23773,N_18238,N_17854);
xor U23774 (N_23774,N_19043,N_18559);
xor U23775 (N_23775,N_17806,N_18734);
nand U23776 (N_23776,N_18538,N_16332);
and U23777 (N_23777,N_18088,N_17178);
nand U23778 (N_23778,N_18522,N_19488);
nor U23779 (N_23779,N_18109,N_17061);
nand U23780 (N_23780,N_16266,N_19082);
nor U23781 (N_23781,N_16294,N_19932);
xor U23782 (N_23782,N_15074,N_18618);
xor U23783 (N_23783,N_15229,N_15854);
nand U23784 (N_23784,N_16538,N_19226);
xnor U23785 (N_23785,N_15714,N_18876);
nor U23786 (N_23786,N_16359,N_16916);
and U23787 (N_23787,N_15809,N_16720);
xnor U23788 (N_23788,N_15838,N_15232);
or U23789 (N_23789,N_16794,N_17583);
or U23790 (N_23790,N_18212,N_18682);
nor U23791 (N_23791,N_16495,N_18744);
or U23792 (N_23792,N_16904,N_17167);
or U23793 (N_23793,N_17763,N_18639);
or U23794 (N_23794,N_15968,N_15911);
and U23795 (N_23795,N_19464,N_18743);
xnor U23796 (N_23796,N_15057,N_17038);
xnor U23797 (N_23797,N_15249,N_18643);
nor U23798 (N_23798,N_19175,N_15494);
nor U23799 (N_23799,N_19174,N_15379);
and U23800 (N_23800,N_16698,N_16153);
nand U23801 (N_23801,N_17397,N_18435);
nand U23802 (N_23802,N_18038,N_17868);
nor U23803 (N_23803,N_16623,N_15737);
nor U23804 (N_23804,N_18347,N_18280);
nand U23805 (N_23805,N_15530,N_15458);
xor U23806 (N_23806,N_19103,N_15394);
xor U23807 (N_23807,N_19364,N_16213);
xor U23808 (N_23808,N_15590,N_15955);
or U23809 (N_23809,N_19388,N_18131);
nand U23810 (N_23810,N_18873,N_18357);
xnor U23811 (N_23811,N_15339,N_17537);
or U23812 (N_23812,N_16031,N_19431);
and U23813 (N_23813,N_15145,N_16218);
or U23814 (N_23814,N_17819,N_18318);
xor U23815 (N_23815,N_18559,N_17767);
xor U23816 (N_23816,N_17407,N_19909);
nor U23817 (N_23817,N_17214,N_19717);
or U23818 (N_23818,N_17175,N_16796);
and U23819 (N_23819,N_19579,N_19391);
nand U23820 (N_23820,N_16518,N_15231);
xnor U23821 (N_23821,N_16419,N_16415);
nand U23822 (N_23822,N_18699,N_18635);
nor U23823 (N_23823,N_18668,N_15039);
or U23824 (N_23824,N_19950,N_15988);
nand U23825 (N_23825,N_18486,N_18267);
nor U23826 (N_23826,N_19528,N_16144);
xnor U23827 (N_23827,N_17470,N_18714);
and U23828 (N_23828,N_15804,N_17823);
xor U23829 (N_23829,N_16279,N_16781);
or U23830 (N_23830,N_15044,N_18620);
nor U23831 (N_23831,N_18867,N_15029);
nor U23832 (N_23832,N_19938,N_16816);
and U23833 (N_23833,N_19110,N_17244);
or U23834 (N_23834,N_15277,N_18299);
and U23835 (N_23835,N_19533,N_19111);
and U23836 (N_23836,N_19970,N_16636);
nand U23837 (N_23837,N_19307,N_16002);
nand U23838 (N_23838,N_19312,N_17097);
and U23839 (N_23839,N_15683,N_16767);
or U23840 (N_23840,N_19378,N_17540);
nand U23841 (N_23841,N_15990,N_19112);
xnor U23842 (N_23842,N_15470,N_17875);
nand U23843 (N_23843,N_18688,N_19677);
xnor U23844 (N_23844,N_18006,N_18827);
nand U23845 (N_23845,N_15810,N_16756);
or U23846 (N_23846,N_15156,N_16475);
and U23847 (N_23847,N_17381,N_17128);
nand U23848 (N_23848,N_15355,N_15741);
or U23849 (N_23849,N_17434,N_17239);
or U23850 (N_23850,N_17285,N_15622);
nand U23851 (N_23851,N_18304,N_17681);
or U23852 (N_23852,N_19230,N_16347);
or U23853 (N_23853,N_18645,N_17595);
xnor U23854 (N_23854,N_16500,N_15283);
nor U23855 (N_23855,N_17076,N_16115);
xnor U23856 (N_23856,N_17020,N_16027);
nand U23857 (N_23857,N_18253,N_17193);
nand U23858 (N_23858,N_18483,N_16496);
nand U23859 (N_23859,N_15073,N_19667);
xor U23860 (N_23860,N_18716,N_16397);
nand U23861 (N_23861,N_15658,N_16874);
and U23862 (N_23862,N_15604,N_15249);
xnor U23863 (N_23863,N_17138,N_18221);
nor U23864 (N_23864,N_16092,N_15410);
nand U23865 (N_23865,N_16035,N_16942);
or U23866 (N_23866,N_16503,N_18257);
and U23867 (N_23867,N_19132,N_16551);
and U23868 (N_23868,N_16677,N_15676);
or U23869 (N_23869,N_15143,N_17520);
nand U23870 (N_23870,N_15676,N_15528);
nand U23871 (N_23871,N_18420,N_17987);
or U23872 (N_23872,N_15750,N_15174);
or U23873 (N_23873,N_19395,N_16944);
and U23874 (N_23874,N_18301,N_15056);
and U23875 (N_23875,N_17697,N_16416);
and U23876 (N_23876,N_19996,N_15918);
nor U23877 (N_23877,N_19372,N_18772);
nor U23878 (N_23878,N_18173,N_16320);
xnor U23879 (N_23879,N_16866,N_16205);
nor U23880 (N_23880,N_18100,N_17964);
nor U23881 (N_23881,N_15462,N_16151);
xor U23882 (N_23882,N_19969,N_16074);
or U23883 (N_23883,N_19761,N_18576);
and U23884 (N_23884,N_17281,N_17924);
and U23885 (N_23885,N_15827,N_16461);
nand U23886 (N_23886,N_16809,N_18366);
and U23887 (N_23887,N_18092,N_16089);
xor U23888 (N_23888,N_15741,N_18351);
and U23889 (N_23889,N_16394,N_15747);
xor U23890 (N_23890,N_19298,N_15245);
xnor U23891 (N_23891,N_15238,N_18591);
xnor U23892 (N_23892,N_16818,N_15477);
nand U23893 (N_23893,N_16807,N_15609);
nor U23894 (N_23894,N_17916,N_18468);
nand U23895 (N_23895,N_18853,N_19748);
or U23896 (N_23896,N_17372,N_18565);
nand U23897 (N_23897,N_16472,N_15452);
nand U23898 (N_23898,N_19815,N_16272);
nor U23899 (N_23899,N_17712,N_15132);
or U23900 (N_23900,N_17402,N_19000);
xnor U23901 (N_23901,N_18949,N_15471);
and U23902 (N_23902,N_17244,N_19109);
nand U23903 (N_23903,N_17042,N_18905);
nor U23904 (N_23904,N_16789,N_17512);
or U23905 (N_23905,N_18792,N_19748);
and U23906 (N_23906,N_16633,N_19071);
nor U23907 (N_23907,N_19018,N_17227);
or U23908 (N_23908,N_15785,N_15058);
or U23909 (N_23909,N_16726,N_17646);
nand U23910 (N_23910,N_19253,N_17710);
or U23911 (N_23911,N_17885,N_19071);
or U23912 (N_23912,N_16241,N_15908);
nand U23913 (N_23913,N_15965,N_15216);
nor U23914 (N_23914,N_17575,N_15442);
or U23915 (N_23915,N_19997,N_19898);
and U23916 (N_23916,N_15192,N_18463);
or U23917 (N_23917,N_17062,N_15718);
or U23918 (N_23918,N_16876,N_16575);
or U23919 (N_23919,N_19586,N_16091);
xnor U23920 (N_23920,N_15811,N_16140);
xor U23921 (N_23921,N_15947,N_15139);
nand U23922 (N_23922,N_15034,N_17614);
and U23923 (N_23923,N_18664,N_16175);
nand U23924 (N_23924,N_16746,N_17258);
or U23925 (N_23925,N_18877,N_15691);
and U23926 (N_23926,N_18998,N_18833);
xnor U23927 (N_23927,N_16226,N_19039);
xor U23928 (N_23928,N_17136,N_19512);
nor U23929 (N_23929,N_16700,N_16695);
nor U23930 (N_23930,N_19262,N_17677);
and U23931 (N_23931,N_16401,N_16019);
xnor U23932 (N_23932,N_17562,N_19740);
nand U23933 (N_23933,N_15425,N_19785);
xnor U23934 (N_23934,N_17184,N_19891);
or U23935 (N_23935,N_15541,N_16666);
and U23936 (N_23936,N_16963,N_18035);
nor U23937 (N_23937,N_17659,N_18164);
or U23938 (N_23938,N_15931,N_18852);
and U23939 (N_23939,N_15117,N_17455);
nand U23940 (N_23940,N_16471,N_15185);
or U23941 (N_23941,N_18619,N_18248);
and U23942 (N_23942,N_15517,N_17765);
nand U23943 (N_23943,N_19959,N_18738);
and U23944 (N_23944,N_15536,N_15703);
xnor U23945 (N_23945,N_16698,N_16898);
nor U23946 (N_23946,N_19862,N_19912);
xor U23947 (N_23947,N_18739,N_17739);
nand U23948 (N_23948,N_17628,N_15962);
and U23949 (N_23949,N_16562,N_15009);
or U23950 (N_23950,N_18581,N_19324);
nand U23951 (N_23951,N_15696,N_18699);
and U23952 (N_23952,N_18743,N_19744);
nand U23953 (N_23953,N_19975,N_19432);
nor U23954 (N_23954,N_19227,N_15862);
nand U23955 (N_23955,N_17998,N_17441);
and U23956 (N_23956,N_19998,N_15306);
nand U23957 (N_23957,N_15997,N_18759);
xnor U23958 (N_23958,N_15089,N_18474);
nand U23959 (N_23959,N_19088,N_18041);
xnor U23960 (N_23960,N_19110,N_18315);
or U23961 (N_23961,N_19302,N_17885);
or U23962 (N_23962,N_18660,N_18865);
xor U23963 (N_23963,N_15338,N_16681);
or U23964 (N_23964,N_18458,N_18454);
and U23965 (N_23965,N_18323,N_15115);
and U23966 (N_23966,N_18533,N_18577);
xnor U23967 (N_23967,N_16348,N_18951);
nand U23968 (N_23968,N_19483,N_16237);
nand U23969 (N_23969,N_19306,N_15718);
and U23970 (N_23970,N_19476,N_16985);
or U23971 (N_23971,N_19028,N_19126);
or U23972 (N_23972,N_16728,N_15018);
or U23973 (N_23973,N_17146,N_19373);
and U23974 (N_23974,N_16095,N_19249);
nand U23975 (N_23975,N_15609,N_15235);
xor U23976 (N_23976,N_16399,N_18138);
xor U23977 (N_23977,N_19093,N_16835);
and U23978 (N_23978,N_18313,N_19542);
and U23979 (N_23979,N_15407,N_15609);
and U23980 (N_23980,N_19969,N_18596);
nand U23981 (N_23981,N_17985,N_19904);
nor U23982 (N_23982,N_15312,N_15736);
xnor U23983 (N_23983,N_18724,N_18099);
nor U23984 (N_23984,N_18257,N_19532);
and U23985 (N_23985,N_17996,N_19867);
nor U23986 (N_23986,N_19158,N_19986);
xnor U23987 (N_23987,N_18227,N_18706);
xnor U23988 (N_23988,N_17670,N_15965);
and U23989 (N_23989,N_18977,N_18488);
nand U23990 (N_23990,N_17531,N_18753);
and U23991 (N_23991,N_18111,N_16788);
nand U23992 (N_23992,N_17878,N_16532);
nand U23993 (N_23993,N_19229,N_18358);
nand U23994 (N_23994,N_15934,N_15197);
and U23995 (N_23995,N_15503,N_18833);
and U23996 (N_23996,N_18590,N_18490);
and U23997 (N_23997,N_19840,N_16942);
xor U23998 (N_23998,N_19832,N_15998);
nor U23999 (N_23999,N_19740,N_15400);
xor U24000 (N_24000,N_18280,N_15929);
nor U24001 (N_24001,N_16520,N_18368);
xor U24002 (N_24002,N_18652,N_15519);
or U24003 (N_24003,N_19093,N_18226);
xor U24004 (N_24004,N_18109,N_19071);
and U24005 (N_24005,N_15312,N_15695);
or U24006 (N_24006,N_16666,N_16879);
or U24007 (N_24007,N_17356,N_16544);
nor U24008 (N_24008,N_18634,N_15189);
xnor U24009 (N_24009,N_19618,N_15113);
or U24010 (N_24010,N_18708,N_16064);
nand U24011 (N_24011,N_19165,N_17934);
nand U24012 (N_24012,N_19629,N_16330);
xor U24013 (N_24013,N_16076,N_15898);
xnor U24014 (N_24014,N_17322,N_18392);
or U24015 (N_24015,N_18229,N_16523);
nor U24016 (N_24016,N_15950,N_15727);
nor U24017 (N_24017,N_19872,N_18311);
or U24018 (N_24018,N_18846,N_16990);
nor U24019 (N_24019,N_16153,N_15100);
nand U24020 (N_24020,N_18690,N_18018);
nor U24021 (N_24021,N_19033,N_16733);
xnor U24022 (N_24022,N_16123,N_16928);
and U24023 (N_24023,N_19906,N_16302);
nand U24024 (N_24024,N_16569,N_18650);
nand U24025 (N_24025,N_15761,N_17506);
nor U24026 (N_24026,N_17754,N_19358);
xor U24027 (N_24027,N_18959,N_19076);
nand U24028 (N_24028,N_19899,N_18733);
or U24029 (N_24029,N_18984,N_17323);
nand U24030 (N_24030,N_18729,N_19217);
and U24031 (N_24031,N_17226,N_19697);
nand U24032 (N_24032,N_17645,N_18227);
xor U24033 (N_24033,N_17442,N_17049);
and U24034 (N_24034,N_19569,N_18131);
and U24035 (N_24035,N_18821,N_15615);
and U24036 (N_24036,N_17979,N_16688);
xor U24037 (N_24037,N_15433,N_17728);
and U24038 (N_24038,N_16373,N_16164);
nand U24039 (N_24039,N_17212,N_16879);
xnor U24040 (N_24040,N_16224,N_15037);
nor U24041 (N_24041,N_16138,N_17077);
nand U24042 (N_24042,N_17733,N_16981);
nand U24043 (N_24043,N_19633,N_17808);
nand U24044 (N_24044,N_15636,N_15487);
nor U24045 (N_24045,N_15695,N_16297);
and U24046 (N_24046,N_19877,N_16696);
nand U24047 (N_24047,N_15527,N_19151);
and U24048 (N_24048,N_15264,N_16050);
nand U24049 (N_24049,N_16524,N_19623);
nor U24050 (N_24050,N_18205,N_16559);
xor U24051 (N_24051,N_19817,N_15681);
or U24052 (N_24052,N_16013,N_18906);
and U24053 (N_24053,N_18567,N_16843);
nor U24054 (N_24054,N_16925,N_19618);
xnor U24055 (N_24055,N_18579,N_18602);
or U24056 (N_24056,N_16477,N_19022);
xnor U24057 (N_24057,N_19285,N_17552);
xor U24058 (N_24058,N_16604,N_19660);
nand U24059 (N_24059,N_15775,N_16061);
nand U24060 (N_24060,N_19825,N_16061);
or U24061 (N_24061,N_18662,N_19802);
and U24062 (N_24062,N_18845,N_18957);
or U24063 (N_24063,N_15677,N_19786);
xnor U24064 (N_24064,N_19957,N_17650);
nor U24065 (N_24065,N_19748,N_15542);
and U24066 (N_24066,N_16021,N_18672);
nand U24067 (N_24067,N_18032,N_16442);
and U24068 (N_24068,N_17890,N_16212);
nor U24069 (N_24069,N_15987,N_19932);
and U24070 (N_24070,N_19064,N_18574);
and U24071 (N_24071,N_16267,N_19548);
or U24072 (N_24072,N_17792,N_17871);
nand U24073 (N_24073,N_19084,N_18020);
nand U24074 (N_24074,N_16779,N_15607);
or U24075 (N_24075,N_17309,N_15754);
and U24076 (N_24076,N_19974,N_18685);
and U24077 (N_24077,N_16648,N_16982);
xor U24078 (N_24078,N_17960,N_15138);
xnor U24079 (N_24079,N_16463,N_15654);
or U24080 (N_24080,N_15494,N_19722);
and U24081 (N_24081,N_15121,N_15807);
nor U24082 (N_24082,N_19768,N_15407);
nand U24083 (N_24083,N_18479,N_19790);
nand U24084 (N_24084,N_16996,N_19569);
or U24085 (N_24085,N_17721,N_19691);
nand U24086 (N_24086,N_19712,N_17931);
xnor U24087 (N_24087,N_18422,N_16029);
xnor U24088 (N_24088,N_18184,N_16485);
xor U24089 (N_24089,N_18825,N_15574);
nor U24090 (N_24090,N_18895,N_18669);
xor U24091 (N_24091,N_19888,N_16101);
or U24092 (N_24092,N_16599,N_15117);
xnor U24093 (N_24093,N_16155,N_17556);
nand U24094 (N_24094,N_16181,N_16328);
nor U24095 (N_24095,N_16677,N_19192);
and U24096 (N_24096,N_15161,N_15163);
nand U24097 (N_24097,N_19402,N_18693);
nor U24098 (N_24098,N_18744,N_17133);
and U24099 (N_24099,N_19614,N_15874);
nor U24100 (N_24100,N_16788,N_16807);
nor U24101 (N_24101,N_18977,N_18844);
or U24102 (N_24102,N_18408,N_18264);
nand U24103 (N_24103,N_15058,N_16847);
or U24104 (N_24104,N_16163,N_15419);
or U24105 (N_24105,N_18262,N_19014);
xor U24106 (N_24106,N_15955,N_19398);
and U24107 (N_24107,N_16676,N_18248);
xnor U24108 (N_24108,N_18931,N_17363);
and U24109 (N_24109,N_18442,N_17798);
nand U24110 (N_24110,N_15125,N_18666);
nand U24111 (N_24111,N_15195,N_15084);
xnor U24112 (N_24112,N_15955,N_17523);
and U24113 (N_24113,N_19796,N_17885);
nand U24114 (N_24114,N_15454,N_18361);
nor U24115 (N_24115,N_15658,N_18667);
and U24116 (N_24116,N_16209,N_19102);
nor U24117 (N_24117,N_19551,N_17200);
or U24118 (N_24118,N_18576,N_18553);
and U24119 (N_24119,N_15197,N_16963);
and U24120 (N_24120,N_16975,N_17994);
or U24121 (N_24121,N_16586,N_17350);
xor U24122 (N_24122,N_18886,N_16563);
nand U24123 (N_24123,N_16514,N_16993);
or U24124 (N_24124,N_15894,N_19668);
or U24125 (N_24125,N_18336,N_16555);
or U24126 (N_24126,N_15544,N_16860);
and U24127 (N_24127,N_15208,N_18502);
nand U24128 (N_24128,N_16323,N_15545);
nor U24129 (N_24129,N_17963,N_19917);
and U24130 (N_24130,N_16335,N_18500);
and U24131 (N_24131,N_17067,N_15616);
or U24132 (N_24132,N_17978,N_16534);
or U24133 (N_24133,N_18754,N_19014);
xnor U24134 (N_24134,N_19487,N_18276);
nand U24135 (N_24135,N_18828,N_18479);
nand U24136 (N_24136,N_17751,N_16947);
nor U24137 (N_24137,N_19673,N_16954);
or U24138 (N_24138,N_19189,N_18021);
nand U24139 (N_24139,N_19704,N_17566);
or U24140 (N_24140,N_16256,N_17642);
xnor U24141 (N_24141,N_18952,N_16842);
nand U24142 (N_24142,N_19521,N_17838);
nor U24143 (N_24143,N_16511,N_16632);
or U24144 (N_24144,N_15517,N_17280);
nand U24145 (N_24145,N_15819,N_19432);
nor U24146 (N_24146,N_18764,N_17185);
nand U24147 (N_24147,N_18162,N_19767);
nor U24148 (N_24148,N_19983,N_17777);
xnor U24149 (N_24149,N_18007,N_18982);
or U24150 (N_24150,N_17928,N_15290);
and U24151 (N_24151,N_17768,N_15596);
or U24152 (N_24152,N_17544,N_17274);
nand U24153 (N_24153,N_18353,N_18555);
nor U24154 (N_24154,N_16777,N_15149);
nand U24155 (N_24155,N_18911,N_17688);
and U24156 (N_24156,N_16039,N_18422);
xnor U24157 (N_24157,N_16123,N_19154);
nor U24158 (N_24158,N_17650,N_19581);
or U24159 (N_24159,N_18761,N_15206);
and U24160 (N_24160,N_18744,N_17891);
and U24161 (N_24161,N_17727,N_16249);
or U24162 (N_24162,N_17047,N_16586);
xnor U24163 (N_24163,N_16882,N_18002);
and U24164 (N_24164,N_17622,N_18077);
nor U24165 (N_24165,N_15783,N_17302);
nand U24166 (N_24166,N_19093,N_18751);
or U24167 (N_24167,N_15229,N_16331);
and U24168 (N_24168,N_17907,N_16300);
or U24169 (N_24169,N_18575,N_16549);
and U24170 (N_24170,N_17477,N_15848);
and U24171 (N_24171,N_19211,N_16912);
nor U24172 (N_24172,N_16708,N_19909);
or U24173 (N_24173,N_17316,N_15941);
xor U24174 (N_24174,N_17464,N_18356);
nor U24175 (N_24175,N_16696,N_18401);
nand U24176 (N_24176,N_18993,N_18859);
and U24177 (N_24177,N_18186,N_19162);
xor U24178 (N_24178,N_19390,N_15768);
nor U24179 (N_24179,N_15943,N_16507);
or U24180 (N_24180,N_18186,N_17794);
or U24181 (N_24181,N_18349,N_15608);
xor U24182 (N_24182,N_18538,N_19798);
and U24183 (N_24183,N_17478,N_18592);
nand U24184 (N_24184,N_16647,N_15374);
and U24185 (N_24185,N_19805,N_18549);
or U24186 (N_24186,N_15576,N_19290);
nor U24187 (N_24187,N_19145,N_17158);
and U24188 (N_24188,N_17034,N_15246);
and U24189 (N_24189,N_17534,N_18813);
or U24190 (N_24190,N_18059,N_19090);
nor U24191 (N_24191,N_19593,N_19851);
nand U24192 (N_24192,N_15424,N_17906);
nand U24193 (N_24193,N_15951,N_17273);
or U24194 (N_24194,N_19213,N_18356);
nor U24195 (N_24195,N_16467,N_18433);
and U24196 (N_24196,N_18839,N_17766);
and U24197 (N_24197,N_16616,N_19665);
nand U24198 (N_24198,N_18069,N_15477);
or U24199 (N_24199,N_16740,N_17880);
and U24200 (N_24200,N_18957,N_17881);
xnor U24201 (N_24201,N_16808,N_15204);
nor U24202 (N_24202,N_19632,N_19754);
and U24203 (N_24203,N_15834,N_18244);
and U24204 (N_24204,N_19442,N_18731);
nor U24205 (N_24205,N_15908,N_15219);
nor U24206 (N_24206,N_15210,N_19106);
or U24207 (N_24207,N_19024,N_17635);
nand U24208 (N_24208,N_18548,N_19574);
and U24209 (N_24209,N_18741,N_17765);
nand U24210 (N_24210,N_17498,N_17265);
nand U24211 (N_24211,N_17833,N_15775);
nand U24212 (N_24212,N_15046,N_18707);
nor U24213 (N_24213,N_15547,N_17236);
nor U24214 (N_24214,N_18652,N_17629);
xnor U24215 (N_24215,N_19161,N_16593);
xnor U24216 (N_24216,N_18896,N_19296);
and U24217 (N_24217,N_19425,N_15919);
xor U24218 (N_24218,N_17412,N_19591);
xnor U24219 (N_24219,N_15059,N_17111);
nand U24220 (N_24220,N_16521,N_17459);
nand U24221 (N_24221,N_16215,N_18633);
nand U24222 (N_24222,N_15329,N_17142);
or U24223 (N_24223,N_18200,N_19889);
or U24224 (N_24224,N_17934,N_19557);
nor U24225 (N_24225,N_15937,N_15305);
nor U24226 (N_24226,N_19069,N_15416);
and U24227 (N_24227,N_19781,N_19313);
or U24228 (N_24228,N_19754,N_15024);
or U24229 (N_24229,N_19814,N_17052);
xnor U24230 (N_24230,N_15751,N_19916);
and U24231 (N_24231,N_16207,N_16599);
nor U24232 (N_24232,N_16342,N_19939);
or U24233 (N_24233,N_19500,N_16369);
nand U24234 (N_24234,N_15351,N_15885);
or U24235 (N_24235,N_16741,N_15261);
or U24236 (N_24236,N_18241,N_18851);
nor U24237 (N_24237,N_17175,N_19464);
nor U24238 (N_24238,N_19324,N_15892);
nand U24239 (N_24239,N_17548,N_18279);
and U24240 (N_24240,N_16728,N_16318);
xor U24241 (N_24241,N_18069,N_19651);
nand U24242 (N_24242,N_17337,N_19585);
or U24243 (N_24243,N_15612,N_17803);
nand U24244 (N_24244,N_16919,N_17701);
and U24245 (N_24245,N_18290,N_16411);
or U24246 (N_24246,N_16952,N_19366);
or U24247 (N_24247,N_18476,N_19759);
or U24248 (N_24248,N_18097,N_17945);
xnor U24249 (N_24249,N_19957,N_17068);
nor U24250 (N_24250,N_17509,N_18687);
xnor U24251 (N_24251,N_16315,N_19699);
or U24252 (N_24252,N_16818,N_19720);
or U24253 (N_24253,N_17095,N_16521);
nor U24254 (N_24254,N_16983,N_19116);
and U24255 (N_24255,N_18943,N_19419);
or U24256 (N_24256,N_15015,N_17070);
and U24257 (N_24257,N_17561,N_19352);
nand U24258 (N_24258,N_15948,N_16745);
or U24259 (N_24259,N_15742,N_16848);
xor U24260 (N_24260,N_15056,N_16717);
nor U24261 (N_24261,N_17020,N_16744);
nand U24262 (N_24262,N_15774,N_19917);
nor U24263 (N_24263,N_18482,N_16916);
xnor U24264 (N_24264,N_16293,N_15201);
xnor U24265 (N_24265,N_15443,N_17680);
or U24266 (N_24266,N_17261,N_15237);
nand U24267 (N_24267,N_17220,N_15022);
xor U24268 (N_24268,N_16365,N_18440);
xnor U24269 (N_24269,N_17841,N_15079);
or U24270 (N_24270,N_17501,N_18389);
and U24271 (N_24271,N_16527,N_16399);
and U24272 (N_24272,N_15764,N_18086);
or U24273 (N_24273,N_17334,N_15250);
nor U24274 (N_24274,N_16793,N_18797);
nor U24275 (N_24275,N_18036,N_17574);
nor U24276 (N_24276,N_15456,N_16489);
and U24277 (N_24277,N_18622,N_15749);
nor U24278 (N_24278,N_16875,N_17531);
xor U24279 (N_24279,N_18612,N_17854);
or U24280 (N_24280,N_17950,N_16751);
or U24281 (N_24281,N_17553,N_17261);
nor U24282 (N_24282,N_15012,N_17366);
and U24283 (N_24283,N_15992,N_19194);
xnor U24284 (N_24284,N_18567,N_16155);
nor U24285 (N_24285,N_19194,N_18900);
and U24286 (N_24286,N_19463,N_19294);
and U24287 (N_24287,N_15903,N_16850);
xor U24288 (N_24288,N_16159,N_15318);
and U24289 (N_24289,N_17325,N_15267);
nor U24290 (N_24290,N_16706,N_19672);
or U24291 (N_24291,N_17835,N_18548);
and U24292 (N_24292,N_16965,N_19201);
nor U24293 (N_24293,N_16800,N_15919);
or U24294 (N_24294,N_19756,N_17167);
xnor U24295 (N_24295,N_18386,N_17555);
and U24296 (N_24296,N_16644,N_15758);
nand U24297 (N_24297,N_18459,N_16603);
or U24298 (N_24298,N_17813,N_19624);
nor U24299 (N_24299,N_18971,N_15113);
xor U24300 (N_24300,N_18092,N_16962);
nand U24301 (N_24301,N_17041,N_16221);
xor U24302 (N_24302,N_18854,N_17012);
nand U24303 (N_24303,N_15432,N_17410);
nand U24304 (N_24304,N_16159,N_19984);
or U24305 (N_24305,N_18203,N_19237);
nand U24306 (N_24306,N_17865,N_18045);
and U24307 (N_24307,N_19758,N_15504);
nor U24308 (N_24308,N_19660,N_17458);
and U24309 (N_24309,N_17464,N_17572);
nand U24310 (N_24310,N_17237,N_19464);
or U24311 (N_24311,N_19625,N_16685);
and U24312 (N_24312,N_15028,N_16389);
xor U24313 (N_24313,N_18809,N_19255);
nand U24314 (N_24314,N_18292,N_15519);
or U24315 (N_24315,N_19988,N_16326);
xnor U24316 (N_24316,N_16423,N_18262);
and U24317 (N_24317,N_17777,N_15433);
or U24318 (N_24318,N_19165,N_15875);
nor U24319 (N_24319,N_15684,N_17742);
nand U24320 (N_24320,N_16470,N_17758);
nor U24321 (N_24321,N_16159,N_19222);
nor U24322 (N_24322,N_15281,N_16025);
nand U24323 (N_24323,N_18147,N_19134);
nor U24324 (N_24324,N_18075,N_19873);
and U24325 (N_24325,N_18085,N_15443);
nor U24326 (N_24326,N_15594,N_17927);
and U24327 (N_24327,N_17546,N_19615);
and U24328 (N_24328,N_18333,N_18450);
xnor U24329 (N_24329,N_16953,N_16127);
xnor U24330 (N_24330,N_15360,N_16048);
nor U24331 (N_24331,N_17684,N_18102);
xor U24332 (N_24332,N_18850,N_19554);
nor U24333 (N_24333,N_16290,N_17214);
xnor U24334 (N_24334,N_17980,N_19891);
xnor U24335 (N_24335,N_17865,N_17102);
or U24336 (N_24336,N_15705,N_18161);
or U24337 (N_24337,N_18075,N_15793);
xnor U24338 (N_24338,N_15996,N_16059);
xor U24339 (N_24339,N_15275,N_18263);
nor U24340 (N_24340,N_17310,N_15488);
and U24341 (N_24341,N_19504,N_17576);
and U24342 (N_24342,N_19429,N_19914);
and U24343 (N_24343,N_17319,N_17659);
nor U24344 (N_24344,N_19389,N_15947);
nor U24345 (N_24345,N_17991,N_17083);
xnor U24346 (N_24346,N_19672,N_16880);
xor U24347 (N_24347,N_16688,N_17317);
nand U24348 (N_24348,N_15779,N_16807);
and U24349 (N_24349,N_15756,N_15394);
and U24350 (N_24350,N_18595,N_16280);
and U24351 (N_24351,N_19857,N_19052);
nand U24352 (N_24352,N_17611,N_17590);
nand U24353 (N_24353,N_18205,N_17377);
nand U24354 (N_24354,N_15831,N_16004);
and U24355 (N_24355,N_18362,N_16054);
xor U24356 (N_24356,N_15599,N_19854);
or U24357 (N_24357,N_17013,N_15346);
xnor U24358 (N_24358,N_19907,N_17792);
and U24359 (N_24359,N_17349,N_18045);
nand U24360 (N_24360,N_19993,N_17342);
xnor U24361 (N_24361,N_16749,N_17960);
nor U24362 (N_24362,N_17781,N_18230);
xor U24363 (N_24363,N_19158,N_16186);
nor U24364 (N_24364,N_16896,N_16479);
nand U24365 (N_24365,N_17009,N_19047);
nor U24366 (N_24366,N_18274,N_17517);
nand U24367 (N_24367,N_17624,N_15744);
nor U24368 (N_24368,N_18690,N_17870);
xnor U24369 (N_24369,N_16975,N_15378);
nand U24370 (N_24370,N_15049,N_18425);
nand U24371 (N_24371,N_19710,N_18366);
or U24372 (N_24372,N_19143,N_15546);
nand U24373 (N_24373,N_16834,N_18464);
and U24374 (N_24374,N_15384,N_17549);
nor U24375 (N_24375,N_16440,N_15610);
nor U24376 (N_24376,N_18246,N_16822);
nor U24377 (N_24377,N_18313,N_18698);
nand U24378 (N_24378,N_16868,N_16276);
xor U24379 (N_24379,N_15053,N_19726);
xor U24380 (N_24380,N_19235,N_15762);
and U24381 (N_24381,N_18354,N_15870);
and U24382 (N_24382,N_19730,N_19747);
xor U24383 (N_24383,N_18424,N_17638);
nand U24384 (N_24384,N_17337,N_15124);
xnor U24385 (N_24385,N_19535,N_16538);
xnor U24386 (N_24386,N_18609,N_15905);
nor U24387 (N_24387,N_15812,N_17175);
nor U24388 (N_24388,N_16616,N_16655);
nor U24389 (N_24389,N_18688,N_19809);
or U24390 (N_24390,N_18045,N_18276);
nand U24391 (N_24391,N_19158,N_18632);
nor U24392 (N_24392,N_17410,N_15839);
nor U24393 (N_24393,N_19277,N_15820);
or U24394 (N_24394,N_19254,N_19367);
and U24395 (N_24395,N_17690,N_16087);
or U24396 (N_24396,N_16013,N_18066);
or U24397 (N_24397,N_19949,N_17690);
xor U24398 (N_24398,N_19808,N_18570);
nor U24399 (N_24399,N_16085,N_17068);
nor U24400 (N_24400,N_16962,N_15643);
nand U24401 (N_24401,N_18864,N_19514);
or U24402 (N_24402,N_15662,N_17645);
nor U24403 (N_24403,N_15609,N_15799);
and U24404 (N_24404,N_17212,N_16584);
xnor U24405 (N_24405,N_18326,N_19746);
and U24406 (N_24406,N_18478,N_16797);
nand U24407 (N_24407,N_17038,N_16648);
xor U24408 (N_24408,N_19951,N_16692);
xnor U24409 (N_24409,N_19522,N_15351);
or U24410 (N_24410,N_17554,N_19458);
xnor U24411 (N_24411,N_18901,N_19325);
or U24412 (N_24412,N_18943,N_19423);
xor U24413 (N_24413,N_16334,N_17151);
or U24414 (N_24414,N_18000,N_16467);
or U24415 (N_24415,N_18566,N_15527);
or U24416 (N_24416,N_18174,N_15288);
or U24417 (N_24417,N_16433,N_16000);
xor U24418 (N_24418,N_15216,N_15688);
nand U24419 (N_24419,N_19892,N_17633);
or U24420 (N_24420,N_18939,N_16669);
and U24421 (N_24421,N_15235,N_15847);
xor U24422 (N_24422,N_17447,N_16953);
xnor U24423 (N_24423,N_19781,N_17429);
nor U24424 (N_24424,N_19934,N_16650);
xnor U24425 (N_24425,N_19847,N_16758);
xor U24426 (N_24426,N_18769,N_19762);
nand U24427 (N_24427,N_16617,N_19665);
nor U24428 (N_24428,N_17118,N_17334);
or U24429 (N_24429,N_16610,N_15442);
and U24430 (N_24430,N_16477,N_15090);
nand U24431 (N_24431,N_19928,N_16417);
nand U24432 (N_24432,N_17341,N_15032);
nor U24433 (N_24433,N_16431,N_17320);
nand U24434 (N_24434,N_16944,N_17960);
or U24435 (N_24435,N_18458,N_15527);
and U24436 (N_24436,N_19740,N_15528);
xor U24437 (N_24437,N_16876,N_16665);
nor U24438 (N_24438,N_19273,N_16037);
and U24439 (N_24439,N_15630,N_18308);
nor U24440 (N_24440,N_17074,N_17429);
xor U24441 (N_24441,N_17154,N_17783);
xnor U24442 (N_24442,N_19692,N_16412);
nor U24443 (N_24443,N_17975,N_16408);
nor U24444 (N_24444,N_19628,N_17889);
nand U24445 (N_24445,N_17077,N_19742);
and U24446 (N_24446,N_16906,N_15151);
xor U24447 (N_24447,N_18214,N_18450);
nor U24448 (N_24448,N_15243,N_19494);
and U24449 (N_24449,N_19942,N_19347);
and U24450 (N_24450,N_15694,N_19769);
and U24451 (N_24451,N_16235,N_17540);
and U24452 (N_24452,N_15132,N_16788);
and U24453 (N_24453,N_16708,N_17508);
nand U24454 (N_24454,N_18971,N_15661);
nor U24455 (N_24455,N_16946,N_16134);
nand U24456 (N_24456,N_17944,N_16769);
xnor U24457 (N_24457,N_16389,N_15053);
and U24458 (N_24458,N_17099,N_16359);
nand U24459 (N_24459,N_18878,N_19023);
and U24460 (N_24460,N_16779,N_19901);
nand U24461 (N_24461,N_17510,N_15726);
nand U24462 (N_24462,N_18926,N_15722);
or U24463 (N_24463,N_17786,N_17566);
or U24464 (N_24464,N_15952,N_15791);
or U24465 (N_24465,N_17946,N_19263);
or U24466 (N_24466,N_19614,N_19409);
and U24467 (N_24467,N_16640,N_16201);
nor U24468 (N_24468,N_18217,N_16149);
and U24469 (N_24469,N_15685,N_17236);
nor U24470 (N_24470,N_17490,N_16310);
nor U24471 (N_24471,N_16573,N_15683);
nand U24472 (N_24472,N_16638,N_17134);
nand U24473 (N_24473,N_17842,N_18617);
xor U24474 (N_24474,N_17649,N_18090);
or U24475 (N_24475,N_18381,N_19262);
xnor U24476 (N_24476,N_18077,N_16376);
xor U24477 (N_24477,N_18396,N_19769);
nor U24478 (N_24478,N_18238,N_18467);
nand U24479 (N_24479,N_16487,N_18855);
nand U24480 (N_24480,N_15545,N_17245);
nor U24481 (N_24481,N_19820,N_16848);
and U24482 (N_24482,N_15700,N_16899);
nand U24483 (N_24483,N_19934,N_19891);
or U24484 (N_24484,N_18222,N_19674);
and U24485 (N_24485,N_17604,N_19217);
or U24486 (N_24486,N_15935,N_18937);
nor U24487 (N_24487,N_16270,N_16609);
xnor U24488 (N_24488,N_16619,N_17462);
and U24489 (N_24489,N_18900,N_17524);
xnor U24490 (N_24490,N_16850,N_16914);
nand U24491 (N_24491,N_17083,N_17421);
or U24492 (N_24492,N_16635,N_17822);
xor U24493 (N_24493,N_15108,N_17611);
and U24494 (N_24494,N_16145,N_19477);
or U24495 (N_24495,N_16645,N_18618);
and U24496 (N_24496,N_18406,N_15600);
xor U24497 (N_24497,N_16769,N_18345);
and U24498 (N_24498,N_18621,N_19786);
nor U24499 (N_24499,N_19278,N_17014);
nand U24500 (N_24500,N_16708,N_17502);
xor U24501 (N_24501,N_17146,N_16561);
xor U24502 (N_24502,N_17406,N_15070);
nor U24503 (N_24503,N_17364,N_18803);
or U24504 (N_24504,N_18617,N_16143);
nor U24505 (N_24505,N_17117,N_18441);
xnor U24506 (N_24506,N_19993,N_19454);
and U24507 (N_24507,N_19397,N_15418);
or U24508 (N_24508,N_19189,N_15273);
nand U24509 (N_24509,N_16672,N_18422);
and U24510 (N_24510,N_17605,N_15325);
or U24511 (N_24511,N_15159,N_19971);
and U24512 (N_24512,N_16621,N_16083);
and U24513 (N_24513,N_15719,N_15609);
or U24514 (N_24514,N_19714,N_16808);
and U24515 (N_24515,N_16120,N_17049);
nor U24516 (N_24516,N_16705,N_17402);
xnor U24517 (N_24517,N_15081,N_16585);
and U24518 (N_24518,N_17173,N_16739);
or U24519 (N_24519,N_18776,N_15063);
nand U24520 (N_24520,N_18564,N_17434);
and U24521 (N_24521,N_16683,N_19795);
or U24522 (N_24522,N_19871,N_18070);
nand U24523 (N_24523,N_15597,N_17568);
nand U24524 (N_24524,N_15034,N_17276);
nand U24525 (N_24525,N_16531,N_19410);
xnor U24526 (N_24526,N_17837,N_16039);
and U24527 (N_24527,N_15510,N_16227);
nand U24528 (N_24528,N_15319,N_18932);
xor U24529 (N_24529,N_18825,N_17058);
xnor U24530 (N_24530,N_19898,N_19617);
or U24531 (N_24531,N_15814,N_19751);
or U24532 (N_24532,N_17749,N_18644);
or U24533 (N_24533,N_15403,N_16134);
or U24534 (N_24534,N_19320,N_19622);
nor U24535 (N_24535,N_15002,N_18721);
nor U24536 (N_24536,N_15504,N_16229);
and U24537 (N_24537,N_17390,N_19531);
xnor U24538 (N_24538,N_17818,N_15923);
or U24539 (N_24539,N_16130,N_15002);
and U24540 (N_24540,N_16424,N_15389);
nor U24541 (N_24541,N_15263,N_18251);
nand U24542 (N_24542,N_18832,N_18117);
and U24543 (N_24543,N_19419,N_19948);
or U24544 (N_24544,N_17129,N_15838);
xor U24545 (N_24545,N_16913,N_19018);
xor U24546 (N_24546,N_15705,N_16577);
nor U24547 (N_24547,N_17055,N_15992);
xor U24548 (N_24548,N_18020,N_19390);
and U24549 (N_24549,N_15572,N_19396);
xor U24550 (N_24550,N_18000,N_15687);
nor U24551 (N_24551,N_18766,N_19797);
nor U24552 (N_24552,N_19632,N_16914);
xnor U24553 (N_24553,N_18597,N_17466);
xor U24554 (N_24554,N_17343,N_17437);
or U24555 (N_24555,N_19312,N_18518);
or U24556 (N_24556,N_19312,N_17409);
nor U24557 (N_24557,N_16957,N_16517);
nor U24558 (N_24558,N_16444,N_16920);
nor U24559 (N_24559,N_17587,N_17028);
and U24560 (N_24560,N_16883,N_15745);
xnor U24561 (N_24561,N_15356,N_18519);
and U24562 (N_24562,N_16858,N_18195);
nor U24563 (N_24563,N_17338,N_18312);
nand U24564 (N_24564,N_17326,N_17583);
or U24565 (N_24565,N_18092,N_16819);
xor U24566 (N_24566,N_16021,N_15324);
and U24567 (N_24567,N_17877,N_15774);
nand U24568 (N_24568,N_17612,N_19529);
nand U24569 (N_24569,N_16626,N_17550);
nand U24570 (N_24570,N_19267,N_18160);
xor U24571 (N_24571,N_15896,N_17754);
xor U24572 (N_24572,N_16604,N_15607);
or U24573 (N_24573,N_17495,N_16373);
nor U24574 (N_24574,N_18957,N_18013);
or U24575 (N_24575,N_16517,N_19058);
and U24576 (N_24576,N_15171,N_17163);
or U24577 (N_24577,N_17942,N_15634);
and U24578 (N_24578,N_15648,N_18307);
xnor U24579 (N_24579,N_18953,N_17733);
nor U24580 (N_24580,N_19576,N_18354);
nor U24581 (N_24581,N_15817,N_16386);
and U24582 (N_24582,N_15678,N_19996);
or U24583 (N_24583,N_17280,N_19573);
nand U24584 (N_24584,N_15220,N_17553);
nor U24585 (N_24585,N_15168,N_15811);
nor U24586 (N_24586,N_18876,N_16387);
nand U24587 (N_24587,N_16934,N_16309);
xnor U24588 (N_24588,N_16120,N_17605);
nor U24589 (N_24589,N_15687,N_15041);
nor U24590 (N_24590,N_19838,N_15301);
and U24591 (N_24591,N_16795,N_18405);
xor U24592 (N_24592,N_18279,N_15138);
nand U24593 (N_24593,N_16416,N_16498);
or U24594 (N_24594,N_16936,N_15168);
nor U24595 (N_24595,N_16521,N_19543);
nand U24596 (N_24596,N_15516,N_18311);
and U24597 (N_24597,N_19907,N_16668);
and U24598 (N_24598,N_17501,N_19273);
nor U24599 (N_24599,N_16903,N_17997);
or U24600 (N_24600,N_18990,N_15612);
nand U24601 (N_24601,N_18499,N_16506);
nor U24602 (N_24602,N_18974,N_16337);
nor U24603 (N_24603,N_17767,N_19159);
nand U24604 (N_24604,N_19054,N_18469);
xor U24605 (N_24605,N_19769,N_15662);
and U24606 (N_24606,N_18117,N_16051);
nand U24607 (N_24607,N_18507,N_16482);
and U24608 (N_24608,N_18873,N_16815);
or U24609 (N_24609,N_19821,N_18764);
xnor U24610 (N_24610,N_18889,N_18169);
or U24611 (N_24611,N_15145,N_18470);
nand U24612 (N_24612,N_19648,N_16974);
nand U24613 (N_24613,N_17237,N_17046);
and U24614 (N_24614,N_19006,N_18633);
nand U24615 (N_24615,N_17513,N_19288);
xnor U24616 (N_24616,N_19032,N_19002);
nand U24617 (N_24617,N_16501,N_18409);
nand U24618 (N_24618,N_15503,N_18099);
or U24619 (N_24619,N_15746,N_16102);
nand U24620 (N_24620,N_19792,N_18202);
or U24621 (N_24621,N_17763,N_16024);
nand U24622 (N_24622,N_17261,N_18084);
nor U24623 (N_24623,N_18917,N_15774);
or U24624 (N_24624,N_15534,N_16556);
nand U24625 (N_24625,N_18946,N_19902);
and U24626 (N_24626,N_16728,N_19485);
nand U24627 (N_24627,N_15531,N_15728);
nor U24628 (N_24628,N_17740,N_17377);
nor U24629 (N_24629,N_18071,N_18983);
and U24630 (N_24630,N_18499,N_16450);
xnor U24631 (N_24631,N_19404,N_18396);
nor U24632 (N_24632,N_17842,N_19790);
or U24633 (N_24633,N_18353,N_19705);
nand U24634 (N_24634,N_19662,N_19275);
xnor U24635 (N_24635,N_19345,N_19890);
nor U24636 (N_24636,N_15276,N_19304);
nand U24637 (N_24637,N_17160,N_15428);
nand U24638 (N_24638,N_15904,N_19257);
nor U24639 (N_24639,N_18503,N_18601);
or U24640 (N_24640,N_19855,N_16117);
xnor U24641 (N_24641,N_16320,N_16712);
or U24642 (N_24642,N_19211,N_17796);
or U24643 (N_24643,N_16169,N_18462);
and U24644 (N_24644,N_18024,N_17002);
or U24645 (N_24645,N_15963,N_17006);
nor U24646 (N_24646,N_17175,N_15488);
or U24647 (N_24647,N_16558,N_15887);
and U24648 (N_24648,N_17187,N_16825);
nand U24649 (N_24649,N_18343,N_17157);
xnor U24650 (N_24650,N_15200,N_17353);
nor U24651 (N_24651,N_17256,N_18483);
nand U24652 (N_24652,N_18741,N_19953);
and U24653 (N_24653,N_19681,N_18361);
nand U24654 (N_24654,N_19325,N_18309);
and U24655 (N_24655,N_17430,N_18801);
nor U24656 (N_24656,N_16216,N_18385);
nand U24657 (N_24657,N_15785,N_15410);
nand U24658 (N_24658,N_18739,N_18628);
nor U24659 (N_24659,N_19472,N_19729);
and U24660 (N_24660,N_16416,N_17263);
or U24661 (N_24661,N_17969,N_19382);
nand U24662 (N_24662,N_16136,N_18252);
nor U24663 (N_24663,N_19261,N_16922);
or U24664 (N_24664,N_15614,N_16518);
nand U24665 (N_24665,N_17809,N_16477);
and U24666 (N_24666,N_18631,N_19912);
and U24667 (N_24667,N_15304,N_15218);
or U24668 (N_24668,N_17489,N_19444);
and U24669 (N_24669,N_18260,N_15459);
xor U24670 (N_24670,N_18246,N_15105);
nor U24671 (N_24671,N_19671,N_16784);
and U24672 (N_24672,N_19820,N_16783);
xnor U24673 (N_24673,N_16477,N_18361);
and U24674 (N_24674,N_19360,N_16243);
nor U24675 (N_24675,N_16211,N_15787);
or U24676 (N_24676,N_18971,N_17667);
nand U24677 (N_24677,N_15919,N_17747);
or U24678 (N_24678,N_19239,N_18828);
and U24679 (N_24679,N_15771,N_15106);
nor U24680 (N_24680,N_18317,N_16704);
or U24681 (N_24681,N_18553,N_19931);
nor U24682 (N_24682,N_18590,N_17953);
xor U24683 (N_24683,N_16121,N_16018);
xor U24684 (N_24684,N_19334,N_19229);
or U24685 (N_24685,N_19146,N_18683);
xnor U24686 (N_24686,N_17529,N_15542);
nor U24687 (N_24687,N_19611,N_19123);
and U24688 (N_24688,N_15060,N_18743);
nor U24689 (N_24689,N_18196,N_17940);
or U24690 (N_24690,N_19866,N_17394);
and U24691 (N_24691,N_18398,N_16773);
or U24692 (N_24692,N_17183,N_15153);
and U24693 (N_24693,N_19789,N_19191);
and U24694 (N_24694,N_17348,N_16316);
nor U24695 (N_24695,N_18516,N_15727);
and U24696 (N_24696,N_16773,N_19958);
xnor U24697 (N_24697,N_15864,N_19056);
nand U24698 (N_24698,N_15153,N_18460);
nand U24699 (N_24699,N_19842,N_16209);
or U24700 (N_24700,N_17251,N_17383);
nor U24701 (N_24701,N_16923,N_15823);
xnor U24702 (N_24702,N_16261,N_17414);
and U24703 (N_24703,N_17868,N_16308);
nor U24704 (N_24704,N_15781,N_17974);
nand U24705 (N_24705,N_18254,N_16424);
and U24706 (N_24706,N_15751,N_15496);
nor U24707 (N_24707,N_16419,N_17181);
nor U24708 (N_24708,N_18187,N_19037);
xnor U24709 (N_24709,N_17870,N_19532);
xnor U24710 (N_24710,N_17554,N_19420);
or U24711 (N_24711,N_15618,N_19147);
and U24712 (N_24712,N_17282,N_19573);
xnor U24713 (N_24713,N_19181,N_17919);
or U24714 (N_24714,N_19579,N_19151);
nand U24715 (N_24715,N_15402,N_16146);
nor U24716 (N_24716,N_19413,N_15199);
or U24717 (N_24717,N_18310,N_19358);
nand U24718 (N_24718,N_19417,N_15745);
and U24719 (N_24719,N_17315,N_18532);
nor U24720 (N_24720,N_18510,N_19872);
nor U24721 (N_24721,N_18689,N_15050);
xor U24722 (N_24722,N_18775,N_16834);
nand U24723 (N_24723,N_17963,N_17603);
xnor U24724 (N_24724,N_16898,N_15340);
nand U24725 (N_24725,N_15656,N_19745);
nor U24726 (N_24726,N_18970,N_17903);
or U24727 (N_24727,N_17890,N_18806);
nor U24728 (N_24728,N_19132,N_17960);
nor U24729 (N_24729,N_15078,N_17266);
nor U24730 (N_24730,N_17630,N_15234);
nand U24731 (N_24731,N_17077,N_18716);
or U24732 (N_24732,N_15167,N_16371);
or U24733 (N_24733,N_16293,N_18903);
xnor U24734 (N_24734,N_17527,N_16445);
nor U24735 (N_24735,N_16114,N_18214);
nor U24736 (N_24736,N_19605,N_17762);
nor U24737 (N_24737,N_16961,N_16275);
nor U24738 (N_24738,N_17081,N_18696);
nor U24739 (N_24739,N_16544,N_18066);
xnor U24740 (N_24740,N_19191,N_15398);
nor U24741 (N_24741,N_16309,N_18662);
nand U24742 (N_24742,N_18814,N_19485);
xnor U24743 (N_24743,N_19673,N_16073);
nor U24744 (N_24744,N_16317,N_16230);
xnor U24745 (N_24745,N_18860,N_17112);
or U24746 (N_24746,N_17588,N_17600);
nand U24747 (N_24747,N_15829,N_19770);
nand U24748 (N_24748,N_19350,N_17698);
and U24749 (N_24749,N_19711,N_18534);
nor U24750 (N_24750,N_19205,N_16446);
and U24751 (N_24751,N_19953,N_15963);
nand U24752 (N_24752,N_19153,N_16626);
xnor U24753 (N_24753,N_18454,N_19014);
and U24754 (N_24754,N_18924,N_17003);
xnor U24755 (N_24755,N_19551,N_18110);
nor U24756 (N_24756,N_18197,N_19872);
or U24757 (N_24757,N_19779,N_19496);
or U24758 (N_24758,N_17372,N_17012);
and U24759 (N_24759,N_19798,N_16758);
xnor U24760 (N_24760,N_17459,N_15504);
and U24761 (N_24761,N_16773,N_15183);
nand U24762 (N_24762,N_16600,N_17152);
or U24763 (N_24763,N_18830,N_17143);
or U24764 (N_24764,N_17328,N_18632);
and U24765 (N_24765,N_15357,N_19830);
nand U24766 (N_24766,N_17215,N_19226);
or U24767 (N_24767,N_17149,N_17190);
and U24768 (N_24768,N_18488,N_18723);
and U24769 (N_24769,N_15157,N_17632);
nand U24770 (N_24770,N_16665,N_15257);
nand U24771 (N_24771,N_17871,N_16466);
nor U24772 (N_24772,N_18078,N_16952);
nand U24773 (N_24773,N_18616,N_15213);
nor U24774 (N_24774,N_19440,N_17963);
or U24775 (N_24775,N_18880,N_18227);
nor U24776 (N_24776,N_19186,N_19255);
nor U24777 (N_24777,N_17561,N_19016);
and U24778 (N_24778,N_16435,N_18001);
or U24779 (N_24779,N_17278,N_15238);
or U24780 (N_24780,N_18324,N_17875);
and U24781 (N_24781,N_16447,N_16093);
nand U24782 (N_24782,N_17524,N_18205);
and U24783 (N_24783,N_15180,N_16987);
nand U24784 (N_24784,N_17548,N_16111);
xnor U24785 (N_24785,N_18122,N_18088);
and U24786 (N_24786,N_17590,N_15204);
and U24787 (N_24787,N_15415,N_18068);
nand U24788 (N_24788,N_18604,N_16840);
xnor U24789 (N_24789,N_17223,N_16218);
xnor U24790 (N_24790,N_18835,N_16355);
nor U24791 (N_24791,N_18216,N_15582);
nand U24792 (N_24792,N_15938,N_18095);
nor U24793 (N_24793,N_18928,N_15424);
and U24794 (N_24794,N_15759,N_18202);
and U24795 (N_24795,N_19518,N_19574);
or U24796 (N_24796,N_18904,N_15996);
and U24797 (N_24797,N_15885,N_17586);
and U24798 (N_24798,N_18717,N_17738);
and U24799 (N_24799,N_17039,N_18017);
nand U24800 (N_24800,N_17510,N_15532);
and U24801 (N_24801,N_15599,N_19789);
xor U24802 (N_24802,N_19537,N_17111);
xnor U24803 (N_24803,N_15504,N_18620);
and U24804 (N_24804,N_18992,N_15493);
xor U24805 (N_24805,N_15939,N_19204);
and U24806 (N_24806,N_15301,N_18714);
xor U24807 (N_24807,N_19225,N_17730);
or U24808 (N_24808,N_17825,N_18985);
and U24809 (N_24809,N_15786,N_15570);
or U24810 (N_24810,N_15958,N_16245);
and U24811 (N_24811,N_19686,N_16816);
xor U24812 (N_24812,N_15384,N_17954);
nand U24813 (N_24813,N_16541,N_19343);
or U24814 (N_24814,N_19991,N_16050);
and U24815 (N_24815,N_18431,N_15005);
nand U24816 (N_24816,N_15537,N_18721);
nor U24817 (N_24817,N_17567,N_18993);
or U24818 (N_24818,N_19744,N_17743);
nor U24819 (N_24819,N_15643,N_17732);
xnor U24820 (N_24820,N_18544,N_15259);
nor U24821 (N_24821,N_15346,N_19154);
or U24822 (N_24822,N_18737,N_18079);
or U24823 (N_24823,N_16145,N_15213);
nand U24824 (N_24824,N_18809,N_17548);
nand U24825 (N_24825,N_17771,N_16222);
nand U24826 (N_24826,N_17897,N_15549);
and U24827 (N_24827,N_18489,N_18400);
and U24828 (N_24828,N_19703,N_16231);
and U24829 (N_24829,N_17091,N_19645);
nand U24830 (N_24830,N_17603,N_15743);
and U24831 (N_24831,N_19541,N_15758);
or U24832 (N_24832,N_17358,N_15217);
and U24833 (N_24833,N_17219,N_17701);
xnor U24834 (N_24834,N_19877,N_15850);
or U24835 (N_24835,N_19966,N_19205);
nand U24836 (N_24836,N_18687,N_18066);
nor U24837 (N_24837,N_16627,N_18775);
or U24838 (N_24838,N_18531,N_15337);
or U24839 (N_24839,N_19554,N_16357);
or U24840 (N_24840,N_18157,N_17373);
xnor U24841 (N_24841,N_15881,N_18314);
nor U24842 (N_24842,N_16048,N_16366);
nand U24843 (N_24843,N_18360,N_19891);
nor U24844 (N_24844,N_15166,N_19252);
nand U24845 (N_24845,N_16517,N_16219);
nor U24846 (N_24846,N_17568,N_18720);
xor U24847 (N_24847,N_17132,N_15134);
and U24848 (N_24848,N_15461,N_15911);
nand U24849 (N_24849,N_19777,N_16851);
nor U24850 (N_24850,N_15388,N_19912);
and U24851 (N_24851,N_17107,N_16258);
and U24852 (N_24852,N_17225,N_19547);
or U24853 (N_24853,N_15148,N_18918);
nand U24854 (N_24854,N_18278,N_17146);
xor U24855 (N_24855,N_17468,N_19097);
or U24856 (N_24856,N_15121,N_19063);
and U24857 (N_24857,N_18766,N_19192);
and U24858 (N_24858,N_19935,N_15491);
xnor U24859 (N_24859,N_15616,N_16760);
nand U24860 (N_24860,N_18632,N_15962);
xnor U24861 (N_24861,N_16692,N_18299);
or U24862 (N_24862,N_16016,N_15307);
or U24863 (N_24863,N_19352,N_15793);
or U24864 (N_24864,N_17489,N_19133);
nor U24865 (N_24865,N_18083,N_17050);
xor U24866 (N_24866,N_17525,N_15215);
nor U24867 (N_24867,N_15141,N_17544);
or U24868 (N_24868,N_19908,N_16599);
nand U24869 (N_24869,N_15403,N_15397);
nand U24870 (N_24870,N_15082,N_17046);
nor U24871 (N_24871,N_19959,N_16584);
or U24872 (N_24872,N_15882,N_17919);
nand U24873 (N_24873,N_15480,N_18526);
xor U24874 (N_24874,N_15141,N_18932);
and U24875 (N_24875,N_19807,N_16532);
nor U24876 (N_24876,N_18950,N_16709);
and U24877 (N_24877,N_18924,N_18026);
or U24878 (N_24878,N_17474,N_18645);
xor U24879 (N_24879,N_18438,N_17485);
nand U24880 (N_24880,N_18791,N_16495);
xor U24881 (N_24881,N_15366,N_18416);
xor U24882 (N_24882,N_15952,N_18503);
or U24883 (N_24883,N_16284,N_17812);
and U24884 (N_24884,N_17002,N_18563);
and U24885 (N_24885,N_16680,N_15294);
or U24886 (N_24886,N_15237,N_15385);
nand U24887 (N_24887,N_17657,N_16053);
nand U24888 (N_24888,N_18634,N_17584);
or U24889 (N_24889,N_15492,N_15056);
nor U24890 (N_24890,N_15699,N_16464);
nand U24891 (N_24891,N_16991,N_19136);
and U24892 (N_24892,N_16187,N_15847);
and U24893 (N_24893,N_17300,N_18812);
xnor U24894 (N_24894,N_19566,N_17070);
nand U24895 (N_24895,N_15987,N_15846);
nor U24896 (N_24896,N_19589,N_18234);
nor U24897 (N_24897,N_16110,N_15798);
xnor U24898 (N_24898,N_19866,N_15478);
nand U24899 (N_24899,N_18038,N_19811);
nand U24900 (N_24900,N_17549,N_15584);
nand U24901 (N_24901,N_16829,N_15588);
or U24902 (N_24902,N_15252,N_17526);
nand U24903 (N_24903,N_17457,N_16168);
nor U24904 (N_24904,N_18204,N_17343);
or U24905 (N_24905,N_17672,N_16510);
or U24906 (N_24906,N_16221,N_18384);
or U24907 (N_24907,N_15709,N_16544);
nor U24908 (N_24908,N_18255,N_19372);
or U24909 (N_24909,N_16153,N_16626);
xor U24910 (N_24910,N_19286,N_17146);
xnor U24911 (N_24911,N_19539,N_18923);
nand U24912 (N_24912,N_15654,N_17986);
nor U24913 (N_24913,N_18370,N_18137);
and U24914 (N_24914,N_19791,N_19259);
nor U24915 (N_24915,N_18684,N_15559);
nor U24916 (N_24916,N_19023,N_18158);
nand U24917 (N_24917,N_15971,N_18467);
nor U24918 (N_24918,N_16589,N_19976);
xor U24919 (N_24919,N_17098,N_19146);
nor U24920 (N_24920,N_19161,N_16984);
nand U24921 (N_24921,N_15457,N_15893);
nor U24922 (N_24922,N_19061,N_17631);
and U24923 (N_24923,N_18071,N_19371);
nand U24924 (N_24924,N_18910,N_18024);
and U24925 (N_24925,N_18119,N_19463);
and U24926 (N_24926,N_17552,N_19309);
or U24927 (N_24927,N_17922,N_18701);
and U24928 (N_24928,N_17947,N_19193);
or U24929 (N_24929,N_15483,N_15023);
nor U24930 (N_24930,N_16814,N_16922);
or U24931 (N_24931,N_16839,N_16681);
nand U24932 (N_24932,N_18620,N_16774);
xor U24933 (N_24933,N_16680,N_17254);
nor U24934 (N_24934,N_17481,N_17883);
or U24935 (N_24935,N_19616,N_18006);
xnor U24936 (N_24936,N_18765,N_17986);
and U24937 (N_24937,N_18827,N_19090);
or U24938 (N_24938,N_19334,N_16295);
nand U24939 (N_24939,N_18602,N_18561);
and U24940 (N_24940,N_18568,N_15113);
and U24941 (N_24941,N_19301,N_17497);
xnor U24942 (N_24942,N_18401,N_19043);
or U24943 (N_24943,N_18096,N_15125);
or U24944 (N_24944,N_17991,N_18944);
or U24945 (N_24945,N_18211,N_18378);
and U24946 (N_24946,N_18817,N_18755);
nor U24947 (N_24947,N_19410,N_16232);
or U24948 (N_24948,N_17452,N_18310);
nor U24949 (N_24949,N_19935,N_18686);
nand U24950 (N_24950,N_17606,N_15056);
or U24951 (N_24951,N_18290,N_16925);
or U24952 (N_24952,N_17429,N_16883);
or U24953 (N_24953,N_19912,N_16522);
or U24954 (N_24954,N_17710,N_18640);
nand U24955 (N_24955,N_17218,N_19465);
nand U24956 (N_24956,N_19332,N_18026);
or U24957 (N_24957,N_19241,N_15273);
and U24958 (N_24958,N_18171,N_16545);
nor U24959 (N_24959,N_15828,N_15198);
nand U24960 (N_24960,N_15874,N_15426);
nor U24961 (N_24961,N_16041,N_19424);
nand U24962 (N_24962,N_15785,N_19450);
xnor U24963 (N_24963,N_15573,N_15043);
xor U24964 (N_24964,N_16500,N_15988);
or U24965 (N_24965,N_17836,N_19464);
xor U24966 (N_24966,N_18322,N_16723);
nand U24967 (N_24967,N_16174,N_17916);
and U24968 (N_24968,N_17977,N_16809);
nor U24969 (N_24969,N_16932,N_16638);
and U24970 (N_24970,N_17402,N_19773);
nand U24971 (N_24971,N_17800,N_19877);
or U24972 (N_24972,N_19697,N_16936);
and U24973 (N_24973,N_15960,N_17965);
nor U24974 (N_24974,N_15310,N_19800);
nand U24975 (N_24975,N_16347,N_18336);
xor U24976 (N_24976,N_16702,N_18244);
or U24977 (N_24977,N_19994,N_19193);
xor U24978 (N_24978,N_16057,N_19534);
or U24979 (N_24979,N_16584,N_18598);
xor U24980 (N_24980,N_19063,N_16935);
or U24981 (N_24981,N_19780,N_16490);
nor U24982 (N_24982,N_17799,N_17090);
nand U24983 (N_24983,N_19917,N_16064);
or U24984 (N_24984,N_18935,N_18145);
nand U24985 (N_24985,N_16291,N_16846);
nor U24986 (N_24986,N_17039,N_17061);
nand U24987 (N_24987,N_19601,N_17115);
and U24988 (N_24988,N_17780,N_17747);
xnor U24989 (N_24989,N_17622,N_19670);
nand U24990 (N_24990,N_16931,N_16021);
xor U24991 (N_24991,N_19749,N_17773);
xor U24992 (N_24992,N_15631,N_17969);
nand U24993 (N_24993,N_18767,N_17582);
nor U24994 (N_24994,N_19995,N_16416);
nand U24995 (N_24995,N_16185,N_15150);
xnor U24996 (N_24996,N_16296,N_16318);
and U24997 (N_24997,N_15610,N_18420);
xor U24998 (N_24998,N_15983,N_19633);
and U24999 (N_24999,N_16544,N_16350);
xnor U25000 (N_25000,N_24789,N_24838);
nor U25001 (N_25001,N_23209,N_20652);
xnor U25002 (N_25002,N_24772,N_22088);
nor U25003 (N_25003,N_24954,N_22734);
xnor U25004 (N_25004,N_20733,N_20262);
xor U25005 (N_25005,N_23668,N_23432);
and U25006 (N_25006,N_22202,N_20893);
and U25007 (N_25007,N_22038,N_23624);
xor U25008 (N_25008,N_22546,N_22595);
xnor U25009 (N_25009,N_24230,N_23660);
xnor U25010 (N_25010,N_22651,N_22116);
or U25011 (N_25011,N_24958,N_23367);
nor U25012 (N_25012,N_23980,N_21392);
nor U25013 (N_25013,N_21642,N_23419);
and U25014 (N_25014,N_20832,N_20810);
and U25015 (N_25015,N_20324,N_23318);
and U25016 (N_25016,N_22872,N_22795);
and U25017 (N_25017,N_23160,N_23170);
nand U25018 (N_25018,N_24743,N_22007);
or U25019 (N_25019,N_20213,N_20927);
nand U25020 (N_25020,N_21566,N_20798);
or U25021 (N_25021,N_22364,N_22189);
nand U25022 (N_25022,N_23255,N_23607);
or U25023 (N_25023,N_22978,N_20092);
or U25024 (N_25024,N_24690,N_24455);
and U25025 (N_25025,N_21699,N_21575);
nand U25026 (N_25026,N_24172,N_20591);
nand U25027 (N_25027,N_20860,N_24408);
nand U25028 (N_25028,N_21875,N_21924);
and U25029 (N_25029,N_20844,N_23133);
or U25030 (N_25030,N_24422,N_23125);
nand U25031 (N_25031,N_23233,N_20751);
nor U25032 (N_25032,N_21960,N_21078);
nor U25033 (N_25033,N_21915,N_23741);
xnor U25034 (N_25034,N_21718,N_24996);
nand U25035 (N_25035,N_21743,N_22145);
xnor U25036 (N_25036,N_23132,N_22353);
nor U25037 (N_25037,N_24178,N_21028);
xnor U25038 (N_25038,N_21665,N_20684);
xor U25039 (N_25039,N_24615,N_24662);
and U25040 (N_25040,N_24607,N_21299);
or U25041 (N_25041,N_23226,N_24805);
and U25042 (N_25042,N_23806,N_23535);
and U25043 (N_25043,N_23533,N_22976);
or U25044 (N_25044,N_22752,N_24327);
or U25045 (N_25045,N_23413,N_20510);
or U25046 (N_25046,N_23162,N_22446);
and U25047 (N_25047,N_22569,N_24765);
nand U25048 (N_25048,N_23642,N_24707);
and U25049 (N_25049,N_21022,N_22264);
or U25050 (N_25050,N_22031,N_24558);
nor U25051 (N_25051,N_21463,N_24596);
nand U25052 (N_25052,N_21710,N_20540);
and U25053 (N_25053,N_21644,N_20706);
nor U25054 (N_25054,N_20284,N_22747);
and U25055 (N_25055,N_20434,N_21577);
nor U25056 (N_25056,N_22653,N_22470);
xnor U25057 (N_25057,N_24913,N_21668);
and U25058 (N_25058,N_21616,N_22713);
nor U25059 (N_25059,N_21885,N_20767);
or U25060 (N_25060,N_24559,N_24293);
or U25061 (N_25061,N_22055,N_24288);
or U25062 (N_25062,N_24198,N_21376);
or U25063 (N_25063,N_24302,N_20368);
nor U25064 (N_25064,N_23789,N_21432);
nor U25065 (N_25065,N_22300,N_21223);
xor U25066 (N_25066,N_20531,N_20218);
nand U25067 (N_25067,N_20567,N_22125);
and U25068 (N_25068,N_20141,N_20574);
nand U25069 (N_25069,N_20665,N_22187);
xnor U25070 (N_25070,N_20010,N_22053);
nor U25071 (N_25071,N_21721,N_24622);
and U25072 (N_25072,N_24507,N_20594);
xnor U25073 (N_25073,N_24991,N_21860);
nand U25074 (N_25074,N_21099,N_20985);
or U25075 (N_25075,N_21568,N_24001);
or U25076 (N_25076,N_21424,N_22958);
nand U25077 (N_25077,N_20124,N_24099);
nand U25078 (N_25078,N_21091,N_20310);
or U25079 (N_25079,N_21853,N_20187);
or U25080 (N_25080,N_21878,N_21595);
or U25081 (N_25081,N_20926,N_24637);
xor U25082 (N_25082,N_20941,N_22244);
or U25083 (N_25083,N_24541,N_21464);
xnor U25084 (N_25084,N_22537,N_20912);
and U25085 (N_25085,N_20204,N_24435);
and U25086 (N_25086,N_21119,N_24668);
nand U25087 (N_25087,N_21156,N_24747);
and U25088 (N_25088,N_22208,N_21285);
nor U25089 (N_25089,N_24856,N_23877);
and U25090 (N_25090,N_22424,N_21708);
nand U25091 (N_25091,N_20461,N_21007);
xor U25092 (N_25092,N_21850,N_21371);
and U25093 (N_25093,N_22362,N_20309);
nor U25094 (N_25094,N_21811,N_22521);
nor U25095 (N_25095,N_23247,N_22603);
xnor U25096 (N_25096,N_21630,N_24732);
nor U25097 (N_25097,N_22731,N_24013);
nor U25098 (N_25098,N_22641,N_21732);
nor U25099 (N_25099,N_20068,N_21106);
nand U25100 (N_25100,N_24487,N_24342);
or U25101 (N_25101,N_23224,N_23951);
nand U25102 (N_25102,N_24227,N_24933);
nor U25103 (N_25103,N_23622,N_24813);
nor U25104 (N_25104,N_24167,N_23055);
and U25105 (N_25105,N_21331,N_20744);
nor U25106 (N_25106,N_24359,N_23331);
or U25107 (N_25107,N_22634,N_22871);
or U25108 (N_25108,N_24523,N_21416);
xor U25109 (N_25109,N_24326,N_22623);
or U25110 (N_25110,N_24225,N_20077);
xor U25111 (N_25111,N_24527,N_24494);
nor U25112 (N_25112,N_22413,N_23589);
xor U25113 (N_25113,N_21641,N_24266);
nand U25114 (N_25114,N_22729,N_22379);
xor U25115 (N_25115,N_22231,N_21681);
xor U25116 (N_25116,N_20763,N_22988);
nor U25117 (N_25117,N_23199,N_22862);
or U25118 (N_25118,N_24875,N_20532);
nor U25119 (N_25119,N_22178,N_21385);
or U25120 (N_25120,N_24185,N_24074);
or U25121 (N_25121,N_23684,N_23575);
nor U25122 (N_25122,N_21417,N_22704);
or U25123 (N_25123,N_24040,N_23458);
or U25124 (N_25124,N_24534,N_21974);
or U25125 (N_25125,N_22482,N_21459);
nor U25126 (N_25126,N_23137,N_24750);
and U25127 (N_25127,N_21343,N_21956);
nor U25128 (N_25128,N_22343,N_23395);
xnor U25129 (N_25129,N_23682,N_22531);
or U25130 (N_25130,N_22973,N_20137);
or U25131 (N_25131,N_21033,N_23591);
and U25132 (N_25132,N_21415,N_24821);
nor U25133 (N_25133,N_23493,N_20935);
and U25134 (N_25134,N_20797,N_23386);
or U25135 (N_25135,N_22776,N_21330);
and U25136 (N_25136,N_20624,N_24539);
nor U25137 (N_25137,N_20539,N_24588);
or U25138 (N_25138,N_20669,N_21023);
xor U25139 (N_25139,N_23011,N_24704);
nand U25140 (N_25140,N_20930,N_20739);
nand U25141 (N_25141,N_20096,N_21748);
xor U25142 (N_25142,N_22811,N_20477);
and U25143 (N_25143,N_21719,N_23586);
nand U25144 (N_25144,N_22585,N_20219);
and U25145 (N_25145,N_20307,N_23345);
nand U25146 (N_25146,N_24763,N_24022);
xnor U25147 (N_25147,N_23737,N_20827);
and U25148 (N_25148,N_22333,N_21972);
xor U25149 (N_25149,N_20809,N_24692);
or U25150 (N_25150,N_20709,N_22104);
xor U25151 (N_25151,N_22403,N_21025);
xor U25152 (N_25152,N_21554,N_22027);
nand U25153 (N_25153,N_22491,N_22937);
or U25154 (N_25154,N_23050,N_20864);
and U25155 (N_25155,N_20344,N_20297);
nand U25156 (N_25156,N_23587,N_21802);
xor U25157 (N_25157,N_23144,N_23521);
or U25158 (N_25158,N_22861,N_23488);
and U25159 (N_25159,N_24702,N_20119);
nand U25160 (N_25160,N_20238,N_20753);
nor U25161 (N_25161,N_24224,N_23970);
xnor U25162 (N_25162,N_24170,N_20590);
xor U25163 (N_25163,N_22063,N_20558);
xor U25164 (N_25164,N_23551,N_21574);
nor U25165 (N_25165,N_22069,N_21856);
nor U25166 (N_25166,N_22559,N_24570);
or U25167 (N_25167,N_23519,N_24263);
nor U25168 (N_25168,N_24300,N_21095);
or U25169 (N_25169,N_21934,N_20794);
nand U25170 (N_25170,N_24749,N_23724);
xor U25171 (N_25171,N_20325,N_23735);
nand U25172 (N_25172,N_22121,N_24072);
and U25173 (N_25173,N_23028,N_22890);
or U25174 (N_25174,N_20750,N_22925);
and U25175 (N_25175,N_21987,N_20494);
and U25176 (N_25176,N_23008,N_22657);
and U25177 (N_25177,N_24552,N_22236);
and U25178 (N_25178,N_24337,N_24365);
and U25179 (N_25179,N_21379,N_22373);
nor U25180 (N_25180,N_21035,N_21100);
xnor U25181 (N_25181,N_22549,N_20755);
nor U25182 (N_25182,N_24656,N_22083);
nand U25183 (N_25183,N_21485,N_20824);
xnor U25184 (N_25184,N_20456,N_20823);
or U25185 (N_25185,N_22773,N_20403);
nand U25186 (N_25186,N_21410,N_22701);
nor U25187 (N_25187,N_20318,N_24754);
and U25188 (N_25188,N_23250,N_20331);
or U25189 (N_25189,N_24751,N_24258);
xnor U25190 (N_25190,N_21542,N_22294);
xnor U25191 (N_25191,N_23872,N_24524);
and U25192 (N_25192,N_21158,N_20192);
and U25193 (N_25193,N_23308,N_24132);
and U25194 (N_25194,N_24910,N_20828);
nand U25195 (N_25195,N_24606,N_22129);
nand U25196 (N_25196,N_20479,N_20766);
nand U25197 (N_25197,N_22859,N_23664);
xnor U25198 (N_25198,N_22676,N_22520);
and U25199 (N_25199,N_20633,N_20547);
xor U25200 (N_25200,N_24629,N_21067);
nand U25201 (N_25201,N_22440,N_24936);
or U25202 (N_25202,N_21524,N_20321);
nand U25203 (N_25203,N_21239,N_24706);
nand U25204 (N_25204,N_23698,N_20134);
and U25205 (N_25205,N_22371,N_22351);
nand U25206 (N_25206,N_20375,N_20432);
nand U25207 (N_25207,N_22665,N_23447);
or U25208 (N_25208,N_22140,N_21923);
or U25209 (N_25209,N_22020,N_20193);
xnor U25210 (N_25210,N_24923,N_20332);
or U25211 (N_25211,N_21725,N_21831);
xor U25212 (N_25212,N_21112,N_20880);
and U25213 (N_25213,N_20518,N_21182);
or U25214 (N_25214,N_23176,N_22718);
or U25215 (N_25215,N_23729,N_20620);
xnor U25216 (N_25216,N_21240,N_24551);
and U25217 (N_25217,N_20184,N_23289);
nand U25218 (N_25218,N_24713,N_21320);
nor U25219 (N_25219,N_21457,N_24906);
or U25220 (N_25220,N_22605,N_20074);
nor U25221 (N_25221,N_24452,N_24195);
nor U25222 (N_25222,N_21068,N_21953);
xor U25223 (N_25223,N_23925,N_20209);
xnor U25224 (N_25224,N_21889,N_23359);
nor U25225 (N_25225,N_21527,N_20362);
nor U25226 (N_25226,N_23175,N_23457);
nand U25227 (N_25227,N_23037,N_23356);
nand U25228 (N_25228,N_20572,N_22152);
nand U25229 (N_25229,N_23506,N_22332);
or U25230 (N_25230,N_21984,N_24222);
nor U25231 (N_25231,N_24152,N_20255);
nand U25232 (N_25232,N_24136,N_23649);
nor U25233 (N_25233,N_22600,N_23006);
or U25234 (N_25234,N_21456,N_22432);
xnor U25235 (N_25235,N_20361,N_23513);
or U25236 (N_25236,N_22015,N_24748);
nor U25237 (N_25237,N_23016,N_23914);
or U25238 (N_25238,N_20185,N_23051);
or U25239 (N_25239,N_23117,N_23888);
xor U25240 (N_25240,N_23992,N_23164);
nor U25241 (N_25241,N_24476,N_24594);
nand U25242 (N_25242,N_24491,N_23296);
and U25243 (N_25243,N_22064,N_22052);
and U25244 (N_25244,N_22710,N_23382);
or U25245 (N_25245,N_23225,N_23288);
or U25246 (N_25246,N_21526,N_22474);
xor U25247 (N_25247,N_22295,N_24636);
nand U25248 (N_25248,N_23675,N_24879);
xnor U25249 (N_25249,N_23343,N_20014);
or U25250 (N_25250,N_20686,N_24961);
or U25251 (N_25251,N_21496,N_21059);
and U25252 (N_25252,N_20708,N_21209);
or U25253 (N_25253,N_20478,N_23929);
xnor U25254 (N_25254,N_21017,N_24047);
xor U25255 (N_25255,N_24686,N_22261);
nor U25256 (N_25256,N_23665,N_20889);
nand U25257 (N_25257,N_21613,N_20314);
nor U25258 (N_25258,N_23362,N_23695);
nor U25259 (N_25259,N_23630,N_24111);
or U25260 (N_25260,N_22891,N_24724);
nor U25261 (N_25261,N_23921,N_21216);
or U25262 (N_25262,N_20037,N_21973);
and U25263 (N_25263,N_20174,N_22283);
xor U25264 (N_25264,N_23310,N_20543);
or U25265 (N_25265,N_23287,N_22277);
or U25266 (N_25266,N_23715,N_21083);
nand U25267 (N_25267,N_20167,N_21257);
and U25268 (N_25268,N_21760,N_23704);
nor U25269 (N_25269,N_21269,N_24519);
and U25270 (N_25270,N_20370,N_21263);
nand U25271 (N_25271,N_20714,N_23400);
nand U25272 (N_25272,N_23663,N_21374);
nand U25273 (N_25273,N_24361,N_22561);
nand U25274 (N_25274,N_20639,N_24148);
and U25275 (N_25275,N_23516,N_23959);
and U25276 (N_25276,N_20021,N_20994);
nor U25277 (N_25277,N_20987,N_20969);
nor U25278 (N_25278,N_21277,N_22366);
or U25279 (N_25279,N_22589,N_23791);
or U25280 (N_25280,N_21809,N_21152);
xor U25281 (N_25281,N_21872,N_23376);
nor U25282 (N_25282,N_21996,N_24912);
or U25283 (N_25283,N_21758,N_24522);
nor U25284 (N_25284,N_21785,N_20788);
xnor U25285 (N_25285,N_20483,N_20413);
nand U25286 (N_25286,N_22649,N_22992);
nand U25287 (N_25287,N_20151,N_22568);
nor U25288 (N_25288,N_24947,N_21284);
nand U25289 (N_25289,N_20188,N_24011);
or U25290 (N_25290,N_20071,N_22968);
nor U25291 (N_25291,N_24461,N_22313);
xor U25292 (N_25292,N_24209,N_21387);
xnor U25293 (N_25293,N_22417,N_22349);
and U25294 (N_25294,N_23350,N_22550);
nor U25295 (N_25295,N_21283,N_20570);
nand U25296 (N_25296,N_24118,N_22818);
nor U25297 (N_25297,N_20923,N_24532);
nor U25298 (N_25298,N_22508,N_20427);
xor U25299 (N_25299,N_24902,N_24369);
nor U25300 (N_25300,N_22042,N_23804);
nor U25301 (N_25301,N_24071,N_24920);
nor U25302 (N_25302,N_21509,N_20537);
or U25303 (N_25303,N_23564,N_21731);
and U25304 (N_25304,N_20300,N_22370);
and U25305 (N_25305,N_21946,N_22009);
and U25306 (N_25306,N_20208,N_20854);
xnor U25307 (N_25307,N_20101,N_24329);
or U25308 (N_25308,N_20953,N_24357);
or U25309 (N_25309,N_21130,N_22211);
xor U25310 (N_25310,N_24826,N_20589);
nor U25311 (N_25311,N_22922,N_24889);
nor U25312 (N_25312,N_22184,N_22302);
nand U25313 (N_25313,N_24809,N_20934);
or U25314 (N_25314,N_22831,N_20961);
nand U25315 (N_25315,N_21167,N_20853);
xnor U25316 (N_25316,N_23555,N_22165);
and U25317 (N_25317,N_23773,N_23627);
nand U25318 (N_25318,N_20999,N_21206);
and U25319 (N_25319,N_23416,N_20785);
or U25320 (N_25320,N_22914,N_22771);
nor U25321 (N_25321,N_22213,N_20446);
and U25322 (N_25322,N_22892,N_23887);
and U25323 (N_25323,N_23529,N_21949);
xnor U25324 (N_25324,N_20177,N_22324);
xor U25325 (N_25325,N_22280,N_23088);
xnor U25326 (N_25326,N_20038,N_20507);
or U25327 (N_25327,N_24579,N_24284);
xor U25328 (N_25328,N_20536,N_24599);
xor U25329 (N_25329,N_21689,N_20227);
nand U25330 (N_25330,N_23934,N_23029);
xor U25331 (N_25331,N_21833,N_24456);
nor U25332 (N_25332,N_24256,N_22374);
or U25333 (N_25333,N_21783,N_24874);
xor U25334 (N_25334,N_21069,N_20269);
and U25335 (N_25335,N_21533,N_20648);
or U25336 (N_25336,N_23845,N_23600);
nor U25337 (N_25337,N_23123,N_22753);
xnor U25338 (N_25338,N_20509,N_24700);
or U25339 (N_25339,N_23520,N_22849);
nor U25340 (N_25340,N_23638,N_20067);
xor U25341 (N_25341,N_23818,N_23942);
and U25342 (N_25342,N_23907,N_24401);
xnor U25343 (N_25343,N_21607,N_20777);
or U25344 (N_25344,N_22781,N_21518);
and U25345 (N_25345,N_20260,N_20399);
and U25346 (N_25346,N_24130,N_24712);
nand U25347 (N_25347,N_20166,N_22777);
nand U25348 (N_25348,N_22635,N_23053);
xnor U25349 (N_25349,N_22198,N_21608);
nand U25350 (N_25350,N_20940,N_20760);
nor U25351 (N_25351,N_23409,N_21324);
nand U25352 (N_25352,N_20820,N_22409);
and U25353 (N_25353,N_23531,N_20691);
xnor U25354 (N_25354,N_23746,N_21704);
xnor U25355 (N_25355,N_22040,N_21862);
nor U25356 (N_25356,N_20380,N_24870);
and U25357 (N_25357,N_21600,N_23384);
nand U25358 (N_25358,N_21629,N_21292);
xnor U25359 (N_25359,N_23222,N_23354);
nor U25360 (N_25360,N_24760,N_22241);
nand U25361 (N_25361,N_24180,N_23126);
nand U25362 (N_25362,N_24984,N_21846);
nand U25363 (N_25363,N_20384,N_20169);
xor U25364 (N_25364,N_23052,N_23389);
or U25365 (N_25365,N_23219,N_21072);
or U25366 (N_25366,N_24880,N_21369);
or U25367 (N_25367,N_24457,N_22043);
nor U25368 (N_25368,N_22131,N_23726);
nand U25369 (N_25369,N_24176,N_20439);
xnor U25370 (N_25370,N_21406,N_23449);
nand U25371 (N_25371,N_24768,N_22199);
nor U25372 (N_25372,N_23728,N_24308);
nand U25373 (N_25373,N_23817,N_23866);
nand U25374 (N_25374,N_21529,N_21306);
xnor U25375 (N_25375,N_23009,N_23254);
or U25376 (N_25376,N_20386,N_20108);
xnor U25377 (N_25377,N_22076,N_21650);
xor U25378 (N_25378,N_23885,N_23709);
nor U25379 (N_25379,N_22656,N_23994);
and U25380 (N_25380,N_20700,N_23539);
nand U25381 (N_25381,N_24972,N_23847);
nand U25382 (N_25382,N_23816,N_24469);
nand U25383 (N_25383,N_23931,N_23046);
xnor U25384 (N_25384,N_20057,N_21649);
xnor U25385 (N_25385,N_20093,N_20086);
and U25386 (N_25386,N_21162,N_23079);
and U25387 (N_25387,N_21786,N_24911);
and U25388 (N_25388,N_20140,N_24628);
nor U25389 (N_25389,N_21453,N_23650);
and U25390 (N_25390,N_23451,N_20319);
xor U25391 (N_25391,N_24776,N_23184);
nand U25392 (N_25392,N_24669,N_20482);
xor U25393 (N_25393,N_24449,N_24841);
xor U25394 (N_25394,N_24943,N_22667);
nor U25395 (N_25395,N_24486,N_21370);
xnor U25396 (N_25396,N_20550,N_22099);
xnor U25397 (N_25397,N_21295,N_20266);
or U25398 (N_25398,N_22994,N_22401);
nand U25399 (N_25399,N_23671,N_21550);
or U25400 (N_25400,N_21976,N_20573);
or U25401 (N_25401,N_22355,N_23238);
nor U25402 (N_25402,N_22462,N_24715);
nor U25403 (N_25403,N_20636,N_24070);
or U25404 (N_25404,N_20869,N_20454);
or U25405 (N_25405,N_24684,N_22932);
nor U25406 (N_25406,N_22532,N_22756);
or U25407 (N_25407,N_24362,N_22322);
nor U25408 (N_25408,N_24246,N_23800);
and U25409 (N_25409,N_20522,N_23111);
xnor U25410 (N_25410,N_23680,N_24535);
nand U25411 (N_25411,N_24305,N_20673);
and U25412 (N_25412,N_23582,N_23163);
and U25413 (N_25413,N_22611,N_20155);
or U25414 (N_25414,N_22722,N_22115);
and U25415 (N_25415,N_24414,N_24793);
nor U25416 (N_25416,N_20857,N_24458);
or U25417 (N_25417,N_20900,N_20581);
nor U25418 (N_25418,N_21683,N_21298);
nand U25419 (N_25419,N_22186,N_24432);
nor U25420 (N_25420,N_24924,N_20775);
xor U25421 (N_25421,N_23999,N_20908);
nand U25422 (N_25422,N_20058,N_21902);
nand U25423 (N_25423,N_22335,N_21246);
xor U25424 (N_25424,N_23057,N_24285);
and U25425 (N_25425,N_23476,N_22049);
xnor U25426 (N_25426,N_21413,N_20222);
xor U25427 (N_25427,N_23372,N_24053);
nand U25428 (N_25428,N_24613,N_20168);
or U25429 (N_25429,N_22796,N_22738);
nand U25430 (N_25430,N_23854,N_21674);
or U25431 (N_25431,N_20270,N_24926);
or U25432 (N_25432,N_21588,N_20317);
xor U25433 (N_25433,N_20156,N_23018);
nand U25434 (N_25434,N_24682,N_22551);
xor U25435 (N_25435,N_21970,N_21790);
xnor U25436 (N_25436,N_20990,N_22279);
nand U25437 (N_25437,N_21691,N_23687);
or U25438 (N_25438,N_20724,N_24799);
and U25439 (N_25439,N_21241,N_21504);
nand U25440 (N_25440,N_22769,N_23782);
nor U25441 (N_25441,N_21037,N_22037);
nand U25442 (N_25442,N_20963,N_22800);
nand U25443 (N_25443,N_23802,N_24925);
nand U25444 (N_25444,N_20924,N_21816);
nand U25445 (N_25445,N_23577,N_23814);
or U25446 (N_25446,N_20385,N_21155);
nor U25447 (N_25447,N_20967,N_22106);
nor U25448 (N_25448,N_23605,N_23455);
xor U25449 (N_25449,N_20833,N_22381);
and U25450 (N_25450,N_23851,N_20299);
nand U25451 (N_25451,N_23060,N_23392);
nor U25452 (N_25452,N_23754,N_22173);
nand U25453 (N_25453,N_24572,N_24908);
xnor U25454 (N_25454,N_20148,N_21061);
nor U25455 (N_25455,N_22350,N_22347);
nand U25456 (N_25456,N_24392,N_24086);
nor U25457 (N_25457,N_21938,N_20275);
and U25458 (N_25458,N_23511,N_22066);
xnor U25459 (N_25459,N_24935,N_20783);
nor U25460 (N_25460,N_22763,N_23646);
or U25461 (N_25461,N_23611,N_24565);
nor U25462 (N_25462,N_21700,N_23861);
xnor U25463 (N_25463,N_22336,N_22552);
and U25464 (N_25464,N_21391,N_23501);
and U25465 (N_25465,N_24377,N_22312);
nor U25466 (N_25466,N_21151,N_21177);
nand U25467 (N_25467,N_22460,N_24159);
or U25468 (N_25468,N_20022,N_22134);
and U25469 (N_25469,N_23251,N_21418);
nor U25470 (N_25470,N_20667,N_21651);
xnor U25471 (N_25471,N_20273,N_24126);
nand U25472 (N_25472,N_20019,N_22919);
and U25473 (N_25473,N_21579,N_20595);
nor U25474 (N_25474,N_20513,N_22748);
or U25475 (N_25475,N_23813,N_23281);
and U25476 (N_25476,N_20933,N_22238);
or U25477 (N_25477,N_20830,N_20748);
and U25478 (N_25478,N_22148,N_20811);
nor U25479 (N_25479,N_20831,N_20678);
nor U25480 (N_25480,N_24459,N_22144);
and U25481 (N_25481,N_22075,N_22119);
or U25482 (N_25482,N_23047,N_20698);
or U25483 (N_25483,N_23049,N_21407);
nor U25484 (N_25484,N_21086,N_23721);
xnor U25485 (N_25485,N_20729,N_20205);
or U25486 (N_25486,N_23243,N_23138);
nor U25487 (N_25487,N_22804,N_24562);
or U25488 (N_25488,N_23810,N_24407);
or U25489 (N_25489,N_22619,N_24802);
or U25490 (N_25490,N_23227,N_20568);
nand U25491 (N_25491,N_23714,N_22608);
and U25492 (N_25492,N_23307,N_21359);
xnor U25493 (N_25493,N_24144,N_20277);
xor U25494 (N_25494,N_20981,N_20789);
xor U25495 (N_25495,N_22930,N_21250);
and U25496 (N_25496,N_22979,N_21012);
xnor U25497 (N_25497,N_22377,N_22624);
nor U25498 (N_25498,N_22288,N_23974);
xnor U25499 (N_25499,N_20463,N_22857);
xor U25500 (N_25500,N_22382,N_23078);
or U25501 (N_25501,N_20158,N_24405);
nor U25502 (N_25502,N_24472,N_20200);
and U25503 (N_25503,N_21036,N_21058);
nand U25504 (N_25504,N_22645,N_22659);
xor U25505 (N_25505,N_20592,N_20770);
nand U25506 (N_25506,N_21672,N_24358);
and U25507 (N_25507,N_24581,N_22766);
nor U25508 (N_25508,N_22516,N_22496);
or U25509 (N_25509,N_23739,N_22828);
and U25510 (N_25510,N_20910,N_20106);
nand U25511 (N_25511,N_21599,N_21892);
xor U25512 (N_25512,N_22404,N_22041);
nor U25513 (N_25513,N_22450,N_22372);
or U25514 (N_25514,N_23487,N_20048);
nor U25515 (N_25515,N_23177,N_24439);
or U25516 (N_25516,N_20852,N_21925);
xor U25517 (N_25517,N_22586,N_24065);
xor U25518 (N_25518,N_24907,N_20932);
nor U25519 (N_25519,N_20867,N_20538);
nand U25520 (N_25520,N_24142,N_24881);
and U25521 (N_25521,N_22019,N_21047);
nand U25522 (N_25522,N_22029,N_23020);
and U25523 (N_25523,N_24382,N_23759);
or U25524 (N_25524,N_21604,N_21558);
xor U25525 (N_25525,N_21888,N_24229);
or U25526 (N_25526,N_21421,N_22393);
and U25527 (N_25527,N_22926,N_23777);
nand U25528 (N_25528,N_23596,N_21800);
nand U25529 (N_25529,N_23290,N_20598);
nand U25530 (N_25530,N_21032,N_23809);
nor U25531 (N_25531,N_20263,N_23062);
nand U25532 (N_25532,N_21729,N_20217);
nand U25533 (N_25533,N_20017,N_22415);
xnor U25534 (N_25534,N_20224,N_23850);
nand U25535 (N_25535,N_23216,N_20781);
or U25536 (N_25536,N_23071,N_21315);
nand U25537 (N_25537,N_23563,N_21601);
and U25538 (N_25538,N_21278,N_22709);
and U25539 (N_25539,N_23231,N_23532);
and U25540 (N_25540,N_24138,N_23565);
or U25541 (N_25541,N_20425,N_21322);
nor U25542 (N_25542,N_21756,N_21940);
nand U25543 (N_25543,N_23156,N_23000);
and U25544 (N_25544,N_21676,N_21513);
nor U25545 (N_25545,N_20303,N_24974);
xnor U25546 (N_25546,N_22412,N_23379);
nor U25547 (N_25547,N_21360,N_21702);
nand U25548 (N_25548,N_24716,N_23106);
xnor U25549 (N_25549,N_21202,N_21762);
nor U25550 (N_25550,N_24343,N_22606);
nand U25551 (N_25551,N_23140,N_24783);
nor U25552 (N_25552,N_21628,N_22384);
and U25553 (N_25553,N_23368,N_24000);
or U25554 (N_25554,N_24739,N_20008);
xnor U25555 (N_25555,N_22061,N_20239);
and U25556 (N_25556,N_22941,N_24427);
nor U25557 (N_25557,N_21362,N_20841);
nand U25558 (N_25558,N_24624,N_23198);
or U25559 (N_25559,N_20256,N_20497);
xnor U25560 (N_25560,N_20237,N_22354);
nand U25561 (N_25561,N_22523,N_21931);
nor U25562 (N_25562,N_23149,N_22894);
nor U25563 (N_25563,N_21325,N_20704);
nand U25564 (N_25564,N_24497,N_23852);
or U25565 (N_25565,N_20225,N_21553);
xnor U25566 (N_25566,N_23193,N_22576);
and U25567 (N_25567,N_23924,N_24653);
nor U25568 (N_25568,N_24355,N_24064);
xor U25569 (N_25569,N_20129,N_20353);
nor U25570 (N_25570,N_24280,N_21521);
and U25571 (N_25571,N_20272,N_20215);
xnor U25572 (N_25572,N_24542,N_22823);
or U25573 (N_25573,N_21750,N_22500);
and U25574 (N_25574,N_21943,N_24390);
nor U25575 (N_25575,N_24137,N_22271);
and U25576 (N_25576,N_20960,N_22755);
or U25577 (N_25577,N_22971,N_22014);
and U25578 (N_25578,N_24325,N_23430);
and U25579 (N_25579,N_23573,N_24987);
xor U25580 (N_25580,N_20954,N_22933);
or U25581 (N_25581,N_20085,N_21001);
or U25582 (N_25582,N_23097,N_22842);
nand U25583 (N_25583,N_24829,N_22151);
nor U25584 (N_25584,N_23127,N_24547);
nand U25585 (N_25585,N_23755,N_23538);
and U25586 (N_25586,N_23636,N_24190);
or U25587 (N_25587,N_24061,N_22180);
or U25588 (N_25588,N_20442,N_20396);
and U25589 (N_25589,N_21687,N_21488);
and U25590 (N_25590,N_23230,N_22130);
or U25591 (N_25591,N_23958,N_24526);
xor U25592 (N_25592,N_22885,N_23223);
xnor U25593 (N_25593,N_21481,N_23964);
nor U25594 (N_25594,N_24386,N_22065);
xnor U25595 (N_25595,N_24129,N_21029);
xor U25596 (N_25596,N_24066,N_21639);
xnor U25597 (N_25597,N_24944,N_24845);
and U25598 (N_25598,N_23168,N_24866);
and U25599 (N_25599,N_21469,N_21571);
and U25600 (N_25600,N_24171,N_22387);
nor U25601 (N_25601,N_24353,N_22345);
and U25602 (N_25602,N_22519,N_23678);
and U25603 (N_25603,N_23207,N_21104);
and U25604 (N_25604,N_22176,N_20993);
and U25605 (N_25605,N_22367,N_20703);
xnor U25606 (N_25606,N_22509,N_22445);
nand U25607 (N_25607,N_21336,N_20627);
xnor U25608 (N_25608,N_23902,N_23574);
nor U25609 (N_25609,N_22607,N_22984);
nor U25610 (N_25610,N_21235,N_20812);
or U25611 (N_25611,N_20046,N_21252);
or U25612 (N_25612,N_20814,N_24504);
xnor U25613 (N_25613,N_21873,N_20944);
and U25614 (N_25614,N_24647,N_20171);
nand U25615 (N_25615,N_21039,N_23489);
and U25616 (N_25616,N_23328,N_22887);
xnor U25617 (N_25617,N_21296,N_23774);
and U25618 (N_25618,N_21722,N_23525);
xnor U25619 (N_25619,N_22207,N_21181);
nand U25620 (N_25620,N_23920,N_24888);
or U25621 (N_25621,N_23656,N_24740);
or U25622 (N_25622,N_21986,N_24234);
nor U25623 (N_25623,N_23712,N_23034);
nor U25624 (N_25624,N_20800,N_23553);
nand U25625 (N_25625,N_24804,N_21844);
and U25626 (N_25626,N_22451,N_23129);
and U25627 (N_25627,N_24801,N_23450);
and U25628 (N_25628,N_21627,N_20444);
xor U25629 (N_25629,N_21855,N_22082);
xnor U25630 (N_25630,N_24521,N_21470);
nand U25631 (N_25631,N_20347,N_22463);
nor U25632 (N_25632,N_21008,N_20615);
nor U25633 (N_25633,N_23437,N_22461);
or U25634 (N_25634,N_24292,N_21774);
xor U25635 (N_25635,N_22917,N_22720);
or U25636 (N_25636,N_24757,N_24951);
or U25637 (N_25637,N_24965,N_21120);
nor U25638 (N_25638,N_22929,N_20525);
nand U25639 (N_25639,N_21903,N_22961);
and U25640 (N_25640,N_21652,N_21137);
or U25641 (N_25641,N_22730,N_23841);
nand U25642 (N_25642,N_21540,N_24151);
nor U25643 (N_25643,N_20040,N_23913);
xnor U25644 (N_25644,N_23056,N_24216);
or U25645 (N_25645,N_23570,N_22767);
xor U25646 (N_25646,N_24871,N_24693);
or U25647 (N_25647,N_22120,N_23448);
nor U25648 (N_25648,N_22678,N_23135);
or U25649 (N_25649,N_24788,N_21757);
or U25650 (N_25650,N_24025,N_23423);
and U25651 (N_25651,N_21980,N_22039);
or U25652 (N_25652,N_21434,N_24106);
xnor U25653 (N_25653,N_23794,N_21005);
xor U25654 (N_25654,N_24169,N_23172);
xor U25655 (N_25655,N_23085,N_23840);
or U25656 (N_25656,N_22931,N_20453);
or U25657 (N_25657,N_24055,N_24276);
and U25658 (N_25658,N_23004,N_21992);
nor U25659 (N_25659,N_22188,N_23462);
nand U25660 (N_25660,N_24219,N_23102);
and U25661 (N_25661,N_20290,N_24398);
xnor U25662 (N_25662,N_21381,N_20561);
and U25663 (N_25663,N_20161,N_24725);
xnor U25664 (N_25664,N_20631,N_21898);
xor U25665 (N_25665,N_20498,N_21189);
and U25666 (N_25666,N_23543,N_20027);
xnor U25667 (N_25667,N_20874,N_21989);
nor U25668 (N_25668,N_21803,N_24135);
nor U25669 (N_25669,N_21132,N_22221);
nor U25670 (N_25670,N_24017,N_22169);
nor U25671 (N_25671,N_22291,N_22564);
xnor U25672 (N_25672,N_22457,N_20500);
or U25673 (N_25673,N_22483,N_21289);
nor U25674 (N_25674,N_23979,N_23859);
xnor U25675 (N_25675,N_23486,N_20146);
or U25676 (N_25676,N_23291,N_22127);
and U25677 (N_25677,N_20136,N_22963);
xor U25678 (N_25678,N_23195,N_21013);
and U25679 (N_25679,N_21562,N_22494);
and U25680 (N_25680,N_20304,N_21784);
or U25681 (N_25681,N_22966,N_22661);
nand U25682 (N_25682,N_20855,N_24164);
xor U25683 (N_25683,N_24566,N_22124);
xor U25684 (N_25684,N_20773,N_21231);
nand U25685 (N_25685,N_23435,N_21670);
nor U25686 (N_25686,N_22594,N_23373);
and U25687 (N_25687,N_20327,N_20523);
nor U25688 (N_25688,N_20122,N_22694);
or U25689 (N_25689,N_23158,N_20529);
and U25690 (N_25690,N_20051,N_20352);
nor U25691 (N_25691,N_22690,N_24567);
nor U25692 (N_25692,N_23470,N_23526);
or U25693 (N_25693,N_22263,N_23558);
xor U25694 (N_25694,N_24182,N_20306);
nor U25695 (N_25695,N_24298,N_22819);
nand U25696 (N_25696,N_21999,N_21864);
or U25697 (N_25697,N_23641,N_21019);
or U25698 (N_25698,N_20836,N_24548);
or U25699 (N_25699,N_22727,N_24425);
and U25700 (N_25700,N_20374,N_23686);
xor U25701 (N_25701,N_23713,N_23962);
xor U25702 (N_25702,N_20196,N_22398);
or U25703 (N_25703,N_24484,N_22171);
xnor U25704 (N_25704,N_24673,N_21895);
and U25705 (N_25705,N_22995,N_22250);
nand U25706 (N_25706,N_23484,N_22081);
or U25707 (N_25707,N_22878,N_24654);
nand U25708 (N_25708,N_20877,N_22522);
and U25709 (N_25709,N_23048,N_23768);
xnor U25710 (N_25710,N_21918,N_24413);
nor U25711 (N_25711,N_24921,N_24928);
xor U25712 (N_25712,N_20722,N_24966);
nor U25713 (N_25713,N_24379,N_20486);
and U25714 (N_25714,N_20131,N_22816);
and U25715 (N_25715,N_24971,N_20717);
and U25716 (N_25716,N_23893,N_22376);
nor U25717 (N_25717,N_21210,N_20407);
nor U25718 (N_25718,N_21088,N_21921);
nor U25719 (N_25719,N_20394,N_22067);
nand U25720 (N_25720,N_22588,N_23072);
nor U25721 (N_25721,N_24741,N_21466);
xor U25722 (N_25722,N_23229,N_24603);
nand U25723 (N_25723,N_23894,N_20162);
xnor U25724 (N_25724,N_21749,N_21807);
xnor U25725 (N_25725,N_22197,N_24247);
xor U25726 (N_25726,N_21911,N_22790);
nand U25727 (N_25727,N_24341,N_20041);
nand U25728 (N_25728,N_24232,N_22426);
and U25729 (N_25729,N_22962,N_21436);
nand U25730 (N_25730,N_21602,N_23261);
nor U25731 (N_25731,N_22737,N_24363);
nand U25732 (N_25732,N_22242,N_20268);
xor U25733 (N_25733,N_24454,N_23613);
xor U25734 (N_25734,N_22468,N_23655);
xnor U25735 (N_25735,N_24964,N_21338);
or U25736 (N_25736,N_23270,N_24490);
or U25737 (N_25737,N_22839,N_22385);
xor U25738 (N_25738,N_24080,N_21841);
nor U25739 (N_25739,N_23321,N_24671);
and U25740 (N_25740,N_22573,N_21706);
or U25741 (N_25741,N_21922,N_24015);
nand U25742 (N_25742,N_24119,N_24346);
or U25743 (N_25743,N_22400,N_20655);
nand U25744 (N_25744,N_24956,N_23131);
or U25745 (N_25745,N_23428,N_23044);
nor U25746 (N_25746,N_22109,N_21408);
and U25747 (N_25747,N_21446,N_21810);
nand U25748 (N_25748,N_24316,N_22910);
and U25749 (N_25749,N_24608,N_21994);
nor U25750 (N_25750,N_22581,N_22498);
nor U25751 (N_25751,N_22967,N_24988);
or U25752 (N_25752,N_24166,N_20416);
nand U25753 (N_25753,N_21146,N_20971);
nand U25754 (N_25754,N_24571,N_24104);
or U25755 (N_25755,N_23453,N_20719);
xor U25756 (N_25756,N_21060,N_22692);
nand U25757 (N_25757,N_24173,N_24212);
and U25758 (N_25758,N_21764,N_24146);
and U25759 (N_25759,N_20947,N_21765);
xnor U25760 (N_25760,N_23976,N_21484);
or U25761 (N_25761,N_20868,N_24893);
xnor U25762 (N_25762,N_22091,N_22072);
nor U25763 (N_25763,N_20422,N_24955);
nand U25764 (N_25764,N_24249,N_22396);
xnor U25765 (N_25765,N_24674,N_22822);
and U25766 (N_25766,N_23349,N_24932);
xor U25767 (N_25767,N_20772,N_23159);
xnor U25768 (N_25768,N_21928,N_24568);
xor U25769 (N_25769,N_24085,N_22691);
and U25770 (N_25770,N_21305,N_22179);
nand U25771 (N_25771,N_21349,N_23842);
xor U25772 (N_25772,N_21661,N_20551);
and U25773 (N_25773,N_23900,N_23228);
and U25774 (N_25774,N_22633,N_23411);
or U25775 (N_25775,N_23477,N_22759);
nand U25776 (N_25776,N_20142,N_21593);
nand U25777 (N_25777,N_20323,N_20713);
or U25778 (N_25778,N_24313,N_22638);
nor U25779 (N_25779,N_22539,N_24197);
xnor U25780 (N_25780,N_20252,N_20579);
nand U25781 (N_25781,N_23892,N_24717);
xnor U25782 (N_25782,N_24975,N_20178);
or U25783 (N_25783,N_21244,N_23927);
and U25784 (N_25784,N_21180,N_22945);
or U25785 (N_25785,N_22380,N_23186);
xor U25786 (N_25786,N_22765,N_20127);
or U25787 (N_25787,N_24718,N_24742);
nor U25788 (N_25788,N_21249,N_21842);
and U25789 (N_25789,N_24934,N_22870);
and U25790 (N_25790,N_24204,N_20281);
xnor U25791 (N_25791,N_23143,N_21804);
nor U25792 (N_25792,N_22684,N_22196);
nand U25793 (N_25793,N_21133,N_22920);
nand U25794 (N_25794,N_22565,N_23708);
xnor U25795 (N_25795,N_21747,N_21632);
and U25796 (N_25796,N_20465,N_24440);
xor U25797 (N_25797,N_24060,N_23292);
or U25798 (N_25798,N_22383,N_20147);
nor U25799 (N_25799,N_21555,N_20493);
nor U25800 (N_25800,N_24556,N_23621);
or U25801 (N_25801,N_21995,N_20411);
nand U25802 (N_25802,N_22079,N_20805);
and U25803 (N_25803,N_23662,N_23946);
nand U25804 (N_25804,N_22886,N_21546);
nor U25805 (N_25805,N_22618,N_23807);
and U25806 (N_25806,N_23042,N_21955);
xnor U25807 (N_25807,N_23275,N_20433);
nor U25808 (N_25808,N_21623,N_24530);
and U25809 (N_25809,N_23578,N_23510);
nor U25810 (N_25810,N_21611,N_20081);
xnor U25811 (N_25811,N_22840,N_24638);
xnor U25812 (N_25812,N_23014,N_23977);
or U25813 (N_25813,N_23808,N_23949);
nor U25814 (N_25814,N_23337,N_21919);
and U25815 (N_25815,N_21212,N_20888);
and U25816 (N_25816,N_22927,N_21397);
nor U25817 (N_25817,N_22918,N_24005);
nand U25818 (N_25818,N_21082,N_22215);
or U25819 (N_25819,N_20555,N_23454);
xnor U25820 (N_25820,N_20992,N_23185);
and U25821 (N_25821,N_21716,N_22143);
nor U25822 (N_25822,N_20641,N_24589);
xnor U25823 (N_25823,N_21089,N_22344);
nor U25824 (N_25824,N_20965,N_20449);
xnor U25825 (N_25825,N_22563,N_22098);
xnor U25826 (N_25826,N_20391,N_20907);
or U25827 (N_25827,N_24217,N_22936);
nand U25828 (N_25828,N_22814,N_23471);
nor U25829 (N_25829,N_22725,N_21002);
nor U25830 (N_25830,N_24777,N_21070);
xor U25831 (N_25831,N_24993,N_21794);
nand U25832 (N_25832,N_24982,N_24762);
nor U25833 (N_25833,N_22274,N_20769);
or U25834 (N_25834,N_22275,N_24174);
or U25835 (N_25835,N_23357,N_22592);
and U25836 (N_25836,N_21113,N_22884);
nand U25837 (N_25837,N_24564,N_21969);
nor U25838 (N_25838,N_22627,N_24372);
or U25839 (N_25839,N_22749,N_21711);
xnor U25840 (N_25840,N_21016,N_21771);
or U25841 (N_25841,N_22325,N_20768);
nand U25842 (N_25842,N_23166,N_24184);
and U25843 (N_25843,N_21551,N_24009);
and U25844 (N_25844,N_23188,N_24899);
nor U25845 (N_25845,N_24127,N_20060);
or U25846 (N_25846,N_21712,N_24641);
nand U25847 (N_25847,N_21703,N_20404);
and U25848 (N_25848,N_23276,N_22921);
xor U25849 (N_25849,N_23001,N_21183);
xnor U25850 (N_25850,N_23544,N_20526);
nand U25851 (N_25851,N_21820,N_20705);
nand U25852 (N_25852,N_21573,N_20813);
and U25853 (N_25853,N_24999,N_24918);
or U25854 (N_25854,N_22566,N_23335);
xnor U25855 (N_25855,N_22954,N_21107);
xor U25856 (N_25856,N_20468,N_22243);
or U25857 (N_25857,N_22062,N_23305);
and U25858 (N_25858,N_20393,N_20747);
xor U25859 (N_25859,N_24631,N_22833);
xor U25860 (N_25860,N_22101,N_23309);
and U25861 (N_25861,N_21309,N_20451);
xnor U25862 (N_25862,N_23799,N_24697);
or U25863 (N_25863,N_23032,N_23113);
xnor U25864 (N_25864,N_22164,N_21044);
xor U25865 (N_25865,N_23835,N_22217);
nand U25866 (N_25866,N_20975,N_21739);
xor U25867 (N_25867,N_20295,N_23099);
nor U25868 (N_25868,N_22880,N_20165);
nor U25869 (N_25869,N_23672,N_21663);
xor U25870 (N_25870,N_23375,N_20983);
and U25871 (N_25871,N_22095,N_20035);
and U25872 (N_25872,N_22025,N_24600);
xor U25873 (N_25873,N_24634,N_24489);
and U25874 (N_25874,N_24163,N_20528);
xor U25875 (N_25875,N_22011,N_23915);
nor U25876 (N_25876,N_21313,N_21525);
nor U25877 (N_25877,N_20274,N_20470);
or U25878 (N_25878,N_22909,N_23990);
and U25879 (N_25879,N_20075,N_20063);
xnor U25880 (N_25880,N_21207,N_23837);
or U25881 (N_25881,N_23583,N_23523);
and U25882 (N_25882,N_20009,N_23282);
nor U25883 (N_25883,N_22159,N_21797);
xnor U25884 (N_25884,N_24904,N_23693);
nor U25885 (N_25885,N_24037,N_21423);
and U25886 (N_25886,N_22392,N_23530);
or U25887 (N_25887,N_21302,N_22306);
nand U25888 (N_25888,N_20409,N_23302);
or U25889 (N_25889,N_23537,N_21709);
xor U25890 (N_25890,N_20746,N_24240);
nand U25891 (N_25891,N_24141,N_20287);
and U25892 (N_25892,N_23167,N_23145);
xnor U25893 (N_25893,N_21982,N_24100);
nand U25894 (N_25894,N_21738,N_24393);
and U25895 (N_25895,N_24851,N_21345);
or U25896 (N_25896,N_23482,N_21165);
nor U25897 (N_25897,N_23811,N_24033);
xor U25898 (N_25898,N_23374,N_22997);
nor U25899 (N_25899,N_21805,N_20929);
xnor U25900 (N_25900,N_20915,N_20905);
or U25901 (N_25901,N_20419,N_22809);
or U25902 (N_25902,N_20476,N_20557);
or U25903 (N_25903,N_21431,N_24555);
nand U25904 (N_25904,N_22219,N_22631);
and U25905 (N_25905,N_24835,N_23725);
and U25906 (N_25906,N_23112,N_20329);
nand U25907 (N_25907,N_22431,N_23679);
xor U25908 (N_25908,N_21859,N_22556);
xor U25909 (N_25909,N_24328,N_24859);
nand U25910 (N_25910,N_24510,N_23363);
nand U25911 (N_25911,N_23824,N_22260);
or U25912 (N_25912,N_21539,N_23606);
or U25913 (N_25913,N_23910,N_24583);
nand U25914 (N_25914,N_20084,N_22492);
xnor U25915 (N_25915,N_20355,N_23905);
or U25916 (N_25916,N_23826,N_23314);
nor U25917 (N_25917,N_21714,N_23258);
nor U25918 (N_25918,N_23495,N_24553);
xor U25919 (N_25919,N_20341,N_21536);
xnor U25920 (N_25920,N_23699,N_21334);
nor U25921 (N_25921,N_22632,N_22660);
and U25922 (N_25922,N_24278,N_21154);
xnor U25923 (N_25923,N_24540,N_23690);
nand U25924 (N_25924,N_24960,N_21822);
xnor U25925 (N_25925,N_20730,N_24063);
nand U25926 (N_25926,N_20006,N_23989);
or U25927 (N_25927,N_24028,N_22679);
or U25928 (N_25928,N_21648,N_23120);
nand U25929 (N_25929,N_21265,N_23710);
nand U25930 (N_25930,N_20053,N_21433);
nand U25931 (N_25931,N_23557,N_22114);
xor U25932 (N_25932,N_24420,N_24095);
or U25933 (N_25933,N_24291,N_22420);
nand U25934 (N_25934,N_24545,N_21115);
or U25935 (N_25935,N_23420,N_22970);
or U25936 (N_25936,N_23107,N_22048);
nor U25937 (N_25937,N_24317,N_22548);
nor U25938 (N_25938,N_21393,N_23405);
and U25939 (N_25939,N_20358,N_22093);
or U25940 (N_25940,N_23466,N_21913);
and U25941 (N_25941,N_22832,N_24092);
nor U25942 (N_25942,N_23490,N_21916);
or U25943 (N_25943,N_22875,N_20359);
nor U25944 (N_25944,N_24665,N_22626);
nor U25945 (N_25945,N_22511,N_23383);
nor U25946 (N_25946,N_22237,N_22299);
nor U25947 (N_25947,N_24529,N_21912);
nand U25948 (N_25948,N_20795,N_22251);
nand U25949 (N_25949,N_22689,N_23200);
nand U25950 (N_25950,N_22318,N_23463);
xor U25951 (N_25951,N_20950,N_23701);
and U25952 (N_25952,N_20937,N_23146);
nor U25953 (N_25953,N_20471,N_22195);
nor U25954 (N_25954,N_24642,N_20230);
and U25955 (N_25955,N_24650,N_21253);
and U25956 (N_25956,N_21971,N_20285);
or U25957 (N_25957,N_22499,N_22399);
nor U25958 (N_25958,N_21153,N_22695);
nand U25959 (N_25959,N_21952,N_23772);
or U25960 (N_25960,N_22174,N_24586);
nand U25961 (N_25961,N_20866,N_24723);
and U25962 (N_25962,N_20376,N_24351);
or U25963 (N_25963,N_21557,N_23733);
nor U25964 (N_25964,N_22640,N_24415);
nor U25965 (N_25965,N_24573,N_22422);
xor U25966 (N_25966,N_21950,N_21092);
nor U25967 (N_25967,N_21175,N_22953);
xor U25968 (N_25968,N_22113,N_22911);
or U25969 (N_25969,N_20906,N_22837);
and U25970 (N_25970,N_20583,N_21621);
and U25971 (N_25971,N_21697,N_23933);
xnor U25972 (N_25972,N_20863,N_20366);
xnor U25973 (N_25973,N_21560,N_22419);
nor U25974 (N_25974,N_23932,N_23517);
xor U25975 (N_25975,N_24625,N_23444);
and U25976 (N_25976,N_20502,N_23017);
or U25977 (N_25977,N_23010,N_24627);
nand U25978 (N_25978,N_22473,N_21876);
nand U25979 (N_25979,N_23380,N_24761);
nand U25980 (N_25980,N_22249,N_24012);
nand U25981 (N_25981,N_22507,N_23504);
and U25982 (N_25982,N_23588,N_20793);
xor U25983 (N_25983,N_24122,N_22784);
nor U25984 (N_25984,N_21564,N_23706);
xor U25985 (N_25985,N_20214,N_20181);
and U25986 (N_25986,N_23805,N_24640);
or U25987 (N_25987,N_22794,N_24480);
nand U25988 (N_25988,N_20996,N_24782);
nor U25989 (N_25989,N_24402,N_21781);
or U25990 (N_25990,N_21399,N_20658);
and U25991 (N_25991,N_22073,N_20223);
or U25992 (N_25992,N_21425,N_20826);
xnor U25993 (N_25993,N_24780,N_24900);
and U25994 (N_25994,N_23334,N_23403);
nor U25995 (N_25995,N_20467,N_20400);
or U25996 (N_25996,N_23597,N_24885);
nor U25997 (N_25997,N_20112,N_21501);
nand U25998 (N_25998,N_22490,N_24334);
nand U25999 (N_25999,N_21268,N_21863);
or U26000 (N_26000,N_23966,N_22575);
and U26001 (N_26001,N_22156,N_20728);
nand U26002 (N_26002,N_22487,N_21894);
xnor U26003 (N_26003,N_23691,N_20552);
xnor U26004 (N_26004,N_22034,N_21799);
xnor U26005 (N_26005,N_24488,N_20128);
nor U26006 (N_26006,N_23426,N_24023);
nand U26007 (N_26007,N_21796,N_23756);
and U26008 (N_26008,N_20278,N_20644);
xnor U26009 (N_26009,N_23881,N_21825);
nor U26010 (N_26010,N_21056,N_24630);
nand U26011 (N_26011,N_21288,N_20312);
or U26012 (N_26012,N_20395,N_22390);
or U26013 (N_26013,N_21908,N_22553);
xnor U26014 (N_26014,N_21227,N_21617);
nor U26015 (N_26015,N_23987,N_21266);
nor U26016 (N_26016,N_24544,N_24937);
nand U26017 (N_26017,N_22855,N_22683);
and U26018 (N_26018,N_21294,N_20668);
nor U26019 (N_26019,N_20005,N_23986);
nand U26020 (N_26020,N_24898,N_22882);
xnor U26021 (N_26021,N_21242,N_24067);
and U26022 (N_26022,N_20865,N_23300);
xnor U26023 (N_26023,N_20245,N_20986);
xor U26024 (N_26024,N_21272,N_24274);
or U26025 (N_26025,N_20725,N_21471);
nand U26026 (N_26026,N_20163,N_21046);
and U26027 (N_26027,N_20819,N_20670);
and U26028 (N_26028,N_24428,N_24868);
nand U26029 (N_26029,N_21186,N_21563);
xnor U26030 (N_26030,N_20556,N_24844);
xor U26031 (N_26031,N_24840,N_22036);
and U26032 (N_26032,N_23838,N_21138);
and U26033 (N_26033,N_20737,N_21053);
nor U26034 (N_26034,N_20420,N_20448);
nor U26035 (N_26035,N_23446,N_20094);
nand U26036 (N_26036,N_21027,N_24259);
and U26037 (N_26037,N_24836,N_24612);
nand U26038 (N_26038,N_22826,N_24520);
or U26039 (N_26039,N_24218,N_24073);
xnor U26040 (N_26040,N_20815,N_21386);
nand U26041 (N_26041,N_22234,N_22741);
or U26042 (N_26042,N_24404,N_21142);
xor U26043 (N_26043,N_23919,N_20757);
nor U26044 (N_26044,N_23654,N_21163);
xor U26045 (N_26045,N_23941,N_23858);
and U26046 (N_26046,N_21755,N_22012);
nor U26047 (N_26047,N_23581,N_22434);
and U26048 (N_26048,N_24307,N_23283);
xnor U26049 (N_26049,N_20438,N_24283);
nand U26050 (N_26050,N_21276,N_22273);
nand U26051 (N_26051,N_23492,N_21377);
nand U26052 (N_26052,N_20778,N_20897);
xnor U26053 (N_26053,N_22510,N_20045);
and U26054 (N_26054,N_24273,N_22464);
or U26055 (N_26055,N_21967,N_22316);
or U26056 (N_26056,N_22406,N_21326);
or U26057 (N_26057,N_22591,N_21232);
xor U26058 (N_26058,N_22815,N_23761);
and U26059 (N_26059,N_23326,N_20194);
xor U26060 (N_26060,N_24254,N_22146);
nor U26061 (N_26061,N_22751,N_20604);
xor U26062 (N_26062,N_21852,N_23911);
xnor U26063 (N_26063,N_21961,N_22948);
and U26064 (N_26064,N_22255,N_20566);
or U26065 (N_26065,N_23147,N_24892);
and U26066 (N_26066,N_22512,N_21658);
and U26067 (N_26067,N_24231,N_23876);
nand U26068 (N_26068,N_20011,N_23378);
or U26069 (N_26069,N_22454,N_21589);
or U26070 (N_26070,N_24116,N_21057);
and U26071 (N_26071,N_20637,N_21310);
and U26072 (N_26072,N_21480,N_24265);
and U26073 (N_26073,N_20365,N_22427);
nand U26074 (N_26074,N_21199,N_24737);
xnor U26075 (N_26075,N_22044,N_20949);
nor U26076 (N_26076,N_21422,N_20701);
xnor U26077 (N_26077,N_20512,N_21448);
and U26078 (N_26078,N_21645,N_22084);
and U26079 (N_26079,N_23961,N_24006);
xor U26080 (N_26080,N_24049,N_24592);
and U26081 (N_26081,N_24896,N_21694);
nand U26082 (N_26082,N_24453,N_22047);
xnor U26083 (N_26083,N_22386,N_24633);
nor U26084 (N_26084,N_23496,N_24304);
xnor U26085 (N_26085,N_22852,N_20379);
or U26086 (N_26086,N_20383,N_24238);
or U26087 (N_26087,N_21440,N_23716);
nor U26088 (N_26088,N_20487,N_24663);
nor U26089 (N_26089,N_22363,N_23311);
nor U26090 (N_26090,N_23263,N_23560);
nand U26091 (N_26091,N_20043,N_22630);
nand U26092 (N_26092,N_21134,N_20886);
or U26093 (N_26093,N_21569,N_23220);
or U26094 (N_26094,N_24977,N_24796);
nand U26095 (N_26095,N_21229,N_21506);
nor U26096 (N_26096,N_21583,N_24462);
and U26097 (N_26097,N_24839,N_24609);
and U26098 (N_26098,N_22181,N_20436);
nor U26099 (N_26099,N_20408,N_24590);
nand U26100 (N_26100,N_24311,N_21519);
or U26101 (N_26101,N_22545,N_21759);
nand U26102 (N_26102,N_21340,N_22256);
xor U26103 (N_26103,N_22200,N_24110);
nor U26104 (N_26104,N_22107,N_20113);
nor U26105 (N_26105,N_22698,N_24412);
nand U26106 (N_26106,N_21565,N_23418);
and U26107 (N_26107,N_24156,N_24601);
or U26108 (N_26108,N_22707,N_24719);
xor U26109 (N_26109,N_22172,N_23388);
nand U26110 (N_26110,N_23190,N_20726);
and U26111 (N_26111,N_24516,N_20354);
or U26112 (N_26112,N_22204,N_22010);
or U26113 (N_26113,N_23434,N_24310);
nor U26114 (N_26114,N_20029,N_24295);
xor U26115 (N_26115,N_21696,N_24752);
nand U26116 (N_26116,N_20424,N_24077);
xor U26117 (N_26117,N_22899,N_21304);
nand U26118 (N_26118,N_23603,N_20247);
xnor U26119 (N_26119,N_24502,N_23853);
nand U26120 (N_26120,N_21441,N_23815);
and U26121 (N_26121,N_21625,N_21121);
or U26122 (N_26122,N_21530,N_22972);
nor U26123 (N_26123,N_20059,N_22758);
or U26124 (N_26124,N_24125,N_22337);
xnor U26125 (N_26125,N_21909,N_24423);
or U26126 (N_26126,N_21917,N_21203);
nor U26127 (N_26127,N_20553,N_23534);
xor U26128 (N_26128,N_23918,N_23196);
and U26129 (N_26129,N_21267,N_22789);
or U26130 (N_26130,N_24691,N_21768);
and U26131 (N_26131,N_22319,N_20241);
nor U26132 (N_26132,N_22391,N_22721);
or U26133 (N_26133,N_23093,N_24378);
nand U26134 (N_26134,N_20978,N_24894);
nand U26135 (N_26135,N_21590,N_20922);
xnor U26136 (N_26136,N_24213,N_22493);
nor U26137 (N_26137,N_24626,N_23912);
nand U26138 (N_26138,N_20609,N_20462);
and U26139 (N_26139,N_23194,N_22442);
nor U26140 (N_26140,N_24433,N_22830);
xor U26141 (N_26141,N_24188,N_23633);
xor U26142 (N_26142,N_24301,N_23827);
or U26143 (N_26143,N_21866,N_22410);
xnor U26144 (N_26144,N_23361,N_21998);
xor U26145 (N_26145,N_21108,N_22326);
nand U26146 (N_26146,N_21899,N_22824);
xnor U26147 (N_26147,N_24774,N_24696);
nand U26148 (N_26148,N_21858,N_22615);
nor U26149 (N_26149,N_22308,N_20050);
or U26150 (N_26150,N_21957,N_20480);
nand U26151 (N_26151,N_22671,N_21404);
or U26152 (N_26152,N_21021,N_23518);
or U26153 (N_26153,N_24436,N_23651);
or U26154 (N_26154,N_21342,N_21084);
or U26155 (N_26155,N_21830,N_21382);
nand U26156 (N_26156,N_24088,N_23926);
nand U26157 (N_26157,N_22613,N_22644);
nor U26158 (N_26158,N_20007,N_21412);
or U26159 (N_26159,N_24332,N_22955);
nand U26160 (N_26160,N_21316,N_20715);
or U26161 (N_26161,N_22673,N_21581);
xor U26162 (N_26162,N_21951,N_21308);
and U26163 (N_26163,N_21818,N_21217);
nor U26164 (N_26164,N_24447,N_23235);
nor U26165 (N_26165,N_22547,N_23742);
nand U26166 (N_26166,N_20904,N_22714);
nor U26167 (N_26167,N_24946,N_24139);
nand U26168 (N_26168,N_21932,N_24419);
nand U26169 (N_26169,N_23313,N_21352);
nor U26170 (N_26170,N_22990,N_24054);
or U26171 (N_26171,N_22303,N_24287);
nor U26172 (N_26172,N_23077,N_20776);
and U26173 (N_26173,N_20942,N_21043);
xor U26174 (N_26174,N_23067,N_23427);
nor U26175 (N_26175,N_21173,N_21079);
xor U26176 (N_26176,N_22949,N_22216);
nand U26177 (N_26177,N_24271,N_22214);
xnor U26178 (N_26178,N_24795,N_23381);
or U26179 (N_26179,N_22108,N_21301);
nor U26180 (N_26180,N_22307,N_24784);
and U26181 (N_26181,N_23645,N_21545);
or U26182 (N_26182,N_21109,N_24998);
and U26183 (N_26183,N_23206,N_24950);
nand U26184 (N_26184,N_20282,N_23889);
or U26185 (N_26185,N_24338,N_21486);
xnor U26186 (N_26186,N_23985,N_23873);
nor U26187 (N_26187,N_22478,N_21467);
nand U26188 (N_26188,N_20628,N_23021);
or U26189 (N_26189,N_23333,N_20316);
and U26190 (N_26190,N_20784,N_23036);
nor U26191 (N_26191,N_21735,N_24245);
nor U26192 (N_26192,N_20333,N_22947);
xor U26193 (N_26193,N_23590,N_24253);
and U26194 (N_26194,N_22888,N_23839);
nor U26195 (N_26195,N_21460,N_23076);
xnor U26196 (N_26196,N_20145,N_22543);
xor U26197 (N_26197,N_22974,N_24756);
or U26198 (N_26198,N_24769,N_24621);
nand U26199 (N_26199,N_21584,N_20072);
nor U26200 (N_26200,N_24192,N_20690);
nor U26201 (N_26201,N_22270,N_22863);
xnor U26202 (N_26202,N_22501,N_23801);
nand U26203 (N_26203,N_24770,N_22330);
or U26204 (N_26204,N_20144,N_20342);
xnor U26205 (N_26205,N_22086,N_23788);
and U26206 (N_26206,N_23836,N_22612);
nor U26207 (N_26207,N_23494,N_24995);
or U26208 (N_26208,N_23764,N_20114);
or U26209 (N_26209,N_23711,N_22981);
or U26210 (N_26210,N_20437,N_20445);
nand U26211 (N_26211,N_20520,N_24659);
and U26212 (N_26212,N_24849,N_20610);
or U26213 (N_26213,N_24467,N_24388);
xnor U26214 (N_26214,N_20601,N_21745);
xnor U26215 (N_26215,N_20503,N_20588);
xor U26216 (N_26216,N_20031,N_21728);
nand U26217 (N_26217,N_23681,N_21062);
nor U26218 (N_26218,N_20659,N_24676);
nand U26219 (N_26219,N_20899,N_22388);
or U26220 (N_26220,N_23483,N_24790);
xor U26221 (N_26221,N_24375,N_20265);
and U26222 (N_26222,N_20244,N_22866);
nand U26223 (N_26223,N_22096,N_21126);
and U26224 (N_26224,N_22449,N_23248);
xnor U26225 (N_26225,N_23864,N_23584);
and U26226 (N_26226,N_22253,N_23398);
or U26227 (N_26227,N_21879,N_21737);
xor U26228 (N_26228,N_24897,N_21965);
nor U26229 (N_26229,N_20634,N_23628);
or U26230 (N_26230,N_22906,N_21274);
or U26231 (N_26231,N_24262,N_22240);
xnor U26232 (N_26232,N_21045,N_23652);
nand U26233 (N_26233,N_20741,N_24981);
and U26234 (N_26234,N_22916,N_20207);
nand U26235 (N_26235,N_22282,N_24399);
xor U26236 (N_26236,N_24196,N_22538);
xnor U26237 (N_26237,N_22652,N_21261);
nor U26238 (N_26238,N_23114,N_21401);
or U26239 (N_26239,N_22024,N_21102);
nor U26240 (N_26240,N_20246,N_23351);
and U26241 (N_26241,N_21690,N_22358);
nor U26242 (N_26242,N_20951,N_24509);
xnor U26243 (N_26243,N_23142,N_22285);
and U26244 (N_26244,N_21222,N_22793);
nor U26245 (N_26245,N_24134,N_23857);
or U26246 (N_26246,N_23433,N_20870);
and U26247 (N_26247,N_24877,N_20621);
and U26248 (N_26248,N_22604,N_21828);
and U26249 (N_26249,N_22192,N_23571);
and U26250 (N_26250,N_20618,N_21398);
nand U26251 (N_26251,N_24969,N_24563);
nand U26252 (N_26252,N_21426,N_24728);
and U26253 (N_26253,N_23771,N_21478);
or U26254 (N_26254,N_21582,N_23595);
nand U26255 (N_26255,N_20822,N_20875);
nor U26256 (N_26256,N_23339,N_22582);
and U26257 (N_26257,N_21117,N_20130);
nor U26258 (N_26258,N_20026,N_21840);
nand U26259 (N_26259,N_23812,N_23909);
or U26260 (N_26260,N_21458,N_21821);
nor U26261 (N_26261,N_24858,N_20170);
xnor U26262 (N_26262,N_24008,N_20491);
xor U26263 (N_26263,N_23747,N_24496);
xnor U26264 (N_26264,N_21935,N_21354);
and U26265 (N_26265,N_23319,N_21314);
or U26266 (N_26266,N_24257,N_21429);
nor U26267 (N_26267,N_24811,N_24666);
nor U26268 (N_26268,N_22836,N_20326);
and U26269 (N_26269,N_21958,N_24336);
nand U26270 (N_26270,N_21686,N_20799);
nand U26271 (N_26271,N_22150,N_22233);
and U26272 (N_26272,N_23087,N_24513);
or U26273 (N_26273,N_21851,N_23385);
and U26274 (N_26274,N_23831,N_21724);
and U26275 (N_26275,N_24680,N_21204);
xnor U26276 (N_26276,N_20569,N_21135);
nand U26277 (N_26277,N_22803,N_21311);
or U26278 (N_26278,N_23139,N_23620);
or U26279 (N_26279,N_22166,N_22744);
or U26280 (N_26280,N_22620,N_22853);
and U26281 (N_26281,N_20879,N_22567);
or U26282 (N_26282,N_23967,N_23792);
or U26283 (N_26283,N_23868,N_23895);
nand U26284 (N_26284,N_23315,N_21522);
and U26285 (N_26285,N_20431,N_23884);
nor U26286 (N_26286,N_23187,N_24771);
xnor U26287 (N_26287,N_20645,N_20619);
xor U26288 (N_26288,N_23245,N_23608);
or U26289 (N_26289,N_21926,N_21041);
nand U26290 (N_26290,N_22293,N_20997);
xnor U26291 (N_26291,N_22421,N_22407);
nor U26292 (N_26292,N_22785,N_24591);
xnor U26293 (N_26293,N_21727,N_24181);
nor U26294 (N_26294,N_22485,N_20787);
nand U26295 (N_26295,N_20710,N_20611);
xnor U26296 (N_26296,N_21208,N_23819);
nand U26297 (N_26297,N_22301,N_21730);
and U26298 (N_26298,N_20121,N_23043);
nand U26299 (N_26299,N_23766,N_21000);
or U26300 (N_26300,N_21798,N_22071);
nor U26301 (N_26301,N_23468,N_22674);
nor U26302 (N_26302,N_24395,N_23903);
and U26303 (N_26303,N_23743,N_22447);
nor U26304 (N_26304,N_20118,N_22021);
and U26305 (N_26305,N_24091,N_23279);
and U26306 (N_26306,N_24620,N_23594);
nand U26307 (N_26307,N_20674,N_20613);
nor U26308 (N_26308,N_20183,N_21225);
nand U26309 (N_26309,N_21947,N_22183);
nand U26310 (N_26310,N_24953,N_20801);
nor U26311 (N_26311,N_22246,N_22662);
or U26312 (N_26312,N_21752,N_22985);
or U26313 (N_26313,N_20211,N_20351);
and U26314 (N_26314,N_20998,N_21827);
xor U26315 (N_26315,N_23975,N_20861);
nand U26316 (N_26316,N_24611,N_23670);
nor U26317 (N_26317,N_23306,N_24543);
nor U26318 (N_26318,N_24233,N_22940);
or U26319 (N_26319,N_22436,N_20233);
xnor U26320 (N_26320,N_23415,N_22411);
xor U26321 (N_26321,N_21215,N_21248);
xor U26322 (N_26322,N_23545,N_21659);
nor U26323 (N_26323,N_24602,N_24909);
nor U26324 (N_26324,N_24746,N_21776);
or U26325 (N_26325,N_24312,N_20735);
nand U26326 (N_26326,N_22964,N_20104);
and U26327 (N_26327,N_23452,N_23456);
nor U26328 (N_26328,N_24807,N_21751);
or U26329 (N_26329,N_22051,N_24417);
nand U26330 (N_26330,N_20984,N_22452);
nand U26331 (N_26331,N_23073,N_23653);
xnor U26332 (N_26332,N_20190,N_22810);
or U26333 (N_26333,N_23744,N_24297);
nor U26334 (N_26334,N_24349,N_20884);
nand U26335 (N_26335,N_23549,N_22716);
or U26336 (N_26336,N_22989,N_22117);
or U26337 (N_26337,N_24905,N_20780);
or U26338 (N_26338,N_24989,N_22369);
or U26339 (N_26339,N_22137,N_24569);
xor U26340 (N_26340,N_20293,N_23246);
nand U26341 (N_26341,N_23442,N_24239);
nand U26342 (N_26342,N_21367,N_23965);
and U26343 (N_26343,N_21671,N_20952);
nor U26344 (N_26344,N_22157,N_24409);
nand U26345 (N_26345,N_21131,N_21264);
nor U26346 (N_26346,N_24681,N_24695);
and U26347 (N_26347,N_24076,N_20020);
and U26348 (N_26348,N_24050,N_24248);
nor U26349 (N_26349,N_23798,N_24597);
and U26350 (N_26350,N_24241,N_21664);
nand U26351 (N_26351,N_23917,N_21287);
and U26352 (N_26352,N_23769,N_23040);
nor U26353 (N_26353,N_24031,N_22252);
and U26354 (N_26354,N_20909,N_24082);
and U26355 (N_26355,N_24878,N_20484);
and U26356 (N_26356,N_20742,N_22334);
or U26357 (N_26357,N_23870,N_20862);
nand U26358 (N_26358,N_22726,N_21449);
or U26359 (N_26359,N_24373,N_22402);
nor U26360 (N_26360,N_22286,N_20079);
and U26361 (N_26361,N_21293,N_20301);
nand U26362 (N_26362,N_20160,N_21420);
or U26363 (N_26363,N_20450,N_22126);
nand U26364 (N_26364,N_22112,N_20683);
nor U26365 (N_26365,N_20417,N_22540);
or U26366 (N_26366,N_23215,N_23268);
xnor U26367 (N_26367,N_22209,N_23522);
or U26368 (N_26368,N_24445,N_23702);
nor U26369 (N_26369,N_22235,N_22503);
xor U26370 (N_26370,N_22788,N_21321);
and U26371 (N_26371,N_20033,N_21904);
or U26372 (N_26372,N_24580,N_21438);
or U26373 (N_26373,N_24617,N_24546);
or U26374 (N_26374,N_22298,N_23080);
and U26375 (N_26375,N_23758,N_21256);
nand U26376 (N_26376,N_21726,N_20414);
or U26377 (N_26377,N_22783,N_21657);
xor U26378 (N_26378,N_24029,N_20036);
xor U26379 (N_26379,N_23736,N_20348);
xnor U26380 (N_26380,N_24448,N_21038);
nand U26381 (N_26381,N_23115,N_23173);
nand U26382 (N_26382,N_21220,N_24729);
and U26383 (N_26383,N_24664,N_24416);
xor U26384 (N_26384,N_21493,N_24200);
xnor U26385 (N_26385,N_21753,N_21051);
nand U26386 (N_26386,N_24778,N_20103);
and U26387 (N_26387,N_23904,N_20322);
xnor U26388 (N_26388,N_22089,N_23973);
nor U26389 (N_26389,N_22975,N_20727);
nor U26390 (N_26390,N_24501,N_20030);
xor U26391 (N_26391,N_24536,N_21978);
or U26392 (N_26392,N_21350,N_22848);
or U26393 (N_26393,N_21640,N_24886);
xor U26394 (N_26394,N_21178,N_23643);
and U26395 (N_26395,N_20015,N_21254);
and U26396 (N_26396,N_24002,N_22629);
nor U26397 (N_26397,N_22820,N_24731);
or U26398 (N_26398,N_20560,N_20938);
or U26399 (N_26399,N_22614,N_23542);
nor U26400 (N_26400,N_21169,N_22321);
and U26401 (N_26401,N_24670,N_22812);
or U26402 (N_26402,N_20816,N_21836);
and U26403 (N_26403,N_20802,N_22524);
xor U26404 (N_26404,N_20109,N_20829);
and U26405 (N_26405,N_23790,N_23891);
or U26406 (N_26406,N_20515,N_20895);
and U26407 (N_26407,N_21615,N_21230);
or U26408 (N_26408,N_21491,N_20334);
or U26409 (N_26409,N_24800,N_20311);
xor U26410 (N_26410,N_24852,N_20013);
and U26411 (N_26411,N_20721,N_23038);
xnor U26412 (N_26412,N_21587,N_22122);
or U26413 (N_26413,N_23377,N_23355);
nand U26414 (N_26414,N_20661,N_23271);
or U26415 (N_26415,N_20720,N_23101);
nor U26416 (N_26416,N_23284,N_23554);
and U26417 (N_26417,N_24103,N_21945);
nand U26418 (N_26418,N_21259,N_22328);
nor U26419 (N_26419,N_21006,N_24368);
or U26420 (N_26420,N_22281,N_22834);
nor U26421 (N_26421,N_20340,N_21190);
nor U26422 (N_26422,N_21452,N_20082);
and U26423 (N_26423,N_22032,N_20172);
nor U26424 (N_26424,N_22465,N_22625);
or U26425 (N_26425,N_22562,N_24315);
nor U26426 (N_26426,N_20903,N_22681);
nand U26427 (N_26427,N_20716,N_22869);
xnor U26428 (N_26428,N_24133,N_20694);
and U26429 (N_26429,N_20519,N_22341);
nand U26430 (N_26430,N_24643,N_23406);
nand U26431 (N_26431,N_23536,N_24764);
or U26432 (N_26432,N_23344,N_21531);
xor U26433 (N_26433,N_24370,N_21592);
nand U26434 (N_26434,N_23353,N_24214);
and U26435 (N_26435,N_24721,N_23631);
or U26436 (N_26436,N_20577,N_24032);
nand U26437 (N_26437,N_20028,N_22059);
nand U26438 (N_26438,N_24794,N_24339);
or U26439 (N_26439,N_21211,N_23752);
nor U26440 (N_26440,N_20294,N_22352);
nor U26441 (N_26441,N_23871,N_24758);
nor U26442 (N_26442,N_23179,N_22980);
nand U26443 (N_26443,N_23502,N_23438);
and U26444 (N_26444,N_22365,N_20850);
xor U26445 (N_26445,N_22477,N_21344);
nor U26446 (N_26446,N_24403,N_20931);
nor U26447 (N_26447,N_24832,N_21769);
xor U26448 (N_26448,N_20707,N_21927);
and U26449 (N_26449,N_24296,N_20089);
and U26450 (N_26450,N_24685,N_24477);
nand U26451 (N_26451,N_24381,N_24861);
xor U26452 (N_26452,N_23875,N_23473);
and U26453 (N_26453,N_22912,N_22923);
xnor U26454 (N_26454,N_22193,N_23012);
xnor U26455 (N_26455,N_24986,N_23183);
or U26456 (N_26456,N_24394,N_23696);
nor U26457 (N_26457,N_20514,N_22708);
xor U26458 (N_26458,N_23041,N_24872);
and U26459 (N_26459,N_21787,N_22327);
nor U26460 (N_26460,N_20549,N_22865);
xor U26461 (N_26461,N_24827,N_21219);
nor U26462 (N_26462,N_22868,N_21461);
nand U26463 (N_26463,N_23061,N_20474);
nor U26464 (N_26464,N_21159,N_23327);
nor U26465 (N_26465,N_21348,N_22998);
or U26466 (N_26466,N_24688,N_21071);
nand U26467 (N_26467,N_20073,N_20123);
nor U26468 (N_26468,N_20367,N_23669);
nor U26469 (N_26469,N_23155,N_21869);
or U26470 (N_26470,N_20943,N_24963);
nor U26471 (N_26471,N_22268,N_20901);
or U26472 (N_26472,N_22481,N_20357);
or U26473 (N_26473,N_22272,N_21196);
nand U26474 (N_26474,N_24244,N_23360);
or U26475 (N_26475,N_20387,N_21403);
nor U26476 (N_26476,N_20052,N_22965);
nand U26477 (N_26477,N_23128,N_22435);
nor U26478 (N_26478,N_24753,N_22950);
nand U26479 (N_26479,N_20065,N_23960);
or U26480 (N_26480,N_22599,N_23485);
or U26481 (N_26481,N_21646,N_22570);
nand U26482 (N_26482,N_22177,N_23512);
xor U26483 (N_26483,N_24177,N_21468);
xor U26484 (N_26484,N_23779,N_21778);
xor U26485 (N_26485,N_24290,N_24478);
xor U26486 (N_26486,N_22397,N_23214);
nor U26487 (N_26487,N_22670,N_24161);
xor U26488 (N_26488,N_20212,N_24397);
or U26489 (N_26489,N_24255,N_20653);
and U26490 (N_26490,N_24818,N_24068);
or U26491 (N_26491,N_21462,N_20774);
and U26492 (N_26492,N_21705,N_21494);
xor U26493 (N_26493,N_21093,N_23707);
nor U26494 (N_26494,N_22368,N_22779);
xor U26495 (N_26495,N_23445,N_24199);
and U26496 (N_26496,N_22530,N_20580);
nor U26497 (N_26497,N_21080,N_20164);
or U26498 (N_26498,N_22799,N_20843);
nor U26499 (N_26499,N_21015,N_24371);
and U26500 (N_26500,N_23481,N_21720);
and U26501 (N_26501,N_20496,N_20392);
nand U26502 (N_26502,N_23293,N_24424);
xnor U26503 (N_26503,N_22514,N_23237);
and U26504 (N_26504,N_22488,N_23396);
nor U26505 (N_26505,N_23528,N_23619);
xor U26506 (N_26506,N_23848,N_21475);
nand U26507 (N_26507,N_20596,N_20473);
or U26508 (N_26508,N_23855,N_24727);
or U26509 (N_26509,N_23623,N_23148);
xnor U26510 (N_26510,N_23953,N_20948);
nand U26511 (N_26511,N_21247,N_23399);
nor U26512 (N_26512,N_23213,N_23832);
nand U26513 (N_26513,N_24500,N_21198);
and U26514 (N_26514,N_21090,N_24709);
nor U26515 (N_26515,N_21777,N_20490);
and U26516 (N_26516,N_20699,N_24389);
or U26517 (N_26517,N_20649,N_24155);
xnor U26518 (N_26518,N_24582,N_24470);
or U26519 (N_26519,N_24578,N_22018);
and U26520 (N_26520,N_24079,N_21801);
nor U26521 (N_26521,N_22827,N_23298);
or U26522 (N_26522,N_20132,N_21594);
or U26523 (N_26523,N_22991,N_22439);
or U26524 (N_26524,N_24493,N_24158);
nand U26525 (N_26525,N_21772,N_23940);
xor U26526 (N_26526,N_22536,N_24069);
xor U26527 (N_26527,N_24584,N_20298);
nand U26528 (N_26528,N_21245,N_22227);
nor U26529 (N_26529,N_20412,N_20988);
xor U26530 (N_26530,N_20847,N_21123);
and U26531 (N_26531,N_24211,N_23169);
and U26532 (N_26532,N_20346,N_21358);
and U26533 (N_26533,N_23467,N_22733);
or U26534 (N_26534,N_23943,N_23882);
nand U26535 (N_26535,N_21307,N_23783);
nand U26536 (N_26536,N_21258,N_22896);
and U26537 (N_26537,N_20466,N_23614);
nand U26538 (N_26538,N_24208,N_23324);
and U26539 (N_26539,N_21597,N_21390);
or U26540 (N_26540,N_22290,N_24515);
and U26541 (N_26541,N_20752,N_22154);
xor U26542 (N_26542,N_23058,N_20803);
and U26543 (N_26543,N_20231,N_23666);
and U26544 (N_26544,N_24773,N_24269);
nor U26545 (N_26545,N_20955,N_23576);
xor U26546 (N_26546,N_24097,N_24518);
or U26547 (N_26547,N_23211,N_20602);
xnor U26548 (N_26548,N_22527,N_23304);
and U26549 (N_26549,N_23297,N_24318);
or U26550 (N_26550,N_22469,N_21197);
nor U26551 (N_26551,N_20220,N_24252);
nand U26552 (N_26552,N_23830,N_24585);
nand U26553 (N_26553,N_22778,N_23781);
nand U26554 (N_26554,N_24121,N_21148);
nand U26555 (N_26555,N_24187,N_22703);
xor U26556 (N_26556,N_21255,N_24632);
nor U26557 (N_26557,N_21541,N_20957);
or U26558 (N_26558,N_20091,N_22935);
xor U26559 (N_26559,N_24128,N_20489);
nor U26560 (N_26560,N_24598,N_21920);
nor U26561 (N_26561,N_20666,N_20616);
nand U26562 (N_26562,N_21933,N_21164);
xnor U26563 (N_26563,N_20098,N_22893);
nor U26564 (N_26564,N_24649,N_21395);
xnor U26565 (N_26565,N_24364,N_23210);
and U26566 (N_26566,N_23901,N_24330);
or U26567 (N_26567,N_20680,N_24863);
or U26568 (N_26568,N_20585,N_22598);
xnor U26569 (N_26569,N_23734,N_24354);
nor U26570 (N_26570,N_22806,N_20782);
or U26571 (N_26571,N_22289,N_23338);
nand U26572 (N_26572,N_23277,N_20995);
xor U26573 (N_26573,N_22320,N_22026);
xnor U26574 (N_26574,N_23330,N_23104);
nand U26575 (N_26575,N_23863,N_24140);
and U26576 (N_26576,N_21010,N_21962);
xor U26577 (N_26577,N_21388,N_21874);
and U26578 (N_26578,N_21291,N_22792);
xnor U26579 (N_26579,N_23192,N_20671);
xor U26580 (N_26580,N_24604,N_24482);
and U26581 (N_26581,N_21896,N_22602);
nand U26582 (N_26582,N_22190,N_21793);
nor U26583 (N_26583,N_22265,N_20834);
and U26584 (N_26584,N_20236,N_24431);
nand U26585 (N_26585,N_21125,N_24983);
nand U26586 (N_26586,N_24915,N_20234);
nor U26587 (N_26587,N_22162,N_20651);
or U26588 (N_26588,N_23610,N_20629);
and U26589 (N_26589,N_24406,N_24922);
nor U26590 (N_26590,N_23540,N_20313);
nor U26591 (N_26591,N_20945,N_21838);
and U26592 (N_26592,N_20152,N_24007);
and U26593 (N_26593,N_24260,N_21609);
nor U26594 (N_26594,N_21191,N_22023);
nand U26595 (N_26595,N_20201,N_23753);
xnor U26596 (N_26596,N_20100,N_23988);
xnor U26597 (N_26597,N_23136,N_21680);
nand U26598 (N_26598,N_23796,N_24096);
nand U26599 (N_26599,N_23499,N_20791);
xor U26600 (N_26600,N_20516,N_24876);
xnor U26601 (N_26601,N_21127,N_20918);
nand U26602 (N_26602,N_23064,N_20771);
or U26603 (N_26603,N_23697,N_22719);
nor U26604 (N_26604,N_23205,N_22757);
or U26605 (N_26605,N_20991,N_21839);
and U26606 (N_26606,N_22486,N_24108);
xnor U26607 (N_26607,N_23421,N_22745);
nor U26608 (N_26608,N_20883,N_22723);
nand U26609 (N_26609,N_22856,N_23969);
xor U26610 (N_26610,N_20330,N_24281);
nand U26611 (N_26611,N_23599,N_22915);
xnor U26612 (N_26612,N_21548,N_23299);
and U26613 (N_26613,N_20388,N_22797);
or U26614 (N_26614,N_21606,N_24864);
or U26615 (N_26615,N_23157,N_21535);
and U26616 (N_26616,N_21273,N_21505);
nand U26617 (N_26617,N_23869,N_22339);
xnor U26618 (N_26618,N_22996,N_21662);
or U26619 (N_26619,N_24812,N_24554);
and U26620 (N_26620,N_24333,N_24272);
nor U26621 (N_26621,N_23667,N_20024);
nor U26622 (N_26622,N_21871,N_23429);
nor U26623 (N_26623,N_21435,N_21677);
nand U26624 (N_26624,N_20712,N_22860);
and U26625 (N_26625,N_24277,N_23464);
and U26626 (N_26626,N_24644,N_21626);
nand U26627 (N_26627,N_21353,N_21364);
or U26628 (N_26628,N_24483,N_23393);
and U26629 (N_26629,N_20264,N_22168);
or U26630 (N_26630,N_20548,N_21773);
and U26631 (N_26631,N_21444,N_23068);
nor U26632 (N_26632,N_22680,N_21834);
nand U26633 (N_26633,N_20890,N_21201);
and U26634 (N_26634,N_22879,N_20576);
nand U26635 (N_26635,N_20821,N_20472);
nand U26636 (N_26636,N_20956,N_22223);
and U26637 (N_26637,N_24084,N_21511);
or U26638 (N_26638,N_24465,N_21954);
and U26639 (N_26639,N_21347,N_20792);
or U26640 (N_26640,N_24010,N_22587);
nand U26641 (N_26641,N_24803,N_22142);
xnor U26642 (N_26642,N_21332,N_24279);
nand U26643 (N_26643,N_24495,N_24931);
xor U26644 (N_26644,N_22712,N_22999);
and U26645 (N_26645,N_22191,N_21375);
and U26646 (N_26646,N_23436,N_20756);
xnor U26647 (N_26647,N_24385,N_22900);
nand U26648 (N_26648,N_21857,N_21907);
xnor U26649 (N_26649,N_24550,N_23593);
nand U26650 (N_26650,N_20743,N_24735);
and U26651 (N_26651,N_20546,N_22908);
xnor U26652 (N_26652,N_20469,N_23787);
nor U26653 (N_26653,N_23825,N_21572);
or U26654 (N_26654,N_22654,N_20838);
and U26655 (N_26655,N_21214,N_21003);
and U26656 (N_26656,N_20695,N_23552);
and U26657 (N_26657,N_22780,N_21040);
and U26658 (N_26658,N_23978,N_21492);
nor U26659 (N_26659,N_23778,N_24862);
or U26660 (N_26660,N_24618,N_22746);
and U26661 (N_26661,N_20149,N_22913);
xnor U26662 (N_26662,N_20443,N_21103);
xor U26663 (N_26663,N_23908,N_23598);
nor U26664 (N_26664,N_22443,N_21715);
or U26665 (N_26665,N_22699,N_23402);
nand U26666 (N_26666,N_24376,N_24087);
or U26667 (N_26667,N_20586,N_24952);
nand U26668 (N_26668,N_20061,N_22647);
and U26669 (N_26669,N_22128,N_22158);
nor U26670 (N_26670,N_21983,N_23694);
nor U26671 (N_26671,N_20440,N_21861);
xor U26672 (N_26672,N_20428,N_20845);
or U26673 (N_26673,N_23253,N_22881);
xor U26674 (N_26674,N_20455,N_21428);
nor U26675 (N_26675,N_22090,N_20761);
nor U26676 (N_26676,N_22637,N_23387);
xnor U26677 (N_26677,N_20457,N_23984);
xor U26678 (N_26678,N_24930,N_21698);
nand U26679 (N_26679,N_21228,N_22437);
and U26680 (N_26680,N_24942,N_22724);
and U26681 (N_26681,N_21556,N_20603);
nand U26682 (N_26682,N_22438,N_22786);
xnor U26683 (N_26683,N_20605,N_24089);
xor U26684 (N_26684,N_24722,N_24306);
or U26685 (N_26685,N_23559,N_20745);
xor U26686 (N_26686,N_21389,N_23141);
and U26687 (N_26687,N_20083,N_24865);
xor U26688 (N_26688,N_20221,N_21414);
nand U26689 (N_26689,N_23303,N_21281);
and U26690 (N_26690,N_20808,N_20654);
or U26691 (N_26691,N_24786,N_21122);
nand U26692 (N_26692,N_21168,N_20430);
and U26693 (N_26693,N_21910,N_23119);
nor U26694 (N_26694,N_20608,N_23204);
or U26695 (N_26695,N_21779,N_21483);
and U26696 (N_26696,N_22429,N_21688);
xnor U26697 (N_26697,N_23615,N_20069);
nor U26698 (N_26698,N_22760,N_21052);
and U26699 (N_26699,N_21561,N_22466);
or U26700 (N_26700,N_24062,N_20369);
nor U26701 (N_26701,N_24679,N_20758);
nand U26702 (N_26702,N_20607,N_24203);
nor U26703 (N_26703,N_21944,N_23366);
nand U26704 (N_26704,N_22802,N_22554);
and U26705 (N_26705,N_22000,N_21442);
nor U26706 (N_26706,N_24531,N_20410);
nor U26707 (N_26707,N_24387,N_21979);
or U26708 (N_26708,N_22658,N_22951);
or U26709 (N_26709,N_23031,N_22092);
or U26710 (N_26710,N_23676,N_23118);
nor U26711 (N_26711,N_23365,N_24237);
or U26712 (N_26712,N_22850,N_21654);
nor U26713 (N_26713,N_24035,N_21224);
or U26714 (N_26714,N_22080,N_24202);
and U26715 (N_26715,N_22087,N_23023);
or U26716 (N_26716,N_24689,N_23459);
or U26717 (N_26717,N_24044,N_22292);
xnor U26718 (N_26718,N_20305,N_21014);
nand U26719 (N_26719,N_22133,N_24042);
nand U26720 (N_26720,N_22050,N_20642);
and U26721 (N_26721,N_24352,N_24179);
or U26722 (N_26722,N_23648,N_22774);
nor U26723 (N_26723,N_23566,N_20505);
nor U26724 (N_26724,N_22682,N_20296);
and U26725 (N_26725,N_21619,N_20345);
nand U26726 (N_26726,N_21605,N_24512);
or U26727 (N_26727,N_21489,N_21829);
nor U26728 (N_26728,N_22609,N_23191);
and U26729 (N_26729,N_23688,N_20349);
xor U26730 (N_26730,N_24623,N_23431);
xor U26731 (N_26731,N_24855,N_20250);
and U26732 (N_26732,N_22229,N_23221);
xnor U26733 (N_26733,N_20232,N_23982);
nand U26734 (N_26734,N_24026,N_21200);
or U26735 (N_26735,N_23569,N_24036);
nand U26736 (N_26736,N_22058,N_21192);
or U26737 (N_26737,N_20630,N_20562);
and U26738 (N_26738,N_22185,N_24101);
or U26739 (N_26739,N_22389,N_20660);
or U26740 (N_26740,N_24226,N_24973);
xnor U26741 (N_26741,N_23390,N_20614);
and U26742 (N_26742,N_21990,N_24051);
or U26743 (N_26743,N_23803,N_24123);
or U26744 (N_26744,N_22664,N_20025);
xnor U26745 (N_26745,N_24744,N_21479);
nand U26746 (N_26746,N_23950,N_23391);
or U26747 (N_26747,N_22455,N_23795);
or U26748 (N_26748,N_22284,N_23939);
nand U26749 (N_26749,N_24380,N_20315);
or U26750 (N_26750,N_20732,N_20663);
nand U26751 (N_26751,N_22266,N_24270);
and U26752 (N_26752,N_24090,N_21066);
and U26753 (N_26753,N_23236,N_20640);
or U26754 (N_26754,N_21510,N_20447);
or U26755 (N_26755,N_22943,N_24168);
xor U26756 (N_26756,N_22987,N_21867);
xnor U26757 (N_26757,N_20622,N_23567);
nand U26758 (N_26758,N_23618,N_22762);
and U26759 (N_26759,N_22359,N_22329);
nand U26760 (N_26760,N_23514,N_24914);
nand U26761 (N_26761,N_20116,N_24471);
xnor U26762 (N_26762,N_22655,N_20764);
and U26763 (N_26763,N_22078,N_21906);
and U26764 (N_26764,N_21948,N_21474);
nand U26765 (N_26765,N_21409,N_22845);
and U26766 (N_26766,N_20105,N_23320);
and U26767 (N_26767,N_20292,N_24779);
and U26768 (N_26768,N_22102,N_23898);
or U26769 (N_26769,N_21643,N_22070);
nor U26770 (N_26770,N_22259,N_20133);
or U26771 (N_26771,N_20806,N_24186);
and U26772 (N_26772,N_24616,N_24658);
xnor U26773 (N_26773,N_21567,N_21160);
nand U26774 (N_26774,N_22346,N_20099);
xor U26775 (N_26775,N_20125,N_23264);
nand U26776 (N_26776,N_22182,N_22666);
nor U26777 (N_26777,N_22103,N_20253);
xnor U26778 (N_26778,N_24384,N_24605);
nor U26779 (N_26779,N_20199,N_23738);
nor U26780 (N_26780,N_24320,N_21445);
and U26781 (N_26781,N_20175,N_21713);
or U26782 (N_26782,N_24703,N_20016);
nor U26783 (N_26783,N_23440,N_21534);
and U26784 (N_26784,N_24720,N_22610);
nor U26785 (N_26785,N_23717,N_22248);
and U26786 (N_26786,N_23417,N_20371);
xnor U26787 (N_26787,N_20001,N_23054);
xor U26788 (N_26788,N_22579,N_21788);
nor U26789 (N_26789,N_24030,N_24410);
xnor U26790 (N_26790,N_20977,N_22060);
nor U26791 (N_26791,N_24506,N_21653);
xor U26792 (N_26792,N_20198,N_23244);
nor U26793 (N_26793,N_20533,N_21323);
or U26794 (N_26794,N_23273,N_23443);
nor U26795 (N_26795,N_23890,N_20976);
or U26796 (N_26796,N_21666,N_24997);
and U26797 (N_26797,N_22356,N_22702);
and U26798 (N_26798,N_22489,N_20939);
and U26799 (N_26799,N_21450,N_23995);
xor U26800 (N_26800,N_21384,N_24475);
and U26801 (N_26801,N_23105,N_22593);
nand U26802 (N_26802,N_24675,N_24980);
or U26803 (N_26803,N_23617,N_20565);
nor U26804 (N_26804,N_20675,N_20873);
or U26805 (N_26805,N_22580,N_24124);
and U26806 (N_26806,N_20946,N_22841);
or U26807 (N_26807,N_24828,N_23461);
xnor U26808 (N_26808,N_22210,N_21701);
xor U26809 (N_26809,N_21166,N_24165);
nor U26810 (N_26810,N_24781,N_24498);
nor U26811 (N_26811,N_24850,N_23005);
or U26812 (N_26812,N_22002,N_22305);
nor U26813 (N_26813,N_24787,N_24109);
or U26814 (N_26814,N_20524,N_22928);
nand U26815 (N_26815,N_24041,N_23422);
nand U26816 (N_26816,N_22022,N_20530);
and U26817 (N_26817,N_23252,N_20039);
nand U26818 (N_26818,N_24418,N_21319);
and U26819 (N_26819,N_20111,N_23740);
nor U26820 (N_26820,N_24444,N_20226);
nand U26821 (N_26821,N_20023,N_24830);
nor U26822 (N_26822,N_22517,N_23325);
xor U26823 (N_26823,N_24710,N_24223);
and U26824 (N_26824,N_22740,N_20702);
xor U26825 (N_26825,N_20681,N_22904);
or U26826 (N_26826,N_24438,N_22686);
or U26827 (N_26827,N_22993,N_20593);
or U26828 (N_26828,N_21598,N_20356);
and U26829 (N_26829,N_23705,N_20689);
and U26830 (N_26830,N_20054,N_22123);
nand U26831 (N_26831,N_20759,N_20397);
nand U26832 (N_26832,N_24561,N_22669);
nor U26833 (N_26833,N_23469,N_21098);
and U26834 (N_26834,N_21096,N_20736);
xnor U26835 (N_26835,N_21780,N_23547);
and U26836 (N_26836,N_23274,N_23833);
nand U26837 (N_26837,N_23341,N_20336);
xor U26838 (N_26838,N_23301,N_20817);
xor U26839 (N_26839,N_22338,N_21939);
or U26840 (N_26840,N_22518,N_24701);
nor U26841 (N_26841,N_20180,N_21891);
and U26842 (N_26842,N_20126,N_21157);
xnor U26843 (N_26843,N_20381,N_21741);
nor U26844 (N_26844,N_21405,N_22475);
xor U26845 (N_26845,N_24034,N_21514);
or U26846 (N_26846,N_21477,N_22677);
and U26847 (N_26847,N_22097,N_24985);
and U26848 (N_26848,N_21678,N_24451);
or U26849 (N_26849,N_23241,N_24059);
nand U26850 (N_26850,N_20974,N_21427);
xor U26851 (N_26851,N_21815,N_21024);
nor U26852 (N_26852,N_21930,N_24822);
xor U26853 (N_26853,N_23084,N_20254);
or U26854 (N_26854,N_24667,N_23749);
nor U26855 (N_26855,N_21596,N_22230);
or U26856 (N_26856,N_22226,N_23218);
or U26857 (N_26857,N_22375,N_21576);
or U26858 (N_26858,N_20692,N_24927);
and U26859 (N_26859,N_21963,N_23580);
nor U26860 (N_26860,N_22764,N_22267);
or U26861 (N_26861,N_20964,N_20308);
xnor U26862 (N_26862,N_20571,N_23272);
or U26863 (N_26863,N_20754,N_24150);
or U26864 (N_26864,N_22572,N_24094);
nand U26865 (N_26865,N_21635,N_21498);
or U26866 (N_26866,N_20554,N_24825);
xnor U26867 (N_26867,N_23295,N_21077);
and U26868 (N_26868,N_23770,N_21454);
nand U26869 (N_26869,N_22902,N_22846);
nor U26870 (N_26870,N_20749,N_21622);
and U26871 (N_26871,N_24492,N_22944);
or U26872 (N_26872,N_21042,N_23509);
or U26873 (N_26873,N_22161,N_23722);
nor U26874 (N_26874,N_23677,N_23723);
or U26875 (N_26875,N_24884,N_23197);
xor U26876 (N_26876,N_20679,N_21193);
or U26877 (N_26877,N_22100,N_20697);
or U26878 (N_26878,N_23063,N_22672);
xor U26879 (N_26879,N_23541,N_22453);
or U26880 (N_26880,N_24360,N_23408);
nand U26881 (N_26881,N_23991,N_20401);
or U26882 (N_26882,N_20150,N_20887);
and U26883 (N_26883,N_21503,N_22471);
and U26884 (N_26884,N_20796,N_22361);
xor U26885 (N_26885,N_21171,N_24808);
and U26886 (N_26886,N_21430,N_24481);
or U26887 (N_26887,N_20289,N_23232);
nand U26888 (N_26888,N_21870,N_24705);
nand U26889 (N_26889,N_21868,N_20765);
and U26890 (N_26890,N_24143,N_23849);
xor U26891 (N_26891,N_23785,N_21900);
or U26892 (N_26892,N_24791,N_23936);
xnor U26893 (N_26893,N_23096,N_23947);
nand U26894 (N_26894,N_24114,N_24466);
nand U26895 (N_26895,N_23030,N_24775);
xor U26896 (N_26896,N_20032,N_24831);
and U26897 (N_26897,N_24411,N_22858);
nor U26898 (N_26898,N_22254,N_23843);
nand U26899 (N_26899,N_22395,N_20962);
or U26900 (N_26900,N_21176,N_21901);
or U26901 (N_26901,N_24210,N_22504);
xnor U26902 (N_26902,N_20936,N_23745);
nand U26903 (N_26903,N_23265,N_21031);
and U26904 (N_26904,N_22459,N_22706);
nand U26905 (N_26905,N_23394,N_24610);
and U26906 (N_26906,N_20159,N_20676);
xor U26907 (N_26907,N_21693,N_21782);
and U26908 (N_26908,N_20677,N_20389);
nor U26909 (N_26909,N_23996,N_22843);
or U26910 (N_26910,N_24286,N_24683);
and U26911 (N_26911,N_21497,N_24714);
nand U26912 (N_26912,N_22642,N_24046);
nor U26913 (N_26913,N_23700,N_21849);
and U26914 (N_26914,N_20597,N_20452);
xnor U26915 (N_26915,N_20475,N_22801);
xor U26916 (N_26916,N_22247,N_20143);
xnor U26917 (N_26917,N_24508,N_20229);
xor U26918 (N_26918,N_22245,N_22340);
xnor U26919 (N_26919,N_21118,N_23632);
xnor U26920 (N_26920,N_21937,N_21129);
or U26921 (N_26921,N_23002,N_24426);
xnor U26922 (N_26922,N_24441,N_23189);
nor U26923 (N_26923,N_24798,N_24154);
xnor U26924 (N_26924,N_22648,N_22035);
or U26925 (N_26925,N_20259,N_22544);
xor U26926 (N_26926,N_23414,N_22541);
nor U26927 (N_26927,N_22946,N_22939);
nor U26928 (N_26928,N_20578,N_23095);
or U26929 (N_26929,N_20360,N_20972);
and U26930 (N_26930,N_23003,N_24528);
or U26931 (N_26931,N_23278,N_24038);
and U26932 (N_26932,N_21030,N_24464);
xor U26933 (N_26933,N_22739,N_22495);
xnor U26934 (N_26934,N_22808,N_21140);
nor U26935 (N_26935,N_23098,N_23371);
nor U26936 (N_26936,N_23846,N_22574);
xnor U26937 (N_26937,N_20859,N_24442);
or U26938 (N_26938,N_23348,N_21843);
xnor U26939 (N_26939,N_21865,N_24303);
xor U26940 (N_26940,N_23015,N_22650);
and U26941 (N_26941,N_22942,N_22697);
xnor U26942 (N_26942,N_24733,N_20650);
nand U26943 (N_26943,N_23323,N_23867);
or U26944 (N_26944,N_23201,N_24460);
nor U26945 (N_26945,N_22938,N_22907);
nand U26946 (N_26946,N_20004,N_20042);
nor U26947 (N_26947,N_22167,N_21128);
nor U26948 (N_26948,N_21612,N_24917);
nand U26949 (N_26949,N_21396,N_23776);
and U26950 (N_26950,N_24335,N_20564);
and U26951 (N_26951,N_20283,N_22877);
or U26952 (N_26952,N_22017,N_22317);
nor U26953 (N_26953,N_24745,N_22094);
or U26954 (N_26954,N_22768,N_20458);
nand U26955 (N_26955,N_23945,N_21673);
or U26956 (N_26956,N_21591,N_22736);
or U26957 (N_26957,N_20718,N_21736);
nor U26958 (N_26958,N_21854,N_21507);
nand U26959 (N_26959,N_24282,N_21357);
nor U26960 (N_26960,N_22405,N_24045);
and U26961 (N_26961,N_22276,N_24105);
nor U26962 (N_26962,N_24820,N_21997);
xnor U26963 (N_26963,N_24131,N_23027);
or U26964 (N_26964,N_20501,N_21552);
nor U26965 (N_26965,N_21482,N_22578);
or U26966 (N_26966,N_24153,N_23242);
nor U26967 (N_26967,N_22873,N_23212);
nor U26968 (N_26968,N_23780,N_23916);
and U26969 (N_26969,N_20835,N_24309);
nor U26970 (N_26970,N_23944,N_24992);
xnor U26971 (N_26971,N_21734,N_20364);
and U26972 (N_26972,N_20902,N_24437);
nor U26973 (N_26973,N_23089,N_24107);
xor U26974 (N_26974,N_22787,N_20837);
nand U26975 (N_26975,N_20186,N_20242);
and U26976 (N_26976,N_20097,N_21048);
nand U26977 (N_26977,N_23820,N_21508);
and U26978 (N_26978,N_21580,N_20210);
nand U26979 (N_26979,N_20000,N_23234);
or U26980 (N_26980,N_23612,N_20435);
nor U26981 (N_26981,N_20405,N_24817);
or U26982 (N_26982,N_23718,N_20892);
or U26983 (N_26983,N_24021,N_23081);
and U26984 (N_26984,N_21124,N_20688);
or U26985 (N_26985,N_22139,N_24189);
or U26986 (N_26986,N_23249,N_21813);
nand U26987 (N_26987,N_23874,N_24699);
nand U26988 (N_26988,N_24730,N_23823);
and U26989 (N_26989,N_20693,N_20291);
and U26990 (N_26990,N_22484,N_24882);
and U26991 (N_26991,N_22003,N_23026);
or U26992 (N_26992,N_24837,N_21795);
nand U26993 (N_26993,N_23100,N_20898);
and U26994 (N_26994,N_20003,N_20896);
xor U26995 (N_26995,N_21419,N_22441);
and U26996 (N_26996,N_21966,N_23086);
xnor U26997 (N_26997,N_22201,N_24429);
or U26998 (N_26998,N_22175,N_22577);
and U26999 (N_26999,N_24962,N_24847);
nand U27000 (N_27000,N_22621,N_21149);
xnor U27001 (N_27001,N_21297,N_21465);
xor U27002 (N_27002,N_20647,N_21634);
nand U27003 (N_27003,N_23404,N_23719);
xor U27004 (N_27004,N_21767,N_24081);
nand U27005 (N_27005,N_22889,N_22897);
xor U27006 (N_27006,N_21685,N_21373);
xor U27007 (N_27007,N_21270,N_22754);
xnor U27008 (N_27008,N_24575,N_20723);
xor U27009 (N_27009,N_23329,N_21655);
nor U27010 (N_27010,N_22770,N_20087);
or U27011 (N_27011,N_23556,N_22497);
and U27012 (N_27012,N_21544,N_21034);
or U27013 (N_27013,N_23763,N_22467);
nand U27014 (N_27014,N_20276,N_21317);
and U27015 (N_27015,N_21614,N_23090);
nand U27016 (N_27016,N_21586,N_24430);
and U27017 (N_27017,N_23410,N_24994);
nand U27018 (N_27018,N_23174,N_21187);
or U27019 (N_27019,N_21394,N_22297);
xnor U27020 (N_27020,N_21011,N_23478);
or U27021 (N_27021,N_21763,N_21009);
or U27022 (N_27022,N_22147,N_24655);
nor U27023 (N_27023,N_22132,N_24577);
nand U27024 (N_27024,N_20286,N_24755);
or U27025 (N_27025,N_24027,N_24112);
or U27026 (N_27026,N_23122,N_20076);
xor U27027 (N_27027,N_21578,N_23640);
or U27028 (N_27028,N_21402,N_21886);
or U27029 (N_27029,N_22456,N_24367);
nor U27030 (N_27030,N_22323,N_24824);
or U27031 (N_27031,N_20390,N_21559);
xor U27032 (N_27032,N_23342,N_23661);
and U27033 (N_27033,N_22798,N_24651);
nor U27034 (N_27034,N_22218,N_22414);
nor U27035 (N_27035,N_22526,N_20320);
or U27036 (N_27036,N_22342,N_22269);
nor U27037 (N_27037,N_23856,N_21476);
or U27038 (N_27038,N_21184,N_23957);
xnor U27039 (N_27039,N_20599,N_23685);
xnor U27040 (N_27040,N_20135,N_23760);
xnor U27041 (N_27041,N_21647,N_23479);
nand U27042 (N_27042,N_24895,N_24957);
nor U27043 (N_27043,N_24537,N_23954);
nand U27044 (N_27044,N_23103,N_22901);
nor U27045 (N_27045,N_20378,N_23202);
nand U27046 (N_27046,N_23358,N_21004);
nor U27047 (N_27047,N_24959,N_22705);
nor U27048 (N_27048,N_23971,N_21075);
nor U27049 (N_27049,N_21516,N_22583);
or U27050 (N_27050,N_23045,N_20423);
xnor U27051 (N_27051,N_21172,N_21087);
xnor U27052 (N_27052,N_23585,N_22905);
nand U27053 (N_27053,N_20240,N_21832);
or U27054 (N_27054,N_22423,N_20970);
and U27055 (N_27055,N_23579,N_20189);
xnor U27056 (N_27056,N_23007,N_22257);
or U27057 (N_27057,N_21147,N_21660);
nor U27058 (N_27058,N_21495,N_20687);
and U27059 (N_27059,N_20682,N_24869);
or U27060 (N_27060,N_23750,N_20626);
or U27061 (N_27061,N_24738,N_22555);
xnor U27062 (N_27062,N_24976,N_23658);
or U27063 (N_27063,N_21439,N_21026);
or U27064 (N_27064,N_22225,N_21985);
nand U27065 (N_27065,N_23091,N_22867);
nand U27066 (N_27066,N_21887,N_22711);
xnor U27067 (N_27067,N_22013,N_23259);
nand U27068 (N_27068,N_22304,N_21633);
nand U27069 (N_27069,N_22472,N_22986);
xor U27070 (N_27070,N_23065,N_20243);
nand U27071 (N_27071,N_24678,N_21517);
and U27072 (N_27072,N_24058,N_22969);
nand U27073 (N_27073,N_24619,N_23257);
and U27074 (N_27074,N_22956,N_23182);
xor U27075 (N_27075,N_21682,N_24039);
and U27076 (N_27076,N_21981,N_23075);
and U27077 (N_27077,N_24221,N_21329);
xor U27078 (N_27078,N_22898,N_24443);
nand U27079 (N_27079,N_21959,N_24319);
or U27080 (N_27080,N_22448,N_20911);
nand U27081 (N_27081,N_22864,N_23108);
xnor U27082 (N_27082,N_20117,N_24901);
xnor U27083 (N_27083,N_20415,N_22006);
or U27084 (N_27084,N_24557,N_23092);
nor U27085 (N_27085,N_24576,N_20849);
and U27086 (N_27086,N_22480,N_23203);
nor U27087 (N_27087,N_23609,N_23505);
nor U27088 (N_27088,N_22688,N_20459);
or U27089 (N_27089,N_21447,N_22458);
nand U27090 (N_27090,N_21789,N_23151);
nand U27091 (N_27091,N_21020,N_22844);
xnor U27092 (N_27092,N_23181,N_24677);
nand U27093 (N_27093,N_24078,N_21400);
xor U27094 (N_27094,N_20779,N_20786);
nor U27095 (N_27095,N_24052,N_23498);
nand U27096 (N_27096,N_23948,N_23312);
nand U27097 (N_27097,N_21318,N_21929);
or U27098 (N_27098,N_24220,N_22224);
nor U27099 (N_27099,N_20377,N_22813);
nor U27100 (N_27100,N_21941,N_24560);
xnor U27101 (N_27101,N_24473,N_24759);
or U27102 (N_27102,N_22310,N_23364);
nand U27103 (N_27103,N_23963,N_21243);
and U27104 (N_27104,N_24854,N_20511);
xor U27105 (N_27105,N_22895,N_20066);
xnor U27106 (N_27106,N_24145,N_21081);
nand U27107 (N_27107,N_22505,N_24391);
or U27108 (N_27108,N_20928,N_20418);
nor U27109 (N_27109,N_22287,N_20279);
nor U27110 (N_27110,N_24236,N_21233);
xor U27111 (N_27111,N_22077,N_20840);
xnor U27112 (N_27112,N_21964,N_22668);
and U27113 (N_27113,N_23775,N_23178);
and U27114 (N_27114,N_24075,N_21890);
or U27115 (N_27115,N_24797,N_24463);
xor U27116 (N_27116,N_24672,N_20921);
nand U27117 (N_27117,N_22296,N_23786);
or U27118 (N_27118,N_22601,N_24261);
nand U27119 (N_27119,N_20989,N_22628);
nand U27120 (N_27120,N_20959,N_22314);
or U27121 (N_27121,N_21337,N_20338);
and U27122 (N_27122,N_24873,N_22715);
or U27123 (N_27123,N_20002,N_24048);
and U27124 (N_27124,N_23647,N_23130);
nand U27125 (N_27125,N_21942,N_24267);
or U27126 (N_27126,N_22542,N_20157);
or U27127 (N_27127,N_22525,N_20206);
nand U27128 (N_27128,N_22170,N_21328);
or U27129 (N_27129,N_23153,N_20871);
or U27130 (N_27130,N_20762,N_22874);
nor U27131 (N_27131,N_24157,N_22571);
xnor U27132 (N_27132,N_21144,N_20337);
and U27133 (N_27133,N_21684,N_21538);
and U27134 (N_27134,N_21327,N_23336);
xor U27135 (N_27135,N_21515,N_23935);
or U27136 (N_27136,N_22074,N_22959);
or U27137 (N_27137,N_22258,N_20790);
nor U27138 (N_27138,N_24228,N_24004);
nor U27139 (N_27139,N_24525,N_24019);
or U27140 (N_27140,N_24823,N_22584);
nand U27141 (N_27141,N_23465,N_23266);
and U27142 (N_27142,N_21018,N_21847);
xor U27143 (N_27143,N_21837,N_21143);
xnor U27144 (N_27144,N_21150,N_22687);
nor U27145 (N_27145,N_23352,N_23370);
nand U27146 (N_27146,N_23059,N_20625);
nand U27147 (N_27147,N_24593,N_22016);
and U27148 (N_27148,N_21251,N_22239);
and U27149 (N_27149,N_24098,N_21085);
nor U27150 (N_27150,N_20107,N_24505);
xor U27151 (N_27151,N_21610,N_23515);
nand U27152 (N_27152,N_20973,N_23240);
xor U27153 (N_27153,N_20426,N_24235);
or U27154 (N_27154,N_20267,N_20110);
xnor U27155 (N_27155,N_20363,N_21845);
nor U27156 (N_27156,N_22416,N_21188);
nand U27157 (N_27157,N_22135,N_24321);
nand U27158 (N_27158,N_21692,N_23834);
and U27159 (N_27159,N_22160,N_24366);
nor U27160 (N_27160,N_20056,N_22743);
and U27161 (N_27161,N_20672,N_24736);
nor U27162 (N_27162,N_23025,N_24344);
and U27163 (N_27163,N_21975,N_20120);
xor U27164 (N_27164,N_22791,N_22761);
and U27165 (N_27165,N_20891,N_20656);
or U27166 (N_27166,N_22360,N_21746);
or U27167 (N_27167,N_21361,N_24646);
or U27168 (N_27168,N_20980,N_21335);
or U27169 (N_27169,N_24967,N_20878);
xor U27170 (N_27170,N_22982,N_22883);
nor U27171 (N_27171,N_20508,N_21049);
and U27172 (N_27172,N_21300,N_21161);
nor U27173 (N_27173,N_22315,N_21372);
xnor U27174 (N_27174,N_23094,N_23035);
nand U27175 (N_27175,N_22141,N_20203);
and U27176 (N_27176,N_23765,N_20968);
and U27177 (N_27177,N_22854,N_21074);
nor U27178 (N_27178,N_24694,N_24919);
or U27179 (N_27179,N_24275,N_24635);
and U27180 (N_27180,N_23472,N_22560);
nor U27181 (N_27181,N_24434,N_23332);
xnor U27182 (N_27182,N_24383,N_23260);
xnor U27183 (N_27183,N_21817,N_23013);
nor U27184 (N_27184,N_23731,N_21792);
nand U27185 (N_27185,N_22203,N_22807);
xor U27186 (N_27186,N_23981,N_22535);
and U27187 (N_27187,N_21064,N_21570);
nand U27188 (N_27188,N_20979,N_20664);
nand U27189 (N_27189,N_24003,N_20064);
or U27190 (N_27190,N_21618,N_20372);
or U27191 (N_27191,N_23082,N_20623);
and U27192 (N_27192,N_23625,N_23878);
nor U27193 (N_27193,N_23150,N_24940);
xnor U27194 (N_27194,N_22728,N_23507);
and U27195 (N_27195,N_23346,N_23626);
nand U27196 (N_27196,N_20441,N_23616);
nor U27197 (N_27197,N_21141,N_24340);
nand U27198 (N_27198,N_22952,N_24661);
nand U27199 (N_27199,N_22825,N_24356);
nand U27200 (N_27200,N_23993,N_20606);
nand U27201 (N_27201,N_20544,N_21195);
or U27202 (N_27202,N_24549,N_20088);
or U27203 (N_27203,N_24323,N_20328);
xor U27204 (N_27204,N_20047,N_24162);
and U27205 (N_27205,N_24149,N_20251);
nand U27206 (N_27206,N_24587,N_24117);
or U27207 (N_27207,N_20738,N_23480);
nor U27208 (N_27208,N_22742,N_24766);
nand U27209 (N_27209,N_20635,N_21234);
nand U27210 (N_27210,N_21333,N_24939);
nand U27211 (N_27211,N_24708,N_24348);
nor U27212 (N_27212,N_21472,N_20429);
nand U27213 (N_27213,N_20517,N_21819);
xnor U27214 (N_27214,N_20406,N_24347);
nor U27215 (N_27215,N_20492,N_22262);
nor U27216 (N_27216,N_23828,N_24833);
nor U27217 (N_27217,N_21170,N_20139);
xor U27218 (N_27218,N_24043,N_20542);
xnor U27219 (N_27219,N_21528,N_23285);
nand U27220 (N_27220,N_23121,N_22663);
nand U27221 (N_27221,N_20807,N_23629);
and U27222 (N_27222,N_21262,N_21076);
or U27223 (N_27223,N_24949,N_24843);
nor U27224 (N_27224,N_24468,N_23955);
or U27225 (N_27225,N_23134,N_23937);
nor U27226 (N_27226,N_20804,N_21537);
or U27227 (N_27227,N_22033,N_24860);
nor U27228 (N_27228,N_20632,N_20179);
xor U27229 (N_27229,N_21549,N_21303);
nand U27230 (N_27230,N_24711,N_22533);
nand U27231 (N_27231,N_20638,N_20534);
nor U27232 (N_27232,N_22479,N_20335);
nor U27233 (N_27233,N_23972,N_23983);
nand U27234 (N_27234,N_21105,N_21808);
nor U27235 (N_27235,N_24614,N_24903);
nand U27236 (N_27236,N_21667,N_24446);
and U27237 (N_27237,N_24867,N_21451);
nor U27238 (N_27238,N_22876,N_23865);
or U27239 (N_27239,N_20842,N_23727);
nor U27240 (N_27240,N_20228,N_21638);
nor U27241 (N_27241,N_21411,N_21378);
or U27242 (N_27242,N_24857,N_24853);
nor U27243 (N_27243,N_23674,N_20846);
and U27244 (N_27244,N_23500,N_22957);
and U27245 (N_27245,N_21740,N_24250);
nor U27246 (N_27246,N_23998,N_22529);
and U27247 (N_27247,N_21679,N_22428);
xnor U27248 (N_27248,N_20216,N_23602);
xnor U27249 (N_27249,N_23124,N_21512);
xor U27250 (N_27250,N_23952,N_24938);
nor U27251 (N_27251,N_21226,N_20018);
nand U27252 (N_27252,N_20138,N_23683);
xnor U27253 (N_27253,N_24645,N_23217);
nor U27254 (N_27254,N_20657,N_21631);
and U27255 (N_27255,N_23070,N_23180);
xor U27256 (N_27256,N_24767,N_20851);
nor U27257 (N_27257,N_20080,N_22924);
or U27258 (N_27258,N_24268,N_23592);
nor U27259 (N_27259,N_24093,N_22639);
xor U27260 (N_27260,N_24421,N_24687);
nand U27261 (N_27261,N_24194,N_23822);
xnor U27262 (N_27262,N_23267,N_20350);
nor U27263 (N_27263,N_20481,N_20527);
and U27264 (N_27264,N_21733,N_21236);
nand U27265 (N_27265,N_22163,N_24816);
and U27266 (N_27266,N_23110,N_21094);
nand U27267 (N_27267,N_20402,N_22433);
nand U27268 (N_27268,N_23503,N_24978);
xor U27269 (N_27269,N_22782,N_23286);
or U27270 (N_27270,N_21848,N_22206);
and U27271 (N_27271,N_20095,N_21624);
nand U27272 (N_27272,N_24517,N_21977);
or U27273 (N_27273,N_20012,N_20643);
nor U27274 (N_27274,N_24215,N_24514);
nor U27275 (N_27275,N_23491,N_20545);
nand U27276 (N_27276,N_21766,N_22136);
nand U27277 (N_27277,N_21669,N_24374);
xnor U27278 (N_27278,N_24016,N_20920);
nor U27279 (N_27279,N_24887,N_22138);
or U27280 (N_27280,N_22528,N_24890);
xor U27281 (N_27281,N_21883,N_24251);
xnor U27282 (N_27282,N_22378,N_24657);
xnor U27283 (N_27283,N_20584,N_20235);
or U27284 (N_27284,N_22028,N_22418);
or U27285 (N_27285,N_21054,N_20034);
nand U27286 (N_27286,N_21707,N_22155);
nor U27287 (N_27287,N_21585,N_24083);
nand U27288 (N_27288,N_22001,N_22057);
and U27289 (N_27289,N_22847,N_23886);
nor U27290 (N_27290,N_21351,N_20646);
and U27291 (N_27291,N_21116,N_23821);
xor U27292 (N_27292,N_22228,N_22534);
or U27293 (N_27293,N_24057,N_23906);
nand U27294 (N_27294,N_23748,N_23844);
nor U27295 (N_27295,N_20506,N_21365);
nand U27296 (N_27296,N_22153,N_24175);
xnor U27297 (N_27297,N_20055,N_20731);
nand U27298 (N_27298,N_21139,N_22622);
xnor U27299 (N_27299,N_21114,N_22309);
xor U27300 (N_27300,N_22590,N_24698);
and U27301 (N_27301,N_23460,N_23527);
nor U27302 (N_27302,N_23601,N_24792);
xnor U27303 (N_27303,N_20339,N_24485);
xnor U27304 (N_27304,N_22008,N_23069);
or U27305 (N_27305,N_21487,N_23757);
nor U27306 (N_27306,N_23956,N_22732);
xor U27307 (N_27307,N_23074,N_23897);
and U27308 (N_27308,N_20062,N_21968);
nand U27309 (N_27309,N_23407,N_22054);
and U27310 (N_27310,N_21547,N_21880);
or U27311 (N_27311,N_20825,N_21221);
nand U27312 (N_27312,N_24806,N_20504);
and U27313 (N_27313,N_20617,N_20302);
or U27314 (N_27314,N_23083,N_22110);
nand U27315 (N_27315,N_21490,N_20197);
and U27316 (N_27316,N_20044,N_20563);
nand U27317 (N_27317,N_22444,N_20696);
and U27318 (N_27318,N_21473,N_23412);
xor U27319 (N_27319,N_22056,N_23152);
and U27320 (N_27320,N_21136,N_22934);
and U27321 (N_27321,N_20885,N_21835);
or U27322 (N_27322,N_23689,N_23024);
nand U27323 (N_27323,N_23441,N_22835);
xnor U27324 (N_27324,N_20248,N_20876);
nor U27325 (N_27325,N_21991,N_22675);
nand U27326 (N_27326,N_24941,N_20343);
nand U27327 (N_27327,N_21882,N_20398);
and U27328 (N_27328,N_20848,N_22149);
xnor U27329 (N_27329,N_23497,N_20280);
nor U27330 (N_27330,N_24014,N_22617);
or U27331 (N_27331,N_21532,N_23280);
and U27332 (N_27332,N_23475,N_23637);
and U27333 (N_27333,N_21455,N_23022);
and U27334 (N_27334,N_21914,N_20872);
nor U27335 (N_27335,N_20913,N_20925);
or U27336 (N_27336,N_20521,N_21286);
and U27337 (N_27337,N_20191,N_24842);
xnor U27338 (N_27338,N_24191,N_24503);
xor U27339 (N_27339,N_23568,N_24726);
or U27340 (N_27340,N_23154,N_24815);
or U27341 (N_27341,N_21185,N_21770);
or U27342 (N_27342,N_21695,N_24324);
or U27343 (N_27343,N_24020,N_21824);
nand U27344 (N_27344,N_21383,N_23208);
or U27345 (N_27345,N_20575,N_22430);
and U27346 (N_27346,N_24350,N_23928);
nor U27347 (N_27347,N_22717,N_23793);
nand U27348 (N_27348,N_21620,N_23880);
xor U27349 (N_27349,N_23938,N_20488);
nand U27350 (N_27350,N_23692,N_20711);
or U27351 (N_27351,N_21754,N_21500);
nand U27352 (N_27352,N_22772,N_24205);
or U27353 (N_27353,N_21341,N_22046);
xnor U27354 (N_27354,N_24299,N_20535);
nor U27355 (N_27355,N_24834,N_20734);
xor U27356 (N_27356,N_20288,N_23369);
and U27357 (N_27357,N_20856,N_21050);
xnor U27358 (N_27358,N_24574,N_24785);
and U27359 (N_27359,N_23703,N_22557);
xor U27360 (N_27360,N_22817,N_22005);
nor U27361 (N_27361,N_21675,N_21368);
nand U27362 (N_27362,N_24056,N_21063);
nand U27363 (N_27363,N_24848,N_24294);
or U27364 (N_27364,N_21145,N_22693);
or U27365 (N_27365,N_20839,N_20916);
or U27366 (N_27366,N_20176,N_23762);
or U27367 (N_27367,N_21111,N_22838);
xor U27368 (N_27368,N_21312,N_22750);
and U27369 (N_27369,N_21380,N_23797);
or U27370 (N_27370,N_23425,N_21290);
or U27371 (N_27371,N_21346,N_22357);
or U27372 (N_27372,N_22476,N_23562);
nor U27373 (N_27373,N_23550,N_20541);
nor U27374 (N_27374,N_20421,N_22829);
and U27375 (N_27375,N_20818,N_22222);
xnor U27376 (N_27376,N_21205,N_22596);
xor U27377 (N_27377,N_24018,N_21363);
xnor U27378 (N_27378,N_21603,N_23317);
nor U27379 (N_27379,N_24979,N_20464);
xnor U27380 (N_27380,N_24479,N_22118);
nor U27381 (N_27381,N_21366,N_23294);
or U27382 (N_27382,N_20257,N_20271);
nand U27383 (N_27383,N_20914,N_23546);
and U27384 (N_27384,N_22506,N_24511);
nor U27385 (N_27385,N_21260,N_24147);
nand U27386 (N_27386,N_24474,N_21812);
and U27387 (N_27387,N_20958,N_21194);
nor U27388 (N_27388,N_20249,N_22205);
or U27389 (N_27389,N_20202,N_21282);
or U27390 (N_27390,N_24120,N_24819);
and U27391 (N_27391,N_21237,N_22700);
xor U27392 (N_27392,N_23171,N_24243);
nand U27393 (N_27393,N_21499,N_22696);
and U27394 (N_27394,N_20154,N_23930);
nor U27395 (N_27395,N_20982,N_23548);
xor U27396 (N_27396,N_20966,N_21520);
xor U27397 (N_27397,N_24345,N_22616);
and U27398 (N_27398,N_22408,N_24916);
nand U27399 (N_27399,N_23604,N_21988);
and U27400 (N_27400,N_20740,N_21717);
and U27401 (N_27401,N_20173,N_22085);
or U27402 (N_27402,N_24207,N_23899);
xnor U27403 (N_27403,N_23340,N_20582);
nand U27404 (N_27404,N_24970,N_22851);
or U27405 (N_27405,N_24289,N_21110);
nor U27406 (N_27406,N_20090,N_23730);
nand U27407 (N_27407,N_23439,N_21823);
xor U27408 (N_27408,N_22977,N_21893);
xor U27409 (N_27409,N_23161,N_22502);
and U27410 (N_27410,N_20382,N_22045);
or U27411 (N_27411,N_23039,N_21543);
and U27412 (N_27412,N_24846,N_22597);
nor U27413 (N_27413,N_23322,N_20258);
nor U27414 (N_27414,N_21355,N_24242);
and U27415 (N_27415,N_21723,N_21437);
xor U27416 (N_27416,N_21275,N_22105);
and U27417 (N_27417,N_20115,N_21791);
or U27418 (N_27418,N_21636,N_23922);
xor U27419 (N_27419,N_23256,N_20559);
nand U27420 (N_27420,N_23524,N_24450);
xor U27421 (N_27421,N_20919,N_22646);
nor U27422 (N_27422,N_24538,N_22425);
xnor U27423 (N_27423,N_23347,N_23116);
nor U27424 (N_27424,N_21806,N_24193);
or U27425 (N_27425,N_21993,N_20587);
nand U27426 (N_27426,N_24810,N_24115);
and U27427 (N_27427,N_23659,N_23829);
or U27428 (N_27428,N_22515,N_23862);
xor U27429 (N_27429,N_23751,N_22232);
or U27430 (N_27430,N_21877,N_23033);
and U27431 (N_27431,N_22394,N_21055);
nand U27432 (N_27432,N_23635,N_22311);
or U27433 (N_27433,N_22220,N_23860);
or U27434 (N_27434,N_21443,N_23474);
nand U27435 (N_27435,N_24945,N_24652);
xor U27436 (N_27436,N_23269,N_23634);
nand U27437 (N_27437,N_21936,N_21073);
nor U27438 (N_27438,N_24990,N_22278);
and U27439 (N_27439,N_24929,N_21884);
or U27440 (N_27440,N_22960,N_24160);
or U27441 (N_27441,N_24595,N_20858);
nor U27442 (N_27442,N_21742,N_23879);
nor U27443 (N_27443,N_23896,N_21905);
xor U27444 (N_27444,N_21502,N_24400);
or U27445 (N_27445,N_24396,N_20153);
or U27446 (N_27446,N_23883,N_21218);
and U27447 (N_27447,N_23767,N_22775);
and U27448 (N_27448,N_24533,N_20685);
and U27449 (N_27449,N_23997,N_23165);
nand U27450 (N_27450,N_24264,N_22004);
or U27451 (N_27451,N_23784,N_24814);
nor U27452 (N_27452,N_20460,N_20495);
nor U27453 (N_27453,N_23644,N_21213);
nor U27454 (N_27454,N_20261,N_22068);
or U27455 (N_27455,N_21101,N_22805);
xnor U27456 (N_27456,N_23239,N_23262);
xnor U27457 (N_27457,N_22636,N_21775);
nor U27458 (N_27458,N_21761,N_21656);
nor U27459 (N_27459,N_20049,N_22558);
nor U27460 (N_27460,N_23572,N_22903);
nor U27461 (N_27461,N_22331,N_24201);
and U27462 (N_27462,N_23508,N_23923);
nand U27463 (N_27463,N_23732,N_21744);
nor U27464 (N_27464,N_22685,N_20499);
and U27465 (N_27465,N_22643,N_22983);
or U27466 (N_27466,N_21174,N_24206);
nor U27467 (N_27467,N_22513,N_21238);
nand U27468 (N_27468,N_23657,N_22821);
nand U27469 (N_27469,N_20195,N_21339);
nor U27470 (N_27470,N_22111,N_23066);
xnor U27471 (N_27471,N_21271,N_20612);
nor U27472 (N_27472,N_21279,N_20894);
nand U27473 (N_27473,N_24024,N_24322);
nand U27474 (N_27474,N_24499,N_24734);
or U27475 (N_27475,N_20078,N_21637);
nand U27476 (N_27476,N_23401,N_23968);
nand U27477 (N_27477,N_23316,N_20882);
xnor U27478 (N_27478,N_20373,N_24648);
and U27479 (N_27479,N_20662,N_21897);
nand U27480 (N_27480,N_20881,N_24883);
or U27481 (N_27481,N_21280,N_23424);
xor U27482 (N_27482,N_24183,N_20182);
or U27483 (N_27483,N_20917,N_20485);
or U27484 (N_27484,N_22348,N_24968);
and U27485 (N_27485,N_24639,N_21814);
or U27486 (N_27486,N_21523,N_22030);
nand U27487 (N_27487,N_21826,N_21065);
or U27488 (N_27488,N_23720,N_23673);
nor U27489 (N_27489,N_20600,N_23397);
or U27490 (N_27490,N_21881,N_24891);
nor U27491 (N_27491,N_22212,N_23019);
nand U27492 (N_27492,N_21179,N_23561);
xor U27493 (N_27493,N_24948,N_22735);
nand U27494 (N_27494,N_24102,N_21097);
nand U27495 (N_27495,N_24660,N_21356);
nand U27496 (N_27496,N_23109,N_24331);
nor U27497 (N_27497,N_20102,N_22194);
or U27498 (N_27498,N_24113,N_23639);
xnor U27499 (N_27499,N_24314,N_20070);
or U27500 (N_27500,N_21223,N_24264);
and U27501 (N_27501,N_22709,N_21483);
nand U27502 (N_27502,N_23715,N_22070);
xor U27503 (N_27503,N_23810,N_20928);
xnor U27504 (N_27504,N_20752,N_22653);
and U27505 (N_27505,N_23685,N_24596);
nand U27506 (N_27506,N_22301,N_24268);
nand U27507 (N_27507,N_21825,N_23441);
xor U27508 (N_27508,N_20464,N_22366);
and U27509 (N_27509,N_21882,N_24865);
nand U27510 (N_27510,N_20203,N_21897);
and U27511 (N_27511,N_23755,N_24796);
xnor U27512 (N_27512,N_23935,N_22098);
xor U27513 (N_27513,N_22901,N_24453);
xnor U27514 (N_27514,N_24805,N_22773);
nand U27515 (N_27515,N_21860,N_22798);
nand U27516 (N_27516,N_21302,N_23341);
xnor U27517 (N_27517,N_22114,N_23621);
and U27518 (N_27518,N_21693,N_22010);
xnor U27519 (N_27519,N_23385,N_23521);
xor U27520 (N_27520,N_24437,N_23518);
nand U27521 (N_27521,N_20314,N_23006);
or U27522 (N_27522,N_22397,N_23067);
xnor U27523 (N_27523,N_24523,N_21285);
or U27524 (N_27524,N_22371,N_24184);
or U27525 (N_27525,N_22260,N_21819);
and U27526 (N_27526,N_24154,N_22459);
nand U27527 (N_27527,N_22417,N_21592);
and U27528 (N_27528,N_24274,N_20385);
nand U27529 (N_27529,N_23218,N_22731);
xor U27530 (N_27530,N_21816,N_23066);
nor U27531 (N_27531,N_22126,N_24517);
nor U27532 (N_27532,N_24959,N_20547);
xnor U27533 (N_27533,N_24700,N_24653);
and U27534 (N_27534,N_24115,N_23193);
xnor U27535 (N_27535,N_24634,N_20339);
nand U27536 (N_27536,N_20172,N_22881);
xnor U27537 (N_27537,N_21208,N_22443);
nand U27538 (N_27538,N_20883,N_24338);
nand U27539 (N_27539,N_20540,N_22816);
nand U27540 (N_27540,N_20077,N_21556);
xnor U27541 (N_27541,N_24469,N_22012);
nand U27542 (N_27542,N_24831,N_21360);
xor U27543 (N_27543,N_22134,N_24545);
xor U27544 (N_27544,N_22377,N_21585);
nand U27545 (N_27545,N_20547,N_21447);
nor U27546 (N_27546,N_22981,N_23415);
nor U27547 (N_27547,N_22108,N_20344);
nand U27548 (N_27548,N_20772,N_21655);
xor U27549 (N_27549,N_20610,N_22862);
or U27550 (N_27550,N_20417,N_23702);
nand U27551 (N_27551,N_24236,N_23715);
nand U27552 (N_27552,N_24936,N_22213);
nand U27553 (N_27553,N_24216,N_24675);
and U27554 (N_27554,N_24092,N_24167);
nand U27555 (N_27555,N_20491,N_20633);
nand U27556 (N_27556,N_22482,N_22182);
or U27557 (N_27557,N_23320,N_21410);
or U27558 (N_27558,N_22631,N_24343);
nand U27559 (N_27559,N_22315,N_22226);
xor U27560 (N_27560,N_24706,N_21957);
or U27561 (N_27561,N_22920,N_24484);
and U27562 (N_27562,N_21590,N_24346);
nor U27563 (N_27563,N_22668,N_24788);
nor U27564 (N_27564,N_22032,N_22279);
nand U27565 (N_27565,N_23717,N_21875);
nor U27566 (N_27566,N_24713,N_20494);
nor U27567 (N_27567,N_22224,N_23109);
or U27568 (N_27568,N_22389,N_22659);
nand U27569 (N_27569,N_23384,N_21058);
nor U27570 (N_27570,N_22104,N_21957);
nor U27571 (N_27571,N_20494,N_24095);
and U27572 (N_27572,N_20685,N_22954);
nand U27573 (N_27573,N_24813,N_22292);
and U27574 (N_27574,N_23771,N_24843);
or U27575 (N_27575,N_22574,N_21590);
nor U27576 (N_27576,N_24256,N_23233);
nor U27577 (N_27577,N_23413,N_23932);
nor U27578 (N_27578,N_22480,N_21531);
nand U27579 (N_27579,N_20512,N_24341);
nor U27580 (N_27580,N_21441,N_21027);
nor U27581 (N_27581,N_21425,N_23699);
or U27582 (N_27582,N_21795,N_23186);
and U27583 (N_27583,N_20180,N_24058);
nand U27584 (N_27584,N_21823,N_22154);
nor U27585 (N_27585,N_22562,N_20130);
nand U27586 (N_27586,N_22627,N_21223);
and U27587 (N_27587,N_22594,N_24243);
nor U27588 (N_27588,N_21405,N_23446);
nor U27589 (N_27589,N_21713,N_24789);
or U27590 (N_27590,N_20763,N_24592);
or U27591 (N_27591,N_21636,N_24382);
and U27592 (N_27592,N_24079,N_22224);
nand U27593 (N_27593,N_20559,N_24934);
nor U27594 (N_27594,N_22278,N_24517);
or U27595 (N_27595,N_20383,N_24458);
nand U27596 (N_27596,N_23707,N_21678);
nor U27597 (N_27597,N_24386,N_22672);
nor U27598 (N_27598,N_21748,N_23265);
nand U27599 (N_27599,N_21494,N_24844);
or U27600 (N_27600,N_22230,N_20775);
nor U27601 (N_27601,N_22267,N_24256);
nand U27602 (N_27602,N_23183,N_21549);
xnor U27603 (N_27603,N_20410,N_21517);
nand U27604 (N_27604,N_21945,N_20251);
nand U27605 (N_27605,N_21953,N_23686);
or U27606 (N_27606,N_22548,N_22268);
xor U27607 (N_27607,N_20556,N_21618);
and U27608 (N_27608,N_22997,N_23361);
or U27609 (N_27609,N_22820,N_21036);
and U27610 (N_27610,N_23119,N_22132);
xnor U27611 (N_27611,N_24695,N_20458);
nand U27612 (N_27612,N_24207,N_21798);
nand U27613 (N_27613,N_21925,N_20163);
nand U27614 (N_27614,N_22082,N_23230);
and U27615 (N_27615,N_24590,N_22377);
and U27616 (N_27616,N_21753,N_22294);
nand U27617 (N_27617,N_23128,N_23777);
xnor U27618 (N_27618,N_23831,N_23913);
and U27619 (N_27619,N_21481,N_24557);
or U27620 (N_27620,N_22846,N_21919);
nand U27621 (N_27621,N_21726,N_23462);
or U27622 (N_27622,N_21917,N_23691);
nand U27623 (N_27623,N_20494,N_24087);
nor U27624 (N_27624,N_24872,N_22796);
nor U27625 (N_27625,N_22789,N_22495);
or U27626 (N_27626,N_24978,N_24716);
nor U27627 (N_27627,N_23126,N_23963);
nand U27628 (N_27628,N_22301,N_24224);
nor U27629 (N_27629,N_20801,N_22353);
nor U27630 (N_27630,N_23302,N_20926);
and U27631 (N_27631,N_22650,N_21800);
nor U27632 (N_27632,N_23187,N_24519);
xor U27633 (N_27633,N_22653,N_21480);
nand U27634 (N_27634,N_24501,N_24193);
xor U27635 (N_27635,N_22104,N_24210);
nand U27636 (N_27636,N_20456,N_22808);
and U27637 (N_27637,N_22100,N_21177);
nor U27638 (N_27638,N_24879,N_22382);
or U27639 (N_27639,N_24851,N_23722);
and U27640 (N_27640,N_24254,N_24746);
nand U27641 (N_27641,N_22127,N_21805);
nand U27642 (N_27642,N_24541,N_22690);
and U27643 (N_27643,N_22859,N_23401);
nor U27644 (N_27644,N_21620,N_23092);
nor U27645 (N_27645,N_20917,N_24080);
nor U27646 (N_27646,N_22871,N_20332);
nand U27647 (N_27647,N_20935,N_20523);
or U27648 (N_27648,N_22339,N_24847);
nor U27649 (N_27649,N_20642,N_24588);
nand U27650 (N_27650,N_23460,N_22147);
nand U27651 (N_27651,N_20412,N_23986);
and U27652 (N_27652,N_24095,N_23565);
xor U27653 (N_27653,N_24941,N_20719);
nor U27654 (N_27654,N_21983,N_24772);
nor U27655 (N_27655,N_22183,N_24764);
xor U27656 (N_27656,N_21864,N_20444);
nor U27657 (N_27657,N_23926,N_20618);
xor U27658 (N_27658,N_22146,N_23552);
xnor U27659 (N_27659,N_22417,N_22364);
and U27660 (N_27660,N_23286,N_23690);
nand U27661 (N_27661,N_22989,N_22032);
nor U27662 (N_27662,N_20685,N_23700);
nand U27663 (N_27663,N_22084,N_21144);
nand U27664 (N_27664,N_23179,N_20857);
xnor U27665 (N_27665,N_23046,N_24077);
xnor U27666 (N_27666,N_20529,N_24019);
nor U27667 (N_27667,N_20861,N_21642);
xnor U27668 (N_27668,N_21952,N_21400);
xor U27669 (N_27669,N_21487,N_21876);
xor U27670 (N_27670,N_21827,N_22260);
or U27671 (N_27671,N_24999,N_24144);
and U27672 (N_27672,N_23363,N_21979);
nand U27673 (N_27673,N_22764,N_23384);
xor U27674 (N_27674,N_20696,N_24977);
and U27675 (N_27675,N_21554,N_23109);
and U27676 (N_27676,N_22267,N_20577);
nand U27677 (N_27677,N_22307,N_20423);
xnor U27678 (N_27678,N_22301,N_24873);
nor U27679 (N_27679,N_22587,N_24052);
nand U27680 (N_27680,N_24545,N_21880);
xor U27681 (N_27681,N_20168,N_20385);
nor U27682 (N_27682,N_24820,N_20465);
or U27683 (N_27683,N_23334,N_24749);
or U27684 (N_27684,N_22959,N_21482);
or U27685 (N_27685,N_21833,N_23618);
xnor U27686 (N_27686,N_23890,N_24448);
or U27687 (N_27687,N_21551,N_21456);
or U27688 (N_27688,N_21409,N_22496);
or U27689 (N_27689,N_23375,N_21381);
or U27690 (N_27690,N_22045,N_20772);
and U27691 (N_27691,N_24646,N_20284);
or U27692 (N_27692,N_20899,N_23208);
xor U27693 (N_27693,N_22236,N_23408);
xnor U27694 (N_27694,N_23076,N_21451);
or U27695 (N_27695,N_20621,N_21517);
xor U27696 (N_27696,N_23639,N_20549);
nand U27697 (N_27697,N_24417,N_24875);
and U27698 (N_27698,N_20166,N_24188);
or U27699 (N_27699,N_20599,N_22699);
nor U27700 (N_27700,N_21518,N_24106);
or U27701 (N_27701,N_20939,N_21488);
nand U27702 (N_27702,N_21491,N_23023);
nand U27703 (N_27703,N_22468,N_22125);
nand U27704 (N_27704,N_21002,N_21871);
xnor U27705 (N_27705,N_20121,N_22091);
and U27706 (N_27706,N_24534,N_20704);
or U27707 (N_27707,N_22435,N_20990);
and U27708 (N_27708,N_20178,N_23443);
or U27709 (N_27709,N_23997,N_22745);
xnor U27710 (N_27710,N_21753,N_24416);
nand U27711 (N_27711,N_24893,N_24356);
nor U27712 (N_27712,N_22449,N_20138);
nor U27713 (N_27713,N_22645,N_22662);
and U27714 (N_27714,N_22356,N_21160);
xnor U27715 (N_27715,N_24042,N_24338);
nand U27716 (N_27716,N_22137,N_22111);
xor U27717 (N_27717,N_22838,N_24182);
and U27718 (N_27718,N_20483,N_22674);
or U27719 (N_27719,N_21276,N_21636);
xnor U27720 (N_27720,N_21073,N_21656);
or U27721 (N_27721,N_20010,N_21524);
and U27722 (N_27722,N_21947,N_20065);
xor U27723 (N_27723,N_24414,N_22493);
or U27724 (N_27724,N_22155,N_24669);
and U27725 (N_27725,N_24031,N_22917);
and U27726 (N_27726,N_24696,N_21363);
xnor U27727 (N_27727,N_20312,N_24474);
and U27728 (N_27728,N_24663,N_21666);
xor U27729 (N_27729,N_21041,N_22676);
and U27730 (N_27730,N_24407,N_22813);
xor U27731 (N_27731,N_22804,N_24712);
xor U27732 (N_27732,N_20114,N_20941);
xnor U27733 (N_27733,N_20916,N_23571);
and U27734 (N_27734,N_22858,N_20635);
and U27735 (N_27735,N_24970,N_20948);
and U27736 (N_27736,N_23221,N_23722);
or U27737 (N_27737,N_21091,N_23703);
and U27738 (N_27738,N_22907,N_21694);
nand U27739 (N_27739,N_24230,N_23016);
nor U27740 (N_27740,N_21082,N_21855);
and U27741 (N_27741,N_24360,N_21275);
nor U27742 (N_27742,N_22669,N_24983);
xor U27743 (N_27743,N_22853,N_21196);
xor U27744 (N_27744,N_22944,N_20085);
or U27745 (N_27745,N_21201,N_22842);
xor U27746 (N_27746,N_23514,N_23885);
or U27747 (N_27747,N_22208,N_20997);
and U27748 (N_27748,N_20019,N_21731);
nand U27749 (N_27749,N_22253,N_23174);
and U27750 (N_27750,N_24405,N_20469);
xor U27751 (N_27751,N_21883,N_23817);
and U27752 (N_27752,N_24681,N_24255);
nand U27753 (N_27753,N_23776,N_21179);
xor U27754 (N_27754,N_20176,N_20716);
nor U27755 (N_27755,N_22117,N_22116);
xnor U27756 (N_27756,N_24254,N_21697);
or U27757 (N_27757,N_22632,N_20371);
xnor U27758 (N_27758,N_23529,N_22010);
and U27759 (N_27759,N_23743,N_23369);
xnor U27760 (N_27760,N_23340,N_24634);
nor U27761 (N_27761,N_20093,N_22389);
xnor U27762 (N_27762,N_23477,N_24785);
xnor U27763 (N_27763,N_24128,N_20384);
or U27764 (N_27764,N_24685,N_23265);
nor U27765 (N_27765,N_23665,N_23770);
nand U27766 (N_27766,N_20955,N_23281);
nand U27767 (N_27767,N_24927,N_21765);
nor U27768 (N_27768,N_20774,N_23937);
nor U27769 (N_27769,N_21009,N_22173);
xor U27770 (N_27770,N_22667,N_22866);
and U27771 (N_27771,N_22869,N_21015);
nand U27772 (N_27772,N_20296,N_20757);
xnor U27773 (N_27773,N_20133,N_24218);
nor U27774 (N_27774,N_23023,N_22634);
nand U27775 (N_27775,N_24249,N_20029);
nor U27776 (N_27776,N_22049,N_24657);
nor U27777 (N_27777,N_23330,N_21086);
nor U27778 (N_27778,N_20261,N_20036);
or U27779 (N_27779,N_21221,N_22603);
nand U27780 (N_27780,N_24479,N_24375);
or U27781 (N_27781,N_24676,N_24957);
nand U27782 (N_27782,N_23890,N_24827);
and U27783 (N_27783,N_20589,N_23356);
and U27784 (N_27784,N_23137,N_24169);
nand U27785 (N_27785,N_20681,N_23014);
xnor U27786 (N_27786,N_23171,N_23367);
nand U27787 (N_27787,N_24643,N_20820);
and U27788 (N_27788,N_21015,N_24434);
and U27789 (N_27789,N_23484,N_22075);
and U27790 (N_27790,N_20417,N_24482);
and U27791 (N_27791,N_24495,N_21438);
or U27792 (N_27792,N_20259,N_21844);
nand U27793 (N_27793,N_20240,N_24712);
or U27794 (N_27794,N_24606,N_21842);
or U27795 (N_27795,N_22581,N_22960);
nor U27796 (N_27796,N_20307,N_24842);
nand U27797 (N_27797,N_22648,N_23522);
or U27798 (N_27798,N_20754,N_23999);
nand U27799 (N_27799,N_22779,N_24399);
and U27800 (N_27800,N_20446,N_22840);
or U27801 (N_27801,N_23323,N_24755);
or U27802 (N_27802,N_22814,N_24540);
xnor U27803 (N_27803,N_22311,N_22575);
xnor U27804 (N_27804,N_23182,N_21846);
nand U27805 (N_27805,N_20508,N_20281);
xnor U27806 (N_27806,N_21969,N_22082);
nor U27807 (N_27807,N_21194,N_23263);
nand U27808 (N_27808,N_23282,N_23795);
and U27809 (N_27809,N_20762,N_24042);
xor U27810 (N_27810,N_22361,N_21281);
xor U27811 (N_27811,N_20319,N_22324);
or U27812 (N_27812,N_21130,N_20811);
nor U27813 (N_27813,N_23307,N_24354);
nor U27814 (N_27814,N_21254,N_20396);
nor U27815 (N_27815,N_23866,N_22705);
and U27816 (N_27816,N_24690,N_24797);
nor U27817 (N_27817,N_24179,N_24592);
and U27818 (N_27818,N_22834,N_20195);
nor U27819 (N_27819,N_23477,N_22112);
nand U27820 (N_27820,N_22215,N_23371);
xnor U27821 (N_27821,N_21854,N_21576);
and U27822 (N_27822,N_23999,N_21313);
or U27823 (N_27823,N_23923,N_24038);
nor U27824 (N_27824,N_20026,N_24721);
or U27825 (N_27825,N_24845,N_21748);
and U27826 (N_27826,N_24275,N_24511);
and U27827 (N_27827,N_20674,N_21961);
xnor U27828 (N_27828,N_24274,N_23086);
and U27829 (N_27829,N_22440,N_22359);
nand U27830 (N_27830,N_22776,N_23422);
nand U27831 (N_27831,N_20778,N_20570);
xor U27832 (N_27832,N_24680,N_22821);
or U27833 (N_27833,N_22912,N_22736);
and U27834 (N_27834,N_22206,N_20855);
or U27835 (N_27835,N_21856,N_24092);
nor U27836 (N_27836,N_24577,N_24060);
nand U27837 (N_27837,N_22746,N_23231);
or U27838 (N_27838,N_21192,N_21452);
nand U27839 (N_27839,N_20703,N_24321);
xnor U27840 (N_27840,N_20446,N_21531);
nor U27841 (N_27841,N_22890,N_20793);
and U27842 (N_27842,N_23721,N_21203);
xnor U27843 (N_27843,N_22391,N_20483);
nor U27844 (N_27844,N_21534,N_22056);
and U27845 (N_27845,N_20634,N_23475);
nand U27846 (N_27846,N_24608,N_21328);
or U27847 (N_27847,N_21313,N_23698);
nand U27848 (N_27848,N_21178,N_22653);
or U27849 (N_27849,N_22442,N_24253);
xnor U27850 (N_27850,N_20252,N_20821);
xor U27851 (N_27851,N_24906,N_23171);
nand U27852 (N_27852,N_24583,N_24971);
nand U27853 (N_27853,N_24425,N_20784);
nor U27854 (N_27854,N_20801,N_21650);
nand U27855 (N_27855,N_21012,N_23216);
or U27856 (N_27856,N_24489,N_21948);
nand U27857 (N_27857,N_23269,N_22744);
or U27858 (N_27858,N_24065,N_20611);
xor U27859 (N_27859,N_20619,N_24564);
xor U27860 (N_27860,N_21228,N_23382);
nand U27861 (N_27861,N_23089,N_22641);
or U27862 (N_27862,N_22489,N_24417);
nand U27863 (N_27863,N_23332,N_24861);
xor U27864 (N_27864,N_21057,N_21413);
and U27865 (N_27865,N_23705,N_20875);
or U27866 (N_27866,N_24062,N_22034);
nor U27867 (N_27867,N_23668,N_20524);
nor U27868 (N_27868,N_24281,N_24163);
nand U27869 (N_27869,N_20366,N_20039);
xnor U27870 (N_27870,N_24743,N_24826);
xor U27871 (N_27871,N_20176,N_24626);
and U27872 (N_27872,N_21232,N_20239);
and U27873 (N_27873,N_20737,N_22511);
nand U27874 (N_27874,N_24804,N_21486);
xnor U27875 (N_27875,N_21739,N_22773);
or U27876 (N_27876,N_24337,N_21205);
or U27877 (N_27877,N_20574,N_21432);
and U27878 (N_27878,N_24983,N_20870);
xnor U27879 (N_27879,N_23920,N_23132);
and U27880 (N_27880,N_23381,N_24183);
xor U27881 (N_27881,N_22396,N_22577);
nor U27882 (N_27882,N_21022,N_22858);
nor U27883 (N_27883,N_23253,N_21130);
nor U27884 (N_27884,N_23635,N_21928);
or U27885 (N_27885,N_23983,N_21959);
nor U27886 (N_27886,N_21784,N_23120);
xor U27887 (N_27887,N_24922,N_24307);
xor U27888 (N_27888,N_22562,N_24774);
nor U27889 (N_27889,N_22956,N_20697);
xnor U27890 (N_27890,N_23632,N_20786);
xor U27891 (N_27891,N_21541,N_24311);
or U27892 (N_27892,N_23674,N_24348);
nor U27893 (N_27893,N_21841,N_23139);
nand U27894 (N_27894,N_21046,N_22708);
or U27895 (N_27895,N_23776,N_21521);
or U27896 (N_27896,N_23613,N_23405);
nand U27897 (N_27897,N_24778,N_23501);
xnor U27898 (N_27898,N_22609,N_21449);
nand U27899 (N_27899,N_20344,N_24917);
xnor U27900 (N_27900,N_20393,N_24232);
nor U27901 (N_27901,N_24621,N_20152);
xnor U27902 (N_27902,N_21765,N_20900);
nor U27903 (N_27903,N_23922,N_23226);
xor U27904 (N_27904,N_23668,N_24373);
nor U27905 (N_27905,N_20480,N_20974);
or U27906 (N_27906,N_21128,N_22154);
xnor U27907 (N_27907,N_23194,N_20241);
nor U27908 (N_27908,N_23005,N_24681);
and U27909 (N_27909,N_21223,N_23780);
xor U27910 (N_27910,N_21008,N_21814);
nand U27911 (N_27911,N_20669,N_21822);
or U27912 (N_27912,N_20485,N_20495);
nand U27913 (N_27913,N_23632,N_23223);
nor U27914 (N_27914,N_21766,N_21684);
or U27915 (N_27915,N_20138,N_20189);
and U27916 (N_27916,N_23671,N_20788);
and U27917 (N_27917,N_22872,N_24231);
or U27918 (N_27918,N_20010,N_23217);
nand U27919 (N_27919,N_21828,N_24796);
nand U27920 (N_27920,N_24456,N_23657);
xor U27921 (N_27921,N_21600,N_22326);
or U27922 (N_27922,N_21267,N_20433);
nor U27923 (N_27923,N_22130,N_22509);
or U27924 (N_27924,N_20639,N_21280);
nand U27925 (N_27925,N_20521,N_24340);
and U27926 (N_27926,N_20880,N_20317);
nand U27927 (N_27927,N_21369,N_21290);
nor U27928 (N_27928,N_20991,N_22226);
and U27929 (N_27929,N_23686,N_23450);
xnor U27930 (N_27930,N_22089,N_21278);
and U27931 (N_27931,N_23449,N_22774);
nand U27932 (N_27932,N_21650,N_21737);
xor U27933 (N_27933,N_20241,N_21811);
or U27934 (N_27934,N_23428,N_23422);
nor U27935 (N_27935,N_24319,N_21382);
nor U27936 (N_27936,N_23041,N_21276);
nand U27937 (N_27937,N_21187,N_23744);
or U27938 (N_27938,N_20001,N_24676);
or U27939 (N_27939,N_22674,N_24443);
nand U27940 (N_27940,N_20849,N_24604);
nor U27941 (N_27941,N_20553,N_20128);
or U27942 (N_27942,N_23499,N_20137);
xor U27943 (N_27943,N_21613,N_21977);
xor U27944 (N_27944,N_20911,N_23468);
nand U27945 (N_27945,N_23029,N_24155);
or U27946 (N_27946,N_20525,N_23985);
nand U27947 (N_27947,N_20902,N_23824);
or U27948 (N_27948,N_23748,N_22219);
xnor U27949 (N_27949,N_22311,N_22179);
nand U27950 (N_27950,N_22350,N_23635);
nand U27951 (N_27951,N_21646,N_21360);
nor U27952 (N_27952,N_21293,N_24400);
nor U27953 (N_27953,N_20321,N_21318);
and U27954 (N_27954,N_22073,N_23273);
nor U27955 (N_27955,N_20854,N_24348);
xor U27956 (N_27956,N_22438,N_24377);
or U27957 (N_27957,N_22280,N_21333);
xnor U27958 (N_27958,N_21462,N_23426);
nor U27959 (N_27959,N_21722,N_24048);
or U27960 (N_27960,N_23354,N_21709);
xnor U27961 (N_27961,N_21110,N_22031);
nand U27962 (N_27962,N_20696,N_20057);
xnor U27963 (N_27963,N_23144,N_21614);
xor U27964 (N_27964,N_21750,N_22114);
xnor U27965 (N_27965,N_22853,N_20799);
nand U27966 (N_27966,N_21892,N_21289);
and U27967 (N_27967,N_22960,N_20980);
xnor U27968 (N_27968,N_24535,N_24973);
xnor U27969 (N_27969,N_21154,N_23090);
nand U27970 (N_27970,N_20234,N_24744);
or U27971 (N_27971,N_24447,N_24556);
or U27972 (N_27972,N_23364,N_24684);
and U27973 (N_27973,N_22899,N_22758);
or U27974 (N_27974,N_20744,N_20619);
or U27975 (N_27975,N_20935,N_22659);
nor U27976 (N_27976,N_21205,N_21138);
or U27977 (N_27977,N_21541,N_21357);
or U27978 (N_27978,N_23882,N_21581);
and U27979 (N_27979,N_24259,N_24816);
xor U27980 (N_27980,N_23161,N_20699);
xnor U27981 (N_27981,N_20766,N_24533);
xor U27982 (N_27982,N_24022,N_23425);
nand U27983 (N_27983,N_22667,N_23517);
xor U27984 (N_27984,N_24638,N_22581);
and U27985 (N_27985,N_21724,N_24305);
xnor U27986 (N_27986,N_21663,N_20723);
nand U27987 (N_27987,N_22931,N_23125);
xnor U27988 (N_27988,N_22585,N_20844);
nand U27989 (N_27989,N_20997,N_22683);
xor U27990 (N_27990,N_20574,N_24218);
nand U27991 (N_27991,N_24400,N_22389);
nand U27992 (N_27992,N_21763,N_22047);
or U27993 (N_27993,N_23733,N_22460);
nand U27994 (N_27994,N_23985,N_23101);
nand U27995 (N_27995,N_24412,N_22594);
xnor U27996 (N_27996,N_23246,N_20958);
or U27997 (N_27997,N_22513,N_24849);
nand U27998 (N_27998,N_22701,N_20202);
nand U27999 (N_27999,N_24831,N_24973);
nand U28000 (N_28000,N_24357,N_24070);
and U28001 (N_28001,N_22611,N_20749);
xor U28002 (N_28002,N_24325,N_24930);
nand U28003 (N_28003,N_24859,N_22781);
and U28004 (N_28004,N_21539,N_22664);
or U28005 (N_28005,N_21248,N_20553);
nor U28006 (N_28006,N_22754,N_22427);
nand U28007 (N_28007,N_23950,N_20932);
and U28008 (N_28008,N_21409,N_24537);
and U28009 (N_28009,N_24454,N_23143);
xnor U28010 (N_28010,N_23002,N_22024);
nand U28011 (N_28011,N_24209,N_22017);
or U28012 (N_28012,N_23949,N_23231);
xor U28013 (N_28013,N_20715,N_20032);
and U28014 (N_28014,N_20020,N_23802);
and U28015 (N_28015,N_20188,N_22186);
nand U28016 (N_28016,N_24163,N_22315);
or U28017 (N_28017,N_21725,N_20317);
nand U28018 (N_28018,N_21891,N_21750);
and U28019 (N_28019,N_23073,N_21947);
nand U28020 (N_28020,N_23670,N_22456);
xor U28021 (N_28021,N_22381,N_20037);
nand U28022 (N_28022,N_23562,N_23784);
xnor U28023 (N_28023,N_20861,N_22444);
or U28024 (N_28024,N_20484,N_20660);
or U28025 (N_28025,N_22637,N_24932);
xor U28026 (N_28026,N_21391,N_22475);
or U28027 (N_28027,N_22022,N_22797);
and U28028 (N_28028,N_21909,N_21440);
nor U28029 (N_28029,N_22706,N_21120);
nand U28030 (N_28030,N_23639,N_24424);
xor U28031 (N_28031,N_20293,N_21453);
nor U28032 (N_28032,N_21083,N_22077);
nor U28033 (N_28033,N_24954,N_21387);
or U28034 (N_28034,N_21123,N_21332);
nand U28035 (N_28035,N_23553,N_21964);
xnor U28036 (N_28036,N_24436,N_24545);
nor U28037 (N_28037,N_24372,N_23516);
and U28038 (N_28038,N_21067,N_21740);
nand U28039 (N_28039,N_24842,N_20825);
xnor U28040 (N_28040,N_22228,N_20000);
nand U28041 (N_28041,N_24721,N_22255);
nor U28042 (N_28042,N_20713,N_22469);
xor U28043 (N_28043,N_20261,N_21762);
nand U28044 (N_28044,N_23753,N_24084);
nand U28045 (N_28045,N_24057,N_20855);
or U28046 (N_28046,N_23448,N_21405);
or U28047 (N_28047,N_24768,N_24650);
or U28048 (N_28048,N_21044,N_20647);
nand U28049 (N_28049,N_21674,N_23834);
and U28050 (N_28050,N_22944,N_20929);
nand U28051 (N_28051,N_23420,N_22741);
and U28052 (N_28052,N_21508,N_21594);
and U28053 (N_28053,N_21798,N_21782);
nand U28054 (N_28054,N_22925,N_23443);
or U28055 (N_28055,N_20449,N_24250);
nor U28056 (N_28056,N_24143,N_22247);
and U28057 (N_28057,N_24354,N_23327);
xor U28058 (N_28058,N_21733,N_24117);
xnor U28059 (N_28059,N_20240,N_23914);
and U28060 (N_28060,N_24616,N_24866);
or U28061 (N_28061,N_20742,N_21432);
or U28062 (N_28062,N_22186,N_24542);
xor U28063 (N_28063,N_24985,N_20638);
xnor U28064 (N_28064,N_20994,N_21022);
xnor U28065 (N_28065,N_23168,N_23854);
or U28066 (N_28066,N_21091,N_21087);
nand U28067 (N_28067,N_22095,N_24536);
xnor U28068 (N_28068,N_21332,N_23823);
xnor U28069 (N_28069,N_24479,N_22129);
and U28070 (N_28070,N_22738,N_22441);
or U28071 (N_28071,N_24932,N_24853);
xnor U28072 (N_28072,N_20716,N_20571);
nor U28073 (N_28073,N_20485,N_22830);
or U28074 (N_28074,N_21745,N_20374);
nor U28075 (N_28075,N_21818,N_23568);
xor U28076 (N_28076,N_22485,N_21669);
nand U28077 (N_28077,N_24587,N_24671);
nand U28078 (N_28078,N_20619,N_21055);
nor U28079 (N_28079,N_22406,N_21792);
nand U28080 (N_28080,N_21472,N_24423);
or U28081 (N_28081,N_20882,N_22625);
or U28082 (N_28082,N_22420,N_21687);
xor U28083 (N_28083,N_21671,N_20356);
nor U28084 (N_28084,N_22336,N_20982);
and U28085 (N_28085,N_21363,N_20939);
xnor U28086 (N_28086,N_23668,N_23115);
and U28087 (N_28087,N_21301,N_22536);
or U28088 (N_28088,N_21295,N_24729);
xor U28089 (N_28089,N_21677,N_21778);
or U28090 (N_28090,N_22104,N_23355);
nand U28091 (N_28091,N_23521,N_24794);
nand U28092 (N_28092,N_23457,N_23909);
xor U28093 (N_28093,N_22305,N_20786);
nand U28094 (N_28094,N_20348,N_22112);
and U28095 (N_28095,N_21853,N_21626);
nand U28096 (N_28096,N_21071,N_21969);
and U28097 (N_28097,N_21645,N_24580);
or U28098 (N_28098,N_24627,N_22736);
nand U28099 (N_28099,N_20910,N_21724);
and U28100 (N_28100,N_22592,N_24073);
and U28101 (N_28101,N_22931,N_24104);
nor U28102 (N_28102,N_21921,N_23322);
or U28103 (N_28103,N_23405,N_24654);
or U28104 (N_28104,N_21834,N_23889);
xnor U28105 (N_28105,N_24961,N_23698);
nor U28106 (N_28106,N_24170,N_24295);
nand U28107 (N_28107,N_21549,N_21360);
or U28108 (N_28108,N_21842,N_24199);
or U28109 (N_28109,N_23430,N_22411);
nor U28110 (N_28110,N_20352,N_20507);
xor U28111 (N_28111,N_22452,N_20589);
xnor U28112 (N_28112,N_21476,N_22334);
or U28113 (N_28113,N_22809,N_24128);
xnor U28114 (N_28114,N_24282,N_20689);
and U28115 (N_28115,N_22844,N_22171);
nor U28116 (N_28116,N_22654,N_22015);
xor U28117 (N_28117,N_21098,N_22582);
xor U28118 (N_28118,N_22705,N_20366);
and U28119 (N_28119,N_20416,N_22790);
or U28120 (N_28120,N_23220,N_20856);
nor U28121 (N_28121,N_21323,N_24430);
xor U28122 (N_28122,N_20554,N_23452);
xnor U28123 (N_28123,N_21687,N_23761);
nor U28124 (N_28124,N_24203,N_24920);
nor U28125 (N_28125,N_21275,N_20632);
nand U28126 (N_28126,N_22977,N_23699);
xor U28127 (N_28127,N_21575,N_23454);
and U28128 (N_28128,N_20115,N_20208);
and U28129 (N_28129,N_23173,N_24896);
or U28130 (N_28130,N_23885,N_22313);
or U28131 (N_28131,N_22416,N_20802);
nand U28132 (N_28132,N_24733,N_24457);
xnor U28133 (N_28133,N_20874,N_24364);
xnor U28134 (N_28134,N_20567,N_20259);
nor U28135 (N_28135,N_20092,N_23818);
nand U28136 (N_28136,N_20222,N_20988);
nor U28137 (N_28137,N_21300,N_22879);
or U28138 (N_28138,N_22011,N_24883);
nor U28139 (N_28139,N_20199,N_23366);
or U28140 (N_28140,N_24003,N_20249);
nand U28141 (N_28141,N_24733,N_20521);
and U28142 (N_28142,N_24611,N_22491);
xnor U28143 (N_28143,N_23482,N_21228);
or U28144 (N_28144,N_23432,N_24988);
nor U28145 (N_28145,N_23593,N_24150);
nor U28146 (N_28146,N_21539,N_21485);
or U28147 (N_28147,N_24465,N_23419);
nor U28148 (N_28148,N_22991,N_23711);
nor U28149 (N_28149,N_20940,N_20478);
or U28150 (N_28150,N_22704,N_21299);
nand U28151 (N_28151,N_20934,N_20927);
and U28152 (N_28152,N_22755,N_23008);
or U28153 (N_28153,N_21655,N_24018);
and U28154 (N_28154,N_22199,N_22170);
xnor U28155 (N_28155,N_24234,N_22167);
and U28156 (N_28156,N_21314,N_22508);
or U28157 (N_28157,N_20963,N_20800);
nand U28158 (N_28158,N_24178,N_24432);
and U28159 (N_28159,N_22356,N_21679);
nor U28160 (N_28160,N_20941,N_22769);
xnor U28161 (N_28161,N_20485,N_22233);
and U28162 (N_28162,N_21756,N_23796);
nor U28163 (N_28163,N_24858,N_24692);
nor U28164 (N_28164,N_21403,N_23418);
nand U28165 (N_28165,N_21988,N_20305);
nor U28166 (N_28166,N_21523,N_24663);
nand U28167 (N_28167,N_20428,N_21915);
or U28168 (N_28168,N_22083,N_22359);
nand U28169 (N_28169,N_23619,N_24192);
nand U28170 (N_28170,N_21472,N_24652);
nor U28171 (N_28171,N_22971,N_22657);
nor U28172 (N_28172,N_24471,N_21362);
and U28173 (N_28173,N_21363,N_20602);
xnor U28174 (N_28174,N_21807,N_23173);
xor U28175 (N_28175,N_20935,N_20855);
nand U28176 (N_28176,N_23036,N_20675);
or U28177 (N_28177,N_20671,N_23542);
or U28178 (N_28178,N_24278,N_23007);
nand U28179 (N_28179,N_21414,N_22546);
and U28180 (N_28180,N_20201,N_24009);
nand U28181 (N_28181,N_24415,N_20008);
xor U28182 (N_28182,N_21153,N_21651);
nand U28183 (N_28183,N_23170,N_22498);
and U28184 (N_28184,N_22679,N_23963);
xor U28185 (N_28185,N_20115,N_24760);
nand U28186 (N_28186,N_23580,N_21611);
xor U28187 (N_28187,N_20212,N_22885);
nor U28188 (N_28188,N_24727,N_22473);
xor U28189 (N_28189,N_22732,N_20773);
and U28190 (N_28190,N_24968,N_21277);
and U28191 (N_28191,N_21202,N_20123);
nand U28192 (N_28192,N_24925,N_23468);
and U28193 (N_28193,N_22301,N_20397);
nand U28194 (N_28194,N_22291,N_22570);
nor U28195 (N_28195,N_21854,N_22956);
xnor U28196 (N_28196,N_21546,N_20595);
or U28197 (N_28197,N_22683,N_22935);
xor U28198 (N_28198,N_23592,N_21696);
and U28199 (N_28199,N_21516,N_20029);
nand U28200 (N_28200,N_22283,N_24407);
or U28201 (N_28201,N_21525,N_22290);
nor U28202 (N_28202,N_21214,N_22089);
nor U28203 (N_28203,N_24080,N_20701);
or U28204 (N_28204,N_23267,N_22725);
xor U28205 (N_28205,N_22271,N_21726);
xnor U28206 (N_28206,N_21616,N_20270);
nand U28207 (N_28207,N_21551,N_22195);
or U28208 (N_28208,N_23666,N_22485);
xor U28209 (N_28209,N_21772,N_24720);
nor U28210 (N_28210,N_24658,N_21555);
and U28211 (N_28211,N_24095,N_22951);
or U28212 (N_28212,N_23584,N_21109);
or U28213 (N_28213,N_22907,N_24706);
nor U28214 (N_28214,N_23066,N_22606);
nand U28215 (N_28215,N_24585,N_21692);
xor U28216 (N_28216,N_22108,N_24155);
xor U28217 (N_28217,N_20199,N_24526);
nand U28218 (N_28218,N_21220,N_23649);
nor U28219 (N_28219,N_20827,N_20931);
or U28220 (N_28220,N_23317,N_21940);
xnor U28221 (N_28221,N_21444,N_24676);
nor U28222 (N_28222,N_23084,N_21903);
xor U28223 (N_28223,N_24054,N_23660);
or U28224 (N_28224,N_20850,N_23217);
nor U28225 (N_28225,N_23812,N_23233);
or U28226 (N_28226,N_24288,N_20812);
nand U28227 (N_28227,N_23863,N_21697);
nand U28228 (N_28228,N_20458,N_23264);
and U28229 (N_28229,N_22117,N_23904);
nand U28230 (N_28230,N_20659,N_24644);
or U28231 (N_28231,N_20279,N_22714);
and U28232 (N_28232,N_20532,N_24525);
and U28233 (N_28233,N_21406,N_20898);
nor U28234 (N_28234,N_20173,N_24622);
nor U28235 (N_28235,N_24796,N_22213);
nor U28236 (N_28236,N_21641,N_20158);
and U28237 (N_28237,N_23086,N_23422);
xnor U28238 (N_28238,N_23508,N_21522);
nand U28239 (N_28239,N_22099,N_20933);
xor U28240 (N_28240,N_23100,N_20220);
or U28241 (N_28241,N_22209,N_23968);
and U28242 (N_28242,N_20365,N_21617);
nor U28243 (N_28243,N_23770,N_22381);
nor U28244 (N_28244,N_24491,N_20839);
nand U28245 (N_28245,N_21241,N_23943);
nor U28246 (N_28246,N_24906,N_22170);
nor U28247 (N_28247,N_23619,N_23902);
and U28248 (N_28248,N_21872,N_21888);
and U28249 (N_28249,N_24319,N_23736);
nand U28250 (N_28250,N_22544,N_22129);
nor U28251 (N_28251,N_23412,N_24751);
nor U28252 (N_28252,N_23300,N_23203);
and U28253 (N_28253,N_23771,N_22754);
and U28254 (N_28254,N_21738,N_21986);
nor U28255 (N_28255,N_21535,N_21858);
or U28256 (N_28256,N_20487,N_20083);
or U28257 (N_28257,N_24779,N_24700);
xor U28258 (N_28258,N_23825,N_20208);
and U28259 (N_28259,N_23904,N_22547);
xor U28260 (N_28260,N_23715,N_21952);
or U28261 (N_28261,N_21188,N_24614);
xor U28262 (N_28262,N_24679,N_23046);
nor U28263 (N_28263,N_22480,N_22477);
nor U28264 (N_28264,N_21976,N_20095);
nand U28265 (N_28265,N_21364,N_20091);
and U28266 (N_28266,N_20984,N_23637);
nand U28267 (N_28267,N_23664,N_23981);
nor U28268 (N_28268,N_20370,N_23998);
xnor U28269 (N_28269,N_24692,N_23860);
xor U28270 (N_28270,N_24951,N_24474);
or U28271 (N_28271,N_22378,N_20410);
xnor U28272 (N_28272,N_24594,N_24960);
nor U28273 (N_28273,N_23691,N_24687);
nor U28274 (N_28274,N_24713,N_23210);
nand U28275 (N_28275,N_20367,N_24912);
or U28276 (N_28276,N_21996,N_22956);
and U28277 (N_28277,N_21395,N_22130);
xor U28278 (N_28278,N_22111,N_21508);
xnor U28279 (N_28279,N_20658,N_24722);
xnor U28280 (N_28280,N_20890,N_20318);
xor U28281 (N_28281,N_20658,N_21418);
or U28282 (N_28282,N_23543,N_20191);
nor U28283 (N_28283,N_24607,N_24884);
and U28284 (N_28284,N_23566,N_23521);
nor U28285 (N_28285,N_23685,N_24019);
and U28286 (N_28286,N_21252,N_23653);
or U28287 (N_28287,N_21245,N_21807);
nand U28288 (N_28288,N_22673,N_23785);
nand U28289 (N_28289,N_22088,N_24770);
nor U28290 (N_28290,N_21056,N_21786);
nor U28291 (N_28291,N_24692,N_22671);
and U28292 (N_28292,N_23935,N_22224);
or U28293 (N_28293,N_23237,N_22040);
and U28294 (N_28294,N_20039,N_24206);
xor U28295 (N_28295,N_21228,N_24446);
nor U28296 (N_28296,N_23793,N_24790);
nand U28297 (N_28297,N_23539,N_20566);
nor U28298 (N_28298,N_20835,N_21084);
or U28299 (N_28299,N_20505,N_22188);
nand U28300 (N_28300,N_22249,N_21601);
xnor U28301 (N_28301,N_21623,N_23841);
or U28302 (N_28302,N_22294,N_22172);
nand U28303 (N_28303,N_20825,N_22378);
or U28304 (N_28304,N_22552,N_22485);
nand U28305 (N_28305,N_21326,N_24829);
and U28306 (N_28306,N_20978,N_22182);
or U28307 (N_28307,N_22001,N_23366);
nand U28308 (N_28308,N_22983,N_24580);
nor U28309 (N_28309,N_20094,N_20283);
and U28310 (N_28310,N_24673,N_21742);
xor U28311 (N_28311,N_21876,N_20694);
or U28312 (N_28312,N_24599,N_20278);
nor U28313 (N_28313,N_23616,N_21911);
or U28314 (N_28314,N_22621,N_22237);
or U28315 (N_28315,N_23688,N_20781);
nor U28316 (N_28316,N_24775,N_23636);
xor U28317 (N_28317,N_23857,N_24237);
or U28318 (N_28318,N_23771,N_20570);
nand U28319 (N_28319,N_23961,N_20293);
nand U28320 (N_28320,N_20281,N_21601);
nor U28321 (N_28321,N_22924,N_20674);
nand U28322 (N_28322,N_20581,N_23965);
and U28323 (N_28323,N_22254,N_20092);
and U28324 (N_28324,N_22249,N_23648);
nand U28325 (N_28325,N_24557,N_24622);
nor U28326 (N_28326,N_22706,N_20104);
and U28327 (N_28327,N_21190,N_21566);
nor U28328 (N_28328,N_22332,N_20176);
and U28329 (N_28329,N_23652,N_22144);
or U28330 (N_28330,N_23829,N_23292);
xnor U28331 (N_28331,N_20596,N_24289);
or U28332 (N_28332,N_20099,N_23308);
nand U28333 (N_28333,N_22329,N_21927);
xor U28334 (N_28334,N_22252,N_20888);
and U28335 (N_28335,N_23092,N_21427);
or U28336 (N_28336,N_23344,N_24802);
nand U28337 (N_28337,N_20924,N_24758);
nor U28338 (N_28338,N_23469,N_23703);
or U28339 (N_28339,N_20538,N_24905);
nand U28340 (N_28340,N_23838,N_20125);
nor U28341 (N_28341,N_20707,N_23285);
xor U28342 (N_28342,N_23443,N_23389);
nor U28343 (N_28343,N_20829,N_21132);
and U28344 (N_28344,N_22556,N_23455);
xor U28345 (N_28345,N_22515,N_24621);
nor U28346 (N_28346,N_23282,N_23545);
xnor U28347 (N_28347,N_20086,N_24642);
nand U28348 (N_28348,N_20807,N_20461);
or U28349 (N_28349,N_22775,N_22936);
and U28350 (N_28350,N_20740,N_22777);
xor U28351 (N_28351,N_21721,N_23210);
or U28352 (N_28352,N_24758,N_24724);
and U28353 (N_28353,N_22299,N_24713);
xnor U28354 (N_28354,N_23169,N_23726);
nand U28355 (N_28355,N_21734,N_21767);
nand U28356 (N_28356,N_23320,N_21397);
and U28357 (N_28357,N_23500,N_21648);
xnor U28358 (N_28358,N_24940,N_21354);
xor U28359 (N_28359,N_22431,N_22648);
and U28360 (N_28360,N_23894,N_23799);
xnor U28361 (N_28361,N_24701,N_23194);
and U28362 (N_28362,N_21047,N_20112);
xor U28363 (N_28363,N_21926,N_22945);
xor U28364 (N_28364,N_21553,N_24058);
nand U28365 (N_28365,N_20863,N_23625);
xnor U28366 (N_28366,N_21451,N_24326);
nand U28367 (N_28367,N_20310,N_20253);
or U28368 (N_28368,N_24249,N_21094);
xnor U28369 (N_28369,N_20665,N_22849);
nand U28370 (N_28370,N_21958,N_24404);
xor U28371 (N_28371,N_23835,N_24527);
nor U28372 (N_28372,N_22139,N_22103);
and U28373 (N_28373,N_20658,N_23725);
and U28374 (N_28374,N_23046,N_23765);
nand U28375 (N_28375,N_23526,N_21019);
and U28376 (N_28376,N_23542,N_20950);
or U28377 (N_28377,N_21680,N_20306);
nand U28378 (N_28378,N_22661,N_22951);
nand U28379 (N_28379,N_21946,N_20381);
or U28380 (N_28380,N_23512,N_21189);
or U28381 (N_28381,N_22981,N_24683);
nand U28382 (N_28382,N_23253,N_22928);
nor U28383 (N_28383,N_22735,N_23264);
xnor U28384 (N_28384,N_21608,N_21833);
nand U28385 (N_28385,N_21401,N_21542);
or U28386 (N_28386,N_20871,N_22174);
nor U28387 (N_28387,N_22916,N_22988);
and U28388 (N_28388,N_22004,N_23063);
xor U28389 (N_28389,N_24948,N_23539);
and U28390 (N_28390,N_24424,N_20132);
nor U28391 (N_28391,N_22696,N_22683);
nand U28392 (N_28392,N_22335,N_20553);
nor U28393 (N_28393,N_22950,N_20119);
xor U28394 (N_28394,N_22382,N_23931);
and U28395 (N_28395,N_21226,N_24266);
or U28396 (N_28396,N_23162,N_20058);
nand U28397 (N_28397,N_20227,N_22591);
nor U28398 (N_28398,N_22950,N_21549);
or U28399 (N_28399,N_21298,N_24284);
or U28400 (N_28400,N_23609,N_24345);
xnor U28401 (N_28401,N_23428,N_23347);
and U28402 (N_28402,N_24005,N_21263);
or U28403 (N_28403,N_20601,N_23814);
xor U28404 (N_28404,N_21110,N_24209);
nor U28405 (N_28405,N_24790,N_24299);
and U28406 (N_28406,N_24292,N_24657);
nand U28407 (N_28407,N_24902,N_20618);
or U28408 (N_28408,N_24047,N_23756);
xnor U28409 (N_28409,N_23517,N_23494);
or U28410 (N_28410,N_23875,N_23216);
and U28411 (N_28411,N_23363,N_22967);
nand U28412 (N_28412,N_24717,N_23040);
and U28413 (N_28413,N_24103,N_20929);
xnor U28414 (N_28414,N_22987,N_20767);
nor U28415 (N_28415,N_24978,N_22641);
nand U28416 (N_28416,N_22011,N_23271);
xor U28417 (N_28417,N_21350,N_22461);
or U28418 (N_28418,N_21543,N_22408);
nor U28419 (N_28419,N_22283,N_21081);
and U28420 (N_28420,N_20866,N_21190);
or U28421 (N_28421,N_22423,N_21260);
or U28422 (N_28422,N_23370,N_24095);
xnor U28423 (N_28423,N_21981,N_21320);
nand U28424 (N_28424,N_20544,N_24603);
xnor U28425 (N_28425,N_22904,N_20182);
xnor U28426 (N_28426,N_22947,N_20382);
nor U28427 (N_28427,N_21819,N_23268);
or U28428 (N_28428,N_20854,N_20786);
and U28429 (N_28429,N_21285,N_20959);
or U28430 (N_28430,N_22562,N_23550);
and U28431 (N_28431,N_24153,N_22817);
or U28432 (N_28432,N_20406,N_20260);
nor U28433 (N_28433,N_21132,N_20976);
nand U28434 (N_28434,N_24115,N_23357);
nand U28435 (N_28435,N_21946,N_22211);
nand U28436 (N_28436,N_20553,N_23804);
xor U28437 (N_28437,N_23712,N_22804);
xor U28438 (N_28438,N_22362,N_23102);
and U28439 (N_28439,N_20101,N_24747);
nor U28440 (N_28440,N_23829,N_20995);
or U28441 (N_28441,N_23631,N_23390);
nand U28442 (N_28442,N_20611,N_23027);
nor U28443 (N_28443,N_20137,N_23075);
nor U28444 (N_28444,N_21558,N_21312);
xnor U28445 (N_28445,N_22847,N_24031);
or U28446 (N_28446,N_24357,N_21343);
or U28447 (N_28447,N_24127,N_22044);
xor U28448 (N_28448,N_23365,N_22459);
or U28449 (N_28449,N_21422,N_20653);
xnor U28450 (N_28450,N_24090,N_24282);
or U28451 (N_28451,N_20879,N_20108);
or U28452 (N_28452,N_22842,N_21499);
nor U28453 (N_28453,N_21838,N_24442);
or U28454 (N_28454,N_22189,N_20805);
nor U28455 (N_28455,N_23364,N_22098);
xor U28456 (N_28456,N_24734,N_24373);
nor U28457 (N_28457,N_22146,N_22027);
or U28458 (N_28458,N_24752,N_22803);
and U28459 (N_28459,N_22326,N_23328);
and U28460 (N_28460,N_21269,N_20362);
nor U28461 (N_28461,N_24708,N_21294);
nor U28462 (N_28462,N_21290,N_24292);
xor U28463 (N_28463,N_22172,N_21927);
or U28464 (N_28464,N_24539,N_20479);
nor U28465 (N_28465,N_23055,N_23357);
xnor U28466 (N_28466,N_22436,N_24265);
nand U28467 (N_28467,N_24347,N_22765);
nor U28468 (N_28468,N_23501,N_23719);
or U28469 (N_28469,N_24776,N_20929);
and U28470 (N_28470,N_22553,N_22583);
or U28471 (N_28471,N_20364,N_22476);
and U28472 (N_28472,N_22114,N_21495);
or U28473 (N_28473,N_23395,N_21350);
nand U28474 (N_28474,N_20988,N_24240);
and U28475 (N_28475,N_23983,N_21053);
nand U28476 (N_28476,N_23311,N_21815);
nor U28477 (N_28477,N_24507,N_22612);
nor U28478 (N_28478,N_22528,N_20000);
and U28479 (N_28479,N_23745,N_20701);
xnor U28480 (N_28480,N_21885,N_23477);
nand U28481 (N_28481,N_23433,N_22455);
nand U28482 (N_28482,N_20029,N_21596);
nor U28483 (N_28483,N_24862,N_23935);
nor U28484 (N_28484,N_21551,N_20487);
or U28485 (N_28485,N_21104,N_20441);
or U28486 (N_28486,N_20880,N_21601);
nor U28487 (N_28487,N_24175,N_23845);
xor U28488 (N_28488,N_22606,N_21403);
nand U28489 (N_28489,N_23171,N_23800);
and U28490 (N_28490,N_24566,N_21779);
and U28491 (N_28491,N_22692,N_21470);
and U28492 (N_28492,N_24018,N_21940);
nor U28493 (N_28493,N_22977,N_24672);
nor U28494 (N_28494,N_20045,N_23010);
and U28495 (N_28495,N_21317,N_20528);
and U28496 (N_28496,N_20385,N_20547);
and U28497 (N_28497,N_24110,N_24633);
or U28498 (N_28498,N_24808,N_23845);
and U28499 (N_28499,N_22118,N_24176);
nand U28500 (N_28500,N_22468,N_23665);
or U28501 (N_28501,N_23192,N_24952);
nor U28502 (N_28502,N_23073,N_22981);
or U28503 (N_28503,N_21152,N_20045);
nor U28504 (N_28504,N_20131,N_20433);
xnor U28505 (N_28505,N_22487,N_23981);
and U28506 (N_28506,N_24926,N_20211);
nor U28507 (N_28507,N_22953,N_23485);
or U28508 (N_28508,N_21051,N_23541);
and U28509 (N_28509,N_24349,N_23844);
and U28510 (N_28510,N_24538,N_22025);
nand U28511 (N_28511,N_21091,N_24470);
xor U28512 (N_28512,N_24346,N_24983);
nor U28513 (N_28513,N_21594,N_20100);
or U28514 (N_28514,N_21994,N_23935);
and U28515 (N_28515,N_23902,N_24551);
xnor U28516 (N_28516,N_23925,N_22649);
nand U28517 (N_28517,N_24119,N_21341);
and U28518 (N_28518,N_21833,N_20492);
or U28519 (N_28519,N_22332,N_22862);
nor U28520 (N_28520,N_24237,N_21439);
xor U28521 (N_28521,N_22672,N_20020);
or U28522 (N_28522,N_22718,N_22861);
xnor U28523 (N_28523,N_21023,N_23054);
or U28524 (N_28524,N_24236,N_20022);
and U28525 (N_28525,N_23264,N_21077);
xnor U28526 (N_28526,N_21850,N_22996);
or U28527 (N_28527,N_21750,N_24846);
nand U28528 (N_28528,N_22816,N_23283);
or U28529 (N_28529,N_24819,N_22316);
xor U28530 (N_28530,N_21779,N_22972);
nor U28531 (N_28531,N_21253,N_24729);
and U28532 (N_28532,N_22437,N_22076);
and U28533 (N_28533,N_20025,N_23242);
xor U28534 (N_28534,N_20095,N_20755);
nand U28535 (N_28535,N_20786,N_21641);
or U28536 (N_28536,N_21157,N_23404);
nor U28537 (N_28537,N_23009,N_21450);
nor U28538 (N_28538,N_23573,N_22705);
xnor U28539 (N_28539,N_20706,N_21636);
xor U28540 (N_28540,N_20507,N_21294);
or U28541 (N_28541,N_20247,N_23170);
or U28542 (N_28542,N_23901,N_22476);
and U28543 (N_28543,N_20292,N_21359);
and U28544 (N_28544,N_24226,N_22932);
xor U28545 (N_28545,N_23365,N_23859);
or U28546 (N_28546,N_23485,N_21177);
xnor U28547 (N_28547,N_22224,N_22085);
and U28548 (N_28548,N_23280,N_21616);
nand U28549 (N_28549,N_22059,N_21479);
nand U28550 (N_28550,N_24291,N_22698);
or U28551 (N_28551,N_22306,N_21174);
or U28552 (N_28552,N_24643,N_21299);
nor U28553 (N_28553,N_22767,N_23668);
xnor U28554 (N_28554,N_21251,N_21493);
and U28555 (N_28555,N_20991,N_21022);
nor U28556 (N_28556,N_22192,N_22749);
nand U28557 (N_28557,N_24320,N_21281);
xnor U28558 (N_28558,N_24715,N_21234);
and U28559 (N_28559,N_21201,N_21487);
nor U28560 (N_28560,N_22427,N_20145);
nor U28561 (N_28561,N_22162,N_23353);
and U28562 (N_28562,N_20682,N_20212);
and U28563 (N_28563,N_24016,N_22598);
xor U28564 (N_28564,N_21688,N_24026);
and U28565 (N_28565,N_20208,N_23681);
and U28566 (N_28566,N_23574,N_21191);
nand U28567 (N_28567,N_24258,N_24408);
xor U28568 (N_28568,N_23538,N_24352);
or U28569 (N_28569,N_24626,N_23975);
or U28570 (N_28570,N_23500,N_21385);
nand U28571 (N_28571,N_24707,N_24011);
nor U28572 (N_28572,N_22254,N_22652);
xnor U28573 (N_28573,N_23874,N_20800);
nand U28574 (N_28574,N_20068,N_22743);
nor U28575 (N_28575,N_24120,N_22116);
and U28576 (N_28576,N_22405,N_21021);
nor U28577 (N_28577,N_23179,N_23010);
xnor U28578 (N_28578,N_24490,N_24954);
and U28579 (N_28579,N_23266,N_23107);
or U28580 (N_28580,N_20443,N_20440);
xnor U28581 (N_28581,N_20339,N_20849);
nor U28582 (N_28582,N_21978,N_24172);
and U28583 (N_28583,N_22232,N_22074);
or U28584 (N_28584,N_20331,N_21972);
or U28585 (N_28585,N_23685,N_21954);
nand U28586 (N_28586,N_20532,N_24340);
or U28587 (N_28587,N_24248,N_21064);
nor U28588 (N_28588,N_24325,N_24655);
xnor U28589 (N_28589,N_24752,N_21894);
nor U28590 (N_28590,N_20144,N_22444);
nor U28591 (N_28591,N_23117,N_21535);
nor U28592 (N_28592,N_23419,N_24952);
xor U28593 (N_28593,N_20545,N_24400);
and U28594 (N_28594,N_22415,N_22314);
or U28595 (N_28595,N_22001,N_22498);
nand U28596 (N_28596,N_24319,N_22400);
or U28597 (N_28597,N_20426,N_20203);
or U28598 (N_28598,N_21130,N_24701);
or U28599 (N_28599,N_23811,N_22820);
xor U28600 (N_28600,N_21404,N_24694);
or U28601 (N_28601,N_24154,N_23293);
nand U28602 (N_28602,N_20984,N_20038);
nand U28603 (N_28603,N_24555,N_22946);
xnor U28604 (N_28604,N_20700,N_20557);
or U28605 (N_28605,N_20937,N_22192);
nand U28606 (N_28606,N_22523,N_22860);
nor U28607 (N_28607,N_21743,N_24151);
nand U28608 (N_28608,N_21908,N_23556);
nand U28609 (N_28609,N_22899,N_21961);
nand U28610 (N_28610,N_24702,N_23977);
nand U28611 (N_28611,N_23608,N_22062);
or U28612 (N_28612,N_24726,N_21501);
or U28613 (N_28613,N_24078,N_24502);
or U28614 (N_28614,N_23221,N_20248);
xnor U28615 (N_28615,N_21524,N_23555);
nand U28616 (N_28616,N_20854,N_22493);
xor U28617 (N_28617,N_22696,N_22326);
nand U28618 (N_28618,N_24785,N_20605);
xor U28619 (N_28619,N_21873,N_20405);
nor U28620 (N_28620,N_23675,N_21172);
xnor U28621 (N_28621,N_20215,N_24647);
nand U28622 (N_28622,N_24176,N_23843);
or U28623 (N_28623,N_24209,N_23102);
or U28624 (N_28624,N_24801,N_20440);
nand U28625 (N_28625,N_21893,N_23005);
or U28626 (N_28626,N_23765,N_22476);
xnor U28627 (N_28627,N_22336,N_20730);
xor U28628 (N_28628,N_20585,N_20667);
nor U28629 (N_28629,N_21613,N_24756);
and U28630 (N_28630,N_21456,N_21641);
nand U28631 (N_28631,N_21582,N_23750);
nor U28632 (N_28632,N_23944,N_24170);
or U28633 (N_28633,N_23958,N_24934);
xnor U28634 (N_28634,N_21429,N_24460);
or U28635 (N_28635,N_24239,N_20588);
nand U28636 (N_28636,N_20049,N_23505);
or U28637 (N_28637,N_20969,N_20510);
nand U28638 (N_28638,N_20600,N_24796);
nand U28639 (N_28639,N_23437,N_21485);
nand U28640 (N_28640,N_24461,N_20717);
nand U28641 (N_28641,N_20129,N_20592);
xor U28642 (N_28642,N_21939,N_24349);
nand U28643 (N_28643,N_24740,N_24690);
or U28644 (N_28644,N_20870,N_24066);
nor U28645 (N_28645,N_22902,N_22259);
and U28646 (N_28646,N_23039,N_21585);
nand U28647 (N_28647,N_21597,N_24761);
xor U28648 (N_28648,N_22258,N_20000);
or U28649 (N_28649,N_24183,N_23816);
and U28650 (N_28650,N_21771,N_22527);
xor U28651 (N_28651,N_24286,N_22124);
and U28652 (N_28652,N_23613,N_22431);
xnor U28653 (N_28653,N_22087,N_20060);
or U28654 (N_28654,N_22252,N_23767);
nand U28655 (N_28655,N_22338,N_24726);
and U28656 (N_28656,N_20755,N_21927);
nand U28657 (N_28657,N_20558,N_24417);
nor U28658 (N_28658,N_21715,N_24865);
or U28659 (N_28659,N_21825,N_24485);
nand U28660 (N_28660,N_24811,N_23651);
xnor U28661 (N_28661,N_21815,N_23466);
or U28662 (N_28662,N_20115,N_24342);
nor U28663 (N_28663,N_22491,N_22830);
nand U28664 (N_28664,N_23171,N_22433);
nand U28665 (N_28665,N_21406,N_23790);
nor U28666 (N_28666,N_21296,N_22230);
or U28667 (N_28667,N_20961,N_24797);
xnor U28668 (N_28668,N_24119,N_21959);
nand U28669 (N_28669,N_22090,N_24435);
and U28670 (N_28670,N_22346,N_20760);
or U28671 (N_28671,N_20204,N_21959);
nand U28672 (N_28672,N_22936,N_21105);
nand U28673 (N_28673,N_20948,N_23979);
xor U28674 (N_28674,N_22250,N_21306);
nand U28675 (N_28675,N_23115,N_20783);
and U28676 (N_28676,N_24801,N_23382);
or U28677 (N_28677,N_22666,N_24801);
nor U28678 (N_28678,N_21453,N_20681);
nor U28679 (N_28679,N_20189,N_20765);
or U28680 (N_28680,N_22813,N_22143);
and U28681 (N_28681,N_23930,N_22580);
and U28682 (N_28682,N_24614,N_24073);
xnor U28683 (N_28683,N_20579,N_20996);
xor U28684 (N_28684,N_21318,N_22852);
xor U28685 (N_28685,N_24670,N_20270);
xor U28686 (N_28686,N_22932,N_21014);
and U28687 (N_28687,N_21810,N_21435);
or U28688 (N_28688,N_23538,N_23054);
xnor U28689 (N_28689,N_22967,N_20842);
nand U28690 (N_28690,N_20989,N_23389);
or U28691 (N_28691,N_24518,N_21155);
and U28692 (N_28692,N_20035,N_22803);
and U28693 (N_28693,N_22141,N_23036);
xor U28694 (N_28694,N_21457,N_23947);
and U28695 (N_28695,N_21190,N_21167);
nand U28696 (N_28696,N_21373,N_23961);
nor U28697 (N_28697,N_24169,N_21265);
nor U28698 (N_28698,N_23952,N_20694);
xnor U28699 (N_28699,N_23744,N_23804);
or U28700 (N_28700,N_21076,N_23412);
nor U28701 (N_28701,N_23581,N_23955);
or U28702 (N_28702,N_22000,N_22570);
and U28703 (N_28703,N_24729,N_23384);
nor U28704 (N_28704,N_22919,N_23923);
nor U28705 (N_28705,N_20177,N_23188);
nand U28706 (N_28706,N_23394,N_24830);
xnor U28707 (N_28707,N_20218,N_22587);
and U28708 (N_28708,N_22310,N_22371);
xor U28709 (N_28709,N_20982,N_22361);
nand U28710 (N_28710,N_23527,N_22206);
nor U28711 (N_28711,N_20218,N_22888);
xor U28712 (N_28712,N_23547,N_23173);
or U28713 (N_28713,N_20455,N_20682);
and U28714 (N_28714,N_22226,N_23635);
nor U28715 (N_28715,N_24046,N_20968);
xnor U28716 (N_28716,N_23298,N_20221);
xor U28717 (N_28717,N_21171,N_20233);
nor U28718 (N_28718,N_24466,N_22850);
and U28719 (N_28719,N_23953,N_20026);
xor U28720 (N_28720,N_20758,N_22440);
nor U28721 (N_28721,N_21253,N_20286);
or U28722 (N_28722,N_20945,N_22731);
nand U28723 (N_28723,N_22751,N_24430);
or U28724 (N_28724,N_20207,N_23178);
nand U28725 (N_28725,N_21438,N_23405);
or U28726 (N_28726,N_20566,N_21195);
or U28727 (N_28727,N_22894,N_24750);
nor U28728 (N_28728,N_20773,N_24900);
or U28729 (N_28729,N_21816,N_23818);
nand U28730 (N_28730,N_21546,N_21059);
nor U28731 (N_28731,N_20618,N_20579);
or U28732 (N_28732,N_22340,N_21377);
nand U28733 (N_28733,N_21877,N_21091);
and U28734 (N_28734,N_20048,N_22743);
xnor U28735 (N_28735,N_20160,N_23729);
xor U28736 (N_28736,N_24091,N_21623);
and U28737 (N_28737,N_21600,N_21052);
nand U28738 (N_28738,N_22010,N_21094);
and U28739 (N_28739,N_20335,N_23008);
xnor U28740 (N_28740,N_21921,N_24388);
nor U28741 (N_28741,N_24290,N_24454);
xnor U28742 (N_28742,N_21909,N_23241);
nor U28743 (N_28743,N_22984,N_22125);
nand U28744 (N_28744,N_23732,N_20003);
or U28745 (N_28745,N_22664,N_21611);
nor U28746 (N_28746,N_20237,N_20132);
nand U28747 (N_28747,N_20173,N_24273);
nor U28748 (N_28748,N_24432,N_21138);
nor U28749 (N_28749,N_24308,N_21774);
or U28750 (N_28750,N_21651,N_20774);
xor U28751 (N_28751,N_24758,N_23765);
and U28752 (N_28752,N_23712,N_22375);
xor U28753 (N_28753,N_24112,N_24931);
nand U28754 (N_28754,N_22352,N_20378);
and U28755 (N_28755,N_23162,N_21128);
xor U28756 (N_28756,N_21185,N_24278);
nor U28757 (N_28757,N_20367,N_23935);
or U28758 (N_28758,N_24420,N_21269);
and U28759 (N_28759,N_20923,N_23264);
xnor U28760 (N_28760,N_24641,N_24084);
nor U28761 (N_28761,N_23994,N_24542);
or U28762 (N_28762,N_24485,N_22620);
nand U28763 (N_28763,N_24579,N_20304);
nor U28764 (N_28764,N_22918,N_20213);
xnor U28765 (N_28765,N_24412,N_21120);
and U28766 (N_28766,N_20976,N_21579);
and U28767 (N_28767,N_22657,N_20945);
and U28768 (N_28768,N_23540,N_22104);
nand U28769 (N_28769,N_20255,N_21691);
nor U28770 (N_28770,N_20197,N_22001);
nand U28771 (N_28771,N_23869,N_21906);
xnor U28772 (N_28772,N_20951,N_21169);
or U28773 (N_28773,N_24240,N_20244);
nand U28774 (N_28774,N_21246,N_20219);
xnor U28775 (N_28775,N_23817,N_24176);
xor U28776 (N_28776,N_22854,N_22619);
nand U28777 (N_28777,N_23770,N_22847);
nand U28778 (N_28778,N_21816,N_20072);
nor U28779 (N_28779,N_21354,N_24417);
nor U28780 (N_28780,N_21319,N_20785);
xor U28781 (N_28781,N_23874,N_21830);
or U28782 (N_28782,N_22861,N_22085);
or U28783 (N_28783,N_21117,N_20350);
xor U28784 (N_28784,N_20229,N_21026);
xnor U28785 (N_28785,N_23052,N_20711);
or U28786 (N_28786,N_24114,N_24090);
nand U28787 (N_28787,N_23599,N_23007);
nand U28788 (N_28788,N_23610,N_24755);
or U28789 (N_28789,N_22526,N_23003);
nor U28790 (N_28790,N_23730,N_23455);
nand U28791 (N_28791,N_21689,N_20010);
or U28792 (N_28792,N_22070,N_24154);
nor U28793 (N_28793,N_24745,N_24209);
nand U28794 (N_28794,N_23739,N_24348);
or U28795 (N_28795,N_23286,N_22491);
and U28796 (N_28796,N_22841,N_21188);
or U28797 (N_28797,N_23545,N_20608);
nand U28798 (N_28798,N_23751,N_22836);
nand U28799 (N_28799,N_20934,N_22181);
and U28800 (N_28800,N_23103,N_20701);
or U28801 (N_28801,N_21641,N_20398);
and U28802 (N_28802,N_23308,N_20600);
xnor U28803 (N_28803,N_20694,N_22611);
or U28804 (N_28804,N_21020,N_23805);
or U28805 (N_28805,N_20585,N_21525);
nor U28806 (N_28806,N_22102,N_22481);
xnor U28807 (N_28807,N_22326,N_21581);
and U28808 (N_28808,N_21249,N_23240);
and U28809 (N_28809,N_21224,N_22142);
or U28810 (N_28810,N_23713,N_21380);
or U28811 (N_28811,N_21413,N_23394);
or U28812 (N_28812,N_24074,N_24813);
nor U28813 (N_28813,N_21396,N_24677);
or U28814 (N_28814,N_22198,N_23647);
nand U28815 (N_28815,N_24909,N_20010);
or U28816 (N_28816,N_24760,N_20314);
nor U28817 (N_28817,N_21140,N_23060);
and U28818 (N_28818,N_24453,N_20809);
nor U28819 (N_28819,N_23809,N_24856);
nor U28820 (N_28820,N_22646,N_21374);
nor U28821 (N_28821,N_22928,N_20629);
and U28822 (N_28822,N_21727,N_23290);
or U28823 (N_28823,N_22966,N_22542);
and U28824 (N_28824,N_20667,N_22410);
and U28825 (N_28825,N_23503,N_22494);
xnor U28826 (N_28826,N_24985,N_21926);
nand U28827 (N_28827,N_21286,N_24014);
nand U28828 (N_28828,N_23413,N_23722);
and U28829 (N_28829,N_22199,N_24993);
and U28830 (N_28830,N_24373,N_22150);
or U28831 (N_28831,N_23906,N_22795);
nand U28832 (N_28832,N_20808,N_21175);
nand U28833 (N_28833,N_21712,N_24366);
nand U28834 (N_28834,N_23635,N_21254);
xor U28835 (N_28835,N_21073,N_20820);
nand U28836 (N_28836,N_23887,N_24078);
xnor U28837 (N_28837,N_21173,N_24575);
and U28838 (N_28838,N_23495,N_22206);
nor U28839 (N_28839,N_23761,N_20169);
and U28840 (N_28840,N_24071,N_20741);
and U28841 (N_28841,N_22162,N_20722);
and U28842 (N_28842,N_23770,N_21406);
xnor U28843 (N_28843,N_21741,N_22701);
xor U28844 (N_28844,N_20103,N_21935);
nand U28845 (N_28845,N_24557,N_20023);
nor U28846 (N_28846,N_20318,N_24481);
or U28847 (N_28847,N_21389,N_24438);
or U28848 (N_28848,N_21349,N_24690);
or U28849 (N_28849,N_21125,N_22980);
nand U28850 (N_28850,N_22903,N_24297);
or U28851 (N_28851,N_22703,N_20990);
and U28852 (N_28852,N_23773,N_23671);
nand U28853 (N_28853,N_23208,N_22214);
or U28854 (N_28854,N_22290,N_24338);
or U28855 (N_28855,N_23262,N_22185);
xnor U28856 (N_28856,N_24581,N_24541);
nand U28857 (N_28857,N_23896,N_21402);
or U28858 (N_28858,N_20168,N_22446);
nor U28859 (N_28859,N_21954,N_22598);
or U28860 (N_28860,N_21771,N_23790);
and U28861 (N_28861,N_21425,N_23318);
or U28862 (N_28862,N_24117,N_21716);
and U28863 (N_28863,N_22987,N_21975);
xnor U28864 (N_28864,N_21006,N_20482);
or U28865 (N_28865,N_21206,N_23503);
or U28866 (N_28866,N_21719,N_24284);
or U28867 (N_28867,N_24915,N_21605);
nor U28868 (N_28868,N_22897,N_20282);
nor U28869 (N_28869,N_20636,N_24341);
nor U28870 (N_28870,N_22177,N_22137);
xor U28871 (N_28871,N_23792,N_20261);
nand U28872 (N_28872,N_21252,N_24569);
xnor U28873 (N_28873,N_21051,N_23575);
or U28874 (N_28874,N_20972,N_20409);
xor U28875 (N_28875,N_22967,N_20832);
and U28876 (N_28876,N_21282,N_23558);
nand U28877 (N_28877,N_24781,N_20596);
nand U28878 (N_28878,N_23653,N_22624);
or U28879 (N_28879,N_24079,N_23153);
or U28880 (N_28880,N_21655,N_23706);
nor U28881 (N_28881,N_24200,N_22358);
nand U28882 (N_28882,N_23309,N_24288);
nor U28883 (N_28883,N_20782,N_21496);
and U28884 (N_28884,N_21359,N_22589);
nand U28885 (N_28885,N_24812,N_20838);
xnor U28886 (N_28886,N_24321,N_22167);
or U28887 (N_28887,N_24807,N_24863);
and U28888 (N_28888,N_23360,N_20437);
or U28889 (N_28889,N_21512,N_20305);
and U28890 (N_28890,N_22819,N_24127);
nor U28891 (N_28891,N_24725,N_20624);
nand U28892 (N_28892,N_22454,N_24738);
and U28893 (N_28893,N_22326,N_23803);
or U28894 (N_28894,N_22554,N_20485);
or U28895 (N_28895,N_24780,N_22303);
or U28896 (N_28896,N_21749,N_21226);
or U28897 (N_28897,N_23994,N_21558);
or U28898 (N_28898,N_23657,N_23762);
nor U28899 (N_28899,N_23879,N_20589);
or U28900 (N_28900,N_23736,N_21391);
and U28901 (N_28901,N_22028,N_23149);
and U28902 (N_28902,N_22778,N_22183);
and U28903 (N_28903,N_24363,N_20851);
nor U28904 (N_28904,N_24498,N_23002);
nand U28905 (N_28905,N_21302,N_22537);
xnor U28906 (N_28906,N_22027,N_21661);
xnor U28907 (N_28907,N_23162,N_22497);
and U28908 (N_28908,N_21185,N_20249);
nand U28909 (N_28909,N_21443,N_22536);
nor U28910 (N_28910,N_24921,N_22852);
or U28911 (N_28911,N_24676,N_22131);
nand U28912 (N_28912,N_21992,N_22215);
nor U28913 (N_28913,N_21024,N_20332);
and U28914 (N_28914,N_21328,N_23353);
nor U28915 (N_28915,N_23252,N_23169);
or U28916 (N_28916,N_20451,N_20147);
nor U28917 (N_28917,N_22679,N_24215);
xnor U28918 (N_28918,N_22131,N_23496);
and U28919 (N_28919,N_23547,N_20275);
nor U28920 (N_28920,N_21941,N_21417);
nand U28921 (N_28921,N_21418,N_22751);
or U28922 (N_28922,N_23895,N_21356);
or U28923 (N_28923,N_23926,N_23185);
xor U28924 (N_28924,N_23674,N_24030);
or U28925 (N_28925,N_22593,N_22264);
nor U28926 (N_28926,N_22083,N_22969);
and U28927 (N_28927,N_23198,N_20356);
nor U28928 (N_28928,N_23572,N_22643);
nand U28929 (N_28929,N_23040,N_20934);
nor U28930 (N_28930,N_23900,N_23054);
nand U28931 (N_28931,N_20040,N_22340);
and U28932 (N_28932,N_22022,N_20940);
and U28933 (N_28933,N_24070,N_20204);
xor U28934 (N_28934,N_21426,N_20407);
or U28935 (N_28935,N_22473,N_20509);
xnor U28936 (N_28936,N_21607,N_22766);
or U28937 (N_28937,N_23335,N_21375);
nor U28938 (N_28938,N_22188,N_23945);
nand U28939 (N_28939,N_23384,N_22957);
or U28940 (N_28940,N_21364,N_23134);
xnor U28941 (N_28941,N_23040,N_21548);
or U28942 (N_28942,N_21054,N_24794);
and U28943 (N_28943,N_21169,N_21712);
or U28944 (N_28944,N_24585,N_24920);
nand U28945 (N_28945,N_24880,N_20179);
nor U28946 (N_28946,N_23043,N_24520);
or U28947 (N_28947,N_24826,N_24291);
and U28948 (N_28948,N_23797,N_22263);
and U28949 (N_28949,N_22711,N_20020);
xor U28950 (N_28950,N_22295,N_24157);
nor U28951 (N_28951,N_22108,N_23383);
or U28952 (N_28952,N_22564,N_20928);
and U28953 (N_28953,N_22483,N_23746);
and U28954 (N_28954,N_22098,N_22967);
xnor U28955 (N_28955,N_23092,N_20880);
nand U28956 (N_28956,N_23321,N_23808);
or U28957 (N_28957,N_21590,N_20652);
nand U28958 (N_28958,N_22572,N_22797);
nor U28959 (N_28959,N_20855,N_24383);
nor U28960 (N_28960,N_24186,N_20696);
xor U28961 (N_28961,N_24074,N_23393);
xor U28962 (N_28962,N_21031,N_20041);
or U28963 (N_28963,N_22845,N_21009);
and U28964 (N_28964,N_22084,N_22094);
nand U28965 (N_28965,N_24691,N_22568);
or U28966 (N_28966,N_20654,N_23503);
nor U28967 (N_28967,N_22553,N_24944);
or U28968 (N_28968,N_23189,N_21418);
xor U28969 (N_28969,N_20361,N_24009);
xor U28970 (N_28970,N_21171,N_20340);
or U28971 (N_28971,N_22199,N_20928);
nor U28972 (N_28972,N_24846,N_21576);
or U28973 (N_28973,N_23674,N_22080);
and U28974 (N_28974,N_22829,N_20264);
and U28975 (N_28975,N_22902,N_24754);
nand U28976 (N_28976,N_23729,N_20563);
or U28977 (N_28977,N_20829,N_22631);
xnor U28978 (N_28978,N_20023,N_22630);
nand U28979 (N_28979,N_20768,N_22535);
nand U28980 (N_28980,N_21843,N_20635);
nor U28981 (N_28981,N_20301,N_22441);
xor U28982 (N_28982,N_20348,N_21883);
nand U28983 (N_28983,N_22827,N_21052);
and U28984 (N_28984,N_22622,N_21141);
or U28985 (N_28985,N_24101,N_23496);
nand U28986 (N_28986,N_22598,N_23485);
and U28987 (N_28987,N_23141,N_22247);
and U28988 (N_28988,N_22057,N_21919);
or U28989 (N_28989,N_21545,N_21983);
xnor U28990 (N_28990,N_24360,N_24346);
nand U28991 (N_28991,N_22630,N_22444);
xor U28992 (N_28992,N_20746,N_24151);
nor U28993 (N_28993,N_24029,N_24057);
or U28994 (N_28994,N_23541,N_22128);
xor U28995 (N_28995,N_23116,N_20245);
nand U28996 (N_28996,N_24228,N_20730);
xnor U28997 (N_28997,N_23482,N_20468);
xor U28998 (N_28998,N_20462,N_20754);
xnor U28999 (N_28999,N_20978,N_23004);
and U29000 (N_29000,N_24141,N_21675);
and U29001 (N_29001,N_24182,N_23523);
and U29002 (N_29002,N_24031,N_23724);
nor U29003 (N_29003,N_20637,N_21007);
and U29004 (N_29004,N_20033,N_21507);
nand U29005 (N_29005,N_22930,N_20183);
xor U29006 (N_29006,N_24069,N_22552);
and U29007 (N_29007,N_23933,N_21473);
or U29008 (N_29008,N_22093,N_21945);
nor U29009 (N_29009,N_21049,N_20998);
xnor U29010 (N_29010,N_21675,N_20790);
xnor U29011 (N_29011,N_24219,N_22547);
and U29012 (N_29012,N_22588,N_23274);
and U29013 (N_29013,N_23742,N_21166);
nand U29014 (N_29014,N_20929,N_22691);
nand U29015 (N_29015,N_23661,N_20839);
nor U29016 (N_29016,N_20598,N_21459);
nor U29017 (N_29017,N_24863,N_22780);
or U29018 (N_29018,N_24598,N_20725);
nand U29019 (N_29019,N_23773,N_20944);
nor U29020 (N_29020,N_22149,N_23713);
nor U29021 (N_29021,N_20676,N_24820);
or U29022 (N_29022,N_23028,N_24990);
xnor U29023 (N_29023,N_23305,N_23749);
nor U29024 (N_29024,N_24799,N_24929);
xor U29025 (N_29025,N_20125,N_24339);
or U29026 (N_29026,N_24191,N_22412);
nor U29027 (N_29027,N_21671,N_24317);
xor U29028 (N_29028,N_24466,N_23809);
or U29029 (N_29029,N_21623,N_21531);
xor U29030 (N_29030,N_24879,N_23621);
or U29031 (N_29031,N_20510,N_20344);
xnor U29032 (N_29032,N_24292,N_23904);
and U29033 (N_29033,N_22387,N_20896);
nand U29034 (N_29034,N_21196,N_24030);
and U29035 (N_29035,N_20798,N_21456);
nor U29036 (N_29036,N_24480,N_20615);
or U29037 (N_29037,N_20140,N_24001);
nor U29038 (N_29038,N_23441,N_21306);
and U29039 (N_29039,N_21504,N_23686);
xor U29040 (N_29040,N_24613,N_21531);
and U29041 (N_29041,N_20358,N_24061);
nand U29042 (N_29042,N_24712,N_20310);
xor U29043 (N_29043,N_20863,N_22115);
and U29044 (N_29044,N_23175,N_21667);
or U29045 (N_29045,N_20379,N_23703);
or U29046 (N_29046,N_21568,N_22416);
xor U29047 (N_29047,N_20717,N_20651);
or U29048 (N_29048,N_21092,N_23796);
and U29049 (N_29049,N_21239,N_21744);
nor U29050 (N_29050,N_23518,N_22291);
xnor U29051 (N_29051,N_23937,N_24568);
nand U29052 (N_29052,N_21006,N_22206);
or U29053 (N_29053,N_24830,N_24883);
nand U29054 (N_29054,N_20863,N_24271);
xnor U29055 (N_29055,N_23305,N_20082);
xor U29056 (N_29056,N_20898,N_24122);
xor U29057 (N_29057,N_23204,N_20387);
and U29058 (N_29058,N_22791,N_22702);
or U29059 (N_29059,N_22387,N_21138);
or U29060 (N_29060,N_21055,N_20092);
or U29061 (N_29061,N_22893,N_20661);
and U29062 (N_29062,N_21325,N_24530);
nand U29063 (N_29063,N_22297,N_22161);
xor U29064 (N_29064,N_22508,N_23281);
and U29065 (N_29065,N_24226,N_24720);
and U29066 (N_29066,N_20742,N_21454);
and U29067 (N_29067,N_21900,N_21919);
and U29068 (N_29068,N_21622,N_24209);
nand U29069 (N_29069,N_21798,N_24300);
nand U29070 (N_29070,N_23306,N_23704);
or U29071 (N_29071,N_24270,N_21767);
or U29072 (N_29072,N_20109,N_23929);
xnor U29073 (N_29073,N_24849,N_23702);
xnor U29074 (N_29074,N_21844,N_24568);
nand U29075 (N_29075,N_20565,N_24167);
xnor U29076 (N_29076,N_24336,N_22925);
or U29077 (N_29077,N_23063,N_22464);
and U29078 (N_29078,N_22358,N_20314);
nand U29079 (N_29079,N_21628,N_24258);
xor U29080 (N_29080,N_20282,N_21332);
or U29081 (N_29081,N_24430,N_22680);
xnor U29082 (N_29082,N_21396,N_22282);
and U29083 (N_29083,N_24015,N_24585);
nor U29084 (N_29084,N_23167,N_20607);
and U29085 (N_29085,N_24859,N_21069);
xor U29086 (N_29086,N_21383,N_22464);
nand U29087 (N_29087,N_23355,N_21490);
xor U29088 (N_29088,N_20908,N_20413);
and U29089 (N_29089,N_23335,N_23720);
or U29090 (N_29090,N_24032,N_20907);
nand U29091 (N_29091,N_24038,N_21693);
and U29092 (N_29092,N_20784,N_23282);
nor U29093 (N_29093,N_23151,N_22719);
nand U29094 (N_29094,N_22519,N_24180);
and U29095 (N_29095,N_21705,N_20811);
nor U29096 (N_29096,N_21306,N_21880);
or U29097 (N_29097,N_20145,N_24308);
or U29098 (N_29098,N_23318,N_21543);
nand U29099 (N_29099,N_22094,N_21101);
and U29100 (N_29100,N_24380,N_21767);
or U29101 (N_29101,N_21979,N_21379);
nand U29102 (N_29102,N_21994,N_21896);
nor U29103 (N_29103,N_24913,N_20779);
nor U29104 (N_29104,N_23377,N_21560);
nor U29105 (N_29105,N_23585,N_24376);
xor U29106 (N_29106,N_24682,N_24948);
nand U29107 (N_29107,N_24576,N_24515);
xor U29108 (N_29108,N_23911,N_21245);
or U29109 (N_29109,N_22303,N_21895);
xor U29110 (N_29110,N_23995,N_23145);
nor U29111 (N_29111,N_21954,N_24812);
or U29112 (N_29112,N_22673,N_22727);
xnor U29113 (N_29113,N_23878,N_21560);
nor U29114 (N_29114,N_20645,N_21947);
nand U29115 (N_29115,N_23169,N_24982);
nor U29116 (N_29116,N_24971,N_21493);
nor U29117 (N_29117,N_20365,N_24267);
xnor U29118 (N_29118,N_24655,N_22443);
nor U29119 (N_29119,N_23369,N_21149);
nor U29120 (N_29120,N_22963,N_23195);
nor U29121 (N_29121,N_20613,N_20436);
and U29122 (N_29122,N_20468,N_21348);
nor U29123 (N_29123,N_23163,N_24156);
nand U29124 (N_29124,N_20988,N_20326);
nor U29125 (N_29125,N_20198,N_21475);
or U29126 (N_29126,N_24041,N_24210);
nor U29127 (N_29127,N_22055,N_24469);
and U29128 (N_29128,N_20548,N_21650);
xnor U29129 (N_29129,N_20362,N_22537);
or U29130 (N_29130,N_22445,N_22127);
or U29131 (N_29131,N_23212,N_20501);
or U29132 (N_29132,N_23204,N_21944);
nand U29133 (N_29133,N_22519,N_24218);
nand U29134 (N_29134,N_21586,N_22904);
or U29135 (N_29135,N_20681,N_21290);
xnor U29136 (N_29136,N_20893,N_20372);
and U29137 (N_29137,N_23521,N_20807);
and U29138 (N_29138,N_24554,N_20924);
and U29139 (N_29139,N_20436,N_21107);
nand U29140 (N_29140,N_21687,N_21294);
nor U29141 (N_29141,N_23361,N_24735);
nand U29142 (N_29142,N_23088,N_23690);
nand U29143 (N_29143,N_22878,N_22481);
or U29144 (N_29144,N_20739,N_23983);
xnor U29145 (N_29145,N_21720,N_21840);
nor U29146 (N_29146,N_22608,N_23255);
and U29147 (N_29147,N_20022,N_24674);
nand U29148 (N_29148,N_20451,N_22676);
nand U29149 (N_29149,N_24629,N_22435);
and U29150 (N_29150,N_22155,N_23516);
and U29151 (N_29151,N_24481,N_22868);
nor U29152 (N_29152,N_24979,N_24724);
nand U29153 (N_29153,N_22296,N_22571);
or U29154 (N_29154,N_22922,N_22926);
nor U29155 (N_29155,N_22738,N_20701);
xnor U29156 (N_29156,N_21105,N_20520);
or U29157 (N_29157,N_21835,N_24829);
or U29158 (N_29158,N_21215,N_23080);
nor U29159 (N_29159,N_22154,N_23293);
nor U29160 (N_29160,N_24947,N_23647);
nor U29161 (N_29161,N_21940,N_23906);
nor U29162 (N_29162,N_22034,N_22077);
nor U29163 (N_29163,N_24228,N_21331);
xor U29164 (N_29164,N_20533,N_22590);
and U29165 (N_29165,N_24104,N_20048);
nor U29166 (N_29166,N_22781,N_24230);
or U29167 (N_29167,N_23572,N_24386);
nand U29168 (N_29168,N_23461,N_20432);
nor U29169 (N_29169,N_22042,N_20230);
nand U29170 (N_29170,N_22411,N_20188);
and U29171 (N_29171,N_21690,N_23817);
nand U29172 (N_29172,N_21013,N_22849);
or U29173 (N_29173,N_20467,N_22288);
or U29174 (N_29174,N_22847,N_20467);
and U29175 (N_29175,N_21998,N_22635);
nand U29176 (N_29176,N_24607,N_21145);
xnor U29177 (N_29177,N_22113,N_21985);
and U29178 (N_29178,N_23728,N_20536);
nor U29179 (N_29179,N_23388,N_22817);
nor U29180 (N_29180,N_22179,N_24347);
nor U29181 (N_29181,N_21544,N_22586);
nand U29182 (N_29182,N_23064,N_22580);
and U29183 (N_29183,N_22224,N_24176);
and U29184 (N_29184,N_23333,N_20625);
nor U29185 (N_29185,N_21133,N_22304);
or U29186 (N_29186,N_21131,N_23590);
xor U29187 (N_29187,N_20867,N_20934);
and U29188 (N_29188,N_23746,N_24687);
and U29189 (N_29189,N_21725,N_23777);
or U29190 (N_29190,N_20524,N_23173);
nor U29191 (N_29191,N_21750,N_24672);
xnor U29192 (N_29192,N_23950,N_23594);
or U29193 (N_29193,N_20197,N_22369);
xor U29194 (N_29194,N_23333,N_24679);
xnor U29195 (N_29195,N_21941,N_20578);
nor U29196 (N_29196,N_22670,N_24525);
nand U29197 (N_29197,N_23302,N_22214);
and U29198 (N_29198,N_23219,N_21280);
nand U29199 (N_29199,N_21474,N_23001);
nor U29200 (N_29200,N_21211,N_21296);
nand U29201 (N_29201,N_23418,N_21157);
xor U29202 (N_29202,N_23222,N_23515);
nand U29203 (N_29203,N_20119,N_22643);
and U29204 (N_29204,N_20904,N_22549);
or U29205 (N_29205,N_24798,N_20828);
nand U29206 (N_29206,N_22490,N_21089);
and U29207 (N_29207,N_23110,N_21475);
xnor U29208 (N_29208,N_23529,N_24885);
nor U29209 (N_29209,N_24521,N_22333);
nand U29210 (N_29210,N_20179,N_23146);
and U29211 (N_29211,N_22825,N_20851);
nand U29212 (N_29212,N_23629,N_23294);
nor U29213 (N_29213,N_20662,N_23994);
nand U29214 (N_29214,N_23397,N_22270);
nor U29215 (N_29215,N_23211,N_21784);
and U29216 (N_29216,N_20666,N_20554);
or U29217 (N_29217,N_20118,N_23880);
or U29218 (N_29218,N_20311,N_20878);
and U29219 (N_29219,N_23515,N_20938);
or U29220 (N_29220,N_24596,N_21661);
nor U29221 (N_29221,N_23015,N_23262);
and U29222 (N_29222,N_21863,N_24639);
and U29223 (N_29223,N_20130,N_20136);
xor U29224 (N_29224,N_24086,N_22945);
nand U29225 (N_29225,N_22779,N_20104);
and U29226 (N_29226,N_20854,N_23895);
and U29227 (N_29227,N_20952,N_23390);
nand U29228 (N_29228,N_24743,N_21262);
or U29229 (N_29229,N_22928,N_21010);
and U29230 (N_29230,N_20118,N_21250);
or U29231 (N_29231,N_22302,N_21294);
nand U29232 (N_29232,N_24408,N_20799);
nor U29233 (N_29233,N_20243,N_22971);
nor U29234 (N_29234,N_24809,N_20321);
and U29235 (N_29235,N_23088,N_23532);
and U29236 (N_29236,N_23321,N_22556);
nor U29237 (N_29237,N_22936,N_23215);
and U29238 (N_29238,N_24826,N_20621);
nand U29239 (N_29239,N_20348,N_24724);
xor U29240 (N_29240,N_21409,N_22520);
nor U29241 (N_29241,N_23792,N_20720);
nor U29242 (N_29242,N_23499,N_24271);
or U29243 (N_29243,N_24891,N_23005);
nor U29244 (N_29244,N_24180,N_21426);
xnor U29245 (N_29245,N_24683,N_20818);
xor U29246 (N_29246,N_22436,N_24484);
nand U29247 (N_29247,N_22311,N_24440);
nor U29248 (N_29248,N_20965,N_23537);
or U29249 (N_29249,N_22897,N_21465);
and U29250 (N_29250,N_22354,N_20191);
nand U29251 (N_29251,N_24739,N_23998);
xnor U29252 (N_29252,N_20092,N_20852);
and U29253 (N_29253,N_24133,N_20033);
xor U29254 (N_29254,N_24944,N_20549);
and U29255 (N_29255,N_23449,N_20305);
nor U29256 (N_29256,N_24418,N_20989);
or U29257 (N_29257,N_23677,N_22832);
and U29258 (N_29258,N_20481,N_24680);
nor U29259 (N_29259,N_24916,N_23966);
and U29260 (N_29260,N_24679,N_20042);
nand U29261 (N_29261,N_24679,N_23987);
xor U29262 (N_29262,N_24496,N_20627);
and U29263 (N_29263,N_23429,N_20201);
nand U29264 (N_29264,N_20217,N_22668);
nor U29265 (N_29265,N_23816,N_20420);
and U29266 (N_29266,N_24104,N_21015);
or U29267 (N_29267,N_23439,N_20420);
or U29268 (N_29268,N_23072,N_22818);
nor U29269 (N_29269,N_22289,N_24681);
or U29270 (N_29270,N_22257,N_24892);
and U29271 (N_29271,N_24790,N_21382);
nor U29272 (N_29272,N_24723,N_20782);
or U29273 (N_29273,N_23711,N_20511);
and U29274 (N_29274,N_23686,N_24988);
xor U29275 (N_29275,N_21198,N_21239);
or U29276 (N_29276,N_24333,N_22016);
or U29277 (N_29277,N_22532,N_22260);
and U29278 (N_29278,N_20250,N_23346);
nor U29279 (N_29279,N_24514,N_23941);
or U29280 (N_29280,N_23543,N_22960);
nand U29281 (N_29281,N_20578,N_21410);
nand U29282 (N_29282,N_24345,N_24841);
nand U29283 (N_29283,N_24072,N_20488);
xnor U29284 (N_29284,N_22703,N_23620);
and U29285 (N_29285,N_20357,N_24361);
nor U29286 (N_29286,N_24818,N_23952);
or U29287 (N_29287,N_22872,N_24345);
nand U29288 (N_29288,N_24610,N_23220);
or U29289 (N_29289,N_22050,N_21718);
nor U29290 (N_29290,N_21787,N_22354);
or U29291 (N_29291,N_24793,N_20419);
and U29292 (N_29292,N_22163,N_24250);
or U29293 (N_29293,N_23341,N_23412);
nor U29294 (N_29294,N_21536,N_24177);
and U29295 (N_29295,N_20400,N_23433);
and U29296 (N_29296,N_20333,N_24547);
and U29297 (N_29297,N_22964,N_21213);
nor U29298 (N_29298,N_22821,N_24322);
or U29299 (N_29299,N_20413,N_23636);
nor U29300 (N_29300,N_22347,N_22659);
or U29301 (N_29301,N_23781,N_22842);
and U29302 (N_29302,N_24918,N_20792);
nand U29303 (N_29303,N_20431,N_22033);
or U29304 (N_29304,N_20194,N_23993);
xor U29305 (N_29305,N_24865,N_20690);
xor U29306 (N_29306,N_23875,N_20992);
nor U29307 (N_29307,N_20318,N_21149);
and U29308 (N_29308,N_24691,N_24951);
xnor U29309 (N_29309,N_24228,N_24818);
or U29310 (N_29310,N_21554,N_21504);
xor U29311 (N_29311,N_24108,N_24403);
or U29312 (N_29312,N_24815,N_23156);
and U29313 (N_29313,N_20883,N_24004);
nand U29314 (N_29314,N_23267,N_20925);
xnor U29315 (N_29315,N_22649,N_21405);
and U29316 (N_29316,N_24679,N_23557);
nor U29317 (N_29317,N_24510,N_23832);
or U29318 (N_29318,N_24599,N_20629);
or U29319 (N_29319,N_20075,N_20250);
and U29320 (N_29320,N_23689,N_22493);
nor U29321 (N_29321,N_21580,N_23914);
nor U29322 (N_29322,N_21999,N_21625);
nor U29323 (N_29323,N_24213,N_23395);
nand U29324 (N_29324,N_20931,N_23809);
nor U29325 (N_29325,N_23767,N_20224);
nand U29326 (N_29326,N_23223,N_21689);
or U29327 (N_29327,N_22737,N_20722);
nand U29328 (N_29328,N_24661,N_24031);
or U29329 (N_29329,N_23784,N_24952);
xor U29330 (N_29330,N_24915,N_24669);
or U29331 (N_29331,N_20574,N_20614);
or U29332 (N_29332,N_20375,N_21095);
xor U29333 (N_29333,N_22196,N_23206);
nand U29334 (N_29334,N_21317,N_24346);
nand U29335 (N_29335,N_22516,N_23935);
xnor U29336 (N_29336,N_22801,N_21689);
or U29337 (N_29337,N_22218,N_23458);
nand U29338 (N_29338,N_22755,N_23046);
or U29339 (N_29339,N_21644,N_24781);
and U29340 (N_29340,N_21184,N_23090);
nand U29341 (N_29341,N_24458,N_20993);
or U29342 (N_29342,N_22641,N_23036);
and U29343 (N_29343,N_24981,N_22831);
nor U29344 (N_29344,N_22523,N_24457);
and U29345 (N_29345,N_23880,N_20632);
xor U29346 (N_29346,N_22885,N_23713);
and U29347 (N_29347,N_20538,N_23462);
nor U29348 (N_29348,N_22850,N_21675);
nand U29349 (N_29349,N_23191,N_24838);
and U29350 (N_29350,N_21288,N_21740);
xor U29351 (N_29351,N_22582,N_20977);
xnor U29352 (N_29352,N_20179,N_24406);
and U29353 (N_29353,N_24999,N_21641);
or U29354 (N_29354,N_23211,N_22333);
nand U29355 (N_29355,N_23638,N_22208);
nand U29356 (N_29356,N_24466,N_23907);
or U29357 (N_29357,N_20462,N_20030);
or U29358 (N_29358,N_20570,N_23959);
and U29359 (N_29359,N_24686,N_23286);
and U29360 (N_29360,N_23035,N_22910);
nand U29361 (N_29361,N_22220,N_20794);
nand U29362 (N_29362,N_20803,N_23212);
and U29363 (N_29363,N_24202,N_20061);
nor U29364 (N_29364,N_24125,N_21787);
and U29365 (N_29365,N_21344,N_22503);
xnor U29366 (N_29366,N_22454,N_20763);
nand U29367 (N_29367,N_23044,N_20573);
and U29368 (N_29368,N_23042,N_21760);
or U29369 (N_29369,N_22828,N_20729);
and U29370 (N_29370,N_23559,N_24724);
nor U29371 (N_29371,N_21976,N_24746);
nor U29372 (N_29372,N_20513,N_20750);
and U29373 (N_29373,N_23832,N_24894);
nor U29374 (N_29374,N_22981,N_23027);
and U29375 (N_29375,N_21122,N_21708);
nand U29376 (N_29376,N_22926,N_20590);
and U29377 (N_29377,N_23059,N_24424);
nand U29378 (N_29378,N_22133,N_22138);
nor U29379 (N_29379,N_23793,N_20020);
nand U29380 (N_29380,N_24689,N_24471);
and U29381 (N_29381,N_20770,N_20848);
xnor U29382 (N_29382,N_24902,N_23667);
xor U29383 (N_29383,N_23833,N_22951);
xnor U29384 (N_29384,N_23431,N_24859);
and U29385 (N_29385,N_22664,N_21591);
xnor U29386 (N_29386,N_22093,N_23839);
and U29387 (N_29387,N_23230,N_23860);
and U29388 (N_29388,N_23611,N_21067);
nor U29389 (N_29389,N_24573,N_22132);
or U29390 (N_29390,N_24317,N_21270);
xor U29391 (N_29391,N_20646,N_20957);
nand U29392 (N_29392,N_21412,N_22231);
or U29393 (N_29393,N_22686,N_24310);
xnor U29394 (N_29394,N_24846,N_23401);
xor U29395 (N_29395,N_23045,N_22253);
and U29396 (N_29396,N_22359,N_20219);
and U29397 (N_29397,N_22401,N_23389);
nor U29398 (N_29398,N_20488,N_24159);
or U29399 (N_29399,N_20303,N_20670);
xor U29400 (N_29400,N_24619,N_21010);
nor U29401 (N_29401,N_21162,N_24997);
xor U29402 (N_29402,N_21711,N_24824);
nor U29403 (N_29403,N_21700,N_20027);
nand U29404 (N_29404,N_23951,N_20889);
and U29405 (N_29405,N_22133,N_20835);
and U29406 (N_29406,N_20235,N_24204);
nor U29407 (N_29407,N_20249,N_20579);
nor U29408 (N_29408,N_22639,N_22811);
and U29409 (N_29409,N_24661,N_20218);
nand U29410 (N_29410,N_23750,N_20586);
and U29411 (N_29411,N_23512,N_22212);
xor U29412 (N_29412,N_22627,N_20446);
or U29413 (N_29413,N_20584,N_20777);
nor U29414 (N_29414,N_24894,N_21112);
and U29415 (N_29415,N_20650,N_23603);
nand U29416 (N_29416,N_21491,N_22807);
or U29417 (N_29417,N_20859,N_24721);
nor U29418 (N_29418,N_20300,N_20200);
nand U29419 (N_29419,N_20553,N_22160);
nor U29420 (N_29420,N_21991,N_20386);
nor U29421 (N_29421,N_24168,N_22618);
and U29422 (N_29422,N_21277,N_24548);
or U29423 (N_29423,N_23546,N_22052);
or U29424 (N_29424,N_22083,N_22335);
xnor U29425 (N_29425,N_22281,N_20889);
and U29426 (N_29426,N_20563,N_23002);
nand U29427 (N_29427,N_21403,N_20100);
xnor U29428 (N_29428,N_22689,N_22113);
or U29429 (N_29429,N_23428,N_20781);
xor U29430 (N_29430,N_20928,N_24087);
xor U29431 (N_29431,N_21951,N_24441);
nand U29432 (N_29432,N_22155,N_22963);
or U29433 (N_29433,N_20836,N_23044);
or U29434 (N_29434,N_22953,N_24377);
xor U29435 (N_29435,N_21034,N_20525);
nand U29436 (N_29436,N_20421,N_20744);
nand U29437 (N_29437,N_24158,N_20992);
nor U29438 (N_29438,N_21726,N_20524);
nand U29439 (N_29439,N_24696,N_20995);
and U29440 (N_29440,N_24471,N_21933);
nand U29441 (N_29441,N_20679,N_21399);
or U29442 (N_29442,N_23695,N_21586);
and U29443 (N_29443,N_23012,N_23285);
and U29444 (N_29444,N_21839,N_20550);
nand U29445 (N_29445,N_22496,N_24806);
xnor U29446 (N_29446,N_21544,N_21951);
xnor U29447 (N_29447,N_23111,N_24301);
xnor U29448 (N_29448,N_20412,N_22433);
xnor U29449 (N_29449,N_21586,N_20045);
or U29450 (N_29450,N_21783,N_24321);
nor U29451 (N_29451,N_24851,N_23383);
or U29452 (N_29452,N_22841,N_22205);
or U29453 (N_29453,N_21682,N_23873);
xnor U29454 (N_29454,N_21524,N_21265);
and U29455 (N_29455,N_23090,N_23875);
and U29456 (N_29456,N_24409,N_21130);
nand U29457 (N_29457,N_20171,N_20029);
and U29458 (N_29458,N_20559,N_21453);
xor U29459 (N_29459,N_23660,N_24929);
nand U29460 (N_29460,N_24101,N_24315);
nor U29461 (N_29461,N_22333,N_20847);
and U29462 (N_29462,N_22032,N_24206);
nor U29463 (N_29463,N_23028,N_23826);
nor U29464 (N_29464,N_21026,N_23676);
nor U29465 (N_29465,N_24674,N_20330);
and U29466 (N_29466,N_21004,N_24271);
xnor U29467 (N_29467,N_20296,N_21646);
or U29468 (N_29468,N_20784,N_22288);
xor U29469 (N_29469,N_22159,N_24900);
nor U29470 (N_29470,N_22577,N_22054);
and U29471 (N_29471,N_20968,N_24123);
nor U29472 (N_29472,N_24622,N_23672);
xor U29473 (N_29473,N_24840,N_23557);
or U29474 (N_29474,N_21726,N_24181);
xor U29475 (N_29475,N_20871,N_20107);
xnor U29476 (N_29476,N_20338,N_22644);
or U29477 (N_29477,N_24877,N_24750);
and U29478 (N_29478,N_21457,N_21076);
nand U29479 (N_29479,N_23536,N_24318);
and U29480 (N_29480,N_21601,N_23359);
nor U29481 (N_29481,N_23114,N_24886);
and U29482 (N_29482,N_22049,N_23871);
or U29483 (N_29483,N_21538,N_20500);
and U29484 (N_29484,N_22503,N_23081);
or U29485 (N_29485,N_21927,N_24471);
xnor U29486 (N_29486,N_22352,N_23622);
nand U29487 (N_29487,N_20747,N_22697);
nand U29488 (N_29488,N_24029,N_21041);
nand U29489 (N_29489,N_20920,N_24300);
or U29490 (N_29490,N_21324,N_21842);
nor U29491 (N_29491,N_21911,N_24859);
and U29492 (N_29492,N_24890,N_21214);
nand U29493 (N_29493,N_22140,N_20825);
or U29494 (N_29494,N_22365,N_20382);
xor U29495 (N_29495,N_20583,N_23605);
xor U29496 (N_29496,N_23407,N_24544);
and U29497 (N_29497,N_23577,N_23395);
nor U29498 (N_29498,N_20674,N_20767);
and U29499 (N_29499,N_20386,N_24160);
or U29500 (N_29500,N_23632,N_20000);
and U29501 (N_29501,N_22457,N_21635);
nor U29502 (N_29502,N_20712,N_21111);
and U29503 (N_29503,N_21721,N_24530);
and U29504 (N_29504,N_21645,N_24830);
and U29505 (N_29505,N_23970,N_20013);
or U29506 (N_29506,N_22673,N_22642);
xor U29507 (N_29507,N_23717,N_22245);
xor U29508 (N_29508,N_20044,N_22302);
nand U29509 (N_29509,N_21250,N_24226);
or U29510 (N_29510,N_20384,N_21328);
nand U29511 (N_29511,N_22781,N_22054);
nand U29512 (N_29512,N_20855,N_22740);
or U29513 (N_29513,N_23761,N_20023);
or U29514 (N_29514,N_23948,N_20200);
nor U29515 (N_29515,N_20607,N_22562);
nor U29516 (N_29516,N_22379,N_22750);
or U29517 (N_29517,N_21330,N_20734);
nor U29518 (N_29518,N_23927,N_24478);
xor U29519 (N_29519,N_22459,N_21665);
and U29520 (N_29520,N_21928,N_21840);
xor U29521 (N_29521,N_22271,N_23539);
or U29522 (N_29522,N_21941,N_21010);
or U29523 (N_29523,N_20185,N_24321);
xnor U29524 (N_29524,N_23942,N_24027);
nor U29525 (N_29525,N_24770,N_22590);
xnor U29526 (N_29526,N_21370,N_22238);
or U29527 (N_29527,N_24830,N_21090);
nand U29528 (N_29528,N_20772,N_21414);
xnor U29529 (N_29529,N_23439,N_23835);
and U29530 (N_29530,N_24566,N_20557);
or U29531 (N_29531,N_21901,N_23036);
xnor U29532 (N_29532,N_23349,N_24738);
and U29533 (N_29533,N_20278,N_23559);
or U29534 (N_29534,N_23984,N_22193);
and U29535 (N_29535,N_22475,N_23191);
nor U29536 (N_29536,N_21188,N_20183);
nor U29537 (N_29537,N_20645,N_21881);
or U29538 (N_29538,N_22060,N_20159);
nand U29539 (N_29539,N_24192,N_20910);
xor U29540 (N_29540,N_23749,N_24361);
and U29541 (N_29541,N_20882,N_20329);
nand U29542 (N_29542,N_20711,N_21130);
nand U29543 (N_29543,N_20060,N_24519);
nor U29544 (N_29544,N_20673,N_22277);
xor U29545 (N_29545,N_22445,N_24210);
nand U29546 (N_29546,N_24525,N_24593);
or U29547 (N_29547,N_22140,N_22956);
nand U29548 (N_29548,N_21031,N_21000);
nor U29549 (N_29549,N_20777,N_21260);
and U29550 (N_29550,N_24698,N_20858);
nor U29551 (N_29551,N_22071,N_23628);
nor U29552 (N_29552,N_23019,N_20378);
or U29553 (N_29553,N_22482,N_20770);
and U29554 (N_29554,N_20949,N_21157);
xor U29555 (N_29555,N_24240,N_22677);
xor U29556 (N_29556,N_21942,N_21947);
and U29557 (N_29557,N_21729,N_23249);
or U29558 (N_29558,N_20465,N_22675);
and U29559 (N_29559,N_24808,N_21248);
or U29560 (N_29560,N_24522,N_24397);
nand U29561 (N_29561,N_20853,N_23391);
nor U29562 (N_29562,N_24357,N_24967);
and U29563 (N_29563,N_22461,N_21529);
xnor U29564 (N_29564,N_22583,N_24235);
or U29565 (N_29565,N_21878,N_21448);
xor U29566 (N_29566,N_23331,N_24081);
and U29567 (N_29567,N_22385,N_23978);
nand U29568 (N_29568,N_20135,N_23021);
xor U29569 (N_29569,N_20674,N_24712);
or U29570 (N_29570,N_23729,N_23892);
xor U29571 (N_29571,N_23316,N_20909);
xnor U29572 (N_29572,N_22258,N_23584);
xnor U29573 (N_29573,N_21455,N_23078);
or U29574 (N_29574,N_21787,N_20169);
and U29575 (N_29575,N_20162,N_21579);
nand U29576 (N_29576,N_22385,N_22072);
nor U29577 (N_29577,N_20730,N_21134);
nand U29578 (N_29578,N_20744,N_22656);
xor U29579 (N_29579,N_20790,N_22591);
and U29580 (N_29580,N_24943,N_21285);
xor U29581 (N_29581,N_22832,N_22017);
nand U29582 (N_29582,N_21430,N_24225);
nor U29583 (N_29583,N_23708,N_23833);
xnor U29584 (N_29584,N_21484,N_23845);
and U29585 (N_29585,N_20145,N_20870);
xor U29586 (N_29586,N_20475,N_21067);
nand U29587 (N_29587,N_24079,N_23985);
and U29588 (N_29588,N_20689,N_23976);
or U29589 (N_29589,N_24422,N_24116);
nand U29590 (N_29590,N_21541,N_20687);
and U29591 (N_29591,N_20626,N_20644);
and U29592 (N_29592,N_23509,N_20159);
and U29593 (N_29593,N_21493,N_20891);
and U29594 (N_29594,N_22805,N_22457);
or U29595 (N_29595,N_21234,N_22192);
nand U29596 (N_29596,N_20258,N_22218);
nor U29597 (N_29597,N_22246,N_22077);
xor U29598 (N_29598,N_23255,N_22166);
nand U29599 (N_29599,N_22449,N_21300);
xor U29600 (N_29600,N_20821,N_23827);
nor U29601 (N_29601,N_21577,N_24729);
nand U29602 (N_29602,N_22988,N_22478);
or U29603 (N_29603,N_20723,N_20564);
xor U29604 (N_29604,N_21992,N_22188);
and U29605 (N_29605,N_21983,N_21162);
xnor U29606 (N_29606,N_22427,N_21890);
xor U29607 (N_29607,N_23222,N_23426);
and U29608 (N_29608,N_23790,N_22514);
or U29609 (N_29609,N_24279,N_22045);
nand U29610 (N_29610,N_21942,N_20115);
and U29611 (N_29611,N_21504,N_22267);
xnor U29612 (N_29612,N_21527,N_22718);
xnor U29613 (N_29613,N_24989,N_20281);
or U29614 (N_29614,N_21613,N_23978);
nor U29615 (N_29615,N_22724,N_22425);
and U29616 (N_29616,N_23023,N_24667);
xor U29617 (N_29617,N_23777,N_22175);
nand U29618 (N_29618,N_22036,N_22914);
and U29619 (N_29619,N_20755,N_24327);
and U29620 (N_29620,N_22263,N_21178);
or U29621 (N_29621,N_20027,N_22674);
and U29622 (N_29622,N_20667,N_22877);
nand U29623 (N_29623,N_20221,N_20194);
nor U29624 (N_29624,N_24444,N_24055);
xor U29625 (N_29625,N_22762,N_20536);
xor U29626 (N_29626,N_24484,N_23738);
nor U29627 (N_29627,N_21693,N_20602);
nor U29628 (N_29628,N_23147,N_21238);
or U29629 (N_29629,N_21126,N_24425);
nand U29630 (N_29630,N_21986,N_22328);
nor U29631 (N_29631,N_24973,N_22082);
or U29632 (N_29632,N_22249,N_22321);
nor U29633 (N_29633,N_22452,N_22542);
or U29634 (N_29634,N_20170,N_24748);
nand U29635 (N_29635,N_20364,N_22783);
nor U29636 (N_29636,N_22414,N_20518);
xor U29637 (N_29637,N_20394,N_20884);
xor U29638 (N_29638,N_23341,N_22415);
nor U29639 (N_29639,N_23757,N_22238);
nand U29640 (N_29640,N_23637,N_22938);
nand U29641 (N_29641,N_24923,N_24870);
nand U29642 (N_29642,N_20955,N_21403);
nor U29643 (N_29643,N_24227,N_23674);
xnor U29644 (N_29644,N_22925,N_22427);
nor U29645 (N_29645,N_20237,N_23640);
xnor U29646 (N_29646,N_22152,N_23410);
xnor U29647 (N_29647,N_20244,N_22800);
nand U29648 (N_29648,N_22799,N_20067);
or U29649 (N_29649,N_21102,N_23969);
or U29650 (N_29650,N_20921,N_21186);
nand U29651 (N_29651,N_20200,N_24102);
nand U29652 (N_29652,N_20262,N_24405);
or U29653 (N_29653,N_24533,N_24594);
or U29654 (N_29654,N_23034,N_20158);
and U29655 (N_29655,N_20329,N_24959);
or U29656 (N_29656,N_20200,N_20542);
and U29657 (N_29657,N_24243,N_22678);
nor U29658 (N_29658,N_20099,N_24143);
nand U29659 (N_29659,N_23947,N_20453);
xor U29660 (N_29660,N_22341,N_23005);
nor U29661 (N_29661,N_23086,N_22358);
xnor U29662 (N_29662,N_24541,N_23147);
nand U29663 (N_29663,N_22097,N_24881);
nor U29664 (N_29664,N_22826,N_23302);
xnor U29665 (N_29665,N_20222,N_21168);
xnor U29666 (N_29666,N_21396,N_23146);
and U29667 (N_29667,N_21172,N_20868);
xor U29668 (N_29668,N_24378,N_24997);
and U29669 (N_29669,N_20878,N_21169);
or U29670 (N_29670,N_24849,N_22455);
nor U29671 (N_29671,N_23781,N_24899);
nand U29672 (N_29672,N_22584,N_22407);
nor U29673 (N_29673,N_23094,N_20275);
xor U29674 (N_29674,N_24125,N_22915);
xor U29675 (N_29675,N_21164,N_24742);
nand U29676 (N_29676,N_21241,N_20978);
or U29677 (N_29677,N_21432,N_24018);
or U29678 (N_29678,N_21829,N_21619);
nand U29679 (N_29679,N_21991,N_21893);
or U29680 (N_29680,N_23696,N_20933);
nand U29681 (N_29681,N_20622,N_20078);
or U29682 (N_29682,N_20295,N_23463);
xor U29683 (N_29683,N_22063,N_24078);
xor U29684 (N_29684,N_24226,N_22541);
nor U29685 (N_29685,N_21297,N_22540);
nor U29686 (N_29686,N_23850,N_23742);
xor U29687 (N_29687,N_21446,N_20849);
and U29688 (N_29688,N_20056,N_21572);
or U29689 (N_29689,N_21728,N_22043);
or U29690 (N_29690,N_20637,N_20088);
nor U29691 (N_29691,N_24338,N_20723);
nand U29692 (N_29692,N_24628,N_23171);
and U29693 (N_29693,N_21257,N_24360);
nor U29694 (N_29694,N_22375,N_20994);
or U29695 (N_29695,N_22930,N_23301);
or U29696 (N_29696,N_24110,N_22705);
and U29697 (N_29697,N_21963,N_21940);
xor U29698 (N_29698,N_21020,N_24766);
nor U29699 (N_29699,N_22049,N_22459);
and U29700 (N_29700,N_20303,N_23250);
xor U29701 (N_29701,N_20195,N_20192);
xor U29702 (N_29702,N_21050,N_20814);
nor U29703 (N_29703,N_22188,N_22858);
nor U29704 (N_29704,N_23833,N_20920);
nand U29705 (N_29705,N_20871,N_21804);
and U29706 (N_29706,N_21700,N_21929);
or U29707 (N_29707,N_20420,N_23935);
or U29708 (N_29708,N_21163,N_22175);
and U29709 (N_29709,N_20310,N_22635);
xor U29710 (N_29710,N_21986,N_22577);
and U29711 (N_29711,N_22197,N_24473);
nor U29712 (N_29712,N_24783,N_20184);
or U29713 (N_29713,N_24889,N_24740);
and U29714 (N_29714,N_24376,N_22448);
and U29715 (N_29715,N_20423,N_23503);
and U29716 (N_29716,N_22832,N_20141);
and U29717 (N_29717,N_24325,N_20379);
xnor U29718 (N_29718,N_21378,N_20407);
or U29719 (N_29719,N_20799,N_22897);
and U29720 (N_29720,N_22898,N_24474);
xor U29721 (N_29721,N_22518,N_20144);
nor U29722 (N_29722,N_20428,N_23867);
nand U29723 (N_29723,N_23945,N_22630);
nand U29724 (N_29724,N_22701,N_23512);
and U29725 (N_29725,N_24836,N_21150);
nand U29726 (N_29726,N_23852,N_21555);
xnor U29727 (N_29727,N_21200,N_23626);
xnor U29728 (N_29728,N_22595,N_22831);
or U29729 (N_29729,N_24904,N_22926);
nand U29730 (N_29730,N_22711,N_22512);
or U29731 (N_29731,N_21803,N_22828);
or U29732 (N_29732,N_22883,N_23373);
nor U29733 (N_29733,N_20261,N_24707);
nand U29734 (N_29734,N_20283,N_23677);
nor U29735 (N_29735,N_23403,N_20296);
nand U29736 (N_29736,N_23970,N_22968);
or U29737 (N_29737,N_21878,N_23989);
or U29738 (N_29738,N_22376,N_24670);
xnor U29739 (N_29739,N_23649,N_23192);
nand U29740 (N_29740,N_24119,N_23531);
or U29741 (N_29741,N_21586,N_21031);
or U29742 (N_29742,N_22163,N_22008);
xor U29743 (N_29743,N_22135,N_22014);
xor U29744 (N_29744,N_24203,N_20250);
nor U29745 (N_29745,N_23043,N_20832);
and U29746 (N_29746,N_20152,N_23115);
nor U29747 (N_29747,N_20330,N_23910);
nand U29748 (N_29748,N_23800,N_22997);
nor U29749 (N_29749,N_21574,N_23086);
xnor U29750 (N_29750,N_22487,N_24451);
or U29751 (N_29751,N_22613,N_24910);
nand U29752 (N_29752,N_23802,N_21344);
xnor U29753 (N_29753,N_23696,N_21584);
and U29754 (N_29754,N_24682,N_20946);
nand U29755 (N_29755,N_24472,N_23988);
or U29756 (N_29756,N_20961,N_20893);
xnor U29757 (N_29757,N_22442,N_20044);
nor U29758 (N_29758,N_23516,N_20786);
xnor U29759 (N_29759,N_20778,N_20989);
and U29760 (N_29760,N_23649,N_23568);
or U29761 (N_29761,N_21073,N_22630);
nand U29762 (N_29762,N_24613,N_23661);
nor U29763 (N_29763,N_23384,N_20419);
nand U29764 (N_29764,N_20600,N_24653);
nand U29765 (N_29765,N_22195,N_20443);
nor U29766 (N_29766,N_23662,N_22265);
xnor U29767 (N_29767,N_20200,N_23511);
nand U29768 (N_29768,N_23933,N_24197);
or U29769 (N_29769,N_21064,N_24728);
nand U29770 (N_29770,N_24314,N_20102);
nand U29771 (N_29771,N_20865,N_21268);
or U29772 (N_29772,N_24473,N_20193);
nand U29773 (N_29773,N_20933,N_21238);
or U29774 (N_29774,N_23175,N_24813);
xnor U29775 (N_29775,N_21712,N_23505);
and U29776 (N_29776,N_21334,N_23378);
and U29777 (N_29777,N_24598,N_23514);
and U29778 (N_29778,N_23056,N_23077);
nand U29779 (N_29779,N_24410,N_22734);
nand U29780 (N_29780,N_23419,N_23161);
xnor U29781 (N_29781,N_23590,N_21378);
nand U29782 (N_29782,N_24430,N_23771);
xnor U29783 (N_29783,N_22650,N_22748);
or U29784 (N_29784,N_22749,N_22070);
or U29785 (N_29785,N_20999,N_20195);
nand U29786 (N_29786,N_23547,N_23623);
or U29787 (N_29787,N_21441,N_21364);
nor U29788 (N_29788,N_23222,N_22537);
or U29789 (N_29789,N_22238,N_21343);
nor U29790 (N_29790,N_22549,N_20939);
and U29791 (N_29791,N_20147,N_24273);
nand U29792 (N_29792,N_22695,N_23548);
xor U29793 (N_29793,N_24292,N_23238);
or U29794 (N_29794,N_24169,N_23895);
nor U29795 (N_29795,N_21374,N_20029);
or U29796 (N_29796,N_22255,N_22961);
nand U29797 (N_29797,N_24663,N_23215);
and U29798 (N_29798,N_24404,N_22038);
nor U29799 (N_29799,N_20862,N_23138);
or U29800 (N_29800,N_20009,N_22137);
and U29801 (N_29801,N_22025,N_24719);
nor U29802 (N_29802,N_22308,N_24890);
xor U29803 (N_29803,N_20018,N_24610);
xor U29804 (N_29804,N_20126,N_22039);
and U29805 (N_29805,N_20557,N_23133);
or U29806 (N_29806,N_21595,N_22271);
and U29807 (N_29807,N_24537,N_20056);
nand U29808 (N_29808,N_22763,N_22098);
nand U29809 (N_29809,N_23990,N_24475);
nand U29810 (N_29810,N_21350,N_24446);
nand U29811 (N_29811,N_20314,N_21143);
or U29812 (N_29812,N_23255,N_24119);
nand U29813 (N_29813,N_23596,N_22254);
and U29814 (N_29814,N_24866,N_22767);
xnor U29815 (N_29815,N_21364,N_24527);
nand U29816 (N_29816,N_24713,N_22389);
nor U29817 (N_29817,N_21334,N_22940);
nand U29818 (N_29818,N_22508,N_23999);
nor U29819 (N_29819,N_21592,N_24199);
nand U29820 (N_29820,N_20564,N_22208);
and U29821 (N_29821,N_24793,N_23089);
nand U29822 (N_29822,N_20697,N_21824);
and U29823 (N_29823,N_20668,N_22452);
or U29824 (N_29824,N_22638,N_22077);
nor U29825 (N_29825,N_20349,N_21099);
xor U29826 (N_29826,N_20621,N_21559);
nand U29827 (N_29827,N_20658,N_24890);
nor U29828 (N_29828,N_23273,N_24303);
nor U29829 (N_29829,N_23893,N_22517);
or U29830 (N_29830,N_24374,N_20613);
and U29831 (N_29831,N_21820,N_20051);
and U29832 (N_29832,N_24388,N_23867);
and U29833 (N_29833,N_22372,N_22735);
xor U29834 (N_29834,N_21171,N_23003);
and U29835 (N_29835,N_21690,N_23538);
or U29836 (N_29836,N_20708,N_20383);
and U29837 (N_29837,N_22595,N_20912);
nor U29838 (N_29838,N_23838,N_22729);
xor U29839 (N_29839,N_22765,N_23280);
xnor U29840 (N_29840,N_23546,N_22364);
xor U29841 (N_29841,N_24236,N_22003);
xnor U29842 (N_29842,N_20736,N_21307);
or U29843 (N_29843,N_23687,N_21276);
or U29844 (N_29844,N_24196,N_20838);
nor U29845 (N_29845,N_20442,N_24675);
or U29846 (N_29846,N_24976,N_21788);
nor U29847 (N_29847,N_20193,N_21118);
nor U29848 (N_29848,N_24619,N_20480);
nand U29849 (N_29849,N_21815,N_22138);
nand U29850 (N_29850,N_21981,N_21757);
nor U29851 (N_29851,N_23670,N_22808);
nor U29852 (N_29852,N_20597,N_20141);
nor U29853 (N_29853,N_22474,N_22493);
or U29854 (N_29854,N_20419,N_23864);
nand U29855 (N_29855,N_21944,N_23225);
xnor U29856 (N_29856,N_22203,N_23896);
xnor U29857 (N_29857,N_23627,N_22217);
and U29858 (N_29858,N_20693,N_20972);
nor U29859 (N_29859,N_22850,N_23049);
nor U29860 (N_29860,N_24382,N_23906);
and U29861 (N_29861,N_22922,N_23632);
xor U29862 (N_29862,N_21574,N_22570);
or U29863 (N_29863,N_20362,N_23497);
xor U29864 (N_29864,N_21508,N_23805);
nand U29865 (N_29865,N_24187,N_22455);
nor U29866 (N_29866,N_22261,N_24918);
and U29867 (N_29867,N_24792,N_23515);
or U29868 (N_29868,N_24253,N_20598);
nor U29869 (N_29869,N_23249,N_22969);
xor U29870 (N_29870,N_24698,N_20777);
nand U29871 (N_29871,N_22543,N_22354);
or U29872 (N_29872,N_22463,N_23995);
xor U29873 (N_29873,N_22304,N_20362);
or U29874 (N_29874,N_23395,N_21394);
or U29875 (N_29875,N_24065,N_24761);
nor U29876 (N_29876,N_23602,N_23541);
nand U29877 (N_29877,N_23541,N_22435);
xor U29878 (N_29878,N_20273,N_23411);
or U29879 (N_29879,N_24527,N_21711);
nor U29880 (N_29880,N_20792,N_23697);
xor U29881 (N_29881,N_20359,N_20629);
xnor U29882 (N_29882,N_22510,N_24580);
nor U29883 (N_29883,N_23002,N_23014);
and U29884 (N_29884,N_23999,N_21016);
or U29885 (N_29885,N_22810,N_23031);
xnor U29886 (N_29886,N_21024,N_20687);
nor U29887 (N_29887,N_23597,N_22123);
xnor U29888 (N_29888,N_24072,N_23496);
and U29889 (N_29889,N_24806,N_24222);
and U29890 (N_29890,N_24106,N_24204);
nor U29891 (N_29891,N_23038,N_24302);
and U29892 (N_29892,N_24275,N_23664);
or U29893 (N_29893,N_21495,N_24025);
nand U29894 (N_29894,N_22216,N_20351);
or U29895 (N_29895,N_20166,N_23379);
and U29896 (N_29896,N_21376,N_22018);
and U29897 (N_29897,N_22006,N_23265);
nand U29898 (N_29898,N_22892,N_22044);
nor U29899 (N_29899,N_21610,N_20755);
nand U29900 (N_29900,N_24024,N_22778);
and U29901 (N_29901,N_22577,N_24884);
or U29902 (N_29902,N_21302,N_23215);
or U29903 (N_29903,N_21099,N_20888);
nor U29904 (N_29904,N_21969,N_21521);
nand U29905 (N_29905,N_21798,N_21712);
xor U29906 (N_29906,N_24687,N_22876);
nor U29907 (N_29907,N_22034,N_20163);
or U29908 (N_29908,N_20652,N_22175);
nor U29909 (N_29909,N_23507,N_20356);
and U29910 (N_29910,N_23153,N_24581);
or U29911 (N_29911,N_20398,N_24160);
nor U29912 (N_29912,N_24326,N_24631);
or U29913 (N_29913,N_22400,N_22417);
or U29914 (N_29914,N_23744,N_21941);
nand U29915 (N_29915,N_22241,N_21077);
nor U29916 (N_29916,N_20069,N_23014);
xnor U29917 (N_29917,N_21752,N_22024);
or U29918 (N_29918,N_23553,N_20086);
nand U29919 (N_29919,N_22288,N_21932);
nand U29920 (N_29920,N_21513,N_22583);
nor U29921 (N_29921,N_20814,N_22815);
xnor U29922 (N_29922,N_21285,N_24510);
xnor U29923 (N_29923,N_23616,N_22247);
xnor U29924 (N_29924,N_20083,N_23361);
nand U29925 (N_29925,N_20472,N_21178);
xnor U29926 (N_29926,N_23720,N_24447);
and U29927 (N_29927,N_24885,N_23120);
and U29928 (N_29928,N_22511,N_24646);
xor U29929 (N_29929,N_21043,N_24345);
and U29930 (N_29930,N_22038,N_23778);
or U29931 (N_29931,N_24133,N_20996);
xnor U29932 (N_29932,N_22786,N_21147);
or U29933 (N_29933,N_20061,N_21304);
nor U29934 (N_29934,N_21459,N_22982);
nor U29935 (N_29935,N_23186,N_21833);
and U29936 (N_29936,N_22204,N_24714);
and U29937 (N_29937,N_22089,N_21055);
or U29938 (N_29938,N_24346,N_23285);
and U29939 (N_29939,N_20777,N_24251);
nand U29940 (N_29940,N_24887,N_24411);
nor U29941 (N_29941,N_20263,N_24329);
and U29942 (N_29942,N_24553,N_23088);
and U29943 (N_29943,N_21189,N_21416);
nor U29944 (N_29944,N_21195,N_24479);
xnor U29945 (N_29945,N_20085,N_21719);
nor U29946 (N_29946,N_24338,N_23989);
or U29947 (N_29947,N_24565,N_22514);
and U29948 (N_29948,N_22860,N_21399);
nand U29949 (N_29949,N_23733,N_20445);
and U29950 (N_29950,N_20545,N_21344);
or U29951 (N_29951,N_22085,N_23272);
and U29952 (N_29952,N_23987,N_20434);
nor U29953 (N_29953,N_20964,N_20860);
nor U29954 (N_29954,N_22391,N_21741);
or U29955 (N_29955,N_23419,N_21982);
xnor U29956 (N_29956,N_23036,N_21335);
and U29957 (N_29957,N_21904,N_24753);
and U29958 (N_29958,N_22141,N_23109);
xor U29959 (N_29959,N_22270,N_20358);
or U29960 (N_29960,N_20349,N_24564);
nand U29961 (N_29961,N_21808,N_22678);
xnor U29962 (N_29962,N_23478,N_21476);
xor U29963 (N_29963,N_23538,N_22719);
and U29964 (N_29964,N_22527,N_21499);
nor U29965 (N_29965,N_20919,N_20504);
nand U29966 (N_29966,N_21729,N_20074);
nand U29967 (N_29967,N_23892,N_23438);
and U29968 (N_29968,N_23347,N_21919);
nor U29969 (N_29969,N_21943,N_24194);
xnor U29970 (N_29970,N_21775,N_24306);
or U29971 (N_29971,N_20909,N_23653);
xnor U29972 (N_29972,N_24032,N_20228);
or U29973 (N_29973,N_20051,N_21569);
and U29974 (N_29974,N_21180,N_23723);
xnor U29975 (N_29975,N_21939,N_23129);
nand U29976 (N_29976,N_20927,N_21687);
or U29977 (N_29977,N_21997,N_24778);
nand U29978 (N_29978,N_21806,N_23051);
nand U29979 (N_29979,N_20799,N_22885);
or U29980 (N_29980,N_24920,N_22575);
and U29981 (N_29981,N_22346,N_20297);
or U29982 (N_29982,N_24670,N_23074);
and U29983 (N_29983,N_24163,N_22843);
xnor U29984 (N_29984,N_23707,N_24786);
xnor U29985 (N_29985,N_20188,N_24700);
and U29986 (N_29986,N_23397,N_23949);
or U29987 (N_29987,N_22429,N_22422);
and U29988 (N_29988,N_24033,N_21564);
and U29989 (N_29989,N_21407,N_24271);
nor U29990 (N_29990,N_23653,N_23039);
nor U29991 (N_29991,N_22616,N_23821);
or U29992 (N_29992,N_20609,N_20716);
and U29993 (N_29993,N_20707,N_21370);
nand U29994 (N_29994,N_20989,N_23747);
nor U29995 (N_29995,N_22420,N_24623);
nor U29996 (N_29996,N_23146,N_21730);
nor U29997 (N_29997,N_23082,N_22449);
or U29998 (N_29998,N_23008,N_22991);
and U29999 (N_29999,N_24219,N_21698);
xnor UO_0 (O_0,N_25953,N_29007);
or UO_1 (O_1,N_28070,N_28088);
xor UO_2 (O_2,N_29947,N_25032);
nor UO_3 (O_3,N_25337,N_25475);
nand UO_4 (O_4,N_27027,N_27283);
and UO_5 (O_5,N_25140,N_27547);
nor UO_6 (O_6,N_28201,N_27537);
nand UO_7 (O_7,N_27707,N_26927);
xor UO_8 (O_8,N_28035,N_27139);
nor UO_9 (O_9,N_25273,N_28658);
nand UO_10 (O_10,N_29418,N_27160);
nor UO_11 (O_11,N_28992,N_27685);
nand UO_12 (O_12,N_28001,N_26162);
xnor UO_13 (O_13,N_25698,N_26269);
nor UO_14 (O_14,N_28863,N_28282);
nor UO_15 (O_15,N_27640,N_26428);
nand UO_16 (O_16,N_27338,N_25990);
nor UO_17 (O_17,N_28140,N_26544);
nor UO_18 (O_18,N_27822,N_27316);
or UO_19 (O_19,N_28570,N_26668);
xnor UO_20 (O_20,N_25454,N_29293);
or UO_21 (O_21,N_27658,N_29073);
xnor UO_22 (O_22,N_25150,N_25925);
xnor UO_23 (O_23,N_29597,N_29942);
nand UO_24 (O_24,N_29816,N_29058);
or UO_25 (O_25,N_27994,N_26849);
nand UO_26 (O_26,N_27300,N_25118);
or UO_27 (O_27,N_29477,N_26375);
and UO_28 (O_28,N_25033,N_25374);
xnor UO_29 (O_29,N_26014,N_29208);
and UO_30 (O_30,N_26785,N_28463);
or UO_31 (O_31,N_25946,N_29632);
or UO_32 (O_32,N_28676,N_27135);
and UO_33 (O_33,N_25270,N_27377);
xor UO_34 (O_34,N_27070,N_27298);
and UO_35 (O_35,N_28410,N_28978);
or UO_36 (O_36,N_29266,N_27981);
nor UO_37 (O_37,N_27986,N_29248);
xnor UO_38 (O_38,N_26638,N_25747);
or UO_39 (O_39,N_29756,N_25806);
xnor UO_40 (O_40,N_29216,N_26391);
xnor UO_41 (O_41,N_28964,N_29669);
xnor UO_42 (O_42,N_26642,N_28232);
and UO_43 (O_43,N_27016,N_29084);
nand UO_44 (O_44,N_26308,N_27617);
xnor UO_45 (O_45,N_28091,N_29228);
xnor UO_46 (O_46,N_25676,N_26692);
and UO_47 (O_47,N_28997,N_29410);
or UO_48 (O_48,N_27169,N_29618);
and UO_49 (O_49,N_29285,N_26527);
nand UO_50 (O_50,N_29015,N_25361);
xnor UO_51 (O_51,N_29503,N_26854);
and UO_52 (O_52,N_27461,N_29000);
and UO_53 (O_53,N_29106,N_28634);
nand UO_54 (O_54,N_29734,N_27832);
nand UO_55 (O_55,N_28283,N_29118);
and UO_56 (O_56,N_28173,N_29358);
or UO_57 (O_57,N_29538,N_29933);
and UO_58 (O_58,N_28860,N_26112);
xnor UO_59 (O_59,N_26604,N_25934);
or UO_60 (O_60,N_25247,N_28223);
nand UO_61 (O_61,N_29414,N_26603);
and UO_62 (O_62,N_25257,N_26369);
xnor UO_63 (O_63,N_29408,N_29970);
xor UO_64 (O_64,N_27337,N_25996);
nor UO_65 (O_65,N_27987,N_26467);
and UO_66 (O_66,N_29067,N_27924);
nand UO_67 (O_67,N_27886,N_26306);
or UO_68 (O_68,N_25711,N_26310);
and UO_69 (O_69,N_29337,N_29724);
nand UO_70 (O_70,N_28249,N_28462);
and UO_71 (O_71,N_26877,N_27155);
and UO_72 (O_72,N_28887,N_29052);
nand UO_73 (O_73,N_25165,N_26730);
nand UO_74 (O_74,N_27144,N_25899);
and UO_75 (O_75,N_29431,N_25442);
or UO_76 (O_76,N_27741,N_26568);
xnor UO_77 (O_77,N_29794,N_27454);
nor UO_78 (O_78,N_29445,N_29561);
and UO_79 (O_79,N_28251,N_29368);
xor UO_80 (O_80,N_27180,N_27747);
xor UO_81 (O_81,N_26647,N_25851);
xnor UO_82 (O_82,N_29577,N_29027);
nand UO_83 (O_83,N_26858,N_25779);
xor UO_84 (O_84,N_26390,N_25773);
or UO_85 (O_85,N_26256,N_29102);
or UO_86 (O_86,N_25269,N_28542);
nor UO_87 (O_87,N_27735,N_28652);
and UO_88 (O_88,N_25804,N_28277);
xor UO_89 (O_89,N_26127,N_28524);
or UO_90 (O_90,N_29547,N_25724);
or UO_91 (O_91,N_26452,N_25687);
nor UO_92 (O_92,N_27087,N_25305);
xor UO_93 (O_93,N_29550,N_26155);
or UO_94 (O_94,N_28981,N_29109);
nand UO_95 (O_95,N_29742,N_28465);
and UO_96 (O_96,N_25323,N_26685);
nor UO_97 (O_97,N_29344,N_26938);
nor UO_98 (O_98,N_28881,N_25670);
nor UO_99 (O_99,N_26423,N_27019);
nand UO_100 (O_100,N_25482,N_25426);
or UO_101 (O_101,N_27616,N_28019);
nor UO_102 (O_102,N_27963,N_26009);
nor UO_103 (O_103,N_28854,N_28016);
xor UO_104 (O_104,N_26096,N_25963);
or UO_105 (O_105,N_25113,N_26050);
nand UO_106 (O_106,N_29423,N_26157);
and UO_107 (O_107,N_26783,N_25436);
xor UO_108 (O_108,N_26817,N_27061);
nand UO_109 (O_109,N_26528,N_28297);
nand UO_110 (O_110,N_28954,N_26305);
xor UO_111 (O_111,N_26278,N_28377);
nor UO_112 (O_112,N_27762,N_28022);
nor UO_113 (O_113,N_28779,N_25631);
nor UO_114 (O_114,N_28559,N_26282);
nor UO_115 (O_115,N_25865,N_26786);
xnor UO_116 (O_116,N_26925,N_28170);
or UO_117 (O_117,N_26864,N_27826);
nor UO_118 (O_118,N_27938,N_29620);
or UO_119 (O_119,N_29973,N_27550);
and UO_120 (O_120,N_27076,N_25610);
or UO_121 (O_121,N_26637,N_26439);
or UO_122 (O_122,N_25285,N_27093);
nor UO_123 (O_123,N_27964,N_28453);
nor UO_124 (O_124,N_26447,N_25137);
nor UO_125 (O_125,N_27580,N_28815);
and UO_126 (O_126,N_27225,N_26116);
or UO_127 (O_127,N_27508,N_29097);
nand UO_128 (O_128,N_27397,N_25288);
and UO_129 (O_129,N_28569,N_29197);
nand UO_130 (O_130,N_27774,N_25885);
or UO_131 (O_131,N_25878,N_27692);
xor UO_132 (O_132,N_26607,N_27715);
nor UO_133 (O_133,N_29772,N_29298);
nand UO_134 (O_134,N_27669,N_28416);
nand UO_135 (O_135,N_25535,N_29617);
nand UO_136 (O_136,N_27293,N_25183);
or UO_137 (O_137,N_29966,N_29643);
nand UO_138 (O_138,N_25438,N_28422);
nor UO_139 (O_139,N_27436,N_27271);
or UO_140 (O_140,N_28608,N_29064);
and UO_141 (O_141,N_27335,N_27411);
and UO_142 (O_142,N_29926,N_25771);
or UO_143 (O_143,N_27635,N_27497);
and UO_144 (O_144,N_27425,N_26865);
nor UO_145 (O_145,N_28871,N_28840);
nand UO_146 (O_146,N_27284,N_27641);
xor UO_147 (O_147,N_28480,N_26911);
nand UO_148 (O_148,N_27967,N_29235);
nor UO_149 (O_149,N_28657,N_27344);
nand UO_150 (O_150,N_28753,N_27888);
and UO_151 (O_151,N_28379,N_27570);
xnor UO_152 (O_152,N_25763,N_27104);
nand UO_153 (O_153,N_27680,N_25427);
and UO_154 (O_154,N_25050,N_26610);
or UO_155 (O_155,N_27127,N_28373);
xnor UO_156 (O_156,N_26807,N_27566);
nor UO_157 (O_157,N_27099,N_26932);
xor UO_158 (O_158,N_27683,N_27805);
nor UO_159 (O_159,N_29232,N_28939);
nor UO_160 (O_160,N_27503,N_25754);
nor UO_161 (O_161,N_26143,N_29493);
xor UO_162 (O_162,N_29206,N_25526);
or UO_163 (O_163,N_27724,N_25404);
and UO_164 (O_164,N_28550,N_29524);
and UO_165 (O_165,N_26242,N_25044);
nand UO_166 (O_166,N_25277,N_29556);
nor UO_167 (O_167,N_29028,N_26502);
and UO_168 (O_168,N_25615,N_27278);
and UO_169 (O_169,N_29744,N_25970);
xnor UO_170 (O_170,N_25845,N_26212);
nand UO_171 (O_171,N_26689,N_29606);
xnor UO_172 (O_172,N_25518,N_29608);
or UO_173 (O_173,N_29051,N_25196);
nor UO_174 (O_174,N_28181,N_26349);
nand UO_175 (O_175,N_27361,N_25149);
and UO_176 (O_176,N_27163,N_26657);
nor UO_177 (O_177,N_28987,N_28663);
xor UO_178 (O_178,N_28213,N_28013);
or UO_179 (O_179,N_26059,N_27068);
nor UO_180 (O_180,N_29122,N_26433);
and UO_181 (O_181,N_28381,N_27460);
xnor UO_182 (O_182,N_28772,N_29726);
nand UO_183 (O_183,N_25406,N_28617);
or UO_184 (O_184,N_28384,N_25449);
xnor UO_185 (O_185,N_27542,N_25370);
nand UO_186 (O_186,N_25081,N_27522);
xor UO_187 (O_187,N_27306,N_26172);
xnor UO_188 (O_188,N_25672,N_28818);
nand UO_189 (O_189,N_26930,N_27304);
xor UO_190 (O_190,N_25998,N_28579);
nand UO_191 (O_191,N_29032,N_29854);
and UO_192 (O_192,N_26379,N_26782);
or UO_193 (O_193,N_25461,N_25551);
or UO_194 (O_194,N_28336,N_27473);
xor UO_195 (O_195,N_29145,N_29143);
xor UO_196 (O_196,N_29584,N_29765);
and UO_197 (O_197,N_26301,N_29335);
and UO_198 (O_198,N_25939,N_26694);
nor UO_199 (O_199,N_26396,N_27389);
nand UO_200 (O_200,N_28185,N_28829);
and UO_201 (O_201,N_26954,N_27329);
nor UO_202 (O_202,N_26843,N_27913);
nand UO_203 (O_203,N_27128,N_25659);
xnor UO_204 (O_204,N_25510,N_29760);
xnor UO_205 (O_205,N_29678,N_27098);
xor UO_206 (O_206,N_25173,N_25625);
or UO_207 (O_207,N_28104,N_26738);
and UO_208 (O_208,N_27631,N_26420);
nor UO_209 (O_209,N_28409,N_25513);
and UO_210 (O_210,N_25757,N_28255);
or UO_211 (O_211,N_28198,N_29317);
and UO_212 (O_212,N_27936,N_28759);
or UO_213 (O_213,N_28599,N_29336);
nand UO_214 (O_214,N_25712,N_26373);
nand UO_215 (O_215,N_27177,N_29177);
nor UO_216 (O_216,N_25046,N_26246);
and UO_217 (O_217,N_26060,N_29277);
and UO_218 (O_218,N_28915,N_26868);
and UO_219 (O_219,N_26011,N_29598);
nand UO_220 (O_220,N_27296,N_28343);
or UO_221 (O_221,N_28413,N_29091);
or UO_222 (O_222,N_27751,N_26523);
or UO_223 (O_223,N_25508,N_29803);
or UO_224 (O_224,N_28315,N_28344);
or UO_225 (O_225,N_28125,N_26389);
xnor UO_226 (O_226,N_28391,N_27840);
nor UO_227 (O_227,N_26268,N_25097);
xor UO_228 (O_228,N_25875,N_29111);
nor UO_229 (O_229,N_25142,N_27749);
or UO_230 (O_230,N_27825,N_25279);
and UO_231 (O_231,N_25221,N_28790);
and UO_232 (O_232,N_27277,N_28655);
and UO_233 (O_233,N_27727,N_29892);
xnor UO_234 (O_234,N_26315,N_25432);
or UO_235 (O_235,N_28946,N_26403);
and UO_236 (O_236,N_28673,N_26804);
and UO_237 (O_237,N_28194,N_28026);
or UO_238 (O_238,N_29735,N_26696);
xnor UO_239 (O_239,N_26431,N_27973);
xnor UO_240 (O_240,N_27555,N_29758);
or UO_241 (O_241,N_25944,N_26613);
and UO_242 (O_242,N_27009,N_27560);
and UO_243 (O_243,N_28156,N_28632);
or UO_244 (O_244,N_26944,N_26294);
xor UO_245 (O_245,N_28087,N_26350);
nand UO_246 (O_246,N_26179,N_25516);
nor UO_247 (O_247,N_25293,N_25419);
and UO_248 (O_248,N_26719,N_27067);
or UO_249 (O_249,N_28124,N_26149);
and UO_250 (O_250,N_25460,N_29108);
xor UO_251 (O_251,N_26630,N_25681);
nor UO_252 (O_252,N_25413,N_26616);
nor UO_253 (O_253,N_28446,N_27213);
nor UO_254 (O_254,N_28182,N_27173);
and UO_255 (O_255,N_28506,N_26825);
or UO_256 (O_256,N_26047,N_28627);
or UO_257 (O_257,N_28802,N_27793);
xor UO_258 (O_258,N_26651,N_28396);
nand UO_259 (O_259,N_29484,N_27063);
xor UO_260 (O_260,N_25844,N_26905);
or UO_261 (O_261,N_26208,N_25394);
xnor UO_262 (O_262,N_28101,N_28591);
nor UO_263 (O_263,N_28784,N_29812);
nor UO_264 (O_264,N_27295,N_25368);
nor UO_265 (O_265,N_29373,N_25231);
and UO_266 (O_266,N_28237,N_25544);
or UO_267 (O_267,N_26987,N_26368);
nand UO_268 (O_268,N_29221,N_26340);
and UO_269 (O_269,N_29021,N_26263);
nand UO_270 (O_270,N_27403,N_29974);
or UO_271 (O_271,N_25410,N_28195);
xnor UO_272 (O_272,N_26254,N_26444);
xnor UO_273 (O_273,N_27201,N_27519);
and UO_274 (O_274,N_25917,N_26205);
xor UO_275 (O_275,N_29976,N_29766);
xnor UO_276 (O_276,N_27999,N_26735);
nor UO_277 (O_277,N_28711,N_27319);
nand UO_278 (O_278,N_28352,N_26820);
nor UO_279 (O_279,N_27034,N_27434);
nand UO_280 (O_280,N_25457,N_27260);
or UO_281 (O_281,N_28024,N_26299);
nand UO_282 (O_282,N_25445,N_26659);
and UO_283 (O_283,N_25600,N_27770);
and UO_284 (O_284,N_26690,N_29242);
nand UO_285 (O_285,N_26290,N_29712);
nand UO_286 (O_286,N_26749,N_28667);
or UO_287 (O_287,N_27120,N_26705);
nand UO_288 (O_288,N_29539,N_29527);
xnor UO_289 (O_289,N_29323,N_29856);
xnor UO_290 (O_290,N_26354,N_28538);
nor UO_291 (O_291,N_29829,N_29708);
nor UO_292 (O_292,N_29488,N_28139);
and UO_293 (O_293,N_25131,N_27352);
nand UO_294 (O_294,N_28012,N_27607);
xor UO_295 (O_295,N_28032,N_28023);
and UO_296 (O_296,N_28965,N_27406);
nor UO_297 (O_297,N_25303,N_26592);
and UO_298 (O_298,N_28495,N_25175);
nand UO_299 (O_299,N_25507,N_27502);
and UO_300 (O_300,N_29065,N_25765);
nor UO_301 (O_301,N_26745,N_26718);
nand UO_302 (O_302,N_25566,N_26995);
or UO_303 (O_303,N_28342,N_28571);
and UO_304 (O_304,N_27970,N_25179);
nand UO_305 (O_305,N_28522,N_28735);
nand UO_306 (O_306,N_29184,N_28848);
nor UO_307 (O_307,N_27465,N_27199);
nor UO_308 (O_308,N_29241,N_27288);
or UO_309 (O_309,N_25799,N_26023);
nor UO_310 (O_310,N_29824,N_26919);
nand UO_311 (O_311,N_28199,N_25876);
nor UO_312 (O_312,N_25123,N_25141);
or UO_313 (O_313,N_25211,N_28970);
and UO_314 (O_314,N_25103,N_25127);
nor UO_315 (O_315,N_27859,N_27515);
xor UO_316 (O_316,N_27317,N_26590);
and UO_317 (O_317,N_29604,N_26139);
xnor UO_318 (O_318,N_28500,N_25941);
or UO_319 (O_319,N_26612,N_27078);
xnor UO_320 (O_320,N_28142,N_29485);
and UO_321 (O_321,N_29462,N_29723);
and UO_322 (O_322,N_29997,N_27212);
nor UO_323 (O_323,N_27846,N_25096);
nor UO_324 (O_324,N_26383,N_26572);
or UO_325 (O_325,N_25995,N_27156);
xor UO_326 (O_326,N_25005,N_25308);
xor UO_327 (O_327,N_28202,N_25655);
nor UO_328 (O_328,N_25776,N_29874);
or UO_329 (O_329,N_29621,N_29403);
xnor UO_330 (O_330,N_28934,N_28841);
or UO_331 (O_331,N_29096,N_26569);
or UO_332 (O_332,N_27387,N_27918);
nand UO_333 (O_333,N_26119,N_28705);
xnor UO_334 (O_334,N_26406,N_25100);
or UO_335 (O_335,N_26240,N_28816);
xnor UO_336 (O_336,N_28947,N_26553);
nor UO_337 (O_337,N_28543,N_26582);
nor UO_338 (O_338,N_29425,N_26704);
nor UO_339 (O_339,N_26534,N_25291);
nor UO_340 (O_340,N_28671,N_27082);
and UO_341 (O_341,N_26888,N_25856);
and UO_342 (O_342,N_27245,N_27065);
nor UO_343 (O_343,N_28021,N_28171);
xor UO_344 (O_344,N_28828,N_28197);
xnor UO_345 (O_345,N_26627,N_29819);
xor UO_346 (O_346,N_28008,N_25207);
nand UO_347 (O_347,N_27270,N_27514);
xnor UO_348 (O_348,N_29993,N_27002);
and UO_349 (O_349,N_26372,N_25592);
or UO_350 (O_350,N_28637,N_28766);
nor UO_351 (O_351,N_27121,N_29001);
nor UO_352 (O_352,N_28487,N_28400);
xor UO_353 (O_353,N_27255,N_26463);
and UO_354 (O_354,N_28364,N_29950);
xor UO_355 (O_355,N_28696,N_28306);
xnor UO_356 (O_356,N_29171,N_28898);
nor UO_357 (O_357,N_27023,N_27141);
xnor UO_358 (O_358,N_26586,N_29653);
and UO_359 (O_359,N_26488,N_26192);
and UO_360 (O_360,N_25967,N_27118);
or UO_361 (O_361,N_28184,N_29502);
xor UO_362 (O_362,N_25067,N_26261);
xnor UO_363 (O_363,N_28212,N_25685);
or UO_364 (O_364,N_27779,N_26537);
nand UO_365 (O_365,N_26330,N_29213);
or UO_366 (O_366,N_29286,N_28015);
nor UO_367 (O_367,N_26065,N_26503);
xnor UO_368 (O_368,N_29009,N_29401);
nor UO_369 (O_369,N_25491,N_27312);
nor UO_370 (O_370,N_28372,N_29398);
or UO_371 (O_371,N_25367,N_28654);
nor UO_372 (O_372,N_28190,N_25721);
and UO_373 (O_373,N_26061,N_27172);
nor UO_374 (O_374,N_26357,N_25471);
xor UO_375 (O_375,N_29240,N_27943);
and UO_376 (O_376,N_27930,N_29563);
nor UO_377 (O_377,N_25292,N_29773);
or UO_378 (O_378,N_26874,N_29890);
and UO_379 (O_379,N_25435,N_27585);
nand UO_380 (O_380,N_29520,N_25420);
or UO_381 (O_381,N_25350,N_27272);
nor UO_382 (O_382,N_28936,N_28767);
and UO_383 (O_383,N_25825,N_25999);
nand UO_384 (O_384,N_25608,N_29438);
nor UO_385 (O_385,N_25272,N_26435);
xnor UO_386 (O_386,N_29302,N_29325);
nor UO_387 (O_387,N_27459,N_26591);
or UO_388 (O_388,N_26230,N_27005);
and UO_389 (O_389,N_26185,N_29370);
xor UO_390 (O_390,N_26797,N_26922);
or UO_391 (O_391,N_25412,N_26184);
nor UO_392 (O_392,N_25762,N_29124);
nand UO_393 (O_393,N_29986,N_28350);
nand UO_394 (O_394,N_25591,N_26988);
or UO_395 (O_395,N_27479,N_26509);
nand UO_396 (O_396,N_27778,N_25278);
xor UO_397 (O_397,N_25360,N_28411);
and UO_398 (O_398,N_29580,N_26387);
xnor UO_399 (O_399,N_25180,N_27699);
nor UO_400 (O_400,N_27442,N_25906);
xor UO_401 (O_401,N_25843,N_29461);
and UO_402 (O_402,N_28847,N_25240);
or UO_403 (O_403,N_29256,N_27391);
or UO_404 (O_404,N_29193,N_27115);
nor UO_405 (O_405,N_26173,N_27196);
or UO_406 (O_406,N_27648,N_26821);
xnor UO_407 (O_407,N_29799,N_26873);
nand UO_408 (O_408,N_27792,N_25198);
and UO_409 (O_409,N_29684,N_25988);
and UO_410 (O_410,N_29641,N_29886);
xor UO_411 (O_411,N_26491,N_27161);
nor UO_412 (O_412,N_28475,N_29720);
nor UO_413 (O_413,N_27148,N_26978);
xor UO_414 (O_414,N_25324,N_29625);
nand UO_415 (O_415,N_28785,N_29603);
or UO_416 (O_416,N_28092,N_27614);
nor UO_417 (O_417,N_28269,N_29375);
nor UO_418 (O_418,N_28387,N_29372);
and UO_419 (O_419,N_26380,N_28683);
and UO_420 (O_420,N_25849,N_28278);
xnor UO_421 (O_421,N_29383,N_26187);
nand UO_422 (O_422,N_28752,N_26459);
nand UO_423 (O_423,N_26174,N_26803);
or UO_424 (O_424,N_26284,N_28192);
nor UO_425 (O_425,N_27765,N_29458);
nand UO_426 (O_426,N_26851,N_26216);
xor UO_427 (O_427,N_25581,N_28856);
nor UO_428 (O_428,N_29806,N_28227);
or UO_429 (O_429,N_27274,N_29770);
or UO_430 (O_430,N_26496,N_29230);
xor UO_431 (O_431,N_27244,N_27200);
nor UO_432 (O_432,N_26664,N_26188);
or UO_433 (O_433,N_28718,N_28361);
and UO_434 (O_434,N_29035,N_29687);
and UO_435 (O_435,N_28425,N_25452);
or UO_436 (O_436,N_26558,N_26840);
and UO_437 (O_437,N_26980,N_25597);
and UO_438 (O_438,N_28743,N_28878);
and UO_439 (O_439,N_27100,N_29865);
nor UO_440 (O_440,N_28773,N_25683);
or UO_441 (O_441,N_26217,N_27054);
and UO_442 (O_442,N_29711,N_27324);
xnor UO_443 (O_443,N_25784,N_27601);
xnor UO_444 (O_444,N_29092,N_28382);
and UO_445 (O_445,N_27572,N_26876);
and UO_446 (O_446,N_29811,N_29328);
or UO_447 (O_447,N_26929,N_25707);
and UO_448 (O_448,N_25866,N_28668);
or UO_449 (O_449,N_27004,N_25794);
and UO_450 (O_450,N_25912,N_28532);
and UO_451 (O_451,N_27787,N_29047);
or UO_452 (O_452,N_25810,N_26231);
nand UO_453 (O_453,N_25927,N_25383);
xor UO_454 (O_454,N_26131,N_27950);
and UO_455 (O_455,N_27224,N_29029);
or UO_456 (O_456,N_27841,N_28044);
xnor UO_457 (O_457,N_28316,N_28548);
nor UO_458 (O_458,N_26405,N_27266);
xnor UO_459 (O_459,N_27866,N_26942);
or UO_460 (O_460,N_27858,N_28941);
nand UO_461 (O_461,N_25644,N_29796);
and UO_462 (O_462,N_29490,N_28492);
nand UO_463 (O_463,N_25229,N_26798);
nand UO_464 (O_464,N_26585,N_28399);
or UO_465 (O_465,N_26319,N_27894);
or UO_466 (O_466,N_29284,N_28996);
nand UO_467 (O_467,N_28963,N_25770);
or UO_468 (O_468,N_25487,N_26244);
nand UO_469 (O_469,N_28460,N_26280);
xor UO_470 (O_470,N_26639,N_28033);
or UO_471 (O_471,N_29350,N_29142);
nor UO_472 (O_472,N_25414,N_27301);
or UO_473 (O_473,N_27719,N_25316);
or UO_474 (O_474,N_29589,N_28741);
and UO_475 (O_475,N_26916,N_28680);
nor UO_476 (O_476,N_27340,N_25647);
or UO_477 (O_477,N_28589,N_28334);
nand UO_478 (O_478,N_27209,N_25634);
nand UO_479 (O_479,N_28980,N_29150);
xor UO_480 (O_480,N_25224,N_25787);
and UO_481 (O_481,N_29879,N_29661);
and UO_482 (O_482,N_27323,N_29070);
nor UO_483 (O_483,N_29848,N_27015);
or UO_484 (O_484,N_29119,N_29554);
nor UO_485 (O_485,N_27539,N_29513);
xnor UO_486 (O_486,N_26728,N_28245);
or UO_487 (O_487,N_26292,N_26159);
xor UO_488 (O_488,N_25287,N_26671);
xnor UO_489 (O_489,N_25528,N_28757);
xnor UO_490 (O_490,N_25819,N_29576);
and UO_491 (O_491,N_25230,N_27875);
nand UO_492 (O_492,N_25380,N_27972);
and UO_493 (O_493,N_25223,N_26731);
or UO_494 (O_494,N_25494,N_29496);
nand UO_495 (O_495,N_25345,N_26609);
nor UO_496 (O_496,N_25107,N_27849);
nand UO_497 (O_497,N_27320,N_26471);
nand UO_498 (O_498,N_29169,N_28517);
and UO_499 (O_499,N_27895,N_26098);
nor UO_500 (O_500,N_29473,N_26846);
nor UO_501 (O_501,N_27638,N_27517);
and UO_502 (O_502,N_27804,N_27872);
or UO_503 (O_503,N_28329,N_28561);
and UO_504 (O_504,N_29982,N_29272);
nand UO_505 (O_505,N_28830,N_27507);
nor UO_506 (O_506,N_29249,N_29568);
or UO_507 (O_507,N_25354,N_25238);
or UO_508 (O_508,N_29449,N_25366);
and UO_509 (O_509,N_28719,N_25766);
or UO_510 (O_510,N_25746,N_26082);
xnor UO_511 (O_511,N_25054,N_25809);
nand UO_512 (O_512,N_25459,N_26074);
or UO_513 (O_513,N_25489,N_27492);
nor UO_514 (O_514,N_28821,N_27611);
and UO_515 (O_515,N_25692,N_27385);
and UO_516 (O_516,N_28169,N_28870);
xor UO_517 (O_517,N_29399,N_27887);
nor UO_518 (O_518,N_28618,N_25929);
nor UO_519 (O_519,N_27702,N_28908);
nor UO_520 (O_520,N_25417,N_26068);
nand UO_521 (O_521,N_27216,N_26358);
or UO_522 (O_522,N_25919,N_27546);
xor UO_523 (O_523,N_25916,N_27903);
nor UO_524 (O_524,N_29957,N_29888);
nor UO_525 (O_525,N_28689,N_27390);
and UO_526 (O_526,N_28215,N_29808);
or UO_527 (O_527,N_29996,N_25108);
xnor UO_528 (O_528,N_25820,N_25674);
and UO_529 (O_529,N_27046,N_27395);
or UO_530 (O_530,N_27829,N_25110);
xnor UO_531 (O_531,N_26344,N_28728);
or UO_532 (O_532,N_26038,N_25042);
xor UO_533 (O_533,N_26364,N_25057);
or UO_534 (O_534,N_26781,N_27264);
or UO_535 (O_535,N_26811,N_26580);
xnor UO_536 (O_536,N_26469,N_25605);
and UO_537 (O_537,N_26475,N_27952);
and UO_538 (O_538,N_29207,N_25318);
or UO_539 (O_539,N_28776,N_29530);
nand UO_540 (O_540,N_29798,N_26796);
xor UO_541 (O_541,N_28216,N_28328);
and UO_542 (O_542,N_27036,N_26450);
xnor UO_543 (O_543,N_29435,N_28990);
xnor UO_544 (O_544,N_28260,N_27080);
and UO_545 (O_545,N_29289,N_27551);
or UO_546 (O_546,N_26577,N_26847);
or UO_547 (O_547,N_28850,N_25547);
xnor UO_548 (O_548,N_28679,N_26741);
nor UO_549 (O_549,N_28271,N_26725);
nor UO_550 (O_550,N_28935,N_28218);
nor UO_551 (O_551,N_29535,N_26165);
or UO_552 (O_552,N_25402,N_27062);
xor UO_553 (O_553,N_27579,N_28903);
xnor UO_554 (O_554,N_29045,N_27518);
and UO_555 (O_555,N_27206,N_27597);
and UO_556 (O_556,N_29075,N_27030);
xor UO_557 (O_557,N_26498,N_27071);
nor UO_558 (O_558,N_29265,N_25983);
and UO_559 (O_559,N_29624,N_27481);
nand UO_560 (O_560,N_28347,N_26224);
and UO_561 (O_561,N_28904,N_29716);
nand UO_562 (O_562,N_27153,N_28299);
nor UO_563 (O_563,N_28452,N_26822);
and UO_564 (O_564,N_27350,N_27268);
or UO_565 (O_565,N_29882,N_25624);
nor UO_566 (O_566,N_25003,N_28154);
nand UO_567 (O_567,N_26989,N_27773);
nor UO_568 (O_568,N_27990,N_29136);
nand UO_569 (O_569,N_29157,N_25009);
or UO_570 (O_570,N_27307,N_28457);
and UO_571 (O_571,N_27985,N_28238);
xor UO_572 (O_572,N_25822,N_28084);
nor UO_573 (O_573,N_27681,N_28090);
or UO_574 (O_574,N_26281,N_25745);
xnor UO_575 (O_575,N_25753,N_26809);
nor UO_576 (O_576,N_27639,N_29276);
nor UO_577 (O_577,N_29695,N_26515);
or UO_578 (O_578,N_27379,N_29471);
or UO_579 (O_579,N_29609,N_26221);
and UO_580 (O_580,N_28619,N_25317);
nand UO_581 (O_581,N_26339,N_29783);
nand UO_582 (O_582,N_26827,N_28180);
and UO_583 (O_583,N_27330,N_25451);
nand UO_584 (O_584,N_28832,N_28765);
nor UO_585 (O_585,N_26275,N_25955);
nand UO_586 (O_586,N_26245,N_28516);
and UO_587 (O_587,N_25931,N_28229);
nor UO_588 (O_588,N_28291,N_25991);
nand UO_589 (O_589,N_27591,N_27509);
or UO_590 (O_590,N_26432,N_27060);
and UO_591 (O_591,N_25467,N_28187);
or UO_592 (O_592,N_28472,N_27339);
nand UO_593 (O_593,N_28905,N_25099);
or UO_594 (O_594,N_26913,N_27035);
or UO_595 (O_595,N_27678,N_25353);
nand UO_596 (O_596,N_27501,N_27520);
nor UO_597 (O_597,N_25264,N_27637);
nand UO_598 (O_598,N_28838,N_29163);
or UO_599 (O_599,N_25177,N_26695);
nand UO_600 (O_600,N_26454,N_27667);
and UO_601 (O_601,N_29316,N_29737);
or UO_602 (O_602,N_25294,N_29779);
and UO_603 (O_603,N_27360,N_27353);
nand UO_604 (O_604,N_29788,N_28157);
or UO_605 (O_605,N_26257,N_29300);
and UO_606 (O_606,N_29478,N_27252);
and UO_607 (O_607,N_25194,N_29836);
or UO_608 (O_608,N_25862,N_25777);
or UO_609 (O_609,N_29688,N_27968);
xor UO_610 (O_610,N_26620,N_25606);
or UO_611 (O_611,N_27784,N_25163);
or UO_612 (O_612,N_25795,N_27309);
nand UO_613 (O_613,N_29498,N_28057);
nand UO_614 (O_614,N_25243,N_27375);
xnor UO_615 (O_615,N_25860,N_26071);
or UO_616 (O_616,N_25302,N_28641);
nand UO_617 (O_617,N_25872,N_27528);
nand UO_618 (O_618,N_26675,N_27447);
xor UO_619 (O_619,N_28161,N_28810);
nor UO_620 (O_620,N_28907,N_27341);
and UO_621 (O_621,N_25846,N_25575);
nand UO_622 (O_622,N_25428,N_26701);
xnor UO_623 (O_623,N_26541,N_29214);
xnor UO_624 (O_624,N_29818,N_28684);
nand UO_625 (O_625,N_25058,N_25650);
nand UO_626 (O_626,N_27901,N_29784);
nand UO_627 (O_627,N_29416,N_28792);
nor UO_628 (O_628,N_26593,N_29935);
and UO_629 (O_629,N_26802,N_29983);
nand UO_630 (O_630,N_27130,N_27851);
nand UO_631 (O_631,N_27256,N_29523);
nor UO_632 (O_632,N_27451,N_25758);
nand UO_633 (O_633,N_27586,N_25456);
nor UO_634 (O_634,N_25691,N_26154);
and UO_635 (O_635,N_29948,N_28099);
nor UO_636 (O_636,N_25079,N_29103);
xnor UO_637 (O_637,N_28011,N_29614);
xnor UO_638 (O_638,N_25598,N_26683);
nor UO_639 (O_639,N_28040,N_27708);
and UO_640 (O_640,N_27410,N_28071);
or UO_641 (O_641,N_29156,N_28262);
or UO_642 (O_642,N_29852,N_25541);
or UO_643 (O_643,N_27558,N_27782);
nor UO_644 (O_644,N_27836,N_26136);
nor UO_645 (O_645,N_29094,N_25994);
nor UO_646 (O_646,N_25045,N_29422);
nor UO_647 (O_647,N_29087,N_25868);
nand UO_648 (O_648,N_25725,N_28899);
xor UO_649 (O_649,N_26133,N_29714);
nor UO_650 (O_650,N_28761,N_27247);
and UO_651 (O_651,N_28606,N_25464);
nand UO_652 (O_652,N_26879,N_28285);
xor UO_653 (O_653,N_27559,N_28603);
nand UO_654 (O_654,N_25728,N_28572);
or UO_655 (O_655,N_26777,N_28482);
nand UO_656 (O_656,N_28913,N_27478);
or UO_657 (O_657,N_27703,N_26891);
and UO_658 (O_658,N_27664,N_27242);
or UO_659 (O_659,N_28222,N_25378);
nor UO_660 (O_660,N_27189,N_27821);
xnor UO_661 (O_661,N_25633,N_29956);
nand UO_662 (O_662,N_27781,N_27364);
nor UO_663 (O_663,N_25673,N_28474);
nand UO_664 (O_664,N_27863,N_27902);
xor UO_665 (O_665,N_25217,N_29220);
nor UO_666 (O_666,N_26239,N_28636);
or UO_667 (O_667,N_27081,N_29729);
or UO_668 (O_668,N_28458,N_29476);
nor UO_669 (O_669,N_28078,N_29089);
or UO_670 (O_670,N_27214,N_27218);
and UO_671 (O_671,N_27310,N_28822);
xnor UO_672 (O_672,N_26012,N_26921);
xnor UO_673 (O_673,N_26138,N_29529);
xnor UO_674 (O_674,N_29288,N_26700);
xor UO_675 (O_675,N_26703,N_25001);
and UO_676 (O_676,N_26323,N_25583);
or UO_677 (O_677,N_25299,N_29987);
xnor UO_678 (O_678,N_28272,N_26977);
and UO_679 (O_679,N_28403,N_29268);
nor UO_680 (O_680,N_27652,N_29279);
and UO_681 (O_681,N_29178,N_25157);
or UO_682 (O_682,N_27622,N_25393);
nand UO_683 (O_683,N_26861,N_27026);
nand UO_684 (O_684,N_28193,N_29273);
nor UO_685 (O_685,N_29778,N_29851);
nand UO_686 (O_686,N_27229,N_27131);
and UO_687 (O_687,N_29651,N_29048);
and UO_688 (O_688,N_25760,N_25181);
and UO_689 (O_689,N_26333,N_27549);
or UO_690 (O_690,N_28900,N_26276);
nand UO_691 (O_691,N_25200,N_26287);
xnor UO_692 (O_692,N_25710,N_26583);
and UO_693 (O_693,N_27124,N_25614);
xor UO_694 (O_694,N_26113,N_28539);
nand UO_695 (O_695,N_27623,N_29750);
nand UO_696 (O_696,N_28281,N_26838);
or UO_697 (O_697,N_29320,N_28496);
nand UO_698 (O_698,N_25164,N_25499);
and UO_699 (O_699,N_28435,N_25347);
nand UO_700 (O_700,N_29385,N_25965);
or UO_701 (O_701,N_28709,N_25922);
and UO_702 (O_702,N_25642,N_27333);
nor UO_703 (O_703,N_27629,N_27565);
xnor UO_704 (O_704,N_29062,N_29980);
or UO_705 (O_705,N_26197,N_25472);
nand UO_706 (O_706,N_26274,N_28800);
nand UO_707 (O_707,N_29738,N_28727);
xnor UO_708 (O_708,N_28536,N_25112);
nand UO_709 (O_709,N_27802,N_28813);
and UO_710 (O_710,N_28988,N_27830);
xnor UO_711 (O_711,N_28700,N_27896);
and UO_712 (O_712,N_29474,N_27351);
nor UO_713 (O_713,N_29510,N_25959);
nand UO_714 (O_714,N_25565,N_26409);
or UO_715 (O_715,N_29448,N_25138);
or UO_716 (O_716,N_29825,N_29710);
nand UO_717 (O_717,N_25358,N_28910);
nand UO_718 (O_718,N_29348,N_27662);
and UO_719 (O_719,N_26660,N_29894);
nor UO_720 (O_720,N_28836,N_26645);
or UO_721 (O_721,N_29718,N_25185);
nand UO_722 (O_722,N_26451,N_27711);
or UO_723 (O_723,N_28942,N_25697);
nand UO_724 (O_724,N_28043,N_27571);
or UO_725 (O_725,N_26016,N_28646);
or UO_726 (O_726,N_25661,N_28060);
xnor UO_727 (O_727,N_28294,N_27359);
or UO_728 (O_728,N_27191,N_29292);
or UO_729 (O_729,N_28498,N_28415);
nor UO_730 (O_730,N_25530,N_25568);
nor UO_731 (O_731,N_25369,N_26397);
and UO_732 (O_732,N_27354,N_29924);
nand UO_733 (O_733,N_26559,N_27521);
nand UO_734 (O_734,N_25826,N_27824);
nor UO_735 (O_735,N_28164,N_25087);
xnor UO_736 (O_736,N_27644,N_28231);
nor UO_737 (O_737,N_29054,N_25663);
nand UO_738 (O_738,N_29139,N_26857);
nor UO_739 (O_739,N_28928,N_26831);
and UO_740 (O_740,N_26758,N_29777);
and UO_741 (O_741,N_26142,N_29713);
nand UO_742 (O_742,N_26293,N_27966);
nand UO_743 (O_743,N_26628,N_27331);
nor UO_744 (O_744,N_29447,N_27495);
or UO_745 (O_745,N_28537,N_29442);
nand UO_746 (O_746,N_25643,N_25684);
or UO_747 (O_747,N_27877,N_29795);
nor UO_748 (O_748,N_27232,N_26321);
xnor UO_749 (O_749,N_29828,N_28805);
xnor UO_750 (O_750,N_26682,N_29578);
nor UO_751 (O_751,N_25029,N_26264);
or UO_752 (O_752,N_26880,N_29334);
and UO_753 (O_753,N_25469,N_26707);
and UO_754 (O_754,N_29364,N_29967);
nand UO_755 (O_755,N_28236,N_28448);
and UO_756 (O_756,N_26562,N_26072);
nand UO_757 (O_757,N_29897,N_29377);
nor UO_758 (O_758,N_25395,N_28775);
xor UO_759 (O_759,N_26359,N_29427);
xor UO_760 (O_760,N_26853,N_26729);
and UO_761 (O_761,N_27421,N_27722);
xor UO_762 (O_762,N_26764,N_25847);
nor UO_763 (O_763,N_29757,N_25429);
or UO_764 (O_764,N_29161,N_29072);
nand UO_765 (O_765,N_26169,N_25559);
or UO_766 (O_766,N_29120,N_27498);
nand UO_767 (O_767,N_29412,N_25159);
xor UO_768 (O_768,N_26856,N_25134);
and UO_769 (O_769,N_26298,N_28534);
nand UO_770 (O_770,N_26044,N_29140);
nand UO_771 (O_771,N_28095,N_25073);
nand UO_772 (O_772,N_28233,N_27910);
or UO_773 (O_773,N_27777,N_25094);
nor UO_774 (O_774,N_28055,N_27612);
and UO_775 (O_775,N_28346,N_29123);
nand UO_776 (O_776,N_29912,N_29867);
xnor UO_777 (O_777,N_25176,N_25904);
nand UO_778 (O_778,N_29246,N_27690);
and UO_779 (O_779,N_26767,N_25124);
xnor UO_780 (O_780,N_27796,N_29514);
xnor UO_781 (O_781,N_28443,N_26543);
xor UO_782 (O_782,N_25083,N_28148);
xnor UO_783 (O_783,N_26347,N_25646);
and UO_784 (O_784,N_29507,N_27055);
nor UO_785 (O_785,N_29199,N_25375);
nand UO_786 (O_786,N_28254,N_27944);
xnor UO_787 (O_787,N_25715,N_29405);
nor UO_788 (O_788,N_27488,N_26105);
and UO_789 (O_789,N_26933,N_29922);
or UO_790 (O_790,N_29932,N_28143);
or UO_791 (O_791,N_29112,N_27746);
xor UO_792 (O_792,N_26968,N_28648);
nor UO_793 (O_793,N_27604,N_27860);
nor UO_794 (O_794,N_25298,N_27223);
or UO_795 (O_795,N_27908,N_25047);
nand UO_796 (O_796,N_25717,N_29105);
xor UO_797 (O_797,N_27464,N_28750);
nand UO_798 (O_798,N_29637,N_29822);
or UO_799 (O_799,N_27136,N_25468);
or UO_800 (O_800,N_26548,N_25567);
xnor UO_801 (O_801,N_28897,N_28429);
nor UO_802 (O_802,N_27856,N_26189);
xor UO_803 (O_803,N_25109,N_28630);
or UO_804 (O_804,N_29844,N_28787);
or UO_805 (O_805,N_25720,N_26427);
xnor UO_806 (O_806,N_29512,N_27032);
nor UO_807 (O_807,N_28451,N_25455);
nand UO_808 (O_808,N_28333,N_29457);
nand UO_809 (O_809,N_26776,N_27596);
xor UO_810 (O_810,N_27091,N_26511);
and UO_811 (O_811,N_29341,N_29080);
nor UO_812 (O_812,N_27424,N_29132);
nor UO_813 (O_813,N_29303,N_25286);
or UO_814 (O_814,N_29146,N_26346);
xor UO_815 (O_815,N_25144,N_29137);
and UO_816 (O_816,N_29203,N_25448);
and UO_817 (O_817,N_25884,N_27991);
nand UO_818 (O_818,N_26519,N_25191);
xor UO_819 (O_819,N_28879,N_25327);
or UO_820 (O_820,N_27534,N_27476);
xor UO_821 (O_821,N_26440,N_28153);
and UO_822 (O_822,N_29313,N_26448);
and UO_823 (O_823,N_26866,N_26975);
xor UO_824 (O_824,N_26640,N_28030);
or UO_825 (O_825,N_29955,N_29701);
nand UO_826 (O_826,N_27813,N_25797);
nand UO_827 (O_827,N_28356,N_25012);
nand UO_828 (O_828,N_26708,N_29934);
xnor UO_829 (O_829,N_27914,N_27095);
or UO_830 (O_830,N_26594,N_28438);
nor UO_831 (O_831,N_27446,N_26756);
and UO_832 (O_832,N_25371,N_26834);
nor UO_833 (O_833,N_26115,N_29730);
nor UO_834 (O_834,N_26236,N_27029);
and UO_835 (O_835,N_29402,N_28027);
or UO_836 (O_836,N_25093,N_29491);
xnor UO_837 (O_837,N_25145,N_28286);
or UO_838 (O_838,N_29371,N_27785);
xnor UO_839 (O_839,N_29915,N_26297);
xor UO_840 (O_840,N_27885,N_29634);
and UO_841 (O_841,N_25801,N_25311);
and UO_842 (O_842,N_25065,N_26304);
or UO_843 (O_843,N_26623,N_27017);
or UO_844 (O_844,N_28314,N_27380);
nor UO_845 (O_845,N_27342,N_29319);
nand UO_846 (O_846,N_28440,N_25792);
nor UO_847 (O_847,N_25082,N_25517);
nor UO_848 (O_848,N_29440,N_26926);
nand UO_849 (O_849,N_28158,N_25686);
or UO_850 (O_850,N_28527,N_29919);
and UO_851 (O_851,N_25926,N_27291);
and UO_852 (O_852,N_29400,N_27941);
nand UO_853 (O_853,N_28163,N_28807);
or UO_854 (O_854,N_28114,N_27971);
nand UO_855 (O_855,N_26806,N_27590);
xor UO_856 (O_856,N_27150,N_26286);
or UO_857 (O_857,N_27625,N_26787);
and UO_858 (O_858,N_27831,N_26947);
nor UO_859 (O_859,N_26644,N_25284);
and UO_860 (O_860,N_28713,N_29861);
or UO_861 (O_861,N_26552,N_27808);
and UO_862 (O_862,N_27097,N_25115);
or UO_863 (O_863,N_29236,N_26992);
nand UO_864 (O_864,N_28645,N_28270);
xor UO_865 (O_865,N_27185,N_26597);
nor UO_866 (O_866,N_27940,N_29098);
or UO_867 (O_867,N_25601,N_25326);
nand UO_868 (O_868,N_28477,N_28541);
and UO_869 (O_869,N_26370,N_29305);
and UO_870 (O_870,N_26900,N_27021);
nand UO_871 (O_871,N_25245,N_26748);
or UO_872 (O_872,N_29441,N_25492);
or UO_873 (O_873,N_25823,N_25562);
nand UO_874 (O_874,N_28771,N_29928);
xnor UO_875 (O_875,N_25538,N_26958);
and UO_876 (O_876,N_29782,N_25063);
xor UO_877 (O_877,N_26058,N_25905);
xor UO_878 (O_878,N_28712,N_27513);
nand UO_879 (O_879,N_26869,N_28651);
and UO_880 (O_880,N_26107,N_25274);
nand UO_881 (O_881,N_26166,N_27182);
nand UO_882 (O_882,N_26130,N_29832);
or UO_883 (O_883,N_28967,N_27730);
or UO_884 (O_884,N_26027,N_26542);
and UO_885 (O_885,N_25102,N_27105);
nand UO_886 (O_886,N_28702,N_27282);
nor UO_887 (O_887,N_27790,N_29805);
xor UO_888 (O_888,N_25027,N_29843);
or UO_889 (O_889,N_28845,N_26727);
nand UO_890 (O_890,N_28715,N_26234);
nand UO_891 (O_891,N_27336,N_26085);
xor UO_892 (O_892,N_26049,N_26124);
nand UO_893 (O_893,N_28330,N_28051);
nand UO_894 (O_894,N_25966,N_25266);
nand UO_895 (O_895,N_26737,N_26407);
nor UO_896 (O_896,N_27705,N_29964);
and UO_897 (O_897,N_29864,N_28100);
nor UO_898 (O_898,N_27373,N_26400);
or UO_899 (O_899,N_29582,N_26676);
or UO_900 (O_900,N_25434,N_26792);
or UO_901 (O_901,N_28473,N_25930);
and UO_902 (O_902,N_29537,N_26872);
nor UO_903 (O_903,N_28433,N_28755);
xor UO_904 (O_904,N_28778,N_27634);
xor UO_905 (O_905,N_28103,N_26480);
nand UO_906 (O_906,N_29753,N_28505);
xnor UO_907 (O_907,N_26500,N_25519);
nor UO_908 (O_908,N_29675,N_27134);
xor UO_909 (O_909,N_25234,N_26260);
nand UO_910 (O_910,N_26249,N_29174);
nand UO_911 (O_911,N_29763,N_25343);
xor UO_912 (O_912,N_28063,N_26393);
and UO_913 (O_913,N_29264,N_25152);
nor UO_914 (O_914,N_25869,N_25791);
or UO_915 (O_915,N_26070,N_29262);
xor UO_916 (O_916,N_25678,N_26093);
xnor UO_917 (O_917,N_25019,N_25533);
xor UO_918 (O_918,N_29775,N_28797);
and UO_919 (O_919,N_26904,N_26976);
or UO_920 (O_920,N_28660,N_28968);
and UO_921 (O_921,N_26110,N_28405);
and UO_922 (O_922,N_29183,N_28769);
or UO_923 (O_923,N_25213,N_29198);
xnor UO_924 (O_924,N_29152,N_25704);
nand UO_925 (O_925,N_25091,N_25397);
nor UO_926 (O_926,N_25811,N_26483);
xor UO_927 (O_927,N_26871,N_25893);
xnor UO_928 (O_928,N_26538,N_29309);
or UO_929 (O_929,N_29382,N_29837);
and UO_930 (O_930,N_27493,N_25622);
xnor UO_931 (O_931,N_28786,N_29715);
nor UO_932 (O_932,N_29042,N_28037);
nor UO_933 (O_933,N_26114,N_28507);
nand UO_934 (O_934,N_25329,N_25485);
xnor UO_935 (O_935,N_25000,N_28986);
and UO_936 (O_936,N_27453,N_26885);
and UO_937 (O_937,N_25219,N_28951);
nand UO_938 (O_938,N_29989,N_27494);
xnor UO_939 (O_939,N_29518,N_27089);
nor UO_940 (O_940,N_25314,N_29467);
or UO_941 (O_941,N_29943,N_28029);
xor UO_942 (O_942,N_28552,N_27527);
nor UO_943 (O_943,N_28688,N_26650);
and UO_944 (O_944,N_25405,N_25956);
and UO_945 (O_945,N_25232,N_27396);
and UO_946 (O_946,N_25004,N_26715);
xnor UO_947 (O_947,N_26171,N_29034);
and UO_948 (O_948,N_28609,N_25129);
xor UO_949 (O_949,N_26522,N_27530);
xor UO_950 (O_950,N_26078,N_26898);
and UO_951 (O_951,N_26366,N_29085);
nor UO_952 (O_952,N_25017,N_27415);
nor UO_953 (O_953,N_27348,N_28803);
and UO_954 (O_954,N_27429,N_25750);
nand UO_955 (O_955,N_25914,N_26832);
or UO_956 (O_956,N_27606,N_26556);
and UO_957 (O_957,N_25014,N_28257);
or UO_958 (O_958,N_29357,N_27438);
and UO_959 (O_959,N_26163,N_28120);
or UO_960 (O_960,N_25236,N_27031);
xnor UO_961 (O_961,N_29433,N_25989);
and UO_962 (O_962,N_27014,N_25935);
nand UO_963 (O_963,N_28626,N_25563);
and UO_964 (O_964,N_26722,N_26026);
nor UO_965 (O_965,N_27110,N_28714);
nor UO_966 (O_966,N_29631,N_28804);
or UO_967 (O_967,N_26884,N_25253);
and UO_968 (O_968,N_28461,N_27798);
and UO_969 (O_969,N_26967,N_27407);
xor UO_970 (O_970,N_25602,N_28025);
nor UO_971 (O_971,N_26076,N_28602);
xor UO_972 (O_972,N_27432,N_25590);
nor UO_973 (O_973,N_29977,N_25986);
xnor UO_974 (O_974,N_26740,N_29116);
nor UO_975 (O_975,N_26908,N_28739);
nor UO_976 (O_976,N_27305,N_29218);
nand UO_977 (O_977,N_25752,N_27598);
and UO_978 (O_978,N_29920,N_27911);
xnor UO_979 (O_979,N_27855,N_29380);
nor UO_980 (O_980,N_26006,N_27961);
or UO_981 (O_981,N_25237,N_25359);
and UO_982 (O_982,N_27696,N_27203);
and UO_983 (O_983,N_25993,N_27152);
nor UO_984 (O_984,N_29281,N_26972);
nand UO_985 (O_985,N_25104,N_26457);
nor UO_986 (O_986,N_28675,N_29940);
nand UO_987 (O_987,N_26329,N_29672);
nor UO_988 (O_988,N_26532,N_26351);
xnor UO_989 (O_989,N_27684,N_25162);
or UO_990 (O_990,N_29658,N_25418);
or UO_991 (O_991,N_29542,N_27490);
nand UO_992 (O_992,N_27186,N_28002);
nor UO_993 (O_993,N_28122,N_25478);
nor UO_994 (O_994,N_27006,N_25473);
xor UO_995 (O_995,N_26215,N_29762);
or UO_996 (O_996,N_29133,N_27717);
nand UO_997 (O_997,N_26844,N_28664);
nor UO_998 (O_998,N_27416,N_27466);
nand UO_999 (O_999,N_28578,N_28895);
or UO_1000 (O_1000,N_28431,N_27632);
and UO_1001 (O_1001,N_28397,N_29764);
or UO_1002 (O_1002,N_26069,N_27733);
and UO_1003 (O_1003,N_26377,N_29244);
xnor UO_1004 (O_1004,N_27868,N_28737);
nor UO_1005 (O_1005,N_25431,N_25249);
nand UO_1006 (O_1006,N_25463,N_26429);
xor UO_1007 (O_1007,N_29068,N_27241);
or UO_1008 (O_1008,N_26763,N_28983);
xor UO_1009 (O_1009,N_28932,N_26575);
or UO_1010 (O_1010,N_29887,N_26652);
nor UO_1011 (O_1011,N_25892,N_28808);
or UO_1012 (O_1012,N_29148,N_27962);
nand UO_1013 (O_1013,N_29434,N_27988);
or UO_1014 (O_1014,N_29165,N_29809);
nand UO_1015 (O_1015,N_27254,N_27117);
nand UO_1016 (O_1016,N_27837,N_28697);
nand UO_1017 (O_1017,N_27775,N_29311);
nor UO_1018 (O_1018,N_28600,N_27240);
nand UO_1019 (O_1019,N_25695,N_26472);
or UO_1020 (O_1020,N_28389,N_29074);
or UO_1021 (O_1021,N_26320,N_29071);
or UO_1022 (O_1022,N_29748,N_29059);
xor UO_1023 (O_1023,N_25074,N_28851);
xor UO_1024 (O_1024,N_26334,N_27603);
nor UO_1025 (O_1025,N_27801,N_28097);
xnor UO_1026 (O_1026,N_27251,N_27732);
xnor UO_1027 (O_1027,N_28146,N_27132);
and UO_1028 (O_1028,N_26041,N_29959);
nand UO_1029 (O_1029,N_25192,N_29114);
nor UO_1030 (O_1030,N_25031,N_28650);
nor UO_1031 (O_1031,N_29786,N_25793);
nand UO_1032 (O_1032,N_26897,N_25049);
nor UO_1033 (O_1033,N_26973,N_28565);
and UO_1034 (O_1034,N_28243,N_27915);
nor UO_1035 (O_1035,N_29880,N_25896);
nand UO_1036 (O_1036,N_26621,N_25969);
nor UO_1037 (O_1037,N_25400,N_27231);
or UO_1038 (O_1038,N_27674,N_25688);
or UO_1039 (O_1039,N_28888,N_28348);
nor UO_1040 (O_1040,N_25553,N_29553);
or UO_1041 (O_1041,N_28605,N_28220);
nor UO_1042 (O_1042,N_26587,N_27145);
and UO_1043 (O_1043,N_28999,N_26028);
nor UO_1044 (O_1044,N_26529,N_27092);
nor UO_1045 (O_1045,N_27651,N_25290);
xnor UO_1046 (O_1046,N_29361,N_29745);
xor UO_1047 (O_1047,N_28098,N_27388);
xor UO_1048 (O_1048,N_28514,N_28484);
nor UO_1049 (O_1049,N_28758,N_27174);
nand UO_1050 (O_1050,N_29823,N_26914);
nor UO_1051 (O_1051,N_25204,N_29925);
and UO_1052 (O_1052,N_26111,N_25018);
nand UO_1053 (O_1053,N_26805,N_25948);
xor UO_1054 (O_1054,N_29395,N_29049);
xnor UO_1055 (O_1055,N_26151,N_29223);
and UO_1056 (O_1056,N_25903,N_28528);
xor UO_1057 (O_1057,N_29958,N_26505);
or UO_1058 (O_1058,N_28625,N_27001);
nor UO_1059 (O_1059,N_28873,N_26120);
nand UO_1060 (O_1060,N_25726,N_28105);
nand UO_1061 (O_1061,N_28911,N_27126);
and UO_1062 (O_1062,N_28882,N_27289);
and UO_1063 (O_1063,N_26813,N_26101);
or UO_1064 (O_1064,N_27047,N_26388);
xnor UO_1065 (O_1065,N_26778,N_25626);
or UO_1066 (O_1066,N_29627,N_26145);
or UO_1067 (O_1067,N_26455,N_29642);
xor UO_1068 (O_1068,N_26546,N_29037);
and UO_1069 (O_1069,N_28145,N_27083);
nor UO_1070 (O_1070,N_28196,N_29562);
or UO_1071 (O_1071,N_29746,N_26812);
or UO_1072 (O_1072,N_29657,N_28647);
xor UO_1073 (O_1073,N_28593,N_25007);
nor UO_1074 (O_1074,N_25982,N_25500);
nand UO_1075 (O_1075,N_26833,N_26443);
nand UO_1076 (O_1076,N_28638,N_29628);
or UO_1077 (O_1077,N_28332,N_28469);
or UO_1078 (O_1078,N_26956,N_26653);
or UO_1079 (O_1079,N_28842,N_25952);
nor UO_1080 (O_1080,N_28659,N_27965);
and UO_1081 (O_1081,N_29482,N_26673);
or UO_1082 (O_1082,N_27075,N_25888);
xor UO_1083 (O_1083,N_28760,N_27883);
or UO_1084 (O_1084,N_29991,N_27455);
or UO_1085 (O_1085,N_28952,N_25557);
or UO_1086 (O_1086,N_28909,N_27553);
xnor UO_1087 (O_1087,N_25790,N_28230);
nor UO_1088 (O_1088,N_26750,N_29509);
nand UO_1089 (O_1089,N_29531,N_28047);
or UO_1090 (O_1090,N_26019,N_25623);
nand UO_1091 (O_1091,N_27954,N_25158);
and UO_1092 (O_1092,N_25671,N_27567);
or UO_1093 (O_1093,N_29175,N_26118);
and UO_1094 (O_1094,N_26147,N_25268);
nand UO_1095 (O_1095,N_25743,N_29517);
nor UO_1096 (O_1096,N_26934,N_27710);
and UO_1097 (O_1097,N_25887,N_27052);
xor UO_1098 (O_1098,N_28160,N_28209);
nor UO_1099 (O_1099,N_27022,N_26494);
xnor UO_1100 (O_1100,N_29549,N_27960);
nand UO_1101 (O_1101,N_28574,N_29921);
or UO_1102 (O_1102,N_25540,N_26536);
and UO_1103 (O_1103,N_26307,N_26337);
or UO_1104 (O_1104,N_28510,N_29685);
and UO_1105 (O_1105,N_28530,N_27328);
nand UO_1106 (O_1106,N_29439,N_28375);
nor UO_1107 (O_1107,N_27864,N_27738);
or UO_1108 (O_1108,N_28295,N_29640);
nor UO_1109 (O_1109,N_29501,N_25594);
or UO_1110 (O_1110,N_27752,N_29906);
and UO_1111 (O_1111,N_26681,N_25220);
nor UO_1112 (O_1112,N_28189,N_29960);
xnor UO_1113 (O_1113,N_27526,N_28094);
nor UO_1114 (O_1114,N_28616,N_28009);
and UO_1115 (O_1115,N_27299,N_25356);
nand UO_1116 (O_1116,N_29069,N_28276);
nand UO_1117 (O_1117,N_29397,N_29754);
or UO_1118 (O_1118,N_29511,N_25377);
xnor UO_1119 (O_1119,N_29212,N_28449);
or UO_1120 (O_1120,N_25641,N_26421);
and UO_1121 (O_1121,N_27706,N_29310);
nand UO_1122 (O_1122,N_27828,N_25960);
nor UO_1123 (O_1123,N_29006,N_28358);
nor UO_1124 (O_1124,N_25466,N_29301);
nand UO_1125 (O_1125,N_27536,N_29002);
nor UO_1126 (O_1126,N_26312,N_28724);
nor UO_1127 (O_1127,N_28901,N_26031);
or UO_1128 (O_1128,N_25423,N_25767);
xnor UO_1129 (O_1129,N_28149,N_28862);
xor UO_1130 (O_1130,N_26545,N_29846);
xor UO_1131 (O_1131,N_29113,N_25008);
nor UO_1132 (O_1132,N_27958,N_29469);
nor UO_1133 (O_1133,N_29905,N_25558);
nand UO_1134 (O_1134,N_25453,N_26974);
nand UO_1135 (O_1135,N_29004,N_29018);
nand UO_1136 (O_1136,N_26931,N_25512);
nand UO_1137 (O_1137,N_28846,N_27982);
nor UO_1138 (O_1138,N_28077,N_26484);
xor UO_1139 (O_1139,N_25837,N_27398);
xor UO_1140 (O_1140,N_26819,N_28573);
and UO_1141 (O_1141,N_25462,N_29839);
or UO_1142 (O_1142,N_25920,N_28814);
or UO_1143 (O_1143,N_26852,N_27404);
or UO_1144 (O_1144,N_29138,N_27619);
and UO_1145 (O_1145,N_27262,N_27610);
xnor UO_1146 (O_1146,N_26134,N_29083);
nand UO_1147 (O_1147,N_28302,N_25915);
and UO_1148 (O_1148,N_27302,N_26362);
nor UO_1149 (O_1149,N_28998,N_27989);
nand UO_1150 (O_1150,N_29984,N_27448);
and UO_1151 (O_1151,N_28994,N_29875);
nand UO_1152 (O_1152,N_27165,N_28521);
nor UO_1153 (O_1153,N_27907,N_29086);
nor UO_1154 (O_1154,N_25078,N_26176);
or UO_1155 (O_1155,N_27757,N_25415);
nor UO_1156 (O_1156,N_25580,N_26924);
nor UO_1157 (O_1157,N_28424,N_25665);
nand UO_1158 (O_1158,N_28685,N_29429);
nand UO_1159 (O_1159,N_29290,N_28107);
xnor UO_1160 (O_1160,N_27334,N_29853);
xnor UO_1161 (O_1161,N_29566,N_26474);
nand UO_1162 (O_1162,N_26709,N_26571);
and UO_1163 (O_1163,N_25942,N_27347);
or UO_1164 (O_1164,N_25038,N_26962);
and UO_1165 (O_1165,N_27891,N_26618);
and UO_1166 (O_1166,N_28639,N_25084);
and UO_1167 (O_1167,N_28974,N_25842);
xor UO_1168 (O_1168,N_29079,N_27011);
nand UO_1169 (O_1169,N_25330,N_25882);
xnor UO_1170 (O_1170,N_26003,N_27955);
or UO_1171 (O_1171,N_28919,N_26446);
and UO_1172 (O_1172,N_27660,N_29944);
and UO_1173 (O_1173,N_29012,N_26691);
xnor UO_1174 (O_1174,N_28501,N_25028);
nor UO_1175 (O_1175,N_28894,N_27780);
or UO_1176 (O_1176,N_29296,N_25778);
and UO_1177 (O_1177,N_26222,N_25586);
and UO_1178 (O_1178,N_28955,N_25187);
xnor UO_1179 (O_1179,N_29063,N_25838);
xnor UO_1180 (O_1180,N_26724,N_28374);
nand UO_1181 (O_1181,N_29662,N_26990);
nor UO_1182 (O_1182,N_27233,N_28327);
and UO_1183 (O_1183,N_27861,N_29831);
and UO_1184 (O_1184,N_29810,N_26547);
xor UO_1185 (O_1185,N_28038,N_26774);
nor UO_1186 (O_1186,N_29158,N_29733);
nand UO_1187 (O_1187,N_27937,N_25430);
nand UO_1188 (O_1188,N_25781,N_28132);
or UO_1189 (O_1189,N_29263,N_29602);
nand UO_1190 (O_1190,N_28263,N_28412);
nor UO_1191 (O_1191,N_29250,N_26674);
or UO_1192 (O_1192,N_29821,N_25632);
xnor UO_1193 (O_1193,N_29797,N_27675);
nand UO_1194 (O_1194,N_28275,N_28780);
or UO_1195 (O_1195,N_26273,N_29953);
and UO_1196 (O_1196,N_29780,N_29842);
and UO_1197 (O_1197,N_29721,N_26196);
and UO_1198 (O_1198,N_29443,N_25840);
or UO_1199 (O_1199,N_26108,N_25813);
or UO_1200 (O_1200,N_28770,N_25874);
nor UO_1201 (O_1201,N_29393,N_25701);
nand UO_1202 (O_1202,N_26422,N_25907);
and UO_1203 (O_1203,N_27642,N_26353);
or UO_1204 (O_1204,N_26946,N_29287);
nor UO_1205 (O_1205,N_28995,N_29480);
or UO_1206 (O_1206,N_26228,N_29061);
xor UO_1207 (O_1207,N_27419,N_25974);
nor UO_1208 (O_1208,N_28731,N_29965);
nand UO_1209 (O_1209,N_27755,N_27679);
xor UO_1210 (O_1210,N_26526,N_28118);
and UO_1211 (O_1211,N_27484,N_28258);
xor UO_1212 (O_1212,N_27898,N_29494);
or UO_1213 (O_1213,N_25498,N_27689);
xnor UO_1214 (O_1214,N_28056,N_25066);
or UO_1215 (O_1215,N_26227,N_28106);
and UO_1216 (O_1216,N_26678,N_25062);
nand UO_1217 (O_1217,N_29426,N_29209);
and UO_1218 (O_1218,N_26994,N_28138);
xnor UO_1219 (O_1219,N_28385,N_28756);
nand UO_1220 (O_1220,N_26434,N_26395);
nand UO_1221 (O_1221,N_28710,N_29691);
or UO_1222 (O_1222,N_29506,N_29437);
and UO_1223 (O_1223,N_29612,N_26206);
nand UO_1224 (O_1224,N_25437,N_29466);
xnor UO_1225 (O_1225,N_27367,N_26300);
or UO_1226 (O_1226,N_26601,N_26859);
xor UO_1227 (O_1227,N_29638,N_26721);
or UO_1228 (O_1228,N_27540,N_28535);
or UO_1229 (O_1229,N_25579,N_27980);
nor UO_1230 (O_1230,N_26327,N_25121);
nand UO_1231 (O_1231,N_25034,N_29564);
nor UO_1232 (O_1232,N_27686,N_27393);
nor UO_1233 (O_1233,N_28825,N_25441);
or UO_1234 (O_1234,N_29559,N_25348);
nand UO_1235 (O_1235,N_28962,N_25574);
nand UO_1236 (O_1236,N_28643,N_28692);
and UO_1237 (O_1237,N_27745,N_25788);
or UO_1238 (O_1238,N_28729,N_26175);
nand UO_1239 (O_1239,N_29472,N_29519);
or UO_1240 (O_1240,N_25545,N_28519);
xnor UO_1241 (O_1241,N_27409,N_25258);
nand UO_1242 (O_1242,N_25521,N_25751);
or UO_1243 (O_1243,N_27545,N_26252);
nor UO_1244 (O_1244,N_25748,N_29107);
nand UO_1245 (O_1245,N_28267,N_25734);
nand UO_1246 (O_1246,N_25325,N_26658);
xor UO_1247 (O_1247,N_26793,N_27064);
nor UO_1248 (O_1248,N_27142,N_26516);
nor UO_1249 (O_1249,N_28959,N_26772);
or UO_1250 (O_1250,N_25020,N_26167);
nor UO_1251 (O_1251,N_25256,N_28366);
nand UO_1252 (O_1252,N_25749,N_29460);
and UO_1253 (O_1253,N_29552,N_26462);
and UO_1254 (O_1254,N_25817,N_28287);
nand UO_1255 (O_1255,N_25209,N_28049);
and UO_1256 (O_1256,N_29914,N_25433);
and UO_1257 (O_1257,N_25950,N_29667);
or UO_1258 (O_1258,N_28812,N_27556);
nor UO_1259 (O_1259,N_25505,N_28383);
and UO_1260 (O_1260,N_25690,N_26007);
xor UO_1261 (O_1261,N_28445,N_28266);
xor UO_1262 (O_1262,N_26697,N_29278);
or UO_1263 (O_1263,N_25520,N_27900);
xnor UO_1264 (O_1264,N_26997,N_28716);
nand UO_1265 (O_1265,N_27926,N_25043);
nor UO_1266 (O_1266,N_28834,N_25889);
nor UO_1267 (O_1267,N_26497,N_28540);
and UO_1268 (O_1268,N_26918,N_26077);
nand UO_1269 (O_1269,N_27248,N_26928);
and UO_1270 (O_1270,N_27797,N_25803);
and UO_1271 (O_1271,N_25244,N_26965);
or UO_1272 (O_1272,N_26479,N_26907);
nor UO_1273 (O_1273,N_29709,N_27613);
xor UO_1274 (O_1274,N_28916,N_29475);
nor UO_1275 (O_1275,N_28545,N_25281);
nand UO_1276 (O_1276,N_28167,N_26801);
nor UO_1277 (O_1277,N_27058,N_29557);
or UO_1278 (O_1278,N_25035,N_26936);
nand UO_1279 (O_1279,N_27931,N_25111);
xor UO_1280 (O_1280,N_27129,N_26698);
nor UO_1281 (O_1281,N_25731,N_27728);
xnor UO_1282 (O_1282,N_27236,N_29961);
and UO_1283 (O_1283,N_25836,N_26289);
xnor UO_1284 (O_1284,N_28623,N_27812);
nor UO_1285 (O_1285,N_29931,N_28795);
nor UO_1286 (O_1286,N_29893,N_26223);
or UO_1287 (O_1287,N_25386,N_26996);
or UO_1288 (O_1288,N_29468,N_28819);
nor UO_1289 (O_1289,N_29594,N_27257);
nand UO_1290 (O_1290,N_28000,N_26384);
or UO_1291 (O_1291,N_26646,N_25918);
nand UO_1292 (O_1292,N_29676,N_26912);
xnor UO_1293 (O_1293,N_27800,N_26636);
or UO_1294 (O_1294,N_25742,N_25511);
and UO_1295 (O_1295,N_29245,N_29121);
and UO_1296 (O_1296,N_29019,N_28365);
nor UO_1297 (O_1297,N_29596,N_27529);
xor UO_1298 (O_1298,N_27953,N_26259);
and UO_1299 (O_1299,N_25664,N_27578);
and UO_1300 (O_1300,N_29201,N_29907);
nor UO_1301 (O_1301,N_27654,N_29404);
or UO_1302 (O_1302,N_26030,N_28628);
and UO_1303 (O_1303,N_26757,N_27392);
nand UO_1304 (O_1304,N_29436,N_25984);
xnor UO_1305 (O_1305,N_29314,N_28206);
nor UO_1306 (O_1306,N_27263,N_29910);
nor UO_1307 (O_1307,N_27137,N_26376);
or UO_1308 (O_1308,N_26109,N_28953);
nor UO_1309 (O_1309,N_25092,N_28874);
and UO_1310 (O_1310,N_27355,N_28508);
xnor UO_1311 (O_1311,N_27090,N_26574);
or UO_1312 (O_1312,N_28891,N_29671);
xnor UO_1313 (O_1313,N_25068,N_25645);
nor UO_1314 (O_1314,N_29860,N_28219);
nand UO_1315 (O_1315,N_27577,N_25101);
nor UO_1316 (O_1316,N_29181,N_25251);
nor UO_1317 (O_1317,N_26870,N_25357);
nor UO_1318 (O_1318,N_26513,N_26437);
and UO_1319 (O_1319,N_25629,N_25987);
nand UO_1320 (O_1320,N_26365,N_25023);
and UO_1321 (O_1321,N_26193,N_25677);
and UO_1322 (O_1322,N_25662,N_27402);
nor UO_1323 (O_1323,N_29607,N_27589);
and UO_1324 (O_1324,N_29505,N_29162);
xor UO_1325 (O_1325,N_28481,N_27709);
xnor UO_1326 (O_1326,N_28730,N_26092);
xor UO_1327 (O_1327,N_25328,N_29858);
xor UO_1328 (O_1328,N_26507,N_25523);
and UO_1329 (O_1329,N_25578,N_26018);
xor UO_1330 (O_1330,N_25372,N_25259);
xor UO_1331 (O_1331,N_26940,N_29269);
nor UO_1332 (O_1332,N_28048,N_27854);
or UO_1333 (O_1333,N_28420,N_26295);
xnor UO_1334 (O_1334,N_25143,N_27028);
nor UO_1335 (O_1335,N_28972,N_25168);
nor UO_1336 (O_1336,N_26867,N_26464);
or UO_1337 (O_1337,N_29291,N_27475);
and UO_1338 (O_1338,N_26296,N_26773);
nand UO_1339 (O_1339,N_27025,N_28034);
nand UO_1340 (O_1340,N_27184,N_25105);
nor UO_1341 (O_1341,N_26784,N_28141);
and UO_1342 (O_1342,N_27676,N_29260);
xnor UO_1343 (O_1343,N_29384,N_29995);
nor UO_1344 (O_1344,N_26056,N_29366);
nor UO_1345 (O_1345,N_26492,N_26086);
or UO_1346 (O_1346,N_26386,N_28922);
or UO_1347 (O_1347,N_26953,N_29187);
or UO_1348 (O_1348,N_25010,N_28872);
nand UO_1349 (O_1349,N_26177,N_27413);
nor UO_1350 (O_1350,N_27865,N_28529);
and UO_1351 (O_1351,N_25582,N_26363);
and UO_1352 (O_1352,N_29239,N_28656);
or UO_1353 (O_1353,N_29979,N_29743);
xor UO_1354 (O_1354,N_29483,N_25022);
nor UO_1355 (O_1355,N_25233,N_25911);
nand UO_1356 (O_1356,N_26207,N_25252);
nor UO_1357 (O_1357,N_29654,N_27489);
nand UO_1358 (O_1358,N_29486,N_28064);
or UO_1359 (O_1359,N_25188,N_26478);
xor UO_1360 (O_1360,N_25703,N_28976);
nor UO_1361 (O_1361,N_27162,N_25714);
and UO_1362 (O_1362,N_25548,N_28615);
or UO_1363 (O_1363,N_28547,N_25216);
nand UO_1364 (O_1364,N_29295,N_25587);
xnor UO_1365 (O_1365,N_29282,N_25560);
nor UO_1366 (O_1366,N_27286,N_26584);
and UO_1367 (O_1367,N_26090,N_26445);
and UO_1368 (O_1368,N_26251,N_27621);
nand UO_1369 (O_1369,N_27951,N_29188);
nor UO_1370 (O_1370,N_29125,N_27666);
or UO_1371 (O_1371,N_26984,N_26662);
nor UO_1372 (O_1372,N_28896,N_27471);
or UO_1373 (O_1373,N_25120,N_26643);
and UO_1374 (O_1374,N_29804,N_26780);
nand UO_1375 (O_1375,N_27167,N_28115);
xnor UO_1376 (O_1376,N_26008,N_27893);
xnor UO_1377 (O_1377,N_29567,N_28666);
nand UO_1378 (O_1378,N_25737,N_29546);
and UO_1379 (O_1379,N_29411,N_29329);
nor UO_1380 (O_1380,N_25584,N_25399);
nor UO_1381 (O_1381,N_28629,N_26209);
nor UO_1382 (O_1382,N_27656,N_29532);
xnor UO_1383 (O_1383,N_25937,N_29525);
or UO_1384 (O_1384,N_26702,N_26841);
nor UO_1385 (O_1385,N_27176,N_27736);
or UO_1386 (O_1386,N_27499,N_29731);
or UO_1387 (O_1387,N_26732,N_25972);
nand UO_1388 (O_1388,N_27600,N_29586);
or UO_1389 (O_1389,N_25390,N_29388);
xor UO_1390 (O_1390,N_25156,N_25089);
or UO_1391 (O_1391,N_25853,N_26487);
or UO_1392 (O_1392,N_25077,N_25320);
nor UO_1393 (O_1393,N_26826,N_28006);
and UO_1394 (O_1394,N_28491,N_27024);
nand UO_1395 (O_1395,N_25858,N_26714);
xor UO_1396 (O_1396,N_28849,N_28703);
and UO_1397 (O_1397,N_28454,N_25241);
xor UO_1398 (O_1398,N_25484,N_25362);
xnor UO_1399 (O_1399,N_25877,N_25669);
nand UO_1400 (O_1400,N_25310,N_26005);
xor UO_1401 (O_1401,N_27511,N_28488);
nand UO_1402 (O_1402,N_26670,N_26083);
nor UO_1403 (O_1403,N_27149,N_26761);
or UO_1404 (O_1404,N_25422,N_26336);
nor UO_1405 (O_1405,N_28274,N_25301);
nand UO_1406 (O_1406,N_26168,N_25346);
xnor UO_1407 (O_1407,N_28221,N_29353);
xnor UO_1408 (O_1408,N_26161,N_27593);
xor UO_1409 (O_1409,N_29630,N_29682);
nand UO_1410 (O_1410,N_25340,N_28768);
or UO_1411 (O_1411,N_27456,N_28061);
or UO_1412 (O_1412,N_27325,N_29376);
and UO_1413 (O_1413,N_25550,N_27500);
nor UO_1414 (O_1414,N_27376,N_25295);
and UO_1415 (O_1415,N_26243,N_27682);
or UO_1416 (O_1416,N_25719,N_29126);
and UO_1417 (O_1417,N_26148,N_29536);
nor UO_1418 (O_1418,N_27806,N_29587);
nand UO_1419 (O_1419,N_28824,N_25902);
or UO_1420 (O_1420,N_26080,N_27823);
nor UO_1421 (O_1421,N_27628,N_26123);
nor UO_1422 (O_1422,N_25332,N_26137);
xnor UO_1423 (O_1423,N_27279,N_28305);
nor UO_1424 (O_1424,N_27208,N_29432);
nor UO_1425 (O_1425,N_27984,N_25401);
xnor UO_1426 (O_1426,N_27042,N_28796);
nand UO_1427 (O_1427,N_25812,N_26617);
and UO_1428 (O_1428,N_29696,N_28611);
and UO_1429 (O_1429,N_29117,N_25891);
and UO_1430 (O_1430,N_25446,N_28806);
or UO_1431 (O_1431,N_27714,N_27544);
or UO_1432 (O_1432,N_26557,N_28930);
nor UO_1433 (O_1433,N_27748,N_27378);
nor UO_1434 (O_1434,N_26121,N_26964);
or UO_1435 (O_1435,N_26426,N_26598);
nor UO_1436 (O_1436,N_28938,N_27947);
or UO_1437 (O_1437,N_29677,N_25577);
xor UO_1438 (O_1438,N_28734,N_26619);
or UO_1439 (O_1439,N_25958,N_27975);
nand UO_1440 (O_1440,N_25364,N_25122);
or UO_1441 (O_1441,N_27181,N_26733);
or UO_1442 (O_1442,N_28493,N_25086);
and UO_1443 (O_1443,N_25276,N_28699);
xnor UO_1444 (O_1444,N_26706,N_29705);
or UO_1445 (O_1445,N_28225,N_28155);
nand UO_1446 (O_1446,N_28553,N_26460);
or UO_1447 (O_1447,N_26518,N_25894);
and UO_1448 (O_1448,N_28736,N_25171);
nand UO_1449 (O_1449,N_27633,N_28791);
or UO_1450 (O_1450,N_26489,N_27923);
and UO_1451 (O_1451,N_27020,N_26937);
nand UO_1452 (O_1452,N_29646,N_26465);
and UO_1453 (O_1453,N_28388,N_25061);
nand UO_1454 (O_1454,N_28144,N_25739);
nand UO_1455 (O_1455,N_28337,N_25255);
or UO_1456 (O_1456,N_28414,N_26848);
nor UO_1457 (O_1457,N_26766,N_26808);
nor UO_1458 (O_1458,N_25689,N_25407);
xor UO_1459 (O_1459,N_27510,N_25132);
nor UO_1460 (O_1460,N_27827,N_26970);
nand UO_1461 (O_1461,N_25977,N_29229);
xor UO_1462 (O_1462,N_25403,N_28109);
or UO_1463 (O_1463,N_28395,N_25556);
nand UO_1464 (O_1464,N_29365,N_26679);
nor UO_1465 (O_1465,N_27791,N_26156);
and UO_1466 (O_1466,N_26589,N_25036);
or UO_1467 (O_1467,N_29565,N_29521);
nor UO_1468 (O_1468,N_29946,N_29160);
nor UO_1469 (O_1469,N_25675,N_27814);
nand UO_1470 (O_1470,N_29871,N_27844);
xnor UO_1471 (O_1471,N_29560,N_28831);
nor UO_1472 (O_1472,N_27133,N_26430);
and UO_1473 (O_1473,N_27704,N_26002);
and UO_1474 (O_1474,N_28177,N_27113);
nor UO_1475 (O_1475,N_27630,N_29419);
or UO_1476 (O_1476,N_27768,N_25722);
or UO_1477 (O_1477,N_26064,N_25821);
nand UO_1478 (O_1478,N_27820,N_26160);
or UO_1479 (O_1479,N_25648,N_26088);
and UO_1480 (O_1480,N_27523,N_26342);
nor UO_1481 (O_1481,N_28523,N_26969);
and UO_1482 (O_1482,N_26486,N_28949);
and UO_1483 (O_1483,N_27368,N_25729);
and UO_1484 (O_1484,N_28502,N_28165);
nand UO_1485 (O_1485,N_26576,N_28007);
xor UO_1486 (O_1486,N_29868,N_25569);
or UO_1487 (O_1487,N_29131,N_27215);
nand UO_1488 (O_1488,N_29911,N_29345);
nor UO_1489 (O_1489,N_26717,N_28738);
xnor UO_1490 (O_1490,N_28732,N_28031);
or UO_1491 (O_1491,N_25352,N_25923);
nand UO_1492 (O_1492,N_26960,N_26381);
and UO_1493 (O_1493,N_26635,N_25411);
xnor UO_1494 (O_1494,N_29938,N_29574);
and UO_1495 (O_1495,N_27107,N_25071);
and UO_1496 (O_1496,N_27983,N_27737);
nor UO_1497 (O_1497,N_25964,N_29771);
xor UO_1498 (O_1498,N_26106,N_25705);
and UO_1499 (O_1499,N_29321,N_28018);
nand UO_1500 (O_1500,N_28747,N_26842);
nand UO_1501 (O_1501,N_26499,N_28855);
nand UO_1502 (O_1502,N_29652,N_27496);
xor UO_1503 (O_1503,N_28045,N_29226);
and UO_1504 (O_1504,N_25928,N_26204);
nand UO_1505 (O_1505,N_29100,N_29155);
nor UO_1506 (O_1506,N_27273,N_28892);
nand UO_1507 (O_1507,N_29374,N_26790);
or UO_1508 (O_1508,N_25490,N_26606);
or UO_1509 (O_1509,N_26860,N_25555);
nor UO_1510 (O_1510,N_25476,N_28917);
and UO_1511 (O_1511,N_27734,N_28354);
xor UO_1512 (O_1512,N_27701,N_28340);
xnor UO_1513 (O_1513,N_26525,N_27957);
nor UO_1514 (O_1514,N_28989,N_28681);
or UO_1515 (O_1515,N_25814,N_28783);
or UO_1516 (O_1516,N_28722,N_29963);
nor UO_1517 (O_1517,N_25225,N_28210);
and UO_1518 (O_1518,N_29937,N_29179);
or UO_1519 (O_1519,N_26882,N_27843);
or UO_1520 (O_1520,N_29900,N_25260);
xnor UO_1521 (O_1521,N_25203,N_29340);
xnor UO_1522 (O_1522,N_27912,N_27147);
nor UO_1523 (O_1523,N_25304,N_27833);
nor UO_1524 (O_1524,N_27742,N_27892);
xor UO_1525 (O_1525,N_27869,N_28127);
nor UO_1526 (O_1526,N_27624,N_28520);
nand UO_1527 (O_1527,N_29869,N_25735);
and UO_1528 (O_1528,N_29144,N_29238);
and UO_1529 (O_1529,N_27543,N_27188);
or UO_1530 (O_1530,N_28312,N_28459);
or UO_1531 (O_1531,N_26476,N_26982);
and UO_1532 (O_1532,N_28742,N_25870);
and UO_1533 (O_1533,N_25833,N_26602);
nand UO_1534 (O_1534,N_27219,N_26815);
and UO_1535 (O_1535,N_25282,N_25708);
nor UO_1536 (O_1536,N_28020,N_27608);
nand UO_1537 (O_1537,N_27217,N_27905);
xor UO_1538 (O_1538,N_28401,N_29135);
nor UO_1539 (O_1539,N_27474,N_27574);
nand UO_1540 (O_1540,N_28082,N_28137);
xnor UO_1541 (O_1541,N_25024,N_29903);
and UO_1542 (O_1542,N_25552,N_26771);
nand UO_1543 (O_1543,N_27033,N_28178);
or UO_1544 (O_1544,N_26181,N_25668);
xnor UO_1545 (O_1545,N_28774,N_28880);
nand UO_1546 (O_1546,N_28494,N_28470);
and UO_1547 (O_1547,N_29044,N_28273);
and UO_1548 (O_1548,N_27932,N_26648);
nand UO_1549 (O_1549,N_29830,N_29908);
nand UO_1550 (O_1550,N_28581,N_27000);
nor UO_1551 (O_1551,N_27935,N_26182);
or UO_1552 (O_1552,N_28073,N_26751);
nor UO_1553 (O_1553,N_29294,N_28597);
and UO_1554 (O_1554,N_29717,N_27525);
xnor UO_1555 (O_1555,N_28556,N_25197);
or UO_1556 (O_1556,N_28214,N_29534);
or UO_1557 (O_1557,N_27220,N_29363);
nor UO_1558 (O_1558,N_27563,N_28723);
nor UO_1559 (O_1559,N_26713,N_27811);
nand UO_1560 (O_1560,N_29346,N_25119);
nor UO_1561 (O_1561,N_27287,N_28402);
nor UO_1562 (O_1562,N_27472,N_26779);
xor UO_1563 (O_1563,N_27048,N_25315);
nand UO_1564 (O_1564,N_27700,N_28466);
nand UO_1565 (O_1565,N_27848,N_28304);
nor UO_1566 (O_1566,N_25242,N_28058);
or UO_1567 (O_1567,N_27468,N_25321);
xnor UO_1568 (O_1568,N_25117,N_25408);
or UO_1569 (O_1569,N_29544,N_27190);
or UO_1570 (O_1570,N_26850,N_26180);
nor UO_1571 (O_1571,N_25639,N_27050);
or UO_1572 (O_1572,N_28386,N_26753);
nor UO_1573 (O_1573,N_25910,N_28351);
nand UO_1574 (O_1574,N_26530,N_26309);
xor UO_1575 (O_1575,N_26600,N_29581);
or UO_1576 (O_1576,N_29969,N_28320);
nand UO_1577 (O_1577,N_26456,N_26029);
nand UO_1578 (O_1578,N_28376,N_28476);
and UO_1579 (O_1579,N_28875,N_25666);
nand UO_1580 (O_1580,N_27198,N_28489);
and UO_1581 (O_1581,N_29801,N_28624);
nand UO_1582 (O_1582,N_25985,N_27114);
nand UO_1583 (O_1583,N_27059,N_27073);
xnor UO_1584 (O_1584,N_25764,N_28677);
xnor UO_1585 (O_1585,N_29369,N_29978);
nor UO_1586 (O_1586,N_28159,N_25381);
nor UO_1587 (O_1587,N_28345,N_27504);
nand UO_1588 (O_1588,N_28744,N_29681);
nor UO_1589 (O_1589,N_27443,N_25246);
nor UO_1590 (O_1590,N_26747,N_28242);
nand UO_1591 (O_1591,N_29224,N_29673);
or UO_1592 (O_1592,N_28564,N_25334);
or UO_1593 (O_1593,N_28649,N_25069);
nor UO_1594 (O_1594,N_27697,N_29499);
nand UO_1595 (O_1595,N_27996,N_26104);
xnor UO_1596 (O_1596,N_28162,N_26210);
xnor UO_1597 (O_1597,N_28835,N_29355);
or UO_1598 (O_1598,N_26661,N_25495);
xnor UO_1599 (O_1599,N_29211,N_28004);
nand UO_1600 (O_1600,N_28585,N_29945);
nand UO_1601 (O_1601,N_26531,N_29834);
and UO_1602 (O_1602,N_27505,N_25824);
xnor UO_1603 (O_1603,N_25524,N_28331);
or UO_1604 (O_1604,N_26326,N_28580);
and UO_1605 (O_1605,N_29095,N_26971);
and UO_1606 (O_1606,N_26335,N_28612);
xnor UO_1607 (O_1607,N_29736,N_27358);
nand UO_1608 (O_1608,N_26830,N_28053);
or UO_1609 (O_1609,N_28074,N_29205);
and UO_1610 (O_1610,N_28076,N_25202);
nand UO_1611 (O_1611,N_27037,N_29020);
nor UO_1612 (O_1612,N_29234,N_25881);
xor UO_1613 (O_1613,N_29659,N_25239);
nor UO_1614 (O_1614,N_27876,N_28958);
or UO_1615 (O_1615,N_28046,N_27672);
or UO_1616 (O_1616,N_26549,N_27230);
or UO_1617 (O_1617,N_25861,N_26622);
or UO_1618 (O_1618,N_26501,N_29650);
and UO_1619 (O_1619,N_28355,N_26608);
nand UO_1620 (O_1620,N_27881,N_25160);
and UO_1621 (O_1621,N_26862,N_25053);
xor UO_1622 (O_1622,N_26979,N_25351);
and UO_1623 (O_1623,N_25416,N_28247);
nand UO_1624 (O_1624,N_25389,N_29615);
nor UO_1625 (O_1625,N_29463,N_25652);
nor UO_1626 (O_1626,N_27079,N_27670);
and UO_1627 (O_1627,N_29930,N_27816);
and UO_1628 (O_1628,N_28586,N_29413);
nand UO_1629 (O_1629,N_28341,N_27088);
xnor UO_1630 (O_1630,N_27512,N_29168);
nor UO_1631 (O_1631,N_25971,N_25867);
nor UO_1632 (O_1632,N_26760,N_26314);
or UO_1633 (O_1633,N_28246,N_28308);
or UO_1634 (O_1634,N_28594,N_27487);
and UO_1635 (O_1635,N_29141,N_26981);
xnor UO_1636 (O_1636,N_29994,N_28940);
xnor UO_1637 (O_1637,N_26316,N_28924);
and UO_1638 (O_1638,N_27917,N_27280);
and UO_1639 (O_1639,N_26461,N_27649);
nand UO_1640 (O_1640,N_29790,N_28419);
or UO_1641 (O_1641,N_29407,N_28211);
xor UO_1642 (O_1642,N_25815,N_26998);
xor UO_1643 (O_1643,N_25954,N_27554);
nor UO_1644 (O_1644,N_27094,N_29381);
or UO_1645 (O_1645,N_29332,N_27677);
xnor UO_1646 (O_1646,N_28301,N_26103);
or UO_1647 (O_1647,N_25226,N_25992);
xnor UO_1648 (O_1648,N_28378,N_27041);
xnor UO_1649 (O_1649,N_28588,N_27524);
nand UO_1650 (O_1650,N_29464,N_25080);
nor UO_1651 (O_1651,N_26939,N_28421);
and UO_1652 (O_1652,N_27008,N_25700);
xor UO_1653 (O_1653,N_27374,N_26039);
nor UO_1654 (O_1654,N_27428,N_29807);
or UO_1655 (O_1655,N_27056,N_26611);
or UO_1656 (O_1656,N_29497,N_25940);
or UO_1657 (O_1657,N_27072,N_26567);
nand UO_1658 (O_1658,N_25379,N_26140);
nand UO_1659 (O_1659,N_26020,N_26034);
or UO_1660 (O_1660,N_28235,N_26596);
or UO_1661 (O_1661,N_25628,N_29038);
and UO_1662 (O_1662,N_26343,N_26886);
nand UO_1663 (O_1663,N_27119,N_28261);
nand UO_1664 (O_1664,N_26198,N_26693);
or UO_1665 (O_1665,N_26199,N_25816);
xor UO_1666 (O_1666,N_27096,N_27151);
nor UO_1667 (O_1667,N_27756,N_28726);
and UO_1668 (O_1668,N_25635,N_28268);
nand UO_1669 (O_1669,N_27870,N_26560);
nand UO_1670 (O_1670,N_27693,N_26144);
xnor UO_1671 (O_1671,N_26075,N_26025);
and UO_1672 (O_1672,N_25201,N_25133);
or UO_1673 (O_1673,N_26768,N_26015);
and UO_1674 (O_1674,N_25595,N_29859);
nor UO_1675 (O_1675,N_29522,N_27469);
nand UO_1676 (O_1676,N_27457,N_29082);
nor UO_1677 (O_1677,N_28208,N_27939);
xor UO_1678 (O_1678,N_29626,N_27003);
and UO_1679 (O_1679,N_27533,N_25002);
and UO_1680 (O_1680,N_27116,N_29354);
nand UO_1681 (O_1681,N_28205,N_27602);
and UO_1682 (O_1682,N_25897,N_29690);
xnor UO_1683 (O_1683,N_28390,N_29387);
xnor UO_1684 (O_1684,N_28079,N_26033);
xor UO_1685 (O_1685,N_27108,N_26413);
nand UO_1686 (O_1686,N_29055,N_29231);
nor UO_1687 (O_1687,N_25660,N_26615);
nand UO_1688 (O_1688,N_27568,N_26961);
nor UO_1689 (O_1689,N_29225,N_25155);
and UO_1690 (O_1690,N_27044,N_29257);
xor UO_1691 (O_1691,N_27313,N_29686);
or UO_1692 (O_1692,N_27483,N_29898);
nor UO_1693 (O_1693,N_28971,N_27418);
xnor UO_1694 (O_1694,N_28014,N_28551);
and UO_1695 (O_1695,N_25613,N_25924);
xnor UO_1696 (O_1696,N_27581,N_28428);
or UO_1697 (O_1697,N_25761,N_28293);
nand UO_1698 (O_1698,N_25015,N_27721);
xnor UO_1699 (O_1699,N_28085,N_26248);
or UO_1700 (O_1700,N_28937,N_26063);
or UO_1701 (O_1701,N_27516,N_26087);
or UO_1702 (O_1702,N_27452,N_25537);
or UO_1703 (O_1703,N_26201,N_26599);
and UO_1704 (O_1704,N_29023,N_25682);
nand UO_1705 (O_1705,N_28497,N_28116);
xor UO_1706 (O_1706,N_26253,N_26097);
nor UO_1707 (O_1707,N_27754,N_29591);
xor UO_1708 (O_1708,N_26986,N_28368);
nor UO_1709 (O_1709,N_26441,N_25030);
nand UO_1710 (O_1710,N_28280,N_29732);
xnor UO_1711 (O_1711,N_27412,N_29601);
or UO_1712 (O_1712,N_28720,N_27720);
nand UO_1713 (O_1713,N_25617,N_28613);
nor UO_1714 (O_1714,N_25978,N_28633);
or UO_1715 (O_1715,N_27103,N_25694);
nand UO_1716 (O_1716,N_28436,N_25898);
nand UO_1717 (O_1717,N_29992,N_29998);
or UO_1718 (O_1718,N_27246,N_27997);
and UO_1719 (O_1719,N_26490,N_29767);
nor UO_1720 (O_1720,N_27154,N_27066);
nor UO_1721 (O_1721,N_26710,N_28518);
nand UO_1722 (O_1722,N_29981,N_25908);
or UO_1723 (O_1723,N_27084,N_29057);
nor UO_1724 (O_1724,N_26520,N_26800);
and UO_1725 (O_1725,N_29017,N_25864);
and UO_1726 (O_1726,N_29470,N_28843);
nand UO_1727 (O_1727,N_29076,N_27650);
and UO_1728 (O_1728,N_29504,N_29360);
or UO_1729 (O_1729,N_26229,N_29129);
xnor UO_1730 (O_1730,N_28883,N_26374);
nand UO_1731 (O_1731,N_26814,N_25313);
or UO_1732 (O_1732,N_25755,N_27197);
nand UO_1733 (O_1733,N_26711,N_27371);
nor UO_1734 (O_1734,N_25503,N_29971);
nand UO_1735 (O_1735,N_29889,N_28966);
xor UO_1736 (O_1736,N_28546,N_25509);
or UO_1737 (O_1737,N_29185,N_29005);
nand UO_1738 (O_1738,N_28450,N_25723);
or UO_1739 (O_1739,N_25392,N_29571);
nand UO_1740 (O_1740,N_26043,N_27318);
nor UO_1741 (O_1741,N_27713,N_25945);
nor UO_1742 (O_1742,N_28503,N_29610);
or UO_1743 (O_1743,N_29204,N_28289);
or UO_1744 (O_1744,N_29481,N_29692);
nand UO_1745 (O_1745,N_28893,N_27729);
xor UO_1746 (O_1746,N_29588,N_28859);
xnor UO_1747 (O_1747,N_26401,N_28674);
nand UO_1748 (O_1748,N_27408,N_26102);
nand UO_1749 (O_1749,N_28307,N_26291);
xnor UO_1750 (O_1750,N_27740,N_29406);
nor UO_1751 (O_1751,N_29929,N_29573);
xnor UO_1752 (O_1752,N_28490,N_29274);
nor UO_1753 (O_1753,N_26054,N_25901);
or UO_1754 (O_1754,N_28217,N_26402);
nor UO_1755 (O_1755,N_27776,N_28456);
xor UO_1756 (O_1756,N_28985,N_27916);
xnor UO_1757 (O_1757,N_29698,N_27010);
nand UO_1758 (O_1758,N_27834,N_28234);
or UO_1759 (O_1759,N_25713,N_26903);
and UO_1760 (O_1760,N_28948,N_29115);
nor UO_1761 (O_1761,N_27871,N_28513);
xor UO_1762 (O_1762,N_27043,N_25775);
or UO_1763 (O_1763,N_29895,N_28610);
and UO_1764 (O_1764,N_25789,N_28975);
nand UO_1765 (O_1765,N_27810,N_27467);
or UO_1766 (O_1766,N_28151,N_29648);
nor UO_1767 (O_1767,N_28929,N_27470);
or UO_1768 (O_1768,N_28592,N_26993);
or UO_1769 (O_1769,N_27051,N_25106);
nor UO_1770 (O_1770,N_25832,N_26948);
nor UO_1771 (O_1771,N_29030,N_27138);
nand UO_1772 (O_1772,N_28717,N_29280);
nand UO_1773 (O_1773,N_28635,N_27789);
or UO_1774 (O_1774,N_29902,N_26392);
nand UO_1775 (O_1775,N_28028,N_29585);
xor UO_1776 (O_1776,N_26578,N_26680);
nand UO_1777 (O_1777,N_25493,N_29789);
xor UO_1778 (O_1778,N_29101,N_28296);
nand UO_1779 (O_1779,N_26046,N_28781);
xnor UO_1780 (O_1780,N_28956,N_27125);
xnor UO_1781 (O_1781,N_26453,N_27480);
xnor UO_1782 (O_1782,N_28693,N_26436);
xnor UO_1783 (O_1783,N_25607,N_26595);
nand UO_1784 (O_1784,N_28360,N_27783);
or UO_1785 (O_1785,N_28324,N_28601);
nand UO_1786 (O_1786,N_28577,N_27441);
nand UO_1787 (O_1787,N_28317,N_27321);
and UO_1788 (O_1788,N_25146,N_26837);
xnor UO_1789 (O_1789,N_29391,N_29222);
or UO_1790 (O_1790,N_26089,N_27668);
and UO_1791 (O_1791,N_29090,N_27250);
and UO_1792 (O_1792,N_29975,N_29845);
nor UO_1793 (O_1793,N_25139,N_29219);
or UO_1794 (O_1794,N_27605,N_26555);
and UO_1795 (O_1795,N_25604,N_27890);
or UO_1796 (O_1796,N_28468,N_25450);
or UO_1797 (O_1797,N_27815,N_26985);
and UO_1798 (O_1798,N_28129,N_28531);
nand UO_1799 (O_1799,N_25921,N_29259);
or UO_1800 (O_1800,N_28067,N_27767);
xnor UO_1801 (O_1801,N_26238,N_29749);
or UO_1802 (O_1802,N_26906,N_27807);
xor UO_1803 (O_1803,N_28512,N_29304);
xor UO_1804 (O_1804,N_27817,N_25424);
and UO_1805 (O_1805,N_27763,N_26225);
or UO_1806 (O_1806,N_26122,N_28558);
nor UO_1807 (O_1807,N_29164,N_28393);
xor UO_1808 (O_1808,N_26895,N_28353);
and UO_1809 (O_1809,N_29927,N_28914);
xnor UO_1810 (O_1810,N_26935,N_25059);
or UO_1811 (O_1811,N_26739,N_28147);
xor UO_1812 (O_1812,N_26132,N_27204);
or UO_1813 (O_1813,N_26010,N_28823);
and UO_1814 (O_1814,N_27819,N_28248);
xnor UO_1815 (O_1815,N_25076,N_26983);
and UO_1816 (O_1816,N_26419,N_28864);
or UO_1817 (O_1817,N_28764,N_27557);
and UO_1818 (O_1818,N_27234,N_29172);
nand UO_1819 (O_1819,N_29540,N_28485);
nor UO_1820 (O_1820,N_29913,N_27427);
and UO_1821 (O_1821,N_26186,N_29855);
nand UO_1822 (O_1822,N_26504,N_26178);
xnor UO_1823 (O_1823,N_26094,N_25483);
or UO_1824 (O_1824,N_26468,N_26267);
and UO_1825 (O_1825,N_26920,N_29774);
and UO_1826 (O_1826,N_27345,N_29857);
nand UO_1827 (O_1827,N_27884,N_25205);
nand UO_1828 (O_1828,N_26052,N_28582);
nand UO_1829 (O_1829,N_27077,N_27588);
and UO_1830 (O_1830,N_27401,N_26540);
nand UO_1831 (O_1831,N_25488,N_27311);
or UO_1832 (O_1832,N_25554,N_26000);
and UO_1833 (O_1833,N_25857,N_25339);
nand UO_1834 (O_1834,N_25829,N_29663);
or UO_1835 (O_1835,N_27919,N_29200);
nor UO_1836 (O_1836,N_28927,N_25126);
and UO_1837 (O_1837,N_29817,N_29330);
xor UO_1838 (O_1838,N_27106,N_28604);
or UO_1839 (O_1839,N_25782,N_29041);
nand UO_1840 (O_1840,N_28590,N_29508);
nand UO_1841 (O_1841,N_28925,N_27221);
nor UO_1842 (O_1842,N_26829,N_29359);
xnor UO_1843 (O_1843,N_28721,N_27040);
nand UO_1844 (O_1844,N_28852,N_25167);
nand UO_1845 (O_1845,N_26219,N_29899);
xnor UO_1846 (O_1846,N_26272,N_29275);
xnor UO_1847 (O_1847,N_27146,N_25039);
or UO_1848 (O_1848,N_26952,N_26036);
nand UO_1849 (O_1849,N_26791,N_29548);
nand UO_1850 (O_1850,N_29704,N_28669);
nor UO_1851 (O_1851,N_25658,N_29078);
nor UO_1852 (O_1852,N_29088,N_27281);
or UO_1853 (O_1853,N_28119,N_28661);
xor UO_1854 (O_1854,N_25184,N_25095);
nor UO_1855 (O_1855,N_25525,N_25169);
xnor UO_1856 (O_1856,N_25531,N_28005);
xor UO_1857 (O_1857,N_26001,N_29127);
and UO_1858 (O_1858,N_26554,N_28857);
and UO_1859 (O_1859,N_29605,N_28653);
nand UO_1860 (O_1860,N_29270,N_26141);
nand UO_1861 (O_1861,N_28833,N_28072);
and UO_1862 (O_1862,N_27867,N_27322);
xnor UO_1863 (O_1863,N_29759,N_28515);
xnor UO_1864 (O_1864,N_27564,N_27039);
and UO_1865 (O_1865,N_29901,N_26032);
or UO_1866 (O_1866,N_29308,N_29660);
nor UO_1867 (O_1867,N_29093,N_26755);
nor UO_1868 (O_1868,N_25938,N_27643);
xnor UO_1869 (O_1869,N_28191,N_27673);
or UO_1870 (O_1870,N_28200,N_25863);
xnor UO_1871 (O_1871,N_26241,N_25859);
nand UO_1872 (O_1872,N_27882,N_29668);
nor UO_1873 (O_1873,N_29036,N_28733);
and UO_1874 (O_1874,N_29838,N_26084);
and UO_1875 (O_1875,N_28672,N_29768);
and UO_1876 (O_1876,N_25398,N_27315);
nand UO_1877 (O_1877,N_28584,N_26633);
nor UO_1878 (O_1878,N_25037,N_25421);
and UO_1879 (O_1879,N_28432,N_27383);
and UO_1880 (O_1880,N_25153,N_27657);
nand UO_1881 (O_1881,N_27422,N_25640);
xor UO_1882 (O_1882,N_28926,N_27101);
xnor UO_1883 (O_1883,N_27979,N_29616);
nor UO_1884 (O_1884,N_29516,N_26270);
or UO_1885 (O_1885,N_29751,N_25444);
and UO_1886 (O_1886,N_29599,N_26632);
xor UO_1887 (O_1887,N_26226,N_26686);
and UO_1888 (O_1888,N_27194,N_28979);
or UO_1889 (O_1889,N_27845,N_27716);
xor UO_1890 (O_1890,N_26022,N_29489);
nor UO_1891 (O_1891,N_29026,N_26902);
nor UO_1892 (O_1892,N_29680,N_29533);
xnor UO_1893 (O_1893,N_26158,N_26190);
nor UO_1894 (O_1894,N_29043,N_25267);
xnor UO_1895 (O_1895,N_26183,N_29347);
nor UO_1896 (O_1896,N_29191,N_28319);
and UO_1897 (O_1897,N_29378,N_26021);
nor UO_1898 (O_1898,N_26067,N_27440);
nand UO_1899 (O_1899,N_27211,N_27873);
and UO_1900 (O_1900,N_27655,N_27007);
nor UO_1901 (O_1901,N_29876,N_25649);
and UO_1902 (O_1902,N_28621,N_29014);
and UO_1903 (O_1903,N_26512,N_29741);
nand UO_1904 (O_1904,N_29820,N_26233);
or UO_1905 (O_1905,N_25439,N_25656);
xor UO_1906 (O_1906,N_29013,N_27207);
nor UO_1907 (O_1907,N_28050,N_28595);
nor UO_1908 (O_1908,N_25090,N_29592);
xnor UO_1909 (O_1909,N_29349,N_27164);
nor UO_1910 (O_1910,N_25618,N_29575);
or UO_1911 (O_1911,N_27587,N_27253);
nand UO_1912 (O_1912,N_25506,N_27803);
nor UO_1913 (O_1913,N_26150,N_29835);
and UO_1914 (O_1914,N_25831,N_29725);
and UO_1915 (O_1915,N_26013,N_29455);
nor UO_1916 (O_1916,N_26117,N_26135);
or UO_1917 (O_1917,N_28447,N_27049);
and UO_1918 (O_1918,N_29104,N_25973);
nand UO_1919 (O_1919,N_27927,N_28339);
or UO_1920 (O_1920,N_26482,N_27688);
nand UO_1921 (O_1921,N_25638,N_29450);
nand UO_1922 (O_1922,N_25680,N_27584);
or UO_1923 (O_1923,N_29827,N_27880);
xor UO_1924 (O_1924,N_25504,N_26759);
nand UO_1925 (O_1925,N_27731,N_26126);
or UO_1926 (O_1926,N_26744,N_26688);
nor UO_1927 (O_1927,N_26893,N_28370);
nor UO_1928 (O_1928,N_29572,N_25189);
and UO_1929 (O_1929,N_27928,N_28439);
or UO_1930 (O_1930,N_27850,N_29011);
nor UO_1931 (O_1931,N_26250,N_29699);
and UO_1932 (O_1932,N_28186,N_28250);
nand UO_1933 (O_1933,N_29558,N_28620);
nand UO_1934 (O_1934,N_28175,N_26458);
xor UO_1935 (O_1935,N_26951,N_29850);
nand UO_1936 (O_1936,N_29645,N_29500);
nand UO_1937 (O_1937,N_27259,N_29202);
nor UO_1938 (O_1938,N_27771,N_27583);
and UO_1939 (O_1939,N_27794,N_25593);
or UO_1940 (O_1940,N_25409,N_28921);
xor UO_1941 (O_1941,N_27847,N_29159);
or UO_1942 (O_1942,N_29420,N_25210);
nand UO_1943 (O_1943,N_29003,N_28642);
or UO_1944 (O_1944,N_28152,N_27653);
nand UO_1945 (O_1945,N_28977,N_27687);
or UO_1946 (O_1946,N_25589,N_28083);
nand UO_1947 (O_1947,N_28886,N_29570);
or UO_1948 (O_1948,N_25839,N_26521);
nor UO_1949 (O_1949,N_25932,N_25657);
xor UO_1950 (O_1950,N_29389,N_26202);
nand UO_1951 (O_1951,N_25855,N_25886);
or UO_1952 (O_1952,N_25654,N_25616);
xnor UO_1953 (O_1953,N_27595,N_26966);
or UO_1954 (O_1954,N_29367,N_29362);
or UO_1955 (O_1955,N_25961,N_27267);
nor UO_1956 (O_1956,N_26835,N_26053);
and UO_1957 (O_1957,N_29877,N_26317);
or UO_1958 (O_1958,N_29153,N_29727);
nor UO_1959 (O_1959,N_29453,N_26770);
nor UO_1960 (O_1960,N_25265,N_29870);
or UO_1961 (O_1961,N_26775,N_25783);
or UO_1962 (O_1962,N_26361,N_28991);
xor UO_1963 (O_1963,N_26878,N_28560);
and UO_1964 (O_1964,N_29237,N_25341);
nor UO_1965 (O_1965,N_26232,N_27695);
or UO_1966 (O_1966,N_28794,N_26588);
nor UO_1967 (O_1967,N_25585,N_29452);
xor UO_1968 (O_1968,N_26631,N_27086);
or UO_1969 (O_1969,N_26910,N_29740);
nand UO_1970 (O_1970,N_29849,N_28311);
nand UO_1971 (O_1971,N_28322,N_28174);
nor UO_1972 (O_1972,N_26551,N_29186);
nand UO_1973 (O_1973,N_25262,N_28323);
nand UO_1974 (O_1974,N_27838,N_26220);
xor UO_1975 (O_1975,N_27400,N_27929);
nand UO_1976 (O_1976,N_25283,N_26414);
xor UO_1977 (O_1977,N_29647,N_28284);
xor UO_1978 (O_1978,N_25098,N_25151);
and UO_1979 (O_1979,N_25289,N_29149);
xnor UO_1980 (O_1980,N_25300,N_28252);
nor UO_1981 (O_1981,N_29904,N_28121);
and UO_1982 (O_1982,N_26153,N_27562);
nor UO_1983 (O_1983,N_28839,N_28349);
nor UO_1984 (O_1984,N_27761,N_27569);
or UO_1985 (O_1985,N_26625,N_26605);
nand UO_1986 (O_1986,N_28583,N_28172);
nand UO_1987 (O_1987,N_25195,N_28313);
nor UO_1988 (O_1988,N_29785,N_27362);
and UO_1989 (O_1989,N_27933,N_25312);
or UO_1990 (O_1990,N_28596,N_27365);
and UO_1991 (O_1991,N_26581,N_27235);
nor UO_1992 (O_1992,N_29343,N_26262);
and UO_1993 (O_1993,N_28695,N_27842);
nand UO_1994 (O_1994,N_28290,N_26302);
and UO_1995 (O_1995,N_25900,N_25740);
and UO_1996 (O_1996,N_27609,N_26901);
and UO_1997 (O_1997,N_28471,N_28499);
or UO_1998 (O_1998,N_28982,N_28890);
or UO_1999 (O_1999,N_27366,N_26655);
nand UO_2000 (O_2000,N_28093,N_28292);
or UO_2001 (O_2001,N_27265,N_27615);
nand UO_2002 (O_2002,N_26579,N_28239);
nand UO_2003 (O_2003,N_27799,N_27698);
and UO_2004 (O_2004,N_26418,N_25199);
nand UO_2005 (O_2005,N_27205,N_26720);
xnor UO_2006 (O_2006,N_27238,N_27535);
and UO_2007 (O_2007,N_25344,N_27433);
nor UO_2008 (O_2008,N_26255,N_28112);
nand UO_2009 (O_2009,N_25830,N_25040);
nor UO_2010 (O_2010,N_25611,N_27786);
and UO_2011 (O_2011,N_26723,N_29379);
nand UO_2012 (O_2012,N_26508,N_29451);
and UO_2013 (O_2013,N_27897,N_27195);
and UO_2014 (O_2014,N_25732,N_27978);
nand UO_2015 (O_2015,N_28931,N_29707);
or UO_2016 (O_2016,N_28751,N_27618);
or UO_2017 (O_2017,N_27370,N_27179);
or UO_2018 (O_2018,N_27764,N_26917);
or UO_2019 (O_2019,N_25542,N_25798);
xor UO_2020 (O_2020,N_27477,N_27297);
nor UO_2021 (O_2021,N_28407,N_28555);
or UO_2022 (O_2022,N_27175,N_29077);
xnor UO_2023 (O_2023,N_26412,N_27998);
nor UO_2024 (O_2024,N_25254,N_25571);
or UO_2025 (O_2025,N_28691,N_26810);
nor UO_2026 (O_2026,N_25135,N_28042);
xnor UO_2027 (O_2027,N_25596,N_28369);
or UO_2028 (O_2028,N_28690,N_28135);
and UO_2029 (O_2029,N_28111,N_25309);
and UO_2030 (O_2030,N_26667,N_29555);
nor UO_2031 (O_2031,N_29099,N_25769);
or UO_2032 (O_2032,N_29936,N_28054);
nor UO_2033 (O_2033,N_28740,N_29623);
nand UO_2034 (O_2034,N_25222,N_27531);
or UO_2035 (O_2035,N_29173,N_25880);
xnor UO_2036 (O_2036,N_28300,N_29190);
nor UO_2037 (O_2037,N_28110,N_27292);
or UO_2038 (O_2038,N_27417,N_29210);
and UO_2039 (O_2039,N_29644,N_25549);
nand UO_2040 (O_2040,N_25026,N_29008);
or UO_2041 (O_2041,N_27013,N_25733);
xnor UO_2042 (O_2042,N_25543,N_29166);
nand UO_2043 (O_2043,N_28066,N_27326);
or UO_2044 (O_2044,N_29972,N_26896);
xnor UO_2045 (O_2045,N_27766,N_27661);
or UO_2046 (O_2046,N_26816,N_28357);
or UO_2047 (O_2047,N_25976,N_25263);
and UO_2048 (O_2048,N_26341,N_25744);
and UO_2049 (O_2049,N_26909,N_26352);
xor UO_2050 (O_2050,N_25786,N_26626);
nor UO_2051 (O_2051,N_25873,N_28631);
nand UO_2052 (O_2052,N_26665,N_25479);
nand UO_2053 (O_2053,N_29342,N_29444);
xnor UO_2054 (O_2054,N_26892,N_29761);
nor UO_2055 (O_2055,N_28698,N_29866);
nand UO_2056 (O_2056,N_28920,N_29255);
xnor UO_2057 (O_2057,N_28256,N_29728);
and UO_2058 (O_2058,N_27170,N_29040);
or UO_2059 (O_2059,N_27969,N_26328);
and UO_2060 (O_2060,N_27386,N_27906);
nor UO_2061 (O_2061,N_27541,N_29465);
or UO_2062 (O_2062,N_27946,N_28204);
nand UO_2063 (O_2063,N_25619,N_28441);
and UO_2064 (O_2064,N_25154,N_26415);
and UO_2065 (O_2065,N_27974,N_29243);
and UO_2066 (O_2066,N_26404,N_25227);
or UO_2067 (O_2067,N_28969,N_28259);
or UO_2068 (O_2068,N_25125,N_28801);
and UO_2069 (O_2069,N_26889,N_29390);
nor UO_2070 (O_2070,N_26955,N_27314);
and UO_2071 (O_2071,N_25396,N_27491);
nand UO_2072 (O_2072,N_28188,N_27889);
and UO_2073 (O_2073,N_26332,N_29180);
nand UO_2074 (O_2074,N_25730,N_26170);
and UO_2075 (O_2075,N_27123,N_28309);
or UO_2076 (O_2076,N_28394,N_25363);
xnor UO_2077 (O_2077,N_25834,N_25854);
nor UO_2078 (O_2078,N_28224,N_28442);
nor UO_2079 (O_2079,N_26004,N_27753);
nand UO_2080 (O_2080,N_27691,N_25636);
nand UO_2081 (O_2081,N_29396,N_27308);
nor UO_2082 (O_2082,N_28131,N_27538);
xor UO_2083 (O_2083,N_29254,N_29526);
nor UO_2084 (O_2084,N_28068,N_27158);
and UO_2085 (O_2085,N_26712,N_29683);
nand UO_2086 (O_2086,N_25828,N_25727);
nor UO_2087 (O_2087,N_28123,N_28701);
or UO_2088 (O_2088,N_28837,N_29954);
nand UO_2089 (O_2089,N_27210,N_28575);
or UO_2090 (O_2090,N_26470,N_29297);
nor UO_2091 (O_2091,N_25333,N_25718);
xor UO_2092 (O_2092,N_26881,N_25166);
nand UO_2093 (O_2093,N_25736,N_29883);
nand UO_2094 (O_2094,N_28176,N_25297);
xnor UO_2095 (O_2095,N_26382,N_27874);
xnor UO_2096 (O_2096,N_26062,N_28096);
nor UO_2097 (O_2097,N_26099,N_26152);
nand UO_2098 (O_2098,N_27294,N_28075);
and UO_2099 (O_2099,N_27636,N_29694);
nor UO_2100 (O_2100,N_25576,N_27956);
xnor UO_2101 (O_2101,N_29700,N_27249);
nand UO_2102 (O_2102,N_27992,N_27977);
nor UO_2103 (O_2103,N_28166,N_26959);
nor UO_2104 (O_2104,N_26663,N_25841);
nand UO_2105 (O_2105,N_26795,N_29545);
or UO_2106 (O_2106,N_28065,N_27290);
and UO_2107 (O_2107,N_29884,N_29492);
nand UO_2108 (O_2108,N_25021,N_25890);
nor UO_2109 (O_2109,N_26360,N_29258);
or UO_2110 (O_2110,N_29307,N_27852);
and UO_2111 (O_2111,N_27112,N_29639);
xnor UO_2112 (O_2112,N_26945,N_29595);
nand UO_2113 (O_2113,N_28568,N_28566);
xnor UO_2114 (O_2114,N_28253,N_29252);
xor UO_2115 (O_2115,N_25796,N_27430);
and UO_2116 (O_2116,N_28486,N_25772);
nor UO_2117 (O_2117,N_26399,N_29755);
or UO_2118 (O_2118,N_26091,N_29424);
xnor UO_2119 (O_2119,N_26146,N_28809);
xnor UO_2120 (O_2120,N_26125,N_25055);
nor UO_2121 (O_2121,N_25962,N_29025);
xor UO_2122 (O_2122,N_27922,N_26794);
and UO_2123 (O_2123,N_27166,N_25759);
and UO_2124 (O_2124,N_26378,N_26677);
nor UO_2125 (O_2125,N_28003,N_29039);
xnor UO_2126 (O_2126,N_29066,N_27920);
or UO_2127 (O_2127,N_26017,N_29446);
xnor UO_2128 (O_2128,N_27835,N_28228);
xnor UO_2129 (O_2129,N_28640,N_26324);
xor UO_2130 (O_2130,N_28326,N_25235);
and UO_2131 (O_2131,N_28207,N_29697);
or UO_2132 (O_2132,N_29833,N_26999);
and UO_2133 (O_2133,N_29192,N_27769);
or UO_2134 (O_2134,N_29147,N_25679);
xor UO_2135 (O_2135,N_28827,N_26824);
or UO_2136 (O_2136,N_28363,N_26788);
and UO_2137 (O_2137,N_25331,N_28557);
nor UO_2138 (O_2138,N_29814,N_25933);
and UO_2139 (O_2139,N_25261,N_26561);
xor UO_2140 (O_2140,N_29326,N_27712);
nor UO_2141 (O_2141,N_28614,N_25336);
nand UO_2142 (O_2142,N_29031,N_28226);
nand UO_2143 (O_2143,N_29515,N_26288);
nand UO_2144 (O_2144,N_26839,N_29046);
nor UO_2145 (O_2145,N_29949,N_25818);
and UO_2146 (O_2146,N_28010,N_29324);
or UO_2147 (O_2147,N_27934,N_26890);
and UO_2148 (O_2148,N_28117,N_29600);
nor UO_2149 (O_2149,N_28817,N_27904);
and UO_2150 (O_2150,N_26398,N_27726);
nand UO_2151 (O_2151,N_26442,N_26345);
nor UO_2152 (O_2152,N_25883,N_25527);
nor UO_2153 (O_2153,N_26040,N_26510);
and UO_2154 (O_2154,N_27921,N_29917);
and UO_2155 (O_2155,N_26634,N_27140);
nor UO_2156 (O_2156,N_28408,N_25280);
and UO_2157 (O_2157,N_26957,N_25693);
or UO_2158 (O_2158,N_26672,N_25425);
nand UO_2159 (O_2159,N_26765,N_26493);
or UO_2160 (O_2160,N_27384,N_25627);
and UO_2161 (O_2161,N_29306,N_26754);
nor UO_2162 (O_2162,N_25075,N_29247);
xor UO_2163 (O_2163,N_27795,N_29167);
nor UO_2164 (O_2164,N_28708,N_28081);
and UO_2165 (O_2165,N_28678,N_25612);
and UO_2166 (O_2166,N_29622,N_27561);
nor UO_2167 (O_2167,N_28318,N_25052);
or UO_2168 (O_2168,N_26743,N_29430);
and UO_2169 (O_2169,N_25979,N_27122);
nand UO_2170 (O_2170,N_25936,N_27942);
nand UO_2171 (O_2171,N_27486,N_29409);
or UO_2172 (O_2172,N_25534,N_27485);
or UO_2173 (O_2173,N_26438,N_26641);
nor UO_2174 (O_2174,N_28957,N_29196);
and UO_2175 (O_2175,N_27111,N_26235);
or UO_2176 (O_2176,N_26203,N_29312);
xor UO_2177 (O_2177,N_26894,N_27275);
nor UO_2178 (O_2178,N_25850,N_28745);
xor UO_2179 (O_2179,N_25570,N_28525);
nand UO_2180 (O_2180,N_28798,N_28725);
or UO_2181 (O_2181,N_25546,N_28134);
nor UO_2182 (O_2182,N_29227,N_29665);
or UO_2183 (O_2183,N_29339,N_28662);
or UO_2184 (O_2184,N_28844,N_25322);
xnor UO_2185 (O_2185,N_29769,N_26258);
xnor UO_2186 (O_2186,N_26565,N_25338);
nand UO_2187 (O_2187,N_29110,N_27012);
nor UO_2188 (O_2188,N_27057,N_25011);
nand UO_2189 (O_2189,N_28335,N_27382);
and UO_2190 (O_2190,N_25909,N_29195);
or UO_2191 (O_2191,N_25391,N_28130);
xnor UO_2192 (O_2192,N_27646,N_28943);
nand UO_2193 (O_2193,N_26055,N_28950);
nor UO_2194 (O_2194,N_28973,N_28241);
xnor UO_2195 (O_2195,N_27346,N_25871);
nand UO_2196 (O_2196,N_28960,N_26845);
and UO_2197 (O_2197,N_28544,N_29154);
nor UO_2198 (O_2198,N_28944,N_29454);
nand UO_2199 (O_2199,N_29613,N_25637);
nor UO_2200 (O_2200,N_29636,N_25599);
xor UO_2201 (O_2201,N_28746,N_25515);
nand UO_2202 (O_2202,N_29896,N_25706);
xor UO_2203 (O_2203,N_29593,N_29333);
nor UO_2204 (O_2204,N_29495,N_26654);
or UO_2205 (O_2205,N_28563,N_29878);
nor UO_2206 (O_2206,N_26081,N_28763);
xor UO_2207 (O_2207,N_27414,N_25768);
nand UO_2208 (O_2208,N_25248,N_28762);
nor UO_2209 (O_2209,N_27439,N_26411);
nor UO_2210 (O_2210,N_27548,N_25275);
nand UO_2211 (O_2211,N_29941,N_26573);
nor UO_2212 (O_2212,N_25349,N_28799);
or UO_2213 (O_2213,N_28179,N_25307);
nor UO_2214 (O_2214,N_26416,N_25808);
nand UO_2215 (O_2215,N_29674,N_27399);
nor UO_2216 (O_2216,N_25470,N_27760);
or UO_2217 (O_2217,N_27949,N_25800);
nand UO_2218 (O_2218,N_28876,N_27369);
or UO_2219 (O_2219,N_28359,N_27435);
nand UO_2220 (O_2220,N_25603,N_25709);
xnor UO_2221 (O_2221,N_25651,N_26408);
xor UO_2222 (O_2222,N_29541,N_28670);
nor UO_2223 (O_2223,N_25190,N_28126);
nor UO_2224 (O_2224,N_26485,N_27725);
or UO_2225 (O_2225,N_26024,N_28889);
nor UO_2226 (O_2226,N_27450,N_29990);
or UO_2227 (O_2227,N_26211,N_26481);
nand UO_2228 (O_2228,N_27552,N_26863);
xnor UO_2229 (O_2229,N_26200,N_28884);
or UO_2230 (O_2230,N_25070,N_25006);
xor UO_2231 (O_2231,N_27592,N_27227);
or UO_2232 (O_2232,N_27069,N_25474);
or UO_2233 (O_2233,N_25072,N_27038);
or UO_2234 (O_2234,N_25306,N_28437);
nand UO_2235 (O_2235,N_26836,N_25522);
xnor UO_2236 (O_2236,N_29693,N_25514);
xor UO_2237 (O_2237,N_28984,N_27349);
nand UO_2238 (O_2238,N_28325,N_26734);
nor UO_2239 (O_2239,N_26915,N_28820);
and UO_2240 (O_2240,N_26191,N_28754);
nor UO_2241 (O_2241,N_28748,N_26649);
nor UO_2242 (O_2242,N_29415,N_29752);
and UO_2243 (O_2243,N_25025,N_25136);
xor UO_2244 (O_2244,N_26266,N_26699);
xor UO_2245 (O_2245,N_26570,N_28789);
nand UO_2246 (O_2246,N_25827,N_28906);
nor UO_2247 (O_2247,N_25193,N_29569);
xor UO_2248 (O_2248,N_27053,N_29840);
nand UO_2249 (O_2249,N_26394,N_26355);
and UO_2250 (O_2250,N_28417,N_25497);
or UO_2251 (O_2251,N_28303,N_26218);
xnor UO_2252 (O_2252,N_28398,N_25696);
and UO_2253 (O_2253,N_26789,N_25186);
or UO_2254 (O_2254,N_25741,N_29988);
nor UO_2255 (O_2255,N_26331,N_26348);
nand UO_2256 (O_2256,N_27193,N_27532);
nor UO_2257 (O_2257,N_26410,N_29781);
nor UO_2258 (O_2258,N_26214,N_29456);
xor UO_2259 (O_2259,N_27303,N_29962);
nor UO_2260 (O_2260,N_27853,N_29543);
and UO_2261 (O_2261,N_28598,N_26473);
nand UO_2262 (O_2262,N_27482,N_25957);
nor UO_2263 (O_2263,N_28371,N_26823);
nand UO_2264 (O_2264,N_25215,N_25949);
or UO_2265 (O_2265,N_29847,N_27269);
xor UO_2266 (O_2266,N_29722,N_29611);
or UO_2267 (O_2267,N_29386,N_26742);
or UO_2268 (O_2268,N_26883,N_25342);
and UO_2269 (O_2269,N_29033,N_25148);
and UO_2270 (O_2270,N_29331,N_29428);
nor UO_2271 (O_2271,N_29551,N_26128);
xor UO_2272 (O_2272,N_26684,N_26564);
and UO_2273 (O_2273,N_25335,N_26129);
nand UO_2274 (O_2274,N_28264,N_28244);
nor UO_2275 (O_2275,N_28509,N_25532);
xor UO_2276 (O_2276,N_27327,N_28866);
and UO_2277 (O_2277,N_28444,N_29338);
nand UO_2278 (O_2278,N_28587,N_27394);
nand UO_2279 (O_2279,N_25481,N_28080);
nand UO_2280 (O_2280,N_28865,N_29787);
nor UO_2281 (O_2281,N_25214,N_29635);
and UO_2282 (O_2282,N_26716,N_27226);
and UO_2283 (O_2283,N_28036,N_25913);
nor UO_2284 (O_2284,N_29327,N_29267);
nor UO_2285 (O_2285,N_27759,N_29253);
nor UO_2286 (O_2286,N_26035,N_28567);
nand UO_2287 (O_2287,N_27665,N_26539);
nand UO_2288 (O_2288,N_28310,N_27363);
nand UO_2289 (O_2289,N_27993,N_28423);
nor UO_2290 (O_2290,N_27626,N_26726);
nand UO_2291 (O_2291,N_29619,N_29968);
or UO_2292 (O_2292,N_26449,N_29583);
nor UO_2293 (O_2293,N_26371,N_29703);
and UO_2294 (O_2294,N_25486,N_25161);
or UO_2295 (O_2295,N_28885,N_25114);
xnor UO_2296 (O_2296,N_29656,N_25128);
nand UO_2297 (O_2297,N_26943,N_25365);
xor UO_2298 (O_2298,N_26277,N_27381);
and UO_2299 (O_2299,N_25943,N_28240);
nand UO_2300 (O_2300,N_28607,N_25529);
and UO_2301 (O_2301,N_26746,N_28464);
nor UO_2302 (O_2302,N_28203,N_28869);
xor UO_2303 (O_2303,N_29459,N_27839);
nor UO_2304 (O_2304,N_26048,N_27948);
and UO_2305 (O_2305,N_29421,N_26949);
xor UO_2306 (O_2306,N_28511,N_27285);
or UO_2307 (O_2307,N_28059,N_25182);
and UO_2308 (O_2308,N_29417,N_26271);
or UO_2309 (O_2309,N_26495,N_28707);
nor UO_2310 (O_2310,N_28902,N_29215);
nand UO_2311 (O_2311,N_27444,N_29923);
or UO_2312 (O_2312,N_26057,N_27228);
nor UO_2313 (O_2313,N_25564,N_29056);
nand UO_2314 (O_2314,N_28826,N_28069);
nor UO_2315 (O_2315,N_28406,N_29702);
and UO_2316 (O_2316,N_27879,N_25130);
xor UO_2317 (O_2317,N_26687,N_25443);
and UO_2318 (O_2318,N_25387,N_25997);
nor UO_2319 (O_2319,N_28062,N_28136);
nor UO_2320 (O_2320,N_26367,N_25172);
nand UO_2321 (O_2321,N_27018,N_27243);
nor UO_2322 (O_2322,N_25480,N_26624);
or UO_2323 (O_2323,N_27862,N_25064);
nor UO_2324 (O_2324,N_29670,N_26669);
nor UO_2325 (O_2325,N_26950,N_25048);
nand UO_2326 (O_2326,N_27168,N_27258);
or UO_2327 (O_2327,N_27178,N_26045);
and UO_2328 (O_2328,N_27332,N_26899);
nor UO_2329 (O_2329,N_28554,N_27187);
and UO_2330 (O_2330,N_27239,N_27909);
nand UO_2331 (O_2331,N_25572,N_27627);
nand UO_2332 (O_2332,N_29392,N_27857);
nor UO_2333 (O_2333,N_28392,N_28993);
or UO_2334 (O_2334,N_26769,N_25465);
or UO_2335 (O_2335,N_29351,N_26666);
and UO_2336 (O_2336,N_26079,N_29633);
xnor UO_2337 (O_2337,N_25968,N_28288);
nand UO_2338 (O_2338,N_28102,N_29881);
and UO_2339 (O_2339,N_27744,N_25609);
nand UO_2340 (O_2340,N_29679,N_27463);
or UO_2341 (O_2341,N_27222,N_29590);
xnor UO_2342 (O_2342,N_25056,N_29792);
nor UO_2343 (O_2343,N_28418,N_28706);
or UO_2344 (O_2344,N_25561,N_27458);
or UO_2345 (O_2345,N_27743,N_27694);
or UO_2346 (O_2346,N_29194,N_27506);
or UO_2347 (O_2347,N_29951,N_29130);
and UO_2348 (O_2348,N_27074,N_28338);
or UO_2349 (O_2349,N_27718,N_25630);
xor UO_2350 (O_2350,N_25116,N_25250);
xor UO_2351 (O_2351,N_25780,N_25212);
and UO_2352 (O_2352,N_29918,N_28877);
xnor UO_2353 (O_2353,N_26247,N_29318);
xnor UO_2354 (O_2354,N_29487,N_25447);
nand UO_2355 (O_2355,N_29739,N_25805);
nor UO_2356 (O_2356,N_27959,N_28622);
or UO_2357 (O_2357,N_28479,N_26524);
and UO_2358 (O_2358,N_29182,N_26313);
or UO_2359 (O_2359,N_28682,N_29939);
xnor UO_2360 (O_2360,N_26195,N_26736);
and UO_2361 (O_2361,N_28665,N_28504);
xor UO_2362 (O_2362,N_28811,N_28150);
nand UO_2363 (O_2363,N_26828,N_28183);
or UO_2364 (O_2364,N_25218,N_26799);
and UO_2365 (O_2365,N_29024,N_25271);
xor UO_2366 (O_2366,N_26535,N_29826);
nor UO_2367 (O_2367,N_25573,N_29873);
nand UO_2368 (O_2368,N_25041,N_28687);
xor UO_2369 (O_2369,N_29985,N_27899);
nand UO_2370 (O_2370,N_29776,N_25501);
or UO_2371 (O_2371,N_27573,N_28562);
nand UO_2372 (O_2372,N_25477,N_26424);
and UO_2373 (O_2373,N_27809,N_25385);
and UO_2374 (O_2374,N_27818,N_29352);
and UO_2375 (O_2375,N_25208,N_27582);
or UO_2376 (O_2376,N_28430,N_29916);
xnor UO_2377 (O_2377,N_28867,N_27085);
xor UO_2378 (O_2378,N_27945,N_27599);
and UO_2379 (O_2379,N_28039,N_28279);
and UO_2380 (O_2380,N_29010,N_26311);
nand UO_2381 (O_2381,N_25738,N_27372);
and UO_2382 (O_2382,N_29271,N_26818);
xnor UO_2383 (O_2383,N_29060,N_28961);
xor UO_2384 (O_2384,N_26100,N_26385);
nand UO_2385 (O_2385,N_27045,N_26875);
and UO_2386 (O_2386,N_25975,N_27261);
or UO_2387 (O_2387,N_26265,N_25296);
xor UO_2388 (O_2388,N_26923,N_26303);
and UO_2389 (O_2389,N_27878,N_26941);
nand UO_2390 (O_2390,N_29802,N_26963);
xnor UO_2391 (O_2391,N_27276,N_28108);
nand UO_2392 (O_2392,N_29706,N_25539);
xnor UO_2393 (O_2393,N_29719,N_25174);
and UO_2394 (O_2394,N_29299,N_28644);
xnor UO_2395 (O_2395,N_28052,N_28749);
or UO_2396 (O_2396,N_29793,N_25756);
and UO_2397 (O_2397,N_26037,N_26325);
nor UO_2398 (O_2398,N_28868,N_27645);
nor UO_2399 (O_2399,N_27750,N_28686);
xor UO_2400 (O_2400,N_25319,N_29664);
nand UO_2401 (O_2401,N_27171,N_26318);
xor UO_2402 (O_2402,N_29863,N_26042);
xor UO_2403 (O_2403,N_25178,N_29747);
and UO_2404 (O_2404,N_29579,N_27739);
and UO_2405 (O_2405,N_28918,N_25536);
and UO_2406 (O_2406,N_26991,N_29189);
xor UO_2407 (O_2407,N_26417,N_28777);
xor UO_2408 (O_2408,N_28912,N_28933);
nor UO_2409 (O_2409,N_28455,N_28265);
xor UO_2410 (O_2410,N_25206,N_29649);
nor UO_2411 (O_2411,N_27183,N_27192);
nor UO_2412 (O_2412,N_27159,N_27594);
and UO_2413 (O_2413,N_25016,N_25807);
or UO_2414 (O_2414,N_25980,N_28113);
nand UO_2415 (O_2415,N_28426,N_26629);
and UO_2416 (O_2416,N_25947,N_27659);
and UO_2417 (O_2417,N_25785,N_26237);
nand UO_2418 (O_2418,N_25699,N_28549);
and UO_2419 (O_2419,N_25835,N_29053);
and UO_2420 (O_2420,N_26477,N_29170);
xnor UO_2421 (O_2421,N_25951,N_28017);
nand UO_2422 (O_2422,N_27431,N_29356);
or UO_2423 (O_2423,N_27723,N_29885);
nor UO_2424 (O_2424,N_29022,N_26566);
nand UO_2425 (O_2425,N_27109,N_26614);
nand UO_2426 (O_2426,N_28858,N_29655);
nor UO_2427 (O_2427,N_27356,N_26517);
nand UO_2428 (O_2428,N_27788,N_29176);
nand UO_2429 (O_2429,N_27423,N_25051);
xnor UO_2430 (O_2430,N_26279,N_26752);
nand UO_2431 (O_2431,N_26506,N_26762);
and UO_2432 (O_2432,N_29689,N_27671);
nand UO_2433 (O_2433,N_25702,N_26533);
and UO_2434 (O_2434,N_25382,N_29629);
nor UO_2435 (O_2435,N_28788,N_28380);
nor UO_2436 (O_2436,N_28483,N_26356);
nand UO_2437 (O_2437,N_29261,N_26283);
xor UO_2438 (O_2438,N_27449,N_29233);
nor UO_2439 (O_2439,N_28923,N_28089);
nand UO_2440 (O_2440,N_26095,N_29016);
or UO_2441 (O_2441,N_29841,N_26550);
nor UO_2442 (O_2442,N_29909,N_25716);
xnor UO_2443 (O_2443,N_29999,N_29151);
or UO_2444 (O_2444,N_26338,N_27445);
or UO_2445 (O_2445,N_25496,N_29050);
xor UO_2446 (O_2446,N_27663,N_28782);
or UO_2447 (O_2447,N_26285,N_28704);
and UO_2448 (O_2448,N_25170,N_27976);
and UO_2449 (O_2449,N_26656,N_29081);
or UO_2450 (O_2450,N_25228,N_25895);
and UO_2451 (O_2451,N_27143,N_25355);
and UO_2452 (O_2452,N_27995,N_29791);
nor UO_2453 (O_2453,N_25373,N_25667);
xnor UO_2454 (O_2454,N_28298,N_25013);
xor UO_2455 (O_2455,N_29283,N_25879);
and UO_2456 (O_2456,N_25060,N_25852);
nor UO_2457 (O_2457,N_28945,N_25981);
nand UO_2458 (O_2458,N_29891,N_27575);
nand UO_2459 (O_2459,N_28168,N_28362);
or UO_2460 (O_2460,N_28694,N_25440);
nand UO_2461 (O_2461,N_25774,N_29528);
nor UO_2462 (O_2462,N_25848,N_26073);
and UO_2463 (O_2463,N_29315,N_27620);
and UO_2464 (O_2464,N_27437,N_27426);
and UO_2465 (O_2465,N_28367,N_27647);
nor UO_2466 (O_2466,N_27462,N_26425);
xor UO_2467 (O_2467,N_26322,N_28478);
nor UO_2468 (O_2468,N_26213,N_29479);
and UO_2469 (O_2469,N_29872,N_27102);
nand UO_2470 (O_2470,N_25653,N_29134);
xnor UO_2471 (O_2471,N_29800,N_25147);
nor UO_2472 (O_2472,N_28467,N_27357);
xor UO_2473 (O_2473,N_25620,N_25588);
nor UO_2474 (O_2474,N_27237,N_25085);
or UO_2475 (O_2475,N_26164,N_28434);
xor UO_2476 (O_2476,N_29815,N_26887);
or UO_2477 (O_2477,N_25384,N_29251);
and UO_2478 (O_2478,N_28404,N_26194);
xor UO_2479 (O_2479,N_26066,N_27576);
nor UO_2480 (O_2480,N_26051,N_28427);
or UO_2481 (O_2481,N_27202,N_28533);
and UO_2482 (O_2482,N_29952,N_29217);
nand UO_2483 (O_2483,N_25621,N_25802);
or UO_2484 (O_2484,N_28086,N_27772);
xnor UO_2485 (O_2485,N_27343,N_29394);
xor UO_2486 (O_2486,N_28576,N_29862);
xor UO_2487 (O_2487,N_28526,N_25388);
and UO_2488 (O_2488,N_28041,N_25376);
nand UO_2489 (O_2489,N_25458,N_29813);
or UO_2490 (O_2490,N_27405,N_27420);
or UO_2491 (O_2491,N_28128,N_26855);
nor UO_2492 (O_2492,N_27925,N_28133);
and UO_2493 (O_2493,N_28853,N_28321);
nor UO_2494 (O_2494,N_27758,N_28793);
nand UO_2495 (O_2495,N_28861,N_25502);
xnor UO_2496 (O_2496,N_26563,N_26466);
or UO_2497 (O_2497,N_27157,N_25088);
nor UO_2498 (O_2498,N_26514,N_29322);
or UO_2499 (O_2499,N_29128,N_29666);
and UO_2500 (O_2500,N_27185,N_29589);
nand UO_2501 (O_2501,N_29985,N_28878);
and UO_2502 (O_2502,N_28558,N_28313);
nor UO_2503 (O_2503,N_29222,N_26700);
xor UO_2504 (O_2504,N_25694,N_26535);
nor UO_2505 (O_2505,N_27986,N_27225);
xnor UO_2506 (O_2506,N_26224,N_26198);
or UO_2507 (O_2507,N_29205,N_28047);
or UO_2508 (O_2508,N_28825,N_29834);
xnor UO_2509 (O_2509,N_27423,N_25152);
nor UO_2510 (O_2510,N_25745,N_27816);
nor UO_2511 (O_2511,N_26909,N_25549);
or UO_2512 (O_2512,N_26779,N_29278);
or UO_2513 (O_2513,N_28371,N_25434);
and UO_2514 (O_2514,N_26519,N_25316);
nand UO_2515 (O_2515,N_25560,N_27033);
nor UO_2516 (O_2516,N_28438,N_29701);
nor UO_2517 (O_2517,N_25899,N_28497);
xnor UO_2518 (O_2518,N_25465,N_27633);
nor UO_2519 (O_2519,N_26559,N_25002);
xnor UO_2520 (O_2520,N_28796,N_28390);
nor UO_2521 (O_2521,N_28940,N_28178);
and UO_2522 (O_2522,N_28305,N_27352);
or UO_2523 (O_2523,N_29104,N_27982);
nor UO_2524 (O_2524,N_25638,N_29553);
nor UO_2525 (O_2525,N_29658,N_27792);
and UO_2526 (O_2526,N_25474,N_29902);
nor UO_2527 (O_2527,N_26392,N_28212);
nor UO_2528 (O_2528,N_25142,N_28774);
xnor UO_2529 (O_2529,N_25593,N_25998);
nor UO_2530 (O_2530,N_26580,N_29732);
nand UO_2531 (O_2531,N_26635,N_25086);
xnor UO_2532 (O_2532,N_28035,N_26958);
nor UO_2533 (O_2533,N_26638,N_26038);
nand UO_2534 (O_2534,N_28537,N_26153);
xnor UO_2535 (O_2535,N_27399,N_26008);
nor UO_2536 (O_2536,N_28432,N_25975);
nor UO_2537 (O_2537,N_25919,N_28655);
xor UO_2538 (O_2538,N_28908,N_28667);
xnor UO_2539 (O_2539,N_25301,N_29826);
or UO_2540 (O_2540,N_29522,N_27346);
nand UO_2541 (O_2541,N_27219,N_29467);
nand UO_2542 (O_2542,N_29464,N_26045);
nand UO_2543 (O_2543,N_25665,N_26811);
xnor UO_2544 (O_2544,N_25163,N_27629);
and UO_2545 (O_2545,N_28577,N_28681);
nand UO_2546 (O_2546,N_28914,N_27106);
nor UO_2547 (O_2547,N_25335,N_29843);
nor UO_2548 (O_2548,N_29235,N_26961);
xnor UO_2549 (O_2549,N_25180,N_25315);
nand UO_2550 (O_2550,N_27501,N_29649);
xor UO_2551 (O_2551,N_29931,N_25760);
or UO_2552 (O_2552,N_26726,N_26648);
or UO_2553 (O_2553,N_29409,N_29658);
nor UO_2554 (O_2554,N_29304,N_29901);
nand UO_2555 (O_2555,N_26008,N_27786);
nor UO_2556 (O_2556,N_26900,N_28085);
nand UO_2557 (O_2557,N_26544,N_26836);
nor UO_2558 (O_2558,N_27224,N_27855);
nor UO_2559 (O_2559,N_29393,N_28310);
nand UO_2560 (O_2560,N_25082,N_26674);
nor UO_2561 (O_2561,N_28325,N_26433);
xor UO_2562 (O_2562,N_26866,N_25701);
xnor UO_2563 (O_2563,N_26620,N_28075);
nand UO_2564 (O_2564,N_25561,N_29139);
nor UO_2565 (O_2565,N_26079,N_27730);
nand UO_2566 (O_2566,N_28115,N_29329);
nor UO_2567 (O_2567,N_28496,N_28429);
nor UO_2568 (O_2568,N_25102,N_25539);
nand UO_2569 (O_2569,N_29764,N_28478);
nor UO_2570 (O_2570,N_26258,N_28220);
nor UO_2571 (O_2571,N_27497,N_27503);
nand UO_2572 (O_2572,N_25084,N_26811);
nand UO_2573 (O_2573,N_27925,N_29432);
xor UO_2574 (O_2574,N_29932,N_27579);
xor UO_2575 (O_2575,N_26994,N_29618);
xnor UO_2576 (O_2576,N_29951,N_28735);
and UO_2577 (O_2577,N_27326,N_26115);
and UO_2578 (O_2578,N_27567,N_25274);
nor UO_2579 (O_2579,N_26086,N_25873);
or UO_2580 (O_2580,N_29811,N_28126);
nand UO_2581 (O_2581,N_25572,N_28785);
nor UO_2582 (O_2582,N_29986,N_28004);
nor UO_2583 (O_2583,N_26151,N_26734);
nor UO_2584 (O_2584,N_27059,N_28800);
nor UO_2585 (O_2585,N_25203,N_27511);
and UO_2586 (O_2586,N_29032,N_28716);
or UO_2587 (O_2587,N_28192,N_27978);
xnor UO_2588 (O_2588,N_29061,N_28397);
xnor UO_2589 (O_2589,N_25541,N_28321);
nor UO_2590 (O_2590,N_26428,N_27535);
or UO_2591 (O_2591,N_28659,N_26216);
nand UO_2592 (O_2592,N_28243,N_25503);
nor UO_2593 (O_2593,N_29306,N_25745);
nand UO_2594 (O_2594,N_27785,N_28376);
or UO_2595 (O_2595,N_26588,N_26946);
xnor UO_2596 (O_2596,N_27754,N_27472);
xor UO_2597 (O_2597,N_28670,N_25038);
xor UO_2598 (O_2598,N_25610,N_27546);
xor UO_2599 (O_2599,N_29857,N_25565);
and UO_2600 (O_2600,N_28806,N_27778);
xnor UO_2601 (O_2601,N_29082,N_27378);
or UO_2602 (O_2602,N_27489,N_28355);
xnor UO_2603 (O_2603,N_28807,N_26375);
or UO_2604 (O_2604,N_28729,N_28302);
nor UO_2605 (O_2605,N_29793,N_25368);
or UO_2606 (O_2606,N_29954,N_28007);
nand UO_2607 (O_2607,N_27784,N_28886);
xnor UO_2608 (O_2608,N_27046,N_29603);
nor UO_2609 (O_2609,N_29491,N_25102);
nor UO_2610 (O_2610,N_27507,N_27402);
nor UO_2611 (O_2611,N_28405,N_29092);
nand UO_2612 (O_2612,N_29658,N_29983);
xor UO_2613 (O_2613,N_25330,N_29084);
nand UO_2614 (O_2614,N_26941,N_28818);
and UO_2615 (O_2615,N_27407,N_27375);
nand UO_2616 (O_2616,N_29501,N_27617);
nand UO_2617 (O_2617,N_26908,N_28486);
nand UO_2618 (O_2618,N_25125,N_29364);
and UO_2619 (O_2619,N_28586,N_27440);
nand UO_2620 (O_2620,N_28380,N_27310);
nand UO_2621 (O_2621,N_28748,N_28749);
nand UO_2622 (O_2622,N_28752,N_25311);
xor UO_2623 (O_2623,N_26484,N_27669);
xnor UO_2624 (O_2624,N_29800,N_28412);
or UO_2625 (O_2625,N_27680,N_27178);
or UO_2626 (O_2626,N_26545,N_26164);
and UO_2627 (O_2627,N_27227,N_25568);
nor UO_2628 (O_2628,N_29766,N_29762);
nor UO_2629 (O_2629,N_29414,N_28238);
or UO_2630 (O_2630,N_27911,N_27993);
nand UO_2631 (O_2631,N_27369,N_28336);
nand UO_2632 (O_2632,N_25176,N_27318);
nand UO_2633 (O_2633,N_29375,N_26151);
nand UO_2634 (O_2634,N_25392,N_29955);
and UO_2635 (O_2635,N_26524,N_27974);
or UO_2636 (O_2636,N_27970,N_29359);
or UO_2637 (O_2637,N_28444,N_26516);
and UO_2638 (O_2638,N_27448,N_29908);
or UO_2639 (O_2639,N_29528,N_28952);
xor UO_2640 (O_2640,N_25492,N_28000);
or UO_2641 (O_2641,N_27337,N_29798);
nor UO_2642 (O_2642,N_27184,N_27089);
xor UO_2643 (O_2643,N_29386,N_28839);
xnor UO_2644 (O_2644,N_25237,N_28979);
nand UO_2645 (O_2645,N_26009,N_25696);
nor UO_2646 (O_2646,N_26405,N_29490);
and UO_2647 (O_2647,N_25563,N_26625);
nor UO_2648 (O_2648,N_27563,N_29378);
or UO_2649 (O_2649,N_25383,N_29469);
nor UO_2650 (O_2650,N_26006,N_26079);
and UO_2651 (O_2651,N_27108,N_29684);
and UO_2652 (O_2652,N_27241,N_26501);
and UO_2653 (O_2653,N_26966,N_27810);
nor UO_2654 (O_2654,N_25215,N_28958);
nand UO_2655 (O_2655,N_26852,N_28562);
nand UO_2656 (O_2656,N_28922,N_29793);
or UO_2657 (O_2657,N_27568,N_29288);
and UO_2658 (O_2658,N_28788,N_27537);
and UO_2659 (O_2659,N_26545,N_25711);
or UO_2660 (O_2660,N_29021,N_29337);
and UO_2661 (O_2661,N_26155,N_28167);
xor UO_2662 (O_2662,N_29156,N_26228);
nand UO_2663 (O_2663,N_28873,N_25224);
and UO_2664 (O_2664,N_25864,N_27828);
or UO_2665 (O_2665,N_29107,N_26230);
nor UO_2666 (O_2666,N_28406,N_25236);
or UO_2667 (O_2667,N_27403,N_27376);
or UO_2668 (O_2668,N_27339,N_27317);
or UO_2669 (O_2669,N_29837,N_26268);
xnor UO_2670 (O_2670,N_26465,N_25014);
xor UO_2671 (O_2671,N_25904,N_27940);
nor UO_2672 (O_2672,N_25764,N_29932);
or UO_2673 (O_2673,N_26415,N_27701);
or UO_2674 (O_2674,N_29899,N_27141);
and UO_2675 (O_2675,N_27515,N_27208);
nand UO_2676 (O_2676,N_25112,N_26597);
and UO_2677 (O_2677,N_27510,N_26503);
nor UO_2678 (O_2678,N_28824,N_29698);
or UO_2679 (O_2679,N_25054,N_27298);
nor UO_2680 (O_2680,N_29084,N_28856);
xnor UO_2681 (O_2681,N_28705,N_26747);
or UO_2682 (O_2682,N_27256,N_29320);
nand UO_2683 (O_2683,N_28715,N_29030);
nor UO_2684 (O_2684,N_26195,N_27081);
and UO_2685 (O_2685,N_26156,N_25894);
nand UO_2686 (O_2686,N_26319,N_27102);
nor UO_2687 (O_2687,N_27597,N_26233);
nand UO_2688 (O_2688,N_29005,N_29544);
nand UO_2689 (O_2689,N_28661,N_26477);
and UO_2690 (O_2690,N_28909,N_27739);
or UO_2691 (O_2691,N_25114,N_29329);
xor UO_2692 (O_2692,N_25577,N_26921);
and UO_2693 (O_2693,N_29665,N_28787);
and UO_2694 (O_2694,N_25200,N_26632);
or UO_2695 (O_2695,N_26886,N_27356);
nand UO_2696 (O_2696,N_25994,N_27926);
nand UO_2697 (O_2697,N_26514,N_28200);
or UO_2698 (O_2698,N_28400,N_26256);
or UO_2699 (O_2699,N_28297,N_25290);
xor UO_2700 (O_2700,N_27419,N_29998);
or UO_2701 (O_2701,N_28010,N_26170);
or UO_2702 (O_2702,N_28204,N_28086);
nor UO_2703 (O_2703,N_25854,N_25654);
nand UO_2704 (O_2704,N_26677,N_28713);
xor UO_2705 (O_2705,N_26371,N_26757);
xor UO_2706 (O_2706,N_28674,N_29031);
or UO_2707 (O_2707,N_26637,N_28366);
nor UO_2708 (O_2708,N_28681,N_26990);
and UO_2709 (O_2709,N_28038,N_27205);
nor UO_2710 (O_2710,N_25251,N_26278);
nor UO_2711 (O_2711,N_29616,N_29571);
or UO_2712 (O_2712,N_27213,N_25803);
nand UO_2713 (O_2713,N_27665,N_27034);
nand UO_2714 (O_2714,N_28294,N_25900);
xnor UO_2715 (O_2715,N_26445,N_26414);
or UO_2716 (O_2716,N_27670,N_27693);
nand UO_2717 (O_2717,N_26077,N_29211);
nand UO_2718 (O_2718,N_29902,N_28973);
and UO_2719 (O_2719,N_28521,N_26061);
nand UO_2720 (O_2720,N_27592,N_27709);
and UO_2721 (O_2721,N_26691,N_25316);
nor UO_2722 (O_2722,N_28287,N_26518);
nand UO_2723 (O_2723,N_27940,N_27816);
or UO_2724 (O_2724,N_25226,N_27272);
xor UO_2725 (O_2725,N_25895,N_27102);
or UO_2726 (O_2726,N_25947,N_26031);
xor UO_2727 (O_2727,N_25428,N_25831);
xor UO_2728 (O_2728,N_25596,N_28869);
or UO_2729 (O_2729,N_27458,N_25124);
and UO_2730 (O_2730,N_25038,N_28467);
and UO_2731 (O_2731,N_25171,N_28973);
or UO_2732 (O_2732,N_26419,N_26868);
or UO_2733 (O_2733,N_27834,N_28075);
or UO_2734 (O_2734,N_27099,N_26025);
xor UO_2735 (O_2735,N_28666,N_27060);
nor UO_2736 (O_2736,N_29167,N_28094);
nor UO_2737 (O_2737,N_29041,N_26589);
nor UO_2738 (O_2738,N_29931,N_25981);
nand UO_2739 (O_2739,N_29156,N_25200);
and UO_2740 (O_2740,N_27501,N_26214);
xnor UO_2741 (O_2741,N_28424,N_28976);
nor UO_2742 (O_2742,N_27524,N_28579);
and UO_2743 (O_2743,N_28827,N_28980);
nand UO_2744 (O_2744,N_27639,N_29505);
nand UO_2745 (O_2745,N_26355,N_26653);
xnor UO_2746 (O_2746,N_27226,N_28289);
xnor UO_2747 (O_2747,N_29971,N_28401);
and UO_2748 (O_2748,N_27095,N_28809);
or UO_2749 (O_2749,N_28035,N_28920);
or UO_2750 (O_2750,N_26806,N_29268);
or UO_2751 (O_2751,N_28074,N_25682);
xor UO_2752 (O_2752,N_28453,N_29567);
nor UO_2753 (O_2753,N_28007,N_29170);
or UO_2754 (O_2754,N_26174,N_26390);
nor UO_2755 (O_2755,N_28001,N_29025);
and UO_2756 (O_2756,N_29896,N_26076);
xnor UO_2757 (O_2757,N_29401,N_27037);
xnor UO_2758 (O_2758,N_26836,N_29302);
and UO_2759 (O_2759,N_27645,N_26018);
nand UO_2760 (O_2760,N_28233,N_25695);
or UO_2761 (O_2761,N_26524,N_28330);
nor UO_2762 (O_2762,N_27919,N_26065);
and UO_2763 (O_2763,N_28119,N_27459);
nor UO_2764 (O_2764,N_29308,N_29459);
xor UO_2765 (O_2765,N_26757,N_28157);
nand UO_2766 (O_2766,N_29554,N_27484);
xor UO_2767 (O_2767,N_26826,N_29582);
or UO_2768 (O_2768,N_27467,N_27629);
or UO_2769 (O_2769,N_26148,N_27371);
and UO_2770 (O_2770,N_27208,N_25789);
nand UO_2771 (O_2771,N_26751,N_29181);
nor UO_2772 (O_2772,N_27403,N_26029);
and UO_2773 (O_2773,N_27691,N_25939);
or UO_2774 (O_2774,N_29179,N_25315);
nor UO_2775 (O_2775,N_26335,N_25452);
xnor UO_2776 (O_2776,N_27473,N_28420);
xor UO_2777 (O_2777,N_28552,N_28508);
and UO_2778 (O_2778,N_28515,N_26116);
xnor UO_2779 (O_2779,N_29387,N_28297);
nand UO_2780 (O_2780,N_25956,N_28192);
nand UO_2781 (O_2781,N_27465,N_25291);
nand UO_2782 (O_2782,N_29656,N_27448);
xor UO_2783 (O_2783,N_29839,N_29364);
xor UO_2784 (O_2784,N_27455,N_27828);
nand UO_2785 (O_2785,N_26388,N_29962);
xor UO_2786 (O_2786,N_28226,N_25206);
and UO_2787 (O_2787,N_27312,N_25936);
xnor UO_2788 (O_2788,N_25238,N_28046);
and UO_2789 (O_2789,N_28392,N_27116);
nor UO_2790 (O_2790,N_28288,N_29025);
nand UO_2791 (O_2791,N_27726,N_25718);
nand UO_2792 (O_2792,N_28282,N_26300);
nor UO_2793 (O_2793,N_26235,N_25334);
and UO_2794 (O_2794,N_26717,N_27173);
nor UO_2795 (O_2795,N_28777,N_29956);
nor UO_2796 (O_2796,N_26526,N_26202);
nand UO_2797 (O_2797,N_26315,N_27003);
or UO_2798 (O_2798,N_25551,N_25286);
or UO_2799 (O_2799,N_26547,N_28175);
nand UO_2800 (O_2800,N_29021,N_29354);
nor UO_2801 (O_2801,N_27759,N_26398);
nor UO_2802 (O_2802,N_28496,N_27432);
or UO_2803 (O_2803,N_25606,N_28708);
or UO_2804 (O_2804,N_28108,N_28743);
or UO_2805 (O_2805,N_29420,N_26475);
or UO_2806 (O_2806,N_27937,N_25615);
and UO_2807 (O_2807,N_29759,N_25415);
and UO_2808 (O_2808,N_28034,N_28355);
xor UO_2809 (O_2809,N_25098,N_28372);
or UO_2810 (O_2810,N_27242,N_27795);
nor UO_2811 (O_2811,N_27891,N_26436);
nand UO_2812 (O_2812,N_26557,N_26492);
xnor UO_2813 (O_2813,N_26175,N_25645);
nand UO_2814 (O_2814,N_29492,N_28630);
nand UO_2815 (O_2815,N_25233,N_25597);
xnor UO_2816 (O_2816,N_26495,N_28051);
xnor UO_2817 (O_2817,N_28626,N_28738);
and UO_2818 (O_2818,N_29756,N_28468);
nand UO_2819 (O_2819,N_28789,N_25777);
and UO_2820 (O_2820,N_28540,N_25748);
xor UO_2821 (O_2821,N_28044,N_27291);
and UO_2822 (O_2822,N_27524,N_29723);
nand UO_2823 (O_2823,N_25541,N_26224);
nor UO_2824 (O_2824,N_28381,N_26943);
nor UO_2825 (O_2825,N_29284,N_26569);
nand UO_2826 (O_2826,N_27467,N_26285);
nor UO_2827 (O_2827,N_28501,N_29001);
xor UO_2828 (O_2828,N_29304,N_27910);
nor UO_2829 (O_2829,N_29217,N_27628);
xor UO_2830 (O_2830,N_26354,N_29018);
xnor UO_2831 (O_2831,N_27547,N_29865);
nor UO_2832 (O_2832,N_29925,N_29786);
nand UO_2833 (O_2833,N_27236,N_29665);
or UO_2834 (O_2834,N_26881,N_25793);
xor UO_2835 (O_2835,N_26765,N_28455);
xnor UO_2836 (O_2836,N_29386,N_28841);
xnor UO_2837 (O_2837,N_27407,N_27556);
or UO_2838 (O_2838,N_27106,N_27271);
xor UO_2839 (O_2839,N_25390,N_28722);
nand UO_2840 (O_2840,N_25716,N_26204);
or UO_2841 (O_2841,N_26861,N_25295);
xnor UO_2842 (O_2842,N_26529,N_25004);
or UO_2843 (O_2843,N_26464,N_28301);
xnor UO_2844 (O_2844,N_29396,N_26325);
xor UO_2845 (O_2845,N_26999,N_29651);
or UO_2846 (O_2846,N_25856,N_28134);
nand UO_2847 (O_2847,N_26735,N_26082);
nand UO_2848 (O_2848,N_26186,N_25758);
and UO_2849 (O_2849,N_29683,N_26196);
nand UO_2850 (O_2850,N_25120,N_27934);
nand UO_2851 (O_2851,N_28656,N_29290);
and UO_2852 (O_2852,N_29190,N_26670);
nor UO_2853 (O_2853,N_28622,N_28720);
nor UO_2854 (O_2854,N_26285,N_28888);
xor UO_2855 (O_2855,N_26043,N_26875);
xor UO_2856 (O_2856,N_28201,N_26525);
nand UO_2857 (O_2857,N_28312,N_29797);
nand UO_2858 (O_2858,N_29276,N_26866);
nor UO_2859 (O_2859,N_29123,N_26930);
nor UO_2860 (O_2860,N_26798,N_29907);
and UO_2861 (O_2861,N_28575,N_28054);
or UO_2862 (O_2862,N_26726,N_27692);
xnor UO_2863 (O_2863,N_28999,N_27124);
and UO_2864 (O_2864,N_28008,N_29936);
xor UO_2865 (O_2865,N_26376,N_29649);
or UO_2866 (O_2866,N_26116,N_25928);
nand UO_2867 (O_2867,N_27809,N_25655);
xnor UO_2868 (O_2868,N_28394,N_26248);
xor UO_2869 (O_2869,N_25758,N_25486);
xor UO_2870 (O_2870,N_27013,N_25548);
or UO_2871 (O_2871,N_25053,N_26615);
or UO_2872 (O_2872,N_27107,N_27378);
xnor UO_2873 (O_2873,N_26287,N_27846);
xor UO_2874 (O_2874,N_28608,N_26118);
nand UO_2875 (O_2875,N_25884,N_28401);
or UO_2876 (O_2876,N_29265,N_27356);
or UO_2877 (O_2877,N_27821,N_26377);
xnor UO_2878 (O_2878,N_26347,N_27004);
nor UO_2879 (O_2879,N_28426,N_28616);
xnor UO_2880 (O_2880,N_29359,N_26142);
nand UO_2881 (O_2881,N_27536,N_27041);
xor UO_2882 (O_2882,N_29887,N_27489);
and UO_2883 (O_2883,N_26870,N_25329);
nor UO_2884 (O_2884,N_27862,N_25898);
xor UO_2885 (O_2885,N_28092,N_28351);
nor UO_2886 (O_2886,N_27995,N_26594);
nor UO_2887 (O_2887,N_26909,N_26772);
nor UO_2888 (O_2888,N_27798,N_25082);
xor UO_2889 (O_2889,N_28800,N_28040);
xnor UO_2890 (O_2890,N_26956,N_29539);
xnor UO_2891 (O_2891,N_25716,N_28059);
and UO_2892 (O_2892,N_29795,N_26869);
and UO_2893 (O_2893,N_28969,N_29853);
nor UO_2894 (O_2894,N_26834,N_25971);
xor UO_2895 (O_2895,N_28529,N_29894);
and UO_2896 (O_2896,N_29947,N_28682);
nor UO_2897 (O_2897,N_28266,N_26067);
and UO_2898 (O_2898,N_28165,N_28769);
or UO_2899 (O_2899,N_28656,N_27799);
or UO_2900 (O_2900,N_26691,N_26621);
nor UO_2901 (O_2901,N_26845,N_27467);
and UO_2902 (O_2902,N_27499,N_27928);
and UO_2903 (O_2903,N_29229,N_26311);
xnor UO_2904 (O_2904,N_25958,N_29712);
and UO_2905 (O_2905,N_29208,N_25600);
xor UO_2906 (O_2906,N_29591,N_25818);
or UO_2907 (O_2907,N_27274,N_28330);
nand UO_2908 (O_2908,N_29178,N_27774);
and UO_2909 (O_2909,N_25969,N_26199);
xnor UO_2910 (O_2910,N_28254,N_29662);
nand UO_2911 (O_2911,N_28057,N_27697);
and UO_2912 (O_2912,N_29292,N_25916);
xnor UO_2913 (O_2913,N_26747,N_29467);
nand UO_2914 (O_2914,N_25173,N_25729);
nor UO_2915 (O_2915,N_28396,N_27390);
nor UO_2916 (O_2916,N_28429,N_29369);
xor UO_2917 (O_2917,N_25026,N_25701);
or UO_2918 (O_2918,N_26611,N_27233);
and UO_2919 (O_2919,N_27802,N_26905);
nand UO_2920 (O_2920,N_29801,N_29264);
nand UO_2921 (O_2921,N_28331,N_26482);
or UO_2922 (O_2922,N_28112,N_25661);
nand UO_2923 (O_2923,N_28690,N_29745);
nand UO_2924 (O_2924,N_27930,N_29036);
or UO_2925 (O_2925,N_26940,N_29498);
or UO_2926 (O_2926,N_26613,N_26289);
and UO_2927 (O_2927,N_29022,N_25562);
and UO_2928 (O_2928,N_26315,N_27080);
or UO_2929 (O_2929,N_27994,N_29868);
nor UO_2930 (O_2930,N_26609,N_28026);
nand UO_2931 (O_2931,N_26883,N_25765);
nor UO_2932 (O_2932,N_27631,N_25520);
xnor UO_2933 (O_2933,N_26161,N_25301);
and UO_2934 (O_2934,N_25560,N_26462);
nand UO_2935 (O_2935,N_27743,N_27781);
nor UO_2936 (O_2936,N_26559,N_25819);
nor UO_2937 (O_2937,N_27134,N_28016);
xnor UO_2938 (O_2938,N_27107,N_29609);
nor UO_2939 (O_2939,N_25033,N_26320);
xnor UO_2940 (O_2940,N_25838,N_26873);
nor UO_2941 (O_2941,N_29813,N_29139);
nand UO_2942 (O_2942,N_25082,N_29043);
xnor UO_2943 (O_2943,N_29787,N_27301);
xor UO_2944 (O_2944,N_28162,N_29681);
xnor UO_2945 (O_2945,N_27014,N_27842);
nor UO_2946 (O_2946,N_27961,N_26363);
nor UO_2947 (O_2947,N_27929,N_26642);
or UO_2948 (O_2948,N_25734,N_28587);
xor UO_2949 (O_2949,N_26753,N_26973);
nor UO_2950 (O_2950,N_27880,N_27822);
nor UO_2951 (O_2951,N_26294,N_26987);
nand UO_2952 (O_2952,N_29121,N_29260);
and UO_2953 (O_2953,N_27441,N_29656);
xor UO_2954 (O_2954,N_27310,N_27347);
or UO_2955 (O_2955,N_26169,N_29485);
and UO_2956 (O_2956,N_25203,N_27950);
nand UO_2957 (O_2957,N_27397,N_28774);
xnor UO_2958 (O_2958,N_26135,N_28138);
nor UO_2959 (O_2959,N_25101,N_26210);
xor UO_2960 (O_2960,N_27133,N_27969);
nor UO_2961 (O_2961,N_29080,N_29766);
xor UO_2962 (O_2962,N_27774,N_25103);
xor UO_2963 (O_2963,N_27004,N_29516);
xor UO_2964 (O_2964,N_25940,N_25038);
nor UO_2965 (O_2965,N_27173,N_28731);
nor UO_2966 (O_2966,N_25013,N_29136);
or UO_2967 (O_2967,N_29080,N_29844);
or UO_2968 (O_2968,N_25199,N_28697);
xor UO_2969 (O_2969,N_29906,N_25497);
nor UO_2970 (O_2970,N_28167,N_25273);
and UO_2971 (O_2971,N_25295,N_26183);
xnor UO_2972 (O_2972,N_25400,N_28705);
or UO_2973 (O_2973,N_27827,N_26722);
or UO_2974 (O_2974,N_25354,N_27557);
and UO_2975 (O_2975,N_29748,N_29675);
nand UO_2976 (O_2976,N_28427,N_28716);
nand UO_2977 (O_2977,N_28099,N_26097);
xnor UO_2978 (O_2978,N_29805,N_26906);
nor UO_2979 (O_2979,N_27575,N_29003);
nand UO_2980 (O_2980,N_26850,N_26051);
nor UO_2981 (O_2981,N_28471,N_28984);
nor UO_2982 (O_2982,N_26713,N_29296);
xor UO_2983 (O_2983,N_27051,N_29753);
nand UO_2984 (O_2984,N_25736,N_26796);
and UO_2985 (O_2985,N_27036,N_26837);
and UO_2986 (O_2986,N_28686,N_25720);
xor UO_2987 (O_2987,N_29668,N_26424);
xor UO_2988 (O_2988,N_26044,N_25397);
xnor UO_2989 (O_2989,N_28413,N_27454);
nor UO_2990 (O_2990,N_29276,N_29243);
and UO_2991 (O_2991,N_29826,N_26916);
nor UO_2992 (O_2992,N_29851,N_27190);
nand UO_2993 (O_2993,N_25279,N_26177);
and UO_2994 (O_2994,N_27715,N_28971);
or UO_2995 (O_2995,N_27302,N_29724);
or UO_2996 (O_2996,N_28331,N_29024);
nor UO_2997 (O_2997,N_28416,N_29020);
xnor UO_2998 (O_2998,N_26677,N_29355);
and UO_2999 (O_2999,N_26615,N_26406);
and UO_3000 (O_3000,N_25953,N_26827);
nand UO_3001 (O_3001,N_29671,N_27757);
nand UO_3002 (O_3002,N_27415,N_26895);
nor UO_3003 (O_3003,N_28912,N_26323);
and UO_3004 (O_3004,N_28698,N_25922);
and UO_3005 (O_3005,N_25971,N_29987);
and UO_3006 (O_3006,N_28065,N_26774);
nor UO_3007 (O_3007,N_27178,N_29869);
xnor UO_3008 (O_3008,N_28583,N_26034);
and UO_3009 (O_3009,N_27476,N_26416);
nand UO_3010 (O_3010,N_29409,N_29784);
nor UO_3011 (O_3011,N_26125,N_27856);
and UO_3012 (O_3012,N_28725,N_27714);
nand UO_3013 (O_3013,N_28780,N_27722);
nor UO_3014 (O_3014,N_25376,N_29987);
nor UO_3015 (O_3015,N_25162,N_26113);
nand UO_3016 (O_3016,N_27704,N_25186);
and UO_3017 (O_3017,N_26614,N_27049);
nor UO_3018 (O_3018,N_28794,N_25673);
and UO_3019 (O_3019,N_25274,N_28214);
nand UO_3020 (O_3020,N_28395,N_29618);
or UO_3021 (O_3021,N_25566,N_29330);
xnor UO_3022 (O_3022,N_26261,N_28769);
nor UO_3023 (O_3023,N_28201,N_28475);
nor UO_3024 (O_3024,N_25050,N_27608);
and UO_3025 (O_3025,N_26359,N_29385);
or UO_3026 (O_3026,N_25099,N_29904);
nand UO_3027 (O_3027,N_29143,N_28300);
nand UO_3028 (O_3028,N_25911,N_26733);
and UO_3029 (O_3029,N_25542,N_25599);
xnor UO_3030 (O_3030,N_26163,N_26427);
nand UO_3031 (O_3031,N_25564,N_25155);
nand UO_3032 (O_3032,N_25414,N_26073);
xor UO_3033 (O_3033,N_26204,N_28690);
nand UO_3034 (O_3034,N_28777,N_28042);
or UO_3035 (O_3035,N_27439,N_27159);
xnor UO_3036 (O_3036,N_28230,N_27175);
nor UO_3037 (O_3037,N_25315,N_28751);
xor UO_3038 (O_3038,N_25764,N_29996);
nor UO_3039 (O_3039,N_26391,N_25355);
or UO_3040 (O_3040,N_26077,N_29111);
xnor UO_3041 (O_3041,N_29196,N_27388);
nor UO_3042 (O_3042,N_29305,N_25223);
xnor UO_3043 (O_3043,N_26994,N_28375);
or UO_3044 (O_3044,N_26326,N_27239);
nor UO_3045 (O_3045,N_25002,N_28337);
nand UO_3046 (O_3046,N_26262,N_26681);
xnor UO_3047 (O_3047,N_28084,N_27413);
xor UO_3048 (O_3048,N_26273,N_27202);
or UO_3049 (O_3049,N_29789,N_25018);
and UO_3050 (O_3050,N_25527,N_26088);
nand UO_3051 (O_3051,N_26635,N_29202);
xnor UO_3052 (O_3052,N_28427,N_27460);
nand UO_3053 (O_3053,N_27003,N_27449);
or UO_3054 (O_3054,N_26461,N_27688);
nand UO_3055 (O_3055,N_29508,N_26995);
or UO_3056 (O_3056,N_27876,N_27496);
or UO_3057 (O_3057,N_25787,N_25072);
xnor UO_3058 (O_3058,N_26753,N_27235);
xnor UO_3059 (O_3059,N_28118,N_26531);
xnor UO_3060 (O_3060,N_28395,N_27185);
and UO_3061 (O_3061,N_29731,N_25458);
and UO_3062 (O_3062,N_29415,N_25245);
nor UO_3063 (O_3063,N_29101,N_27302);
or UO_3064 (O_3064,N_25613,N_28651);
and UO_3065 (O_3065,N_26250,N_27395);
or UO_3066 (O_3066,N_25330,N_28435);
nand UO_3067 (O_3067,N_28268,N_29919);
and UO_3068 (O_3068,N_25233,N_28184);
nor UO_3069 (O_3069,N_26393,N_27267);
and UO_3070 (O_3070,N_25970,N_28514);
and UO_3071 (O_3071,N_28206,N_29922);
nand UO_3072 (O_3072,N_26532,N_29268);
or UO_3073 (O_3073,N_26172,N_27802);
and UO_3074 (O_3074,N_27145,N_27138);
nand UO_3075 (O_3075,N_25193,N_28371);
nor UO_3076 (O_3076,N_26545,N_29771);
nand UO_3077 (O_3077,N_27364,N_27998);
nor UO_3078 (O_3078,N_29734,N_28172);
nand UO_3079 (O_3079,N_28889,N_29287);
xor UO_3080 (O_3080,N_25670,N_25733);
or UO_3081 (O_3081,N_26690,N_25474);
or UO_3082 (O_3082,N_29137,N_27455);
xor UO_3083 (O_3083,N_29247,N_26959);
nor UO_3084 (O_3084,N_28699,N_27111);
nand UO_3085 (O_3085,N_27056,N_28024);
and UO_3086 (O_3086,N_28908,N_28230);
and UO_3087 (O_3087,N_27500,N_25665);
or UO_3088 (O_3088,N_25398,N_29870);
and UO_3089 (O_3089,N_25869,N_28045);
nand UO_3090 (O_3090,N_26887,N_25367);
nor UO_3091 (O_3091,N_26288,N_29086);
or UO_3092 (O_3092,N_28369,N_28385);
nor UO_3093 (O_3093,N_28892,N_28403);
and UO_3094 (O_3094,N_29492,N_26863);
and UO_3095 (O_3095,N_26154,N_29835);
nand UO_3096 (O_3096,N_29061,N_27606);
xnor UO_3097 (O_3097,N_28650,N_26786);
nand UO_3098 (O_3098,N_29796,N_27186);
and UO_3099 (O_3099,N_25528,N_27864);
nor UO_3100 (O_3100,N_26404,N_27964);
xor UO_3101 (O_3101,N_29767,N_25754);
xor UO_3102 (O_3102,N_28967,N_29965);
xnor UO_3103 (O_3103,N_26835,N_26967);
xnor UO_3104 (O_3104,N_29556,N_28252);
or UO_3105 (O_3105,N_25281,N_29527);
and UO_3106 (O_3106,N_29328,N_29661);
or UO_3107 (O_3107,N_25432,N_29011);
nor UO_3108 (O_3108,N_25126,N_26679);
xnor UO_3109 (O_3109,N_26404,N_26226);
nor UO_3110 (O_3110,N_27416,N_29704);
nand UO_3111 (O_3111,N_27299,N_28324);
nor UO_3112 (O_3112,N_29569,N_25935);
nor UO_3113 (O_3113,N_29793,N_25369);
and UO_3114 (O_3114,N_28429,N_26210);
nand UO_3115 (O_3115,N_27882,N_27788);
and UO_3116 (O_3116,N_25659,N_28774);
and UO_3117 (O_3117,N_27816,N_28917);
nor UO_3118 (O_3118,N_26348,N_27552);
nand UO_3119 (O_3119,N_25927,N_29603);
or UO_3120 (O_3120,N_27678,N_25603);
and UO_3121 (O_3121,N_27115,N_27522);
or UO_3122 (O_3122,N_27083,N_28209);
nor UO_3123 (O_3123,N_28330,N_29635);
or UO_3124 (O_3124,N_26937,N_27774);
xnor UO_3125 (O_3125,N_25077,N_28624);
xnor UO_3126 (O_3126,N_29324,N_27550);
nand UO_3127 (O_3127,N_29993,N_25998);
nand UO_3128 (O_3128,N_26473,N_28634);
xnor UO_3129 (O_3129,N_29981,N_28214);
nand UO_3130 (O_3130,N_29832,N_28336);
xnor UO_3131 (O_3131,N_27414,N_27629);
nand UO_3132 (O_3132,N_26909,N_27068);
nand UO_3133 (O_3133,N_29284,N_28700);
nand UO_3134 (O_3134,N_27655,N_25165);
and UO_3135 (O_3135,N_28900,N_29690);
nor UO_3136 (O_3136,N_26334,N_27730);
nand UO_3137 (O_3137,N_28496,N_26677);
xnor UO_3138 (O_3138,N_27754,N_29178);
nand UO_3139 (O_3139,N_27118,N_28175);
nor UO_3140 (O_3140,N_26050,N_26680);
nor UO_3141 (O_3141,N_26701,N_25339);
or UO_3142 (O_3142,N_27804,N_26499);
or UO_3143 (O_3143,N_28878,N_25931);
and UO_3144 (O_3144,N_25505,N_28299);
nor UO_3145 (O_3145,N_29407,N_27384);
or UO_3146 (O_3146,N_25903,N_25946);
xor UO_3147 (O_3147,N_25796,N_28461);
or UO_3148 (O_3148,N_26620,N_27101);
and UO_3149 (O_3149,N_29756,N_28603);
nor UO_3150 (O_3150,N_27992,N_29096);
or UO_3151 (O_3151,N_28272,N_27722);
nor UO_3152 (O_3152,N_27414,N_28680);
and UO_3153 (O_3153,N_27131,N_27052);
nor UO_3154 (O_3154,N_27279,N_25478);
xnor UO_3155 (O_3155,N_26889,N_27374);
nor UO_3156 (O_3156,N_25639,N_27389);
nand UO_3157 (O_3157,N_26438,N_25227);
or UO_3158 (O_3158,N_26204,N_27081);
nand UO_3159 (O_3159,N_25619,N_25988);
nand UO_3160 (O_3160,N_25628,N_29637);
xor UO_3161 (O_3161,N_29721,N_25490);
xnor UO_3162 (O_3162,N_25662,N_27029);
xor UO_3163 (O_3163,N_28706,N_27536);
nand UO_3164 (O_3164,N_29304,N_26089);
and UO_3165 (O_3165,N_28189,N_27112);
xnor UO_3166 (O_3166,N_27554,N_29305);
or UO_3167 (O_3167,N_29163,N_28067);
and UO_3168 (O_3168,N_25202,N_26821);
nand UO_3169 (O_3169,N_27982,N_26522);
nand UO_3170 (O_3170,N_27673,N_26908);
and UO_3171 (O_3171,N_25049,N_27357);
or UO_3172 (O_3172,N_26171,N_27976);
or UO_3173 (O_3173,N_29655,N_28324);
nor UO_3174 (O_3174,N_27009,N_26334);
or UO_3175 (O_3175,N_28523,N_28688);
nand UO_3176 (O_3176,N_25263,N_27884);
nand UO_3177 (O_3177,N_26259,N_28147);
xnor UO_3178 (O_3178,N_28874,N_25922);
or UO_3179 (O_3179,N_29065,N_26890);
nand UO_3180 (O_3180,N_28482,N_27706);
nor UO_3181 (O_3181,N_29316,N_28646);
xnor UO_3182 (O_3182,N_25926,N_28768);
nor UO_3183 (O_3183,N_29455,N_29317);
or UO_3184 (O_3184,N_27250,N_29065);
xor UO_3185 (O_3185,N_29300,N_27361);
or UO_3186 (O_3186,N_25379,N_29831);
or UO_3187 (O_3187,N_29038,N_27265);
nor UO_3188 (O_3188,N_29083,N_27431);
xnor UO_3189 (O_3189,N_25492,N_27806);
or UO_3190 (O_3190,N_27159,N_28623);
and UO_3191 (O_3191,N_27990,N_26662);
or UO_3192 (O_3192,N_26635,N_25157);
and UO_3193 (O_3193,N_28289,N_26423);
nand UO_3194 (O_3194,N_28652,N_28312);
xor UO_3195 (O_3195,N_29122,N_28421);
xor UO_3196 (O_3196,N_26574,N_28189);
nor UO_3197 (O_3197,N_29320,N_25943);
or UO_3198 (O_3198,N_29365,N_28206);
and UO_3199 (O_3199,N_25541,N_28697);
nor UO_3200 (O_3200,N_27985,N_29773);
and UO_3201 (O_3201,N_25776,N_27297);
nor UO_3202 (O_3202,N_29046,N_25533);
or UO_3203 (O_3203,N_26220,N_25968);
nand UO_3204 (O_3204,N_25084,N_29382);
xor UO_3205 (O_3205,N_27827,N_28895);
nor UO_3206 (O_3206,N_26120,N_28566);
or UO_3207 (O_3207,N_26803,N_29578);
or UO_3208 (O_3208,N_28739,N_27179);
nand UO_3209 (O_3209,N_27333,N_25432);
or UO_3210 (O_3210,N_28544,N_26508);
xor UO_3211 (O_3211,N_26459,N_28372);
nand UO_3212 (O_3212,N_28688,N_27580);
nand UO_3213 (O_3213,N_28178,N_29503);
nand UO_3214 (O_3214,N_29230,N_28679);
and UO_3215 (O_3215,N_28114,N_25433);
nor UO_3216 (O_3216,N_26420,N_25398);
and UO_3217 (O_3217,N_25493,N_27719);
and UO_3218 (O_3218,N_27860,N_28494);
xor UO_3219 (O_3219,N_26345,N_27896);
xnor UO_3220 (O_3220,N_26145,N_29651);
xnor UO_3221 (O_3221,N_27312,N_27470);
xor UO_3222 (O_3222,N_29896,N_25304);
or UO_3223 (O_3223,N_26049,N_27529);
xnor UO_3224 (O_3224,N_28358,N_29783);
nand UO_3225 (O_3225,N_25372,N_28779);
xnor UO_3226 (O_3226,N_27602,N_29795);
xnor UO_3227 (O_3227,N_28911,N_27376);
or UO_3228 (O_3228,N_29177,N_25919);
nor UO_3229 (O_3229,N_28405,N_29999);
nand UO_3230 (O_3230,N_28007,N_26532);
nand UO_3231 (O_3231,N_27986,N_25444);
and UO_3232 (O_3232,N_25817,N_29745);
nor UO_3233 (O_3233,N_29911,N_28898);
xnor UO_3234 (O_3234,N_25320,N_29177);
and UO_3235 (O_3235,N_29844,N_27424);
and UO_3236 (O_3236,N_26221,N_28867);
or UO_3237 (O_3237,N_26610,N_27518);
xnor UO_3238 (O_3238,N_28146,N_27880);
or UO_3239 (O_3239,N_29475,N_28488);
or UO_3240 (O_3240,N_29708,N_27214);
nor UO_3241 (O_3241,N_29826,N_27957);
and UO_3242 (O_3242,N_26798,N_27896);
xnor UO_3243 (O_3243,N_29996,N_27244);
nor UO_3244 (O_3244,N_28233,N_26195);
or UO_3245 (O_3245,N_29135,N_25076);
and UO_3246 (O_3246,N_27550,N_29485);
nor UO_3247 (O_3247,N_25866,N_26746);
or UO_3248 (O_3248,N_29014,N_26764);
and UO_3249 (O_3249,N_26437,N_28894);
nand UO_3250 (O_3250,N_29551,N_29092);
nand UO_3251 (O_3251,N_26422,N_25154);
nand UO_3252 (O_3252,N_27474,N_29560);
or UO_3253 (O_3253,N_26942,N_29741);
xor UO_3254 (O_3254,N_26556,N_29690);
nand UO_3255 (O_3255,N_28742,N_28578);
and UO_3256 (O_3256,N_29487,N_27596);
xnor UO_3257 (O_3257,N_26099,N_26230);
nand UO_3258 (O_3258,N_28132,N_28249);
xor UO_3259 (O_3259,N_28939,N_29857);
nand UO_3260 (O_3260,N_25742,N_29085);
xor UO_3261 (O_3261,N_27750,N_27793);
or UO_3262 (O_3262,N_29882,N_27022);
xnor UO_3263 (O_3263,N_27492,N_27790);
or UO_3264 (O_3264,N_26704,N_29770);
or UO_3265 (O_3265,N_28257,N_28820);
nor UO_3266 (O_3266,N_29532,N_25364);
nor UO_3267 (O_3267,N_25382,N_28669);
xnor UO_3268 (O_3268,N_29088,N_25471);
nor UO_3269 (O_3269,N_25978,N_25294);
or UO_3270 (O_3270,N_25023,N_29818);
nand UO_3271 (O_3271,N_27845,N_28850);
and UO_3272 (O_3272,N_26814,N_25776);
or UO_3273 (O_3273,N_28272,N_25290);
nand UO_3274 (O_3274,N_29560,N_28599);
or UO_3275 (O_3275,N_26177,N_26351);
nand UO_3276 (O_3276,N_29118,N_29642);
nand UO_3277 (O_3277,N_27261,N_25455);
xnor UO_3278 (O_3278,N_29841,N_25831);
and UO_3279 (O_3279,N_26929,N_27079);
and UO_3280 (O_3280,N_26909,N_29622);
nor UO_3281 (O_3281,N_28282,N_29369);
nand UO_3282 (O_3282,N_25512,N_27765);
and UO_3283 (O_3283,N_26644,N_29520);
or UO_3284 (O_3284,N_25991,N_29710);
and UO_3285 (O_3285,N_29002,N_28082);
xor UO_3286 (O_3286,N_25986,N_26890);
nor UO_3287 (O_3287,N_29368,N_26182);
and UO_3288 (O_3288,N_29197,N_25787);
or UO_3289 (O_3289,N_26182,N_27885);
or UO_3290 (O_3290,N_25967,N_28234);
or UO_3291 (O_3291,N_25587,N_25904);
xor UO_3292 (O_3292,N_25443,N_26308);
xnor UO_3293 (O_3293,N_26318,N_28966);
nand UO_3294 (O_3294,N_27526,N_25304);
nor UO_3295 (O_3295,N_25586,N_28054);
or UO_3296 (O_3296,N_29219,N_29119);
nor UO_3297 (O_3297,N_26323,N_28894);
xnor UO_3298 (O_3298,N_27938,N_26222);
or UO_3299 (O_3299,N_27902,N_25181);
and UO_3300 (O_3300,N_28537,N_29549);
nand UO_3301 (O_3301,N_26086,N_26337);
and UO_3302 (O_3302,N_25136,N_28626);
nand UO_3303 (O_3303,N_29552,N_29166);
nor UO_3304 (O_3304,N_29286,N_28196);
xor UO_3305 (O_3305,N_25506,N_27682);
nand UO_3306 (O_3306,N_26262,N_27759);
xor UO_3307 (O_3307,N_25179,N_27062);
xnor UO_3308 (O_3308,N_29835,N_26668);
and UO_3309 (O_3309,N_28876,N_28492);
xor UO_3310 (O_3310,N_25516,N_26360);
or UO_3311 (O_3311,N_29868,N_29587);
or UO_3312 (O_3312,N_28872,N_25565);
nand UO_3313 (O_3313,N_29778,N_27139);
xnor UO_3314 (O_3314,N_25434,N_28608);
xor UO_3315 (O_3315,N_27897,N_26796);
and UO_3316 (O_3316,N_27032,N_27540);
and UO_3317 (O_3317,N_29554,N_27688);
or UO_3318 (O_3318,N_28408,N_25896);
nand UO_3319 (O_3319,N_29841,N_25999);
xor UO_3320 (O_3320,N_27288,N_26731);
and UO_3321 (O_3321,N_26994,N_27245);
or UO_3322 (O_3322,N_27414,N_29291);
nor UO_3323 (O_3323,N_29277,N_28031);
or UO_3324 (O_3324,N_27123,N_29197);
or UO_3325 (O_3325,N_29457,N_29255);
nand UO_3326 (O_3326,N_29277,N_25082);
or UO_3327 (O_3327,N_26476,N_28464);
nor UO_3328 (O_3328,N_26792,N_27207);
xnor UO_3329 (O_3329,N_27352,N_28405);
or UO_3330 (O_3330,N_28017,N_27237);
nand UO_3331 (O_3331,N_25245,N_29999);
nand UO_3332 (O_3332,N_25096,N_28649);
and UO_3333 (O_3333,N_28163,N_25227);
nor UO_3334 (O_3334,N_26913,N_25397);
xor UO_3335 (O_3335,N_25651,N_26159);
xor UO_3336 (O_3336,N_27259,N_26194);
nand UO_3337 (O_3337,N_29142,N_26750);
nand UO_3338 (O_3338,N_27637,N_26773);
nand UO_3339 (O_3339,N_28459,N_28386);
or UO_3340 (O_3340,N_28947,N_27358);
nand UO_3341 (O_3341,N_27919,N_29637);
and UO_3342 (O_3342,N_28417,N_27755);
and UO_3343 (O_3343,N_29259,N_25336);
nor UO_3344 (O_3344,N_26641,N_26801);
nand UO_3345 (O_3345,N_28271,N_25002);
nand UO_3346 (O_3346,N_25685,N_29568);
or UO_3347 (O_3347,N_27578,N_25789);
or UO_3348 (O_3348,N_28143,N_26499);
nand UO_3349 (O_3349,N_29986,N_29512);
nor UO_3350 (O_3350,N_28283,N_27884);
and UO_3351 (O_3351,N_26226,N_27558);
and UO_3352 (O_3352,N_29300,N_26282);
and UO_3353 (O_3353,N_26747,N_29166);
nand UO_3354 (O_3354,N_29118,N_27421);
nor UO_3355 (O_3355,N_26327,N_27130);
nor UO_3356 (O_3356,N_26029,N_27406);
nand UO_3357 (O_3357,N_26718,N_27399);
or UO_3358 (O_3358,N_26542,N_29213);
or UO_3359 (O_3359,N_26974,N_28965);
xnor UO_3360 (O_3360,N_28676,N_25971);
nand UO_3361 (O_3361,N_27781,N_25884);
nand UO_3362 (O_3362,N_28461,N_25320);
and UO_3363 (O_3363,N_26812,N_28487);
or UO_3364 (O_3364,N_25767,N_27686);
xnor UO_3365 (O_3365,N_29389,N_28383);
nand UO_3366 (O_3366,N_25434,N_29478);
or UO_3367 (O_3367,N_26456,N_29808);
nand UO_3368 (O_3368,N_25648,N_28778);
or UO_3369 (O_3369,N_29995,N_25553);
or UO_3370 (O_3370,N_28486,N_27994);
nand UO_3371 (O_3371,N_26650,N_29752);
and UO_3372 (O_3372,N_28098,N_25505);
xor UO_3373 (O_3373,N_26806,N_27216);
xor UO_3374 (O_3374,N_28303,N_28666);
nor UO_3375 (O_3375,N_25960,N_25543);
nand UO_3376 (O_3376,N_25928,N_27541);
and UO_3377 (O_3377,N_25239,N_29893);
nand UO_3378 (O_3378,N_27646,N_25881);
or UO_3379 (O_3379,N_29335,N_29448);
nor UO_3380 (O_3380,N_25227,N_29376);
or UO_3381 (O_3381,N_25049,N_29596);
nand UO_3382 (O_3382,N_29572,N_26158);
nor UO_3383 (O_3383,N_25208,N_25896);
nand UO_3384 (O_3384,N_28008,N_26123);
nand UO_3385 (O_3385,N_28393,N_28595);
nand UO_3386 (O_3386,N_29253,N_29091);
and UO_3387 (O_3387,N_28568,N_25163);
and UO_3388 (O_3388,N_27206,N_29787);
and UO_3389 (O_3389,N_28578,N_28539);
and UO_3390 (O_3390,N_27981,N_29165);
xor UO_3391 (O_3391,N_29327,N_27046);
xor UO_3392 (O_3392,N_26967,N_29155);
nand UO_3393 (O_3393,N_26663,N_25632);
or UO_3394 (O_3394,N_25769,N_29939);
and UO_3395 (O_3395,N_29513,N_29413);
and UO_3396 (O_3396,N_25293,N_28673);
nand UO_3397 (O_3397,N_26348,N_28360);
and UO_3398 (O_3398,N_26397,N_29651);
xnor UO_3399 (O_3399,N_25554,N_25572);
nand UO_3400 (O_3400,N_25672,N_26855);
or UO_3401 (O_3401,N_26366,N_29885);
and UO_3402 (O_3402,N_25519,N_29952);
xnor UO_3403 (O_3403,N_29508,N_25948);
and UO_3404 (O_3404,N_25779,N_29349);
nor UO_3405 (O_3405,N_26141,N_25870);
nor UO_3406 (O_3406,N_29571,N_27165);
or UO_3407 (O_3407,N_29370,N_25112);
xor UO_3408 (O_3408,N_28544,N_25619);
nand UO_3409 (O_3409,N_29272,N_26765);
and UO_3410 (O_3410,N_28736,N_28953);
xnor UO_3411 (O_3411,N_26636,N_29827);
xnor UO_3412 (O_3412,N_26330,N_29676);
and UO_3413 (O_3413,N_26555,N_29062);
nor UO_3414 (O_3414,N_28788,N_27112);
xor UO_3415 (O_3415,N_25962,N_28046);
nand UO_3416 (O_3416,N_28688,N_29722);
nand UO_3417 (O_3417,N_27972,N_25550);
nor UO_3418 (O_3418,N_27004,N_28842);
and UO_3419 (O_3419,N_27226,N_25504);
and UO_3420 (O_3420,N_26533,N_28996);
nand UO_3421 (O_3421,N_26253,N_26630);
xor UO_3422 (O_3422,N_25923,N_29424);
and UO_3423 (O_3423,N_27024,N_29069);
nand UO_3424 (O_3424,N_26231,N_25427);
or UO_3425 (O_3425,N_29281,N_29580);
nand UO_3426 (O_3426,N_26335,N_29719);
and UO_3427 (O_3427,N_27485,N_25725);
nand UO_3428 (O_3428,N_26445,N_29827);
xnor UO_3429 (O_3429,N_25910,N_26784);
nand UO_3430 (O_3430,N_26096,N_26327);
and UO_3431 (O_3431,N_29747,N_27968);
or UO_3432 (O_3432,N_29853,N_27422);
nand UO_3433 (O_3433,N_29487,N_26397);
nand UO_3434 (O_3434,N_26052,N_25798);
and UO_3435 (O_3435,N_27020,N_29259);
or UO_3436 (O_3436,N_26284,N_27568);
nor UO_3437 (O_3437,N_27606,N_25335);
or UO_3438 (O_3438,N_26613,N_26739);
xnor UO_3439 (O_3439,N_26381,N_25752);
and UO_3440 (O_3440,N_25057,N_27686);
nor UO_3441 (O_3441,N_25889,N_28897);
or UO_3442 (O_3442,N_28827,N_29024);
nor UO_3443 (O_3443,N_25969,N_29382);
nand UO_3444 (O_3444,N_28099,N_26863);
nand UO_3445 (O_3445,N_26283,N_26590);
nand UO_3446 (O_3446,N_28211,N_29750);
xnor UO_3447 (O_3447,N_25446,N_26022);
nand UO_3448 (O_3448,N_28463,N_27815);
nor UO_3449 (O_3449,N_25354,N_26131);
xnor UO_3450 (O_3450,N_26329,N_27335);
nand UO_3451 (O_3451,N_29627,N_25976);
xnor UO_3452 (O_3452,N_27151,N_25946);
nand UO_3453 (O_3453,N_25867,N_25599);
and UO_3454 (O_3454,N_27781,N_27072);
or UO_3455 (O_3455,N_25132,N_29453);
nand UO_3456 (O_3456,N_25448,N_26130);
nand UO_3457 (O_3457,N_28784,N_26446);
nand UO_3458 (O_3458,N_26268,N_25973);
xor UO_3459 (O_3459,N_27688,N_26986);
and UO_3460 (O_3460,N_27673,N_26959);
nand UO_3461 (O_3461,N_29011,N_29072);
nor UO_3462 (O_3462,N_27168,N_29269);
xnor UO_3463 (O_3463,N_29483,N_26934);
nand UO_3464 (O_3464,N_27135,N_27409);
nor UO_3465 (O_3465,N_28907,N_29257);
xor UO_3466 (O_3466,N_29992,N_26843);
nand UO_3467 (O_3467,N_26126,N_25318);
and UO_3468 (O_3468,N_29541,N_25857);
and UO_3469 (O_3469,N_28891,N_29991);
xor UO_3470 (O_3470,N_29673,N_27875);
nor UO_3471 (O_3471,N_26490,N_29026);
nand UO_3472 (O_3472,N_28821,N_26432);
or UO_3473 (O_3473,N_27417,N_27404);
xnor UO_3474 (O_3474,N_26551,N_26394);
and UO_3475 (O_3475,N_29976,N_28153);
xor UO_3476 (O_3476,N_26516,N_28251);
nand UO_3477 (O_3477,N_26497,N_26298);
nor UO_3478 (O_3478,N_29787,N_26910);
nand UO_3479 (O_3479,N_27552,N_28625);
nand UO_3480 (O_3480,N_26446,N_29391);
nor UO_3481 (O_3481,N_27762,N_26455);
or UO_3482 (O_3482,N_29077,N_26972);
nor UO_3483 (O_3483,N_25111,N_26695);
nand UO_3484 (O_3484,N_29661,N_26716);
nand UO_3485 (O_3485,N_28839,N_27393);
nor UO_3486 (O_3486,N_28929,N_26818);
and UO_3487 (O_3487,N_29335,N_25947);
and UO_3488 (O_3488,N_26965,N_25093);
nand UO_3489 (O_3489,N_29017,N_28143);
nand UO_3490 (O_3490,N_28326,N_29585);
nand UO_3491 (O_3491,N_28646,N_28832);
and UO_3492 (O_3492,N_29713,N_28584);
nand UO_3493 (O_3493,N_27644,N_26129);
nand UO_3494 (O_3494,N_27688,N_28258);
nor UO_3495 (O_3495,N_26685,N_28377);
nand UO_3496 (O_3496,N_27016,N_29263);
or UO_3497 (O_3497,N_27527,N_27755);
nor UO_3498 (O_3498,N_29378,N_26267);
or UO_3499 (O_3499,N_26856,N_28756);
endmodule